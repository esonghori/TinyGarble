
module hamming ( x, y, o );
  input [1023:0] x;
  input [1023:0] y;
  output [10:0] o;
  wire   n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442,
         n24443, n24444, n24445, n24446, n24447, n24448, n24449, n24450,
         n24451, n24452, n24453, n24454, n24455, n24456, n24457, n24458,
         n24459, n24460, n24461, n24462, n24463, n24464, n24465, n24466,
         n24467, n24468, n24469, n24470, n24471, n24472, n24473, n24474,
         n24475, n24476, n24477, n24478, n24479, n24480, n24481, n24482,
         n24483, n24484, n24485, n24486, n24487, n24488, n24489, n24490,
         n24491, n24492, n24493, n24494, n24495, n24496, n24497, n24498,
         n24499, n24500, n24501, n24502, n24503, n24504, n24505, n24506,
         n24507, n24508, n24509, n24510, n24511, n24512, n24513, n24514,
         n24515, n24516, n24517, n24518, n24519, n24520, n24521, n24522,
         n24523, n24524, n24525, n24526, n24527, n24528, n24529, n24530,
         n24531, n24532, n24533, n24534, n24535, n24536, n24537, n24538,
         n24539, n24540, n24541, n24542, n24543, n24544, n24545, n24546,
         n24547, n24548, n24549, n24550, n24551, n24552, n24553, n24554,
         n24555, n24556, n24557, n24558, n24559, n24560, n24561, n24562,
         n24563, n24564, n24565, n24566, n24567, n24568, n24569, n24570,
         n24571, n24572, n24573, n24574, n24575, n24576, n24577, n24578,
         n24579, n24580, n24581, n24582, n24583, n24584, n24585, n24586,
         n24587, n24588, n24589, n24590, n24591, n24592, n24593, n24594,
         n24595, n24596, n24597, n24598, n24599, n24600, n24601, n24602,
         n24603, n24604, n24605, n24606, n24607, n24608, n24609, n24610,
         n24611, n24612, n24613, n24614, n24615, n24616, n24617, n24618,
         n24619, n24620, n24621, n24622, n24623, n24624, n24625, n24626,
         n24627, n24628, n24629, n24630, n24631, n24632, n24633, n24634,
         n24635, n24636, n24637, n24638, n24639, n24640, n24641, n24642,
         n24643, n24644, n24645, n24646, n24647, n24648, n24649, n24650,
         n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658,
         n24659, n24660, n24661, n24662, n24663, n24664, n24665, n24666,
         n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674,
         n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682,
         n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24690,
         n24691, n24692, n24693, n24694, n24695, n24696, n24697, n24698,
         n24699, n24700, n24701, n24702, n24703, n24704, n24705, n24706,
         n24707, n24708, n24709, n24710, n24711, n24712, n24713, n24714,
         n24715, n24716, n24717, n24718, n24719, n24720, n24721, n24722,
         n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730,
         n24731, n24732, n24733, n24734, n24735, n24736, n24737, n24738,
         n24739, n24740, n24741, n24742, n24743, n24744, n24745, n24746,
         n24747, n24748, n24749, n24750, n24751, n24752, n24753, n24754,
         n24755, n24756, n24757, n24758, n24759, n24760, n24761, n24762,
         n24763, n24764, n24765, n24766, n24767, n24768, n24769, n24770,
         n24771, n24772, n24773, n24774, n24775, n24776, n24777, n24778,
         n24779, n24780, n24781, n24782, n24783, n24784, n24785, n24786,
         n24787, n24788, n24789, n24790, n24791, n24792, n24793, n24794,
         n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802,
         n24803, n24804, n24805, n24806, n24807, n24808, n24809, n24810,
         n24811, n24812, n24813, n24814, n24815, n24816, n24817, n24818,
         n24819, n24820, n24821, n24822, n24823, n24824, n24825, n24826,
         n24827, n24828, n24829, n24830, n24831, n24832, n24833, n24834,
         n24835, n24836, n24837, n24838, n24839, n24840, n24841, n24842,
         n24843, n24844, n24845, n24846, n24847, n24848, n24849, n24850,
         n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858,
         n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866,
         n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874,
         n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882,
         n24883, n24884, n24885, n24886, n24887, n24888, n24889, n24890,
         n24891, n24892, n24893, n24894, n24895, n24896, n24897, n24898,
         n24899, n24900, n24901, n24902, n24903, n24904, n24905, n24906,
         n24907, n24908, n24909, n24910, n24911, n24912, n24913, n24914,
         n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922,
         n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930,
         n24931, n24932, n24933, n24934, n24935, n24936, n24937, n24938,
         n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24946,
         n24947, n24948, n24949, n24950, n24951, n24952, n24953, n24954,
         n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962,
         n24963, n24964, n24965, n24966, n24967, n24968, n24969, n24970,
         n24971, n24972, n24973, n24974, n24975, n24976, n24977, n24978,
         n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986,
         n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994,
         n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002,
         n25003, n25004, n25005, n25006, n25007, n25008, n25009, n25010,
         n25011, n25012, n25013, n25014, n25015, n25016, n25017, n25018,
         n25019, n25020, n25021, n25022, n25023, n25024, n25025, n25026,
         n25027, n25028, n25029, n25030, n25031, n25032, n25033, n25034,
         n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25042,
         n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050,
         n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058,
         n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066,
         n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074,
         n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082,
         n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090,
         n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098,
         n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106,
         n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114,
         n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122,
         n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130,
         n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138,
         n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146,
         n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154,
         n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162,
         n25163, n25164, n25165, n25166, n25167, n25168, n25169, n25170,
         n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25178,
         n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186,
         n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194,
         n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202,
         n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210,
         n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218,
         n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226,
         n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234,
         n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242,
         n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250,
         n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258,
         n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266,
         n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274,
         n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282,
         n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290,
         n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298,
         n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306,
         n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314,
         n25315, n25316, n25317, n25318, n25319, n25320, n25321, n25322,
         n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330,
         n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338,
         n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346,
         n25347, n25348, n25349, n25350, n25351, n25352, n25353, n25354,
         n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362,
         n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370,
         n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378,
         n25379, n25380, n25381, n25382, n25383, n25384, n25385, n25386,
         n25387, n25388, n25389, n25390, n25391, n25392, n25393, n25394,
         n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402,
         n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410,
         n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418,
         n25419, n25420, n25421, n25422, n25423, n25424, n25425, n25426,
         n25427, n25428, n25429, n25430, n25431, n25432, n25433, n25434,
         n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442,
         n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450,
         n25451, n25452, n25453, n25454, n25455, n25456, n25457, n25458,
         n25459, n25460, n25461, n25462, n25463, n25464, n25465, n25466,
         n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474,
         n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482,
         n25483, n25484, n25485, n25486, n25487, n25488, n25489, n25490,
         n25491, n25492, n25493, n25494, n25495, n25496, n25497, n25498,
         n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506,
         n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514,
         n25515, n25516, n25517, n25518, n25519, n25520, n25521, n25522,
         n25523, n25524, n25525, n25526, n25527, n25528, n25529, n25530,
         n25531, n25532, n25533, n25534, n25535, n25536, n25537, n25538,
         n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546,
         n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554,
         n25555, n25556, n25557, n25558, n25559, n25560, n25561, n25562,
         n25563, n25564, n25565, n25566, n25567, n25568, n25569, n25570,
         n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578,
         n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586,
         n25587, n25588, n25589, n25590, n25591, n25592, n25593, n25594,
         n25595, n25596, n25597, n25598, n25599, n25600, n25601, n25602,
         n25603, n25604, n25605, n25606, n25607, n25608, n25609, n25610,
         n25611, n25612, n25613, n25614, n25615, n25616, n25617, n25618,
         n25619, n25620, n25621, n25622, n25623, n25624, n25625, n25626,
         n25627, n25628, n25629, n25630, n25631, n25632, n25633, n25634,
         n25635, n25636, n25637, n25638, n25639, n25640, n25641, n25642,
         n25643, n25644, n25645, n25646, n25647, n25648, n25649, n25650,
         n25651, n25652, n25653, n25654, n25655, n25656, n25657, n25658,
         n25659, n25660, n25661, n25662, n25663, n25664, n25665, n25666,
         n25667, n25668, n25669, n25670, n25671, n25672, n25673, n25674,
         n25675, n25676, n25677, n25678, n25679, n25680, n25681, n25682,
         n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690,
         n25691, n25692, n25693, n25694, n25695, n25696, n25697, n25698,
         n25699, n25700, n25701, n25702, n25703, n25704, n25705, n25706,
         n25707, n25708, n25709, n25710, n25711, n25712, n25713, n25714,
         n25715, n25716, n25717, n25718, n25719, n25720, n25721, n25722,
         n25723, n25724, n25725, n25726, n25727, n25728, n25729, n25730,
         n25731, n25732, n25733, n25734, n25735, n25736, n25737, n25738,
         n25739, n25740, n25741, n25742, n25743, n25744, n25745, n25746,
         n25747, n25748, n25749, n25750, n25751, n25752, n25753, n25754,
         n25755, n25756, n25757, n25758, n25759, n25760, n25761, n25762,
         n25763, n25764, n25765, n25766, n25767, n25768, n25769, n25770,
         n25771, n25772, n25773, n25774, n25775, n25776, n25777, n25778,
         n25779, n25780, n25781, n25782, n25783, n25784, n25785, n25786,
         n25787, n25788, n25789, n25790, n25791, n25792, n25793, n25794,
         n25795, n25796, n25797, n25798, n25799, n25800, n25801, n25802,
         n25803, n25804, n25805, n25806, n25807, n25808, n25809, n25810,
         n25811, n25812, n25813, n25814, n25815, n25816, n25817, n25818,
         n25819, n25820, n25821, n25822, n25823, n25824, n25825, n25826,
         n25827, n25828, n25829, n25830, n25831, n25832, n25833, n25834,
         n25835, n25836, n25837, n25838, n25839, n25840, n25841, n25842,
         n25843, n25844, n25845, n25846, n25847, n25848, n25849, n25850,
         n25851, n25852, n25853, n25854, n25855, n25856, n25857, n25858,
         n25859, n25860, n25861, n25862, n25863, n25864, n25865, n25866,
         n25867, n25868, n25869, n25870, n25871, n25872, n25873, n25874,
         n25875, n25876, n25877, n25878, n25879, n25880, n25881, n25882,
         n25883, n25884, n25885, n25886, n25887, n25888, n25889, n25890,
         n25891, n25892, n25893, n25894, n25895, n25896, n25897, n25898,
         n25899, n25900, n25901, n25902, n25903, n25904, n25905, n25906,
         n25907, n25908, n25909, n25910, n25911, n25912, n25913, n25914,
         n25915, n25916, n25917, n25918, n25919, n25920, n25921, n25922,
         n25923, n25924, n25925, n25926, n25927, n25928, n25929, n25930,
         n25931, n25932, n25933, n25934, n25935, n25936, n25937, n25938,
         n25939, n25940, n25941, n25942, n25943, n25944, n25945, n25946,
         n25947, n25948, n25949, n25950, n25951, n25952, n25953, n25954,
         n25955, n25956, n25957, n25958, n25959, n25960, n25961, n25962,
         n25963, n25964, n25965, n25966, n25967, n25968, n25969, n25970,
         n25971, n25972, n25973, n25974, n25975, n25976, n25977, n25978,
         n25979, n25980, n25981, n25982, n25983, n25984, n25985, n25986,
         n25987, n25988, n25989, n25990, n25991, n25992, n25993, n25994,
         n25995, n25996, n25997, n25998, n25999, n26000, n26001, n26002,
         n26003, n26004, n26005, n26006, n26007, n26008, n26009, n26010,
         n26011, n26012, n26013, n26014, n26015, n26016, n26017, n26018,
         n26019, n26020, n26021, n26022, n26023, n26024, n26025, n26026,
         n26027, n26028, n26029, n26030, n26031, n26032, n26033, n26034,
         n26035, n26036, n26037, n26038, n26039, n26040, n26041, n26042,
         n26043, n26044, n26045, n26046, n26047, n26048, n26049, n26050,
         n26051, n26052, n26053, n26054, n26055, n26056, n26057, n26058,
         n26059, n26060, n26061, n26062, n26063, n26064, n26065, n26066,
         n26067, n26068, n26069, n26070, n26071, n26072, n26073, n26074,
         n26075, n26076, n26077, n26078, n26079, n26080, n26081, n26082,
         n26083, n26084, n26085, n26086, n26087, n26088, n26089, n26090,
         n26091, n26092, n26093, n26094, n26095, n26096, n26097, n26098,
         n26099, n26100, n26101, n26102, n26103, n26104, n26105, n26106,
         n26107, n26108, n26109, n26110, n26111, n26112, n26113, n26114,
         n26115, n26116, n26117, n26118, n26119, n26120, n26121, n26122,
         n26123, n26124, n26125, n26126, n26127, n26128, n26129, n26130,
         n26131, n26132, n26133, n26134, n26135, n26136, n26137, n26138,
         n26139, n26140, n26141, n26142, n26143, n26144, n26145, n26146,
         n26147, n26148, n26149, n26150, n26151, n26152, n26153, n26154,
         n26155, n26156, n26157, n26158, n26159, n26160, n26161, n26162,
         n26163, n26164, n26165, n26166, n26167, n26168, n26169, n26170,
         n26171, n26172, n26173, n26174, n26175, n26176, n26177, n26178,
         n26179, n26180, n26181, n26182, n26183, n26184, n26185, n26186,
         n26187, n26188, n26189, n26190, n26191, n26192, n26193, n26194,
         n26195, n26196, n26197, n26198, n26199, n26200, n26201, n26202,
         n26203, n26204, n26205, n26206, n26207, n26208, n26209, n26210,
         n26211, n26212, n26213, n26214, n26215, n26216, n26217, n26218,
         n26219, n26220, n26221, n26222, n26223, n26224, n26225, n26226,
         n26227, n26228, n26229, n26230, n26231, n26232, n26233, n26234,
         n26235, n26236, n26237, n26238, n26239, n26240, n26241, n26242,
         n26243, n26244, n26245, n26246, n26247, n26248, n26249, n26250,
         n26251, n26252, n26253, n26254, n26255, n26256, n26257, n26258,
         n26259, n26260, n26261, n26262, n26263, n26264, n26265, n26266,
         n26267, n26268, n26269, n26270, n26271, n26272, n26273, n26274,
         n26275, n26276, n26277, n26278, n26279, n26280, n26281, n26282,
         n26283, n26284, n26285, n26286, n26287, n26288, n26289, n26290,
         n26291, n26292, n26293, n26294, n26295, n26296, n26297, n26298,
         n26299, n26300, n26301, n26302, n26303, n26304, n26305, n26306,
         n26307, n26308, n26309, n26310, n26311, n26312, n26313, n26314,
         n26315, n26316, n26317, n26318, n26319, n26320, n26321, n26322,
         n26323, n26324, n26325, n26326, n26327, n26328, n26329, n26330,
         n26331, n26332, n26333, n26334, n26335, n26336, n26337, n26338,
         n26339, n26340, n26341, n26342, n26343, n26344, n26345, n26346,
         n26347, n26348, n26349, n26350, n26351, n26352, n26353, n26354,
         n26355, n26356, n26357, n26358, n26359, n26360, n26361, n26362,
         n26363, n26364, n26365, n26366, n26367, n26368, n26369, n26370,
         n26371, n26372, n26373, n26374, n26375, n26376, n26377, n26378,
         n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386,
         n26387, n26388, n26389, n26390, n26391, n26392, n26393, n26394,
         n26395, n26396, n26397, n26398, n26399, n26400, n26401, n26402,
         n26403, n26404, n26405, n26406, n26407, n26408, n26409, n26410,
         n26411, n26412, n26413, n26414, n26415, n26416, n26417, n26418,
         n26419, n26420, n26421, n26422, n26423, n26424, n26425, n26426,
         n26427, n26428, n26429, n26430, n26431, n26432, n26433, n26434,
         n26435, n26436, n26437, n26438, n26439, n26440, n26441, n26442,
         n26443, n26444, n26445, n26446, n26447, n26448, n26449, n26450,
         n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458,
         n26459, n26460, n26461, n26462, n26463, n26464, n26465, n26466,
         n26467, n26468, n26469, n26470, n26471, n26472, n26473, n26474,
         n26475, n26476, n26477, n26478, n26479, n26480, n26481, n26482,
         n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490,
         n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498,
         n26499, n26500, n26501, n26502, n26503, n26504, n26505, n26506,
         n26507, n26508, n26509, n26510, n26511, n26512, n26513, n26514,
         n26515, n26516, n26517, n26518, n26519, n26520, n26521, n26522,
         n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530,
         n26531, n26532, n26533, n26534, n26535, n26536, n26537, n26538,
         n26539, n26540, n26541, n26542, n26543, n26544, n26545, n26546,
         n26547, n26548, n26549, n26550, n26551, n26552, n26553, n26554,
         n26555, n26556, n26557, n26558, n26559, n26560, n26561, n26562,
         n26563, n26564, n26565, n26566, n26567, n26568, n26569, n26570,
         n26571, n26572, n26573, n26574, n26575, n26576, n26577, n26578,
         n26579, n26580, n26581, n26582, n26583, n26584, n26585, n26586,
         n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594,
         n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602,
         n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610,
         n26611, n26612, n26613, n26614, n26615, n26616, n26617, n26618,
         n26619, n26620, n26621, n26622, n26623, n26624, n26625, n26626,
         n26627, n26628, n26629, n26630, n26631, n26632, n26633, n26634,
         n26635, n26636, n26637, n26638, n26639, n26640, n26641, n26642,
         n26643, n26644, n26645, n26646, n26647, n26648, n26649, n26650,
         n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658,
         n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666,
         n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674,
         n26675, n26676, n26677, n26678, n26679, n26680, n26681, n26682,
         n26683, n26684, n26685, n26686, n26687, n26688, n26689, n26690,
         n26691, n26692, n26693, n26694, n26695, n26696, n26697, n26698,
         n26699, n26700, n26701, n26702, n26703, n26704, n26705, n26706,
         n26707, n26708, n26709, n26710, n26711, n26712, n26713, n26714,
         n26715, n26716, n26717, n26718, n26719, n26720, n26721, n26722,
         n26723, n26724, n26725, n26726, n26727, n26728, n26729, n26730,
         n26731, n26732, n26733, n26734, n26735, n26736, n26737, n26738,
         n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746,
         n26747, n26748, n26749, n26750, n26751, n26752, n26753, n26754,
         n26755, n26756, n26757, n26758, n26759, n26760, n26761, n26762,
         n26763, n26764, n26765, n26766, n26767, n26768, n26769, n26770,
         n26771, n26772, n26773, n26774, n26775, n26776, n26777, n26778,
         n26779, n26780, n26781, n26782, n26783, n26784, n26785, n26786,
         n26787, n26788, n26789, n26790, n26791, n26792, n26793, n26794,
         n26795, n26796, n26797, n26798, n26799, n26800, n26801, n26802,
         n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810,
         n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818,
         n26819, n26820, n26821, n26822, n26823, n26824, n26825, n26826,
         n26827, n26828, n26829, n26830, n26831, n26832, n26833, n26834,
         n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842,
         n26843, n26844, n26845, n26846, n26847, n26848, n26849, n26850,
         n26851, n26852, n26853, n26854, n26855, n26856, n26857, n26858,
         n26859, n26860, n26861, n26862, n26863, n26864, n26865, n26866,
         n26867, n26868, n26869, n26870, n26871, n26872, n26873, n26874,
         n26875, n26876, n26877, n26878, n26879, n26880, n26881, n26882,
         n26883, n26884, n26885, n26886, n26887, n26888, n26889, n26890,
         n26891, n26892, n26893, n26894, n26895, n26896, n26897, n26898,
         n26899, n26900, n26901, n26902, n26903, n26904, n26905, n26906,
         n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914,
         n26915, n26916, n26917, n26918, n26919, n26920, n26921, n26922,
         n26923, n26924, n26925, n26926, n26927, n26928, n26929, n26930,
         n26931, n26932, n26933, n26934, n26935, n26936, n26937, n26938,
         n26939, n26940, n26941, n26942, n26943, n26944, n26945, n26946,
         n26947, n26948, n26949, n26950, n26951, n26952, n26953, n26954,
         n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962,
         n26963, n26964, n26965, n26966, n26967, n26968, n26969, n26970,
         n26971, n26972, n26973, n26974, n26975, n26976, n26977, n26978,
         n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986,
         n26987, n26988, n26989, n26990, n26991, n26992, n26993, n26994,
         n26995, n26996, n26997, n26998, n26999, n27000, n27001, n27002,
         n27003, n27004, n27005, n27006, n27007, n27008, n27009, n27010,
         n27011, n27012, n27013, n27014, n27015, n27016, n27017, n27018,
         n27019, n27020, n27021, n27022, n27023, n27024, n27025, n27026,
         n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034,
         n27035, n27036, n27037, n27038, n27039, n27040, n27041, n27042,
         n27043, n27044, n27045, n27046, n27047, n27048, n27049, n27050,
         n27051, n27052, n27053, n27054, n27055, n27056, n27057, n27058,
         n27059, n27060, n27061, n27062, n27063, n27064, n27065, n27066,
         n27067, n27068, n27069, n27070, n27071, n27072, n27073, n27074,
         n27075, n27076, n27077, n27078, n27079, n27080, n27081, n27082,
         n27083, n27084, n27085, n27086, n27087, n27088, n27089, n27090,
         n27091, n27092, n27093, n27094, n27095, n27096, n27097, n27098,
         n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27106,
         n27107, n27108, n27109, n27110, n27111, n27112, n27113, n27114,
         n27115, n27116, n27117, n27118, n27119, n27120, n27121, n27122,
         n27123, n27124, n27125, n27126, n27127, n27128, n27129, n27130,
         n27131, n27132, n27133, n27134, n27135, n27136, n27137, n27138,
         n27139, n27140, n27141, n27142, n27143, n27144, n27145, n27146,
         n27147, n27148, n27149, n27150, n27151, n27152, n27153, n27154,
         n27155, n27156, n27157, n27158, n27159, n27160, n27161, n27162,
         n27163, n27164, n27165, n27166, n27167, n27168, n27169, n27170,
         n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178,
         n27179, n27180, n27181, n27182, n27183, n27184, n27185, n27186,
         n27187, n27188, n27189, n27190, n27191, n27192, n27193, n27194,
         n27195, n27196, n27197, n27198, n27199, n27200, n27201, n27202,
         n27203, n27204, n27205, n27206, n27207, n27208, n27209, n27210,
         n27211, n27212, n27213, n27214, n27215, n27216, n27217, n27218,
         n27219, n27220, n27221, n27222, n27223, n27224, n27225, n27226,
         n27227, n27228, n27229, n27230, n27231, n27232, n27233, n27234,
         n27235, n27236, n27237, n27238, n27239, n27240, n27241, n27242,
         n27243, n27244, n27245, n27246, n27247, n27248, n27249, n27250,
         n27251, n27252, n27253, n27254, n27255, n27256, n27257, n27258,
         n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27266,
         n27267, n27268, n27269, n27270, n27271, n27272, n27273, n27274,
         n27275, n27276, n27277, n27278, n27279, n27280, n27281, n27282,
         n27283, n27284, n27285, n27286, n27287, n27288, n27289, n27290,
         n27291, n27292, n27293, n27294, n27295, n27296, n27297, n27298,
         n27299, n27300, n27301, n27302, n27303, n27304, n27305, n27306,
         n27307, n27308, n27309, n27310, n27311, n27312, n27313, n27314,
         n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27322,
         n27323, n27324, n27325, n27326, n27327, n27328, n27329, n27330,
         n27331, n27332, n27333, n27334, n27335, n27336, n27337, n27338,
         n27339, n27340, n27341, n27342, n27343, n27344, n27345, n27346,
         n27347, n27348, n27349, n27350, n27351, n27352, n27353, n27354,
         n27355, n27356, n27357, n27358, n27359, n27360, n27361, n27362,
         n27363, n27364, n27365, n27366, n27367, n27368, n27369, n27370,
         n27371, n27372, n27373, n27374, n27375, n27376, n27377, n27378,
         n27379, n27380, n27381, n27382, n27383, n27384, n27385, n27386,
         n27387, n27388, n27389, n27390, n27391, n27392, n27393, n27394,
         n27395, n27396, n27397, n27398, n27399, n27400, n27401, n27402,
         n27403, n27404, n27405, n27406, n27407, n27408, n27409, n27410,
         n27411, n27412, n27413, n27414, n27415, n27416, n27417, n27418,
         n27419, n27420, n27421, n27422, n27423, n27424, n27425, n27426,
         n27427, n27428, n27429, n27430, n27431, n27432, n27433, n27434,
         n27435, n27436, n27437, n27438, n27439, n27440, n27441, n27442,
         n27443, n27444, n27445, n27446, n27447, n27448, n27449, n27450,
         n27451, n27452, n27453, n27454, n27455, n27456, n27457, n27458,
         n27459, n27460, n27461, n27462, n27463, n27464, n27465, n27466,
         n27467, n27468, n27469, n27470, n27471, n27472, n27473, n27474,
         n27475, n27476, n27477, n27478, n27479, n27480, n27481, n27482,
         n27483, n27484, n27485, n27486, n27487, n27488, n27489, n27490,
         n27491, n27492, n27493, n27494, n27495, n27496, n27497, n27498,
         n27499, n27500, n27501, n27502, n27503, n27504, n27505, n27506,
         n27507, n27508, n27509, n27510, n27511, n27512, n27513, n27514,
         n27515, n27516, n27517, n27518, n27519, n27520, n27521, n27522,
         n27523, n27524, n27525, n27526, n27527, n27528, n27529, n27530,
         n27531, n27532, n27533, n27534, n27535, n27536, n27537, n27538,
         n27539, n27540, n27541, n27542, n27543, n27544, n27545, n27546,
         n27547, n27548, n27549, n27550, n27551, n27552, n27553, n27554,
         n27555, n27556, n27557, n27558, n27559, n27560, n27561, n27562,
         n27563, n27564, n27565, n27566, n27567, n27568, n27569, n27570,
         n27571, n27572, n27573, n27574, n27575, n27576, n27577, n27578,
         n27579, n27580, n27581, n27582, n27583, n27584, n27585, n27586,
         n27587, n27588, n27589, n27590, n27591, n27592, n27593, n27594,
         n27595, n27596, n27597, n27598, n27599, n27600, n27601, n27602,
         n27603, n27604, n27605, n27606, n27607, n27608, n27609, n27610,
         n27611, n27612, n27613, n27614, n27615, n27616, n27617, n27618,
         n27619, n27620, n27621, n27622, n27623, n27624, n27625, n27626,
         n27627, n27628, n27629, n27630, n27631, n27632, n27633, n27634,
         n27635, n27636, n27637, n27638, n27639, n27640, n27641, n27642,
         n27643, n27644, n27645, n27646, n27647, n27648, n27649, n27650,
         n27651, n27652, n27653, n27654, n27655, n27656, n27657, n27658,
         n27659, n27660, n27661, n27662, n27663, n27664, n27665, n27666,
         n27667, n27668, n27669, n27670, n27671, n27672, n27673, n27674,
         n27675, n27676, n27677, n27678, n27679, n27680, n27681, n27682,
         n27683, n27684, n27685, n27686, n27687, n27688, n27689, n27690,
         n27691, n27692, n27693, n27694, n27695, n27696, n27697, n27698,
         n27699, n27700, n27701, n27702, n27703, n27704, n27705, n27706,
         n27707, n27708, n27709, n27710, n27711, n27712, n27713, n27714,
         n27715, n27716, n27717, n27718, n27719, n27720, n27721, n27722,
         n27723, n27724, n27725, n27726, n27727, n27728, n27729, n27730,
         n27731, n27732, n27733, n27734, n27735, n27736, n27737, n27738,
         n27739, n27740, n27741, n27742, n27743, n27744, n27745, n27746,
         n27747, n27748, n27749, n27750, n27751, n27752, n27753, n27754,
         n27755, n27756, n27757, n27758, n27759, n27760, n27761, n27762,
         n27763, n27764, n27765, n27766, n27767, n27768, n27769, n27770,
         n27771, n27772, n27773, n27774, n27775, n27776, n27777, n27778,
         n27779, n27780, n27781, n27782, n27783, n27784, n27785, n27786,
         n27787, n27788, n27789, n27790, n27791, n27792, n27793, n27794,
         n27795, n27796, n27797, n27798, n27799, n27800, n27801, n27802,
         n27803, n27804, n27805, n27806, n27807, n27808, n27809, n27810,
         n27811, n27812, n27813, n27814, n27815, n27816, n27817, n27818,
         n27819, n27820, n27821, n27822, n27823, n27824, n27825, n27826,
         n27827, n27828, n27829, n27830, n27831, n27832, n27833, n27834,
         n27835, n27836, n27837, n27838, n27839, n27840, n27841, n27842,
         n27843, n27844, n27845, n27846, n27847, n27848, n27849, n27850,
         n27851, n27852, n27853, n27854, n27855, n27856, n27857, n27858,
         n27859, n27860, n27861, n27862, n27863, n27864, n27865, n27866,
         n27867, n27868, n27869, n27870, n27871, n27872, n27873, n27874,
         n27875, n27876, n27877, n27878, n27879, n27880, n27881, n27882,
         n27883, n27884, n27885, n27886, n27887, n27888, n27889, n27890,
         n27891, n27892, n27893, n27894, n27895, n27896, n27897, n27898,
         n27899, n27900, n27901, n27902, n27903, n27904, n27905, n27906,
         n27907, n27908, n27909, n27910, n27911, n27912, n27913, n27914,
         n27915, n27916, n27917, n27918, n27919, n27920, n27921, n27922,
         n27923, n27924, n27925, n27926, n27927, n27928, n27929, n27930,
         n27931, n27932, n27933, n27934, n27935, n27936, n27937, n27938,
         n27939, n27940, n27941, n27942, n27943, n27944, n27945, n27946,
         n27947, n27948, n27949, n27950, n27951, n27952, n27953, n27954,
         n27955, n27956, n27957, n27958, n27959, n27960, n27961, n27962,
         n27963, n27964, n27965, n27966, n27967, n27968, n27969, n27970,
         n27971, n27972, n27973, n27974, n27975, n27976, n27977, n27978,
         n27979, n27980, n27981, n27982, n27983, n27984, n27985, n27986,
         n27987, n27988, n27989, n27990, n27991, n27992, n27993, n27994,
         n27995, n27996, n27997, n27998, n27999, n28000, n28001, n28002,
         n28003, n28004, n28005, n28006, n28007, n28008, n28009, n28010,
         n28011, n28012, n28013, n28014, n28015, n28016, n28017, n28018,
         n28019, n28020, n28021, n28022, n28023, n28024, n28025, n28026,
         n28027, n28028, n28029, n28030, n28031, n28032, n28033, n28034,
         n28035, n28036, n28037, n28038, n28039, n28040, n28041, n28042,
         n28043, n28044, n28045, n28046, n28047, n28048, n28049, n28050,
         n28051, n28052, n28053, n28054, n28055, n28056, n28057, n28058,
         n28059, n28060, n28061, n28062, n28063, n28064, n28065, n28066,
         n28067, n28068, n28069, n28070, n28071, n28072, n28073, n28074,
         n28075, n28076, n28077, n28078, n28079, n28080, n28081, n28082,
         n28083, n28084, n28085, n28086, n28087, n28088, n28089, n28090,
         n28091, n28092, n28093, n28094, n28095, n28096, n28097, n28098,
         n28099, n28100, n28101, n28102, n28103, n28104, n28105, n28106,
         n28107, n28108, n28109, n28110, n28111, n28112, n28113, n28114,
         n28115, n28116, n28117, n28118, n28119, n28120, n28121, n28122,
         n28123, n28124, n28125, n28126, n28127, n28128, n28129, n28130,
         n28131, n28132, n28133, n28134, n28135, n28136, n28137, n28138,
         n28139, n28140, n28141, n28142, n28143, n28144, n28145, n28146,
         n28147, n28148, n28149, n28150, n28151, n28152, n28153, n28154,
         n28155, n28156, n28157, n28158, n28159, n28160, n28161, n28162,
         n28163, n28164, n28165, n28166, n28167, n28168, n28169, n28170,
         n28171, n28172, n28173, n28174, n28175, n28176, n28177, n28178,
         n28179, n28180, n28181, n28182, n28183, n28184, n28185, n28186,
         n28187, n28188, n28189, n28190, n28191, n28192, n28193, n28194,
         n28195, n28196, n28197, n28198, n28199, n28200, n28201, n28202,
         n28203, n28204, n28205, n28206, n28207, n28208, n28209, n28210,
         n28211, n28212, n28213, n28214, n28215, n28216, n28217, n28218,
         n28219, n28220, n28221, n28222, n28223, n28224, n28225, n28226,
         n28227, n28228, n28229, n28230, n28231, n28232, n28233, n28234,
         n28235, n28236, n28237, n28238, n28239, n28240, n28241, n28242,
         n28243, n28244, n28245, n28246, n28247, n28248, n28249, n28250,
         n28251, n28252, n28253, n28254, n28255, n28256, n28257, n28258,
         n28259, n28260, n28261, n28262, n28263, n28264, n28265, n28266,
         n28267, n28268, n28269, n28270, n28271, n28272, n28273, n28274,
         n28275, n28276, n28277, n28278, n28279, n28280, n28281, n28282,
         n28283, n28284, n28285, n28286, n28287, n28288, n28289, n28290,
         n28291, n28292, n28293, n28294, n28295, n28296, n28297, n28298,
         n28299, n28300, n28301, n28302, n28303, n28304, n28305, n28306,
         n28307, n28308, n28309, n28310, n28311, n28312, n28313, n28314,
         n28315, n28316, n28317, n28318, n28319, n28320, n28321, n28322,
         n28323, n28324, n28325, n28326, n28327, n28328, n28329, n28330,
         n28331, n28332, n28333, n28334, n28335, n28336, n28337, n28338,
         n28339, n28340, n28341, n28342, n28343, n28344, n28345, n28346,
         n28347, n28348, n28349, n28350, n28351, n28352, n28353, n28354,
         n28355, n28356, n28357, n28358, n28359, n28360, n28361, n28362,
         n28363, n28364, n28365, n28366, n28367, n28368, n28369, n28370,
         n28371, n28372, n28373, n28374, n28375, n28376, n28377, n28378,
         n28379, n28380, n28381, n28382, n28383, n28384, n28385, n28386,
         n28387, n28388, n28389, n28390, n28391, n28392, n28393, n28394,
         n28395, n28396, n28397, n28398, n28399, n28400, n28401, n28402,
         n28403, n28404, n28405, n28406, n28407, n28408, n28409, n28410,
         n28411, n28412, n28413, n28414, n28415, n28416, n28417, n28418,
         n28419, n28420, n28421, n28422, n28423, n28424, n28425, n28426,
         n28427, n28428, n28429, n28430, n28431, n28432, n28433, n28434,
         n28435, n28436, n28437, n28438, n28439, n28440, n28441, n28442,
         n28443, n28444, n28445, n28446, n28447, n28448, n28449, n28450,
         n28451, n28452, n28453, n28454, n28455, n28456, n28457, n28458,
         n28459, n28460, n28461, n28462, n28463, n28464, n28465, n28466,
         n28467, n28468, n28469, n28470, n28471, n28472, n28473, n28474,
         n28475, n28476, n28477, n28478, n28479, n28480, n28481, n28482,
         n28483, n28484, n28485, n28486, n28487, n28488, n28489, n28490,
         n28491, n28492, n28493, n28494, n28495, n28496, n28497, n28498,
         n28499, n28500, n28501, n28502, n28503, n28504, n28505, n28506,
         n28507, n28508, n28509, n28510, n28511, n28512, n28513, n28514,
         n28515, n28516, n28517, n28518, n28519, n28520, n28521, n28522,
         n28523, n28524, n28525, n28526, n28527, n28528, n28529, n28530,
         n28531, n28532, n28533, n28534, n28535, n28536, n28537, n28538,
         n28539, n28540, n28541, n28542, n28543, n28544, n28545, n28546,
         n28547, n28548, n28549, n28550, n28551, n28552, n28553, n28554,
         n28555, n28556, n28557, n28558, n28559, n28560, n28561, n28562,
         n28563, n28564, n28565, n28566, n28567, n28568, n28569, n28570,
         n28571, n28572, n28573, n28574, n28575, n28576, n28577, n28578,
         n28579, n28580, n28581, n28582, n28583, n28584, n28585, n28586,
         n28587, n28588, n28589, n28590, n28591, n28592, n28593, n28594,
         n28595, n28596, n28597, n28598, n28599, n28600, n28601, n28602,
         n28603, n28604, n28605, n28606, n28607, n28608, n28609, n28610,
         n28611, n28612, n28613, n28614, n28615, n28616, n28617, n28618,
         n28619, n28620, n28621, n28622, n28623, n28624, n28625, n28626,
         n28627, n28628, n28629, n28630, n28631, n28632, n28633, n28634,
         n28635, n28636, n28637, n28638, n28639, n28640, n28641, n28642,
         n28643, n28644, n28645, n28646, n28647, n28648, n28649, n28650,
         n28651, n28652, n28653, n28654, n28655, n28656, n28657, n28658,
         n28659, n28660, n28661, n28662, n28663, n28664, n28665, n28666,
         n28667, n28668, n28669, n28670, n28671, n28672, n28673, n28674,
         n28675, n28676, n28677, n28678, n28679, n28680, n28681, n28682,
         n28683, n28684, n28685, n28686, n28687, n28688, n28689, n28690,
         n28691, n28692, n28693, n28694, n28695, n28696, n28697, n28698,
         n28699, n28700, n28701, n28702, n28703, n28704, n28705, n28706,
         n28707, n28708, n28709, n28710, n28711, n28712, n28713, n28714,
         n28715, n28716, n28717, n28718, n28719, n28720, n28721, n28722,
         n28723, n28724, n28725, n28726, n28727, n28728, n28729, n28730,
         n28731, n28732, n28733, n28734, n28735, n28736, n28737, n28738,
         n28739, n28740, n28741, n28742, n28743, n28744, n28745, n28746,
         n28747, n28748, n28749, n28750, n28751, n28752, n28753, n28754,
         n28755, n28756, n28757, n28758, n28759, n28760, n28761, n28762,
         n28763, n28764, n28765, n28766, n28767, n28768, n28769, n28770,
         n28771, n28772, n28773, n28774, n28775, n28776, n28777, n28778,
         n28779, n28780, n28781, n28782, n28783, n28784, n28785, n28786,
         n28787, n28788, n28789, n28790, n28791, n28792, n28793, n28794,
         n28795, n28796, n28797, n28798, n28799, n28800, n28801, n28802,
         n28803, n28804, n28805, n28806, n28807, n28808, n28809, n28810,
         n28811, n28812, n28813, n28814, n28815, n28816, n28817, n28818,
         n28819, n28820, n28821, n28822, n28823, n28824, n28825, n28826,
         n28827, n28828, n28829, n28830, n28831, n28832, n28833, n28834,
         n28835, n28836, n28837, n28838, n28839, n28840, n28841, n28842,
         n28843, n28844, n28845, n28846, n28847, n28848, n28849, n28850,
         n28851, n28852, n28853, n28854, n28855, n28856, n28857, n28858,
         n28859, n28860, n28861, n28862, n28863, n28864, n28865, n28866,
         n28867, n28868, n28869, n28870, n28871, n28872, n28873, n28874,
         n28875, n28876, n28877, n28878, n28879, n28880, n28881, n28882,
         n28883, n28884, n28885, n28886, n28887, n28888, n28889, n28890,
         n28891, n28892, n28893, n28894, n28895, n28896, n28897, n28898,
         n28899, n28900, n28901, n28902, n28903, n28904, n28905, n28906,
         n28907, n28908, n28909, n28910, n28911, n28912, n28913, n28914,
         n28915, n28916, n28917, n28918, n28919, n28920, n28921, n28922,
         n28923, n28924, n28925, n28926, n28927, n28928, n28929, n28930,
         n28931, n28932, n28933, n28934, n28935, n28936, n28937, n28938,
         n28939, n28940, n28941, n28942, n28943, n28944, n28945, n28946,
         n28947, n28948, n28949, n28950, n28951, n28952, n28953, n28954,
         n28955, n28956, n28957, n28958, n28959, n28960, n28961, n28962,
         n28963, n28964, n28965, n28966, n28967, n28968, n28969, n28970,
         n28971, n28972, n28973, n28974, n28975, n28976, n28977, n28978,
         n28979, n28980, n28981, n28982, n28983, n28984, n28985, n28986,
         n28987, n28988, n28989, n28990, n28991, n28992, n28993, n28994,
         n28995, n28996, n28997, n28998, n28999, n29000, n29001, n29002,
         n29003, n29004, n29005, n29006, n29007, n29008, n29009, n29010,
         n29011, n29012, n29013, n29014, n29015, n29016, n29017, n29018,
         n29019, n29020, n29021, n29022, n29023, n29024, n29025, n29026,
         n29027, n29028, n29029, n29030, n29031, n29032, n29033, n29034,
         n29035, n29036, n29037, n29038, n29039, n29040, n29041, n29042,
         n29043, n29044, n29045, n29046, n29047, n29048, n29049, n29050,
         n29051, n29052, n29053, n29054, n29055, n29056, n29057, n29058,
         n29059, n29060, n29061, n29062, n29063, n29064, n29065, n29066,
         n29067, n29068, n29069, n29070, n29071, n29072, n29073, n29074,
         n29075, n29076, n29077, n29078, n29079, n29080, n29081, n29082,
         n29083, n29084, n29085, n29086, n29087, n29088, n29089, n29090,
         n29091, n29092, n29093, n29094, n29095, n29096, n29097, n29098,
         n29099, n29100, n29101, n29102, n29103, n29104, n29105, n29106,
         n29107, n29108, n29109, n29110, n29111, n29112, n29113, n29114,
         n29115, n29116, n29117, n29118, n29119, n29120, n29121, n29122,
         n29123, n29124, n29125, n29126, n29127, n29128, n29129, n29130,
         n29131, n29132, n29133, n29134, n29135, n29136, n29137, n29138,
         n29139, n29140, n29141, n29142, n29143, n29144, n29145, n29146,
         n29147, n29148, n29149, n29150, n29151, n29152, n29153, n29154,
         n29155, n29156, n29157, n29158, n29159, n29160, n29161, n29162,
         n29163, n29164, n29165, n29166, n29167, n29168, n29169, n29170,
         n29171, n29172, n29173, n29174, n29175, n29176, n29177, n29178,
         n29179, n29180, n29181, n29182, n29183, n29184, n29185, n29186,
         n29187, n29188, n29189, n29190, n29191, n29192, n29193, n29194,
         n29195, n29196, n29197, n29198, n29199, n29200, n29201, n29202,
         n29203, n29204, n29205, n29206, n29207, n29208, n29209, n29210,
         n29211, n29212, n29213, n29214, n29215, n29216, n29217, n29218,
         n29219, n29220, n29221, n29222, n29223, n29224, n29225, n29226,
         n29227, n29228, n29229, n29230, n29231, n29232, n29233, n29234,
         n29235, n29236, n29237, n29238, n29239, n29240, n29241, n29242,
         n29243, n29244, n29245, n29246, n29247, n29248, n29249, n29250,
         n29251, n29252, n29253, n29254, n29255, n29256, n29257, n29258,
         n29259, n29260, n29261, n29262, n29263, n29264, n29265, n29266,
         n29267, n29268, n29269, n29270, n29271, n29272, n29273, n29274,
         n29275, n29276, n29277, n29278, n29279, n29280, n29281, n29282,
         n29283, n29284, n29285, n29286, n29287, n29288, n29289, n29290,
         n29291, n29292, n29293, n29294, n29295, n29296, n29297, n29298,
         n29299, n29300, n29301, n29302, n29303, n29304, n29305, n29306,
         n29307, n29308, n29309, n29310, n29311, n29312, n29313, n29314,
         n29315, n29316, n29317, n29318, n29319, n29320, n29321, n29322,
         n29323, n29324, n29325, n29326, n29327, n29328, n29329, n29330,
         n29331, n29332, n29333, n29334, n29335, n29336, n29337, n29338,
         n29339, n29340, n29341, n29342, n29343, n29344, n29345, n29346,
         n29347, n29348, n29349, n29350, n29351, n29352, n29353, n29354,
         n29355, n29356, n29357, n29358, n29359, n29360, n29361, n29362,
         n29363, n29364, n29365, n29366, n29367, n29368, n29369, n29370,
         n29371, n29372, n29373, n29374, n29375, n29376, n29377, n29378,
         n29379, n29380, n29381, n29382, n29383, n29384, n29385, n29386,
         n29387, n29388, n29389, n29390, n29391, n29392, n29393, n29394,
         n29395, n29396, n29397, n29398, n29399, n29400, n29401, n29402,
         n29403, n29404, n29405, n29406, n29407, n29408, n29409, n29410,
         n29411, n29412, n29413, n29414, n29415, n29416, n29417, n29418,
         n29419, n29420, n29421, n29422, n29423, n29424, n29425, n29426,
         n29427, n29428, n29429, n29430, n29431, n29432, n29433, n29434,
         n29435, n29436, n29437, n29438, n29439, n29440, n29441, n29442,
         n29443, n29444, n29445, n29446, n29447, n29448, n29449, n29450,
         n29451, n29452, n29453, n29454, n29455, n29456, n29457, n29458,
         n29459, n29460, n29461, n29462, n29463, n29464, n29465, n29466,
         n29467, n29468, n29469, n29470, n29471, n29472, n29473, n29474,
         n29475, n29476, n29477, n29478, n29479, n29480, n29481, n29482,
         n29483, n29484, n29485, n29486, n29487, n29488, n29489, n29490,
         n29491, n29492, n29493, n29494, n29495, n29496, n29497, n29498,
         n29499, n29500, n29501, n29502, n29503, n29504, n29505, n29506,
         n29507, n29508, n29509, n29510, n29511, n29512, n29513, n29514,
         n29515, n29516, n29517, n29518, n29519, n29520, n29521, n29522,
         n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530,
         n29531, n29532, n29533, n29534, n29535, n29536, n29537, n29538,
         n29539, n29540, n29541, n29542, n29543, n29544, n29545, n29546,
         n29547, n29548, n29549, n29550, n29551, n29552, n29553, n29554,
         n29555, n29556, n29557, n29558, n29559, n29560, n29561, n29562,
         n29563, n29564, n29565, n29566, n29567, n29568, n29569, n29570,
         n29571, n29572, n29573, n29574, n29575, n29576, n29577, n29578,
         n29579, n29580, n29581, n29582, n29583, n29584, n29585, n29586,
         n29587, n29588, n29589, n29590, n29591, n29592, n29593, n29594,
         n29595, n29596, n29597, n29598, n29599, n29600, n29601, n29602,
         n29603, n29604, n29605, n29606, n29607, n29608, n29609, n29610,
         n29611, n29612, n29613, n29614, n29615, n29616, n29617, n29618,
         n29619, n29620, n29621, n29622, n29623, n29624, n29625, n29626,
         n29627, n29628, n29629, n29630, n29631, n29632, n29633, n29634,
         n29635, n29636, n29637, n29638, n29639, n29640, n29641, n29642,
         n29643, n29644, n29645, n29646, n29647, n29648, n29649, n29650,
         n29651, n29652, n29653, n29654, n29655, n29656, n29657, n29658,
         n29659, n29660, n29661, n29662, n29663, n29664, n29665, n29666,
         n29667, n29668, n29669, n29670, n29671, n29672, n29673, n29674,
         n29675, n29676, n29677, n29678, n29679, n29680, n29681, n29682,
         n29683, n29684, n29685, n29686, n29687, n29688, n29689, n29690,
         n29691, n29692, n29693, n29694, n29695, n29696, n29697, n29698,
         n29699, n29700, n29701, n29702, n29703, n29704, n29705, n29706,
         n29707, n29708, n29709, n29710, n29711, n29712, n29713, n29714,
         n29715, n29716, n29717, n29718, n29719, n29720, n29721, n29722,
         n29723, n29724, n29725, n29726, n29727, n29728, n29729, n29730,
         n29731, n29732, n29733, n29734, n29735, n29736, n29737, n29738,
         n29739, n29740, n29741, n29742, n29743, n29744, n29745, n29746,
         n29747, n29748, n29749, n29750, n29751, n29752, n29753, n29754,
         n29755, n29756, n29757, n29758, n29759, n29760, n29761, n29762,
         n29763, n29764, n29765, n29766, n29767, n29768, n29769, n29770,
         n29771, n29772, n29773, n29774, n29775, n29776, n29777, n29778,
         n29779, n29780, n29781, n29782, n29783, n29784, n29785, n29786,
         n29787, n29788, n29789, n29790, n29791, n29792, n29793, n29794,
         n29795, n29796, n29797, n29798, n29799, n29800, n29801, n29802,
         n29803, n29804, n29805, n29806, n29807, n29808, n29809, n29810,
         n29811, n29812, n29813, n29814, n29815, n29816, n29817, n29818,
         n29819, n29820, n29821, n29822, n29823, n29824, n29825, n29826,
         n29827, n29828, n29829, n29830, n29831, n29832, n29833, n29834,
         n29835, n29836, n29837, n29838, n29839, n29840, n29841, n29842,
         n29843, n29844, n29845, n29846, n29847, n29848, n29849, n29850,
         n29851, n29852, n29853, n29854, n29855, n29856, n29857, n29858,
         n29859, n29860, n29861, n29862, n29863, n29864, n29865, n29866,
         n29867, n29868, n29869, n29870, n29871, n29872, n29873, n29874,
         n29875, n29876, n29877, n29878, n29879, n29880, n29881, n29882,
         n29883, n29884, n29885, n29886, n29887, n29888, n29889, n29890,
         n29891, n29892, n29893, n29894, n29895, n29896, n29897, n29898,
         n29899, n29900, n29901, n29902, n29903, n29904, n29905, n29906,
         n29907, n29908, n29909, n29910, n29911, n29912, n29913, n29914,
         n29915, n29916, n29917, n29918, n29919, n29920, n29921, n29922,
         n29923, n29924, n29925, n29926, n29927, n29928, n29929, n29930,
         n29931, n29932, n29933, n29934, n29935, n29936, n29937, n29938,
         n29939, n29940, n29941, n29942, n29943, n29944, n29945, n29946,
         n29947, n29948, n29949, n29950, n29951, n29952, n29953, n29954,
         n29955, n29956, n29957, n29958, n29959, n29960, n29961, n29962,
         n29963, n29964, n29965, n29966, n29967, n29968, n29969, n29970,
         n29971, n29972, n29973, n29974, n29975, n29976, n29977, n29978,
         n29979, n29980, n29981, n29982, n29983, n29984, n29985, n29986,
         n29987, n29988, n29989, n29990, n29991, n29992, n29993, n29994,
         n29995, n29996, n29997, n29998, n29999, n30000, n30001, n30002,
         n30003, n30004, n30005, n30006, n30007, n30008, n30009, n30010,
         n30011, n30012, n30013, n30014, n30015, n30016, n30017, n30018,
         n30019, n30020, n30021, n30022, n30023, n30024, n30025, n30026,
         n30027, n30028, n30029, n30030, n30031, n30032, n30033, n30034,
         n30035, n30036, n30037, n30038, n30039, n30040, n30041, n30042,
         n30043, n30044, n30045, n30046, n30047, n30048, n30049, n30050,
         n30051, n30052, n30053, n30054, n30055, n30056, n30057, n30058,
         n30059, n30060, n30061, n30062, n30063, n30064, n30065, n30066,
         n30067, n30068, n30069, n30070, n30071, n30072, n30073, n30074,
         n30075, n30076, n30077, n30078, n30079, n30080, n30081, n30082,
         n30083, n30084, n30085, n30086, n30087, n30088, n30089, n30090,
         n30091, n30092, n30093, n30094, n30095, n30096, n30097, n30098,
         n30099, n30100, n30101, n30102, n30103, n30104, n30105, n30106,
         n30107, n30108, n30109, n30110, n30111, n30112, n30113, n30114,
         n30115, n30116, n30117, n30118, n30119, n30120, n30121, n30122,
         n30123, n30124, n30125, n30126, n30127, n30128, n30129, n30130,
         n30131, n30132, n30133, n30134, n30135, n30136, n30137, n30138,
         n30139, n30140, n30141, n30142, n30143, n30144, n30145, n30146,
         n30147, n30148, n30149, n30150, n30151, n30152, n30153, n30154,
         n30155, n30156, n30157, n30158, n30159, n30160, n30161, n30162,
         n30163, n30164, n30165, n30166, n30167, n30168, n30169, n30170,
         n30171, n30172, n30173, n30174, n30175, n30176, n30177, n30178,
         n30179, n30180, n30181, n30182, n30183, n30184, n30185, n30186,
         n30187, n30188, n30189, n30190, n30191, n30192, n30193, n30194,
         n30195, n30196, n30197, n30198, n30199, n30200, n30201, n30202,
         n30203, n30204, n30205, n30206, n30207, n30208, n30209, n30210,
         n30211, n30212, n30213, n30214, n30215, n30216, n30217, n30218,
         n30219, n30220, n30221, n30222, n30223, n30224, n30225, n30226,
         n30227, n30228, n30229, n30230, n30231, n30232, n30233, n30234,
         n30235, n30236, n30237, n30238, n30239, n30240, n30241, n30242,
         n30243, n30244, n30245, n30246, n30247, n30248, n30249, n30250,
         n30251, n30252, n30253, n30254, n30255, n30256, n30257, n30258,
         n30259, n30260, n30261, n30262, n30263, n30264, n30265, n30266,
         n30267, n30268, n30269, n30270, n30271, n30272, n30273, n30274,
         n30275, n30276, n30277, n30278, n30279, n30280, n30281, n30282,
         n30283, n30284, n30285, n30286, n30287, n30288, n30289, n30290,
         n30291, n30292, n30293, n30294, n30295, n30296, n30297, n30298,
         n30299, n30300, n30301, n30302, n30303, n30304, n30305, n30306,
         n30307, n30308, n30309, n30310, n30311, n30312, n30313, n30314,
         n30315, n30316, n30317, n30318, n30319, n30320, n30321, n30322,
         n30323, n30324, n30325, n30326, n30327, n30328, n30329, n30330,
         n30331, n30332, n30333, n30334, n30335, n30336, n30337, n30338,
         n30339, n30340, n30341, n30342, n30343, n30344, n30345, n30346,
         n30347, n30348, n30349, n30350, n30351, n30352, n30353, n30354,
         n30355, n30356, n30357, n30358, n30359, n30360, n30361, n30362,
         n30363, n30364, n30365, n30366, n30367, n30368, n30369, n30370,
         n30371, n30372, n30373, n30374, n30375, n30376, n30377, n30378,
         n30379, n30380, n30381, n30382, n30383, n30384, n30385, n30386,
         n30387, n30388, n30389, n30390, n30391, n30392, n30393, n30394,
         n30395, n30396, n30397, n30398, n30399, n30400, n30401, n30402,
         n30403, n30404, n30405, n30406, n30407, n30408, n30409, n30410,
         n30411, n30412, n30413, n30414, n30415, n30416, n30417, n30418,
         n30419, n30420, n30421, n30422, n30423, n30424, n30425, n30426,
         n30427, n30428, n30429, n30430, n30431, n30432, n30433, n30434,
         n30435, n30436, n30437, n30438, n30439, n30440, n30441, n30442,
         n30443, n30444, n30445, n30446, n30447, n30448, n30449, n30450,
         n30451, n30452, n30453, n30454, n30455, n30456, n30457, n30458,
         n30459, n30460, n30461, n30462, n30463, n30464, n30465, n30466,
         n30467, n30468, n30469, n30470, n30471, n30472, n30473, n30474,
         n30475, n30476, n30477, n30478, n30479, n30480, n30481, n30482,
         n30483, n30484, n30485, n30486, n30487, n30488, n30489, n30490,
         n30491, n30492, n30493, n30494, n30495, n30496, n30497, n30498,
         n30499, n30500, n30501, n30502, n30503, n30504, n30505, n30506,
         n30507, n30508, n30509, n30510, n30511, n30512, n30513, n30514,
         n30515, n30516, n30517, n30518, n30519, n30520, n30521, n30522,
         n30523, n30524, n30525, n30526, n30527, n30528, n30529, n30530,
         n30531, n30532, n30533, n30534, n30535, n30536, n30537, n30538,
         n30539, n30540, n30541, n30542, n30543, n30544, n30545, n30546,
         n30547, n30548, n30549, n30550, n30551, n30552, n30553, n30554,
         n30555, n30556, n30557, n30558, n30559, n30560, n30561, n30562,
         n30563, n30564, n30565, n30566, n30567, n30568, n30569, n30570,
         n30571, n30572, n30573, n30574, n30575, n30576, n30577, n30578,
         n30579, n30580, n30581, n30582, n30583, n30584, n30585, n30586,
         n30587, n30588, n30589, n30590, n30591, n30592, n30593, n30594,
         n30595, n30596, n30597, n30598, n30599, n30600, n30601, n30602,
         n30603, n30604, n30605, n30606, n30607, n30608, n30609, n30610,
         n30611, n30612, n30613, n30614, n30615, n30616, n30617, n30618,
         n30619, n30620, n30621, n30622, n30623, n30624, n30625, n30626,
         n30627, n30628, n30629, n30630, n30631, n30632, n30633, n30634,
         n30635, n30636, n30637, n30638, n30639, n30640, n30641, n30642,
         n30643, n30644, n30645, n30646, n30647, n30648, n30649, n30650,
         n30651, n30652, n30653, n30654, n30655, n30656, n30657, n30658,
         n30659, n30660, n30661, n30662, n30663, n30664, n30665, n30666,
         n30667, n30668, n30669, n30670, n30671, n30672, n30673, n30674,
         n30675, n30676, n30677, n30678, n30679, n30680, n30681, n30682,
         n30683, n30684, n30685, n30686, n30687, n30688, n30689, n30690,
         n30691, n30692, n30693, n30694, n30695, n30696, n30697, n30698,
         n30699, n30700, n30701, n30702, n30703, n30704, n30705, n30706,
         n30707, n30708, n30709, n30710, n30711, n30712, n30713, n30714,
         n30715, n30716, n30717, n30718, n30719, n30720, n30721, n30722,
         n30723, n30724, n30725, n30726, n30727, n30728, n30729, n30730,
         n30731, n30732, n30733, n30734, n30735, n30736, n30737, n30738,
         n30739, n30740, n30741, n30742, n30743, n30744, n30745, n30746,
         n30747, n30748, n30749, n30750, n30751, n30752, n30753, n30754,
         n30755, n30756, n30757, n30758, n30759, n30760, n30761, n30762,
         n30763, n30764, n30765, n30766, n30767, n30768, n30769, n30770,
         n30771, n30772, n30773, n30774, n30775, n30776, n30777, n30778,
         n30779, n30780, n30781, n30782, n30783, n30784, n30785, n30786,
         n30787, n30788, n30789, n30790, n30791, n30792, n30793, n30794,
         n30795, n30796, n30797, n30798, n30799, n30800, n30801, n30802,
         n30803, n30804, n30805, n30806, n30807, n30808, n30809, n30810,
         n30811, n30812, n30813, n30814, n30815, n30816, n30817, n30818,
         n30819, n30820, n30821, n30822, n30823, n30824, n30825, n30826,
         n30827, n30828, n30829, n30830, n30831, n30832, n30833, n30834,
         n30835, n30836, n30837, n30838, n30839, n30840, n30841, n30842,
         n30843, n30844, n30845, n30846, n30847, n30848, n30849, n30850,
         n30851, n30852, n30853, n30854, n30855, n30856, n30857, n30858,
         n30859, n30860, n30861, n30862, n30863, n30864, n30865, n30866,
         n30867, n30868, n30869, n30870, n30871, n30872, n30873, n30874,
         n30875, n30876, n30877, n30878, n30879, n30880, n30881, n30882,
         n30883, n30884, n30885, n30886, n30887, n30888, n30889, n30890,
         n30891, n30892, n30893, n30894, n30895, n30896, n30897, n30898,
         n30899, n30900, n30901, n30902, n30903, n30904, n30905, n30906,
         n30907, n30908, n30909, n30910, n30911, n30912, n30913, n30914,
         n30915, n30916, n30917, n30918, n30919, n30920, n30921, n30922,
         n30923, n30924, n30925, n30926, n30927, n30928, n30929, n30930,
         n30931, n30932, n30933, n30934, n30935, n30936, n30937, n30938,
         n30939, n30940, n30941, n30942, n30943, n30944, n30945, n30946,
         n30947, n30948, n30949, n30950, n30951, n30952, n30953, n30954,
         n30955, n30956, n30957, n30958, n30959, n30960, n30961, n30962,
         n30963, n30964, n30965, n30966, n30967, n30968, n30969, n30970,
         n30971, n30972, n30973, n30974, n30975, n30976, n30977, n30978,
         n30979, n30980, n30981, n30982, n30983, n30984, n30985, n30986,
         n30987, n30988, n30989, n30990, n30991, n30992, n30993, n30994,
         n30995, n30996, n30997, n30998, n30999, n31000, n31001, n31002,
         n31003, n31004, n31005, n31006, n31007, n31008, n31009, n31010,
         n31011, n31012, n31013, n31014, n31015, n31016, n31017, n31018,
         n31019, n31020, n31021, n31022, n31023, n31024, n31025, n31026,
         n31027, n31028, n31029, n31030, n31031, n31032, n31033, n31034,
         n31035, n31036, n31037, n31038, n31039, n31040, n31041, n31042,
         n31043, n31044, n31045, n31046, n31047, n31048, n31049, n31050,
         n31051, n31052, n31053, n31054, n31055, n31056, n31057, n31058,
         n31059, n31060, n31061, n31062, n31063, n31064, n31065, n31066,
         n31067, n31068, n31069, n31070, n31071, n31072, n31073, n31074,
         n31075, n31076, n31077, n31078, n31079, n31080, n31081, n31082,
         n31083, n31084, n31085, n31086, n31087, n31088, n31089, n31090,
         n31091, n31092, n31093, n31094, n31095, n31096, n31097, n31098,
         n31099, n31100, n31101, n31102, n31103, n31104, n31105, n31106,
         n31107, n31108, n31109, n31110, n31111, n31112, n31113, n31114,
         n31115, n31116, n31117, n31118, n31119, n31120, n31121, n31122,
         n31123, n31124, n31125, n31126, n31127, n31128, n31129, n31130,
         n31131, n31132, n31133, n31134, n31135, n31136, n31137, n31138,
         n31139, n31140, n31141, n31142, n31143, n31144, n31145, n31146,
         n31147, n31148, n31149, n31150, n31151, n31152, n31153, n31154,
         n31155, n31156, n31157, n31158, n31159, n31160, n31161, n31162,
         n31163, n31164, n31165, n31166, n31167, n31168, n31169, n31170,
         n31171, n31172, n31173, n31174, n31175, n31176, n31177, n31178,
         n31179, n31180, n31181, n31182, n31183, n31184, n31185, n31186,
         n31187, n31188, n31189, n31190, n31191, n31192, n31193, n31194,
         n31195, n31196, n31197, n31198, n31199, n31200, n31201, n31202,
         n31203, n31204, n31205, n31206, n31207, n31208, n31209, n31210,
         n31211, n31212, n31213, n31214, n31215, n31216, n31217, n31218,
         n31219, n31220, n31221, n31222, n31223, n31224, n31225, n31226,
         n31227, n31228, n31229, n31230, n31231, n31232, n31233, n31234,
         n31235, n31236, n31237, n31238, n31239, n31240, n31241, n31242,
         n31243, n31244, n31245, n31246, n31247, n31248, n31249, n31250,
         n31251, n31252, n31253, n31254, n31255, n31256, n31257, n31258,
         n31259, n31260, n31261, n31262, n31263, n31264, n31265, n31266,
         n31267, n31268, n31269, n31270, n31271, n31272, n31273, n31274,
         n31275, n31276, n31277, n31278, n31279, n31280, n31281, n31282,
         n31283, n31284, n31285, n31286, n31287, n31288, n31289, n31290,
         n31291, n31292, n31293, n31294, n31295, n31296, n31297, n31298,
         n31299, n31300, n31301, n31302, n31303, n31304, n31305, n31306,
         n31307, n31308, n31309, n31310, n31311, n31312, n31313, n31314,
         n31315, n31316, n31317, n31318, n31319, n31320, n31321, n31322,
         n31323, n31324, n31325, n31326, n31327, n31328, n31329, n31330,
         n31331, n31332, n31333, n31334, n31335, n31336, n31337, n31338,
         n31339, n31340, n31341, n31342, n31343, n31344, n31345, n31346,
         n31347, n31348, n31349, n31350, n31351, n31352, n31353, n31354,
         n31355, n31356, n31357, n31358, n31359, n31360, n31361, n31362,
         n31363, n31364, n31365, n31366, n31367, n31368, n31369, n31370,
         n31371, n31372, n31373, n31374, n31375, n31376, n31377, n31378,
         n31379, n31380, n31381, n31382, n31383, n31384, n31385, n31386,
         n31387, n31388, n31389, n31390, n31391, n31392, n31393, n31394,
         n31395, n31396, n31397, n31398, n31399, n31400, n31401, n31402,
         n31403, n31404, n31405, n31406, n31407, n31408, n31409, n31410,
         n31411, n31412, n31413, n31414, n31415, n31416, n31417, n31418,
         n31419, n31420, n31421, n31422, n31423, n31424, n31425, n31426,
         n31427, n31428, n31429, n31430, n31431, n31432, n31433, n31434,
         n31435, n31436, n31437, n31438, n31439, n31440, n31441, n31442,
         n31443, n31444, n31445, n31446, n31447, n31448, n31449, n31450,
         n31451, n31452, n31453, n31454, n31455, n31456, n31457, n31458,
         n31459, n31460, n31461, n31462, n31463, n31464, n31465, n31466,
         n31467, n31468, n31469, n31470, n31471, n31472, n31473, n31474,
         n31475, n31476, n31477, n31478, n31479, n31480, n31481, n31482,
         n31483, n31484, n31485, n31486, n31487, n31488, n31489, n31490,
         n31491, n31492, n31493, n31494, n31495, n31496, n31497, n31498,
         n31499, n31500, n31501, n31502, n31503, n31504, n31505, n31506,
         n31507, n31508, n31509, n31510, n31511, n31512, n31513, n31514,
         n31515, n31516, n31517, n31518, n31519, n31520, n31521, n31522,
         n31523, n31524, n31525, n31526, n31527, n31528, n31529, n31530,
         n31531, n31532, n31533, n31534, n31535, n31536, n31537, n31538,
         n31539, n31540, n31541, n31542, n31543, n31544, n31545, n31546,
         n31547, n31548, n31549, n31550, n31551, n31552, n31553, n31554,
         n31555, n31556, n31557, n31558, n31559, n31560, n31561, n31562,
         n31563, n31564, n31565, n31566, n31567, n31568, n31569, n31570,
         n31571, n31572, n31573, n31574, n31575, n31576, n31577, n31578,
         n31579, n31580, n31581, n31582, n31583, n31584, n31585, n31586,
         n31587, n31588, n31589, n31590, n31591, n31592, n31593, n31594,
         n31595, n31596, n31597, n31598, n31599, n31600, n31601, n31602,
         n31603, n31604, n31605, n31606, n31607, n31608, n31609, n31610,
         n31611, n31612, n31613, n31614, n31615, n31616, n31617, n31618,
         n31619, n31620, n31621, n31622, n31623, n31624, n31625, n31626,
         n31627, n31628, n31629, n31630, n31631, n31632, n31633, n31634,
         n31635, n31636, n31637, n31638, n31639, n31640, n31641, n31642,
         n31643, n31644, n31645, n31646, n31647, n31648, n31649, n31650,
         n31651, n31652, n31653, n31654, n31655, n31656, n31657, n31658,
         n31659, n31660, n31661, n31662, n31663, n31664, n31665, n31666,
         n31667, n31668, n31669, n31670, n31671, n31672, n31673, n31674,
         n31675, n31676, n31677, n31678, n31679, n31680, n31681, n31682,
         n31683, n31684, n31685, n31686, n31687, n31688, n31689, n31690,
         n31691, n31692, n31693, n31694, n31695, n31696, n31697, n31698,
         n31699, n31700, n31701, n31702, n31703, n31704, n31705, n31706,
         n31707, n31708, n31709, n31710, n31711, n31712, n31713, n31714,
         n31715, n31716, n31717, n31718, n31719, n31720, n31721, n31722,
         n31723, n31724, n31725, n31726, n31727, n31728, n31729, n31730,
         n31731, n31732, n31733, n31734, n31735, n31736, n31737, n31738,
         n31739, n31740, n31741, n31742, n31743, n31744, n31745, n31746,
         n31747, n31748, n31749, n31750, n31751, n31752, n31753, n31754,
         n31755, n31756, n31757, n31758, n31759, n31760, n31761, n31762,
         n31763, n31764, n31765, n31766, n31767, n31768, n31769, n31770,
         n31771, n31772, n31773, n31774, n31775, n31776, n31777, n31778,
         n31779, n31780, n31781, n31782, n31783, n31784, n31785, n31786,
         n31787, n31788, n31789, n31790, n31791, n31792, n31793, n31794,
         n31795, n31796, n31797, n31798, n31799, n31800, n31801, n31802,
         n31803, n31804, n31805, n31806, n31807, n31808, n31809, n31810,
         n31811, n31812, n31813, n31814, n31815, n31816, n31817, n31818,
         n31819, n31820, n31821, n31822, n31823, n31824, n31825, n31826,
         n31827, n31828, n31829, n31830, n31831, n31832, n31833, n31834,
         n31835, n31836, n31837, n31838, n31839, n31840, n31841, n31842,
         n31843, n31844, n31845, n31846, n31847, n31848, n31849, n31850,
         n31851, n31852, n31853, n31854, n31855, n31856, n31857, n31858,
         n31859, n31860, n31861, n31862, n31863, n31864, n31865, n31866,
         n31867, n31868, n31869, n31870, n31871, n31872, n31873, n31874,
         n31875, n31876, n31877, n31878, n31879, n31880, n31881, n31882,
         n31883, n31884, n31885, n31886, n31887, n31888, n31889, n31890,
         n31891, n31892, n31893, n31894, n31895, n31896, n31897, n31898,
         n31899, n31900, n31901, n31902, n31903, n31904, n31905, n31906,
         n31907, n31908, n31909, n31910, n31911, n31912, n31913, n31914,
         n31915, n31916, n31917, n31918, n31919, n31920, n31921, n31922,
         n31923, n31924, n31925, n31926, n31927, n31928, n31929, n31930,
         n31931, n31932, n31933, n31934, n31935, n31936, n31937, n31938,
         n31939, n31940, n31941, n31942, n31943, n31944, n31945, n31946,
         n31947, n31948, n31949, n31950, n31951, n31952, n31953, n31954,
         n31955, n31956, n31957, n31958, n31959, n31960, n31961, n31962,
         n31963, n31964, n31965, n31966, n31967, n31968, n31969, n31970,
         n31971, n31972, n31973, n31974, n31975, n31976, n31977, n31978,
         n31979, n31980, n31981, n31982, n31983, n31984, n31985, n31986,
         n31987, n31988, n31989, n31990, n31991, n31992, n31993, n31994,
         n31995, n31996, n31997, n31998, n31999, n32000, n32001, n32002,
         n32003, n32004, n32005, n32006, n32007, n32008, n32009, n32010,
         n32011, n32012, n32013, n32014, n32015, n32016, n32017, n32018,
         n32019, n32020, n32021, n32022, n32023, n32024, n32025, n32026,
         n32027, n32028, n32029, n32030, n32031, n32032, n32033, n32034,
         n32035, n32036, n32037, n32038, n32039, n32040, n32041, n32042,
         n32043, n32044, n32045, n32046, n32047, n32048, n32049, n32050,
         n32051, n32052, n32053, n32054, n32055, n32056, n32057, n32058,
         n32059, n32060, n32061, n32062, n32063, n32064, n32065, n32066,
         n32067, n32068, n32069, n32070, n32071, n32072, n32073, n32074,
         n32075, n32076, n32077, n32078, n32079, n32080, n32081, n32082,
         n32083, n32084, n32085, n32086, n32087, n32088, n32089, n32090,
         n32091, n32092, n32093, n32094, n32095, n32096, n32097, n32098,
         n32099, n32100, n32101, n32102, n32103, n32104, n32105, n32106,
         n32107, n32108, n32109, n32110, n32111, n32112, n32113, n32114,
         n32115, n32116, n32117, n32118, n32119, n32120, n32121, n32122,
         n32123, n32124, n32125, n32126, n32127, n32128, n32129, n32130,
         n32131, n32132, n32133, n32134, n32135, n32136, n32137, n32138,
         n32139, n32140, n32141, n32142, n32143, n32144, n32145, n32146,
         n32147, n32148, n32149, n32150, n32151, n32152, n32153, n32154,
         n32155, n32156, n32157, n32158, n32159, n32160, n32161, n32162,
         n32163, n32164, n32165, n32166, n32167, n32168, n32169, n32170,
         n32171, n32172, n32173, n32174, n32175, n32176, n32177, n32178,
         n32179, n32180, n32181, n32182, n32183, n32184, n32185, n32186,
         n32187, n32188, n32189, n32190, n32191, n32192, n32193, n32194,
         n32195, n32196, n32197, n32198, n32199, n32200, n32201, n32202,
         n32203, n32204, n32205, n32206, n32207, n32208, n32209, n32210,
         n32211, n32212, n32213, n32214, n32215, n32216, n32217, n32218,
         n32219, n32220, n32221, n32222, n32223, n32224, n32225, n32226,
         n32227, n32228, n32229, n32230, n32231, n32232, n32233, n32234,
         n32235, n32236, n32237, n32238, n32239, n32240, n32241, n32242,
         n32243, n32244, n32245, n32246, n32247, n32248, n32249, n32250,
         n32251, n32252, n32253, n32254, n32255, n32256, n32257, n32258,
         n32259, n32260, n32261, n32262, n32263, n32264, n32265, n32266,
         n32267, n32268, n32269, n32270, n32271, n32272, n32273, n32274,
         n32275, n32276, n32277, n32278, n32279, n32280, n32281, n32282,
         n32283, n32284, n32285, n32286, n32287, n32288, n32289, n32290,
         n32291, n32292, n32293, n32294, n32295, n32296, n32297, n32298,
         n32299, n32300, n32301, n32302, n32303, n32304, n32305, n32306,
         n32307, n32308, n32309, n32310, n32311, n32312, n32313, n32314,
         n32315, n32316, n32317, n32318, n32319, n32320, n32321, n32322,
         n32323, n32324, n32325, n32326, n32327, n32328, n32329, n32330,
         n32331, n32332, n32333, n32334, n32335, n32336, n32337, n32338,
         n32339, n32340, n32341, n32342, n32343, n32344, n32345, n32346,
         n32347, n32348, n32349, n32350, n32351, n32352, n32353, n32354,
         n32355, n32356, n32357, n32358, n32359, n32360, n32361, n32362,
         n32363, n32364, n32365, n32366, n32367, n32368, n32369, n32370,
         n32371, n32372, n32373, n32374, n32375, n32376, n32377, n32378,
         n32379, n32380, n32381, n32382, n32383, n32384, n32385, n32386,
         n32387, n32388, n32389, n32390, n32391, n32392, n32393, n32394,
         n32395, n32396, n32397, n32398, n32399, n32400, n32401, n32402,
         n32403, n32404, n32405, n32406, n32407, n32408, n32409, n32410,
         n32411, n32412, n32413, n32414, n32415, n32416, n32417, n32418,
         n32419, n32420, n32421, n32422, n32423, n32424, n32425, n32426,
         n32427, n32428, n32429, n32430, n32431, n32432, n32433, n32434,
         n32435, n32436, n32437, n32438, n32439, n32440, n32441, n32442,
         n32443, n32444, n32445, n32446, n32447, n32448, n32449, n32450,
         n32451, n32452, n32453, n32454, n32455, n32456, n32457, n32458,
         n32459, n32460, n32461, n32462, n32463, n32464, n32465, n32466,
         n32467, n32468, n32469, n32470, n32471, n32472, n32473, n32474,
         n32475, n32476, n32477, n32478, n32479, n32480, n32481, n32482,
         n32483, n32484, n32485, n32486, n32487, n32488, n32489, n32490,
         n32491, n32492, n32493, n32494, n32495, n32496, n32497, n32498,
         n32499, n32500, n32501, n32502, n32503, n32504, n32505, n32506,
         n32507, n32508, n32509, n32510, n32511, n32512, n32513, n32514,
         n32515, n32516, n32517, n32518, n32519, n32520, n32521, n32522,
         n32523, n32524, n32525, n32526, n32527, n32528, n32529, n32530,
         n32531, n32532, n32533, n32534, n32535, n32536, n32537, n32538,
         n32539, n32540, n32541, n32542, n32543, n32544, n32545, n32546,
         n32547, n32548, n32549, n32550, n32551, n32552, n32553, n32554,
         n32555, n32556, n32557, n32558, n32559, n32560, n32561, n32562,
         n32563, n32564, n32565, n32566, n32567, n32568, n32569, n32570,
         n32571, n32572, n32573, n32574, n32575, n32576, n32577, n32578,
         n32579, n32580, n32581, n32582, n32583, n32584, n32585, n32586,
         n32587, n32588, n32589, n32590, n32591, n32592, n32593, n32594,
         n32595, n32596, n32597, n32598, n32599, n32600, n32601, n32602,
         n32603, n32604, n32605, n32606, n32607, n32608, n32609, n32610,
         n32611, n32612, n32613, n32614, n32615, n32616, n32617, n32618,
         n32619, n32620, n32621, n32622, n32623, n32624, n32625, n32626,
         n32627, n32628, n32629, n32630, n32631, n32632, n32633, n32634,
         n32635, n32636, n32637, n32638, n32639, n32640, n32641, n32642,
         n32643, n32644, n32645, n32646, n32647, n32648, n32649, n32650,
         n32651, n32652, n32653, n32654, n32655, n32656, n32657, n32658,
         n32659, n32660, n32661, n32662, n32663, n32664, n32665, n32666,
         n32667, n32668, n32669, n32670, n32671, n32672, n32673, n32674,
         n32675, n32676, n32677, n32678, n32679, n32680, n32681, n32682,
         n32683, n32684, n32685, n32686, n32687, n32688, n32689, n32690,
         n32691, n32692, n32693, n32694, n32695, n32696, n32697, n32698,
         n32699, n32700, n32701, n32702, n32703, n32704, n32705, n32706,
         n32707, n32708, n32709, n32710, n32711, n32712, n32713, n32714,
         n32715, n32716, n32717, n32718, n32719, n32720, n32721, n32722,
         n32723, n32724, n32725, n32726, n32727, n32728, n32729, n32730,
         n32731, n32732, n32733, n32734, n32735, n32736, n32737, n32738,
         n32739, n32740, n32741, n32742, n32743, n32744, n32745, n32746,
         n32747, n32748, n32749, n32750, n32751, n32752, n32753, n32754,
         n32755, n32756, n32757, n32758, n32759, n32760, n32761, n32762,
         n32763, n32764, n32765, n32766, n32767, n32768, n32769, n32770,
         n32771, n32772, n32773, n32774, n32775, n32776, n32777, n32778,
         n32779, n32780, n32781, n32782, n32783, n32784, n32785, n32786,
         n32787, n32788, n32789, n32790, n32791, n32792, n32793, n32794,
         n32795, n32796, n32797, n32798, n32799, n32800, n32801, n32802,
         n32803, n32804, n32805, n32806, n32807, n32808, n32809, n32810,
         n32811, n32812, n32813, n32814, n32815, n32816, n32817, n32818,
         n32819, n32820, n32821, n32822, n32823, n32824, n32825, n32826,
         n32827, n32828, n32829, n32830, n32831, n32832, n32833, n32834,
         n32835, n32836, n32837, n32838, n32839, n32840, n32841, n32842,
         n32843, n32844, n32845, n32846, n32847, n32848, n32849, n32850,
         n32851, n32852, n32853, n32854, n32855, n32856, n32857, n32858,
         n32859, n32860, n32861, n32862, n32863, n32864, n32865, n32866,
         n32867, n32868, n32869, n32870, n32871, n32872, n32873, n32874,
         n32875, n32876, n32877, n32878, n32879, n32880, n32881, n32882,
         n32883, n32884, n32885, n32886, n32887, n32888, n32889, n32890,
         n32891, n32892, n32893, n32894, n32895, n32896, n32897, n32898,
         n32899, n32900, n32901, n32902, n32903, n32904, n32905, n32906,
         n32907, n32908, n32909, n32910, n32911, n32912, n32913, n32914,
         n32915, n32916, n32917, n32918, n32919, n32920, n32921, n32922,
         n32923, n32924, n32925, n32926, n32927, n32928, n32929, n32930,
         n32931, n32932, n32933, n32934, n32935, n32936, n32937, n32938,
         n32939, n32940, n32941, n32942, n32943, n32944, n32945, n32946,
         n32947, n32948, n32949, n32950, n32951, n32952, n32953, n32954,
         n32955, n32956, n32957, n32958, n32959, n32960, n32961, n32962,
         n32963, n32964, n32965, n32966, n32967, n32968, n32969, n32970,
         n32971, n32972, n32973, n32974, n32975, n32976, n32977, n32978,
         n32979, n32980, n32981, n32982, n32983, n32984, n32985, n32986,
         n32987, n32988, n32989, n32990, n32991, n32992, n32993, n32994,
         n32995, n32996, n32997, n32998, n32999, n33000, n33001, n33002,
         n33003, n33004, n33005, n33006, n33007, n33008, n33009, n33010,
         n33011, n33012, n33013, n33014, n33015, n33016, n33017, n33018,
         n33019, n33020, n33021, n33022, n33023, n33024, n33025, n33026,
         n33027, n33028, n33029, n33030, n33031, n33032, n33033, n33034,
         n33035, n33036, n33037, n33038, n33039, n33040, n33041, n33042,
         n33043, n33044, n33045, n33046, n33047, n33048, n33049, n33050,
         n33051, n33052, n33053, n33054, n33055, n33056, n33057, n33058,
         n33059, n33060, n33061, n33062, n33063, n33064, n33065, n33066,
         n33067, n33068, n33069, n33070, n33071, n33072, n33073, n33074,
         n33075, n33076, n33077, n33078, n33079, n33080, n33081, n33082,
         n33083, n33084, n33085, n33086, n33087, n33088, n33089, n33090,
         n33091, n33092, n33093, n33094, n33095, n33096, n33097, n33098,
         n33099, n33100, n33101, n33102, n33103, n33104, n33105, n33106,
         n33107, n33108, n33109, n33110, n33111, n33112, n33113, n33114,
         n33115, n33116, n33117, n33118, n33119, n33120, n33121, n33122,
         n33123, n33124, n33125, n33126, n33127, n33128, n33129, n33130,
         n33131, n33132, n33133, n33134, n33135, n33136, n33137, n33138,
         n33139, n33140, n33141, n33142, n33143, n33144, n33145, n33146,
         n33147, n33148, n33149, n33150, n33151, n33152, n33153, n33154,
         n33155, n33156, n33157, n33158, n33159, n33160, n33161, n33162,
         n33163, n33164, n33165, n33166, n33167, n33168, n33169, n33170,
         n33171, n33172, n33173, n33174, n33175, n33176, n33177, n33178,
         n33179, n33180, n33181, n33182, n33183, n33184, n33185, n33186,
         n33187, n33188, n33189, n33190, n33191, n33192, n33193, n33194,
         n33195, n33196, n33197, n33198, n33199, n33200, n33201, n33202,
         n33203, n33204, n33205, n33206, n33207, n33208, n33209, n33210,
         n33211, n33212, n33213, n33214, n33215, n33216, n33217, n33218,
         n33219, n33220, n33221, n33222, n33223, n33224, n33225, n33226,
         n33227, n33228, n33229, n33230, n33231, n33232, n33233, n33234,
         n33235, n33236, n33237, n33238, n33239, n33240, n33241, n33242,
         n33243, n33244, n33245, n33246, n33247, n33248, n33249, n33250,
         n33251, n33252, n33253, n33254, n33255, n33256, n33257, n33258,
         n33259, n33260, n33261, n33262, n33263, n33264, n33265, n33266,
         n33267, n33268, n33269, n33270, n33271, n33272, n33273, n33274,
         n33275, n33276, n33277, n33278, n33279, n33280, n33281, n33282,
         n33283, n33284, n33285, n33286, n33287, n33288, n33289, n33290,
         n33291, n33292, n33293, n33294, n33295, n33296, n33297, n33298,
         n33299, n33300, n33301, n33302, n33303, n33304, n33305, n33306,
         n33307, n33308, n33309, n33310, n33311, n33312, n33313, n33314,
         n33315, n33316, n33317, n33318, n33319, n33320, n33321, n33322,
         n33323, n33324, n33325, n33326, n33327, n33328, n33329, n33330,
         n33331, n33332, n33333, n33334, n33335, n33336, n33337, n33338,
         n33339, n33340, n33341, n33342, n33343, n33344, n33345, n33346,
         n33347, n33348, n33349, n33350, n33351, n33352, n33353, n33354,
         n33355, n33356, n33357, n33358, n33359, n33360, n33361, n33362,
         n33363, n33364, n33365, n33366, n33367, n33368, n33369, n33370,
         n33371, n33372, n33373, n33374, n33375, n33376, n33377, n33378,
         n33379, n33380, n33381, n33382, n33383, n33384, n33385, n33386,
         n33387, n33388, n33389, n33390, n33391, n33392, n33393, n33394,
         n33395, n33396, n33397, n33398, n33399, n33400, n33401, n33402,
         n33403, n33404, n33405, n33406, n33407, n33408, n33409, n33410,
         n33411, n33412, n33413, n33414, n33415, n33416, n33417, n33418,
         n33419, n33420, n33421, n33422, n33423, n33424, n33425, n33426,
         n33427, n33428, n33429, n33430, n33431, n33432, n33433, n33434,
         n33435, n33436, n33437, n33438, n33439, n33440, n33441, n33442,
         n33443, n33444, n33445, n33446, n33447, n33448, n33449, n33450,
         n33451, n33452, n33453, n33454, n33455, n33456, n33457, n33458,
         n33459, n33460, n33461, n33462, n33463, n33464, n33465, n33466,
         n33467, n33468, n33469, n33470, n33471, n33472, n33473, n33474,
         n33475, n33476, n33477, n33478, n33479, n33480, n33481, n33482,
         n33483, n33484, n33485, n33486, n33487, n33488, n33489, n33490,
         n33491, n33492, n33493, n33494, n33495, n33496, n33497, n33498,
         n33499, n33500, n33501, n33502, n33503, n33504, n33505, n33506,
         n33507, n33508, n33509, n33510, n33511, n33512, n33513, n33514,
         n33515, n33516, n33517, n33518, n33519, n33520, n33521, n33522,
         n33523, n33524, n33525, n33526, n33527, n33528, n33529, n33530,
         n33531, n33532, n33533, n33534, n33535, n33536, n33537, n33538,
         n33539, n33540, n33541, n33542, n33543, n33544, n33545, n33546,
         n33547, n33548, n33549, n33550, n33551, n33552, n33553, n33554,
         n33555, n33556, n33557, n33558, n33559, n33560, n33561, n33562,
         n33563, n33564, n33565, n33566, n33567, n33568, n33569, n33570,
         n33571, n33572, n33573, n33574, n33575, n33576, n33577, n33578,
         n33579, n33580, n33581, n33582, n33583, n33584, n33585, n33586,
         n33587, n33588, n33589, n33590, n33591, n33592, n33593, n33594,
         n33595, n33596, n33597, n33598, n33599, n33600, n33601, n33602,
         n33603, n33604, n33605, n33606, n33607, n33608, n33609, n33610,
         n33611, n33612, n33613, n33614, n33615, n33616, n33617, n33618,
         n33619, n33620, n33621, n33622, n33623, n33624, n33625, n33626,
         n33627, n33628, n33629, n33630, n33631, n33632, n33633, n33634,
         n33635, n33636, n33637, n33638, n33639, n33640, n33641, n33642,
         n33643, n33644, n33645, n33646, n33647, n33648, n33649, n33650,
         n33651, n33652, n33653, n33654, n33655, n33656, n33657, n33658,
         n33659, n33660, n33661, n33662, n33663, n33664, n33665, n33666,
         n33667, n33668, n33669, n33670, n33671, n33672, n33673, n33674,
         n33675, n33676, n33677, n33678, n33679, n33680, n33681, n33682,
         n33683, n33684, n33685, n33686, n33687, n33688, n33689, n33690,
         n33691, n33692, n33693, n33694, n33695, n33696, n33697, n33698,
         n33699, n33700, n33701, n33702, n33703, n33704, n33705, n33706,
         n33707, n33708, n33709, n33710, n33711, n33712, n33713, n33714,
         n33715, n33716, n33717, n33718, n33719, n33720, n33721, n33722,
         n33723, n33724, n33725, n33726, n33727, n33728, n33729, n33730,
         n33731, n33732, n33733, n33734, n33735, n33736, n33737, n33738,
         n33739, n33740, n33741, n33742, n33743, n33744, n33745, n33746,
         n33747, n33748, n33749, n33750, n33751, n33752, n33753, n33754,
         n33755, n33756, n33757, n33758, n33759, n33760, n33761, n33762,
         n33763, n33764, n33765, n33766, n33767, n33768, n33769, n33770,
         n33771, n33772, n33773, n33774, n33775, n33776, n33777, n33778,
         n33779, n33780, n33781, n33782, n33783, n33784, n33785, n33786,
         n33787, n33788, n33789, n33790, n33791, n33792, n33793, n33794,
         n33795, n33796, n33797, n33798, n33799, n33800, n33801, n33802,
         n33803, n33804, n33805, n33806, n33807, n33808, n33809, n33810,
         n33811, n33812, n33813, n33814, n33815, n33816, n33817, n33818,
         n33819, n33820, n33821, n33822, n33823, n33824, n33825, n33826,
         n33827, n33828, n33829, n33830, n33831, n33832, n33833, n33834,
         n33835, n33836, n33837, n33838, n33839, n33840, n33841, n33842,
         n33843, n33844, n33845, n33846, n33847, n33848, n33849, n33850,
         n33851, n33852, n33853, n33854, n33855, n33856, n33857, n33858,
         n33859, n33860, n33861, n33862, n33863, n33864, n33865, n33866,
         n33867, n33868, n33869, n33870, n33871, n33872, n33873, n33874,
         n33875, n33876, n33877, n33878, n33879, n33880, n33881, n33882,
         n33883, n33884, n33885, n33886, n33887, n33888, n33889, n33890,
         n33891, n33892, n33893, n33894, n33895, n33896, n33897, n33898,
         n33899, n33900, n33901, n33902, n33903, n33904, n33905, n33906,
         n33907, n33908, n33909, n33910, n33911, n33912, n33913, n33914,
         n33915, n33916, n33917, n33918, n33919, n33920, n33921, n33922,
         n33923, n33924, n33925, n33926, n33927, n33928, n33929, n33930,
         n33931, n33932, n33933, n33934, n33935, n33936, n33937, n33938,
         n33939, n33940, n33941, n33942, n33943, n33944, n33945, n33946,
         n33947, n33948, n33949, n33950, n33951, n33952, n33953, n33954,
         n33955, n33956, n33957, n33958, n33959, n33960, n33961, n33962,
         n33963, n33964, n33965, n33966, n33967, n33968, n33969, n33970,
         n33971, n33972, n33973, n33974, n33975, n33976, n33977, n33978,
         n33979, n33980, n33981, n33982, n33983, n33984, n33985, n33986,
         n33987, n33988, n33989, n33990, n33991, n33992, n33993, n33994,
         n33995, n33996, n33997, n33998, n33999, n34000, n34001, n34002,
         n34003, n34004, n34005, n34006, n34007, n34008, n34009, n34010,
         n34011, n34012, n34013, n34014, n34015, n34016, n34017, n34018,
         n34019, n34020, n34021, n34022, n34023, n34024, n34025, n34026,
         n34027, n34028, n34029, n34030, n34031, n34032, n34033, n34034,
         n34035, n34036, n34037, n34038, n34039, n34040, n34041, n34042,
         n34043, n34044, n34045, n34046, n34047, n34048, n34049, n34050,
         n34051, n34052, n34053, n34054, n34055, n34056, n34057, n34058,
         n34059, n34060, n34061, n34062, n34063, n34064, n34065, n34066,
         n34067, n34068, n34069, n34070, n34071, n34072, n34073, n34074,
         n34075, n34076, n34077, n34078, n34079, n34080, n34081, n34082,
         n34083, n34084, n34085, n34086, n34087, n34088, n34089, n34090,
         n34091, n34092, n34093, n34094, n34095, n34096, n34097, n34098,
         n34099, n34100, n34101, n34102, n34103, n34104, n34105, n34106,
         n34107, n34108, n34109, n34110, n34111, n34112, n34113, n34114,
         n34115, n34116, n34117, n34118, n34119, n34120, n34121, n34122,
         n34123, n34124, n34125, n34126, n34127, n34128, n34129, n34130,
         n34131, n34132, n34133, n34134, n34135, n34136, n34137, n34138,
         n34139, n34140, n34141, n34142, n34143, n34144, n34145, n34146,
         n34147, n34148, n34149, n34150, n34151, n34152, n34153, n34154,
         n34155, n34156, n34157, n34158, n34159, n34160, n34161, n34162,
         n34163, n34164, n34165, n34166, n34167, n34168, n34169, n34170,
         n34171, n34172, n34173, n34174, n34175, n34176, n34177, n34178,
         n34179, n34180, n34181, n34182, n34183, n34184, n34185, n34186,
         n34187, n34188, n34189, n34190, n34191, n34192, n34193, n34194,
         n34195, n34196, n34197, n34198, n34199, n34200, n34201, n34202,
         n34203, n34204, n34205, n34206, n34207, n34208, n34209, n34210,
         n34211, n34212, n34213, n34214, n34215, n34216, n34217, n34218,
         n34219, n34220, n34221, n34222, n34223, n34224, n34225, n34226,
         n34227, n34228, n34229, n34230, n34231, n34232, n34233, n34234,
         n34235, n34236, n34237, n34238, n34239, n34240, n34241, n34242,
         n34243, n34244, n34245, n34246, n34247, n34248, n34249, n34250,
         n34251, n34252, n34253, n34254, n34255, n34256, n34257, n34258,
         n34259, n34260, n34261, n34262, n34263, n34264, n34265, n34266,
         n34267, n34268, n34269, n34270, n34271, n34272, n34273, n34274,
         n34275, n34276, n34277, n34278, n34279, n34280, n34281, n34282,
         n34283, n34284, n34285, n34286, n34287, n34288, n34289, n34290,
         n34291, n34292, n34293, n34294, n34295, n34296, n34297, n34298,
         n34299, n34300, n34301, n34302, n34303, n34304, n34305, n34306,
         n34307, n34308, n34309, n34310, n34311, n34312, n34313, n34314,
         n34315, n34316, n34317, n34318, n34319, n34320, n34321, n34322,
         n34323, n34324, n34325, n34326, n34327, n34328, n34329, n34330,
         n34331, n34332, n34333, n34334, n34335, n34336, n34337, n34338,
         n34339, n34340, n34341, n34342, n34343, n34344, n34345, n34346,
         n34347, n34348, n34349, n34350, n34351, n34352, n34353, n34354,
         n34355, n34356, n34357, n34358, n34359, n34360, n34361, n34362,
         n34363, n34364, n34365, n34366, n34367, n34368, n34369, n34370,
         n34371, n34372, n34373, n34374, n34375, n34376, n34377, n34378,
         n34379, n34380, n34381, n34382, n34383, n34384, n34385, n34386,
         n34387, n34388, n34389, n34390, n34391, n34392, n34393, n34394,
         n34395, n34396, n34397, n34398, n34399, n34400, n34401, n34402,
         n34403, n34404, n34405, n34406, n34407, n34408, n34409, n34410,
         n34411, n34412, n34413, n34414, n34415, n34416, n34417, n34418,
         n34419, n34420, n34421, n34422, n34423, n34424, n34425, n34426,
         n34427, n34428, n34429, n34430, n34431, n34432, n34433, n34434,
         n34435, n34436, n34437, n34438, n34439, n34440, n34441, n34442,
         n34443, n34444, n34445, n34446, n34447, n34448, n34449, n34450,
         n34451, n34452, n34453, n34454, n34455, n34456, n34457, n34458,
         n34459, n34460, n34461, n34462, n34463, n34464, n34465, n34466,
         n34467, n34468, n34469, n34470, n34471, n34472, n34473, n34474,
         n34475, n34476, n34477, n34478, n34479, n34480, n34481, n34482,
         n34483, n34484, n34485, n34486, n34487, n34488, n34489, n34490,
         n34491, n34492, n34493, n34494, n34495, n34496, n34497, n34498,
         n34499, n34500, n34501, n34502, n34503, n34504, n34505, n34506,
         n34507, n34508, n34509, n34510, n34511, n34512, n34513, n34514,
         n34515, n34516, n34517, n34518, n34519, n34520, n34521, n34522,
         n34523, n34524, n34525, n34526, n34527, n34528, n34529, n34530,
         n34531, n34532, n34533, n34534, n34535, n34536, n34537, n34538,
         n34539, n34540, n34541, n34542, n34543, n34544, n34545, n34546,
         n34547, n34548, n34549, n34550, n34551, n34552, n34553, n34554,
         n34555, n34556, n34557, n34558, n34559, n34560, n34561, n34562,
         n34563, n34564, n34565, n34566, n34567, n34568, n34569, n34570,
         n34571, n34572, n34573, n34574, n34575, n34576, n34577, n34578,
         n34579, n34580, n34581, n34582, n34583, n34584, n34585, n34586,
         n34587, n34588, n34589, n34590, n34591, n34592, n34593, n34594,
         n34595, n34596, n34597, n34598, n34599, n34600, n34601, n34602,
         n34603, n34604, n34605, n34606, n34607, n34608, n34609, n34610,
         n34611, n34612, n34613, n34614, n34615, n34616, n34617, n34618,
         n34619, n34620, n34621, n34622, n34623, n34624, n34625, n34626,
         n34627, n34628, n34629, n34630, n34631, n34632, n34633, n34634,
         n34635, n34636, n34637, n34638, n34639, n34640, n34641, n34642,
         n34643, n34644, n34645, n34646, n34647, n34648, n34649, n34650,
         n34651, n34652, n34653, n34654, n34655, n34656, n34657, n34658,
         n34659, n34660, n34661, n34662, n34663, n34664, n34665, n34666,
         n34667, n34668, n34669, n34670, n34671, n34672, n34673, n34674,
         n34675, n34676, n34677, n34678, n34679, n34680, n34681, n34682,
         n34683, n34684, n34685, n34686, n34687, n34688, n34689, n34690,
         n34691, n34692, n34693, n34694, n34695, n34696, n34697, n34698,
         n34699, n34700, n34701, n34702, n34703, n34704, n34705, n34706,
         n34707, n34708, n34709, n34710, n34711, n34712, n34713, n34714,
         n34715, n34716, n34717, n34718, n34719, n34720, n34721, n34722,
         n34723, n34724, n34725, n34726, n34727, n34728, n34729, n34730,
         n34731, n34732, n34733, n34734, n34735, n34736, n34737, n34738,
         n34739, n34740, n34741, n34742, n34743, n34744, n34745, n34746,
         n34747, n34748, n34749, n34750, n34751, n34752, n34753, n34754,
         n34755, n34756, n34757, n34758, n34759, n34760, n34761, n34762,
         n34763, n34764, n34765, n34766, n34767, n34768, n34769, n34770,
         n34771, n34772, n34773, n34774, n34775, n34776, n34777, n34778,
         n34779, n34780, n34781, n34782, n34783, n34784, n34785, n34786,
         n34787, n34788, n34789, n34790, n34791, n34792, n34793, n34794,
         n34795, n34796, n34797, n34798, n34799, n34800, n34801, n34802,
         n34803, n34804, n34805, n34806, n34807, n34808, n34809, n34810,
         n34811, n34812, n34813, n34814, n34815, n34816, n34817, n34818,
         n34819, n34820, n34821, n34822, n34823, n34824, n34825, n34826,
         n34827, n34828, n34829, n34830, n34831, n34832, n34833, n34834,
         n34835, n34836, n34837, n34838, n34839, n34840, n34841, n34842,
         n34843, n34844, n34845, n34846, n34847, n34848, n34849, n34850,
         n34851, n34852, n34853, n34854, n34855, n34856, n34857, n34858,
         n34859, n34860, n34861, n34862, n34863, n34864, n34865, n34866,
         n34867, n34868, n34869, n34870, n34871, n34872, n34873, n34874,
         n34875, n34876, n34877, n34878, n34879, n34880, n34881, n34882,
         n34883, n34884, n34885, n34886, n34887, n34888, n34889, n34890,
         n34891, n34892, n34893, n34894, n34895, n34896, n34897, n34898,
         n34899, n34900, n34901, n34902, n34903, n34904, n34905, n34906,
         n34907, n34908, n34909, n34910, n34911, n34912, n34913, n34914,
         n34915, n34916, n34917, n34918, n34919, n34920, n34921, n34922,
         n34923, n34924, n34925, n34926, n34927, n34928, n34929, n34930,
         n34931, n34932, n34933, n34934, n34935, n34936, n34937, n34938,
         n34939, n34940, n34941, n34942, n34943, n34944, n34945, n34946,
         n34947, n34948, n34949, n34950, n34951, n34952, n34953, n34954,
         n34955, n34956, n34957, n34958, n34959, n34960, n34961, n34962,
         n34963, n34964, n34965, n34966, n34967, n34968, n34969, n34970,
         n34971, n34972, n34973, n34974, n34975, n34976, n34977, n34978,
         n34979, n34980, n34981, n34982, n34983, n34984, n34985, n34986,
         n34987, n34988, n34989, n34990, n34991, n34992, n34993, n34994,
         n34995, n34996, n34997, n34998, n34999, n35000, n35001, n35002,
         n35003, n35004, n35005, n35006, n35007, n35008, n35009, n35010,
         n35011, n35012, n35013, n35014, n35015, n35016, n35017, n35018,
         n35019, n35020, n35021, n35022, n35023, n35024, n35025, n35026,
         n35027, n35028, n35029, n35030, n35031, n35032, n35033, n35034,
         n35035, n35036, n35037, n35038, n35039, n35040, n35041, n35042,
         n35043, n35044, n35045, n35046, n35047, n35048, n35049, n35050,
         n35051, n35052, n35053, n35054, n35055, n35056, n35057, n35058,
         n35059, n35060, n35061, n35062, n35063, n35064, n35065, n35066,
         n35067, n35068, n35069, n35070, n35071, n35072, n35073, n35074,
         n35075, n35076, n35077, n35078, n35079, n35080, n35081, n35082,
         n35083, n35084, n35085, n35086, n35087, n35088, n35089, n35090,
         n35091, n35092, n35093, n35094, n35095, n35096, n35097, n35098,
         n35099, n35100, n35101, n35102, n35103, n35104, n35105, n35106,
         n35107, n35108, n35109, n35110, n35111, n35112, n35113, n35114,
         n35115, n35116, n35117, n35118, n35119, n35120, n35121, n35122,
         n35123, n35124, n35125, n35126, n35127, n35128, n35129, n35130,
         n35131, n35132, n35133, n35134, n35135, n35136, n35137, n35138,
         n35139, n35140, n35141, n35142, n35143, n35144, n35145, n35146,
         n35147, n35148, n35149, n35150, n35151, n35152, n35153, n35154,
         n35155, n35156, n35157, n35158, n35159, n35160, n35161, n35162,
         n35163, n35164, n35165, n35166, n35167, n35168, n35169, n35170,
         n35171, n35172, n35173, n35174, n35175, n35176, n35177, n35178,
         n35179, n35180, n35181, n35182, n35183, n35184, n35185, n35186,
         n35187, n35188, n35189, n35190, n35191, n35192, n35193, n35194,
         n35195, n35196, n35197, n35198, n35199, n35200, n35201, n35202,
         n35203, n35204, n35205, n35206, n35207, n35208, n35209, n35210,
         n35211, n35212, n35213, n35214, n35215, n35216, n35217, n35218,
         n35219, n35220, n35221, n35222, n35223, n35224, n35225, n35226,
         n35227, n35228, n35229, n35230, n35231, n35232, n35233, n35234,
         n35235, n35236, n35237, n35238, n35239, n35240, n35241, n35242,
         n35243, n35244, n35245, n35246, n35247, n35248, n35249, n35250,
         n35251, n35252, n35253, n35254, n35255, n35256, n35257, n35258,
         n35259, n35260, n35261, n35262, n35263, n35264, n35265, n35266,
         n35267, n35268, n35269, n35270, n35271, n35272, n35273, n35274,
         n35275, n35276, n35277, n35278, n35279, n35280, n35281, n35282,
         n35283, n35284, n35285, n35286, n35287, n35288, n35289, n35290,
         n35291, n35292, n35293, n35294, n35295, n35296, n35297, n35298,
         n35299, n35300, n35301, n35302, n35303, n35304, n35305, n35306,
         n35307, n35308, n35309, n35310, n35311, n35312, n35313, n35314,
         n35315, n35316, n35317, n35318, n35319, n35320, n35321, n35322,
         n35323, n35324, n35325, n35326, n35327, n35328, n35329, n35330,
         n35331, n35332, n35333, n35334, n35335, n35336, n35337, n35338,
         n35339, n35340, n35341, n35342, n35343, n35344, n35345, n35346,
         n35347, n35348, n35349, n35350, n35351, n35352, n35353, n35354,
         n35355, n35356, n35357, n35358, n35359, n35360, n35361, n35362,
         n35363, n35364, n35365, n35366, n35367, n35368, n35369, n35370,
         n35371, n35372, n35373, n35374, n35375, n35376, n35377, n35378,
         n35379, n35380, n35381, n35382, n35383, n35384, n35385, n35386,
         n35387, n35388, n35389, n35390, n35391, n35392, n35393, n35394,
         n35395, n35396, n35397, n35398, n35399, n35400, n35401, n35402,
         n35403, n35404, n35405, n35406, n35407, n35408, n35409, n35410,
         n35411, n35412, n35413, n35414, n35415, n35416, n35417, n35418,
         n35419, n35420, n35421, n35422, n35423, n35424, n35425, n35426,
         n35427, n35428, n35429, n35430, n35431, n35432, n35433, n35434,
         n35435, n35436, n35437, n35438, n35439, n35440, n35441, n35442,
         n35443, n35444, n35445, n35446, n35447, n35448, n35449, n35450,
         n35451, n35452, n35453, n35454, n35455, n35456, n35457, n35458,
         n35459, n35460, n35461, n35462, n35463, n35464, n35465, n35466,
         n35467, n35468, n35469, n35470, n35471, n35472, n35473, n35474,
         n35475, n35476, n35477, n35478, n35479, n35480, n35481, n35482,
         n35483, n35484, n35485, n35486, n35487, n35488, n35489, n35490,
         n35491, n35492, n35493, n35494, n35495, n35496, n35497, n35498,
         n35499, n35500, n35501, n35502, n35503, n35504, n35505, n35506,
         n35507, n35508, n35509, n35510, n35511, n35512, n35513, n35514,
         n35515, n35516, n35517, n35518, n35519, n35520, n35521, n35522,
         n35523, n35524, n35525, n35526, n35527, n35528, n35529, n35530,
         n35531, n35532, n35533, n35534, n35535, n35536, n35537, n35538,
         n35539, n35540, n35541, n35542, n35543, n35544, n35545, n35546,
         n35547, n35548, n35549, n35550, n35551, n35552, n35553, n35554,
         n35555, n35556, n35557, n35558, n35559, n35560, n35561, n35562,
         n35563, n35564, n35565, n35566, n35567, n35568, n35569, n35570,
         n35571, n35572, n35573, n35574, n35575, n35576, n35577, n35578,
         n35579, n35580, n35581, n35582, n35583, n35584, n35585, n35586,
         n35587, n35588, n35589, n35590, n35591, n35592, n35593, n35594,
         n35595, n35596, n35597, n35598, n35599, n35600, n35601, n35602,
         n35603, n35604, n35605, n35606, n35607, n35608, n35609, n35610,
         n35611, n35612, n35613, n35614, n35615, n35616, n35617, n35618,
         n35619, n35620, n35621, n35622, n35623, n35624, n35625, n35626,
         n35627, n35628, n35629, n35630, n35631, n35632, n35633, n35634,
         n35635, n35636, n35637, n35638, n35639, n35640, n35641, n35642,
         n35643, n35644, n35645, n35646, n35647, n35648, n35649, n35650,
         n35651, n35652, n35653, n35654, n35655, n35656, n35657, n35658,
         n35659, n35660, n35661, n35662, n35663, n35664, n35665, n35666,
         n35667, n35668, n35669, n35670, n35671, n35672, n35673, n35674,
         n35675, n35676, n35677, n35678, n35679, n35680, n35681, n35682,
         n35683, n35684, n35685, n35686, n35687, n35688, n35689, n35690,
         n35691, n35692, n35693, n35694, n35695, n35696, n35697, n35698,
         n35699, n35700, n35701, n35702, n35703, n35704, n35705, n35706,
         n35707, n35708, n35709, n35710, n35711, n35712, n35713, n35714,
         n35715, n35716, n35717, n35718, n35719, n35720, n35721, n35722,
         n35723, n35724, n35725, n35726, n35727, n35728, n35729, n35730,
         n35731, n35732, n35733, n35734, n35735, n35736, n35737, n35738,
         n35739, n35740, n35741, n35742, n35743, n35744, n35745, n35746,
         n35747, n35748, n35749, n35750, n35751, n35752, n35753, n35754,
         n35755, n35756, n35757, n35758, n35759, n35760, n35761, n35762,
         n35763, n35764, n35765, n35766, n35767, n35768, n35769, n35770,
         n35771, n35772, n35773, n35774, n35775, n35776, n35777, n35778,
         n35779, n35780, n35781, n35782, n35783, n35784, n35785, n35786,
         n35787, n35788, n35789, n35790, n35791, n35792, n35793, n35794,
         n35795, n35796, n35797, n35798, n35799, n35800, n35801, n35802,
         n35803, n35804, n35805, n35806, n35807, n35808, n35809, n35810,
         n35811, n35812, n35813, n35814, n35815, n35816, n35817, n35818,
         n35819, n35820, n35821, n35822, n35823, n35824, n35825, n35826,
         n35827, n35828, n35829, n35830, n35831, n35832, n35833, n35834,
         n35835, n35836, n35837, n35838, n35839, n35840, n35841, n35842,
         n35843, n35844, n35845, n35846, n35847, n35848, n35849, n35850,
         n35851, n35852, n35853, n35854, n35855, n35856, n35857, n35858,
         n35859, n35860, n35861, n35862, n35863, n35864, n35865, n35866,
         n35867, n35868, n35869, n35870, n35871, n35872, n35873, n35874,
         n35875, n35876, n35877, n35878, n35879, n35880, n35881, n35882,
         n35883, n35884, n35885, n35886, n35887, n35888, n35889, n35890,
         n35891, n35892, n35893, n35894, n35895, n35896, n35897, n35898,
         n35899, n35900, n35901, n35902, n35903, n35904, n35905, n35906,
         n35907, n35908, n35909, n35910, n35911, n35912, n35913, n35914,
         n35915, n35916, n35917, n35918, n35919, n35920, n35921, n35922,
         n35923, n35924, n35925, n35926, n35927, n35928, n35929, n35930,
         n35931, n35932, n35933, n35934, n35935, n35936, n35937, n35938,
         n35939, n35940, n35941, n35942, n35943, n35944, n35945, n35946,
         n35947, n35948, n35949, n35950, n35951, n35952, n35953, n35954,
         n35955, n35956, n35957, n35958, n35959, n35960, n35961, n35962,
         n35963, n35964, n35965, n35966, n35967, n35968, n35969, n35970,
         n35971, n35972, n35973, n35974, n35975, n35976, n35977, n35978,
         n35979, n35980, n35981, n35982, n35983, n35984, n35985, n35986,
         n35987, n35988, n35989, n35990, n35991, n35992, n35993, n35994,
         n35995, n35996, n35997, n35998, n35999, n36000, n36001, n36002,
         n36003, n36004, n36005, n36006, n36007, n36008, n36009, n36010,
         n36011, n36012, n36013, n36014, n36015, n36016, n36017, n36018,
         n36019, n36020, n36021, n36022, n36023, n36024, n36025, n36026,
         n36027, n36028, n36029, n36030, n36031, n36032, n36033, n36034,
         n36035, n36036, n36037, n36038, n36039, n36040, n36041, n36042,
         n36043, n36044, n36045, n36046, n36047, n36048, n36049, n36050,
         n36051, n36052, n36053, n36054, n36055, n36056, n36057, n36058,
         n36059, n36060, n36061, n36062, n36063, n36064, n36065, n36066,
         n36067, n36068, n36069, n36070, n36071, n36072, n36073, n36074,
         n36075, n36076, n36077, n36078, n36079, n36080, n36081, n36082,
         n36083, n36084, n36085, n36086, n36087, n36088, n36089, n36090,
         n36091, n36092, n36093, n36094, n36095, n36096, n36097, n36098,
         n36099, n36100, n36101, n36102, n36103, n36104, n36105, n36106,
         n36107, n36108, n36109, n36110, n36111, n36112, n36113, n36114,
         n36115, n36116, n36117, n36118, n36119, n36120, n36121, n36122,
         n36123, n36124, n36125, n36126, n36127, n36128, n36129, n36130,
         n36131, n36132, n36133, n36134, n36135, n36136, n36137, n36138,
         n36139, n36140, n36141, n36142, n36143, n36144, n36145, n36146,
         n36147, n36148, n36149, n36150, n36151, n36152, n36153, n36154,
         n36155, n36156, n36157, n36158, n36159, n36160, n36161, n36162,
         n36163, n36164, n36165, n36166, n36167, n36168, n36169, n36170,
         n36171, n36172, n36173, n36174, n36175, n36176, n36177, n36178,
         n36179, n36180, n36181, n36182, n36183, n36184, n36185, n36186,
         n36187, n36188, n36189, n36190, n36191, n36192, n36193, n36194,
         n36195, n36196, n36197, n36198, n36199, n36200, n36201, n36202,
         n36203, n36204, n36205, n36206, n36207, n36208, n36209, n36210,
         n36211, n36212, n36213, n36214, n36215, n36216, n36217, n36218,
         n36219, n36220, n36221, n36222, n36223, n36224, n36225, n36226,
         n36227, n36228, n36229, n36230, n36231, n36232, n36233, n36234,
         n36235, n36236, n36237, n36238, n36239, n36240, n36241, n36242,
         n36243, n36244, n36245, n36246, n36247, n36248, n36249, n36250,
         n36251, n36252, n36253, n36254, n36255, n36256, n36257, n36258,
         n36259, n36260, n36261, n36262, n36263, n36264, n36265, n36266,
         n36267, n36268, n36269, n36270, n36271, n36272, n36273, n36274,
         n36275, n36276, n36277, n36278, n36279, n36280, n36281, n36282,
         n36283, n36284, n36285, n36286, n36287, n36288, n36289, n36290,
         n36291, n36292, n36293, n36294, n36295, n36296, n36297, n36298,
         n36299, n36300, n36301, n36302, n36303, n36304, n36305, n36306,
         n36307, n36308, n36309, n36310, n36311, n36312, n36313, n36314,
         n36315, n36316, n36317, n36318, n36319, n36320, n36321, n36322,
         n36323, n36324, n36325, n36326, n36327, n36328, n36329, n36330,
         n36331, n36332, n36333, n36334, n36335, n36336, n36337, n36338,
         n36339, n36340, n36341, n36342, n36343, n36344, n36345, n36346,
         n36347, n36348, n36349, n36350, n36351, n36352, n36353, n36354,
         n36355, n36356, n36357, n36358, n36359, n36360, n36361, n36362,
         n36363, n36364, n36365, n36366, n36367, n36368, n36369, n36370,
         n36371, n36372, n36373, n36374, n36375, n36376, n36377, n36378,
         n36379, n36380, n36381, n36382, n36383, n36384, n36385, n36386,
         n36387, n36388, n36389, n36390, n36391, n36392, n36393, n36394,
         n36395, n36396, n36397, n36398, n36399, n36400, n36401, n36402,
         n36403, n36404, n36405, n36406, n36407, n36408, n36409, n36410,
         n36411, n36412, n36413, n36414, n36415, n36416, n36417, n36418,
         n36419, n36420, n36421, n36422, n36423, n36424, n36425, n36426,
         n36427, n36428, n36429, n36430, n36431, n36432, n36433, n36434,
         n36435, n36436, n36437, n36438, n36439, n36440, n36441, n36442,
         n36443, n36444, n36445, n36446, n36447, n36448, n36449, n36450,
         n36451, n36452, n36453, n36454, n36455, n36456, n36457, n36458,
         n36459, n36460, n36461, n36462, n36463, n36464, n36465, n36466,
         n36467, n36468, n36469, n36470, n36471, n36472, n36473, n36474,
         n36475, n36476, n36477, n36478, n36479, n36480, n36481, n36482,
         n36483, n36484, n36485, n36486, n36487, n36488, n36489, n36490,
         n36491, n36492, n36493, n36494, n36495, n36496, n36497, n36498,
         n36499, n36500, n36501, n36502, n36503, n36504, n36505, n36506,
         n36507, n36508, n36509, n36510, n36511, n36512, n36513, n36514,
         n36515, n36516, n36517, n36518, n36519, n36520, n36521, n36522,
         n36523, n36524, n36525, n36526, n36527, n36528, n36529, n36530,
         n36531, n36532, n36533, n36534, n36535, n36536, n36537, n36538,
         n36539, n36540, n36541, n36542, n36543, n36544, n36545, n36546,
         n36547, n36548, n36549, n36550, n36551, n36552, n36553, n36554,
         n36555, n36556, n36557, n36558, n36559, n36560, n36561, n36562,
         n36563, n36564, n36565, n36566, n36567, n36568, n36569, n36570,
         n36571, n36572, n36573, n36574, n36575, n36576, n36577, n36578,
         n36579, n36580, n36581, n36582, n36583, n36584, n36585, n36586,
         n36587, n36588, n36589, n36590, n36591, n36592, n36593, n36594,
         n36595, n36596, n36597, n36598, n36599, n36600, n36601, n36602,
         n36603, n36604, n36605, n36606, n36607, n36608, n36609, n36610,
         n36611, n36612, n36613, n36614, n36615, n36616, n36617, n36618,
         n36619, n36620, n36621, n36622, n36623, n36624, n36625, n36626,
         n36627, n36628, n36629, n36630, n36631, n36632, n36633, n36634,
         n36635, n36636, n36637, n36638, n36639, n36640, n36641, n36642,
         n36643, n36644, n36645, n36646, n36647, n36648, n36649, n36650,
         n36651, n36652, n36653, n36654, n36655, n36656, n36657, n36658,
         n36659, n36660, n36661, n36662, n36663, n36664, n36665, n36666,
         n36667, n36668, n36669, n36670, n36671, n36672, n36673, n36674,
         n36675, n36676, n36677, n36678, n36679, n36680, n36681, n36682,
         n36683, n36684, n36685, n36686, n36687, n36688, n36689, n36690,
         n36691, n36692, n36693, n36694, n36695, n36696, n36697, n36698,
         n36699, n36700, n36701, n36702, n36703, n36704, n36705, n36706,
         n36707, n36708, n36709, n36710, n36711, n36712, n36713, n36714,
         n36715, n36716, n36717, n36718, n36719, n36720, n36721, n36722,
         n36723, n36724, n36725, n36726, n36727, n36728, n36729, n36730,
         n36731, n36732, n36733, n36734, n36735, n36736, n36737, n36738,
         n36739, n36740, n36741, n36742, n36743, n36744, n36745, n36746,
         n36747, n36748, n36749, n36750, n36751, n36752, n36753, n36754,
         n36755, n36756, n36757, n36758, n36759, n36760, n36761, n36762,
         n36763, n36764, n36765, n36766, n36767, n36768, n36769, n36770,
         n36771, n36772, n36773, n36774, n36775, n36776, n36777, n36778,
         n36779, n36780, n36781, n36782, n36783, n36784, n36785, n36786,
         n36787, n36788, n36789, n36790, n36791, n36792, n36793, n36794,
         n36795, n36796, n36797, n36798, n36799, n36800, n36801, n36802,
         n36803, n36804, n36805, n36806, n36807, n36808, n36809, n36810,
         n36811, n36812, n36813, n36814, n36815, n36816, n36817, n36818,
         n36819, n36820, n36821, n36822, n36823, n36824, n36825, n36826,
         n36827, n36828, n36829, n36830, n36831, n36832, n36833, n36834,
         n36835, n36836, n36837, n36838, n36839, n36840, n36841, n36842,
         n36843, n36844, n36845, n36846, n36847, n36848, n36849, n36850,
         n36851, n36852, n36853, n36854, n36855, n36856, n36857, n36858,
         n36859, n36860, n36861, n36862, n36863, n36864, n36865, n36866,
         n36867, n36868, n36869, n36870, n36871, n36872, n36873, n36874,
         n36875, n36876, n36877, n36878, n36879, n36880, n36881, n36882,
         n36883, n36884, n36885, n36886, n36887, n36888, n36889, n36890,
         n36891, n36892, n36893, n36894, n36895, n36896, n36897, n36898,
         n36899, n36900, n36901, n36902, n36903, n36904, n36905, n36906,
         n36907, n36908, n36909, n36910, n36911, n36912, n36913, n36914,
         n36915, n36916, n36917, n36918, n36919, n36920, n36921, n36922,
         n36923, n36924, n36925, n36926, n36927, n36928, n36929, n36930,
         n36931, n36932, n36933, n36934, n36935, n36936, n36937, n36938,
         n36939, n36940, n36941, n36942, n36943, n36944, n36945, n36946,
         n36947, n36948, n36949, n36950, n36951, n36952, n36953, n36954,
         n36955, n36956, n36957, n36958, n36959, n36960, n36961, n36962,
         n36963, n36964, n36965, n36966, n36967, n36968, n36969, n36970,
         n36971, n36972, n36973, n36974, n36975, n36976, n36977, n36978,
         n36979, n36980, n36981, n36982, n36983, n36984, n36985, n36986,
         n36987, n36988, n36989, n36990, n36991, n36992, n36993, n36994,
         n36995, n36996, n36997, n36998, n36999, n37000, n37001, n37002,
         n37003, n37004, n37005, n37006, n37007, n37008, n37009, n37010,
         n37011, n37012, n37013, n37014, n37015, n37016, n37017, n37018,
         n37019, n37020, n37021, n37022, n37023, n37024, n37025, n37026,
         n37027, n37028, n37029, n37030, n37031, n37032, n37033, n37034,
         n37035, n37036, n37037, n37038, n37039, n37040, n37041, n37042,
         n37043, n37044, n37045, n37046, n37047, n37048, n37049, n37050,
         n37051, n37052, n37053, n37054, n37055, n37056, n37057, n37058,
         n37059, n37060, n37061, n37062, n37063, n37064, n37065, n37066,
         n37067, n37068, n37069, n37070, n37071, n37072, n37073, n37074,
         n37075, n37076, n37077, n37078, n37079, n37080, n37081, n37082,
         n37083, n37084, n37085, n37086, n37087, n37088, n37089, n37090,
         n37091, n37092, n37093, n37094, n37095, n37096, n37097, n37098,
         n37099, n37100, n37101, n37102, n37103, n37104, n37105, n37106,
         n37107, n37108, n37109, n37110, n37111, n37112, n37113, n37114,
         n37115, n37116, n37117, n37118, n37119, n37120, n37121, n37122,
         n37123, n37124, n37125, n37126, n37127, n37128, n37129, n37130,
         n37131, n37132, n37133, n37134, n37135, n37136, n37137, n37138,
         n37139, n37140, n37141, n37142, n37143, n37144, n37145, n37146,
         n37147, n37148, n37149, n37150, n37151, n37152, n37153, n37154,
         n37155, n37156, n37157, n37158, n37159, n37160, n37161, n37162,
         n37163, n37164, n37165, n37166, n37167, n37168, n37169, n37170,
         n37171, n37172, n37173, n37174, n37175, n37176, n37177, n37178,
         n37179, n37180, n37181, n37182, n37183, n37184, n37185, n37186,
         n37187, n37188, n37189, n37190, n37191, n37192, n37193, n37194,
         n37195, n37196, n37197, n37198, n37199, n37200, n37201, n37202,
         n37203, n37204, n37205, n37206, n37207, n37208, n37209, n37210,
         n37211, n37212, n37213, n37214, n37215, n37216, n37217, n37218,
         n37219, n37220, n37221, n37222, n37223, n37224, n37225, n37226,
         n37227, n37228, n37229, n37230, n37231, n37232, n37233, n37234,
         n37235, n37236, n37237, n37238, n37239, n37240, n37241, n37242,
         n37243, n37244, n37245, n37246, n37247, n37248, n37249, n37250,
         n37251, n37252, n37253, n37254, n37255, n37256, n37257, n37258,
         n37259, n37260, n37261, n37262, n37263, n37264, n37265, n37266,
         n37267, n37268, n37269, n37270, n37271, n37272, n37273, n37274,
         n37275, n37276, n37277, n37278, n37279, n37280, n37281, n37282,
         n37283, n37284, n37285, n37286, n37287, n37288, n37289, n37290,
         n37291, n37292, n37293, n37294, n37295, n37296, n37297, n37298,
         n37299, n37300, n37301, n37302, n37303, n37304, n37305, n37306,
         n37307, n37308, n37309, n37310, n37311, n37312, n37313, n37314,
         n37315, n37316, n37317, n37318, n37319, n37320, n37321, n37322,
         n37323, n37324, n37325, n37326, n37327, n37328, n37329, n37330,
         n37331, n37332, n37333, n37334, n37335, n37336, n37337, n37338,
         n37339, n37340, n37341, n37342, n37343, n37344, n37345, n37346,
         n37347, n37348, n37349, n37350, n37351, n37352, n37353, n37354,
         n37355, n37356, n37357, n37358, n37359, n37360, n37361, n37362,
         n37363, n37364, n37365, n37366, n37367, n37368, n37369, n37370,
         n37371, n37372, n37373, n37374, n37375, n37376, n37377, n37378,
         n37379, n37380, n37381, n37382, n37383, n37384, n37385, n37386,
         n37387, n37388, n37389, n37390, n37391, n37392, n37393, n37394,
         n37395, n37396, n37397, n37398, n37399, n37400, n37401, n37402,
         n37403, n37404, n37405, n37406, n37407, n37408, n37409, n37410,
         n37411, n37412, n37413, n37414, n37415, n37416, n37417, n37418,
         n37419, n37420, n37421, n37422, n37423, n37424, n37425, n37426,
         n37427, n37428, n37429, n37430, n37431, n37432, n37433, n37434,
         n37435, n37436, n37437, n37438, n37439, n37440, n37441, n37442,
         n37443, n37444, n37445, n37446, n37447, n37448, n37449, n37450,
         n37451, n37452, n37453, n37454, n37455, n37456, n37457, n37458,
         n37459, n37460, n37461, n37462, n37463, n37464, n37465, n37466,
         n37467, n37468, n37469, n37470, n37471, n37472, n37473, n37474,
         n37475, n37476, n37477, n37478, n37479, n37480, n37481, n37482,
         n37483, n37484, n37485, n37486, n37487, n37488, n37489, n37490,
         n37491, n37492, n37493, n37494, n37495, n37496, n37497, n37498,
         n37499, n37500, n37501, n37502, n37503, n37504, n37505, n37506,
         n37507, n37508, n37509, n37510, n37511, n37512, n37513, n37514,
         n37515, n37516, n37517, n37518, n37519, n37520, n37521, n37522,
         n37523, n37524, n37525, n37526, n37527, n37528, n37529, n37530,
         n37531, n37532, n37533, n37534, n37535, n37536, n37537, n37538,
         n37539, n37540, n37541, n37542, n37543, n37544, n37545, n37546,
         n37547, n37548, n37549, n37550, n37551, n37552, n37553, n37554,
         n37555, n37556, n37557, n37558, n37559, n37560, n37561, n37562,
         n37563, n37564, n37565, n37566, n37567, n37568, n37569, n37570,
         n37571, n37572, n37573, n37574, n37575, n37576, n37577, n37578,
         n37579, n37580, n37581, n37582, n37583, n37584, n37585, n37586,
         n37587, n37588, n37589, n37590, n37591, n37592, n37593, n37594,
         n37595, n37596, n37597, n37598, n37599, n37600, n37601, n37602,
         n37603, n37604, n37605, n37606, n37607, n37608, n37609, n37610,
         n37611, n37612, n37613, n37614, n37615, n37616, n37617, n37618,
         n37619, n37620, n37621, n37622, n37623, n37624, n37625, n37626,
         n37627, n37628, n37629, n37630, n37631, n37632, n37633, n37634,
         n37635, n37636, n37637, n37638, n37639, n37640, n37641, n37642,
         n37643, n37644, n37645, n37646, n37647, n37648, n37649, n37650,
         n37651, n37652, n37653, n37654, n37655, n37656, n37657, n37658,
         n37659, n37660, n37661, n37662, n37663, n37664, n37665, n37666,
         n37667, n37668, n37669, n37670, n37671, n37672, n37673, n37674,
         n37675, n37676, n37677, n37678, n37679, n37680, n37681, n37682,
         n37683, n37684, n37685, n37686, n37687, n37688, n37689, n37690,
         n37691, n37692, n37693, n37694, n37695, n37696, n37697, n37698,
         n37699, n37700, n37701, n37702, n37703, n37704, n37705, n37706,
         n37707, n37708, n37709, n37710, n37711, n37712, n37713, n37714,
         n37715, n37716, n37717, n37718, n37719, n37720, n37721, n37722,
         n37723, n37724, n37725, n37726, n37727, n37728, n37729, n37730,
         n37731, n37732, n37733, n37734, n37735, n37736, n37737, n37738,
         n37739, n37740, n37741, n37742, n37743, n37744, n37745, n37746,
         n37747, n37748, n37749, n37750, n37751, n37752, n37753, n37754,
         n37755, n37756, n37757, n37758, n37759, n37760, n37761, n37762,
         n37763, n37764, n37765, n37766, n37767, n37768, n37769, n37770,
         n37771, n37772, n37773, n37774, n37775, n37776, n37777, n37778,
         n37779, n37780, n37781, n37782, n37783, n37784, n37785, n37786,
         n37787, n37788, n37789, n37790, n37791, n37792, n37793, n37794,
         n37795, n37796, n37797, n37798, n37799, n37800, n37801, n37802,
         n37803, n37804, n37805, n37806, n37807, n37808, n37809, n37810,
         n37811, n37812, n37813, n37814, n37815, n37816, n37817, n37818,
         n37819, n37820, n37821, n37822, n37823, n37824, n37825, n37826,
         n37827, n37828, n37829, n37830, n37831, n37832, n37833, n37834,
         n37835, n37836, n37837, n37838, n37839, n37840, n37841, n37842,
         n37843, n37844, n37845, n37846, n37847, n37848, n37849, n37850,
         n37851, n37852, n37853, n37854, n37855, n37856, n37857, n37858,
         n37859, n37860, n37861, n37862, n37863, n37864, n37865, n37866,
         n37867, n37868, n37869, n37870, n37871, n37872, n37873, n37874,
         n37875, n37876, n37877, n37878, n37879, n37880, n37881, n37882,
         n37883, n37884, n37885, n37886, n37887, n37888, n37889, n37890,
         n37891, n37892, n37893, n37894, n37895, n37896, n37897, n37898,
         n37899, n37900, n37901, n37902, n37903, n37904, n37905, n37906,
         n37907, n37908, n37909, n37910, n37911, n37912, n37913, n37914,
         n37915, n37916, n37917, n37918, n37919, n37920, n37921, n37922,
         n37923, n37924, n37925, n37926, n37927, n37928, n37929, n37930,
         n37931, n37932, n37933, n37934, n37935, n37936, n37937, n37938,
         n37939, n37940, n37941, n37942, n37943, n37944, n37945, n37946,
         n37947, n37948, n37949, n37950, n37951, n37952, n37953, n37954,
         n37955, n37956, n37957, n37958, n37959, n37960, n37961, n37962,
         n37963, n37964, n37965, n37966, n37967, n37968, n37969, n37970,
         n37971, n37972, n37973, n37974, n37975, n37976, n37977, n37978,
         n37979, n37980, n37981, n37982, n37983, n37984, n37985, n37986,
         n37987, n37988, n37989, n37990, n37991, n37992, n37993, n37994,
         n37995, n37996, n37997, n37998, n37999, n38000, n38001, n38002,
         n38003, n38004, n38005, n38006, n38007, n38008, n38009, n38010,
         n38011, n38012, n38013, n38014, n38015, n38016, n38017, n38018,
         n38019, n38020, n38021, n38022, n38023, n38024, n38025, n38026,
         n38027, n38028, n38029, n38030, n38031, n38032, n38033, n38034,
         n38035, n38036, n38037, n38038, n38039, n38040, n38041, n38042,
         n38043, n38044, n38045, n38046, n38047, n38048, n38049, n38050,
         n38051, n38052, n38053, n38054, n38055, n38056, n38057, n38058,
         n38059, n38060, n38061, n38062, n38063, n38064, n38065, n38066,
         n38067, n38068, n38069, n38070, n38071, n38072, n38073, n38074,
         n38075, n38076, n38077, n38078, n38079, n38080, n38081, n38082,
         n38083, n38084, n38085, n38086, n38087, n38088, n38089, n38090,
         n38091, n38092, n38093, n38094, n38095, n38096, n38097, n38098,
         n38099, n38100, n38101, n38102, n38103, n38104, n38105, n38106,
         n38107, n38108, n38109, n38110, n38111, n38112, n38113, n38114,
         n38115, n38116, n38117, n38118, n38119, n38120, n38121, n38122,
         n38123, n38124, n38125, n38126, n38127, n38128, n38129, n38130,
         n38131, n38132, n38133, n38134, n38135, n38136, n38137, n38138,
         n38139, n38140, n38141, n38142, n38143, n38144, n38145, n38146,
         n38147, n38148, n38149, n38150, n38151, n38152, n38153, n38154,
         n38155, n38156, n38157, n38158, n38159, n38160, n38161, n38162,
         n38163, n38164, n38165, n38166, n38167, n38168, n38169, n38170,
         n38171, n38172, n38173, n38174, n38175, n38176, n38177, n38178,
         n38179, n38180, n38181, n38182, n38183, n38184, n38185, n38186,
         n38187, n38188, n38189, n38190, n38191, n38192, n38193, n38194,
         n38195, n38196, n38197, n38198, n38199, n38200, n38201, n38202,
         n38203, n38204, n38205, n38206, n38207, n38208, n38209, n38210,
         n38211, n38212, n38213, n38214, n38215, n38216, n38217, n38218,
         n38219, n38220, n38221, n38222, n38223, n38224, n38225, n38226,
         n38227, n38228, n38229, n38230, n38231, n38232, n38233, n38234,
         n38235, n38236, n38237, n38238, n38239, n38240, n38241, n38242,
         n38243, n38244, n38245, n38246, n38247, n38248, n38249, n38250,
         n38251, n38252, n38253, n38254, n38255, n38256, n38257, n38258,
         n38259, n38260, n38261, n38262, n38263, n38264, n38265, n38266,
         n38267, n38268, n38269, n38270, n38271, n38272, n38273, n38274,
         n38275, n38276, n38277, n38278, n38279, n38280, n38281, n38282,
         n38283, n38284, n38285, n38286, n38287, n38288, n38289, n38290,
         n38291, n38292, n38293, n38294, n38295, n38296, n38297, n38298,
         n38299, n38300, n38301, n38302, n38303, n38304, n38305, n38306,
         n38307, n38308, n38309, n38310, n38311, n38312, n38313, n38314,
         n38315, n38316, n38317, n38318, n38319, n38320, n38321, n38322,
         n38323, n38324, n38325, n38326, n38327, n38328, n38329, n38330,
         n38331, n38332, n38333, n38334, n38335, n38336, n38337, n38338,
         n38339, n38340, n38341, n38342, n38343, n38344, n38345, n38346,
         n38347, n38348, n38349, n38350, n38351, n38352, n38353, n38354,
         n38355, n38356, n38357, n38358, n38359, n38360, n38361, n38362,
         n38363, n38364, n38365, n38366, n38367, n38368, n38369, n38370,
         n38371, n38372, n38373, n38374, n38375, n38376, n38377, n38378,
         n38379, n38380, n38381, n38382, n38383, n38384, n38385, n38386,
         n38387, n38388, n38389, n38390, n38391, n38392, n38393, n38394,
         n38395, n38396, n38397, n38398, n38399, n38400, n38401, n38402,
         n38403, n38404, n38405, n38406, n38407, n38408, n38409, n38410,
         n38411, n38412, n38413, n38414, n38415, n38416, n38417, n38418,
         n38419, n38420, n38421, n38422, n38423, n38424, n38425, n38426,
         n38427, n38428, n38429, n38430, n38431, n38432, n38433, n38434,
         n38435, n38436, n38437, n38438, n38439, n38440, n38441, n38442,
         n38443, n38444, n38445, n38446, n38447, n38448, n38449, n38450,
         n38451, n38452, n38453, n38454, n38455, n38456, n38457, n38458,
         n38459, n38460, n38461, n38462, n38463, n38464, n38465, n38466,
         n38467, n38468, n38469, n38470, n38471, n38472, n38473, n38474,
         n38475, n38476, n38477, n38478, n38479, n38480, n38481, n38482,
         n38483, n38484, n38485, n38486, n38487, n38488, n38489, n38490,
         n38491, n38492, n38493, n38494, n38495, n38496, n38497, n38498,
         n38499, n38500, n38501, n38502, n38503, n38504, n38505, n38506,
         n38507, n38508, n38509, n38510, n38511, n38512, n38513, n38514,
         n38515, n38516, n38517, n38518, n38519, n38520, n38521, n38522,
         n38523, n38524, n38525, n38526, n38527, n38528, n38529, n38530,
         n38531, n38532, n38533, n38534, n38535, n38536, n38537, n38538,
         n38539, n38540, n38541, n38542, n38543, n38544, n38545, n38546,
         n38547, n38548, n38549, n38550, n38551, n38552, n38553, n38554,
         n38555, n38556, n38557, n38558, n38559, n38560, n38561, n38562,
         n38563, n38564, n38565, n38566, n38567, n38568, n38569, n38570,
         n38571, n38572, n38573, n38574, n38575, n38576, n38577, n38578,
         n38579, n38580, n38581, n38582, n38583, n38584, n38585, n38586,
         n38587, n38588, n38589, n38590, n38591, n38592, n38593, n38594,
         n38595, n38596, n38597, n38598, n38599, n38600, n38601, n38602,
         n38603, n38604, n38605, n38606, n38607, n38608, n38609, n38610,
         n38611, n38612, n38613, n38614, n38615, n38616, n38617, n38618,
         n38619, n38620, n38621, n38622, n38623, n38624, n38625, n38626,
         n38627, n38628, n38629, n38630, n38631, n38632, n38633, n38634,
         n38635, n38636, n38637, n38638, n38639, n38640, n38641, n38642,
         n38643, n38644, n38645, n38646, n38647, n38648, n38649, n38650,
         n38651, n38652, n38653, n38654, n38655, n38656, n38657, n38658,
         n38659, n38660, n38661, n38662, n38663, n38664, n38665, n38666,
         n38667, n38668, n38669, n38670, n38671, n38672, n38673, n38674,
         n38675, n38676, n38677, n38678, n38679, n38680, n38681, n38682,
         n38683, n38684, n38685, n38686, n38687, n38688, n38689, n38690,
         n38691, n38692, n38693, n38694, n38695, n38696, n38697, n38698,
         n38699, n38700, n38701, n38702, n38703, n38704, n38705, n38706,
         n38707, n38708, n38709, n38710, n38711, n38712, n38713, n38714,
         n38715, n38716, n38717, n38718, n38719, n38720, n38721, n38722,
         n38723, n38724, n38725, n38726, n38727, n38728, n38729, n38730,
         n38731, n38732, n38733, n38734, n38735, n38736, n38737, n38738,
         n38739, n38740, n38741, n38742, n38743, n38744, n38745, n38746,
         n38747, n38748, n38749, n38750, n38751, n38752, n38753, n38754,
         n38755, n38756, n38757, n38758, n38759, n38760, n38761, n38762,
         n38763, n38764, n38765, n38766, n38767, n38768, n38769, n38770,
         n38771, n38772, n38773, n38774, n38775, n38776, n38777, n38778,
         n38779, n38780, n38781, n38782, n38783, n38784, n38785, n38786,
         n38787, n38788, n38789, n38790, n38791, n38792, n38793, n38794,
         n38795, n38796, n38797, n38798, n38799, n38800, n38801, n38802,
         n38803, n38804, n38805, n38806, n38807, n38808, n38809, n38810,
         n38811, n38812, n38813, n38814, n38815, n38816, n38817, n38818,
         n38819, n38820, n38821, n38822, n38823, n38824, n38825, n38826,
         n38827, n38828, n38829, n38830, n38831, n38832, n38833, n38834,
         n38835, n38836, n38837, n38838, n38839, n38840, n38841, n38842,
         n38843, n38844, n38845, n38846, n38847, n38848, n38849, n38850,
         n38851, n38852, n38853, n38854, n38855, n38856, n38857, n38858,
         n38859, n38860, n38861, n38862, n38863, n38864, n38865, n38866,
         n38867, n38868, n38869, n38870, n38871, n38872, n38873, n38874,
         n38875, n38876, n38877, n38878, n38879, n38880, n38881, n38882,
         n38883, n38884, n38885, n38886, n38887, n38888, n38889, n38890,
         n38891, n38892, n38893, n38894, n38895, n38896, n38897, n38898,
         n38899, n38900, n38901, n38902, n38903, n38904, n38905, n38906,
         n38907, n38908, n38909, n38910, n38911, n38912, n38913, n38914,
         n38915, n38916, n38917, n38918, n38919, n38920, n38921, n38922,
         n38923, n38924, n38925, n38926, n38927, n38928, n38929, n38930,
         n38931, n38932, n38933, n38934, n38935, n38936, n38937, n38938,
         n38939, n38940, n38941, n38942, n38943, n38944, n38945, n38946,
         n38947, n38948, n38949, n38950, n38951, n38952, n38953, n38954,
         n38955, n38956, n38957, n38958, n38959, n38960, n38961, n38962,
         n38963, n38964, n38965, n38966, n38967, n38968, n38969, n38970,
         n38971, n38972, n38973, n38974, n38975, n38976, n38977, n38978,
         n38979, n38980, n38981, n38982, n38983, n38984, n38985, n38986,
         n38987, n38988, n38989, n38990, n38991, n38992, n38993, n38994,
         n38995, n38996, n38997, n38998, n38999, n39000, n39001, n39002,
         n39003, n39004, n39005, n39006, n39007, n39008, n39009, n39010,
         n39011, n39012, n39013, n39014, n39015, n39016, n39017, n39018,
         n39019, n39020, n39021, n39022, n39023, n39024, n39025, n39026,
         n39027, n39028, n39029, n39030, n39031, n39032, n39033, n39034,
         n39035, n39036, n39037, n39038, n39039, n39040, n39041, n39042,
         n39043, n39044, n39045, n39046, n39047, n39048, n39049, n39050,
         n39051, n39052, n39053, n39054, n39055, n39056, n39057, n39058,
         n39059, n39060, n39061, n39062, n39063, n39064, n39065, n39066,
         n39067, n39068, n39069, n39070, n39071, n39072, n39073, n39074,
         n39075, n39076, n39077, n39078, n39079, n39080, n39081, n39082,
         n39083, n39084, n39085, n39086, n39087, n39088, n39089, n39090,
         n39091, n39092, n39093, n39094, n39095, n39096, n39097, n39098,
         n39099, n39100, n39101, n39102, n39103, n39104, n39105, n39106,
         n39107, n39108, n39109, n39110, n39111, n39112, n39113, n39114,
         n39115, n39116, n39117, n39118, n39119, n39120, n39121, n39122,
         n39123, n39124, n39125, n39126, n39127, n39128, n39129, n39130,
         n39131, n39132, n39133, n39134, n39135, n39136, n39137, n39138,
         n39139, n39140, n39141, n39142, n39143, n39144, n39145, n39146,
         n39147, n39148, n39149, n39150, n39151, n39152, n39153, n39154,
         n39155, n39156, n39157, n39158, n39159, n39160, n39161, n39162,
         n39163, n39164, n39165, n39166, n39167, n39168, n39169, n39170,
         n39171, n39172, n39173, n39174, n39175, n39176, n39177, n39178,
         n39179, n39180, n39181, n39182, n39183, n39184, n39185, n39186,
         n39187, n39188, n39189, n39190, n39191, n39192, n39193, n39194,
         n39195, n39196, n39197, n39198, n39199, n39200, n39201, n39202,
         n39203, n39204, n39205, n39206, n39207, n39208, n39209, n39210,
         n39211, n39212, n39213, n39214, n39215, n39216, n39217, n39218,
         n39219, n39220, n39221, n39222, n39223, n39224, n39225, n39226,
         n39227, n39228, n39229, n39230, n39231, n39232, n39233, n39234,
         n39235, n39236, n39237, n39238, n39239, n39240, n39241, n39242,
         n39243, n39244, n39245, n39246, n39247, n39248, n39249, n39250,
         n39251, n39252, n39253, n39254, n39255, n39256, n39257, n39258,
         n39259, n39260, n39261, n39262, n39263, n39264, n39265, n39266,
         n39267, n39268, n39269, n39270, n39271, n39272, n39273, n39274,
         n39275, n39276, n39277, n39278, n39279, n39280, n39281, n39282,
         n39283, n39284, n39285, n39286, n39287, n39288, n39289, n39290,
         n39291, n39292, n39293, n39294, n39295, n39296, n39297, n39298,
         n39299, n39300, n39301, n39302, n39303, n39304, n39305, n39306,
         n39307, n39308, n39309, n39310, n39311, n39312, n39313, n39314,
         n39315, n39316, n39317, n39318, n39319, n39320, n39321, n39322,
         n39323, n39324, n39325, n39326, n39327, n39328, n39329, n39330,
         n39331, n39332, n39333, n39334, n39335, n39336, n39337, n39338,
         n39339, n39340, n39341, n39342, n39343, n39344, n39345, n39346,
         n39347, n39348, n39349, n39350, n39351, n39352, n39353, n39354,
         n39355, n39356, n39357, n39358, n39359, n39360, n39361, n39362,
         n39363, n39364, n39365, n39366, n39367, n39368, n39369, n39370,
         n39371, n39372, n39373, n39374, n39375, n39376, n39377, n39378,
         n39379, n39380, n39381, n39382, n39383, n39384, n39385, n39386,
         n39387, n39388, n39389, n39390, n39391, n39392, n39393, n39394,
         n39395, n39396, n39397, n39398, n39399, n39400, n39401, n39402,
         n39403, n39404, n39405, n39406, n39407, n39408, n39409, n39410,
         n39411, n39412, n39413, n39414, n39415, n39416, n39417, n39418,
         n39419, n39420, n39421, n39422, n39423, n39424, n39425, n39426,
         n39427, n39428, n39429, n39430, n39431, n39432, n39433, n39434,
         n39435, n39436, n39437, n39438, n39439, n39440, n39441, n39442,
         n39443, n39444, n39445, n39446, n39447, n39448, n39449, n39450,
         n39451, n39452, n39453, n39454, n39455, n39456, n39457, n39458,
         n39459, n39460, n39461, n39462, n39463, n39464, n39465, n39466,
         n39467, n39468, n39469, n39470, n39471, n39472, n39473, n39474,
         n39475, n39476, n39477, n39478, n39479, n39480, n39481, n39482,
         n39483, n39484, n39485, n39486, n39487, n39488, n39489, n39490,
         n39491, n39492, n39493, n39494, n39495, n39496, n39497, n39498,
         n39499, n39500, n39501, n39502, n39503, n39504, n39505, n39506,
         n39507, n39508, n39509, n39510, n39511, n39512, n39513, n39514,
         n39515, n39516, n39517, n39518, n39519, n39520, n39521, n39522,
         n39523, n39524, n39525, n39526, n39527, n39528, n39529, n39530,
         n39531, n39532, n39533, n39534, n39535, n39536, n39537, n39538,
         n39539, n39540, n39541, n39542, n39543, n39544, n39545, n39546,
         n39547, n39548, n39549, n39550, n39551, n39552, n39553, n39554,
         n39555, n39556, n39557, n39558, n39559, n39560, n39561, n39562,
         n39563, n39564, n39565, n39566, n39567, n39568, n39569, n39570,
         n39571, n39572, n39573, n39574, n39575, n39576, n39577, n39578,
         n39579, n39580, n39581, n39582, n39583, n39584, n39585, n39586,
         n39587, n39588, n39589, n39590, n39591, n39592, n39593, n39594,
         n39595, n39596, n39597, n39598, n39599, n39600, n39601, n39602,
         n39603, n39604, n39605, n39606, n39607, n39608, n39609, n39610,
         n39611, n39612, n39613, n39614, n39615, n39616, n39617, n39618,
         n39619, n39620, n39621, n39622, n39623, n39624, n39625, n39626,
         n39627, n39628, n39629, n39630, n39631, n39632, n39633, n39634,
         n39635, n39636, n39637, n39638, n39639, n39640, n39641, n39642,
         n39643, n39644, n39645, n39646, n39647, n39648, n39649, n39650,
         n39651, n39652, n39653, n39654, n39655, n39656, n39657, n39658,
         n39659, n39660, n39661, n39662, n39663, n39664, n39665, n39666,
         n39667, n39668, n39669, n39670, n39671, n39672, n39673, n39674,
         n39675, n39676, n39677, n39678, n39679, n39680, n39681, n39682,
         n39683, n39684, n39685, n39686, n39687, n39688, n39689, n39690,
         n39691, n39692, n39693, n39694, n39695, n39696, n39697, n39698,
         n39699, n39700, n39701, n39702, n39703, n39704, n39705, n39706,
         n39707, n39708, n39709, n39710, n39711, n39712, n39713, n39714,
         n39715, n39716, n39717, n39718, n39719, n39720, n39721, n39722,
         n39723, n39724, n39725, n39726, n39727, n39728, n39729, n39730,
         n39731, n39732, n39733, n39734, n39735, n39736, n39737, n39738,
         n39739, n39740, n39741, n39742, n39743, n39744, n39745, n39746,
         n39747, n39748, n39749, n39750, n39751, n39752, n39753, n39754,
         n39755, n39756, n39757, n39758, n39759, n39760, n39761, n39762,
         n39763, n39764, n39765, n39766, n39767, n39768, n39769, n39770,
         n39771, n39772, n39773, n39774, n39775, n39776, n39777, n39778,
         n39779, n39780, n39781, n39782, n39783, n39784, n39785, n39786,
         n39787, n39788, n39789, n39790, n39791, n39792, n39793, n39794,
         n39795, n39796, n39797, n39798, n39799, n39800, n39801, n39802,
         n39803, n39804, n39805, n39806, n39807, n39808, n39809, n39810,
         n39811, n39812, n39813, n39814, n39815, n39816, n39817, n39818,
         n39819, n39820, n39821, n39822, n39823, n39824, n39825, n39826,
         n39827, n39828, n39829, n39830, n39831, n39832, n39833, n39834,
         n39835, n39836, n39837, n39838, n39839, n39840, n39841, n39842,
         n39843, n39844, n39845, n39846, n39847, n39848, n39849, n39850,
         n39851, n39852, n39853, n39854, n39855, n39856, n39857, n39858,
         n39859, n39860, n39861, n39862, n39863, n39864, n39865, n39866,
         n39867, n39868, n39869, n39870, n39871, n39872, n39873, n39874,
         n39875, n39876, n39877, n39878, n39879, n39880, n39881, n39882,
         n39883, n39884, n39885, n39886, n39887, n39888, n39889, n39890,
         n39891, n39892, n39893, n39894, n39895, n39896, n39897, n39898,
         n39899, n39900, n39901, n39902, n39903, n39904, n39905, n39906,
         n39907, n39908, n39909, n39910, n39911, n39912, n39913, n39914,
         n39915, n39916, n39917, n39918, n39919, n39920, n39921, n39922,
         n39923, n39924, n39925, n39926, n39927, n39928, n39929, n39930,
         n39931, n39932, n39933, n39934, n39935, n39936, n39937, n39938,
         n39939, n39940, n39941, n39942, n39943, n39944, n39945, n39946,
         n39947, n39948, n39949, n39950, n39951, n39952, n39953, n39954,
         n39955, n39956, n39957, n39958, n39959, n39960, n39961, n39962,
         n39963, n39964, n39965, n39966, n39967, n39968, n39969, n39970,
         n39971, n39972, n39973, n39974, n39975, n39976, n39977, n39978,
         n39979, n39980, n39981, n39982, n39983, n39984, n39985, n39986,
         n39987, n39988, n39989, n39990, n39991, n39992, n39993, n39994,
         n39995, n39996, n39997, n39998, n39999, n40000, n40001, n40002,
         n40003, n40004, n40005, n40006, n40007, n40008, n40009, n40010,
         n40011, n40012, n40013, n40014, n40015, n40016, n40017, n40018,
         n40019, n40020, n40021, n40022, n40023, n40024, n40025, n40026,
         n40027, n40028, n40029, n40030, n40031, n40032, n40033, n40034,
         n40035, n40036, n40037, n40038, n40039, n40040, n40041, n40042,
         n40043, n40044, n40045, n40046, n40047, n40048, n40049, n40050,
         n40051, n40052, n40053, n40054, n40055, n40056, n40057, n40058,
         n40059, n40060, n40061, n40062, n40063, n40064, n40065, n40066,
         n40067, n40068, n40069, n40070, n40071, n40072, n40073, n40074,
         n40075, n40076, n40077, n40078, n40079, n40080, n40081, n40082,
         n40083, n40084, n40085, n40086, n40087, n40088, n40089, n40090,
         n40091, n40092, n40093, n40094, n40095, n40096, n40097, n40098,
         n40099, n40100, n40101, n40102, n40103, n40104, n40105, n40106,
         n40107, n40108, n40109, n40110, n40111, n40112, n40113, n40114,
         n40115, n40116, n40117, n40118, n40119, n40120, n40121, n40122,
         n40123, n40124, n40125, n40126, n40127, n40128, n40129, n40130,
         n40131, n40132, n40133, n40134, n40135, n40136, n40137, n40138,
         n40139, n40140, n40141, n40142, n40143, n40144, n40145, n40146,
         n40147, n40148, n40149, n40150, n40151, n40152, n40153, n40154,
         n40155, n40156, n40157, n40158, n40159, n40160, n40161, n40162,
         n40163, n40164, n40165, n40166, n40167, n40168, n40169, n40170,
         n40171, n40172, n40173, n40174, n40175, n40176, n40177, n40178,
         n40179, n40180, n40181, n40182, n40183, n40184, n40185, n40186,
         n40187, n40188, n40189, n40190, n40191, n40192, n40193, n40194,
         n40195, n40196, n40197, n40198, n40199, n40200, n40201, n40202,
         n40203, n40204, n40205, n40206, n40207, n40208, n40209, n40210,
         n40211, n40212, n40213, n40214, n40215, n40216, n40217, n40218,
         n40219, n40220, n40221, n40222, n40223, n40224, n40225, n40226,
         n40227, n40228, n40229, n40230, n40231, n40232, n40233, n40234,
         n40235, n40236, n40237, n40238, n40239, n40240, n40241, n40242,
         n40243, n40244, n40245, n40246, n40247, n40248, n40249, n40250,
         n40251, n40252, n40253, n40254, n40255, n40256, n40257, n40258,
         n40259, n40260, n40261, n40262, n40263, n40264, n40265, n40266,
         n40267, n40268, n40269, n40270, n40271, n40272, n40273, n40274,
         n40275, n40276, n40277, n40278, n40279, n40280, n40281, n40282,
         n40283, n40284, n40285, n40286, n40287, n40288, n40289, n40290,
         n40291, n40292, n40293, n40294, n40295, n40296, n40297, n40298,
         n40299, n40300, n40301, n40302, n40303, n40304, n40305, n40306,
         n40307, n40308, n40309, n40310, n40311, n40312, n40313, n40314,
         n40315, n40316, n40317, n40318, n40319, n40320, n40321, n40322,
         n40323, n40324, n40325, n40326, n40327, n40328, n40329, n40330,
         n40331, n40332, n40333, n40334, n40335, n40336, n40337, n40338,
         n40339, n40340, n40341, n40342, n40343, n40344, n40345, n40346,
         n40347, n40348, n40349, n40350, n40351, n40352, n40353, n40354,
         n40355, n40356, n40357, n40358, n40359, n40360, n40361, n40362,
         n40363, n40364, n40365, n40366, n40367, n40368, n40369, n40370,
         n40371, n40372, n40373, n40374, n40375, n40376, n40377, n40378,
         n40379, n40380, n40381, n40382, n40383, n40384, n40385, n40386,
         n40387, n40388, n40389, n40390, n40391, n40392, n40393, n40394,
         n40395, n40396, n40397, n40398, n40399, n40400, n40401, n40402,
         n40403, n40404, n40405, n40406, n40407, n40408, n40409, n40410,
         n40411, n40412, n40413, n40414, n40415, n40416, n40417, n40418,
         n40419, n40420, n40421, n40422, n40423, n40424, n40425, n40426,
         n40427, n40428, n40429, n40430, n40431, n40432, n40433, n40434,
         n40435, n40436, n40437, n40438, n40439, n40440, n40441, n40442,
         n40443, n40444, n40445, n40446, n40447, n40448, n40449, n40450,
         n40451, n40452, n40453, n40454, n40455, n40456, n40457, n40458,
         n40459, n40460, n40461, n40462, n40463, n40464, n40465, n40466,
         n40467, n40468, n40469, n40470, n40471, n40472, n40473, n40474,
         n40475, n40476, n40477, n40478, n40479, n40480, n40481, n40482,
         n40483, n40484, n40485, n40486, n40487, n40488, n40489, n40490,
         n40491, n40492, n40493, n40494, n40495, n40496, n40497, n40498,
         n40499, n40500, n40501, n40502, n40503, n40504, n40505, n40506,
         n40507, n40508, n40509, n40510, n40511, n40512, n40513, n40514,
         n40515, n40516, n40517, n40518, n40519, n40520, n40521, n40522,
         n40523, n40524, n40525, n40526, n40527, n40528, n40529, n40530,
         n40531, n40532, n40533, n40534, n40535, n40536, n40537, n40538,
         n40539, n40540, n40541, n40542, n40543, n40544, n40545, n40546,
         n40547, n40548, n40549, n40550, n40551, n40552, n40553, n40554,
         n40555, n40556, n40557, n40558, n40559, n40560, n40561, n40562,
         n40563, n40564, n40565, n40566, n40567, n40568, n40569, n40570,
         n40571, n40572, n40573, n40574, n40575, n40576, n40577, n40578,
         n40579, n40580, n40581, n40582, n40583, n40584, n40585, n40586,
         n40587, n40588, n40589, n40590, n40591, n40592, n40593, n40594,
         n40595, n40596, n40597, n40598, n40599, n40600, n40601, n40602,
         n40603, n40604, n40605, n40606, n40607, n40608, n40609, n40610,
         n40611, n40612, n40613, n40614, n40615, n40616, n40617, n40618,
         n40619, n40620, n40621, n40622, n40623, n40624, n40625, n40626,
         n40627, n40628, n40629, n40630, n40631, n40632, n40633, n40634,
         n40635, n40636, n40637, n40638, n40639, n40640, n40641, n40642,
         n40643, n40644, n40645, n40646, n40647, n40648, n40649, n40650,
         n40651, n40652, n40653, n40654, n40655, n40656, n40657, n40658,
         n40659, n40660, n40661, n40662, n40663, n40664, n40665, n40666,
         n40667, n40668, n40669, n40670, n40671, n40672, n40673, n40674,
         n40675, n40676, n40677, n40678, n40679, n40680, n40681, n40682,
         n40683, n40684, n40685, n40686, n40687, n40688, n40689, n40690,
         n40691, n40692, n40693, n40694, n40695, n40696, n40697, n40698,
         n40699, n40700, n40701, n40702, n40703, n40704, n40705, n40706,
         n40707, n40708, n40709, n40710, n40711, n40712, n40713, n40714,
         n40715, n40716, n40717, n40718, n40719, n40720, n40721, n40722,
         n40723, n40724, n40725, n40726, n40727, n40728, n40729, n40730,
         n40731, n40732, n40733, n40734, n40735, n40736, n40737, n40738,
         n40739, n40740, n40741, n40742, n40743, n40744, n40745, n40746,
         n40747, n40748, n40749, n40750, n40751, n40752, n40753, n40754,
         n40755, n40756, n40757, n40758, n40759, n40760, n40761, n40762,
         n40763, n40764, n40765, n40766, n40767, n40768, n40769, n40770,
         n40771, n40772, n40773, n40774, n40775, n40776, n40777, n40778,
         n40779, n40780, n40781, n40782, n40783, n40784, n40785, n40786,
         n40787, n40788, n40789, n40790, n40791, n40792, n40793, n40794,
         n40795, n40796, n40797, n40798, n40799, n40800, n40801, n40802,
         n40803, n40804, n40805, n40806, n40807, n40808, n40809, n40810,
         n40811, n40812, n40813, n40814, n40815, n40816, n40817, n40818,
         n40819, n40820, n40821, n40822, n40823, n40824, n40825, n40826,
         n40827, n40828, n40829, n40830, n40831, n40832, n40833, n40834,
         n40835, n40836, n40837, n40838, n40839, n40840, n40841, n40842,
         n40843, n40844, n40845, n40846, n40847, n40848, n40849, n40850,
         n40851, n40852, n40853, n40854, n40855, n40856, n40857, n40858,
         n40859, n40860, n40861, n40862, n40863, n40864, n40865, n40866,
         n40867, n40868, n40869, n40870, n40871, n40872, n40873, n40874,
         n40875, n40876, n40877, n40878, n40879, n40880, n40881, n40882,
         n40883, n40884, n40885, n40886, n40887, n40888, n40889, n40890,
         n40891, n40892, n40893, n40894, n40895, n40896, n40897, n40898,
         n40899, n40900, n40901, n40902, n40903, n40904, n40905, n40906,
         n40907, n40908, n40909, n40910, n40911, n40912, n40913, n40914,
         n40915, n40916, n40917, n40918, n40919, n40920, n40921, n40922,
         n40923, n40924, n40925, n40926, n40927, n40928, n40929, n40930,
         n40931, n40932, n40933, n40934, n40935, n40936, n40937, n40938,
         n40939, n40940, n40941, n40942, n40943, n40944, n40945, n40946,
         n40947, n40948, n40949, n40950, n40951, n40952, n40953, n40954,
         n40955, n40956, n40957, n40958, n40959, n40960, n40961, n40962,
         n40963, n40964, n40965, n40966, n40967, n40968, n40969, n40970,
         n40971, n40972, n40973, n40974, n40975, n40976, n40977, n40978,
         n40979, n40980, n40981, n40982, n40983, n40984, n40985, n40986,
         n40987, n40988, n40989, n40990, n40991, n40992, n40993, n40994,
         n40995, n40996, n40997, n40998, n40999, n41000, n41001, n41002,
         n41003, n41004, n41005, n41006, n41007, n41008, n41009, n41010,
         n41011, n41012, n41013, n41014, n41015, n41016, n41017, n41018,
         n41019, n41020, n41021, n41022, n41023, n41024, n41025, n41026,
         n41027, n41028, n41029, n41030, n41031, n41032, n41033, n41034,
         n41035, n41036, n41037, n41038, n41039, n41040, n41041, n41042,
         n41043, n41044, n41045, n41046, n41047, n41048, n41049, n41050,
         n41051, n41052, n41053, n41054, n41055, n41056, n41057, n41058,
         n41059, n41060, n41061, n41062, n41063, n41064, n41065, n41066,
         n41067, n41068, n41069, n41070, n41071, n41072, n41073, n41074,
         n41075, n41076, n41077, n41078, n41079, n41080, n41081, n41082,
         n41083, n41084, n41085, n41086, n41087, n41088, n41089, n41090,
         n41091, n41092, n41093, n41094, n41095, n41096, n41097, n41098,
         n41099, n41100, n41101, n41102, n41103, n41104, n41105, n41106,
         n41107, n41108, n41109, n41110, n41111, n41112, n41113, n41114,
         n41115, n41116, n41117, n41118, n41119, n41120, n41121, n41122,
         n41123, n41124, n41125, n41126, n41127, n41128, n41129, n41130,
         n41131, n41132, n41133, n41134, n41135, n41136, n41137, n41138,
         n41139, n41140, n41141, n41142, n41143, n41144, n41145, n41146,
         n41147, n41148, n41149, n41150, n41151, n41152, n41153, n41154,
         n41155, n41156, n41157, n41158, n41159, n41160, n41161, n41162,
         n41163, n41164, n41165, n41166, n41167, n41168, n41169, n41170,
         n41171, n41172, n41173, n41174, n41175, n41176, n41177, n41178,
         n41179, n41180, n41181, n41182, n41183, n41184, n41185, n41186,
         n41187, n41188, n41189, n41190, n41191, n41192, n41193, n41194,
         n41195, n41196, n41197, n41198, n41199, n41200, n41201, n41202,
         n41203, n41204, n41205, n41206, n41207, n41208, n41209, n41210,
         n41211, n41212, n41213, n41214, n41215, n41216, n41217, n41218,
         n41219, n41220, n41221, n41222, n41223, n41224, n41225, n41226,
         n41227, n41228, n41229, n41230, n41231, n41232, n41233, n41234,
         n41235, n41236, n41237, n41238, n41239, n41240, n41241, n41242,
         n41243, n41244, n41245, n41246, n41247, n41248, n41249, n41250,
         n41251, n41252, n41253, n41254, n41255, n41256, n41257, n41258,
         n41259, n41260, n41261, n41262, n41263, n41264, n41265, n41266,
         n41267, n41268, n41269, n41270, n41271, n41272, n41273, n41274,
         n41275, n41276, n41277, n41278, n41279, n41280, n41281, n41282,
         n41283, n41284, n41285, n41286, n41287, n41288, n41289, n41290,
         n41291, n41292, n41293, n41294, n41295, n41296, n41297, n41298,
         n41299, n41300, n41301, n41302, n41303, n41304, n41305, n41306,
         n41307, n41308, n41309, n41310, n41311, n41312, n41313, n41314,
         n41315, n41316, n41317, n41318, n41319, n41320, n41321, n41322,
         n41323, n41324, n41325, n41326, n41327, n41328, n41329, n41330,
         n41331, n41332, n41333, n41334, n41335, n41336, n41337, n41338,
         n41339, n41340, n41341, n41342, n41343, n41344, n41345, n41346,
         n41347, n41348, n41349, n41350, n41351, n41352, n41353, n41354,
         n41355, n41356, n41357, n41358, n41359, n41360, n41361, n41362,
         n41363, n41364, n41365, n41366, n41367, n41368, n41369, n41370,
         n41371, n41372, n41373, n41374, n41375, n41376, n41377, n41378,
         n41379, n41380, n41381, n41382, n41383, n41384, n41385, n41386,
         n41387, n41388, n41389, n41390, n41391, n41392, n41393, n41394,
         n41395, n41396, n41397, n41398, n41399, n41400, n41401, n41402,
         n41403, n41404, n41405, n41406, n41407, n41408, n41409, n41410,
         n41411, n41412, n41413, n41414, n41415, n41416, n41417, n41418,
         n41419, n41420, n41421, n41422, n41423, n41424, n41425, n41426,
         n41427, n41428, n41429, n41430, n41431, n41432, n41433, n41434,
         n41435, n41436, n41437, n41438, n41439, n41440, n41441, n41442,
         n41443, n41444, n41445, n41446, n41447, n41448, n41449, n41450,
         n41451, n41452, n41453, n41454, n41455, n41456, n41457, n41458,
         n41459, n41460, n41461, n41462, n41463, n41464, n41465, n41466,
         n41467, n41468, n41469, n41470, n41471, n41472, n41473, n41474,
         n41475, n41476, n41477, n41478, n41479, n41480, n41481, n41482,
         n41483, n41484, n41485, n41486, n41487, n41488, n41489, n41490,
         n41491, n41492, n41493, n41494, n41495, n41496, n41497, n41498,
         n41499, n41500, n41501, n41502, n41503, n41504, n41505, n41506,
         n41507, n41508, n41509, n41510, n41511, n41512, n41513, n41514,
         n41515, n41516, n41517, n41518, n41519, n41520, n41521, n41522,
         n41523, n41524, n41525, n41526, n41527, n41528, n41529, n41530,
         n41531, n41532, n41533, n41534, n41535, n41536, n41537, n41538,
         n41539, n41540, n41541, n41542, n41543, n41544, n41545, n41546,
         n41547, n41548, n41549, n41550, n41551, n41552, n41553, n41554,
         n41555, n41556, n41557, n41558, n41559, n41560, n41561, n41562,
         n41563, n41564, n41565, n41566, n41567, n41568, n41569, n41570,
         n41571, n41572, n41573, n41574, n41575, n41576, n41577, n41578,
         n41579, n41580, n41581, n41582, n41583, n41584, n41585, n41586,
         n41587, n41588, n41589, n41590, n41591, n41592, n41593, n41594,
         n41595, n41596, n41597, n41598, n41599, n41600, n41601, n41602,
         n41603, n41604, n41605, n41606, n41607, n41608, n41609, n41610,
         n41611, n41612, n41613, n41614, n41615, n41616, n41617, n41618,
         n41619, n41620, n41621, n41622, n41623, n41624, n41625, n41626,
         n41627, n41628, n41629, n41630, n41631, n41632, n41633, n41634,
         n41635, n41636, n41637, n41638, n41639, n41640, n41641, n41642,
         n41643, n41644, n41645, n41646, n41647, n41648, n41649, n41650,
         n41651, n41652, n41653, n41654, n41655, n41656, n41657, n41658,
         n41659, n41660, n41661, n41662, n41663, n41664, n41665, n41666,
         n41667, n41668, n41669, n41670, n41671, n41672, n41673, n41674,
         n41675, n41676, n41677, n41678, n41679, n41680, n41681, n41682,
         n41683, n41684, n41685, n41686, n41687, n41688, n41689, n41690,
         n41691, n41692, n41693, n41694, n41695, n41696, n41697, n41698,
         n41699, n41700, n41701, n41702, n41703, n41704, n41705, n41706,
         n41707, n41708, n41709, n41710, n41711, n41712, n41713, n41714,
         n41715, n41716, n41717, n41718, n41719, n41720, n41721, n41722,
         n41723, n41724, n41725, n41726, n41727, n41728, n41729, n41730,
         n41731, n41732, n41733, n41734, n41735, n41736, n41737, n41738,
         n41739, n41740, n41741, n41742, n41743, n41744, n41745, n41746,
         n41747, n41748, n41749, n41750, n41751, n41752, n41753, n41754,
         n41755, n41756, n41757, n41758, n41759, n41760, n41761, n41762,
         n41763, n41764, n41765, n41766, n41767, n41768, n41769, n41770,
         n41771, n41772, n41773, n41774, n41775, n41776, n41777, n41778,
         n41779, n41780, n41781, n41782, n41783, n41784, n41785, n41786,
         n41787, n41788, n41789, n41790, n41791, n41792, n41793, n41794,
         n41795, n41796, n41797, n41798, n41799, n41800, n41801, n41802,
         n41803, n41804, n41805, n41806, n41807, n41808, n41809, n41810,
         n41811, n41812, n41813, n41814, n41815, n41816, n41817, n41818,
         n41819, n41820, n41821, n41822, n41823, n41824, n41825, n41826,
         n41827, n41828, n41829, n41830, n41831, n41832, n41833, n41834,
         n41835, n41836, n41837, n41838, n41839, n41840, n41841, n41842,
         n41843, n41844, n41845, n41846, n41847, n41848, n41849, n41850,
         n41851, n41852, n41853, n41854, n41855, n41856, n41857, n41858,
         n41859, n41860, n41861, n41862, n41863, n41864, n41865, n41866,
         n41867, n41868, n41869, n41870, n41871, n41872, n41873, n41874,
         n41875, n41876, n41877, n41878, n41879, n41880, n41881, n41882,
         n41883, n41884, n41885, n41886, n41887, n41888, n41889, n41890,
         n41891, n41892, n41893, n41894, n41895, n41896, n41897, n41898,
         n41899, n41900, n41901, n41902, n41903, n41904, n41905, n41906,
         n41907, n41908, n41909, n41910, n41911, n41912, n41913, n41914,
         n41915, n41916, n41917, n41918, n41919, n41920, n41921, n41922,
         n41923, n41924, n41925, n41926, n41927, n41928, n41929, n41930,
         n41931, n41932, n41933, n41934, n41935, n41936, n41937, n41938,
         n41939, n41940, n41941, n41942, n41943, n41944, n41945, n41946,
         n41947, n41948, n41949, n41950, n41951, n41952, n41953, n41954,
         n41955, n41956, n41957, n41958, n41959, n41960, n41961, n41962,
         n41963, n41964, n41965, n41966, n41967, n41968, n41969, n41970,
         n41971, n41972, n41973, n41974, n41975, n41976, n41977, n41978,
         n41979, n41980, n41981, n41982, n41983, n41984, n41985, n41986,
         n41987, n41988, n41989, n41990, n41991, n41992, n41993, n41994,
         n41995, n41996, n41997, n41998, n41999, n42000, n42001, n42002,
         n42003, n42004, n42005, n42006, n42007, n42008, n42009, n42010,
         n42011, n42012, n42013, n42014, n42015, n42016, n42017, n42018,
         n42019, n42020, n42021, n42022, n42023, n42024, n42025, n42026,
         n42027, n42028, n42029, n42030, n42031, n42032, n42033, n42034,
         n42035, n42036, n42037, n42038, n42039, n42040, n42041, n42042,
         n42043, n42044, n42045, n42046, n42047, n42048, n42049, n42050,
         n42051, n42052, n42053, n42054, n42055, n42056, n42057, n42058,
         n42059, n42060, n42061, n42062, n42063, n42064, n42065, n42066,
         n42067, n42068, n42069, n42070, n42071, n42072, n42073, n42074,
         n42075, n42076, n42077, n42078, n42079, n42080, n42081, n42082,
         n42083, n42084, n42085, n42086, n42087, n42088, n42089, n42090,
         n42091, n42092, n42093, n42094, n42095, n42096, n42097, n42098,
         n42099, n42100, n42101, n42102, n42103, n42104, n42105, n42106,
         n42107, n42108, n42109, n42110, n42111, n42112, n42113, n42114,
         n42115, n42116, n42117, n42118, n42119, n42120, n42121, n42122,
         n42123, n42124, n42125, n42126, n42127, n42128, n42129, n42130,
         n42131, n42132, n42133, n42134, n42135, n42136, n42137, n42138,
         n42139, n42140, n42141, n42142, n42143, n42144, n42145, n42146,
         n42147, n42148, n42149, n42150, n42151, n42152, n42153, n42154,
         n42155, n42156, n42157, n42158, n42159, n42160, n42161, n42162,
         n42163, n42164, n42165, n42166, n42167, n42168, n42169, n42170,
         n42171, n42172, n42173, n42174, n42175, n42176, n42177, n42178,
         n42179, n42180, n42181, n42182, n42183, n42184, n42185, n42186,
         n42187, n42188, n42189, n42190, n42191, n42192, n42193, n42194,
         n42195, n42196, n42197, n42198, n42199, n42200, n42201, n42202,
         n42203, n42204, n42205, n42206, n42207, n42208, n42209, n42210,
         n42211, n42212, n42213, n42214, n42215, n42216, n42217, n42218,
         n42219, n42220, n42221, n42222, n42223, n42224, n42225, n42226,
         n42227, n42228, n42229, n42230, n42231, n42232, n42233, n42234,
         n42235, n42236, n42237, n42238, n42239, n42240, n42241, n42242,
         n42243, n42244, n42245, n42246, n42247, n42248, n42249, n42250,
         n42251, n42252, n42253, n42254, n42255, n42256, n42257, n42258,
         n42259, n42260, n42261, n42262, n42263, n42264, n42265, n42266,
         n42267, n42268, n42269, n42270, n42271, n42272, n42273, n42274,
         n42275, n42276, n42277, n42278, n42279, n42280, n42281, n42282,
         n42283, n42284, n42285, n42286, n42287, n42288, n42289, n42290,
         n42291, n42292, n42293, n42294, n42295, n42296, n42297, n42298,
         n42299, n42300, n42301, n42302, n42303, n42304, n42305, n42306,
         n42307, n42308, n42309, n42310, n42311, n42312, n42313, n42314,
         n42315, n42316, n42317, n42318, n42319, n42320, n42321, n42322,
         n42323, n42324, n42325, n42326, n42327, n42328, n42329, n42330,
         n42331, n42332, n42333, n42334, n42335, n42336, n42337, n42338,
         n42339, n42340, n42341, n42342, n42343, n42344, n42345, n42346,
         n42347, n42348, n42349, n42350, n42351, n42352, n42353, n42354,
         n42355, n42356, n42357, n42358, n42359, n42360, n42361, n42362,
         n42363, n42364, n42365, n42366, n42367, n42368, n42369, n42370,
         n42371, n42372, n42373, n42374, n42375, n42376, n42377, n42378,
         n42379, n42380, n42381, n42382, n42383, n42384, n42385, n42386,
         n42387, n42388, n42389, n42390, n42391, n42392, n42393, n42394,
         n42395, n42396, n42397, n42398, n42399, n42400, n42401, n42402,
         n42403, n42404, n42405, n42406, n42407, n42408, n42409, n42410,
         n42411, n42412, n42413, n42414, n42415, n42416, n42417, n42418,
         n42419, n42420, n42421, n42422, n42423, n42424, n42425, n42426,
         n42427, n42428, n42429, n42430, n42431, n42432, n42433, n42434,
         n42435, n42436, n42437, n42438, n42439, n42440, n42441, n42442,
         n42443, n42444, n42445, n42446, n42447, n42448, n42449, n42450,
         n42451, n42452, n42453, n42454, n42455, n42456, n42457, n42458,
         n42459, n42460, n42461, n42462, n42463, n42464, n42465, n42466,
         n42467, n42468, n42469, n42470, n42471, n42472, n42473, n42474,
         n42475, n42476, n42477, n42478, n42479, n42480, n42481, n42482,
         n42483, n42484, n42485, n42486, n42487, n42488, n42489, n42490,
         n42491, n42492, n42493, n42494, n42495, n42496, n42497, n42498,
         n42499, n42500, n42501, n42502, n42503, n42504, n42505, n42506,
         n42507, n42508, n42509, n42510, n42511, n42512, n42513, n42514,
         n42515, n42516, n42517, n42518, n42519, n42520, n42521, n42522,
         n42523, n42524, n42525, n42526, n42527, n42528, n42529, n42530,
         n42531, n42532, n42533, n42534, n42535, n42536, n42537, n42538,
         n42539, n42540, n42541, n42542, n42543, n42544, n42545, n42546,
         n42547, n42548, n42549, n42550, n42551, n42552, n42553, n42554,
         n42555, n42556, n42557, n42558, n42559, n42560, n42561, n42562,
         n42563, n42564, n42565, n42566, n42567, n42568, n42569, n42570,
         n42571, n42572, n42573, n42574, n42575, n42576, n42577, n42578,
         n42579, n42580, n42581, n42582, n42583, n42584, n42585, n42586,
         n42587, n42588, n42589, n42590, n42591, n42592, n42593, n42594,
         n42595, n42596, n42597, n42598, n42599, n42600, n42601, n42602,
         n42603, n42604, n42605, n42606, n42607, n42608, n42609, n42610,
         n42611, n42612, n42613, n42614, n42615, n42616, n42617, n42618,
         n42619, n42620, n42621, n42622, n42623, n42624, n42625, n42626,
         n42627, n42628, n42629, n42630, n42631, n42632, n42633, n42634,
         n42635, n42636, n42637, n42638, n42639, n42640, n42641, n42642,
         n42643, n42644, n42645, n42646, n42647, n42648, n42649, n42650,
         n42651, n42652, n42653, n42654, n42655, n42656, n42657, n42658,
         n42659, n42660, n42661, n42662, n42663, n42664, n42665, n42666,
         n42667, n42668, n42669, n42670, n42671, n42672, n42673, n42674,
         n42675, n42676, n42677, n42678, n42679, n42680, n42681, n42682,
         n42683, n42684, n42685, n42686, n42687, n42688, n42689, n42690,
         n42691, n42692, n42693, n42694, n42695, n42696, n42697, n42698,
         n42699, n42700, n42701, n42702, n42703, n42704, n42705, n42706,
         n42707, n42708, n42709, n42710, n42711, n42712, n42713, n42714,
         n42715, n42716, n42717, n42718, n42719, n42720, n42721, n42722,
         n42723, n42724, n42725, n42726, n42727, n42728, n42729, n42730,
         n42731, n42732, n42733, n42734, n42735, n42736, n42737, n42738,
         n42739, n42740, n42741, n42742, n42743, n42744, n42745, n42746,
         n42747, n42748, n42749, n42750, n42751, n42752, n42753, n42754,
         n42755, n42756, n42757, n42758, n42759, n42760, n42761, n42762,
         n42763, n42764, n42765, n42766, n42767, n42768, n42769, n42770,
         n42771, n42772, n42773, n42774, n42775, n42776, n42777, n42778,
         n42779, n42780, n42781, n42782, n42783, n42784, n42785, n42786,
         n42787, n42788, n42789, n42790, n42791, n42792, n42793, n42794,
         n42795, n42796, n42797, n42798, n42799, n42800, n42801, n42802,
         n42803, n42804, n42805, n42806, n42807, n42808, n42809, n42810,
         n42811, n42812, n42813, n42814, n42815, n42816, n42817, n42818,
         n42819, n42820, n42821, n42822, n42823, n42824, n42825, n42826,
         n42827, n42828, n42829, n42830, n42831, n42832, n42833, n42834,
         n42835, n42836, n42837, n42838, n42839, n42840, n42841, n42842,
         n42843, n42844, n42845, n42846, n42847, n42848, n42849, n42850,
         n42851, n42852, n42853, n42854, n42855, n42856, n42857, n42858,
         n42859, n42860, n42861, n42862, n42863, n42864, n42865, n42866,
         n42867, n42868, n42869, n42870, n42871, n42872, n42873, n42874,
         n42875, n42876, n42877, n42878, n42879, n42880, n42881, n42882,
         n42883, n42884, n42885, n42886, n42887, n42888, n42889, n42890,
         n42891, n42892, n42893, n42894, n42895, n42896, n42897, n42898,
         n42899, n42900, n42901, n42902, n42903, n42904, n42905, n42906,
         n42907, n42908, n42909, n42910, n42911, n42912, n42913, n42914,
         n42915, n42916, n42917, n42918, n42919, n42920, n42921, n42922,
         n42923, n42924, n42925, n42926, n42927, n42928, n42929, n42930,
         n42931, n42932, n42933, n42934, n42935, n42936, n42937, n42938,
         n42939, n42940, n42941, n42942, n42943, n42944, n42945, n42946,
         n42947, n42948, n42949, n42950, n42951, n42952, n42953, n42954,
         n42955, n42956, n42957, n42958, n42959, n42960, n42961, n42962,
         n42963, n42964, n42965, n42966, n42967, n42968, n42969, n42970,
         n42971, n42972, n42973, n42974, n42975, n42976, n42977, n42978,
         n42979, n42980, n42981, n42982, n42983, n42984, n42985, n42986,
         n42987, n42988, n42989, n42990, n42991, n42992, n42993, n42994,
         n42995, n42996, n42997, n42998, n42999, n43000, n43001, n43002,
         n43003, n43004, n43005, n43006, n43007, n43008, n43009, n43010,
         n43011, n43012, n43013, n43014, n43015, n43016, n43017, n43018,
         n43019, n43020, n43021, n43022, n43023, n43024, n43025, n43026,
         n43027, n43028, n43029, n43030, n43031, n43032, n43033, n43034,
         n43035, n43036, n43037, n43038, n43039, n43040, n43041, n43042,
         n43043, n43044, n43045, n43046, n43047, n43048, n43049, n43050,
         n43051, n43052, n43053, n43054, n43055, n43056, n43057, n43058,
         n43059, n43060, n43061, n43062, n43063, n43064, n43065, n43066,
         n43067, n43068, n43069, n43070, n43071, n43072, n43073, n43074,
         n43075, n43076, n43077, n43078, n43079, n43080, n43081, n43082,
         n43083, n43084, n43085, n43086, n43087, n43088, n43089, n43090,
         n43091, n43092, n43093, n43094, n43095, n43096, n43097, n43098,
         n43099, n43100, n43101, n43102, n43103, n43104, n43105, n43106,
         n43107, n43108, n43109, n43110, n43111, n43112, n43113, n43114,
         n43115, n43116, n43117, n43118, n43119, n43120, n43121, n43122,
         n43123, n43124, n43125, n43126, n43127, n43128, n43129, n43130,
         n43131, n43132, n43133, n43134, n43135, n43136, n43137, n43138,
         n43139, n43140, n43141, n43142, n43143, n43144, n43145, n43146,
         n43147, n43148, n43149, n43150, n43151, n43152, n43153, n43154,
         n43155, n43156, n43157, n43158, n43159, n43160, n43161, n43162,
         n43163, n43164, n43165, n43166, n43167, n43168, n43169, n43170,
         n43171, n43172, n43173, n43174, n43175, n43176, n43177, n43178,
         n43179, n43180, n43181, n43182, n43183, n43184, n43185, n43186,
         n43187, n43188, n43189, n43190, n43191, n43192, n43193, n43194,
         n43195, n43196, n43197, n43198, n43199, n43200, n43201, n43202,
         n43203, n43204, n43205, n43206, n43207, n43208, n43209, n43210,
         n43211, n43212, n43213, n43214, n43215, n43216, n43217, n43218,
         n43219, n43220, n43221, n43222, n43223, n43224, n43225, n43226,
         n43227, n43228, n43229, n43230, n43231, n43232, n43233, n43234,
         n43235, n43236, n43237, n43238, n43239, n43240, n43241, n43242,
         n43243, n43244, n43245, n43246, n43247, n43248, n43249, n43250,
         n43251, n43252, n43253, n43254, n43255, n43256, n43257, n43258,
         n43259, n43260, n43261, n43262, n43263, n43264, n43265, n43266,
         n43267, n43268, n43269, n43270, n43271, n43272, n43273, n43274,
         n43275, n43276, n43277, n43278, n43279, n43280, n43281, n43282,
         n43283, n43284, n43285, n43286, n43287, n43288, n43289, n43290,
         n43291, n43292, n43293, n43294, n43295, n43296, n43297, n43298,
         n43299, n43300, n43301, n43302, n43303, n43304, n43305, n43306,
         n43307, n43308, n43309, n43310, n43311, n43312, n43313, n43314,
         n43315, n43316, n43317, n43318, n43319, n43320, n43321, n43322,
         n43323, n43324, n43325, n43326, n43327, n43328, n43329, n43330,
         n43331, n43332, n43333, n43334, n43335, n43336, n43337, n43338,
         n43339, n43340, n43341, n43342, n43343, n43344, n43345, n43346,
         n43347, n43348, n43349, n43350, n43351, n43352, n43353, n43354,
         n43355, n43356, n43357, n43358, n43359, n43360, n43361, n43362,
         n43363, n43364, n43365, n43366, n43367, n43368, n43369, n43370,
         n43371, n43372, n43373, n43374, n43375, n43376, n43377, n43378,
         n43379, n43380, n43381, n43382, n43383, n43384, n43385, n43386,
         n43387, n43388, n43389, n43390, n43391, n43392, n43393, n43394,
         n43395, n43396, n43397, n43398, n43399, n43400, n43401, n43402,
         n43403, n43404, n43405, n43406, n43407, n43408, n43409, n43410,
         n43411, n43412, n43413, n43414, n43415, n43416, n43417, n43418,
         n43419, n43420, n43421, n43422, n43423, n43424, n43425, n43426,
         n43427, n43428, n43429, n43430, n43431, n43432, n43433, n43434,
         n43435, n43436, n43437, n43438, n43439, n43440, n43441, n43442,
         n43443, n43444, n43445, n43446, n43447, n43448, n43449, n43450,
         n43451, n43452, n43453, n43454, n43455, n43456, n43457, n43458,
         n43459, n43460, n43461, n43462, n43463, n43464, n43465, n43466,
         n43467, n43468, n43469, n43470, n43471, n43472, n43473, n43474,
         n43475, n43476, n43477, n43478, n43479, n43480, n43481, n43482,
         n43483, n43484, n43485, n43486, n43487, n43488, n43489, n43490,
         n43491, n43492, n43493, n43494, n43495, n43496, n43497, n43498,
         n43499, n43500, n43501, n43502, n43503, n43504, n43505, n43506,
         n43507, n43508, n43509, n43510, n43511, n43512, n43513, n43514,
         n43515, n43516, n43517, n43518, n43519, n43520, n43521, n43522,
         n43523, n43524, n43525, n43526, n43527, n43528, n43529, n43530,
         n43531, n43532, n43533, n43534, n43535, n43536, n43537, n43538,
         n43539, n43540, n43541, n43542, n43543, n43544, n43545, n43546,
         n43547, n43548, n43549, n43550, n43551, n43552, n43553, n43554,
         n43555, n43556, n43557, n43558, n43559, n43560, n43561, n43562,
         n43563, n43564, n43565, n43566, n43567, n43568, n43569, n43570,
         n43571, n43572, n43573, n43574, n43575, n43576, n43577, n43578,
         n43579, n43580, n43581, n43582, n43583, n43584, n43585, n43586,
         n43587, n43588, n43589, n43590, n43591, n43592, n43593, n43594,
         n43595, n43596, n43597, n43598, n43599, n43600, n43601, n43602,
         n43603, n43604, n43605, n43606, n43607, n43608, n43609, n43610,
         n43611, n43612, n43613, n43614, n43615, n43616, n43617, n43618,
         n43619, n43620, n43621, n43622, n43623, n43624, n43625, n43626,
         n43627, n43628, n43629, n43630, n43631, n43632, n43633, n43634,
         n43635, n43636, n43637, n43638, n43639, n43640, n43641, n43642,
         n43643, n43644, n43645, n43646, n43647, n43648, n43649, n43650,
         n43651, n43652, n43653, n43654, n43655, n43656, n43657, n43658,
         n43659, n43660, n43661, n43662, n43663, n43664, n43665, n43666,
         n43667, n43668, n43669, n43670, n43671, n43672, n43673, n43674,
         n43675, n43676, n43677, n43678, n43679, n43680, n43681, n43682,
         n43683, n43684, n43685, n43686, n43687, n43688, n43689, n43690,
         n43691, n43692, n43693, n43694, n43695, n43696, n43697, n43698,
         n43699, n43700, n43701, n43702, n43703, n43704, n43705, n43706,
         n43707, n43708, n43709, n43710, n43711, n43712, n43713, n43714,
         n43715, n43716, n43717, n43718, n43719, n43720, n43721, n43722,
         n43723, n43724, n43725, n43726, n43727, n43728, n43729, n43730,
         n43731, n43732, n43733, n43734, n43735, n43736, n43737, n43738,
         n43739, n43740, n43741, n43742, n43743, n43744, n43745, n43746,
         n43747, n43748, n43749, n43750, n43751, n43752, n43753, n43754,
         n43755, n43756, n43757, n43758, n43759, n43760, n43761, n43762,
         n43763, n43764, n43765, n43766, n43767, n43768, n43769, n43770,
         n43771, n43772, n43773, n43774, n43775, n43776, n43777, n43778,
         n43779, n43780, n43781, n43782, n43783, n43784, n43785, n43786,
         n43787, n43788, n43789, n43790, n43791, n43792, n43793, n43794,
         n43795, n43796, n43797, n43798, n43799, n43800, n43801, n43802,
         n43803, n43804, n43805, n43806, n43807, n43808, n43809, n43810,
         n43811, n43812, n43813, n43814, n43815, n43816, n43817, n43818,
         n43819, n43820, n43821, n43822, n43823, n43824, n43825, n43826,
         n43827, n43828, n43829, n43830, n43831, n43832, n43833, n43834,
         n43835, n43836, n43837, n43838, n43839, n43840, n43841, n43842,
         n43843, n43844, n43845, n43846, n43847, n43848, n43849, n43850,
         n43851, n43852, n43853, n43854, n43855, n43856, n43857, n43858,
         n43859, n43860, n43861, n43862, n43863, n43864, n43865, n43866,
         n43867, n43868, n43869, n43870, n43871, n43872, n43873, n43874,
         n43875, n43876, n43877, n43878, n43879, n43880, n43881, n43882,
         n43883, n43884, n43885, n43886, n43887, n43888, n43889, n43890,
         n43891, n43892, n43893, n43894, n43895, n43896, n43897, n43898,
         n43899, n43900, n43901, n43902, n43903, n43904, n43905, n43906,
         n43907, n43908, n43909, n43910, n43911, n43912, n43913, n43914,
         n43915, n43916, n43917, n43918, n43919, n43920, n43921, n43922,
         n43923, n43924, n43925, n43926, n43927, n43928, n43929, n43930,
         n43931, n43932, n43933, n43934, n43935, n43936, n43937, n43938,
         n43939, n43940, n43941, n43942, n43943, n43944, n43945, n43946,
         n43947, n43948, n43949, n43950, n43951, n43952, n43953, n43954,
         n43955, n43956, n43957, n43958, n43959, n43960, n43961, n43962,
         n43963, n43964, n43965, n43966, n43967, n43968, n43969, n43970,
         n43971, n43972, n43973, n43974, n43975, n43976, n43977, n43978,
         n43979, n43980, n43981, n43982, n43983, n43984, n43985, n43986,
         n43987, n43988, n43989, n43990, n43991, n43992, n43993, n43994,
         n43995, n43996, n43997, n43998, n43999, n44000, n44001, n44002,
         n44003, n44004, n44005, n44006, n44007, n44008, n44009, n44010,
         n44011, n44012, n44013, n44014, n44015, n44016, n44017, n44018,
         n44019, n44020, n44021, n44022, n44023, n44024, n44025, n44026,
         n44027, n44028, n44029, n44030, n44031, n44032, n44033, n44034,
         n44035, n44036, n44037, n44038, n44039, n44040, n44041, n44042,
         n44043, n44044, n44045, n44046, n44047, n44048, n44049, n44050,
         n44051, n44052, n44053, n44054, n44055, n44056, n44057, n44058,
         n44059, n44060, n44061, n44062, n44063, n44064, n44065, n44066,
         n44067, n44068, n44069, n44070, n44071, n44072, n44073, n44074,
         n44075, n44076, n44077, n44078, n44079, n44080, n44081, n44082,
         n44083, n44084, n44085, n44086, n44087, n44088, n44089, n44090,
         n44091, n44092, n44093, n44094, n44095, n44096, n44097, n44098,
         n44099, n44100, n44101, n44102, n44103, n44104, n44105, n44106,
         n44107, n44108, n44109, n44110, n44111, n44112, n44113, n44114,
         n44115, n44116, n44117, n44118, n44119, n44120, n44121, n44122,
         n44123, n44124, n44125, n44126, n44127, n44128, n44129, n44130,
         n44131, n44132, n44133, n44134, n44135, n44136, n44137, n44138,
         n44139, n44140, n44141, n44142, n44143, n44144, n44145, n44146,
         n44147, n44148, n44149, n44150, n44151, n44152, n44153, n44154,
         n44155, n44156, n44157, n44158, n44159, n44160, n44161, n44162,
         n44163, n44164, n44165, n44166, n44167, n44168, n44169, n44170,
         n44171, n44172, n44173, n44174, n44175, n44176, n44177, n44178,
         n44179, n44180, n44181, n44182, n44183, n44184, n44185, n44186,
         n44187, n44188, n44189, n44190, n44191, n44192, n44193, n44194,
         n44195, n44196, n44197, n44198, n44199, n44200, n44201, n44202,
         n44203, n44204, n44205, n44206, n44207, n44208, n44209, n44210,
         n44211, n44212, n44213, n44214, n44215, n44216, n44217, n44218,
         n44219, n44220, n44221, n44222, n44223, n44224, n44225, n44226,
         n44227, n44228, n44229, n44230, n44231, n44232, n44233, n44234,
         n44235, n44236, n44237, n44238, n44239, n44240, n44241, n44242,
         n44243, n44244, n44245, n44246, n44247, n44248, n44249, n44250,
         n44251, n44252, n44253, n44254, n44255, n44256, n44257, n44258,
         n44259, n44260, n44261, n44262, n44263, n44264, n44265, n44266,
         n44267, n44268, n44269, n44270, n44271, n44272, n44273, n44274,
         n44275, n44276, n44277, n44278, n44279, n44280, n44281, n44282,
         n44283, n44284, n44285, n44286, n44287, n44288, n44289, n44290,
         n44291, n44292, n44293, n44294, n44295, n44296, n44297, n44298,
         n44299, n44300, n44301, n44302, n44303, n44304, n44305, n44306,
         n44307, n44308, n44309, n44310, n44311, n44312, n44313, n44314,
         n44315, n44316, n44317, n44318, n44319, n44320, n44321, n44322,
         n44323, n44324, n44325, n44326, n44327, n44328, n44329, n44330,
         n44331, n44332, n44333, n44334, n44335, n44336, n44337, n44338,
         n44339, n44340, n44341, n44342, n44343, n44344, n44345, n44346,
         n44347, n44348, n44349, n44350, n44351, n44352, n44353, n44354,
         n44355, n44356, n44357, n44358, n44359, n44360, n44361, n44362,
         n44363, n44364, n44365, n44366, n44367, n44368, n44369, n44370,
         n44371, n44372, n44373, n44374, n44375, n44376, n44377, n44378,
         n44379, n44380, n44381, n44382, n44383, n44384, n44385, n44386,
         n44387, n44388, n44389, n44390, n44391, n44392, n44393, n44394,
         n44395, n44396, n44397, n44398, n44399, n44400, n44401, n44402,
         n44403, n44404, n44405, n44406, n44407, n44408, n44409, n44410,
         n44411, n44412, n44413, n44414, n44415, n44416, n44417, n44418,
         n44419, n44420, n44421, n44422, n44423, n44424, n44425, n44426,
         n44427, n44428, n44429, n44430, n44431, n44432, n44433, n44434,
         n44435, n44436, n44437, n44438, n44439, n44440, n44441, n44442,
         n44443, n44444, n44445, n44446, n44447, n44448, n44449, n44450,
         n44451, n44452, n44453, n44454, n44455, n44456, n44457, n44458,
         n44459, n44460, n44461, n44462, n44463, n44464, n44465, n44466,
         n44467, n44468, n44469, n44470, n44471, n44472, n44473, n44474,
         n44475, n44476, n44477, n44478, n44479, n44480, n44481, n44482,
         n44483, n44484, n44485, n44486, n44487, n44488, n44489, n44490,
         n44491, n44492, n44493, n44494, n44495, n44496, n44497, n44498,
         n44499, n44500, n44501, n44502, n44503, n44504, n44505, n44506,
         n44507, n44508, n44509, n44510, n44511, n44512, n44513, n44514,
         n44515, n44516, n44517, n44518, n44519, n44520, n44521, n44522,
         n44523, n44524, n44525, n44526, n44527, n44528, n44529, n44530,
         n44531, n44532, n44533, n44534, n44535, n44536, n44537, n44538,
         n44539, n44540, n44541, n44542, n44543, n44544, n44545, n44546,
         n44547, n44548, n44549, n44550, n44551, n44552, n44553, n44554,
         n44555, n44556, n44557, n44558, n44559, n44560, n44561, n44562,
         n44563, n44564, n44565, n44566, n44567, n44568, n44569, n44570,
         n44571, n44572, n44573, n44574, n44575, n44576, n44577, n44578,
         n44579, n44580, n44581, n44582, n44583, n44584, n44585, n44586,
         n44587, n44588, n44589, n44590, n44591, n44592, n44593, n44594,
         n44595, n44596, n44597, n44598, n44599, n44600, n44601, n44602,
         n44603, n44604, n44605, n44606, n44607, n44608, n44609, n44610,
         n44611, n44612, n44613, n44614, n44615, n44616, n44617, n44618,
         n44619, n44620, n44621, n44622, n44623, n44624, n44625, n44626,
         n44627, n44628, n44629, n44630, n44631, n44632, n44633, n44634,
         n44635, n44636, n44637, n44638, n44639, n44640, n44641, n44642,
         n44643, n44644, n44645, n44646, n44647, n44648, n44649, n44650,
         n44651, n44652, n44653, n44654, n44655, n44656, n44657, n44658,
         n44659, n44660, n44661, n44662, n44663, n44664, n44665, n44666,
         n44667, n44668, n44669, n44670, n44671, n44672, n44673, n44674,
         n44675, n44676, n44677, n44678, n44679, n44680, n44681, n44682,
         n44683, n44684, n44685, n44686, n44687, n44688, n44689, n44690,
         n44691, n44692, n44693, n44694, n44695, n44696, n44697, n44698,
         n44699, n44700, n44701, n44702, n44703, n44704, n44705, n44706,
         n44707, n44708, n44709, n44710, n44711, n44712, n44713, n44714,
         n44715, n44716, n44717, n44718, n44719, n44720, n44721, n44722,
         n44723, n44724, n44725, n44726, n44727, n44728, n44729, n44730,
         n44731, n44732, n44733, n44734, n44735, n44736, n44737, n44738,
         n44739, n44740, n44741, n44742, n44743, n44744, n44745, n44746,
         n44747, n44748, n44749, n44750, n44751, n44752, n44753, n44754,
         n44755, n44756, n44757, n44758, n44759, n44760, n44761, n44762,
         n44763, n44764, n44765, n44766, n44767, n44768, n44769, n44770,
         n44771, n44772, n44773, n44774, n44775, n44776, n44777, n44778,
         n44779, n44780, n44781, n44782, n44783, n44784, n44785, n44786,
         n44787, n44788, n44789, n44790, n44791, n44792, n44793, n44794,
         n44795, n44796, n44797, n44798, n44799, n44800, n44801, n44802,
         n44803, n44804, n44805, n44806, n44807, n44808, n44809, n44810,
         n44811, n44812, n44813, n44814, n44815, n44816, n44817, n44818,
         n44819, n44820, n44821, n44822, n44823, n44824, n44825, n44826,
         n44827, n44828, n44829, n44830, n44831, n44832, n44833, n44834,
         n44835, n44836, n44837, n44838, n44839, n44840, n44841, n44842,
         n44843, n44844, n44845, n44846, n44847, n44848, n44849, n44850,
         n44851, n44852, n44853, n44854, n44855, n44856, n44857, n44858,
         n44859, n44860, n44861, n44862, n44863, n44864, n44865, n44866,
         n44867, n44868, n44869, n44870, n44871, n44872, n44873, n44874,
         n44875, n44876, n44877, n44878, n44879, n44880, n44881, n44882,
         n44883, n44884, n44885, n44886, n44887, n44888, n44889, n44890,
         n44891, n44892, n44893, n44894, n44895, n44896, n44897, n44898,
         n44899, n44900, n44901, n44902, n44903, n44904, n44905, n44906,
         n44907, n44908, n44909, n44910, n44911, n44912, n44913, n44914,
         n44915, n44916, n44917, n44918, n44919, n44920, n44921, n44922,
         n44923, n44924, n44925, n44926, n44927, n44928, n44929, n44930,
         n44931, n44932, n44933, n44934, n44935, n44936, n44937, n44938,
         n44939, n44940, n44941, n44942, n44943, n44944, n44945, n44946,
         n44947, n44948, n44949, n44950, n44951, n44952, n44953, n44954,
         n44955, n44956, n44957, n44958, n44959, n44960, n44961, n44962,
         n44963, n44964, n44965, n44966, n44967, n44968, n44969, n44970,
         n44971, n44972, n44973, n44974, n44975, n44976, n44977, n44978,
         n44979, n44980, n44981, n44982, n44983, n44984, n44985, n44986,
         n44987, n44988, n44989, n44990, n44991, n44992, n44993, n44994,
         n44995, n44996, n44997, n44998, n44999, n45000, n45001, n45002,
         n45003, n45004, n45005, n45006, n45007, n45008, n45009, n45010,
         n45011, n45012, n45013, n45014, n45015, n45016, n45017, n45018,
         n45019, n45020, n45021, n45022, n45023, n45024, n45025, n45026,
         n45027, n45028, n45029, n45030, n45031, n45032, n45033, n45034,
         n45035, n45036, n45037, n45038, n45039, n45040, n45041, n45042,
         n45043, n45044, n45045, n45046, n45047, n45048, n45049, n45050,
         n45051, n45052, n45053, n45054, n45055, n45056, n45057, n45058,
         n45059, n45060, n45061, n45062, n45063, n45064, n45065, n45066,
         n45067, n45068, n45069, n45070, n45071, n45072, n45073, n45074,
         n45075, n45076, n45077, n45078, n45079, n45080, n45081, n45082,
         n45083, n45084, n45085, n45086, n45087, n45088, n45089, n45090,
         n45091, n45092, n45093, n45094, n45095, n45096, n45097, n45098,
         n45099, n45100, n45101, n45102, n45103, n45104, n45105, n45106,
         n45107, n45108, n45109, n45110, n45111, n45112, n45113, n45114,
         n45115, n45116, n45117, n45118, n45119, n45120, n45121, n45122,
         n45123, n45124, n45125, n45126, n45127, n45128, n45129, n45130,
         n45131, n45132, n45133, n45134, n45135, n45136, n45137, n45138,
         n45139, n45140, n45141, n45142, n45143, n45144, n45145, n45146,
         n45147, n45148, n45149, n45150, n45151, n45152, n45153, n45154,
         n45155, n45156, n45157, n45158, n45159, n45160, n45161, n45162,
         n45163, n45164, n45165, n45166, n45167, n45168, n45169, n45170,
         n45171, n45172, n45173, n45174, n45175, n45176, n45177, n45178,
         n45179, n45180, n45181, n45182, n45183, n45184, n45185, n45186,
         n45187, n45188, n45189, n45190, n45191, n45192, n45193, n45194,
         n45195, n45196, n45197, n45198, n45199, n45200, n45201, n45202,
         n45203, n45204, n45205, n45206, n45207, n45208, n45209, n45210,
         n45211, n45212, n45213, n45214, n45215, n45216, n45217, n45218,
         n45219, n45220, n45221, n45222, n45223, n45224, n45225, n45226,
         n45227, n45228, n45229, n45230, n45231, n45232, n45233, n45234,
         n45235, n45236, n45237, n45238, n45239, n45240, n45241, n45242,
         n45243, n45244, n45245, n45246, n45247, n45248, n45249, n45250,
         n45251, n45252, n45253, n45254, n45255, n45256, n45257, n45258,
         n45259, n45260, n45261, n45262, n45263, n45264, n45265, n45266,
         n45267, n45268, n45269, n45270, n45271, n45272, n45273, n45274,
         n45275, n45276, n45277, n45278, n45279, n45280, n45281, n45282,
         n45283, n45284, n45285, n45286, n45287, n45288, n45289, n45290,
         n45291, n45292, n45293, n45294, n45295, n45296, n45297, n45298,
         n45299, n45300, n45301, n45302, n45303, n45304, n45305, n45306,
         n45307, n45308, n45309, n45310, n45311, n45312, n45313, n45314,
         n45315, n45316, n45317, n45318, n45319, n45320, n45321, n45322,
         n45323, n45324, n45325, n45326, n45327, n45328, n45329, n45330,
         n45331, n45332, n45333, n45334, n45335, n45336, n45337, n45338,
         n45339, n45340, n45341, n45342, n45343, n45344, n45345, n45346,
         n45347, n45348, n45349, n45350, n45351, n45352, n45353, n45354,
         n45355, n45356, n45357, n45358, n45359, n45360, n45361, n45362,
         n45363, n45364, n45365, n45366, n45367, n45368, n45369, n45370,
         n45371, n45372, n45373, n45374, n45375, n45376, n45377, n45378,
         n45379, n45380, n45381, n45382, n45383, n45384, n45385, n45386,
         n45387, n45388, n45389, n45390, n45391, n45392, n45393, n45394,
         n45395, n45396, n45397, n45398, n45399, n45400, n45401, n45402,
         n45403, n45404, n45405, n45406, n45407, n45408, n45409, n45410,
         n45411, n45412, n45413, n45414, n45415, n45416, n45417, n45418,
         n45419, n45420, n45421, n45422, n45423, n45424, n45425, n45426,
         n45427, n45428, n45429, n45430, n45431, n45432, n45433, n45434,
         n45435, n45436, n45437, n45438, n45439, n45440, n45441, n45442,
         n45443, n45444, n45445, n45446, n45447, n45448, n45449, n45450,
         n45451, n45452, n45453, n45454, n45455, n45456, n45457, n45458,
         n45459, n45460, n45461, n45462, n45463, n45464, n45465, n45466,
         n45467, n45468, n45469, n45470, n45471, n45472, n45473, n45474,
         n45475, n45476, n45477, n45478, n45479, n45480, n45481, n45482,
         n45483, n45484, n45485, n45486, n45487, n45488, n45489, n45490,
         n45491, n45492, n45493, n45494, n45495, n45496, n45497, n45498,
         n45499, n45500, n45501, n45502, n45503, n45504, n45505, n45506,
         n45507, n45508, n45509, n45510, n45511, n45512, n45513, n45514,
         n45515, n45516, n45517, n45518, n45519, n45520, n45521, n45522,
         n45523, n45524, n45525, n45526, n45527, n45528, n45529, n45530,
         n45531, n45532, n45533, n45534, n45535, n45536, n45537, n45538,
         n45539, n45540, n45541, n45542, n45543, n45544, n45545, n45546,
         n45547, n45548, n45549, n45550, n45551, n45552, n45553, n45554,
         n45555, n45556, n45557, n45558, n45559, n45560, n45561, n45562,
         n45563, n45564, n45565, n45566, n45567, n45568, n45569, n45570,
         n45571, n45572, n45573, n45574, n45575, n45576, n45577, n45578,
         n45579, n45580, n45581, n45582, n45583, n45584, n45585, n45586,
         n45587, n45588, n45589, n45590, n45591, n45592, n45593, n45594,
         n45595, n45596, n45597, n45598, n45599, n45600, n45601, n45602,
         n45603, n45604, n45605, n45606, n45607, n45608, n45609, n45610,
         n45611, n45612, n45613, n45614, n45615, n45616, n45617, n45618,
         n45619, n45620, n45621, n45622, n45623, n45624, n45625, n45626,
         n45627, n45628, n45629, n45630, n45631, n45632, n45633, n45634,
         n45635, n45636, n45637, n45638, n45639, n45640, n45641, n45642,
         n45643, n45644, n45645, n45646, n45647, n45648, n45649, n45650,
         n45651, n45652, n45653, n45654, n45655, n45656, n45657, n45658,
         n45659, n45660, n45661, n45662, n45663, n45664, n45665, n45666,
         n45667, n45668, n45669, n45670, n45671, n45672, n45673, n45674,
         n45675, n45676, n45677, n45678, n45679, n45680, n45681, n45682,
         n45683, n45684, n45685, n45686, n45687, n45688, n45689, n45690,
         n45691, n45692, n45693, n45694, n45695, n45696, n45697, n45698,
         n45699, n45700, n45701, n45702, n45703, n45704, n45705, n45706,
         n45707, n45708, n45709, n45710, n45711, n45712, n45713, n45714,
         n45715, n45716, n45717, n45718, n45719, n45720, n45721, n45722,
         n45723, n45724, n45725, n45726, n45727, n45728, n45729, n45730,
         n45731, n45732, n45733, n45734, n45735, n45736, n45737, n45738,
         n45739, n45740, n45741, n45742, n45743, n45744, n45745, n45746,
         n45747, n45748, n45749, n45750, n45751, n45752, n45753, n45754,
         n45755, n45756, n45757, n45758, n45759, n45760, n45761, n45762,
         n45763, n45764, n45765, n45766, n45767, n45768, n45769, n45770,
         n45771, n45772, n45773, n45774, n45775, n45776, n45777, n45778,
         n45779, n45780, n45781, n45782, n45783, n45784, n45785, n45786,
         n45787, n45788, n45789, n45790, n45791, n45792, n45793, n45794,
         n45795, n45796, n45797, n45798, n45799, n45800, n45801, n45802,
         n45803, n45804, n45805, n45806, n45807, n45808, n45809, n45810,
         n45811, n45812, n45813, n45814, n45815, n45816, n45817, n45818,
         n45819, n45820, n45821, n45822, n45823, n45824, n45825, n45826,
         n45827, n45828, n45829, n45830, n45831, n45832, n45833, n45834,
         n45835, n45836, n45837, n45838, n45839, n45840, n45841, n45842,
         n45843, n45844, n45845, n45846, n45847, n45848, n45849, n45850,
         n45851, n45852, n45853, n45854, n45855, n45856, n45857, n45858,
         n45859, n45860, n45861, n45862, n45863, n45864, n45865, n45866,
         n45867, n45868, n45869, n45870, n45871, n45872, n45873, n45874,
         n45875, n45876, n45877, n45878, n45879, n45880, n45881, n45882,
         n45883, n45884, n45885, n45886, n45887, n45888, n45889, n45890,
         n45891, n45892, n45893, n45894, n45895, n45896, n45897, n45898,
         n45899, n45900, n45901, n45902, n45903, n45904, n45905, n45906,
         n45907, n45908, n45909, n45910, n45911, n45912, n45913, n45914,
         n45915, n45916, n45917, n45918, n45919, n45920, n45921, n45922,
         n45923, n45924, n45925, n45926, n45927, n45928, n45929, n45930,
         n45931, n45932, n45933, n45934, n45935, n45936, n45937, n45938,
         n45939, n45940, n45941, n45942, n45943, n45944, n45945, n45946,
         n45947, n45948, n45949, n45950, n45951, n45952, n45953, n45954,
         n45955, n45956, n45957, n45958, n45959, n45960, n45961, n45962,
         n45963, n45964, n45965, n45966, n45967, n45968, n45969, n45970,
         n45971, n45972, n45973, n45974, n45975, n45976, n45977, n45978,
         n45979, n45980, n45981, n45982, n45983, n45984, n45985, n45986,
         n45987, n45988, n45989, n45990, n45991, n45992, n45993, n45994,
         n45995, n45996, n45997, n45998, n45999, n46000, n46001, n46002,
         n46003, n46004, n46005, n46006, n46007, n46008, n46009, n46010,
         n46011, n46012, n46013, n46014, n46015, n46016, n46017, n46018,
         n46019, n46020, n46021, n46022, n46023, n46024, n46025, n46026,
         n46027, n46028, n46029, n46030, n46031, n46032, n46033, n46034,
         n46035, n46036, n46037, n46038, n46039, n46040, n46041, n46042,
         n46043, n46044, n46045, n46046, n46047, n46048, n46049, n46050,
         n46051, n46052, n46053, n46054, n46055, n46056, n46057, n46058,
         n46059, n46060, n46061, n46062, n46063, n46064, n46065, n46066,
         n46067, n46068, n46069, n46070, n46071, n46072, n46073, n46074,
         n46075, n46076, n46077, n46078, n46079, n46080, n46081, n46082,
         n46083, n46084, n46085, n46086, n46087, n46088, n46089, n46090,
         n46091, n46092, n46093, n46094, n46095, n46096, n46097, n46098,
         n46099, n46100, n46101, n46102, n46103, n46104, n46105, n46106,
         n46107, n46108, n46109, n46110, n46111, n46112, n46113, n46114,
         n46115, n46116, n46117, n46118, n46119, n46120, n46121, n46122,
         n46123, n46124, n46125, n46126, n46127, n46128, n46129, n46130,
         n46131, n46132, n46133, n46134, n46135, n46136, n46137, n46138,
         n46139, n46140, n46141, n46142, n46143, n46144, n46145, n46146,
         n46147, n46148, n46149, n46150, n46151, n46152, n46153, n46154,
         n46155, n46156, n46157, n46158, n46159, n46160, n46161, n46162,
         n46163, n46164, n46165, n46166, n46167, n46168, n46169, n46170,
         n46171, n46172, n46173, n46174, n46175, n46176, n46177, n46178,
         n46179, n46180, n46181, n46182, n46183, n46184, n46185, n46186,
         n46187, n46188, n46189, n46190, n46191, n46192, n46193, n46194,
         n46195, n46196, n46197, n46198, n46199, n46200, n46201, n46202,
         n46203, n46204, n46205, n46206, n46207, n46208, n46209, n46210,
         n46211, n46212, n46213, n46214, n46215, n46216, n46217, n46218,
         n46219, n46220, n46221, n46222, n46223, n46224, n46225, n46226,
         n46227, n46228, n46229, n46230, n46231, n46232, n46233, n46234,
         n46235, n46236, n46237, n46238, n46239, n46240, n46241, n46242,
         n46243, n46244, n46245, n46246, n46247, n46248, n46249, n46250,
         n46251, n46252, n46253, n46254, n46255, n46256, n46257, n46258,
         n46259, n46260, n46261, n46262, n46263, n46264, n46265, n46266,
         n46267, n46268, n46269, n46270, n46271, n46272, n46273, n46274,
         n46275, n46276, n46277, n46278, n46279, n46280, n46281, n46282,
         n46283, n46284, n46285, n46286, n46287, n46288, n46289, n46290,
         n46291, n46292, n46293, n46294, n46295, n46296, n46297, n46298,
         n46299, n46300, n46301, n46302, n46303, n46304, n46305, n46306,
         n46307, n46308, n46309, n46310, n46311, n46312, n46313, n46314,
         n46315, n46316, n46317, n46318, n46319, n46320, n46321, n46322,
         n46323, n46324, n46325, n46326, n46327, n46328, n46329, n46330,
         n46331, n46332, n46333, n46334, n46335, n46336, n46337, n46338,
         n46339, n46340, n46341, n46342, n46343, n46344, n46345, n46346,
         n46347, n46348, n46349, n46350, n46351, n46352, n46353, n46354,
         n46355, n46356, n46357, n46358, n46359, n46360, n46361, n46362,
         n46363, n46364, n46365, n46366, n46367, n46368, n46369, n46370,
         n46371, n46372, n46373, n46374, n46375, n46376, n46377, n46378,
         n46379, n46380, n46381, n46382, n46383, n46384, n46385, n46386,
         n46387, n46388, n46389, n46390, n46391, n46392, n46393, n46394,
         n46395, n46396, n46397, n46398, n46399, n46400, n46401, n46402,
         n46403, n46404, n46405, n46406, n46407, n46408, n46409, n46410,
         n46411, n46412, n46413, n46414, n46415, n46416, n46417, n46418,
         n46419, n46420, n46421, n46422, n46423, n46424, n46425, n46426,
         n46427, n46428, n46429, n46430, n46431, n46432, n46433, n46434,
         n46435, n46436, n46437, n46438, n46439, n46440, n46441, n46442,
         n46443, n46444, n46445, n46446, n46447, n46448, n46449, n46450,
         n46451, n46452, n46453, n46454, n46455, n46456, n46457, n46458,
         n46459, n46460, n46461, n46462, n46463, n46464, n46465, n46466,
         n46467, n46468, n46469, n46470, n46471, n46472, n46473, n46474,
         n46475, n46476, n46477, n46478, n46479, n46480, n46481, n46482,
         n46483, n46484, n46485, n46486, n46487, n46488, n46489, n46490,
         n46491, n46492, n46493, n46494, n46495, n46496, n46497, n46498,
         n46499, n46500, n46501, n46502, n46503, n46504, n46505, n46506,
         n46507, n46508, n46509, n46510, n46511, n46512, n46513, n46514,
         n46515, n46516, n46517, n46518, n46519, n46520, n46521, n46522,
         n46523, n46524, n46525, n46526, n46527, n46528, n46529, n46530,
         n46531, n46532, n46533, n46534, n46535, n46536, n46537, n46538,
         n46539, n46540, n46541, n46542, n46543, n46544, n46545, n46546,
         n46547, n46548, n46549, n46550, n46551, n46552, n46553, n46554,
         n46555, n46556, n46557, n46558, n46559, n46560, n46561, n46562,
         n46563, n46564, n46565, n46566, n46567, n46568, n46569, n46570,
         n46571, n46572, n46573, n46574, n46575, n46576, n46577, n46578,
         n46579, n46580, n46581, n46582, n46583, n46584, n46585, n46586,
         n46587, n46588, n46589, n46590, n46591, n46592, n46593, n46594,
         n46595, n46596, n46597, n46598, n46599, n46600, n46601, n46602,
         n46603, n46604, n46605, n46606, n46607, n46608, n46609, n46610,
         n46611, n46612, n46613, n46614, n46615, n46616, n46617, n46618,
         n46619, n46620, n46621, n46622, n46623, n46624, n46625, n46626,
         n46627, n46628, n46629, n46630, n46631, n46632, n46633, n46634,
         n46635, n46636, n46637, n46638, n46639, n46640, n46641, n46642,
         n46643, n46644, n46645, n46646, n46647, n46648, n46649, n46650,
         n46651, n46652, n46653, n46654, n46655, n46656, n46657, n46658,
         n46659, n46660, n46661, n46662, n46663, n46664, n46665, n46666,
         n46667, n46668, n46669, n46670, n46671, n46672, n46673, n46674,
         n46675, n46676, n46677, n46678, n46679, n46680, n46681, n46682,
         n46683, n46684, n46685, n46686, n46687, n46688, n46689, n46690,
         n46691, n46692, n46693, n46694, n46695, n46696, n46697, n46698,
         n46699, n46700, n46701, n46702, n46703, n46704, n46705, n46706,
         n46707, n46708, n46709, n46710, n46711, n46712, n46713, n46714,
         n46715, n46716, n46717, n46718, n46719, n46720, n46721, n46722,
         n46723, n46724, n46725, n46726, n46727, n46728, n46729, n46730,
         n46731, n46732, n46733, n46734, n46735, n46736, n46737, n46738,
         n46739, n46740, n46741, n46742, n46743, n46744, n46745, n46746,
         n46747, n46748, n46749, n46750, n46751, n46752, n46753, n46754,
         n46755, n46756, n46757, n46758, n46759, n46760, n46761, n46762,
         n46763, n46764, n46765, n46766, n46767, n46768, n46769, n46770,
         n46771, n46772, n46773, n46774, n46775, n46776, n46777, n46778,
         n46779, n46780, n46781, n46782, n46783, n46784, n46785, n46786,
         n46787, n46788, n46789, n46790, n46791, n46792, n46793, n46794,
         n46795, n46796, n46797, n46798, n46799, n46800, n46801, n46802,
         n46803, n46804, n46805, n46806, n46807, n46808, n46809, n46810,
         n46811, n46812, n46813, n46814, n46815, n46816, n46817, n46818,
         n46819, n46820, n46821, n46822, n46823, n46824, n46825, n46826,
         n46827, n46828, n46829, n46830, n46831, n46832, n46833, n46834,
         n46835, n46836, n46837, n46838, n46839, n46840, n46841, n46842,
         n46843, n46844, n46845, n46846, n46847, n46848, n46849, n46850,
         n46851, n46852, n46853, n46854, n46855, n46856, n46857, n46858,
         n46859, n46860, n46861, n46862, n46863, n46864, n46865, n46866,
         n46867, n46868, n46869, n46870, n46871, n46872, n46873, n46874,
         n46875, n46876, n46877, n46878, n46879, n46880, n46881, n46882,
         n46883, n46884, n46885, n46886, n46887, n46888, n46889, n46890,
         n46891, n46892, n46893, n46894, n46895, n46896, n46897, n46898,
         n46899, n46900, n46901, n46902, n46903, n46904, n46905, n46906,
         n46907, n46908, n46909, n46910, n46911, n46912, n46913, n46914,
         n46915, n46916, n46917, n46918, n46919, n46920, n46921, n46922,
         n46923, n46924, n46925, n46926, n46927, n46928, n46929, n46930,
         n46931, n46932, n46933, n46934, n46935, n46936, n46937, n46938,
         n46939, n46940, n46941, n46942, n46943, n46944, n46945, n46946,
         n46947, n46948, n46949, n46950, n46951, n46952, n46953, n46954,
         n46955, n46956, n46957, n46958, n46959, n46960, n46961, n46962,
         n46963, n46964, n46965, n46966, n46967, n46968, n46969, n46970,
         n46971, n46972, n46973, n46974, n46975, n46976, n46977, n46978,
         n46979, n46980, n46981, n46982, n46983, n46984, n46985, n46986,
         n46987, n46988, n46989, n46990, n46991, n46992, n46993, n46994,
         n46995, n46996, n46997, n46998, n46999, n47000, n47001, n47002,
         n47003, n47004, n47005, n47006, n47007, n47008, n47009, n47010,
         n47011, n47012, n47013, n47014, n47015, n47016, n47017, n47018,
         n47019, n47020, n47021, n47022, n47023, n47024, n47025, n47026,
         n47027, n47028, n47029, n47030, n47031, n47032, n47033, n47034,
         n47035, n47036, n47037, n47038, n47039, n47040, n47041, n47042,
         n47043, n47044, n47045, n47046, n47047, n47048, n47049, n47050,
         n47051, n47052, n47053, n47054, n47055, n47056, n47057, n47058,
         n47059, n47060, n47061, n47062, n47063, n47064, n47065, n47066,
         n47067, n47068, n47069, n47070, n47071, n47072, n47073, n47074,
         n47075, n47076, n47077, n47078, n47079, n47080, n47081, n47082,
         n47083, n47084, n47085, n47086, n47087, n47088, n47089, n47090,
         n47091, n47092, n47093, n47094, n47095, n47096, n47097, n47098,
         n47099, n47100, n47101, n47102, n47103, n47104, n47105, n47106,
         n47107, n47108, n47109, n47110, n47111, n47112, n47113, n47114,
         n47115, n47116, n47117, n47118, n47119, n47120, n47121, n47122,
         n47123, n47124, n47125, n47126, n47127, n47128, n47129, n47130,
         n47131, n47132, n47133, n47134, n47135, n47136, n47137, n47138,
         n47139, n47140, n47141, n47142, n47143, n47144, n47145, n47146,
         n47147, n47148, n47149, n47150, n47151, n47152, n47153, n47154,
         n47155, n47156, n47157, n47158, n47159, n47160, n47161, n47162,
         n47163, n47164, n47165, n47166, n47167, n47168, n47169, n47170,
         n47171, n47172, n47173, n47174, n47175, n47176, n47177, n47178,
         n47179, n47180, n47181, n47182, n47183, n47184, n47185, n47186,
         n47187, n47188, n47189, n47190, n47191, n47192, n47193, n47194,
         n47195, n47196, n47197, n47198, n47199, n47200, n47201, n47202,
         n47203, n47204, n47205, n47206, n47207, n47208, n47209, n47210,
         n47211, n47212, n47213, n47214, n47215, n47216, n47217, n47218,
         n47219, n47220, n47221, n47222, n47223, n47224, n47225, n47226,
         n47227, n47228, n47229, n47230, n47231, n47232, n47233, n47234,
         n47235, n47236, n47237, n47238, n47239, n47240, n47241, n47242,
         n47243, n47244, n47245, n47246, n47247, n47248, n47249, n47250,
         n47251, n47252, n47253, n47254, n47255, n47256, n47257, n47258,
         n47259, n47260, n47261, n47262, n47263, n47264, n47265, n47266,
         n47267, n47268, n47269, n47270, n47271, n47272, n47273, n47274,
         n47275, n47276, n47277, n47278, n47279, n47280, n47281, n47282,
         n47283, n47284, n47285, n47286, n47287, n47288, n47289, n47290,
         n47291, n47292, n47293, n47294, n47295, n47296, n47297, n47298,
         n47299, n47300, n47301, n47302, n47303, n47304, n47305, n47306,
         n47307, n47308, n47309, n47310, n47311, n47312, n47313, n47314,
         n47315, n47316, n47317, n47318, n47319, n47320, n47321, n47322,
         n47323, n47324, n47325, n47326, n47327, n47328, n47329, n47330,
         n47331, n47332, n47333, n47334, n47335, n47336, n47337, n47338,
         n47339, n47340, n47341, n47342, n47343, n47344, n47345, n47346,
         n47347, n47348, n47349, n47350, n47351, n47352, n47353, n47354,
         n47355, n47356, n47357, n47358, n47359, n47360, n47361, n47362,
         n47363, n47364, n47365, n47366, n47367, n47368, n47369, n47370,
         n47371, n47372, n47373, n47374, n47375, n47376, n47377, n47378,
         n47379, n47380, n47381, n47382, n47383, n47384, n47385, n47386,
         n47387, n47388, n47389, n47390, n47391, n47392, n47393, n47394,
         n47395, n47396, n47397, n47398, n47399, n47400, n47401, n47402,
         n47403, n47404, n47405, n47406, n47407, n47408, n47409, n47410,
         n47411, n47412, n47413, n47414, n47415, n47416, n47417, n47418,
         n47419, n47420, n47421, n47422, n47423, n47424, n47425, n47426,
         n47427, n47428, n47429, n47430, n47431, n47432, n47433, n47434,
         n47435, n47436, n47437, n47438, n47439, n47440, n47441, n47442,
         n47443, n47444, n47445, n47446, n47447, n47448, n47449, n47450,
         n47451, n47452, n47453, n47454, n47455, n47456, n47457, n47458,
         n47459, n47460, n47461, n47462, n47463, n47464, n47465, n47466,
         n47467, n47468, n47469, n47470, n47471, n47472, n47473, n47474,
         n47475, n47476, n47477, n47478, n47479, n47480, n47481, n47482,
         n47483, n47484, n47485, n47486, n47487, n47488, n47489, n47490,
         n47491, n47492, n47493, n47494, n47495, n47496, n47497, n47498,
         n47499, n47500, n47501, n47502, n47503, n47504, n47505, n47506,
         n47507, n47508, n47509, n47510, n47511, n47512, n47513, n47514,
         n47515, n47516, n47517, n47518, n47519, n47520, n47521, n47522,
         n47523, n47524, n47525, n47526, n47527, n47528, n47529, n47530,
         n47531, n47532, n47533, n47534, n47535, n47536, n47537, n47538,
         n47539, n47540, n47541, n47542, n47543, n47544, n47545, n47546,
         n47547, n47548, n47549, n47550, n47551, n47552, n47553, n47554,
         n47555, n47556, n47557, n47558, n47559, n47560, n47561, n47562,
         n47563, n47564, n47565, n47566, n47567, n47568, n47569, n47570,
         n47571, n47572, n47573, n47574, n47575, n47576, n47577, n47578,
         n47579, n47580, n47581, n47582, n47583, n47584, n47585, n47586,
         n47587, n47588, n47589, n47590, n47591, n47592, n47593, n47594,
         n47595, n47596, n47597, n47598, n47599, n47600, n47601, n47602,
         n47603, n47604, n47605, n47606, n47607, n47608, n47609, n47610,
         n47611, n47612, n47613, n47614, n47615, n47616, n47617, n47618,
         n47619, n47620, n47621, n47622, n47623, n47624, n47625, n47626,
         n47627, n47628, n47629, n47630, n47631, n47632, n47633, n47634,
         n47635, n47636, n47637, n47638, n47639, n47640, n47641, n47642,
         n47643, n47644, n47645, n47646, n47647, n47648, n47649, n47650,
         n47651, n47652, n47653, n47654, n47655, n47656, n47657, n47658,
         n47659, n47660, n47661, n47662, n47663, n47664, n47665, n47666,
         n47667, n47668, n47669, n47670, n47671, n47672, n47673, n47674,
         n47675, n47676, n47677, n47678, n47679, n47680, n47681, n47682,
         n47683, n47684, n47685, n47686, n47687, n47688, n47689, n47690,
         n47691, n47692, n47693, n47694, n47695, n47696, n47697, n47698,
         n47699, n47700, n47701, n47702, n47703, n47704, n47705, n47706,
         n47707, n47708, n47709, n47710, n47711, n47712, n47713, n47714,
         n47715, n47716, n47717, n47718, n47719, n47720, n47721, n47722,
         n47723, n47724, n47725, n47726, n47727, n47728, n47729, n47730,
         n47731, n47732, n47733, n47734, n47735, n47736, n47737, n47738,
         n47739, n47740, n47741, n47742, n47743, n47744, n47745, n47746,
         n47747, n47748, n47749, n47750, n47751, n47752, n47753, n47754,
         n47755, n47756, n47757, n47758, n47759, n47760, n47761, n47762,
         n47763, n47764, n47765, n47766, n47767, n47768, n47769, n47770,
         n47771, n47772, n47773, n47774, n47775, n47776, n47777, n47778,
         n47779, n47780, n47781, n47782, n47783, n47784, n47785, n47786,
         n47787, n47788, n47789, n47790, n47791, n47792, n47793, n47794,
         n47795, n47796, n47797, n47798, n47799, n47800, n47801, n47802,
         n47803, n47804, n47805, n47806, n47807, n47808, n47809, n47810,
         n47811, n47812, n47813, n47814, n47815, n47816, n47817, n47818,
         n47819, n47820, n47821, n47822, n47823, n47824, n47825, n47826,
         n47827, n47828, n47829, n47830, n47831, n47832, n47833, n47834,
         n47835, n47836, n47837, n47838, n47839, n47840, n47841, n47842,
         n47843, n47844, n47845, n47846, n47847, n47848, n47849, n47850,
         n47851, n47852, n47853, n47854, n47855, n47856, n47857, n47858,
         n47859, n47860, n47861, n47862, n47863, n47864, n47865, n47866,
         n47867, n47868, n47869, n47870, n47871, n47872, n47873, n47874,
         n47875, n47876, n47877, n47878, n47879, n47880, n47881, n47882,
         n47883, n47884, n47885, n47886, n47887, n47888, n47889, n47890,
         n47891, n47892, n47893, n47894, n47895, n47896, n47897, n47898,
         n47899, n47900, n47901, n47902, n47903, n47904, n47905, n47906,
         n47907, n47908, n47909, n47910, n47911, n47912, n47913, n47914,
         n47915, n47916, n47917, n47918, n47919, n47920, n47921, n47922,
         n47923, n47924, n47925, n47926, n47927, n47928, n47929, n47930,
         n47931, n47932, n47933, n47934, n47935, n47936, n47937, n47938,
         n47939, n47940, n47941, n47942, n47943, n47944, n47945, n47946,
         n47947, n47948, n47949, n47950, n47951, n47952, n47953, n47954,
         n47955, n47956, n47957, n47958, n47959, n47960, n47961, n47962,
         n47963, n47964, n47965, n47966, n47967, n47968, n47969, n47970,
         n47971, n47972, n47973, n47974, n47975, n47976, n47977, n47978,
         n47979, n47980, n47981, n47982, n47983, n47984, n47985, n47986,
         n47987, n47988, n47989, n47990, n47991, n47992, n47993, n47994,
         n47995, n47996, n47997, n47998, n47999, n48000, n48001, n48002,
         n48003, n48004, n48005, n48006, n48007, n48008, n48009, n48010,
         n48011, n48012, n48013, n48014, n48015, n48016, n48017, n48018,
         n48019, n48020, n48021, n48022, n48023, n48024, n48025, n48026,
         n48027, n48028, n48029, n48030, n48031, n48032, n48033, n48034,
         n48035, n48036, n48037, n48038, n48039, n48040, n48041, n48042,
         n48043, n48044, n48045, n48046, n48047, n48048, n48049, n48050,
         n48051, n48052, n48053, n48054, n48055, n48056, n48057, n48058,
         n48059, n48060, n48061, n48062, n48063, n48064, n48065, n48066,
         n48067, n48068, n48069, n48070, n48071, n48072, n48073, n48074,
         n48075, n48076, n48077, n48078, n48079, n48080, n48081, n48082,
         n48083, n48084, n48085, n48086, n48087, n48088, n48089, n48090,
         n48091, n48092, n48093, n48094, n48095, n48096, n48097, n48098,
         n48099, n48100, n48101, n48102, n48103, n48104, n48105, n48106,
         n48107, n48108, n48109, n48110, n48111, n48112, n48113, n48114,
         n48115, n48116, n48117, n48118, n48119, n48120, n48121, n48122,
         n48123, n48124, n48125, n48126, n48127, n48128, n48129, n48130,
         n48131, n48132, n48133, n48134, n48135, n48136, n48137, n48138,
         n48139, n48140, n48141, n48142, n48143, n48144, n48145, n48146,
         n48147, n48148, n48149, n48150, n48151, n48152, n48153, n48154,
         n48155, n48156, n48157, n48158, n48159, n48160, n48161, n48162,
         n48163, n48164, n48165, n48166, n48167, n48168, n48169, n48170,
         n48171, n48172, n48173, n48174, n48175, n48176, n48177, n48178,
         n48179, n48180, n48181, n48182, n48183, n48184, n48185, n48186,
         n48187, n48188, n48189, n48190, n48191, n48192, n48193, n48194,
         n48195, n48196, n48197, n48198, n48199, n48200, n48201, n48202,
         n48203, n48204, n48205, n48206, n48207, n48208, n48209, n48210,
         n48211, n48212, n48213, n48214, n48215, n48216, n48217, n48218,
         n48219, n48220, n48221, n48222, n48223, n48224, n48225, n48226,
         n48227, n48228, n48229, n48230, n48231, n48232, n48233, n48234,
         n48235, n48236, n48237, n48238, n48239, n48240, n48241, n48242,
         n48243, n48244, n48245, n48246, n48247, n48248, n48249, n48250,
         n48251, n48252, n48253, n48254, n48255, n48256, n48257, n48258,
         n48259, n48260, n48261, n48262, n48263, n48264, n48265, n48266,
         n48267, n48268, n48269, n48270, n48271, n48272, n48273, n48274,
         n48275, n48276, n48277, n48278, n48279, n48280, n48281, n48282,
         n48283, n48284, n48285, n48286, n48287, n48288, n48289, n48290,
         n48291, n48292, n48293, n48294, n48295, n48296, n48297, n48298,
         n48299, n48300, n48301, n48302, n48303, n48304, n48305, n48306,
         n48307, n48308, n48309, n48310, n48311, n48312, n48313, n48314,
         n48315, n48316, n48317, n48318, n48319, n48320, n48321, n48322,
         n48323, n48324, n48325, n48326, n48327, n48328, n48329, n48330,
         n48331, n48332, n48333, n48334, n48335, n48336, n48337, n48338,
         n48339, n48340, n48341, n48342, n48343, n48344, n48345, n48346,
         n48347, n48348, n48349, n48350, n48351, n48352, n48353, n48354,
         n48355, n48356, n48357, n48358, n48359, n48360, n48361, n48362,
         n48363, n48364, n48365, n48366, n48367, n48368, n48369, n48370,
         n48371, n48372, n48373, n48374, n48375, n48376, n48377, n48378,
         n48379, n48380, n48381, n48382, n48383, n48384, n48385, n48386,
         n48387, n48388, n48389, n48390, n48391, n48392, n48393, n48394,
         n48395, n48396, n48397, n48398, n48399, n48400, n48401, n48402,
         n48403, n48404, n48405, n48406, n48407, n48408, n48409, n48410,
         n48411, n48412, n48413, n48414, n48415, n48416, n48417, n48418,
         n48419, n48420, n48421, n48422, n48423, n48424, n48425, n48426,
         n48427, n48428, n48429, n48430, n48431, n48432, n48433, n48434,
         n48435, n48436, n48437, n48438, n48439, n48440, n48441, n48442,
         n48443, n48444, n48445, n48446, n48447, n48448, n48449, n48450,
         n48451, n48452, n48453, n48454, n48455, n48456, n48457, n48458,
         n48459, n48460, n48461, n48462, n48463, n48464, n48465, n48466,
         n48467, n48468, n48469, n48470, n48471, n48472, n48473, n48474,
         n48475, n48476, n48477, n48478, n48479, n48480, n48481, n48482,
         n48483, n48484, n48485, n48486, n48487, n48488, n48489, n48490,
         n48491, n48492, n48493, n48494, n48495, n48496, n48497, n48498,
         n48499, n48500, n48501, n48502, n48503, n48504, n48505, n48506,
         n48507, n48508, n48509, n48510, n48511, n48512, n48513, n48514,
         n48515, n48516, n48517, n48518, n48519, n48520, n48521, n48522,
         n48523, n48524, n48525, n48526, n48527, n48528, n48529, n48530,
         n48531, n48532, n48533, n48534, n48535, n48536, n48537, n48538,
         n48539, n48540, n48541, n48542, n48543, n48544, n48545, n48546,
         n48547, n48548, n48549, n48550, n48551, n48552, n48553, n48554,
         n48555, n48556, n48557, n48558, n48559, n48560, n48561, n48562,
         n48563, n48564, n48565, n48566, n48567, n48568, n48569, n48570,
         n48571, n48572, n48573, n48574, n48575, n48576, n48577, n48578,
         n48579, n48580, n48581, n48582, n48583, n48584, n48585, n48586,
         n48587, n48588, n48589, n48590, n48591, n48592, n48593, n48594,
         n48595, n48596, n48597, n48598, n48599, n48600, n48601, n48602,
         n48603, n48604, n48605, n48606, n48607, n48608, n48609, n48610,
         n48611, n48612, n48613, n48614, n48615, n48616, n48617, n48618,
         n48619, n48620, n48621, n48622, n48623, n48624, n48625, n48626,
         n48627, n48628, n48629, n48630, n48631, n48632, n48633, n48634,
         n48635, n48636, n48637, n48638, n48639, n48640, n48641, n48642,
         n48643, n48644, n48645, n48646, n48647, n48648, n48649, n48650,
         n48651, n48652, n48653, n48654, n48655, n48656, n48657, n48658,
         n48659, n48660, n48661, n48662, n48663, n48664, n48665, n48666,
         n48667, n48668, n48669, n48670, n48671, n48672, n48673, n48674,
         n48675, n48676, n48677, n48678, n48679, n48680, n48681, n48682,
         n48683, n48684, n48685, n48686, n48687, n48688, n48689, n48690,
         n48691, n48692, n48693, n48694, n48695, n48696, n48697, n48698,
         n48699, n48700, n48701, n48702, n48703, n48704, n48705, n48706,
         n48707, n48708, n48709, n48710, n48711, n48712, n48713, n48714,
         n48715, n48716, n48717, n48718, n48719, n48720, n48721, n48722,
         n48723, n48724, n48725, n48726, n48727, n48728, n48729, n48730,
         n48731, n48732, n48733, n48734, n48735, n48736, n48737, n48738,
         n48739, n48740, n48741, n48742, n48743, n48744, n48745, n48746,
         n48747, n48748, n48749, n48750, n48751, n48752, n48753, n48754,
         n48755, n48756, n48757, n48758, n48759, n48760, n48761, n48762,
         n48763, n48764, n48765, n48766, n48767, n48768, n48769, n48770,
         n48771, n48772, n48773, n48774, n48775, n48776, n48777, n48778,
         n48779, n48780, n48781, n48782, n48783, n48784, n48785, n48786,
         n48787, n48788, n48789, n48790, n48791, n48792, n48793, n48794,
         n48795, n48796, n48797, n48798, n48799, n48800, n48801, n48802,
         n48803, n48804, n48805, n48806, n48807, n48808, n48809, n48810,
         n48811, n48812, n48813, n48814, n48815, n48816, n48817, n48818,
         n48819, n48820, n48821, n48822, n48823, n48824, n48825, n48826,
         n48827, n48828, n48829, n48830, n48831, n48832, n48833, n48834,
         n48835, n48836, n48837, n48838, n48839, n48840, n48841, n48842,
         n48843, n48844, n48845, n48846, n48847, n48848, n48849, n48850,
         n48851, n48852, n48853, n48854, n48855, n48856, n48857, n48858,
         n48859, n48860, n48861, n48862, n48863, n48864, n48865, n48866,
         n48867, n48868, n48869, n48870, n48871, n48872, n48873, n48874,
         n48875, n48876, n48877, n48878, n48879, n48880, n48881, n48882,
         n48883, n48884, n48885, n48886, n48887, n48888, n48889, n48890,
         n48891, n48892, n48893, n48894, n48895, n48896, n48897, n48898,
         n48899, n48900, n48901, n48902, n48903, n48904, n48905, n48906,
         n48907, n48908, n48909, n48910, n48911, n48912, n48913, n48914,
         n48915, n48916, n48917, n48918, n48919, n48920, n48921, n48922,
         n48923, n48924, n48925, n48926, n48927, n48928, n48929, n48930,
         n48931, n48932, n48933, n48934, n48935, n48936, n48937, n48938,
         n48939, n48940, n48941, n48942, n48943, n48944, n48945, n48946,
         n48947, n48948, n48949, n48950, n48951, n48952, n48953, n48954,
         n48955, n48956, n48957, n48958, n48959, n48960, n48961, n48962,
         n48963, n48964, n48965, n48966, n48967, n48968, n48969, n48970,
         n48971, n48972, n48973, n48974, n48975, n48976, n48977, n48978,
         n48979, n48980, n48981, n48982, n48983, n48984, n48985, n48986,
         n48987, n48988, n48989, n48990, n48991, n48992, n48993, n48994,
         n48995, n48996, n48997, n48998, n48999, n49000, n49001, n49002,
         n49003, n49004, n49005, n49006, n49007, n49008, n49009, n49010,
         n49011, n49012, n49013, n49014, n49015, n49016, n49017, n49018,
         n49019, n49020, n49021, n49022, n49023, n49024, n49025, n49026,
         n49027, n49028, n49029, n49030, n49031, n49032, n49033, n49034,
         n49035, n49036, n49037, n49038, n49039, n49040, n49041, n49042,
         n49043, n49044, n49045, n49046, n49047, n49048, n49049, n49050,
         n49051, n49052, n49053, n49054, n49055, n49056, n49057, n49058,
         n49059, n49060, n49061, n49062, n49063, n49064, n49065, n49066,
         n49067, n49068, n49069, n49070, n49071, n49072, n49073, n49074,
         n49075, n49076, n49077, n49078, n49079, n49080, n49081, n49082,
         n49083, n49084, n49085, n49086, n49087, n49088, n49089, n49090,
         n49091, n49092, n49093, n49094, n49095, n49096, n49097, n49098,
         n49099, n49100, n49101, n49102, n49103, n49104, n49105, n49106,
         n49107, n49108, n49109, n49110, n49111, n49112, n49113, n49114,
         n49115, n49116, n49117, n49118, n49119, n49120, n49121, n49122,
         n49123, n49124, n49125, n49126, n49127, n49128, n49129, n49130,
         n49131, n49132, n49133, n49134, n49135, n49136, n49137, n49138,
         n49139, n49140, n49141, n49142, n49143, n49144, n49145, n49146,
         n49147, n49148, n49149, n49150, n49151, n49152, n49153, n49154,
         n49155, n49156, n49157, n49158, n49159, n49160, n49161, n49162,
         n49163, n49164, n49165, n49166, n49167, n49168, n49169, n49170,
         n49171, n49172, n49173, n49174, n49175, n49176, n49177, n49178,
         n49179, n49180, n49181, n49182, n49183, n49184, n49185, n49186,
         n49187, n49188, n49189, n49190, n49191, n49192, n49193, n49194,
         n49195, n49196, n49197, n49198, n49199, n49200, n49201, n49202,
         n49203, n49204, n49205, n49206, n49207, n49208, n49209, n49210,
         n49211, n49212, n49213, n49214, n49215, n49216, n49217, n49218,
         n49219, n49220, n49221, n49222, n49223, n49224, n49225, n49226,
         n49227, n49228, n49229, n49230, n49231, n49232, n49233, n49234,
         n49235, n49236, n49237, n49238, n49239, n49240, n49241, n49242,
         n49243, n49244, n49245, n49246, n49247, n49248, n49249, n49250,
         n49251, n49252, n49253, n49254, n49255, n49256, n49257, n49258,
         n49259, n49260, n49261, n49262, n49263, n49264, n49265, n49266,
         n49267, n49268, n49269, n49270, n49271, n49272, n49273, n49274,
         n49275, n49276, n49277, n49278, n49279, n49280, n49281, n49282,
         n49283, n49284, n49285, n49286, n49287, n49288, n49289, n49290,
         n49291, n49292, n49293, n49294, n49295, n49296, n49297, n49298,
         n49299, n49300, n49301, n49302, n49303, n49304, n49305, n49306,
         n49307, n49308, n49309, n49310, n49311, n49312, n49313, n49314,
         n49315, n49316, n49317, n49318, n49319, n49320, n49321, n49322,
         n49323, n49324, n49325, n49326, n49327, n49328, n49329, n49330,
         n49331, n49332, n49333, n49334, n49335, n49336, n49337, n49338,
         n49339, n49340, n49341, n49342, n49343, n49344, n49345, n49346,
         n49347, n49348, n49349, n49350, n49351, n49352, n49353, n49354,
         n49355, n49356, n49357, n49358, n49359, n49360, n49361, n49362,
         n49363, n49364, n49365, n49366, n49367, n49368, n49369, n49370,
         n49371, n49372, n49373, n49374, n49375, n49376, n49377, n49378,
         n49379, n49380, n49381, n49382, n49383, n49384, n49385, n49386,
         n49387, n49388, n49389, n49390, n49391, n49392, n49393, n49394,
         n49395, n49396, n49397, n49398, n49399, n49400, n49401, n49402,
         n49403, n49404, n49405, n49406, n49407, n49408, n49409, n49410,
         n49411, n49412, n49413, n49414, n49415, n49416, n49417, n49418,
         n49419, n49420, n49421, n49422, n49423, n49424, n49425, n49426,
         n49427, n49428, n49429, n49430, n49431, n49432, n49433, n49434,
         n49435, n49436, n49437, n49438, n49439, n49440, n49441, n49442,
         n49443, n49444, n49445, n49446, n49447, n49448, n49449, n49450,
         n49451, n49452, n49453, n49454, n49455, n49456, n49457, n49458,
         n49459, n49460, n49461, n49462, n49463, n49464, n49465, n49466,
         n49467, n49468, n49469, n49470, n49471, n49472, n49473, n49474,
         n49475, n49476, n49477, n49478, n49479, n49480, n49481, n49482,
         n49483, n49484, n49485, n49486, n49487, n49488, n49489, n49490,
         n49491, n49492, n49493, n49494, n49495, n49496, n49497, n49498,
         n49499, n49500, n49501, n49502, n49503, n49504, n49505, n49506,
         n49507, n49508, n49509, n49510, n49511, n49512, n49513, n49514,
         n49515, n49516, n49517, n49518, n49519, n49520, n49521, n49522,
         n49523, n49524, n49525, n49526, n49527, n49528, n49529, n49530,
         n49531, n49532, n49533, n49534, n49535, n49536, n49537, n49538,
         n49539, n49540, n49541, n49542, n49543, n49544, n49545, n49546,
         n49547, n49548, n49549, n49550, n49551, n49552, n49553, n49554,
         n49555, n49556, n49557, n49558, n49559, n49560, n49561, n49562,
         n49563, n49564, n49565, n49566, n49567, n49568, n49569, n49570,
         n49571, n49572, n49573, n49574, n49575, n49576, n49577, n49578,
         n49579, n49580, n49581, n49582, n49583, n49584, n49585, n49586,
         n49587, n49588, n49589, n49590, n49591, n49592, n49593, n49594,
         n49595, n49596, n49597, n49598, n49599, n49600, n49601, n49602,
         n49603, n49604, n49605, n49606, n49607, n49608, n49609, n49610,
         n49611, n49612, n49613, n49614, n49615, n49616, n49617, n49618,
         n49619, n49620, n49621, n49622, n49623, n49624, n49625, n49626,
         n49627, n49628, n49629, n49630, n49631, n49632, n49633, n49634,
         n49635, n49636, n49637, n49638, n49639, n49640, n49641, n49642,
         n49643, n49644, n49645, n49646, n49647, n49648, n49649, n49650,
         n49651, n49652, n49653, n49654, n49655, n49656, n49657, n49658,
         n49659, n49660, n49661, n49662, n49663, n49664, n49665, n49666,
         n49667, n49668, n49669, n49670, n49671, n49672, n49673, n49674,
         n49675, n49676, n49677, n49678, n49679, n49680, n49681, n49682,
         n49683, n49684, n49685, n49686, n49687, n49688, n49689, n49690,
         n49691, n49692, n49693, n49694, n49695, n49696, n49697, n49698,
         n49699, n49700, n49701, n49702, n49703, n49704, n49705, n49706,
         n49707, n49708, n49709, n49710, n49711, n49712, n49713, n49714,
         n49715, n49716, n49717, n49718, n49719, n49720, n49721, n49722,
         n49723, n49724, n49725, n49726, n49727, n49728, n49729, n49730,
         n49731, n49732, n49733, n49734, n49735, n49736, n49737, n49738,
         n49739, n49740, n49741, n49742, n49743, n49744, n49745, n49746,
         n49747, n49748, n49749, n49750, n49751, n49752, n49753, n49754,
         n49755, n49756, n49757, n49758, n49759, n49760, n49761, n49762,
         n49763, n49764, n49765, n49766, n49767, n49768, n49769, n49770,
         n49771, n49772, n49773, n49774, n49775, n49776, n49777, n49778,
         n49779, n49780, n49781, n49782, n49783, n49784, n49785, n49786,
         n49787, n49788, n49789, n49790, n49791, n49792, n49793, n49794,
         n49795, n49796, n49797, n49798, n49799, n49800, n49801, n49802,
         n49803, n49804, n49805, n49806, n49807, n49808, n49809, n49810,
         n49811, n49812, n49813, n49814, n49815, n49816, n49817, n49818,
         n49819, n49820, n49821, n49822, n49823, n49824, n49825, n49826,
         n49827, n49828, n49829, n49830, n49831, n49832, n49833, n49834,
         n49835, n49836, n49837, n49838, n49839, n49840, n49841, n49842,
         n49843, n49844, n49845, n49846, n49847, n49848, n49849, n49850,
         n49851, n49852, n49853, n49854, n49855, n49856, n49857, n49858,
         n49859, n49860, n49861, n49862, n49863, n49864, n49865, n49866,
         n49867, n49868, n49869, n49870, n49871, n49872, n49873, n49874,
         n49875, n49876, n49877, n49878, n49879, n49880, n49881, n49882,
         n49883, n49884, n49885, n49886, n49887, n49888, n49889, n49890,
         n49891, n49892, n49893, n49894, n49895, n49896, n49897, n49898,
         n49899, n49900, n49901, n49902, n49903, n49904, n49905, n49906,
         n49907, n49908, n49909, n49910, n49911, n49912, n49913, n49914,
         n49915, n49916, n49917, n49918, n49919, n49920, n49921, n49922,
         n49923, n49924, n49925, n49926, n49927, n49928, n49929, n49930,
         n49931, n49932, n49933, n49934, n49935, n49936, n49937, n49938,
         n49939, n49940, n49941, n49942, n49943, n49944, n49945, n49946,
         n49947, n49948, n49949, n49950, n49951, n49952, n49953, n49954,
         n49955, n49956, n49957, n49958, n49959, n49960, n49961, n49962,
         n49963, n49964, n49965, n49966, n49967, n49968, n49969, n49970,
         n49971, n49972, n49973, n49974, n49975, n49976, n49977, n49978,
         n49979, n49980, n49981, n49982, n49983, n49984, n49985, n49986,
         n49987, n49988, n49989, n49990, n49991, n49992, n49993, n49994,
         n49995, n49996, n49997, n49998, n49999, n50000, n50001, n50002,
         n50003, n50004, n50005, n50006, n50007, n50008, n50009, n50010,
         n50011, n50012, n50013, n50014, n50015, n50016, n50017, n50018,
         n50019, n50020, n50021, n50022, n50023, n50024, n50025, n50026,
         n50027, n50028, n50029, n50030, n50031, n50032, n50033, n50034,
         n50035, n50036, n50037, n50038, n50039, n50040, n50041, n50042,
         n50043, n50044, n50045, n50046, n50047, n50048, n50049, n50050,
         n50051, n50052, n50053, n50054, n50055, n50056, n50057, n50058,
         n50059, n50060, n50061, n50062, n50063, n50064, n50065, n50066,
         n50067, n50068, n50069, n50070, n50071, n50072, n50073, n50074,
         n50075, n50076, n50077, n50078, n50079, n50080, n50081, n50082,
         n50083, n50084, n50085, n50086, n50087, n50088, n50089, n50090,
         n50091, n50092, n50093, n50094, n50095, n50096, n50097, n50098,
         n50099, n50100, n50101, n50102, n50103, n50104, n50105, n50106,
         n50107, n50108, n50109, n50110, n50111, n50112, n50113, n50114,
         n50115, n50116, n50117, n50118, n50119, n50120, n50121, n50122,
         n50123, n50124, n50125, n50126, n50127, n50128, n50129, n50130,
         n50131, n50132, n50133, n50134, n50135, n50136, n50137, n50138,
         n50139, n50140, n50141, n50142, n50143, n50144, n50145, n50146,
         n50147, n50148, n50149, n50150, n50151, n50152, n50153, n50154,
         n50155, n50156, n50157, n50158, n50159, n50160, n50161, n50162,
         n50163, n50164, n50165, n50166, n50167, n50168, n50169, n50170,
         n50171, n50172, n50173, n50174, n50175, n50176, n50177, n50178,
         n50179, n50180, n50181, n50182, n50183, n50184, n50185, n50186,
         n50187, n50188, n50189, n50190, n50191, n50192, n50193, n50194,
         n50195, n50196, n50197, n50198, n50199, n50200, n50201, n50202,
         n50203, n50204, n50205, n50206, n50207, n50208, n50209, n50210,
         n50211, n50212, n50213, n50214, n50215, n50216, n50217, n50218,
         n50219, n50220, n50221, n50222, n50223, n50224, n50225, n50226,
         n50227, n50228, n50229, n50230, n50231, n50232, n50233, n50234,
         n50235, n50236, n50237, n50238, n50239, n50240, n50241, n50242,
         n50243, n50244, n50245, n50246, n50247, n50248, n50249, n50250,
         n50251, n50252, n50253, n50254, n50255, n50256, n50257, n50258,
         n50259, n50260, n50261, n50262, n50263, n50264, n50265, n50266,
         n50267, n50268, n50269, n50270, n50271, n50272, n50273, n50274,
         n50275, n50276, n50277, n50278, n50279, n50280, n50281, n50282,
         n50283, n50284, n50285, n50286, n50287, n50288, n50289, n50290,
         n50291, n50292, n50293, n50294, n50295, n50296, n50297, n50298,
         n50299, n50300, n50301, n50302, n50303, n50304, n50305, n50306,
         n50307, n50308, n50309, n50310, n50311, n50312, n50313, n50314,
         n50315, n50316, n50317, n50318, n50319, n50320, n50321, n50322,
         n50323, n50324, n50325, n50326, n50327, n50328, n50329, n50330,
         n50331, n50332, n50333, n50334, n50335, n50336, n50337, n50338,
         n50339, n50340, n50341, n50342, n50343, n50344, n50345, n50346,
         n50347, n50348, n50349, n50350, n50351, n50352, n50353, n50354,
         n50355, n50356, n50357, n50358, n50359, n50360, n50361, n50362,
         n50363, n50364, n50365, n50366, n50367, n50368, n50369, n50370,
         n50371, n50372, n50373, n50374, n50375, n50376, n50377, n50378,
         n50379, n50380, n50381, n50382, n50383, n50384, n50385, n50386,
         n50387, n50388, n50389, n50390, n50391, n50392, n50393, n50394,
         n50395, n50396, n50397, n50398, n50399, n50400, n50401, n50402,
         n50403, n50404, n50405, n50406, n50407, n50408, n50409, n50410,
         n50411, n50412, n50413, n50414, n50415, n50416, n50417, n50418,
         n50419, n50420, n50421, n50422, n50423, n50424, n50425, n50426,
         n50427, n50428, n50429, n50430, n50431, n50432, n50433, n50434,
         n50435, n50436, n50437, n50438, n50439, n50440, n50441, n50442,
         n50443, n50444, n50445, n50446, n50447, n50448, n50449, n50450,
         n50451, n50452, n50453, n50454, n50455, n50456, n50457, n50458,
         n50459, n50460, n50461, n50462, n50463, n50464, n50465, n50466,
         n50467, n50468, n50469, n50470, n50471, n50472, n50473, n50474,
         n50475, n50476, n50477, n50478, n50479, n50480, n50481, n50482,
         n50483, n50484, n50485, n50486, n50487, n50488, n50489, n50490,
         n50491, n50492, n50493, n50494, n50495, n50496, n50497, n50498,
         n50499, n50500, n50501, n50502, n50503, n50504, n50505, n50506,
         n50507, n50508, n50509, n50510, n50511, n50512, n50513, n50514,
         n50515, n50516, n50517, n50518, n50519, n50520, n50521, n50522,
         n50523, n50524, n50525, n50526, n50527, n50528, n50529, n50530,
         n50531, n50532, n50533, n50534, n50535, n50536, n50537, n50538,
         n50539, n50540, n50541, n50542, n50543, n50544, n50545, n50546,
         n50547, n50548, n50549, n50550, n50551, n50552, n50553, n50554,
         n50555, n50556, n50557, n50558, n50559, n50560, n50561, n50562,
         n50563, n50564, n50565, n50566, n50567, n50568, n50569, n50570,
         n50571, n50572, n50573, n50574, n50575, n50576, n50577, n50578,
         n50579, n50580, n50581, n50582, n50583, n50584, n50585, n50586,
         n50587, n50588, n50589, n50590, n50591, n50592, n50593, n50594,
         n50595, n50596, n50597, n50598, n50599, n50600, n50601, n50602,
         n50603, n50604, n50605, n50606, n50607, n50608, n50609, n50610,
         n50611, n50612, n50613, n50614, n50615, n50616, n50617, n50618,
         n50619, n50620, n50621, n50622, n50623, n50624, n50625, n50626,
         n50627, n50628, n50629, n50630, n50631, n50632, n50633, n50634,
         n50635, n50636, n50637, n50638, n50639, n50640, n50641, n50642,
         n50643, n50644, n50645, n50646, n50647, n50648, n50649, n50650,
         n50651, n50652, n50653, n50654, n50655, n50656, n50657, n50658,
         n50659, n50660, n50661, n50662, n50663, n50664, n50665, n50666,
         n50667, n50668, n50669, n50670, n50671, n50672, n50673, n50674,
         n50675, n50676, n50677, n50678, n50679, n50680, n50681, n50682,
         n50683, n50684, n50685, n50686, n50687, n50688, n50689, n50690,
         n50691, n50692, n50693, n50694, n50695, n50696, n50697, n50698,
         n50699, n50700, n50701, n50702, n50703, n50704, n50705, n50706,
         n50707, n50708, n50709, n50710, n50711, n50712, n50713, n50714,
         n50715, n50716, n50717, n50718, n50719, n50720, n50721, n50722,
         n50723, n50724, n50725, n50726, n50727, n50728, n50729, n50730,
         n50731, n50732, n50733, n50734, n50735, n50736, n50737, n50738,
         n50739, n50740, n50741, n50742, n50743, n50744, n50745, n50746,
         n50747, n50748, n50749, n50750, n50751, n50752, n50753, n50754,
         n50755, n50756, n50757, n50758, n50759, n50760, n50761, n50762,
         n50763, n50764, n50765, n50766, n50767, n50768, n50769, n50770,
         n50771, n50772, n50773, n50774, n50775, n50776, n50777, n50778,
         n50779, n50780, n50781, n50782, n50783, n50784, n50785, n50786,
         n50787, n50788, n50789, n50790, n50791, n50792, n50793, n50794,
         n50795, n50796, n50797, n50798, n50799, n50800, n50801, n50802,
         n50803, n50804, n50805, n50806, n50807, n50808, n50809, n50810,
         n50811, n50812, n50813, n50814, n50815, n50816, n50817, n50818,
         n50819, n50820, n50821, n50822, n50823, n50824, n50825, n50826,
         n50827, n50828, n50829, n50830, n50831, n50832, n50833, n50834,
         n50835, n50836, n50837, n50838, n50839, n50840, n50841, n50842,
         n50843, n50844, n50845, n50846, n50847, n50848, n50849, n50850,
         n50851, n50852, n50853, n50854, n50855, n50856, n50857, n50858,
         n50859, n50860, n50861, n50862, n50863, n50864, n50865, n50866,
         n50867, n50868, n50869, n50870, n50871, n50872, n50873, n50874,
         n50875, n50876, n50877, n50878, n50879, n50880, n50881, n50882,
         n50883, n50884, n50885, n50886, n50887, n50888, n50889, n50890,
         n50891, n50892, n50893, n50894, n50895, n50896, n50897, n50898,
         n50899, n50900, n50901, n50902, n50903, n50904, n50905, n50906,
         n50907, n50908, n50909, n50910, n50911, n50912, n50913, n50914,
         n50915, n50916, n50917, n50918, n50919, n50920, n50921, n50922,
         n50923, n50924, n50925, n50926, n50927, n50928, n50929, n50930,
         n50931, n50932, n50933, n50934, n50935, n50936, n50937, n50938,
         n50939, n50940, n50941, n50942, n50943, n50944, n50945, n50946,
         n50947, n50948, n50949, n50950, n50951, n50952, n50953, n50954,
         n50955, n50956, n50957, n50958, n50959, n50960, n50961, n50962,
         n50963, n50964, n50965, n50966, n50967, n50968, n50969, n50970,
         n50971, n50972, n50973, n50974, n50975, n50976, n50977, n50978,
         n50979, n50980, n50981, n50982, n50983, n50984, n50985, n50986,
         n50987, n50988, n50989, n50990, n50991, n50992, n50993, n50994,
         n50995, n50996, n50997, n50998, n50999, n51000, n51001, n51002,
         n51003, n51004, n51005, n51006, n51007, n51008, n51009, n51010,
         n51011, n51012, n51013, n51014, n51015, n51016, n51017, n51018,
         n51019, n51020, n51021, n51022, n51023, n51024, n51025, n51026,
         n51027, n51028, n51029, n51030, n51031, n51032, n51033, n51034,
         n51035, n51036, n51037, n51038, n51039, n51040, n51041, n51042,
         n51043, n51044, n51045, n51046, n51047, n51048, n51049, n51050,
         n51051, n51052, n51053, n51054, n51055, n51056, n51057, n51058,
         n51059, n51060, n51061, n51062, n51063, n51064, n51065, n51066,
         n51067, n51068, n51069, n51070, n51071, n51072, n51073, n51074,
         n51075, n51076, n51077, n51078, n51079, n51080, n51081, n51082,
         n51083, n51084, n51085, n51086, n51087, n51088, n51089, n51090,
         n51091, n51092, n51093, n51094, n51095, n51096, n51097, n51098,
         n51099, n51100, n51101, n51102, n51103, n51104, n51105, n51106,
         n51107, n51108, n51109, n51110, n51111, n51112, n51113, n51114,
         n51115, n51116, n51117, n51118, n51119, n51120, n51121, n51122,
         n51123, n51124, n51125, n51126, n51127, n51128, n51129, n51130,
         n51131, n51132, n51133, n51134, n51135, n51136, n51137, n51138,
         n51139, n51140, n51141, n51142, n51143, n51144, n51145, n51146,
         n51147, n51148, n51149, n51150, n51151, n51152, n51153, n51154,
         n51155, n51156, n51157, n51158, n51159, n51160, n51161, n51162,
         n51163, n51164, n51165, n51166, n51167, n51168, n51169, n51170,
         n51171, n51172, n51173, n51174, n51175, n51176, n51177, n51178,
         n51179, n51180, n51181, n51182, n51183, n51184, n51185, n51186,
         n51187, n51188, n51189, n51190, n51191, n51192, n51193, n51194,
         n51195, n51196, n51197, n51198, n51199, n51200, n51201, n51202,
         n51203, n51204, n51205, n51206, n51207, n51208, n51209, n51210,
         n51211, n51212, n51213, n51214, n51215, n51216, n51217, n51218,
         n51219, n51220, n51221, n51222, n51223, n51224, n51225, n51226,
         n51227, n51228, n51229, n51230, n51231, n51232, n51233, n51234,
         n51235, n51236, n51237, n51238, n51239, n51240, n51241, n51242,
         n51243, n51244, n51245, n51246, n51247, n51248, n51249, n51250,
         n51251, n51252, n51253, n51254, n51255, n51256, n51257, n51258,
         n51259, n51260, n51261, n51262, n51263, n51264, n51265, n51266,
         n51267, n51268, n51269, n51270, n51271, n51272, n51273, n51274,
         n51275, n51276, n51277, n51278, n51279, n51280, n51281, n51282,
         n51283, n51284, n51285, n51286, n51287, n51288, n51289, n51290,
         n51291, n51292, n51293, n51294, n51295, n51296, n51297, n51298,
         n51299, n51300, n51301, n51302, n51303, n51304, n51305, n51306,
         n51307, n51308, n51309, n51310, n51311, n51312, n51313, n51314,
         n51315, n51316, n51317, n51318, n51319, n51320, n51321, n51322,
         n51323, n51324, n51325, n51326, n51327, n51328, n51329, n51330,
         n51331, n51332, n51333, n51334, n51335, n51336, n51337, n51338,
         n51339, n51340, n51341, n51342, n51343, n51344, n51345, n51346,
         n51347, n51348, n51349, n51350, n51351, n51352, n51353, n51354,
         n51355, n51356, n51357, n51358, n51359, n51360, n51361, n51362,
         n51363, n51364, n51365, n51366, n51367, n51368, n51369, n51370,
         n51371, n51372, n51373, n51374, n51375, n51376, n51377, n51378,
         n51379, n51380, n51381, n51382, n51383, n51384, n51385, n51386,
         n51387, n51388, n51389, n51390, n51391, n51392, n51393, n51394,
         n51395, n51396, n51397, n51398, n51399, n51400, n51401, n51402,
         n51403, n51404, n51405, n51406, n51407, n51408, n51409, n51410,
         n51411, n51412, n51413, n51414, n51415, n51416, n51417, n51418,
         n51419, n51420, n51421, n51422, n51423, n51424, n51425, n51426,
         n51427, n51428, n51429, n51430, n51431, n51432, n51433, n51434,
         n51435, n51436, n51437, n51438, n51439, n51440, n51441, n51442,
         n51443, n51444, n51445, n51446, n51447, n51448, n51449, n51450,
         n51451, n51452, n51453, n51454, n51455, n51456, n51457, n51458,
         n51459, n51460, n51461, n51462, n51463, n51464, n51465, n51466,
         n51467, n51468, n51469, n51470, n51471, n51472, n51473, n51474,
         n51475, n51476, n51477, n51478, n51479, n51480, n51481, n51482,
         n51483, n51484, n51485, n51486, n51487, n51488, n51489, n51490,
         n51491, n51492, n51493, n51494, n51495, n51496, n51497, n51498,
         n51499, n51500, n51501, n51502, n51503, n51504, n51505, n51506,
         n51507, n51508, n51509, n51510, n51511, n51512, n51513, n51514,
         n51515, n51516, n51517, n51518, n51519, n51520, n51521, n51522,
         n51523, n51524, n51525, n51526, n51527, n51528, n51529, n51530,
         n51531, n51532, n51533, n51534, n51535, n51536, n51537, n51538,
         n51539, n51540, n51541, n51542, n51543, n51544, n51545, n51546,
         n51547, n51548, n51549, n51550, n51551, n51552, n51553, n51554,
         n51555, n51556, n51557, n51558, n51559, n51560, n51561, n51562,
         n51563, n51564, n51565, n51566, n51567, n51568, n51569, n51570,
         n51571, n51572, n51573, n51574, n51575, n51576, n51577, n51578,
         n51579, n51580, n51581, n51582, n51583, n51584, n51585, n51586,
         n51587, n51588, n51589, n51590, n51591, n51592, n51593, n51594,
         n51595, n51596, n51597, n51598, n51599, n51600, n51601, n51602,
         n51603, n51604, n51605, n51606, n51607, n51608, n51609, n51610,
         n51611, n51612, n51613, n51614, n51615, n51616, n51617, n51618,
         n51619, n51620, n51621, n51622, n51623, n51624, n51625, n51626,
         n51627, n51628, n51629, n51630, n51631, n51632, n51633, n51634,
         n51635, n51636, n51637, n51638, n51639, n51640, n51641, n51642,
         n51643, n51644, n51645, n51646, n51647, n51648, n51649, n51650,
         n51651, n51652, n51653, n51654, n51655, n51656, n51657, n51658,
         n51659, n51660, n51661, n51662, n51663, n51664, n51665, n51666,
         n51667, n51668, n51669, n51670, n51671, n51672, n51673, n51674,
         n51675, n51676, n51677, n51678, n51679, n51680, n51681, n51682,
         n51683, n51684, n51685, n51686, n51687, n51688, n51689, n51690,
         n51691, n51692, n51693, n51694, n51695, n51696, n51697, n51698,
         n51699, n51700, n51701, n51702, n51703, n51704, n51705, n51706,
         n51707, n51708, n51709, n51710, n51711, n51712, n51713, n51714,
         n51715, n51716, n51717, n51718, n51719, n51720, n51721, n51722,
         n51723, n51724, n51725, n51726, n51727, n51728, n51729, n51730,
         n51731, n51732, n51733, n51734, n51735, n51736, n51737, n51738,
         n51739, n51740, n51741, n51742, n51743, n51744, n51745, n51746,
         n51747, n51748, n51749, n51750, n51751, n51752, n51753, n51754,
         n51755, n51756, n51757, n51758, n51759, n51760, n51761, n51762,
         n51763, n51764, n51765, n51766, n51767, n51768, n51769, n51770,
         n51771, n51772, n51773, n51774, n51775, n51776, n51777, n51778,
         n51779, n51780, n51781, n51782, n51783, n51784, n51785, n51786,
         n51787, n51788, n51789, n51790, n51791, n51792, n51793, n51794,
         n51795, n51796, n51797, n51798, n51799, n51800, n51801, n51802,
         n51803, n51804, n51805, n51806, n51807, n51808, n51809, n51810,
         n51811, n51812, n51813, n51814, n51815, n51816, n51817, n51818,
         n51819, n51820, n51821, n51822, n51823, n51824, n51825, n51826,
         n51827, n51828, n51829, n51830, n51831, n51832, n51833, n51834,
         n51835, n51836, n51837, n51838, n51839, n51840, n51841, n51842,
         n51843, n51844, n51845, n51846, n51847, n51848, n51849, n51850,
         n51851, n51852, n51853, n51854, n51855, n51856, n51857, n51858,
         n51859, n51860, n51861, n51862, n51863, n51864, n51865, n51866,
         n51867, n51868, n51869, n51870, n51871, n51872, n51873, n51874,
         n51875, n51876, n51877, n51878, n51879, n51880, n51881, n51882,
         n51883, n51884, n51885, n51886, n51887, n51888, n51889, n51890,
         n51891, n51892, n51893, n51894, n51895, n51896, n51897, n51898,
         n51899, n51900, n51901, n51902, n51903, n51904, n51905, n51906,
         n51907, n51908, n51909, n51910, n51911, n51912, n51913, n51914,
         n51915, n51916, n51917, n51918, n51919, n51920, n51921, n51922,
         n51923, n51924, n51925, n51926, n51927, n51928, n51929, n51930,
         n51931, n51932, n51933, n51934, n51935, n51936, n51937, n51938,
         n51939, n51940, n51941, n51942, n51943, n51944, n51945, n51946,
         n51947, n51948, n51949, n51950, n51951, n51952, n51953, n51954,
         n51955, n51956, n51957, n51958, n51959, n51960, n51961, n51962,
         n51963, n51964, n51965, n51966, n51967, n51968, n51969, n51970,
         n51971, n51972, n51973, n51974, n51975, n51976, n51977, n51978,
         n51979, n51980, n51981, n51982, n51983, n51984, n51985, n51986,
         n51987, n51988, n51989, n51990, n51991, n51992, n51993, n51994,
         n51995, n51996, n51997, n51998, n51999, n52000, n52001, n52002,
         n52003, n52004, n52005, n52006, n52007, n52008, n52009, n52010,
         n52011, n52012, n52013, n52014, n52015, n52016, n52017, n52018,
         n52019, n52020, n52021, n52022, n52023, n52024, n52025, n52026,
         n52027, n52028, n52029, n52030, n52031, n52032, n52033, n52034,
         n52035, n52036, n52037, n52038, n52039, n52040, n52041, n52042,
         n52043, n52044, n52045, n52046, n52047, n52048, n52049, n52050,
         n52051, n52052, n52053, n52054, n52055, n52056, n52057, n52058,
         n52059, n52060, n52061, n52062, n52063, n52064, n52065, n52066,
         n52067, n52068, n52069, n52070, n52071, n52072, n52073, n52074,
         n52075, n52076, n52077, n52078, n52079, n52080, n52081, n52082,
         n52083, n52084, n52085, n52086, n52087, n52088, n52089, n52090,
         n52091, n52092, n52093, n52094, n52095, n52096, n52097, n52098,
         n52099, n52100, n52101, n52102, n52103, n52104, n52105, n52106,
         n52107, n52108, n52109, n52110, n52111, n52112, n52113, n52114,
         n52115, n52116, n52117, n52118, n52119, n52120, n52121, n52122,
         n52123, n52124, n52125, n52126, n52127, n52128, n52129, n52130,
         n52131, n52132, n52133, n52134, n52135, n52136, n52137, n52138,
         n52139, n52140, n52141, n52142, n52143, n52144, n52145, n52146,
         n52147, n52148, n52149, n52150, n52151, n52152, n52153, n52154,
         n52155, n52156, n52157, n52158, n52159, n52160, n52161, n52162,
         n52163, n52164, n52165, n52166, n52167, n52168, n52169, n52170,
         n52171, n52172, n52173, n52174, n52175, n52176, n52177, n52178,
         n52179, n52180, n52181, n52182, n52183, n52184, n52185, n52186,
         n52187, n52188, n52189, n52190, n52191, n52192, n52193, n52194,
         n52195, n52196, n52197, n52198, n52199, n52200, n52201, n52202,
         n52203, n52204, n52205, n52206, n52207, n52208, n52209, n52210,
         n52211, n52212, n52213, n52214, n52215, n52216, n52217, n52218,
         n52219, n52220, n52221, n52222, n52223, n52224, n52225, n52226,
         n52227, n52228, n52229, n52230, n52231, n52232, n52233, n52234,
         n52235, n52236, n52237, n52238, n52239, n52240, n52241, n52242,
         n52243, n52244, n52245, n52246, n52247, n52248, n52249, n52250,
         n52251, n52252, n52253, n52254, n52255, n52256, n52257, n52258,
         n52259, n52260, n52261, n52262, n52263, n52264, n52265, n52266,
         n52267, n52268, n52269, n52270, n52271, n52272, n52273, n52274,
         n52275, n52276, n52277, n52278, n52279, n52280, n52281, n52282,
         n52283, n52284, n52285, n52286, n52287, n52288, n52289, n52290,
         n52291, n52292, n52293, n52294, n52295, n52296, n52297, n52298,
         n52299, n52300, n52301, n52302, n52303, n52304, n52305, n52306,
         n52307, n52308, n52309, n52310, n52311, n52312, n52313, n52314,
         n52315, n52316, n52317, n52318, n52319, n52320, n52321, n52322,
         n52323, n52324, n52325, n52326, n52327, n52328, n52329, n52330,
         n52331, n52332, n52333, n52334, n52335, n52336, n52337, n52338,
         n52339, n52340, n52341, n52342, n52343, n52344, n52345, n52346,
         n52347, n52348, n52349, n52350, n52351, n52352, n52353, n52354,
         n52355, n52356, n52357, n52358, n52359, n52360, n52361, n52362,
         n52363, n52364, n52365, n52366, n52367, n52368, n52369, n52370,
         n52371, n52372, n52373, n52374, n52375, n52376, n52377, n52378,
         n52379, n52380, n52381, n52382, n52383, n52384, n52385, n52386,
         n52387, n52388, n52389, n52390, n52391, n52392, n52393, n52394,
         n52395, n52396, n52397, n52398, n52399, n52400, n52401, n52402,
         n52403, n52404, n52405, n52406, n52407, n52408, n52409, n52410,
         n52411, n52412, n52413, n52414, n52415, n52416, n52417, n52418,
         n52419, n52420, n52421, n52422, n52423, n52424, n52425, n52426,
         n52427, n52428, n52429, n52430, n52431, n52432, n52433, n52434,
         n52435, n52436, n52437, n52438, n52439, n52440, n52441, n52442,
         n52443, n52444, n52445, n52446, n52447, n52448, n52449, n52450,
         n52451, n52452, n52453, n52454, n52455, n52456, n52457, n52458,
         n52459, n52460, n52461, n52462, n52463, n52464, n52465, n52466,
         n52467, n52468, n52469, n52470, n52471, n52472, n52473, n52474,
         n52475, n52476, n52477, n52478, n52479, n52480, n52481, n52482,
         n52483, n52484, n52485, n52486, n52487, n52488, n52489, n52490,
         n52491, n52492, n52493, n52494, n52495, n52496, n52497, n52498,
         n52499, n52500, n52501, n52502, n52503, n52504, n52505, n52506,
         n52507, n52508, n52509, n52510, n52511, n52512, n52513, n52514,
         n52515, n52516, n52517, n52518, n52519, n52520, n52521, n52522,
         n52523, n52524, n52525, n52526, n52527, n52528, n52529, n52530,
         n52531, n52532, n52533, n52534, n52535, n52536, n52537, n52538,
         n52539, n52540, n52541, n52542, n52543, n52544, n52545, n52546,
         n52547, n52548, n52549, n52550, n52551, n52552, n52553, n52554,
         n52555, n52556, n52557, n52558, n52559, n52560, n52561, n52562,
         n52563, n52564, n52565, n52566, n52567, n52568, n52569, n52570,
         n52571, n52572, n52573, n52574, n52575, n52576, n52577, n52578,
         n52579, n52580, n52581, n52582, n52583, n52584, n52585, n52586,
         n52587, n52588, n52589, n52590, n52591, n52592, n52593, n52594,
         n52595, n52596, n52597, n52598, n52599, n52600, n52601, n52602,
         n52603, n52604, n52605, n52606, n52607, n52608, n52609, n52610,
         n52611, n52612, n52613, n52614, n52615, n52616, n52617, n52618,
         n52619, n52620, n52621, n52622, n52623, n52624, n52625, n52626,
         n52627, n52628, n52629, n52630, n52631, n52632, n52633, n52634,
         n52635, n52636, n52637, n52638, n52639, n52640, n52641, n52642,
         n52643, n52644, n52645, n52646, n52647, n52648, n52649, n52650,
         n52651, n52652, n52653, n52654, n52655, n52656, n52657, n52658,
         n52659, n52660, n52661, n52662, n52663, n52664, n52665, n52666,
         n52667, n52668, n52669, n52670, n52671, n52672, n52673, n52674,
         n52675, n52676, n52677, n52678, n52679, n52680, n52681, n52682,
         n52683, n52684, n52685, n52686, n52687, n52688, n52689, n52690,
         n52691, n52692, n52693, n52694, n52695, n52696, n52697, n52698,
         n52699, n52700, n52701, n52702, n52703, n52704, n52705, n52706,
         n52707, n52708, n52709, n52710, n52711, n52712, n52713, n52714,
         n52715, n52716, n52717, n52718, n52719, n52720, n52721, n52722,
         n52723, n52724, n52725, n52726, n52727, n52728, n52729, n52730,
         n52731, n52732, n52733, n52734, n52735, n52736, n52737, n52738,
         n52739, n52740, n52741, n52742, n52743, n52744, n52745, n52746,
         n52747, n52748, n52749, n52750, n52751, n52752, n52753, n52754,
         n52755, n52756, n52757, n52758, n52759, n52760, n52761, n52762,
         n52763, n52764, n52765, n52766, n52767, n52768, n52769, n52770,
         n52771, n52772, n52773, n52774, n52775, n52776, n52777, n52778,
         n52779, n52780, n52781, n52782, n52783, n52784, n52785, n52786,
         n52787, n52788, n52789, n52790, n52791, n52792, n52793, n52794,
         n52795, n52796, n52797, n52798, n52799, n52800, n52801, n52802,
         n52803, n52804, n52805, n52806, n52807, n52808, n52809, n52810,
         n52811, n52812, n52813, n52814, n52815, n52816, n52817, n52818,
         n52819, n52820, n52821, n52822, n52823, n52824, n52825, n52826,
         n52827, n52828, n52829, n52830, n52831, n52832, n52833, n52834,
         n52835, n52836, n52837, n52838, n52839, n52840, n52841, n52842,
         n52843, n52844, n52845, n52846, n52847, n52848, n52849, n52850,
         n52851, n52852, n52853, n52854, n52855, n52856, n52857, n52858,
         n52859, n52860, n52861, n52862, n52863, n52864, n52865, n52866,
         n52867, n52868, n52869, n52870, n52871, n52872, n52873, n52874,
         n52875, n52876, n52877, n52878, n52879, n52880, n52881, n52882,
         n52883, n52884, n52885, n52886, n52887, n52888, n52889, n52890,
         n52891, n52892, n52893, n52894, n52895, n52896, n52897, n52898,
         n52899, n52900, n52901, n52902, n52903, n52904, n52905, n52906,
         n52907, n52908, n52909, n52910, n52911, n52912, n52913, n52914,
         n52915, n52916, n52917, n52918, n52919, n52920, n52921, n52922,
         n52923, n52924, n52925, n52926, n52927, n52928, n52929, n52930,
         n52931, n52932, n52933, n52934, n52935, n52936, n52937, n52938,
         n52939, n52940, n52941, n52942, n52943, n52944, n52945, n52946,
         n52947, n52948, n52949, n52950, n52951, n52952, n52953, n52954,
         n52955, n52956, n52957, n52958, n52959, n52960, n52961, n52962,
         n52963, n52964, n52965, n52966, n52967, n52968, n52969, n52970,
         n52971, n52972, n52973, n52974, n52975, n52976, n52977, n52978,
         n52979, n52980, n52981, n52982, n52983, n52984, n52985, n52986,
         n52987, n52988, n52989, n52990, n52991, n52992, n52993, n52994,
         n52995, n52996, n52997, n52998, n52999, n53000, n53001, n53002,
         n53003, n53004, n53005, n53006, n53007, n53008, n53009, n53010,
         n53011, n53012, n53013, n53014, n53015, n53016, n53017, n53018,
         n53019, n53020, n53021, n53022, n53023, n53024, n53025, n53026,
         n53027, n53028, n53029, n53030, n53031, n53032, n53033, n53034,
         n53035, n53036, n53037, n53038, n53039, n53040, n53041, n53042,
         n53043, n53044, n53045, n53046, n53047, n53048, n53049, n53050,
         n53051, n53052, n53053, n53054, n53055, n53056, n53057, n53058,
         n53059, n53060, n53061, n53062, n53063, n53064, n53065, n53066,
         n53067, n53068, n53069, n53070, n53071, n53072, n53073, n53074,
         n53075, n53076, n53077, n53078, n53079, n53080, n53081, n53082,
         n53083, n53084, n53085, n53086, n53087, n53088, n53089, n53090,
         n53091, n53092, n53093, n53094, n53095, n53096, n53097, n53098,
         n53099, n53100, n53101, n53102, n53103, n53104, n53105, n53106,
         n53107, n53108, n53109, n53110, n53111, n53112, n53113, n53114,
         n53115, n53116, n53117, n53118, n53119, n53120, n53121, n53122,
         n53123, n53124, n53125, n53126, n53127, n53128, n53129, n53130,
         n53131, n53132, n53133, n53134, n53135, n53136, n53137, n53138,
         n53139, n53140, n53141, n53142, n53143, n53144, n53145, n53146,
         n53147, n53148, n53149, n53150, n53151, n53152, n53153, n53154,
         n53155, n53156, n53157, n53158, n53159, n53160, n53161, n53162,
         n53163, n53164, n53165, n53166, n53167, n53168, n53169, n53170,
         n53171, n53172, n53173, n53174, n53175, n53176, n53177, n53178,
         n53179, n53180, n53181, n53182, n53183, n53184, n53185, n53186,
         n53187, n53188, n53189, n53190, n53191, n53192, n53193, n53194,
         n53195, n53196, n53197, n53198, n53199, n53200, n53201, n53202,
         n53203, n53204, n53205, n53206, n53207, n53208, n53209, n53210,
         n53211, n53212, n53213, n53214, n53215, n53216, n53217, n53218,
         n53219, n53220, n53221, n53222, n53223, n53224, n53225, n53226,
         n53227, n53228, n53229, n53230, n53231, n53232, n53233, n53234,
         n53235, n53236, n53237, n53238, n53239, n53240, n53241, n53242,
         n53243, n53244, n53245, n53246, n53247, n53248, n53249, n53250,
         n53251, n53252, n53253, n53254, n53255, n53256, n53257, n53258,
         n53259, n53260, n53261, n53262, n53263, n53264, n53265, n53266,
         n53267, n53268, n53269, n53270, n53271, n53272, n53273, n53274,
         n53275, n53276, n53277, n53278, n53279, n53280, n53281, n53282,
         n53283, n53284, n53285, n53286, n53287, n53288, n53289, n53290,
         n53291, n53292, n53293, n53294, n53295, n53296, n53297, n53298,
         n53299, n53300, n53301, n53302, n53303, n53304, n53305, n53306,
         n53307, n53308, n53309, n53310, n53311, n53312, n53313, n53314,
         n53315, n53316, n53317, n53318, n53319, n53320, n53321, n53322,
         n53323, n53324, n53325, n53326, n53327, n53328, n53329, n53330,
         n53331, n53332, n53333, n53334, n53335, n53336, n53337, n53338,
         n53339, n53340, n53341, n53342, n53343, n53344, n53345, n53346,
         n53347, n53348, n53349, n53350, n53351, n53352, n53353, n53354,
         n53355, n53356, n53357, n53358, n53359, n53360, n53361, n53362,
         n53363, n53364, n53365, n53366, n53367, n53368, n53369, n53370,
         n53371, n53372, n53373, n53374, n53375, n53376, n53377, n53378,
         n53379, n53380, n53381, n53382, n53383, n53384, n53385, n53386,
         n53387, n53388, n53389, n53390, n53391, n53392, n53393, n53394,
         n53395, n53396, n53397, n53398, n53399, n53400, n53401, n53402,
         n53403, n53404, n53405, n53406, n53407, n53408, n53409, n53410,
         n53411, n53412, n53413, n53414, n53415, n53416, n53417, n53418,
         n53419, n53420, n53421, n53422, n53423, n53424, n53425, n53426,
         n53427, n53428, n53429, n53430, n53431, n53432, n53433, n53434,
         n53435, n53436, n53437, n53438, n53439, n53440, n53441, n53442,
         n53443, n53444, n53445, n53446, n53447, n53448, n53449, n53450,
         n53451, n53452, n53453, n53454, n53455, n53456, n53457, n53458,
         n53459, n53460, n53461, n53462, n53463, n53464, n53465, n53466,
         n53467, n53468, n53469, n53470, n53471, n53472, n53473, n53474,
         n53475, n53476, n53477, n53478, n53479, n53480, n53481, n53482,
         n53483, n53484, n53485, n53486, n53487, n53488, n53489, n53490,
         n53491, n53492, n53493, n53494, n53495, n53496, n53497, n53498,
         n53499, n53500, n53501, n53502, n53503, n53504, n53505, n53506,
         n53507, n53508, n53509, n53510, n53511, n53512, n53513, n53514,
         n53515, n53516, n53517, n53518, n53519, n53520, n53521, n53522,
         n53523, n53524, n53525, n53526, n53527, n53528, n53529, n53530,
         n53531, n53532, n53533, n53534, n53535, n53536, n53537, n53538,
         n53539, n53540, n53541, n53542, n53543, n53544, n53545, n53546,
         n53547, n53548, n53549, n53550, n53551, n53552, n53553, n53554,
         n53555, n53556, n53557, n53558, n53559, n53560, n53561, n53562,
         n53563, n53564, n53565, n53566, n53567, n53568, n53569, n53570,
         n53571, n53572, n53573, n53574, n53575, n53576, n53577, n53578,
         n53579, n53580, n53581, n53582, n53583, n53584, n53585, n53586,
         n53587, n53588, n53589, n53590, n53591, n53592, n53593, n53594,
         n53595, n53596, n53597, n53598, n53599, n53600, n53601, n53602,
         n53603, n53604, n53605, n53606, n53607, n53608, n53609, n53610,
         n53611, n53612, n53613, n53614, n53615, n53616, n53617, n53618,
         n53619, n53620, n53621, n53622, n53623, n53624, n53625, n53626,
         n53627, n53628, n53629, n53630, n53631, n53632, n53633, n53634,
         n53635, n53636, n53637, n53638, n53639, n53640, n53641, n53642,
         n53643, n53644, n53645, n53646, n53647, n53648, n53649, n53650,
         n53651, n53652, n53653, n53654, n53655, n53656, n53657, n53658,
         n53659, n53660, n53661, n53662, n53663, n53664, n53665, n53666,
         n53667, n53668, n53669, n53670, n53671, n53672, n53673, n53674,
         n53675, n53676, n53677, n53678, n53679, n53680, n53681, n53682,
         n53683, n53684, n53685, n53686, n53687, n53688, n53689, n53690,
         n53691, n53692, n53693, n53694, n53695, n53696, n53697, n53698,
         n53699, n53700, n53701, n53702, n53703, n53704, n53705, n53706,
         n53707, n53708, n53709, n53710, n53711, n53712, n53713, n53714,
         n53715, n53716, n53717, n53718, n53719, n53720, n53721, n53722,
         n53723, n53724, n53725, n53726, n53727, n53728, n53729, n53730,
         n53731, n53732, n53733, n53734, n53735, n53736, n53737, n53738,
         n53739, n53740, n53741, n53742, n53743, n53744, n53745, n53746,
         n53747, n53748, n53749, n53750, n53751, n53752, n53753, n53754,
         n53755, n53756, n53757, n53758, n53759, n53760, n53761, n53762,
         n53763, n53764, n53765, n53766, n53767, n53768, n53769, n53770,
         n53771, n53772, n53773, n53774, n53775, n53776, n53777, n53778,
         n53779, n53780, n53781, n53782, n53783, n53784, n53785, n53786,
         n53787, n53788, n53789, n53790, n53791, n53792, n53793, n53794,
         n53795, n53796, n53797, n53798, n53799, n53800, n53801, n53802,
         n53803, n53804, n53805, n53806, n53807, n53808, n53809, n53810,
         n53811, n53812, n53813, n53814, n53815, n53816, n53817, n53818,
         n53819, n53820, n53821, n53822, n53823, n53824, n53825, n53826,
         n53827, n53828, n53829, n53830, n53831, n53832, n53833, n53834,
         n53835, n53836, n53837, n53838, n53839, n53840, n53841, n53842,
         n53843, n53844, n53845, n53846, n53847, n53848, n53849, n53850,
         n53851, n53852, n53853, n53854, n53855, n53856, n53857, n53858,
         n53859, n53860, n53861, n53862, n53863, n53864, n53865, n53866,
         n53867, n53868, n53869, n53870, n53871, n53872, n53873, n53874,
         n53875, n53876, n53877, n53878, n53879, n53880, n53881, n53882,
         n53883, n53884, n53885, n53886, n53887, n53888, n53889, n53890,
         n53891, n53892, n53893, n53894, n53895, n53896, n53897, n53898,
         n53899, n53900, n53901, n53902, n53903, n53904, n53905, n53906,
         n53907, n53908, n53909, n53910, n53911, n53912, n53913, n53914,
         n53915, n53916, n53917, n53918, n53919, n53920, n53921, n53922,
         n53923, n53924, n53925, n53926, n53927, n53928, n53929, n53930,
         n53931, n53932, n53933, n53934, n53935, n53936, n53937, n53938,
         n53939, n53940, n53941, n53942, n53943, n53944, n53945, n53946,
         n53947, n53948, n53949, n53950, n53951, n53952, n53953, n53954,
         n53955, n53956, n53957, n53958, n53959, n53960, n53961, n53962,
         n53963, n53964, n53965, n53966, n53967, n53968, n53969, n53970,
         n53971, n53972, n53973, n53974, n53975, n53976, n53977, n53978,
         n53979, n53980, n53981, n53982, n53983, n53984, n53985, n53986,
         n53987, n53988, n53989, n53990, n53991, n53992, n53993, n53994,
         n53995, n53996, n53997, n53998, n53999, n54000, n54001, n54002,
         n54003, n54004, n54005, n54006, n54007, n54008, n54009, n54010,
         n54011, n54012, n54013, n54014, n54015, n54016, n54017, n54018,
         n54019, n54020, n54021, n54022, n54023, n54024, n54025, n54026,
         n54027, n54028, n54029, n54030, n54031, n54032, n54033, n54034,
         n54035, n54036, n54037, n54038, n54039, n54040, n54041, n54042,
         n54043, n54044, n54045, n54046, n54047, n54048, n54049, n54050,
         n54051, n54052, n54053, n54054, n54055, n54056, n54057, n54058,
         n54059, n54060, n54061, n54062, n54063, n54064, n54065, n54066,
         n54067, n54068, n54069, n54070, n54071, n54072, n54073, n54074,
         n54075, n54076, n54077, n54078, n54079, n54080, n54081, n54082,
         n54083, n54084, n54085, n54086, n54087, n54088, n54089, n54090,
         n54091, n54092, n54093, n54094, n54095, n54096, n54097, n54098,
         n54099, n54100, n54101, n54102, n54103, n54104, n54105, n54106,
         n54107, n54108, n54109, n54110, n54111, n54112, n54113, n54114,
         n54115, n54116, n54117, n54118, n54119, n54120, n54121, n54122,
         n54123, n54124, n54125, n54126, n54127, n54128, n54129, n54130,
         n54131, n54132, n54133, n54134, n54135, n54136, n54137, n54138,
         n54139, n54140, n54141, n54142, n54143, n54144, n54145, n54146,
         n54147, n54148, n54149, n54150, n54151, n54152, n54153, n54154,
         n54155, n54156, n54157, n54158, n54159, n54160, n54161, n54162,
         n54163, n54164, n54165, n54166, n54167, n54168, n54169, n54170,
         n54171, n54172, n54173, n54174, n54175, n54176, n54177, n54178,
         n54179, n54180, n54181, n54182, n54183, n54184, n54185, n54186,
         n54187, n54188, n54189, n54190, n54191, n54192, n54193, n54194,
         n54195, n54196, n54197, n54198, n54199, n54200, n54201, n54202,
         n54203, n54204, n54205, n54206, n54207, n54208, n54209, n54210,
         n54211, n54212, n54213, n54214, n54215, n54216, n54217, n54218,
         n54219, n54220, n54221, n54222, n54223, n54224, n54225, n54226,
         n54227, n54228, n54229, n54230, n54231, n54232, n54233, n54234,
         n54235, n54236, n54237, n54238, n54239, n54240, n54241, n54242,
         n54243, n54244, n54245, n54246, n54247, n54248, n54249, n54250,
         n54251, n54252, n54253, n54254, n54255, n54256, n54257, n54258,
         n54259, n54260, n54261, n54262, n54263, n54264, n54265, n54266,
         n54267, n54268, n54269, n54270, n54271, n54272, n54273, n54274,
         n54275, n54276, n54277, n54278, n54279, n54280, n54281, n54282,
         n54283, n54284, n54285, n54286, n54287, n54288, n54289, n54290,
         n54291, n54292, n54293, n54294, n54295, n54296, n54297, n54298,
         n54299, n54300, n54301, n54302, n54303, n54304, n54305, n54306,
         n54307, n54308, n54309, n54310, n54311, n54312, n54313, n54314,
         n54315, n54316, n54317, n54318, n54319, n54320, n54321, n54322,
         n54323, n54324, n54325, n54326, n54327, n54328, n54329, n54330,
         n54331, n54332, n54333, n54334, n54335, n54336, n54337, n54338,
         n54339, n54340, n54341, n54342, n54343, n54344, n54345, n54346,
         n54347, n54348, n54349, n54350, n54351, n54352, n54353, n54354,
         n54355, n54356, n54357, n54358, n54359, n54360, n54361, n54362,
         n54363, n54364, n54365, n54366, n54367, n54368, n54369, n54370,
         n54371, n54372, n54373, n54374, n54375, n54376, n54377, n54378,
         n54379, n54380, n54381, n54382, n54383, n54384, n54385, n54386,
         n54387, n54388, n54389, n54390, n54391, n54392, n54393, n54394,
         n54395, n54396, n54397, n54398, n54399, n54400, n54401, n54402,
         n54403, n54404, n54405, n54406, n54407, n54408, n54409, n54410,
         n54411, n54412, n54413, n54414, n54415, n54416, n54417, n54418,
         n54419, n54420, n54421, n54422, n54423, n54424, n54425, n54426,
         n54427, n54428, n54429, n54430, n54431, n54432, n54433, n54434,
         n54435, n54436, n54437, n54438, n54439, n54440, n54441, n54442,
         n54443, n54444, n54445, n54446, n54447, n54448, n54449, n54450,
         n54451, n54452, n54453, n54454, n54455, n54456, n54457, n54458,
         n54459, n54460, n54461, n54462, n54463, n54464, n54465, n54466,
         n54467, n54468, n54469, n54470, n54471, n54472, n54473, n54474,
         n54475, n54476, n54477, n54478, n54479, n54480, n54481, n54482,
         n54483, n54484, n54485, n54486, n54487, n54488, n54489, n54490,
         n54491, n54492, n54493, n54494, n54495, n54496, n54497, n54498,
         n54499, n54500, n54501, n54502, n54503, n54504, n54505, n54506,
         n54507, n54508, n54509, n54510, n54511, n54512, n54513, n54514,
         n54515, n54516, n54517, n54518, n54519, n54520, n54521, n54522,
         n54523, n54524, n54525, n54526, n54527, n54528, n54529, n54530,
         n54531, n54532, n54533, n54534, n54535, n54536, n54537, n54538,
         n54539, n54540, n54541, n54542, n54543, n54544, n54545, n54546,
         n54547, n54548, n54549, n54550, n54551, n54552, n54553, n54554,
         n54555, n54556, n54557, n54558, n54559, n54560, n54561, n54562,
         n54563, n54564, n54565, n54566, n54567, n54568, n54569, n54570,
         n54571, n54572, n54573, n54574, n54575, n54576, n54577, n54578,
         n54579, n54580, n54581, n54582, n54583, n54584, n54585, n54586,
         n54587, n54588, n54589, n54590, n54591, n54592, n54593, n54594,
         n54595, n54596, n54597, n54598, n54599, n54600, n54601, n54602,
         n54603, n54604, n54605, n54606, n54607, n54608, n54609, n54610,
         n54611, n54612, n54613, n54614, n54615, n54616, n54617, n54618,
         n54619, n54620, n54621, n54622, n54623, n54624, n54625, n54626,
         n54627, n54628, n54629, n54630, n54631, n54632, n54633, n54634,
         n54635, n54636, n54637, n54638, n54639, n54640, n54641, n54642,
         n54643, n54644, n54645, n54646, n54647, n54648, n54649, n54650,
         n54651, n54652, n54653, n54654, n54655, n54656, n54657, n54658,
         n54659, n54660, n54661, n54662, n54663, n54664, n54665, n54666,
         n54667, n54668, n54669, n54670, n54671, n54672, n54673, n54674,
         n54675, n54676, n54677, n54678, n54679, n54680, n54681, n54682,
         n54683, n54684, n54685, n54686, n54687, n54688, n54689, n54690,
         n54691, n54692, n54693, n54694, n54695, n54696, n54697, n54698,
         n54699, n54700, n54701, n54702, n54703, n54704, n54705, n54706,
         n54707, n54708, n54709, n54710, n54711, n54712, n54713, n54714,
         n54715, n54716, n54717, n54718, n54719, n54720, n54721, n54722,
         n54723, n54724, n54725, n54726, n54727, n54728, n54729, n54730,
         n54731, n54732, n54733, n54734, n54735, n54736, n54737, n54738,
         n54739, n54740, n54741, n54742, n54743, n54744, n54745, n54746,
         n54747, n54748, n54749, n54750, n54751, n54752, n54753, n54754,
         n54755, n54756, n54757, n54758, n54759, n54760, n54761, n54762,
         n54763, n54764, n54765, n54766, n54767, n54768, n54769, n54770,
         n54771, n54772, n54773, n54774, n54775, n54776, n54777, n54778,
         n54779, n54780, n54781, n54782, n54783, n54784, n54785, n54786,
         n54787, n54788, n54789, n54790, n54791, n54792, n54793, n54794,
         n54795, n54796, n54797, n54798, n54799, n54800, n54801, n54802,
         n54803, n54804, n54805, n54806, n54807, n54808, n54809, n54810,
         n54811, n54812, n54813, n54814, n54815, n54816, n54817, n54818,
         n54819, n54820, n54821, n54822, n54823, n54824, n54825, n54826,
         n54827, n54828, n54829, n54830, n54831, n54832, n54833, n54834,
         n54835, n54836, n54837, n54838, n54839, n54840, n54841, n54842,
         n54843, n54844, n54845, n54846, n54847, n54848, n54849, n54850,
         n54851, n54852, n54853, n54854, n54855, n54856, n54857, n54858,
         n54859, n54860, n54861, n54862, n54863, n54864, n54865, n54866,
         n54867, n54868, n54869, n54870, n54871, n54872, n54873, n54874,
         n54875, n54876, n54877, n54878, n54879, n54880, n54881, n54882,
         n54883, n54884, n54885, n54886, n54887, n54888, n54889, n54890,
         n54891, n54892, n54893, n54894, n54895, n54896, n54897, n54898,
         n54899, n54900, n54901, n54902, n54903, n54904, n54905, n54906,
         n54907, n54908, n54909, n54910, n54911, n54912, n54913, n54914,
         n54915, n54916, n54917, n54918, n54919, n54920, n54921, n54922,
         n54923, n54924, n54925, n54926, n54927, n54928, n54929, n54930,
         n54931, n54932, n54933, n54934, n54935, n54936, n54937, n54938,
         n54939, n54940, n54941, n54942, n54943, n54944, n54945, n54946,
         n54947, n54948, n54949, n54950, n54951, n54952, n54953, n54954,
         n54955, n54956, n54957, n54958, n54959, n54960, n54961, n54962,
         n54963, n54964, n54965, n54966, n54967, n54968, n54969, n54970,
         n54971, n54972, n54973, n54974, n54975, n54976, n54977, n54978,
         n54979, n54980, n54981, n54982, n54983, n54984, n54985, n54986,
         n54987, n54988, n54989, n54990, n54991, n54992, n54993, n54994,
         n54995, n54996, n54997, n54998, n54999, n55000, n55001, n55002,
         n55003, n55004, n55005, n55006, n55007, n55008, n55009, n55010,
         n55011, n55012, n55013, n55014, n55015, n55016, n55017, n55018,
         n55019, n55020, n55021, n55022, n55023, n55024, n55025, n55026,
         n55027, n55028, n55029, n55030, n55031, n55032, n55033, n55034,
         n55035, n55036, n55037, n55038, n55039, n55040, n55041, n55042,
         n55043, n55044, n55045, n55046, n55047, n55048, n55049, n55050,
         n55051, n55052, n55053, n55054, n55055, n55056, n55057, n55058,
         n55059, n55060, n55061, n55062, n55063, n55064, n55065, n55066,
         n55067, n55068, n55069, n55070, n55071, n55072, n55073, n55074,
         n55075, n55076, n55077, n55078, n55079, n55080, n55081, n55082,
         n55083, n55084, n55085, n55086, n55087, n55088, n55089, n55090,
         n55091, n55092, n55093, n55094, n55095, n55096, n55097, n55098,
         n55099, n55100, n55101, n55102, n55103, n55104, n55105, n55106,
         n55107, n55108, n55109, n55110, n55111, n55112, n55113, n55114,
         n55115, n55116, n55117, n55118, n55119, n55120, n55121, n55122,
         n55123, n55124, n55125, n55126, n55127, n55128, n55129, n55130,
         n55131, n55132, n55133, n55134, n55135, n55136, n55137, n55138,
         n55139, n55140, n55141, n55142, n55143, n55144, n55145, n55146,
         n55147, n55148, n55149, n55150, n55151, n55152, n55153, n55154,
         n55155, n55156, n55157, n55158, n55159, n55160, n55161, n55162,
         n55163, n55164, n55165, n55166, n55167, n55168, n55169, n55170,
         n55171, n55172, n55173, n55174, n55175, n55176, n55177, n55178,
         n55179, n55180, n55181, n55182, n55183, n55184, n55185, n55186,
         n55187, n55188, n55189, n55190, n55191, n55192, n55193, n55194,
         n55195, n55196, n55197, n55198, n55199, n55200, n55201, n55202,
         n55203, n55204, n55205, n55206, n55207, n55208, n55209, n55210,
         n55211, n55212, n55213, n55214, n55215, n55216, n55217, n55218,
         n55219, n55220, n55221, n55222, n55223, n55224, n55225, n55226,
         n55227, n55228, n55229, n55230, n55231, n55232, n55233, n55234,
         n55235, n55236, n55237, n55238, n55239, n55240, n55241, n55242,
         n55243, n55244, n55245, n55246, n55247, n55248, n55249, n55250,
         n55251, n55252, n55253, n55254, n55255, n55256, n55257, n55258,
         n55259, n55260, n55261, n55262, n55263, n55264, n55265, n55266,
         n55267, n55268, n55269, n55270, n55271, n55272, n55273, n55274,
         n55275, n55276, n55277, n55278, n55279, n55280, n55281, n55282,
         n55283, n55284, n55285, n55286, n55287, n55288, n55289, n55290,
         n55291, n55292, n55293, n55294, n55295, n55296, n55297, n55298,
         n55299, n55300, n55301, n55302, n55303, n55304, n55305, n55306,
         n55307, n55308, n55309, n55310, n55311, n55312, n55313, n55314,
         n55315, n55316, n55317, n55318, n55319, n55320, n55321, n55322,
         n55323, n55324, n55325, n55326, n55327, n55328, n55329, n55330,
         n55331, n55332, n55333, n55334, n55335, n55336, n55337, n55338,
         n55339, n55340, n55341, n55342, n55343, n55344, n55345, n55346,
         n55347, n55348, n55349, n55350, n55351, n55352, n55353, n55354,
         n55355, n55356, n55357, n55358, n55359, n55360, n55361, n55362,
         n55363, n55364, n55365, n55366, n55367, n55368, n55369, n55370,
         n55371, n55372, n55373, n55374, n55375, n55376, n55377, n55378,
         n55379, n55380, n55381, n55382, n55383, n55384, n55385, n55386,
         n55387, n55388, n55389, n55390, n55391, n55392, n55393, n55394,
         n55395, n55396, n55397, n55398, n55399, n55400, n55401, n55402,
         n55403, n55404, n55405, n55406, n55407, n55408, n55409, n55410,
         n55411, n55412, n55413, n55414, n55415, n55416, n55417, n55418,
         n55419, n55420, n55421, n55422, n55423, n55424, n55425, n55426,
         n55427, n55428, n55429, n55430, n55431, n55432, n55433, n55434,
         n55435, n55436, n55437, n55438, n55439, n55440, n55441, n55442,
         n55443, n55444, n55445, n55446, n55447, n55448, n55449, n55450,
         n55451, n55452, n55453, n55454, n55455, n55456, n55457, n55458,
         n55459, n55460, n55461, n55462, n55463, n55464, n55465, n55466,
         n55467, n55468, n55469, n55470, n55471, n55472, n55473, n55474,
         n55475, n55476, n55477, n55478, n55479, n55480, n55481, n55482,
         n55483, n55484, n55485, n55486, n55487, n55488, n55489, n55490,
         n55491, n55492, n55493, n55494, n55495, n55496, n55497, n55498,
         n55499, n55500, n55501, n55502, n55503, n55504, n55505, n55506,
         n55507, n55508, n55509, n55510, n55511, n55512, n55513, n55514,
         n55515, n55516, n55517, n55518, n55519, n55520, n55521, n55522,
         n55523, n55524, n55525, n55526, n55527, n55528, n55529, n55530,
         n55531, n55532, n55533, n55534, n55535, n55536, n55537, n55538,
         n55539, n55540, n55541, n55542, n55543, n55544, n55545, n55546,
         n55547, n55548, n55549, n55550, n55551, n55552, n55553, n55554,
         n55555, n55556, n55557, n55558, n55559, n55560, n55561, n55562,
         n55563, n55564, n55565, n55566, n55567, n55568, n55569, n55570,
         n55571, n55572, n55573, n55574, n55575, n55576, n55577, n55578,
         n55579, n55580, n55581, n55582, n55583, n55584, n55585, n55586,
         n55587, n55588, n55589, n55590, n55591, n55592, n55593, n55594,
         n55595, n55596, n55597, n55598, n55599, n55600, n55601, n55602,
         n55603, n55604, n55605, n55606, n55607, n55608, n55609, n55610,
         n55611, n55612, n55613, n55614, n55615, n55616, n55617, n55618,
         n55619, n55620, n55621, n55622, n55623, n55624, n55625, n55626,
         n55627, n55628, n55629, n55630, n55631, n55632, n55633, n55634,
         n55635, n55636, n55637, n55638, n55639, n55640, n55641, n55642,
         n55643, n55644, n55645, n55646, n55647, n55648, n55649, n55650,
         n55651, n55652, n55653, n55654, n55655, n55656, n55657, n55658,
         n55659, n55660, n55661, n55662, n55663, n55664, n55665, n55666,
         n55667, n55668, n55669, n55670, n55671, n55672, n55673, n55674,
         n55675, n55676, n55677, n55678, n55679, n55680, n55681, n55682,
         n55683, n55684, n55685, n55686, n55687, n55688, n55689, n55690,
         n55691, n55692, n55693, n55694, n55695, n55696, n55697, n55698,
         n55699, n55700, n55701, n55702, n55703, n55704, n55705, n55706,
         n55707, n55708, n55709, n55710, n55711, n55712, n55713, n55714,
         n55715, n55716, n55717, n55718, n55719, n55720, n55721, n55722,
         n55723, n55724, n55725, n55726, n55727, n55728, n55729, n55730,
         n55731, n55732, n55733, n55734, n55735, n55736, n55737, n55738,
         n55739, n55740, n55741, n55742, n55743, n55744, n55745, n55746,
         n55747, n55748, n55749, n55750, n55751, n55752, n55753, n55754,
         n55755, n55756, n55757, n55758, n55759, n55760, n55761, n55762,
         n55763, n55764, n55765, n55766, n55767, n55768, n55769, n55770,
         n55771, n55772, n55773, n55774, n55775, n55776, n55777, n55778,
         n55779, n55780, n55781, n55782, n55783, n55784, n55785, n55786,
         n55787, n55788, n55789, n55790, n55791, n55792, n55793, n55794,
         n55795, n55796, n55797, n55798, n55799, n55800, n55801, n55802,
         n55803, n55804, n55805, n55806, n55807, n55808, n55809, n55810,
         n55811, n55812, n55813, n55814, n55815, n55816, n55817, n55818,
         n55819, n55820, n55821, n55822, n55823, n55824, n55825, n55826,
         n55827, n55828, n55829, n55830, n55831, n55832, n55833, n55834,
         n55835, n55836, n55837, n55838, n55839, n55840, n55841, n55842,
         n55843, n55844, n55845, n55846, n55847, n55848, n55849, n55850,
         n55851, n55852, n55853, n55854, n55855, n55856, n55857, n55858,
         n55859, n55860, n55861, n55862, n55863, n55864, n55865, n55866,
         n55867, n55868, n55869, n55870, n55871, n55872, n55873, n55874,
         n55875, n55876, n55877, n55878, n55879, n55880, n55881, n55882,
         n55883, n55884, n55885, n55886, n55887, n55888, n55889, n55890,
         n55891, n55892, n55893, n55894, n55895, n55896, n55897, n55898,
         n55899, n55900, n55901, n55902, n55903, n55904, n55905, n55906,
         n55907, n55908, n55909, n55910, n55911, n55912, n55913, n55914,
         n55915, n55916, n55917, n55918, n55919, n55920, n55921, n55922,
         n55923, n55924, n55925, n55926, n55927, n55928, n55929, n55930,
         n55931, n55932, n55933, n55934, n55935, n55936, n55937, n55938,
         n55939, n55940, n55941, n55942, n55943, n55944, n55945, n55946,
         n55947, n55948, n55949, n55950, n55951, n55952, n55953, n55954,
         n55955, n55956, n55957, n55958, n55959, n55960, n55961, n55962,
         n55963, n55964, n55965, n55966, n55967, n55968, n55969, n55970,
         n55971, n55972, n55973, n55974, n55975, n55976, n55977, n55978,
         n55979, n55980, n55981, n55982, n55983, n55984, n55985, n55986,
         n55987, n55988, n55989, n55990, n55991, n55992, n55993, n55994,
         n55995, n55996, n55997, n55998, n55999, n56000, n56001, n56002,
         n56003, n56004, n56005, n56006, n56007, n56008, n56009, n56010,
         n56011, n56012, n56013, n56014, n56015, n56016, n56017, n56018,
         n56019, n56020, n56021, n56022, n56023, n56024, n56025, n56026,
         n56027, n56028, n56029, n56030, n56031, n56032, n56033, n56034,
         n56035, n56036, n56037, n56038, n56039, n56040, n56041, n56042,
         n56043, n56044, n56045, n56046, n56047, n56048, n56049, n56050,
         n56051, n56052, n56053, n56054, n56055, n56056, n56057, n56058,
         n56059, n56060, n56061, n56062, n56063, n56064, n56065, n56066,
         n56067, n56068, n56069, n56070, n56071, n56072, n56073, n56074,
         n56075, n56076, n56077, n56078, n56079, n56080, n56081, n56082,
         n56083, n56084, n56085, n56086, n56087, n56088, n56089, n56090,
         n56091, n56092, n56093, n56094, n56095, n56096, n56097, n56098,
         n56099, n56100, n56101, n56102, n56103, n56104, n56105, n56106,
         n56107, n56108, n56109, n56110, n56111, n56112, n56113, n56114,
         n56115, n56116, n56117, n56118, n56119, n56120, n56121, n56122,
         n56123, n56124, n56125, n56126, n56127, n56128, n56129, n56130,
         n56131, n56132, n56133, n56134, n56135, n56136, n56137, n56138,
         n56139, n56140, n56141, n56142, n56143, n56144, n56145, n56146,
         n56147, n56148, n56149, n56150, n56151, n56152, n56153, n56154,
         n56155, n56156, n56157, n56158, n56159, n56160, n56161, n56162,
         n56163, n56164, n56165, n56166, n56167, n56168, n56169, n56170,
         n56171, n56172, n56173, n56174, n56175, n56176, n56177, n56178,
         n56179, n56180, n56181, n56182, n56183, n56184, n56185, n56186,
         n56187, n56188, n56189, n56190, n56191, n56192, n56193, n56194,
         n56195, n56196, n56197, n56198, n56199, n56200, n56201, n56202,
         n56203, n56204, n56205, n56206, n56207, n56208, n56209, n56210,
         n56211, n56212, n56213, n56214, n56215, n56216, n56217, n56218,
         n56219, n56220, n56221, n56222, n56223, n56224, n56225, n56226,
         n56227, n56228, n56229, n56230, n56231, n56232, n56233, n56234,
         n56235, n56236, n56237, n56238, n56239, n56240, n56241, n56242,
         n56243, n56244, n56245, n56246, n56247, n56248, n56249, n56250,
         n56251, n56252, n56253, n56254, n56255, n56256, n56257, n56258,
         n56259, n56260, n56261, n56262, n56263, n56264, n56265, n56266,
         n56267, n56268, n56269, n56270, n56271, n56272, n56273, n56274,
         n56275, n56276, n56277, n56278, n56279, n56280, n56281, n56282,
         n56283, n56284, n56285, n56286, n56287, n56288, n56289, n56290,
         n56291, n56292, n56293, n56294, n56295, n56296, n56297, n56298,
         n56299, n56300, n56301, n56302, n56303, n56304, n56305, n56306,
         n56307, n56308, n56309, n56310, n56311, n56312, n56313, n56314,
         n56315, n56316, n56317, n56318, n56319, n56320, n56321, n56322,
         n56323, n56324, n56325, n56326, n56327, n56328, n56329, n56330,
         n56331, n56332, n56333, n56334, n56335, n56336, n56337, n56338,
         n56339, n56340, n56341, n56342, n56343, n56344, n56345, n56346,
         n56347, n56348, n56349, n56350, n56351, n56352, n56353, n56354,
         n56355, n56356, n56357, n56358, n56359, n56360, n56361, n56362,
         n56363, n56364, n56365, n56366, n56367, n56368, n56369, n56370,
         n56371, n56372, n56373, n56374, n56375, n56376, n56377, n56378,
         n56379, n56380, n56381, n56382, n56383, n56384, n56385, n56386,
         n56387, n56388, n56389, n56390, n56391, n56392, n56393, n56394,
         n56395, n56396, n56397, n56398, n56399, n56400, n56401, n56402,
         n56403, n56404, n56405, n56406, n56407, n56408, n56409, n56410,
         n56411, n56412, n56413, n56414, n56415, n56416, n56417, n56418,
         n56419, n56420, n56421, n56422, n56423, n56424, n56425, n56426,
         n56427, n56428, n56429, n56430, n56431, n56432, n56433, n56434,
         n56435, n56436, n56437, n56438, n56439, n56440, n56441, n56442,
         n56443, n56444, n56445, n56446, n56447, n56448, n56449, n56450,
         n56451, n56452, n56453, n56454, n56455, n56456, n56457, n56458,
         n56459, n56460, n56461, n56462, n56463, n56464, n56465, n56466,
         n56467, n56468, n56469, n56470, n56471, n56472, n56473, n56474,
         n56475, n56476, n56477, n56478, n56479, n56480, n56481, n56482,
         n56483, n56484, n56485, n56486, n56487, n56488, n56489, n56490,
         n56491, n56492, n56493, n56494, n56495, n56496, n56497, n56498,
         n56499, n56500, n56501, n56502, n56503, n56504, n56505, n56506,
         n56507, n56508, n56509, n56510, n56511, n56512, n56513, n56514,
         n56515, n56516, n56517, n56518, n56519, n56520, n56521, n56522,
         n56523, n56524, n56525, n56526, n56527, n56528, n56529, n56530,
         n56531, n56532, n56533, n56534, n56535, n56536, n56537, n56538,
         n56539, n56540, n56541, n56542, n56543, n56544, n56545, n56546,
         n56547, n56548, n56549, n56550, n56551, n56552, n56553, n56554,
         n56555, n56556, n56557, n56558, n56559, n56560, n56561, n56562,
         n56563, n56564, n56565, n56566, n56567, n56568, n56569, n56570,
         n56571, n56572, n56573, n56574, n56575, n56576, n56577, n56578,
         n56579, n56580, n56581, n56582, n56583, n56584, n56585, n56586,
         n56587, n56588, n56589, n56590, n56591, n56592, n56593, n56594,
         n56595, n56596, n56597, n56598, n56599, n56600, n56601, n56602,
         n56603, n56604, n56605, n56606, n56607, n56608, n56609, n56610,
         n56611, n56612, n56613, n56614, n56615, n56616, n56617, n56618,
         n56619, n56620, n56621, n56622, n56623, n56624, n56625, n56626,
         n56627, n56628, n56629, n56630, n56631, n56632, n56633, n56634,
         n56635, n56636, n56637, n56638, n56639, n56640, n56641, n56642,
         n56643, n56644, n56645, n56646, n56647, n56648, n56649, n56650,
         n56651, n56652, n56653, n56654, n56655, n56656, n56657, n56658,
         n56659, n56660, n56661, n56662, n56663, n56664, n56665, n56666,
         n56667, n56668, n56669, n56670, n56671, n56672, n56673, n56674,
         n56675, n56676, n56677, n56678, n56679, n56680, n56681, n56682,
         n56683, n56684, n56685, n56686, n56687, n56688, n56689, n56690,
         n56691, n56692, n56693, n56694, n56695, n56696, n56697, n56698,
         n56699, n56700, n56701, n56702, n56703, n56704, n56705, n56706,
         n56707, n56708, n56709, n56710, n56711, n56712, n56713, n56714,
         n56715, n56716, n56717, n56718, n56719, n56720, n56721, n56722,
         n56723, n56724, n56725, n56726, n56727, n56728, n56729, n56730,
         n56731, n56732, n56733, n56734, n56735, n56736, n56737, n56738,
         n56739, n56740, n56741, n56742, n56743, n56744, n56745, n56746,
         n56747, n56748, n56749, n56750, n56751, n56752, n56753, n56754,
         n56755, n56756, n56757, n56758, n56759, n56760, n56761, n56762,
         n56763, n56764, n56765, n56766, n56767, n56768, n56769, n56770,
         n56771, n56772, n56773, n56774, n56775, n56776, n56777, n56778,
         n56779, n56780, n56781, n56782, n56783, n56784, n56785, n56786,
         n56787, n56788, n56789, n56790, n56791, n56792, n56793, n56794,
         n56795, n56796, n56797, n56798, n56799, n56800, n56801, n56802,
         n56803, n56804, n56805, n56806, n56807, n56808, n56809, n56810,
         n56811, n56812, n56813, n56814, n56815, n56816, n56817, n56818,
         n56819, n56820, n56821, n56822, n56823, n56824, n56825, n56826,
         n56827, n56828, n56829, n56830, n56831, n56832, n56833, n56834,
         n56835, n56836, n56837, n56838, n56839, n56840, n56841, n56842,
         n56843, n56844, n56845, n56846, n56847, n56848, n56849, n56850,
         n56851, n56852, n56853, n56854, n56855, n56856, n56857, n56858,
         n56859, n56860, n56861, n56862, n56863, n56864, n56865, n56866,
         n56867, n56868, n56869, n56870, n56871, n56872, n56873, n56874,
         n56875, n56876, n56877, n56878, n56879, n56880, n56881, n56882,
         n56883, n56884, n56885, n56886, n56887, n56888, n56889, n56890,
         n56891, n56892, n56893, n56894, n56895, n56896, n56897, n56898,
         n56899, n56900, n56901, n56902, n56903, n56904, n56905, n56906,
         n56907, n56908, n56909, n56910, n56911, n56912, n56913, n56914,
         n56915, n56916, n56917, n56918, n56919, n56920, n56921, n56922,
         n56923, n56924, n56925, n56926, n56927, n56928, n56929, n56930,
         n56931, n56932, n56933, n56934, n56935, n56936, n56937, n56938,
         n56939, n56940, n56941, n56942, n56943, n56944, n56945, n56946,
         n56947, n56948, n56949, n56950, n56951, n56952, n56953, n56954,
         n56955, n56956, n56957, n56958, n56959, n56960, n56961, n56962,
         n56963, n56964, n56965, n56966, n56967, n56968, n56969, n56970,
         n56971, n56972, n56973, n56974, n56975, n56976, n56977, n56978,
         n56979, n56980, n56981, n56982, n56983, n56984, n56985, n56986,
         n56987, n56988, n56989, n56990, n56991, n56992, n56993, n56994,
         n56995, n56996, n56997, n56998, n56999, n57000, n57001, n57002,
         n57003, n57004, n57005, n57006, n57007, n57008, n57009, n57010,
         n57011, n57012, n57013, n57014, n57015, n57016, n57017, n57018,
         n57019, n57020, n57021, n57022, n57023, n57024, n57025, n57026,
         n57027, n57028, n57029, n57030, n57031, n57032, n57033, n57034,
         n57035, n57036, n57037, n57038, n57039, n57040, n57041, n57042,
         n57043, n57044, n57045, n57046, n57047, n57048, n57049, n57050,
         n57051, n57052, n57053, n57054, n57055, n57056, n57057, n57058,
         n57059, n57060, n57061, n57062, n57063, n57064, n57065, n57066,
         n57067, n57068, n57069, n57070, n57071, n57072, n57073, n57074,
         n57075, n57076, n57077, n57078, n57079, n57080, n57081, n57082,
         n57083, n57084, n57085, n57086, n57087, n57088, n57089, n57090,
         n57091, n57092, n57093, n57094, n57095, n57096, n57097, n57098,
         n57099, n57100, n57101, n57102, n57103, n57104, n57105, n57106,
         n57107, n57108, n57109, n57110, n57111, n57112, n57113, n57114,
         n57115, n57116, n57117, n57118, n57119, n57120, n57121, n57122,
         n57123, n57124, n57125, n57126, n57127, n57128, n57129, n57130,
         n57131, n57132, n57133, n57134, n57135, n57136, n57137, n57138,
         n57139, n57140, n57141, n57142, n57143, n57144, n57145, n57146,
         n57147, n57148, n57149, n57150, n57151, n57152, n57153, n57154,
         n57155, n57156, n57157, n57158, n57159, n57160, n57161, n57162,
         n57163, n57164, n57165, n57166, n57167, n57168, n57169, n57170,
         n57171, n57172, n57173, n57174, n57175, n57176, n57177, n57178,
         n57179, n57180, n57181, n57182, n57183, n57184, n57185, n57186,
         n57187, n57188, n57189, n57190, n57191, n57192, n57193, n57194,
         n57195, n57196, n57197, n57198, n57199, n57200, n57201, n57202,
         n57203, n57204, n57205, n57206, n57207, n57208, n57209, n57210,
         n57211, n57212, n57213, n57214, n57215, n57216, n57217, n57218,
         n57219, n57220, n57221, n57222, n57223, n57224, n57225, n57226,
         n57227, n57228, n57229, n57230, n57231, n57232, n57233, n57234,
         n57235, n57236, n57237, n57238, n57239, n57240, n57241, n57242,
         n57243, n57244, n57245, n57246, n57247, n57248, n57249, n57250,
         n57251, n57252, n57253, n57254, n57255, n57256, n57257, n57258,
         n57259, n57260, n57261, n57262, n57263, n57264, n57265, n57266,
         n57267, n57268, n57269, n57270, n57271, n57272, n57273, n57274,
         n57275, n57276, n57277, n57278, n57279, n57280, n57281, n57282,
         n57283, n57284, n57285, n57286, n57287, n57288, n57289, n57290,
         n57291, n57292, n57293, n57294, n57295, n57296, n57297, n57298,
         n57299, n57300, n57301, n57302, n57303, n57304, n57305, n57306,
         n57307, n57308, n57309, n57310, n57311, n57312, n57313, n57314,
         n57315, n57316, n57317, n57318, n57319, n57320, n57321, n57322,
         n57323, n57324, n57325, n57326, n57327, n57328, n57329, n57330,
         n57331, n57332, n57333, n57334, n57335, n57336, n57337, n57338,
         n57339, n57340, n57341, n57342, n57343, n57344, n57345, n57346,
         n57347, n57348, n57349, n57350, n57351, n57352, n57353, n57354,
         n57355, n57356, n57357, n57358, n57359, n57360, n57361, n57362,
         n57363, n57364, n57365, n57366, n57367, n57368, n57369, n57370,
         n57371, n57372, n57373, n57374, n57375, n57376, n57377, n57378,
         n57379, n57380, n57381, n57382, n57383, n57384, n57385, n57386,
         n57387, n57388, n57389, n57390, n57391, n57392, n57393, n57394,
         n57395, n57396, n57397, n57398, n57399, n57400, n57401, n57402,
         n57403, n57404, n57405, n57406, n57407, n57408, n57409, n57410,
         n57411, n57412, n57413, n57414, n57415, n57416, n57417, n57418,
         n57419, n57420, n57421, n57422, n57423, n57424, n57425, n57426,
         n57427, n57428, n57429, n57430, n57431, n57432, n57433, n57434,
         n57435, n57436, n57437, n57438, n57439, n57440, n57441, n57442,
         n57443, n57444, n57445, n57446, n57447, n57448, n57449, n57450,
         n57451, n57452, n57453, n57454, n57455, n57456, n57457, n57458,
         n57459, n57460, n57461, n57462, n57463, n57464, n57465, n57466,
         n57467, n57468, n57469, n57470, n57471, n57472, n57473, n57474,
         n57475, n57476, n57477, n57478, n57479, n57480, n57481, n57482,
         n57483, n57484, n57485, n57486, n57487, n57488, n57489, n57490,
         n57491, n57492, n57493, n57494, n57495, n57496, n57497, n57498,
         n57499, n57500, n57501, n57502, n57503, n57504, n57505, n57506,
         n57507, n57508, n57509, n57510, n57511, n57512, n57513, n57514,
         n57515, n57516, n57517, n57518, n57519, n57520, n57521, n57522,
         n57523, n57524, n57525, n57526, n57527, n57528, n57529, n57530,
         n57531, n57532, n57533, n57534, n57535, n57536, n57537, n57538,
         n57539, n57540, n57541, n57542, n57543, n57544, n57545, n57546,
         n57547, n57548, n57549, n57550, n57551, n57552, n57553, n57554,
         n57555, n57556, n57557, n57558, n57559, n57560, n57561, n57562,
         n57563, n57564, n57565, n57566, n57567, n57568, n57569, n57570,
         n57571, n57572, n57573, n57574, n57575, n57576, n57577, n57578,
         n57579, n57580, n57581, n57582, n57583, n57584, n57585, n57586,
         n57587, n57588, n57589, n57590, n57591, n57592, n57593, n57594,
         n57595, n57596, n57597, n57598, n57599, n57600, n57601, n57602,
         n57603, n57604, n57605, n57606, n57607, n57608, n57609, n57610,
         n57611, n57612, n57613, n57614, n57615, n57616, n57617, n57618,
         n57619, n57620, n57621, n57622, n57623, n57624, n57625, n57626,
         n57627, n57628, n57629, n57630, n57631, n57632, n57633, n57634,
         n57635, n57636, n57637, n57638, n57639, n57640, n57641, n57642,
         n57643, n57644, n57645, n57646, n57647, n57648, n57649, n57650,
         n57651, n57652, n57653, n57654, n57655, n57656, n57657, n57658,
         n57659, n57660, n57661, n57662, n57663, n57664, n57665, n57666,
         n57667, n57668, n57669, n57670, n57671, n57672, n57673, n57674,
         n57675, n57676, n57677, n57678, n57679, n57680, n57681, n57682,
         n57683, n57684, n57685, n57686, n57687, n57688, n57689, n57690,
         n57691, n57692, n57693, n57694, n57695, n57696, n57697, n57698,
         n57699, n57700, n57701, n57702, n57703, n57704, n57705, n57706,
         n57707, n57708, n57709, n57710, n57711, n57712, n57713, n57714,
         n57715, n57716, n57717, n57718, n57719, n57720, n57721, n57722,
         n57723, n57724, n57725, n57726, n57727, n57728, n57729, n57730,
         n57731, n57732, n57733, n57734, n57735, n57736, n57737, n57738,
         n57739, n57740, n57741, n57742, n57743, n57744, n57745, n57746,
         n57747, n57748, n57749, n57750, n57751, n57752, n57753, n57754,
         n57755, n57756, n57757, n57758, n57759, n57760, n57761, n57762,
         n57763, n57764, n57765, n57766, n57767, n57768, n57769, n57770,
         n57771, n57772, n57773, n57774, n57775, n57776, n57777, n57778,
         n57779, n57780, n57781, n57782, n57783, n57784, n57785, n57786,
         n57787, n57788, n57789, n57790, n57791, n57792, n57793, n57794,
         n57795, n57796, n57797, n57798, n57799, n57800, n57801, n57802,
         n57803, n57804, n57805, n57806, n57807, n57808, n57809, n57810,
         n57811, n57812, n57813, n57814, n57815, n57816, n57817, n57818,
         n57819, n57820, n57821, n57822, n57823, n57824, n57825, n57826,
         n57827, n57828, n57829, n57830, n57831, n57832, n57833, n57834,
         n57835, n57836, n57837, n57838, n57839, n57840, n57841, n57842,
         n57843, n57844, n57845, n57846, n57847, n57848, n57849, n57850,
         n57851, n57852, n57853, n57854, n57855, n57856, n57857, n57858,
         n57859, n57860, n57861, n57862, n57863, n57864, n57865, n57866,
         n57867, n57868, n57869, n57870, n57871, n57872, n57873, n57874,
         n57875, n57876, n57877, n57878, n57879, n57880, n57881, n57882,
         n57883, n57884, n57885, n57886, n57887, n57888, n57889, n57890,
         n57891, n57892, n57893, n57894, n57895, n57896, n57897, n57898,
         n57899, n57900, n57901, n57902, n57903, n57904, n57905, n57906,
         n57907, n57908, n57909, n57910, n57911, n57912, n57913, n57914,
         n57915, n57916, n57917, n57918, n57919, n57920, n57921, n57922,
         n57923, n57924, n57925, n57926, n57927, n57928, n57929, n57930,
         n57931, n57932, n57933, n57934, n57935, n57936, n57937, n57938,
         n57939, n57940, n57941, n57942, n57943, n57944, n57945, n57946,
         n57947, n57948, n57949, n57950, n57951, n57952, n57953, n57954,
         n57955, n57956, n57957, n57958, n57959, n57960, n57961, n57962,
         n57963, n57964, n57965, n57966, n57967, n57968, n57969, n57970,
         n57971, n57972, n57973, n57974, n57975, n57976, n57977, n57978,
         n57979, n57980, n57981, n57982, n57983, n57984, n57985, n57986,
         n57987, n57988, n57989, n57990, n57991, n57992, n57993, n57994,
         n57995, n57996, n57997, n57998, n57999, n58000, n58001, n58002,
         n58003, n58004, n58005, n58006, n58007, n58008, n58009, n58010,
         n58011, n58012, n58013, n58014, n58015, n58016, n58017, n58018,
         n58019, n58020, n58021, n58022, n58023, n58024, n58025, n58026,
         n58027, n58028, n58029, n58030, n58031, n58032, n58033, n58034,
         n58035, n58036, n58037, n58038, n58039, n58040, n58041, n58042,
         n58043, n58044, n58045, n58046, n58047, n58048, n58049, n58050,
         n58051, n58052, n58053, n58054, n58055, n58056, n58057, n58058,
         n58059, n58060, n58061, n58062, n58063, n58064, n58065, n58066,
         n58067, n58068, n58069, n58070, n58071, n58072, n58073, n58074,
         n58075, n58076, n58077, n58078, n58079, n58080, n58081, n58082,
         n58083, n58084, n58085, n58086, n58087, n58088, n58089, n58090,
         n58091, n58092, n58093, n58094, n58095, n58096, n58097, n58098,
         n58099, n58100, n58101, n58102, n58103, n58104, n58105, n58106,
         n58107, n58108, n58109, n58110, n58111, n58112, n58113, n58114,
         n58115, n58116, n58117, n58118, n58119, n58120, n58121, n58122,
         n58123, n58124, n58125, n58126, n58127, n58128, n58129, n58130,
         n58131, n58132, n58133, n58134, n58135, n58136, n58137, n58138,
         n58139, n58140, n58141, n58142, n58143, n58144, n58145, n58146,
         n58147, n58148, n58149, n58150, n58151, n58152, n58153, n58154,
         n58155, n58156, n58157, n58158, n58159, n58160, n58161, n58162,
         n58163, n58164, n58165, n58166, n58167, n58168, n58169, n58170,
         n58171, n58172, n58173, n58174, n58175, n58176, n58177, n58178,
         n58179, n58180, n58181, n58182, n58183, n58184, n58185, n58186,
         n58187, n58188, n58189, n58190, n58191, n58192, n58193, n58194,
         n58195, n58196, n58197, n58198, n58199, n58200, n58201, n58202,
         n58203, n58204, n58205, n58206, n58207, n58208, n58209, n58210,
         n58211, n58212, n58213, n58214, n58215, n58216, n58217, n58218,
         n58219, n58220, n58221, n58222, n58223, n58224, n58225, n58226,
         n58227, n58228, n58229, n58230, n58231, n58232, n58233, n58234,
         n58235, n58236, n58237, n58238, n58239, n58240, n58241, n58242,
         n58243, n58244, n58245, n58246, n58247, n58248, n58249, n58250,
         n58251, n58252, n58253, n58254, n58255, n58256, n58257, n58258,
         n58259, n58260, n58261, n58262, n58263, n58264, n58265, n58266,
         n58267, n58268, n58269, n58270, n58271, n58272, n58273, n58274,
         n58275, n58276, n58277, n58278, n58279, n58280, n58281, n58282,
         n58283, n58284, n58285, n58286, n58287, n58288, n58289, n58290,
         n58291, n58292, n58293, n58294, n58295, n58296, n58297, n58298,
         n58299, n58300, n58301, n58302, n58303, n58304, n58305, n58306,
         n58307, n58308, n58309, n58310, n58311, n58312, n58313, n58314,
         n58315, n58316, n58317, n58318, n58319, n58320, n58321, n58322,
         n58323, n58324, n58325, n58326, n58327, n58328, n58329, n58330,
         n58331, n58332, n58333, n58334, n58335, n58336, n58337, n58338,
         n58339, n58340, n58341, n58342, n58343, n58344, n58345, n58346,
         n58347, n58348, n58349, n58350, n58351, n58352, n58353, n58354,
         n58355, n58356, n58357, n58358, n58359, n58360, n58361, n58362,
         n58363, n58364, n58365, n58366, n58367, n58368, n58369, n58370,
         n58371, n58372, n58373, n58374, n58375, n58376, n58377, n58378,
         n58379, n58380, n58381, n58382, n58383, n58384, n58385, n58386,
         n58387, n58388, n58389, n58390, n58391, n58392, n58393, n58394,
         n58395, n58396, n58397, n58398, n58399, n58400, n58401, n58402,
         n58403, n58404, n58405, n58406, n58407, n58408, n58409, n58410,
         n58411, n58412, n58413, n58414, n58415, n58416, n58417, n58418,
         n58419, n58420, n58421, n58422, n58423, n58424, n58425, n58426,
         n58427, n58428, n58429, n58430, n58431, n58432, n58433, n58434,
         n58435, n58436, n58437, n58438, n58439, n58440, n58441, n58442,
         n58443, n58444, n58445, n58446, n58447, n58448, n58449, n58450,
         n58451, n58452, n58453, n58454, n58455, n58456, n58457, n58458,
         n58459, n58460, n58461, n58462, n58463, n58464, n58465, n58466,
         n58467, n58468, n58469, n58470, n58471, n58472, n58473, n58474,
         n58475, n58476, n58477, n58478, n58479, n58480, n58481, n58482,
         n58483, n58484, n58485, n58486, n58487, n58488, n58489, n58490,
         n58491, n58492, n58493, n58494, n58495, n58496, n58497, n58498,
         n58499, n58500, n58501, n58502, n58503, n58504, n58505, n58506,
         n58507, n58508, n58509, n58510, n58511, n58512, n58513, n58514,
         n58515, n58516, n58517, n58518, n58519, n58520, n58521, n58522,
         n58523, n58524, n58525, n58526, n58527, n58528, n58529, n58530,
         n58531, n58532, n58533, n58534, n58535, n58536, n58537, n58538,
         n58539, n58540, n58541, n58542, n58543, n58544, n58545, n58546,
         n58547, n58548, n58549, n58550, n58551, n58552, n58553, n58554,
         n58555, n58556, n58557, n58558, n58559, n58560, n58561, n58562,
         n58563, n58564, n58565, n58566, n58567, n58568, n58569, n58570,
         n58571, n58572, n58573, n58574, n58575, n58576, n58577, n58578,
         n58579, n58580, n58581, n58582, n58583, n58584, n58585, n58586,
         n58587, n58588, n58589, n58590, n58591, n58592, n58593, n58594,
         n58595, n58596, n58597, n58598, n58599, n58600, n58601, n58602,
         n58603, n58604, n58605, n58606, n58607, n58608, n58609, n58610,
         n58611, n58612, n58613, n58614, n58615, n58616, n58617, n58618,
         n58619, n58620, n58621, n58622, n58623, n58624, n58625, n58626,
         n58627, n58628, n58629, n58630, n58631, n58632, n58633, n58634,
         n58635, n58636, n58637, n58638, n58639, n58640, n58641, n58642,
         n58643, n58644, n58645, n58646, n58647, n58648, n58649, n58650,
         n58651, n58652, n58653, n58654, n58655, n58656, n58657, n58658,
         n58659, n58660, n58661, n58662, n58663, n58664, n58665, n58666,
         n58667, n58668, n58669, n58670, n58671, n58672, n58673, n58674,
         n58675, n58676, n58677, n58678, n58679, n58680, n58681, n58682,
         n58683, n58684, n58685, n58686, n58687, n58688, n58689, n58690,
         n58691, n58692, n58693, n58694, n58695, n58696, n58697, n58698,
         n58699, n58700, n58701, n58702, n58703, n58704, n58705, n58706,
         n58707, n58708, n58709, n58710, n58711, n58712, n58713, n58714,
         n58715, n58716, n58717, n58718;

  NOR U35632 ( .A(n32612), .B(n32614), .Z(n24435) );
  XOR U35633 ( .A(n32614), .B(n32613), .Z(n24436) );
  NOR U35634 ( .A(n32615), .B(n24436), .Z(n24437) );
  NOR U35635 ( .A(n24435), .B(n24437), .Z(n24438) );
  IV U35636 ( .A(n24438), .Z(n24439) );
  NOR U35637 ( .A(n32610), .B(n24439), .Z(n24440) );
  NOR U35638 ( .A(n32611), .B(n24439), .Z(n24441) );
  NOR U35639 ( .A(n24440), .B(n24441), .Z(n35971) );
  IV U35640 ( .A(n32602), .Z(n24442) );
  NOR U35641 ( .A(n32602), .B(n32601), .Z(n24443) );
  NOR U35642 ( .A(n32600), .B(n24442), .Z(n24444) );
  NOR U35643 ( .A(n32603), .B(n24444), .Z(n24445) );
  NOR U35644 ( .A(n24443), .B(n24445), .Z(n35974) );
  IV U35645 ( .A(n45995), .Z(n24446) );
  IV U35646 ( .A(n45997), .Z(n24447) );
  NOR U35647 ( .A(n24447), .B(n24446), .Z(n24448) );
  NOR U35648 ( .A(n45997), .B(n45995), .Z(n24449) );
  NOR U35649 ( .A(n45996), .B(n24449), .Z(n24450) );
  NOR U35650 ( .A(n24448), .B(n24450), .Z(n49546) );
  NOR U35651 ( .A(n49769), .B(n49768), .Z(n24451) );
  NOR U35652 ( .A(n49770), .B(n24451), .Z(n24452) );
  IV U35653 ( .A(n24452), .Z(n49773) );
  IV U35654 ( .A(n53542), .Z(n24453) );
  IV U35655 ( .A(n53544), .Z(n24454) );
  IV U35656 ( .A(n53539), .Z(n24455) );
  NOR U35657 ( .A(n53539), .B(n53540), .Z(n24456) );
  NOR U35658 ( .A(n53538), .B(n24455), .Z(n24457) );
  NOR U35659 ( .A(n53541), .B(n24457), .Z(n24458) );
  NOR U35660 ( .A(n24456), .B(n24458), .Z(n24459) );
  NOR U35661 ( .A(n24453), .B(n24454), .Z(n24460) );
  NOR U35662 ( .A(n24460), .B(n24459), .Z(n56618) );
  NOR U35663 ( .A(n57338), .B(n57339), .Z(n24461) );
  IV U35664 ( .A(n57340), .Z(n24462) );
  NOR U35665 ( .A(n24461), .B(n24462), .Z(n24463) );
  NOR U35666 ( .A(n57337), .B(n57336), .Z(n24464) );
  NOR U35667 ( .A(n57340), .B(n24464), .Z(n24465) );
  NOR U35668 ( .A(n24463), .B(n24465), .Z(n24466) );
  IV U35669 ( .A(n24466), .Z(n57353) );
  IV U35670 ( .A(n57428), .Z(n24467) );
  IV U35671 ( .A(n57433), .Z(n24468) );
  NOR U35672 ( .A(n57434), .B(n24468), .Z(n24469) );
  IV U35673 ( .A(n57430), .Z(n24470) );
  IV U35674 ( .A(n57432), .Z(n24471) );
  NOR U35675 ( .A(n57432), .B(n24470), .Z(n24472) );
  NOR U35676 ( .A(n57431), .B(n24472), .Z(n24473) );
  NOR U35677 ( .A(n57430), .B(n24471), .Z(n24474) );
  NOR U35678 ( .A(n24473), .B(n24474), .Z(n24475) );
  NOR U35679 ( .A(n24469), .B(n24475), .Z(n24476) );
  NOR U35680 ( .A(n57429), .B(n24467), .Z(n24477) );
  XOR U35681 ( .A(n24476), .B(n24477), .Z(n57435) );
  IV U35682 ( .A(n58020), .Z(n24478) );
  NOR U35683 ( .A(n58023), .B(n58022), .Z(n24479) );
  NOR U35684 ( .A(n24478), .B(n58021), .Z(n24480) );
  NOR U35685 ( .A(n24479), .B(n24480), .Z(n24481) );
  NOR U35686 ( .A(n58025), .B(n58024), .Z(n24482) );
  XOR U35687 ( .A(n58026), .B(n58025), .Z(n24483) );
  NOR U35688 ( .A(n58028), .B(n24483), .Z(n24484) );
  NOR U35689 ( .A(n24482), .B(n24484), .Z(n24485) );
  NOR U35690 ( .A(n24485), .B(n58027), .Z(n24486) );
  XOR U35691 ( .A(n24481), .B(n24486), .Z(n24487) );
  IV U35692 ( .A(n24487), .Z(n58029) );
  IV U35693 ( .A(n55807), .Z(n24488) );
  NOR U35694 ( .A(n55808), .B(n55807), .Z(n24489) );
  NOR U35695 ( .A(n55808), .B(n55806), .Z(n24490) );
  XOR U35696 ( .A(n55809), .B(n24490), .Z(n24491) );
  NOR U35697 ( .A(n24488), .B(n24491), .Z(n24492) );
  NOR U35698 ( .A(n24489), .B(n24492), .Z(n55810) );
  IV U35699 ( .A(n58341), .Z(n24493) );
  NOR U35700 ( .A(n58344), .B(n58343), .Z(n24494) );
  NOR U35701 ( .A(n58345), .B(n24494), .Z(n24495) );
  NOR U35702 ( .A(n24493), .B(n58342), .Z(n24496) );
  NOR U35703 ( .A(n24496), .B(n24495), .Z(n58346) );
  NOR U35704 ( .A(n54914), .B(n54913), .Z(n24497) );
  NOR U35705 ( .A(n54916), .B(n24497), .Z(n24498) );
  IV U35706 ( .A(n24498), .Z(n54912) );
  IV U35707 ( .A(x[1023]), .Z(n24499) );
  XOR U35708 ( .A(n24499), .B(y[1023]), .Z(n55074) );
  XOR U35709 ( .A(x[1022]), .B(y[1022]), .Z(n55038) );
  XOR U35710 ( .A(x[1021]), .B(y[1021]), .Z(n55009) );
  XOR U35711 ( .A(x[1020]), .B(y[1020]), .Z(n54983) );
  XOR U35712 ( .A(x[1019]), .B(y[1019]), .Z(n54955) );
  XOR U35713 ( .A(x[1018]), .B(y[1018]), .Z(n54932) );
  XOR U35714 ( .A(x[1017]), .B(y[1017]), .Z(n48092) );
  XOR U35715 ( .A(x[1016]), .B(y[1016]), .Z(n48064) );
  XOR U35716 ( .A(x[1015]), .B(y[1015]), .Z(n44677) );
  XOR U35717 ( .A(x[1014]), .B(y[1014]), .Z(n44659) );
  XOR U35718 ( .A(x[1013]), .B(y[1013]), .Z(n44643) );
  XOR U35719 ( .A(x[1012]), .B(y[1012]), .Z(n44615) );
  XOR U35720 ( .A(x[1011]), .B(y[1011]), .Z(n44597) );
  XOR U35721 ( .A(x[1010]), .B(y[1010]), .Z(n44572) );
  XOR U35722 ( .A(x[1009]), .B(y[1009]), .Z(n44554) );
  XOR U35723 ( .A(x[1008]), .B(y[1008]), .Z(n37936) );
  XOR U35724 ( .A(x[1007]), .B(y[1007]), .Z(n37930) );
  XOR U35725 ( .A(x[1006]), .B(y[1006]), .Z(n37926) );
  XOR U35726 ( .A(x[1005]), .B(y[1005]), .Z(n37909) );
  XOR U35727 ( .A(x[1004]), .B(y[1004]), .Z(n37901) );
  XOR U35728 ( .A(x[1003]), .B(y[1003]), .Z(n37889) );
  XOR U35729 ( .A(x[1002]), .B(y[1002]), .Z(n37870) );
  XOR U35730 ( .A(x[1001]), .B(y[1001]), .Z(n37858) );
  XOR U35731 ( .A(x[1000]), .B(y[1000]), .Z(n37839) );
  XOR U35732 ( .A(x[999]), .B(y[999]), .Z(n37819) );
  XOR U35733 ( .A(x[998]), .B(y[998]), .Z(n37824) );
  XOR U35734 ( .A(x[997]), .B(y[997]), .Z(n37798) );
  XOR U35735 ( .A(x[996]), .B(y[996]), .Z(n37791) );
  XOR U35736 ( .A(x[995]), .B(y[995]), .Z(n34385) );
  XOR U35737 ( .A(x[994]), .B(y[994]), .Z(n34379) );
  XOR U35738 ( .A(x[993]), .B(y[993]), .Z(n34372) );
  XOR U35739 ( .A(x[992]), .B(y[992]), .Z(n31185) );
  XOR U35740 ( .A(x[991]), .B(y[991]), .Z(n28069) );
  XOR U35741 ( .A(x[990]), .B(y[990]), .Z(n28066) );
  XOR U35742 ( .A(x[989]), .B(y[989]), .Z(n37962) );
  XOR U35743 ( .A(x[988]), .B(y[988]), .Z(n28060) );
  IV U35744 ( .A(n28060), .Z(n28062) );
  XOR U35745 ( .A(x[987]), .B(y[987]), .Z(n24500) );
  IV U35746 ( .A(n24500), .Z(n28053) );
  XOR U35747 ( .A(x[986]), .B(y[986]), .Z(n28044) );
  XOR U35748 ( .A(x[985]), .B(y[985]), .Z(n24502) );
  XOR U35749 ( .A(x[984]), .B(y[984]), .Z(n28039) );
  XOR U35750 ( .A(x[983]), .B(y[983]), .Z(n24508) );
  XOR U35751 ( .A(x[982]), .B(y[982]), .Z(n24505) );
  XOR U35752 ( .A(x[981]), .B(y[981]), .Z(n24511) );
  XOR U35753 ( .A(x[980]), .B(y[980]), .Z(n28032) );
  XOR U35754 ( .A(x[979]), .B(y[979]), .Z(n28029) );
  XOR U35755 ( .A(x[978]), .B(y[978]), .Z(n24514) );
  XOR U35756 ( .A(x[977]), .B(y[977]), .Z(n24520) );
  XOR U35757 ( .A(x[976]), .B(y[976]), .Z(n24517) );
  XOR U35758 ( .A(x[975]), .B(y[975]), .Z(n28024) );
  XOR U35759 ( .A(x[974]), .B(y[974]), .Z(n28021) );
  XOR U35760 ( .A(x[973]), .B(y[973]), .Z(n24526) );
  XOR U35761 ( .A(x[972]), .B(y[972]), .Z(n24523) );
  XOR U35762 ( .A(x[971]), .B(y[971]), .Z(n24532) );
  XOR U35763 ( .A(x[970]), .B(y[970]), .Z(n24529) );
  XOR U35764 ( .A(x[969]), .B(y[969]), .Z(n24538) );
  XOR U35765 ( .A(x[968]), .B(y[968]), .Z(n24535) );
  XOR U35766 ( .A(x[967]), .B(y[967]), .Z(n28017) );
  XOR U35767 ( .A(x[966]), .B(y[966]), .Z(n28014) );
  XOR U35768 ( .A(x[965]), .B(y[965]), .Z(n28011) );
  XOR U35769 ( .A(x[964]), .B(y[964]), .Z(n28008) );
  XOR U35770 ( .A(x[963]), .B(y[963]), .Z(n28004) );
  XOR U35771 ( .A(x[962]), .B(y[962]), .Z(n28001) );
  XOR U35772 ( .A(x[961]), .B(y[961]), .Z(n24541) );
  XOR U35773 ( .A(x[960]), .B(y[960]), .Z(n27995) );
  XOR U35774 ( .A(x[959]), .B(y[959]), .Z(n24544) );
  XOR U35775 ( .A(x[958]), .B(y[958]), .Z(n27988) );
  XOR U35776 ( .A(x[957]), .B(y[957]), .Z(n27985) );
  XOR U35777 ( .A(x[956]), .B(y[956]), .Z(n24547) );
  XOR U35778 ( .A(x[955]), .B(y[955]), .Z(n27981) );
  XOR U35779 ( .A(x[954]), .B(y[954]), .Z(n27978) );
  XOR U35780 ( .A(x[953]), .B(y[953]), .Z(n27974) );
  XOR U35781 ( .A(x[952]), .B(y[952]), .Z(n27971) );
  XOR U35782 ( .A(x[951]), .B(y[951]), .Z(n27968) );
  XOR U35783 ( .A(x[950]), .B(y[950]), .Z(n27965) );
  XOR U35784 ( .A(x[949]), .B(y[949]), .Z(n27961) );
  XOR U35785 ( .A(x[948]), .B(y[948]), .Z(n27958) );
  XOR U35786 ( .A(x[947]), .B(y[947]), .Z(n27954) );
  XOR U35787 ( .A(x[946]), .B(y[946]), .Z(n27951) );
  XOR U35788 ( .A(x[945]), .B(y[945]), .Z(n27947) );
  XOR U35789 ( .A(x[944]), .B(y[944]), .Z(n27944) );
  XOR U35790 ( .A(x[943]), .B(y[943]), .Z(n24553) );
  XOR U35791 ( .A(x[942]), .B(y[942]), .Z(n24550) );
  XOR U35792 ( .A(x[941]), .B(y[941]), .Z(n24559) );
  XOR U35793 ( .A(x[940]), .B(y[940]), .Z(n24556) );
  XOR U35794 ( .A(x[939]), .B(y[939]), .Z(n24565) );
  XOR U35795 ( .A(x[938]), .B(y[938]), .Z(n24562) );
  XOR U35796 ( .A(x[937]), .B(y[937]), .Z(n24571) );
  XOR U35797 ( .A(x[936]), .B(y[936]), .Z(n24568) );
  XOR U35798 ( .A(x[935]), .B(y[935]), .Z(n27939) );
  XOR U35799 ( .A(x[934]), .B(y[934]), .Z(n27936) );
  XOR U35800 ( .A(x[933]), .B(y[933]), .Z(n27932) );
  XOR U35801 ( .A(x[932]), .B(y[932]), .Z(n27929) );
  XOR U35802 ( .A(x[931]), .B(y[931]), .Z(n24575) );
  XOR U35803 ( .A(x[930]), .B(y[930]), .Z(n24581) );
  XOR U35804 ( .A(x[929]), .B(y[929]), .Z(n24578) );
  XOR U35805 ( .A(x[928]), .B(y[928]), .Z(n27916) );
  XOR U35806 ( .A(x[927]), .B(y[927]), .Z(n27912) );
  XOR U35807 ( .A(x[926]), .B(y[926]), .Z(n27920) );
  XOR U35808 ( .A(x[925]), .B(y[925]), .Z(n27908) );
  XOR U35809 ( .A(x[924]), .B(y[924]), .Z(n27905) );
  XOR U35810 ( .A(x[923]), .B(y[923]), .Z(n24587) );
  XOR U35811 ( .A(x[922]), .B(y[922]), .Z(n24584) );
  XOR U35812 ( .A(x[921]), .B(y[921]), .Z(n27901) );
  XOR U35813 ( .A(x[920]), .B(y[920]), .Z(n27898) );
  XOR U35814 ( .A(x[919]), .B(y[919]), .Z(n24593) );
  XOR U35815 ( .A(x[918]), .B(y[918]), .Z(n24590) );
  XOR U35816 ( .A(x[917]), .B(y[917]), .Z(n27895) );
  XOR U35817 ( .A(x[916]), .B(y[916]), .Z(n27892) );
  XOR U35818 ( .A(x[915]), .B(y[915]), .Z(n24599) );
  XOR U35819 ( .A(x[914]), .B(y[914]), .Z(n24596) );
  XOR U35820 ( .A(x[913]), .B(y[913]), .Z(n27888) );
  XOR U35821 ( .A(x[912]), .B(y[912]), .Z(n27885) );
  XOR U35822 ( .A(x[911]), .B(y[911]), .Z(n27881) );
  XOR U35823 ( .A(x[910]), .B(y[910]), .Z(n27878) );
  XOR U35824 ( .A(x[909]), .B(y[909]), .Z(n27874) );
  XOR U35825 ( .A(x[908]), .B(y[908]), .Z(n27871) );
  XOR U35826 ( .A(x[907]), .B(y[907]), .Z(n24602) );
  XOR U35827 ( .A(x[906]), .B(y[906]), .Z(n27867) );
  XOR U35828 ( .A(x[905]), .B(y[905]), .Z(n27864) );
  XOR U35829 ( .A(x[904]), .B(y[904]), .Z(n27860) );
  XOR U35830 ( .A(x[903]), .B(y[903]), .Z(n27857) );
  XOR U35831 ( .A(x[902]), .B(y[902]), .Z(n24605) );
  XOR U35832 ( .A(x[901]), .B(y[901]), .Z(n24611) );
  XOR U35833 ( .A(x[900]), .B(y[900]), .Z(n24608) );
  XOR U35834 ( .A(x[899]), .B(y[899]), .Z(n27852) );
  XOR U35835 ( .A(x[898]), .B(y[898]), .Z(n27849) );
  XOR U35836 ( .A(x[897]), .B(y[897]), .Z(n24617) );
  XOR U35837 ( .A(x[896]), .B(y[896]), .Z(n24614) );
  XOR U35838 ( .A(x[895]), .B(y[895]), .Z(n24623) );
  XOR U35839 ( .A(x[894]), .B(y[894]), .Z(n24620) );
  XOR U35840 ( .A(x[893]), .B(y[893]), .Z(n24629) );
  XOR U35841 ( .A(x[892]), .B(y[892]), .Z(n24626) );
  XOR U35842 ( .A(x[891]), .B(y[891]), .Z(n24632) );
  XOR U35843 ( .A(x[890]), .B(y[890]), .Z(n27842) );
  XOR U35844 ( .A(x[889]), .B(y[889]), .Z(n27839) );
  XOR U35845 ( .A(x[888]), .B(y[888]), .Z(n24635) );
  XOR U35846 ( .A(x[887]), .B(y[887]), .Z(n24641) );
  XOR U35847 ( .A(x[886]), .B(y[886]), .Z(n24638) );
  XOR U35848 ( .A(x[885]), .B(y[885]), .Z(n27836) );
  XOR U35849 ( .A(x[884]), .B(y[884]), .Z(n27833) );
  XOR U35850 ( .A(x[883]), .B(y[883]), .Z(n24647) );
  XOR U35851 ( .A(x[882]), .B(y[882]), .Z(n24644) );
  XOR U35852 ( .A(x[881]), .B(y[881]), .Z(n24653) );
  XOR U35853 ( .A(x[880]), .B(y[880]), .Z(n24650) );
  XOR U35854 ( .A(x[879]), .B(y[879]), .Z(n24659) );
  XOR U35855 ( .A(x[878]), .B(y[878]), .Z(n24656) );
  XOR U35856 ( .A(x[877]), .B(y[877]), .Z(n24665) );
  XOR U35857 ( .A(x[876]), .B(y[876]), .Z(n24662) );
  XOR U35858 ( .A(x[875]), .B(y[875]), .Z(n24671) );
  XOR U35859 ( .A(x[874]), .B(y[874]), .Z(n24668) );
  XOR U35860 ( .A(x[873]), .B(y[873]), .Z(n24674) );
  XOR U35861 ( .A(x[872]), .B(y[872]), .Z(n27826) );
  XOR U35862 ( .A(x[871]), .B(y[871]), .Z(n27823) );
  XOR U35863 ( .A(x[870]), .B(y[870]), .Z(n27819) );
  XOR U35864 ( .A(x[869]), .B(y[869]), .Z(n27816) );
  XOR U35865 ( .A(x[868]), .B(y[868]), .Z(n27812) );
  XOR U35866 ( .A(x[867]), .B(y[867]), .Z(n27809) );
  XOR U35867 ( .A(x[866]), .B(y[866]), .Z(n24678) );
  XOR U35868 ( .A(x[865]), .B(y[865]), .Z(n27805) );
  XOR U35869 ( .A(x[864]), .B(y[864]), .Z(n27802) );
  XOR U35870 ( .A(x[863]), .B(y[863]), .Z(n27798) );
  XOR U35871 ( .A(x[862]), .B(y[862]), .Z(n27795) );
  XOR U35872 ( .A(x[861]), .B(y[861]), .Z(n24681) );
  XOR U35873 ( .A(x[860]), .B(y[860]), .Z(n27792) );
  XOR U35874 ( .A(x[859]), .B(y[859]), .Z(n27789) );
  XOR U35875 ( .A(x[858]), .B(y[858]), .Z(n27785) );
  XOR U35876 ( .A(x[857]), .B(y[857]), .Z(n27782) );
  XOR U35877 ( .A(x[856]), .B(y[856]), .Z(n24684) );
  XOR U35878 ( .A(x[855]), .B(y[855]), .Z(n24690) );
  XOR U35879 ( .A(x[854]), .B(y[854]), .Z(n24687) );
  XOR U35880 ( .A(x[853]), .B(y[853]), .Z(n24696) );
  XOR U35881 ( .A(x[852]), .B(y[852]), .Z(n24693) );
  XOR U35882 ( .A(x[851]), .B(y[851]), .Z(n24702) );
  XOR U35883 ( .A(x[850]), .B(y[850]), .Z(n24699) );
  XOR U35884 ( .A(x[849]), .B(y[849]), .Z(n24706) );
  XOR U35885 ( .A(x[848]), .B(y[848]), .Z(n24712) );
  XOR U35886 ( .A(x[847]), .B(y[847]), .Z(n24709) );
  XOR U35887 ( .A(x[846]), .B(y[846]), .Z(n24718) );
  XOR U35888 ( .A(x[845]), .B(y[845]), .Z(n24715) );
  XOR U35889 ( .A(x[844]), .B(y[844]), .Z(n27775) );
  XOR U35890 ( .A(x[843]), .B(y[843]), .Z(n27772) );
  XOR U35891 ( .A(x[842]), .B(y[842]), .Z(n24721) );
  XOR U35892 ( .A(x[841]), .B(y[841]), .Z(n27763) );
  XOR U35893 ( .A(x[840]), .B(y[840]), .Z(n27760) );
  XOR U35894 ( .A(x[839]), .B(y[839]), .Z(n24727) );
  XOR U35895 ( .A(x[838]), .B(y[838]), .Z(n24724) );
  XOR U35896 ( .A(x[837]), .B(y[837]), .Z(n24733) );
  XOR U35897 ( .A(x[836]), .B(y[836]), .Z(n24730) );
  XOR U35898 ( .A(x[835]), .B(y[835]), .Z(n24739) );
  XOR U35899 ( .A(x[834]), .B(y[834]), .Z(n24736) );
  XOR U35900 ( .A(x[833]), .B(y[833]), .Z(n24745) );
  XOR U35901 ( .A(x[832]), .B(y[832]), .Z(n24742) );
  XOR U35902 ( .A(x[831]), .B(y[831]), .Z(n24748) );
  XOR U35903 ( .A(x[830]), .B(y[830]), .Z(n27752) );
  XOR U35904 ( .A(x[829]), .B(y[829]), .Z(n27749) );
  XOR U35905 ( .A(x[828]), .B(y[828]), .Z(n27736) );
  XOR U35906 ( .A(x[827]), .B(y[827]), .Z(n27733) );
  XOR U35907 ( .A(x[826]), .B(y[826]), .Z(n24751) );
  XOR U35908 ( .A(x[825]), .B(y[825]), .Z(n24757) );
  XOR U35909 ( .A(x[824]), .B(y[824]), .Z(n24754) );
  XOR U35910 ( .A(x[823]), .B(y[823]), .Z(n27727) );
  XOR U35911 ( .A(x[822]), .B(y[822]), .Z(n27724) );
  XOR U35912 ( .A(x[821]), .B(y[821]), .Z(n24763) );
  XOR U35913 ( .A(x[820]), .B(y[820]), .Z(n24760) );
  XOR U35914 ( .A(x[819]), .B(y[819]), .Z(n24767) );
  XOR U35915 ( .A(x[818]), .B(y[818]), .Z(n24773) );
  XOR U35916 ( .A(x[817]), .B(y[817]), .Z(n24770) );
  XOR U35917 ( .A(x[816]), .B(y[816]), .Z(n24779) );
  XOR U35918 ( .A(x[815]), .B(y[815]), .Z(n24776) );
  XOR U35919 ( .A(x[814]), .B(y[814]), .Z(n24785) );
  XOR U35920 ( .A(x[813]), .B(y[813]), .Z(n24782) );
  XOR U35921 ( .A(x[812]), .B(y[812]), .Z(n24791) );
  XOR U35922 ( .A(x[811]), .B(y[811]), .Z(n24788) );
  XOR U35923 ( .A(x[810]), .B(y[810]), .Z(n24794) );
  XOR U35924 ( .A(x[809]), .B(y[809]), .Z(n24801) );
  XOR U35925 ( .A(x[808]), .B(y[808]), .Z(n24798) );
  XOR U35926 ( .A(x[807]), .B(y[807]), .Z(n24807) );
  XOR U35927 ( .A(x[806]), .B(y[806]), .Z(n24804) );
  XOR U35928 ( .A(x[805]), .B(y[805]), .Z(n24813) );
  XOR U35929 ( .A(x[804]), .B(y[804]), .Z(n24810) );
  XOR U35930 ( .A(x[803]), .B(y[803]), .Z(n24819) );
  XOR U35931 ( .A(x[802]), .B(y[802]), .Z(n24816) );
  XOR U35932 ( .A(x[801]), .B(y[801]), .Z(n24822) );
  XOR U35933 ( .A(x[800]), .B(y[800]), .Z(n27711) );
  XOR U35934 ( .A(x[799]), .B(y[799]), .Z(n24825) );
  XOR U35935 ( .A(x[798]), .B(y[798]), .Z(n24831) );
  XOR U35936 ( .A(x[797]), .B(y[797]), .Z(n24828) );
  XOR U35937 ( .A(x[796]), .B(y[796]), .Z(n24837) );
  XOR U35938 ( .A(x[795]), .B(y[795]), .Z(n24834) );
  XOR U35939 ( .A(x[794]), .B(y[794]), .Z(n24840) );
  XOR U35940 ( .A(x[793]), .B(y[793]), .Z(n27705) );
  XOR U35941 ( .A(x[792]), .B(y[792]), .Z(n27702) );
  XOR U35942 ( .A(x[791]), .B(y[791]), .Z(n27699) );
  XOR U35943 ( .A(x[790]), .B(y[790]), .Z(n27696) );
  XOR U35944 ( .A(x[789]), .B(y[789]), .Z(n27692) );
  XOR U35945 ( .A(x[788]), .B(y[788]), .Z(n27689) );
  XOR U35946 ( .A(x[787]), .B(y[787]), .Z(n24846) );
  XOR U35947 ( .A(x[786]), .B(y[786]), .Z(n24843) );
  XOR U35948 ( .A(x[785]), .B(y[785]), .Z(n27684) );
  XOR U35949 ( .A(x[784]), .B(y[784]), .Z(n27681) );
  XOR U35950 ( .A(x[783]), .B(y[783]), .Z(n24852) );
  XOR U35951 ( .A(x[782]), .B(y[782]), .Z(n24849) );
  XOR U35952 ( .A(x[781]), .B(y[781]), .Z(n24858) );
  XOR U35953 ( .A(x[780]), .B(y[780]), .Z(n24855) );
  XOR U35954 ( .A(x[779]), .B(y[779]), .Z(n24864) );
  XOR U35955 ( .A(x[778]), .B(y[778]), .Z(n24861) );
  XOR U35956 ( .A(x[777]), .B(y[777]), .Z(n24871) );
  XOR U35957 ( .A(x[776]), .B(y[776]), .Z(n24868) );
  XOR U35958 ( .A(x[775]), .B(y[775]), .Z(n24878) );
  XOR U35959 ( .A(x[774]), .B(y[774]), .Z(n24875) );
  XOR U35960 ( .A(x[773]), .B(y[773]), .Z(n24884) );
  XOR U35961 ( .A(x[772]), .B(y[772]), .Z(n24881) );
  XOR U35962 ( .A(x[771]), .B(y[771]), .Z(n24890) );
  XOR U35963 ( .A(x[770]), .B(y[770]), .Z(n24887) );
  XOR U35964 ( .A(x[769]), .B(y[769]), .Z(n27676) );
  XOR U35965 ( .A(x[768]), .B(y[768]), .Z(n27673) );
  XOR U35966 ( .A(x[767]), .B(y[767]), .Z(n24893) );
  XOR U35967 ( .A(x[766]), .B(y[766]), .Z(n27669) );
  XOR U35968 ( .A(x[765]), .B(y[765]), .Z(n27666) );
  XOR U35969 ( .A(x[764]), .B(y[764]), .Z(n24899) );
  XOR U35970 ( .A(x[763]), .B(y[763]), .Z(n24896) );
  XOR U35971 ( .A(x[762]), .B(y[762]), .Z(n24902) );
  XOR U35972 ( .A(x[761]), .B(y[761]), .Z(n27662) );
  XOR U35973 ( .A(x[760]), .B(y[760]), .Z(n27659) );
  XOR U35974 ( .A(x[759]), .B(y[759]), .Z(n27655) );
  XOR U35975 ( .A(x[758]), .B(y[758]), .Z(n27652) );
  XOR U35976 ( .A(x[757]), .B(y[757]), .Z(n24908) );
  XOR U35977 ( .A(x[756]), .B(y[756]), .Z(n24905) );
  XOR U35978 ( .A(x[755]), .B(y[755]), .Z(n24914) );
  XOR U35979 ( .A(x[754]), .B(y[754]), .Z(n24911) );
  XOR U35980 ( .A(x[753]), .B(y[753]), .Z(n24920) );
  XOR U35981 ( .A(x[752]), .B(y[752]), .Z(n24917) );
  XOR U35982 ( .A(x[751]), .B(y[751]), .Z(n24926) );
  XOR U35983 ( .A(x[750]), .B(y[750]), .Z(n24923) );
  XOR U35984 ( .A(x[749]), .B(y[749]), .Z(n27646) );
  XOR U35985 ( .A(x[748]), .B(y[748]), .Z(n27643) );
  XOR U35986 ( .A(x[747]), .B(y[747]), .Z(n27639) );
  XOR U35987 ( .A(x[746]), .B(y[746]), .Z(n27636) );
  XOR U35988 ( .A(x[745]), .B(y[745]), .Z(n24932) );
  XOR U35989 ( .A(x[744]), .B(y[744]), .Z(n24929) );
  XOR U35990 ( .A(x[743]), .B(y[743]), .Z(n24938) );
  XOR U35991 ( .A(x[742]), .B(y[742]), .Z(n24935) );
  XOR U35992 ( .A(x[741]), .B(y[741]), .Z(n24944) );
  XOR U35993 ( .A(x[740]), .B(y[740]), .Z(n24941) );
  XOR U35994 ( .A(x[739]), .B(y[739]), .Z(n24947) );
  XOR U35995 ( .A(x[738]), .B(y[738]), .Z(n24951) );
  XOR U35996 ( .A(x[737]), .B(y[737]), .Z(n27624) );
  XOR U35997 ( .A(x[736]), .B(y[736]), .Z(n27621) );
  XOR U35998 ( .A(x[735]), .B(y[735]), .Z(n24957) );
  XOR U35999 ( .A(x[734]), .B(y[734]), .Z(n24954) );
  XOR U36000 ( .A(x[733]), .B(y[733]), .Z(n24963) );
  XOR U36001 ( .A(x[732]), .B(y[732]), .Z(n24960) );
  XOR U36002 ( .A(x[731]), .B(y[731]), .Z(n24966) );
  XOR U36003 ( .A(x[730]), .B(y[730]), .Z(n27616) );
  XOR U36004 ( .A(x[729]), .B(y[729]), .Z(n27613) );
  XOR U36005 ( .A(x[728]), .B(y[728]), .Z(n24972) );
  XOR U36006 ( .A(x[727]), .B(y[727]), .Z(n24969) );
  XOR U36007 ( .A(x[726]), .B(y[726]), .Z(n27609) );
  XOR U36008 ( .A(x[725]), .B(y[725]), .Z(n27606) );
  XOR U36009 ( .A(x[724]), .B(y[724]), .Z(n24978) );
  XOR U36010 ( .A(x[723]), .B(y[723]), .Z(n24975) );
  XOR U36011 ( .A(x[722]), .B(y[722]), .Z(n27602) );
  XOR U36012 ( .A(x[721]), .B(y[721]), .Z(n27599) );
  XOR U36013 ( .A(x[720]), .B(y[720]), .Z(n24984) );
  XOR U36014 ( .A(x[719]), .B(y[719]), .Z(n24981) );
  XOR U36015 ( .A(x[718]), .B(y[718]), .Z(n24990) );
  XOR U36016 ( .A(x[717]), .B(y[717]), .Z(n24987) );
  XOR U36017 ( .A(x[716]), .B(y[716]), .Z(n24996) );
  XOR U36018 ( .A(x[715]), .B(y[715]), .Z(n24993) );
  XOR U36019 ( .A(x[714]), .B(y[714]), .Z(n25002) );
  XOR U36020 ( .A(x[713]), .B(y[713]), .Z(n24999) );
  XOR U36021 ( .A(x[712]), .B(y[712]), .Z(n27586) );
  XOR U36022 ( .A(x[711]), .B(y[711]), .Z(n25005) );
  XOR U36023 ( .A(x[710]), .B(y[710]), .Z(n27590) );
  XOR U36024 ( .A(x[709]), .B(y[709]), .Z(n25009) );
  XOR U36025 ( .A(x[708]), .B(y[708]), .Z(n25015) );
  XOR U36026 ( .A(x[707]), .B(y[707]), .Z(n25012) );
  XOR U36027 ( .A(x[706]), .B(y[706]), .Z(n25021) );
  XOR U36028 ( .A(x[705]), .B(y[705]), .Z(n25018) );
  XOR U36029 ( .A(x[704]), .B(y[704]), .Z(n25024) );
  XOR U36030 ( .A(x[703]), .B(y[703]), .Z(n25030) );
  XOR U36031 ( .A(x[702]), .B(y[702]), .Z(n25027) );
  XOR U36032 ( .A(x[701]), .B(y[701]), .Z(n25037) );
  XOR U36033 ( .A(x[700]), .B(y[700]), .Z(n25034) );
  XOR U36034 ( .A(x[699]), .B(y[699]), .Z(n27567) );
  XOR U36035 ( .A(x[698]), .B(y[698]), .Z(n27570) );
  XOR U36036 ( .A(x[697]), .B(y[697]), .Z(n25040) );
  XOR U36037 ( .A(x[696]), .B(y[696]), .Z(n27556) );
  XOR U36038 ( .A(x[695]), .B(y[695]), .Z(n25043) );
  XOR U36039 ( .A(x[694]), .B(y[694]), .Z(n27547) );
  XOR U36040 ( .A(x[693]), .B(y[693]), .Z(n25046) );
  XOR U36041 ( .A(x[692]), .B(y[692]), .Z(n27541) );
  XOR U36042 ( .A(x[691]), .B(y[691]), .Z(n27538) );
  XOR U36043 ( .A(x[690]), .B(y[690]), .Z(n27533) );
  XOR U36044 ( .A(x[689]), .B(y[689]), .Z(n27530) );
  XOR U36045 ( .A(x[688]), .B(y[688]), .Z(n25049) );
  XOR U36046 ( .A(x[687]), .B(y[687]), .Z(n25055) );
  XOR U36047 ( .A(x[686]), .B(y[686]), .Z(n25052) );
  XOR U36048 ( .A(x[685]), .B(y[685]), .Z(n25061) );
  XOR U36049 ( .A(x[684]), .B(y[684]), .Z(n25058) );
  XOR U36050 ( .A(x[683]), .B(y[683]), .Z(n25067) );
  XOR U36051 ( .A(x[682]), .B(y[682]), .Z(n25064) );
  XOR U36052 ( .A(x[681]), .B(y[681]), .Z(n25073) );
  XOR U36053 ( .A(x[680]), .B(y[680]), .Z(n25070) );
  XOR U36054 ( .A(x[679]), .B(y[679]), .Z(n25079) );
  XOR U36055 ( .A(x[678]), .B(y[678]), .Z(n25076) );
  XOR U36056 ( .A(x[677]), .B(y[677]), .Z(n25082) );
  XOR U36057 ( .A(x[676]), .B(y[676]), .Z(n27521) );
  XOR U36058 ( .A(x[675]), .B(y[675]), .Z(n27518) );
  XOR U36059 ( .A(x[674]), .B(y[674]), .Z(n25085) );
  XOR U36060 ( .A(x[673]), .B(y[673]), .Z(n25091) );
  XOR U36061 ( .A(x[672]), .B(y[672]), .Z(n25088) );
  XOR U36062 ( .A(x[671]), .B(y[671]), .Z(n27513) );
  XOR U36063 ( .A(x[670]), .B(y[670]), .Z(n27510) );
  XOR U36064 ( .A(x[669]), .B(y[669]), .Z(n25094) );
  XOR U36065 ( .A(x[668]), .B(y[668]), .Z(n25100) );
  XOR U36066 ( .A(x[667]), .B(y[667]), .Z(n25097) );
  XOR U36067 ( .A(x[666]), .B(y[666]), .Z(n25103) );
  XOR U36068 ( .A(x[665]), .B(y[665]), .Z(n25109) );
  XOR U36069 ( .A(x[664]), .B(y[664]), .Z(n25106) );
  XOR U36070 ( .A(x[663]), .B(y[663]), .Z(n25115) );
  XOR U36071 ( .A(x[662]), .B(y[662]), .Z(n25112) );
  XOR U36072 ( .A(x[661]), .B(y[661]), .Z(n25121) );
  XOR U36073 ( .A(x[660]), .B(y[660]), .Z(n25118) );
  XOR U36074 ( .A(x[659]), .B(y[659]), .Z(n25127) );
  XOR U36075 ( .A(x[658]), .B(y[658]), .Z(n25124) );
  XOR U36076 ( .A(x[657]), .B(y[657]), .Z(n27501) );
  XOR U36077 ( .A(x[656]), .B(y[656]), .Z(n27498) );
  XOR U36078 ( .A(x[655]), .B(y[655]), .Z(n27486) );
  XOR U36079 ( .A(x[654]), .B(y[654]), .Z(n27482) );
  XOR U36080 ( .A(x[653]), .B(y[653]), .Z(n25130) );
  XOR U36081 ( .A(x[652]), .B(y[652]), .Z(n25133) );
  XOR U36082 ( .A(x[651]), .B(y[651]), .Z(n25140) );
  XOR U36083 ( .A(x[650]), .B(y[650]), .Z(n25137) );
  XOR U36084 ( .A(x[649]), .B(y[649]), .Z(n27478) );
  XOR U36085 ( .A(x[648]), .B(y[648]), .Z(n27475) );
  XOR U36086 ( .A(x[647]), .B(y[647]), .Z(n25146) );
  XOR U36087 ( .A(x[646]), .B(y[646]), .Z(n25143) );
  XOR U36088 ( .A(x[645]), .B(y[645]), .Z(n25152) );
  XOR U36089 ( .A(x[644]), .B(y[644]), .Z(n25149) );
  XOR U36090 ( .A(x[643]), .B(y[643]), .Z(n25158) );
  XOR U36091 ( .A(x[642]), .B(y[642]), .Z(n25155) );
  XOR U36092 ( .A(x[641]), .B(y[641]), .Z(n27470) );
  XOR U36093 ( .A(x[640]), .B(y[640]), .Z(n27467) );
  XOR U36094 ( .A(x[639]), .B(y[639]), .Z(n25164) );
  XOR U36095 ( .A(x[638]), .B(y[638]), .Z(n25161) );
  XOR U36096 ( .A(x[637]), .B(y[637]), .Z(n27464) );
  XOR U36097 ( .A(x[636]), .B(y[636]), .Z(n27461) );
  XOR U36098 ( .A(x[635]), .B(y[635]), .Z(n27458) );
  XOR U36099 ( .A(x[634]), .B(y[634]), .Z(n27455) );
  XOR U36100 ( .A(x[633]), .B(y[633]), .Z(n27451) );
  XOR U36101 ( .A(x[632]), .B(y[632]), .Z(n27448) );
  XOR U36102 ( .A(x[631]), .B(y[631]), .Z(n25170) );
  XOR U36103 ( .A(x[630]), .B(y[630]), .Z(n25167) );
  XOR U36104 ( .A(x[629]), .B(y[629]), .Z(n25176) );
  XOR U36105 ( .A(x[628]), .B(y[628]), .Z(n25173) );
  XOR U36106 ( .A(x[627]), .B(y[627]), .Z(n25182) );
  XOR U36107 ( .A(x[626]), .B(y[626]), .Z(n25179) );
  XOR U36108 ( .A(x[625]), .B(y[625]), .Z(n25185) );
  XOR U36109 ( .A(x[624]), .B(y[624]), .Z(n27441) );
  XOR U36110 ( .A(x[623]), .B(y[623]), .Z(n25188) );
  XOR U36111 ( .A(x[622]), .B(y[622]), .Z(n25194) );
  XOR U36112 ( .A(x[621]), .B(y[621]), .Z(n25191) );
  XOR U36113 ( .A(x[620]), .B(y[620]), .Z(n25200) );
  XOR U36114 ( .A(x[619]), .B(y[619]), .Z(n25197) );
  XOR U36115 ( .A(x[618]), .B(y[618]), .Z(n25203) );
  XOR U36116 ( .A(x[617]), .B(y[617]), .Z(n25209) );
  XOR U36117 ( .A(x[616]), .B(y[616]), .Z(n25206) );
  XOR U36118 ( .A(x[615]), .B(y[615]), .Z(n25215) );
  XOR U36119 ( .A(x[614]), .B(y[614]), .Z(n25212) );
  XOR U36120 ( .A(x[613]), .B(y[613]), .Z(n25218) );
  XOR U36121 ( .A(x[612]), .B(y[612]), .Z(n27430) );
  XOR U36122 ( .A(x[611]), .B(y[611]), .Z(n27427) );
  XOR U36123 ( .A(x[610]), .B(y[610]), .Z(n25221) );
  XOR U36124 ( .A(x[609]), .B(y[609]), .Z(n25227) );
  XOR U36125 ( .A(x[608]), .B(y[608]), .Z(n25224) );
  XOR U36126 ( .A(x[607]), .B(y[607]), .Z(n25230) );
  XOR U36127 ( .A(x[606]), .B(y[606]), .Z(n27416) );
  XOR U36128 ( .A(x[605]), .B(y[605]), .Z(n25233) );
  XOR U36129 ( .A(x[604]), .B(y[604]), .Z(n27410) );
  XOR U36130 ( .A(x[603]), .B(y[603]), .Z(n27407) );
  XOR U36131 ( .A(x[602]), .B(y[602]), .Z(n27404) );
  XOR U36132 ( .A(x[601]), .B(y[601]), .Z(n27401) );
  XOR U36133 ( .A(x[600]), .B(y[600]), .Z(n27397) );
  XOR U36134 ( .A(x[599]), .B(y[599]), .Z(n27394) );
  XOR U36135 ( .A(x[598]), .B(y[598]), .Z(n25237) );
  XOR U36136 ( .A(x[597]), .B(y[597]), .Z(n25243) );
  XOR U36137 ( .A(x[596]), .B(y[596]), .Z(n25240) );
  XOR U36138 ( .A(x[595]), .B(y[595]), .Z(n27389) );
  XOR U36139 ( .A(x[594]), .B(y[594]), .Z(n27386) );
  XOR U36140 ( .A(x[593]), .B(y[593]), .Z(n27382) );
  XOR U36141 ( .A(x[592]), .B(y[592]), .Z(n27379) );
  XOR U36142 ( .A(x[591]), .B(y[591]), .Z(n27375) );
  XOR U36143 ( .A(x[590]), .B(y[590]), .Z(n27372) );
  XOR U36144 ( .A(x[589]), .B(y[589]), .Z(n25246) );
  XOR U36145 ( .A(x[588]), .B(y[588]), .Z(n27362) );
  XOR U36146 ( .A(x[587]), .B(y[587]), .Z(n27356) );
  XOR U36147 ( .A(x[586]), .B(y[586]), .Z(n27353) );
  XOR U36148 ( .A(x[585]), .B(y[585]), .Z(n25252) );
  XOR U36149 ( .A(x[584]), .B(y[584]), .Z(n25249) );
  XOR U36150 ( .A(x[583]), .B(y[583]), .Z(n27350) );
  XOR U36151 ( .A(x[582]), .B(y[582]), .Z(n27347) );
  XOR U36152 ( .A(x[581]), .B(y[581]), .Z(n25258) );
  XOR U36153 ( .A(x[580]), .B(y[580]), .Z(n25255) );
  XOR U36154 ( .A(x[579]), .B(y[579]), .Z(n27343) );
  XOR U36155 ( .A(x[578]), .B(y[578]), .Z(n27340) );
  XOR U36156 ( .A(x[577]), .B(y[577]), .Z(n27336) );
  XOR U36157 ( .A(x[576]), .B(y[576]), .Z(n27333) );
  XOR U36158 ( .A(x[575]), .B(y[575]), .Z(n27329) );
  XOR U36159 ( .A(x[574]), .B(y[574]), .Z(n27326) );
  XOR U36160 ( .A(x[573]), .B(y[573]), .Z(n25264) );
  XOR U36161 ( .A(x[572]), .B(y[572]), .Z(n25261) );
  XOR U36162 ( .A(x[571]), .B(y[571]), .Z(n27322) );
  XOR U36163 ( .A(x[570]), .B(y[570]), .Z(n27319) );
  XOR U36164 ( .A(x[569]), .B(y[569]), .Z(n25270) );
  XOR U36165 ( .A(x[568]), .B(y[568]), .Z(n25267) );
  XOR U36166 ( .A(x[567]), .B(y[567]), .Z(n25276) );
  XOR U36167 ( .A(x[566]), .B(y[566]), .Z(n25273) );
  XOR U36168 ( .A(x[565]), .B(y[565]), .Z(n25282) );
  XOR U36169 ( .A(x[564]), .B(y[564]), .Z(n25279) );
  XOR U36170 ( .A(x[563]), .B(y[563]), .Z(n25285) );
  XOR U36171 ( .A(x[562]), .B(y[562]), .Z(n27307) );
  XOR U36172 ( .A(x[561]), .B(y[561]), .Z(n27301) );
  XOR U36173 ( .A(x[560]), .B(y[560]), .Z(n27298) );
  XOR U36174 ( .A(x[559]), .B(y[559]), .Z(n25291) );
  XOR U36175 ( .A(x[558]), .B(y[558]), .Z(n25288) );
  XOR U36176 ( .A(x[557]), .B(y[557]), .Z(n25297) );
  XOR U36177 ( .A(x[556]), .B(y[556]), .Z(n25294) );
  XOR U36178 ( .A(x[555]), .B(y[555]), .Z(n25303) );
  XOR U36179 ( .A(x[554]), .B(y[554]), .Z(n25300) );
  XOR U36180 ( .A(x[553]), .B(y[553]), .Z(n25309) );
  XOR U36181 ( .A(x[552]), .B(y[552]), .Z(n25306) );
  XOR U36182 ( .A(x[551]), .B(y[551]), .Z(n25312) );
  XOR U36183 ( .A(x[550]), .B(y[550]), .Z(n25318) );
  XOR U36184 ( .A(x[549]), .B(y[549]), .Z(n25315) );
  XOR U36185 ( .A(x[548]), .B(y[548]), .Z(n25324) );
  XOR U36186 ( .A(x[547]), .B(y[547]), .Z(n25321) );
  XOR U36187 ( .A(x[546]), .B(y[546]), .Z(n25330) );
  XOR U36188 ( .A(x[545]), .B(y[545]), .Z(n25327) );
  XOR U36189 ( .A(x[544]), .B(y[544]), .Z(n27285) );
  XOR U36190 ( .A(x[543]), .B(y[543]), .Z(n25333) );
  XOR U36191 ( .A(x[542]), .B(y[542]), .Z(n27289) );
  XOR U36192 ( .A(x[541]), .B(y[541]), .Z(n27282) );
  XOR U36193 ( .A(x[540]), .B(y[540]), .Z(n27279) );
  XOR U36194 ( .A(x[539]), .B(y[539]), .Z(n25340) );
  XOR U36195 ( .A(x[538]), .B(y[538]), .Z(n25337) );
  XOR U36196 ( .A(x[537]), .B(y[537]), .Z(n27274) );
  XOR U36197 ( .A(x[536]), .B(y[536]), .Z(n27271) );
  XOR U36198 ( .A(x[535]), .B(y[535]), .Z(n25346) );
  XOR U36199 ( .A(x[534]), .B(y[534]), .Z(n25343) );
  XOR U36200 ( .A(x[533]), .B(y[533]), .Z(n27267) );
  XOR U36201 ( .A(x[532]), .B(y[532]), .Z(n27264) );
  XOR U36202 ( .A(x[531]), .B(y[531]), .Z(n25352) );
  XOR U36203 ( .A(x[530]), .B(y[530]), .Z(n25349) );
  XOR U36204 ( .A(x[529]), .B(y[529]), .Z(n25355) );
  XOR U36205 ( .A(x[528]), .B(y[528]), .Z(n27257) );
  XOR U36206 ( .A(x[527]), .B(y[527]), .Z(n25358) );
  XOR U36207 ( .A(x[526]), .B(y[526]), .Z(n27250) );
  XOR U36208 ( .A(x[525]), .B(y[525]), .Z(n27247) );
  XOR U36209 ( .A(x[524]), .B(y[524]), .Z(n25364) );
  XOR U36210 ( .A(x[523]), .B(y[523]), .Z(n25361) );
  XOR U36211 ( .A(x[522]), .B(y[522]), .Z(n25370) );
  XOR U36212 ( .A(x[521]), .B(y[521]), .Z(n25367) );
  XOR U36213 ( .A(x[520]), .B(y[520]), .Z(n25374) );
  XOR U36214 ( .A(x[519]), .B(y[519]), .Z(n27243) );
  XOR U36215 ( .A(x[518]), .B(y[518]), .Z(n27240) );
  XOR U36216 ( .A(x[517]), .B(y[517]), .Z(n27236) );
  XOR U36217 ( .A(x[516]), .B(y[516]), .Z(n27233) );
  XOR U36218 ( .A(x[515]), .B(y[515]), .Z(n25377) );
  XOR U36219 ( .A(x[514]), .B(y[514]), .Z(n25383) );
  XOR U36220 ( .A(x[513]), .B(y[513]), .Z(n25380) );
  XOR U36221 ( .A(x[512]), .B(y[512]), .Z(n25389) );
  XOR U36222 ( .A(x[511]), .B(y[511]), .Z(n25386) );
  XOR U36223 ( .A(x[510]), .B(y[510]), .Z(n25395) );
  XOR U36224 ( .A(x[509]), .B(y[509]), .Z(n25392) );
  XOR U36225 ( .A(x[508]), .B(y[508]), .Z(n25401) );
  XOR U36226 ( .A(x[507]), .B(y[507]), .Z(n25398) );
  XOR U36227 ( .A(x[506]), .B(y[506]), .Z(n25404) );
  XOR U36228 ( .A(x[505]), .B(y[505]), .Z(n25410) );
  XOR U36229 ( .A(x[504]), .B(y[504]), .Z(n25407) );
  XOR U36230 ( .A(x[503]), .B(y[503]), .Z(n25416) );
  XOR U36231 ( .A(x[502]), .B(y[502]), .Z(n25413) );
  XOR U36232 ( .A(x[501]), .B(y[501]), .Z(n25422) );
  XOR U36233 ( .A(x[500]), .B(y[500]), .Z(n25419) );
  XOR U36234 ( .A(x[499]), .B(y[499]), .Z(n25426) );
  XOR U36235 ( .A(x[498]), .B(y[498]), .Z(n25432) );
  XOR U36236 ( .A(x[497]), .B(y[497]), .Z(n25429) );
  XOR U36237 ( .A(x[496]), .B(y[496]), .Z(n25438) );
  XOR U36238 ( .A(x[495]), .B(y[495]), .Z(n25435) );
  XOR U36239 ( .A(x[494]), .B(y[494]), .Z(n25441) );
  XOR U36240 ( .A(x[493]), .B(y[493]), .Z(n25445) );
  XOR U36241 ( .A(x[492]), .B(y[492]), .Z(n27219) );
  XOR U36242 ( .A(x[491]), .B(y[491]), .Z(n27213) );
  XOR U36243 ( .A(x[490]), .B(y[490]), .Z(n27210) );
  XOR U36244 ( .A(x[489]), .B(y[489]), .Z(n25451) );
  XOR U36245 ( .A(x[488]), .B(y[488]), .Z(n25448) );
  XOR U36246 ( .A(x[487]), .B(y[487]), .Z(n25457) );
  XOR U36247 ( .A(x[486]), .B(y[486]), .Z(n25454) );
  XOR U36248 ( .A(x[485]), .B(y[485]), .Z(n25463) );
  XOR U36249 ( .A(x[484]), .B(y[484]), .Z(n25460) );
  XOR U36250 ( .A(x[483]), .B(y[483]), .Z(n25470) );
  XOR U36251 ( .A(x[482]), .B(y[482]), .Z(n25467) );
  XOR U36252 ( .A(x[481]), .B(y[481]), .Z(n25476) );
  XOR U36253 ( .A(x[480]), .B(y[480]), .Z(n25473) );
  XOR U36254 ( .A(x[479]), .B(y[479]), .Z(n27196) );
  XOR U36255 ( .A(x[478]), .B(y[478]), .Z(n25479) );
  XOR U36256 ( .A(x[477]), .B(y[477]), .Z(n27200) );
  XOR U36257 ( .A(x[476]), .B(y[476]), .Z(n25486) );
  XOR U36258 ( .A(x[475]), .B(y[475]), .Z(n25483) );
  XOR U36259 ( .A(x[474]), .B(y[474]), .Z(n25492) );
  XOR U36260 ( .A(x[473]), .B(y[473]), .Z(n25489) );
  XOR U36261 ( .A(x[472]), .B(y[472]), .Z(n25495) );
  XOR U36262 ( .A(x[471]), .B(y[471]), .Z(n27192) );
  XOR U36263 ( .A(x[470]), .B(y[470]), .Z(n27189) );
  XOR U36264 ( .A(x[469]), .B(y[469]), .Z(n25501) );
  XOR U36265 ( .A(x[468]), .B(y[468]), .Z(n25498) );
  XOR U36266 ( .A(x[467]), .B(y[467]), .Z(n25504) );
  XOR U36267 ( .A(x[466]), .B(y[466]), .Z(n25510) );
  XOR U36268 ( .A(x[465]), .B(y[465]), .Z(n25507) );
  XOR U36269 ( .A(x[464]), .B(y[464]), .Z(n25516) );
  XOR U36270 ( .A(x[463]), .B(y[463]), .Z(n25513) );
  XOR U36271 ( .A(x[462]), .B(y[462]), .Z(n27183) );
  XOR U36272 ( .A(x[461]), .B(y[461]), .Z(n27180) );
  XOR U36273 ( .A(x[460]), .B(y[460]), .Z(n25522) );
  XOR U36274 ( .A(x[459]), .B(y[459]), .Z(n25519) );
  XOR U36275 ( .A(x[458]), .B(y[458]), .Z(n25529) );
  XOR U36276 ( .A(x[457]), .B(y[457]), .Z(n25526) );
  XOR U36277 ( .A(x[456]), .B(y[456]), .Z(n27167) );
  XOR U36278 ( .A(x[455]), .B(y[455]), .Z(n25532) );
  XOR U36279 ( .A(x[454]), .B(y[454]), .Z(n27171) );
  XOR U36280 ( .A(x[453]), .B(y[453]), .Z(n25536) );
  XOR U36281 ( .A(x[452]), .B(y[452]), .Z(n27163) );
  XOR U36282 ( .A(x[451]), .B(y[451]), .Z(n27160) );
  XOR U36283 ( .A(x[450]), .B(y[450]), .Z(n27157) );
  XOR U36284 ( .A(x[449]), .B(y[449]), .Z(n27154) );
  XOR U36285 ( .A(x[448]), .B(y[448]), .Z(n27150) );
  XOR U36286 ( .A(x[447]), .B(y[447]), .Z(n27147) );
  XOR U36287 ( .A(x[446]), .B(y[446]), .Z(n25542) );
  XOR U36288 ( .A(x[445]), .B(y[445]), .Z(n25539) );
  XOR U36289 ( .A(x[444]), .B(y[444]), .Z(n25548) );
  XOR U36290 ( .A(x[443]), .B(y[443]), .Z(n25545) );
  XOR U36291 ( .A(x[442]), .B(y[442]), .Z(n25554) );
  XOR U36292 ( .A(x[441]), .B(y[441]), .Z(n25551) );
  XOR U36293 ( .A(x[440]), .B(y[440]), .Z(n25557) );
  XOR U36294 ( .A(x[439]), .B(y[439]), .Z(n27142) );
  XOR U36295 ( .A(x[438]), .B(y[438]), .Z(n27139) );
  XOR U36296 ( .A(x[437]), .B(y[437]), .Z(n25563) );
  XOR U36297 ( .A(x[436]), .B(y[436]), .Z(n25560) );
  XOR U36298 ( .A(x[435]), .B(y[435]), .Z(n25566) );
  XOR U36299 ( .A(x[434]), .B(y[434]), .Z(n27128) );
  XOR U36300 ( .A(x[433]), .B(y[433]), .Z(n25569) );
  XOR U36301 ( .A(x[432]), .B(y[432]), .Z(n27123) );
  XOR U36302 ( .A(x[431]), .B(y[431]), .Z(n27120) );
  XOR U36303 ( .A(x[430]), .B(y[430]), .Z(n25575) );
  XOR U36304 ( .A(x[429]), .B(y[429]), .Z(n25572) );
  XOR U36305 ( .A(x[428]), .B(y[428]), .Z(n27116) );
  XOR U36306 ( .A(x[427]), .B(y[427]), .Z(n27113) );
  XOR U36307 ( .A(x[426]), .B(y[426]), .Z(n25581) );
  XOR U36308 ( .A(x[425]), .B(y[425]), .Z(n25578) );
  XOR U36309 ( .A(x[424]), .B(y[424]), .Z(n27108) );
  XOR U36310 ( .A(x[423]), .B(y[423]), .Z(n27105) );
  XOR U36311 ( .A(x[422]), .B(y[422]), .Z(n25587) );
  XOR U36312 ( .A(x[421]), .B(y[421]), .Z(n25584) );
  XOR U36313 ( .A(x[420]), .B(y[420]), .Z(n25593) );
  XOR U36314 ( .A(x[419]), .B(y[419]), .Z(n25590) );
  XOR U36315 ( .A(x[418]), .B(y[418]), .Z(n25599) );
  XOR U36316 ( .A(x[417]), .B(y[417]), .Z(n25596) );
  XOR U36317 ( .A(x[416]), .B(y[416]), .Z(n27099) );
  XOR U36318 ( .A(x[415]), .B(y[415]), .Z(n27096) );
  XOR U36319 ( .A(x[414]), .B(y[414]), .Z(n25605) );
  XOR U36320 ( .A(x[413]), .B(y[413]), .Z(n25602) );
  XOR U36321 ( .A(x[412]), .B(y[412]), .Z(n25611) );
  XOR U36322 ( .A(x[411]), .B(y[411]), .Z(n25608) );
  XOR U36323 ( .A(x[410]), .B(y[410]), .Z(n27091) );
  XOR U36324 ( .A(x[409]), .B(y[409]), .Z(n27088) );
  XOR U36325 ( .A(x[408]), .B(y[408]), .Z(n27084) );
  XOR U36326 ( .A(x[407]), .B(y[407]), .Z(n27081) );
  XOR U36327 ( .A(x[406]), .B(y[406]), .Z(n27078) );
  XOR U36328 ( .A(x[405]), .B(y[405]), .Z(n27075) );
  XOR U36329 ( .A(x[404]), .B(y[404]), .Z(n27071) );
  XOR U36330 ( .A(x[403]), .B(y[403]), .Z(n27068) );
  XOR U36331 ( .A(x[402]), .B(y[402]), .Z(n25614) );
  XOR U36332 ( .A(x[401]), .B(y[401]), .Z(n25620) );
  XOR U36333 ( .A(x[400]), .B(y[400]), .Z(n25617) );
  XOR U36334 ( .A(x[399]), .B(y[399]), .Z(n27064) );
  XOR U36335 ( .A(x[398]), .B(y[398]), .Z(n27061) );
  XOR U36336 ( .A(x[397]), .B(y[397]), .Z(n27057) );
  XOR U36337 ( .A(x[396]), .B(y[396]), .Z(n27054) );
  XOR U36338 ( .A(x[395]), .B(y[395]), .Z(n27051) );
  XOR U36339 ( .A(x[394]), .B(y[394]), .Z(n27048) );
  XOR U36340 ( .A(x[393]), .B(y[393]), .Z(n25623) );
  XOR U36341 ( .A(x[392]), .B(y[392]), .Z(n25629) );
  XOR U36342 ( .A(x[391]), .B(y[391]), .Z(n25626) );
  XOR U36343 ( .A(x[390]), .B(y[390]), .Z(n27043) );
  XOR U36344 ( .A(x[389]), .B(y[389]), .Z(n27040) );
  XOR U36345 ( .A(x[388]), .B(y[388]), .Z(n25632) );
  XOR U36346 ( .A(x[387]), .B(y[387]), .Z(n27032) );
  XOR U36347 ( .A(x[386]), .B(y[386]), .Z(n25635) );
  XOR U36348 ( .A(x[385]), .B(y[385]), .Z(n27027) );
  XOR U36349 ( .A(x[384]), .B(y[384]), .Z(n27024) );
  XOR U36350 ( .A(x[383]), .B(y[383]), .Z(n25641) );
  XOR U36351 ( .A(x[382]), .B(y[382]), .Z(n25638) );
  XOR U36352 ( .A(x[381]), .B(y[381]), .Z(n27021) );
  XOR U36353 ( .A(x[380]), .B(y[380]), .Z(n27018) );
  XOR U36354 ( .A(x[379]), .B(y[379]), .Z(n27015) );
  XOR U36355 ( .A(x[378]), .B(y[378]), .Z(n27012) );
  XOR U36356 ( .A(x[377]), .B(y[377]), .Z(n25647) );
  XOR U36357 ( .A(x[376]), .B(y[376]), .Z(n25644) );
  XOR U36358 ( .A(x[375]), .B(y[375]), .Z(n25650) );
  XOR U36359 ( .A(x[374]), .B(y[374]), .Z(n25656) );
  XOR U36360 ( .A(x[373]), .B(y[373]), .Z(n25653) );
  XOR U36361 ( .A(x[372]), .B(y[372]), .Z(n26999) );
  XOR U36362 ( .A(x[371]), .B(y[371]), .Z(n26996) );
  XOR U36363 ( .A(x[370]), .B(y[370]), .Z(n26992) );
  XOR U36364 ( .A(x[369]), .B(y[369]), .Z(n26989) );
  XOR U36365 ( .A(x[368]), .B(y[368]), .Z(n26985) );
  XOR U36366 ( .A(x[367]), .B(y[367]), .Z(n26982) );
  XOR U36367 ( .A(x[366]), .B(y[366]), .Z(n26978) );
  XOR U36368 ( .A(x[365]), .B(y[365]), .Z(n26975) );
  XOR U36369 ( .A(x[364]), .B(y[364]), .Z(n26971) );
  XOR U36370 ( .A(x[363]), .B(y[363]), .Z(n26968) );
  XOR U36371 ( .A(x[362]), .B(y[362]), .Z(n25659) );
  XOR U36372 ( .A(x[361]), .B(y[361]), .Z(n26964) );
  XOR U36373 ( .A(x[360]), .B(y[360]), .Z(n26961) );
  XOR U36374 ( .A(x[359]), .B(y[359]), .Z(n26957) );
  XOR U36375 ( .A(x[358]), .B(y[358]), .Z(n26954) );
  XOR U36376 ( .A(x[357]), .B(y[357]), .Z(n25662) );
  XOR U36377 ( .A(x[356]), .B(y[356]), .Z(n26951) );
  XOR U36378 ( .A(x[355]), .B(y[355]), .Z(n26948) );
  XOR U36379 ( .A(x[354]), .B(y[354]), .Z(n26944) );
  XOR U36380 ( .A(x[353]), .B(y[353]), .Z(n26941) );
  XOR U36381 ( .A(x[352]), .B(y[352]), .Z(n25665) );
  XOR U36382 ( .A(x[351]), .B(y[351]), .Z(n25671) );
  XOR U36383 ( .A(x[350]), .B(y[350]), .Z(n25668) );
  XOR U36384 ( .A(x[349]), .B(y[349]), .Z(n26935) );
  XOR U36385 ( .A(x[348]), .B(y[348]), .Z(n26932) );
  XOR U36386 ( .A(x[347]), .B(y[347]), .Z(n26928) );
  XOR U36387 ( .A(x[346]), .B(y[346]), .Z(n26925) );
  XOR U36388 ( .A(x[345]), .B(y[345]), .Z(n26921) );
  XOR U36389 ( .A(x[344]), .B(y[344]), .Z(n26918) );
  XOR U36390 ( .A(x[343]), .B(y[343]), .Z(n25674) );
  XOR U36391 ( .A(x[342]), .B(y[342]), .Z(n26912) );
  XOR U36392 ( .A(x[341]), .B(y[341]), .Z(n25677) );
  XOR U36393 ( .A(x[340]), .B(y[340]), .Z(n25683) );
  XOR U36394 ( .A(x[339]), .B(y[339]), .Z(n25680) );
  XOR U36395 ( .A(x[338]), .B(y[338]), .Z(n25689) );
  XOR U36396 ( .A(x[337]), .B(y[337]), .Z(n25686) );
  XOR U36397 ( .A(x[336]), .B(y[336]), .Z(n25692) );
  XOR U36398 ( .A(x[335]), .B(y[335]), .Z(n26905) );
  XOR U36399 ( .A(x[334]), .B(y[334]), .Z(n26902) );
  XOR U36400 ( .A(x[333]), .B(y[333]), .Z(n25698) );
  XOR U36401 ( .A(x[332]), .B(y[332]), .Z(n25695) );
  XOR U36402 ( .A(x[331]), .B(y[331]), .Z(n25704) );
  XOR U36403 ( .A(x[330]), .B(y[330]), .Z(n25701) );
  XOR U36404 ( .A(x[329]), .B(y[329]), .Z(n25710) );
  XOR U36405 ( .A(x[328]), .B(y[328]), .Z(n25707) );
  XOR U36406 ( .A(x[327]), .B(y[327]), .Z(n25716) );
  XOR U36407 ( .A(x[326]), .B(y[326]), .Z(n25713) );
  XOR U36408 ( .A(x[325]), .B(y[325]), .Z(n26896) );
  XOR U36409 ( .A(x[324]), .B(y[324]), .Z(n26893) );
  XOR U36410 ( .A(x[323]), .B(y[323]), .Z(n25719) );
  XOR U36411 ( .A(x[322]), .B(y[322]), .Z(n25725) );
  XOR U36412 ( .A(x[321]), .B(y[321]), .Z(n25722) );
  XOR U36413 ( .A(x[320]), .B(y[320]), .Z(n25731) );
  XOR U36414 ( .A(x[319]), .B(y[319]), .Z(n25728) );
  XOR U36415 ( .A(x[318]), .B(y[318]), .Z(n25734) );
  XOR U36416 ( .A(x[317]), .B(y[317]), .Z(n26889) );
  XOR U36417 ( .A(x[316]), .B(y[316]), .Z(n26886) );
  XOR U36418 ( .A(x[315]), .B(y[315]), .Z(n26882) );
  XOR U36419 ( .A(x[314]), .B(y[314]), .Z(n26879) );
  XOR U36420 ( .A(x[313]), .B(y[313]), .Z(n26875) );
  XOR U36421 ( .A(x[312]), .B(y[312]), .Z(n26872) );
  XOR U36422 ( .A(x[311]), .B(y[311]), .Z(n25738) );
  XOR U36423 ( .A(x[310]), .B(y[310]), .Z(n25744) );
  XOR U36424 ( .A(x[309]), .B(y[309]), .Z(n25741) );
  XOR U36425 ( .A(x[308]), .B(y[308]), .Z(n26866) );
  XOR U36426 ( .A(x[307]), .B(y[307]), .Z(n26863) );
  XOR U36427 ( .A(x[306]), .B(y[306]), .Z(n26860) );
  XOR U36428 ( .A(x[305]), .B(y[305]), .Z(n26857) );
  XOR U36429 ( .A(x[304]), .B(y[304]), .Z(n26853) );
  XOR U36430 ( .A(x[303]), .B(y[303]), .Z(n26850) );
  XOR U36431 ( .A(x[302]), .B(y[302]), .Z(n26846) );
  XOR U36432 ( .A(x[301]), .B(y[301]), .Z(n26843) );
  XOR U36433 ( .A(x[300]), .B(y[300]), .Z(n26839) );
  XOR U36434 ( .A(x[299]), .B(y[299]), .Z(n26836) );
  XOR U36435 ( .A(x[298]), .B(y[298]), .Z(n25747) );
  XOR U36436 ( .A(x[297]), .B(y[297]), .Z(n26830) );
  XOR U36437 ( .A(x[296]), .B(y[296]), .Z(n25750) );
  XOR U36438 ( .A(x[295]), .B(y[295]), .Z(n26824) );
  XOR U36439 ( .A(x[294]), .B(y[294]), .Z(n26821) );
  XOR U36440 ( .A(x[293]), .B(y[293]), .Z(n25756) );
  XOR U36441 ( .A(x[292]), .B(y[292]), .Z(n25753) );
  XOR U36442 ( .A(x[291]), .B(y[291]), .Z(n25762) );
  XOR U36443 ( .A(x[290]), .B(y[290]), .Z(n25759) );
  XOR U36444 ( .A(x[289]), .B(y[289]), .Z(n25769) );
  XOR U36445 ( .A(x[288]), .B(y[288]), .Z(n25766) );
  XOR U36446 ( .A(x[287]), .B(y[287]), .Z(n25772) );
  XOR U36447 ( .A(x[286]), .B(y[286]), .Z(n26816) );
  XOR U36448 ( .A(x[285]), .B(y[285]), .Z(n25778) );
  XOR U36449 ( .A(x[284]), .B(y[284]), .Z(n25775) );
  XOR U36450 ( .A(x[283]), .B(y[283]), .Z(n25784) );
  XOR U36451 ( .A(x[282]), .B(y[282]), .Z(n25781) );
  XOR U36452 ( .A(x[281]), .B(y[281]), .Z(n26809) );
  XOR U36453 ( .A(x[280]), .B(y[280]), .Z(n26806) );
  XOR U36454 ( .A(x[279]), .B(y[279]), .Z(n26802) );
  XOR U36455 ( .A(x[278]), .B(y[278]), .Z(n26799) );
  XOR U36456 ( .A(x[277]), .B(y[277]), .Z(n26795) );
  XOR U36457 ( .A(x[276]), .B(y[276]), .Z(n26792) );
  XOR U36458 ( .A(x[275]), .B(y[275]), .Z(n25787) );
  XOR U36459 ( .A(x[274]), .B(y[274]), .Z(n26786) );
  XOR U36460 ( .A(x[273]), .B(y[273]), .Z(n25790) );
  XOR U36461 ( .A(x[272]), .B(y[272]), .Z(n25796) );
  XOR U36462 ( .A(x[271]), .B(y[271]), .Z(n25793) );
  XOR U36463 ( .A(x[270]), .B(y[270]), .Z(n25802) );
  XOR U36464 ( .A(x[269]), .B(y[269]), .Z(n25799) );
  XOR U36465 ( .A(x[268]), .B(y[268]), .Z(n25808) );
  XOR U36466 ( .A(x[267]), .B(y[267]), .Z(n25805) );
  XOR U36467 ( .A(x[266]), .B(y[266]), .Z(n25814) );
  XOR U36468 ( .A(x[265]), .B(y[265]), .Z(n25811) );
  XOR U36469 ( .A(x[264]), .B(y[264]), .Z(n25817) );
  XOR U36470 ( .A(x[263]), .B(y[263]), .Z(n26778) );
  XOR U36471 ( .A(x[262]), .B(y[262]), .Z(n26775) );
  XOR U36472 ( .A(x[261]), .B(y[261]), .Z(n25823) );
  XOR U36473 ( .A(x[260]), .B(y[260]), .Z(n25820) );
  XOR U36474 ( .A(x[259]), .B(y[259]), .Z(n26772) );
  XOR U36475 ( .A(x[258]), .B(y[258]), .Z(n26769) );
  XOR U36476 ( .A(x[257]), .B(y[257]), .Z(n25826) );
  XOR U36477 ( .A(x[256]), .B(y[256]), .Z(n26758) );
  XOR U36478 ( .A(x[255]), .B(y[255]), .Z(n25829) );
  XOR U36479 ( .A(x[254]), .B(y[254]), .Z(n25836) );
  XOR U36480 ( .A(x[253]), .B(y[253]), .Z(n25833) );
  XOR U36481 ( .A(x[252]), .B(y[252]), .Z(n26752) );
  XOR U36482 ( .A(x[251]), .B(y[251]), .Z(n26749) );
  XOR U36483 ( .A(x[250]), .B(y[250]), .Z(n25839) );
  XOR U36484 ( .A(x[249]), .B(y[249]), .Z(n26745) );
  XOR U36485 ( .A(x[248]), .B(y[248]), .Z(n26742) );
  XOR U36486 ( .A(x[247]), .B(y[247]), .Z(n26739) );
  XOR U36487 ( .A(x[246]), .B(y[246]), .Z(n26736) );
  XOR U36488 ( .A(x[245]), .B(y[245]), .Z(n26732) );
  XOR U36489 ( .A(x[244]), .B(y[244]), .Z(n26729) );
  XOR U36490 ( .A(x[243]), .B(y[243]), .Z(n25843) );
  XOR U36491 ( .A(x[242]), .B(y[242]), .Z(n26726) );
  XOR U36492 ( .A(x[241]), .B(y[241]), .Z(n26723) );
  XOR U36493 ( .A(x[240]), .B(y[240]), .Z(n26719) );
  XOR U36494 ( .A(x[239]), .B(y[239]), .Z(n26716) );
  XOR U36495 ( .A(x[238]), .B(y[238]), .Z(n25848) );
  XOR U36496 ( .A(x[237]), .B(y[237]), .Z(n25845) );
  XOR U36497 ( .A(x[236]), .B(y[236]), .Z(n25854) );
  XOR U36498 ( .A(x[235]), .B(y[235]), .Z(n25851) );
  XOR U36499 ( .A(x[234]), .B(y[234]), .Z(n25860) );
  XOR U36500 ( .A(x[233]), .B(y[233]), .Z(n25857) );
  XOR U36501 ( .A(x[232]), .B(y[232]), .Z(n25863) );
  XOR U36502 ( .A(x[231]), .B(y[231]), .Z(n26709) );
  XOR U36503 ( .A(x[230]), .B(y[230]), .Z(n26706) );
  XOR U36504 ( .A(x[229]), .B(y[229]), .Z(n26703) );
  XOR U36505 ( .A(x[228]), .B(y[228]), .Z(n26700) );
  XOR U36506 ( .A(x[227]), .B(y[227]), .Z(n26696) );
  XOR U36507 ( .A(x[226]), .B(y[226]), .Z(n26693) );
  XOR U36508 ( .A(x[225]), .B(y[225]), .Z(n26689) );
  XOR U36509 ( .A(x[224]), .B(y[224]), .Z(n26686) );
  XOR U36510 ( .A(x[223]), .B(y[223]), .Z(n26682) );
  XOR U36511 ( .A(x[222]), .B(y[222]), .Z(n26679) );
  XOR U36512 ( .A(x[221]), .B(y[221]), .Z(n26666) );
  XOR U36513 ( .A(x[220]), .B(y[220]), .Z(n26663) );
  XOR U36514 ( .A(x[219]), .B(y[219]), .Z(n25866) );
  XOR U36515 ( .A(x[218]), .B(y[218]), .Z(n25872) );
  XOR U36516 ( .A(x[217]), .B(y[217]), .Z(n25869) );
  XOR U36517 ( .A(x[216]), .B(y[216]), .Z(n25878) );
  XOR U36518 ( .A(x[215]), .B(y[215]), .Z(n25875) );
  XOR U36519 ( .A(x[214]), .B(y[214]), .Z(n26658) );
  XOR U36520 ( .A(x[213]), .B(y[213]), .Z(n26655) );
  XOR U36521 ( .A(x[212]), .B(y[212]), .Z(n26651) );
  XOR U36522 ( .A(x[211]), .B(y[211]), .Z(n26648) );
  XOR U36523 ( .A(x[210]), .B(y[210]), .Z(n25881) );
  XOR U36524 ( .A(x[209]), .B(y[209]), .Z(n26642) );
  XOR U36525 ( .A(x[208]), .B(y[208]), .Z(n25884) );
  XOR U36526 ( .A(x[207]), .B(y[207]), .Z(n25890) );
  XOR U36527 ( .A(x[206]), .B(y[206]), .Z(n25887) );
  XOR U36528 ( .A(x[205]), .B(y[205]), .Z(n25896) );
  XOR U36529 ( .A(x[204]), .B(y[204]), .Z(n25893) );
  XOR U36530 ( .A(x[203]), .B(y[203]), .Z(n25899) );
  XOR U36531 ( .A(x[202]), .B(y[202]), .Z(n25905) );
  XOR U36532 ( .A(x[201]), .B(y[201]), .Z(n25902) );
  XOR U36533 ( .A(x[200]), .B(y[200]), .Z(n25911) );
  XOR U36534 ( .A(x[199]), .B(y[199]), .Z(n25908) );
  XOR U36535 ( .A(x[198]), .B(y[198]), .Z(n25914) );
  XOR U36536 ( .A(x[197]), .B(y[197]), .Z(n26634) );
  XOR U36537 ( .A(x[196]), .B(y[196]), .Z(n26631) );
  XOR U36538 ( .A(x[195]), .B(y[195]), .Z(n25920) );
  XOR U36539 ( .A(x[194]), .B(y[194]), .Z(n25917) );
  XOR U36540 ( .A(x[193]), .B(y[193]), .Z(n25926) );
  XOR U36541 ( .A(x[192]), .B(y[192]), .Z(n25923) );
  XOR U36542 ( .A(x[191]), .B(y[191]), .Z(n25932) );
  XOR U36543 ( .A(x[190]), .B(y[190]), .Z(n25929) );
  XOR U36544 ( .A(x[189]), .B(y[189]), .Z(n26625) );
  XOR U36545 ( .A(x[188]), .B(y[188]), .Z(n26622) );
  XOR U36546 ( .A(x[187]), .B(y[187]), .Z(n26618) );
  XOR U36547 ( .A(x[186]), .B(y[186]), .Z(n26615) );
  XOR U36548 ( .A(x[185]), .B(y[185]), .Z(n26610) );
  XOR U36549 ( .A(x[184]), .B(y[184]), .Z(n26607) );
  XOR U36550 ( .A(x[183]), .B(y[183]), .Z(n25938) );
  XOR U36551 ( .A(x[182]), .B(y[182]), .Z(n25935) );
  XOR U36552 ( .A(x[181]), .B(y[181]), .Z(n25944) );
  XOR U36553 ( .A(x[180]), .B(y[180]), .Z(n25941) );
  XOR U36554 ( .A(x[179]), .B(y[179]), .Z(n25950) );
  XOR U36555 ( .A(x[178]), .B(y[178]), .Z(n25947) );
  XOR U36556 ( .A(x[177]), .B(y[177]), .Z(n26601) );
  XOR U36557 ( .A(x[176]), .B(y[176]), .Z(n26598) );
  XOR U36558 ( .A(x[175]), .B(y[175]), .Z(n26594) );
  XOR U36559 ( .A(x[174]), .B(y[174]), .Z(n26591) );
  XOR U36560 ( .A(x[173]), .B(y[173]), .Z(n26587) );
  XOR U36561 ( .A(x[172]), .B(y[172]), .Z(n26584) );
  XOR U36562 ( .A(x[171]), .B(y[171]), .Z(n25953) );
  XOR U36563 ( .A(x[170]), .B(y[170]), .Z(n26580) );
  XOR U36564 ( .A(x[169]), .B(y[169]), .Z(n26577) );
  XOR U36565 ( .A(x[168]), .B(y[168]), .Z(n26573) );
  XOR U36566 ( .A(x[167]), .B(y[167]), .Z(n26570) );
  XOR U36567 ( .A(x[166]), .B(y[166]), .Z(n25956) );
  XOR U36568 ( .A(x[165]), .B(y[165]), .Z(n25962) );
  XOR U36569 ( .A(x[164]), .B(y[164]), .Z(n25959) );
  XOR U36570 ( .A(x[163]), .B(y[163]), .Z(n25969) );
  XOR U36571 ( .A(x[162]), .B(y[162]), .Z(n25966) );
  XOR U36572 ( .A(x[161]), .B(y[161]), .Z(n25976) );
  XOR U36573 ( .A(x[160]), .B(y[160]), .Z(n25973) );
  XOR U36574 ( .A(x[159]), .B(y[159]), .Z(n25979) );
  XOR U36575 ( .A(x[158]), .B(y[158]), .Z(n26563) );
  XOR U36576 ( .A(x[157]), .B(y[157]), .Z(n26560) );
  XOR U36577 ( .A(x[156]), .B(y[156]), .Z(n25985) );
  XOR U36578 ( .A(x[155]), .B(y[155]), .Z(n25982) );
  XOR U36579 ( .A(x[154]), .B(y[154]), .Z(n25991) );
  XOR U36580 ( .A(x[153]), .B(y[153]), .Z(n25988) );
  XOR U36581 ( .A(x[152]), .B(y[152]), .Z(n25998) );
  XOR U36582 ( .A(x[151]), .B(y[151]), .Z(n25995) );
  XOR U36583 ( .A(x[150]), .B(y[150]), .Z(n26001) );
  XOR U36584 ( .A(x[149]), .B(y[149]), .Z(n26007) );
  XOR U36585 ( .A(x[148]), .B(y[148]), .Z(n26004) );
  XOR U36586 ( .A(x[147]), .B(y[147]), .Z(n26013) );
  XOR U36587 ( .A(x[146]), .B(y[146]), .Z(n26010) );
  XOR U36588 ( .A(x[145]), .B(y[145]), .Z(n26019) );
  XOR U36589 ( .A(x[144]), .B(y[144]), .Z(n26016) );
  XOR U36590 ( .A(x[143]), .B(y[143]), .Z(n26025) );
  XOR U36591 ( .A(x[142]), .B(y[142]), .Z(n26022) );
  XOR U36592 ( .A(x[141]), .B(y[141]), .Z(n26028) );
  XOR U36593 ( .A(x[140]), .B(y[140]), .Z(n26550) );
  XOR U36594 ( .A(x[139]), .B(y[139]), .Z(n26547) );
  XOR U36595 ( .A(x[138]), .B(y[138]), .Z(n26031) );
  XOR U36596 ( .A(x[137]), .B(y[137]), .Z(n26034) );
  XOR U36597 ( .A(x[136]), .B(y[136]), .Z(n26040) );
  XOR U36598 ( .A(x[135]), .B(y[135]), .Z(n26037) );
  XOR U36599 ( .A(x[134]), .B(y[134]), .Z(n26046) );
  XOR U36600 ( .A(x[133]), .B(y[133]), .Z(n26043) );
  XOR U36601 ( .A(x[132]), .B(y[132]), .Z(n26052) );
  XOR U36602 ( .A(x[131]), .B(y[131]), .Z(n26049) );
  XOR U36603 ( .A(x[130]), .B(y[130]), .Z(n26540) );
  XOR U36604 ( .A(x[129]), .B(y[129]), .Z(n26537) );
  XOR U36605 ( .A(x[128]), .B(y[128]), .Z(n26058) );
  XOR U36606 ( .A(x[127]), .B(y[127]), .Z(n26055) );
  XOR U36607 ( .A(x[126]), .B(y[126]), .Z(n26064) );
  XOR U36608 ( .A(x[125]), .B(y[125]), .Z(n26061) );
  XOR U36609 ( .A(x[124]), .B(y[124]), .Z(n26070) );
  XOR U36610 ( .A(x[123]), .B(y[123]), .Z(n26067) );
  XOR U36611 ( .A(x[122]), .B(y[122]), .Z(n26073) );
  XOR U36612 ( .A(x[121]), .B(y[121]), .Z(n26530) );
  XOR U36613 ( .A(x[120]), .B(y[120]), .Z(n26527) );
  XOR U36614 ( .A(x[119]), .B(y[119]), .Z(n26079) );
  XOR U36615 ( .A(x[118]), .B(y[118]), .Z(n26076) );
  XOR U36616 ( .A(x[117]), .B(y[117]), .Z(n26524) );
  XOR U36617 ( .A(x[116]), .B(y[116]), .Z(n26521) );
  XOR U36618 ( .A(x[115]), .B(y[115]), .Z(n26518) );
  XOR U36619 ( .A(x[114]), .B(y[114]), .Z(n26515) );
  XOR U36620 ( .A(x[113]), .B(y[113]), .Z(n26510) );
  XOR U36621 ( .A(x[112]), .B(y[112]), .Z(n26507) );
  XOR U36622 ( .A(x[111]), .B(y[111]), .Z(n26503) );
  XOR U36623 ( .A(x[110]), .B(y[110]), .Z(n26500) );
  XOR U36624 ( .A(x[109]), .B(y[109]), .Z(n26496) );
  XOR U36625 ( .A(x[108]), .B(y[108]), .Z(n26493) );
  XOR U36626 ( .A(x[107]), .B(y[107]), .Z(n26489) );
  XOR U36627 ( .A(x[106]), .B(y[106]), .Z(n26486) );
  XOR U36628 ( .A(x[105]), .B(y[105]), .Z(n26482) );
  XOR U36629 ( .A(x[104]), .B(y[104]), .Z(n26479) );
  XOR U36630 ( .A(x[103]), .B(y[103]), .Z(n26085) );
  XOR U36631 ( .A(x[102]), .B(y[102]), .Z(n26082) );
  XOR U36632 ( .A(x[101]), .B(y[101]), .Z(n26091) );
  XOR U36633 ( .A(x[100]), .B(y[100]), .Z(n26088) );
  XOR U36634 ( .A(x[99]), .B(y[99]), .Z(n26097) );
  XOR U36635 ( .A(x[98]), .B(y[98]), .Z(n26094) );
  XOR U36636 ( .A(x[97]), .B(y[97]), .Z(n26475) );
  XOR U36637 ( .A(x[96]), .B(y[96]), .Z(n26472) );
  XOR U36638 ( .A(x[95]), .B(y[95]), .Z(n26469) );
  XOR U36639 ( .A(x[94]), .B(y[94]), .Z(n26466) );
  XOR U36640 ( .A(x[93]), .B(y[93]), .Z(n26462) );
  XOR U36641 ( .A(x[92]), .B(y[92]), .Z(n26459) );
  XOR U36642 ( .A(x[91]), .B(y[91]), .Z(n26103) );
  XOR U36643 ( .A(x[90]), .B(y[90]), .Z(n26100) );
  XOR U36644 ( .A(x[89]), .B(y[89]), .Z(n26454) );
  XOR U36645 ( .A(x[88]), .B(y[88]), .Z(n26451) );
  XOR U36646 ( .A(x[87]), .B(y[87]), .Z(n26447) );
  XOR U36647 ( .A(x[86]), .B(y[86]), .Z(n26444) );
  XOR U36648 ( .A(x[85]), .B(y[85]), .Z(n26440) );
  XOR U36649 ( .A(x[84]), .B(y[84]), .Z(n26437) );
  XOR U36650 ( .A(x[83]), .B(y[83]), .Z(n26109) );
  XOR U36651 ( .A(x[82]), .B(y[82]), .Z(n26106) );
  XOR U36652 ( .A(x[81]), .B(y[81]), .Z(n26433) );
  XOR U36653 ( .A(x[80]), .B(y[80]), .Z(n26430) );
  XOR U36654 ( .A(x[79]), .B(y[79]), .Z(n26426) );
  XOR U36655 ( .A(x[78]), .B(y[78]), .Z(n26423) );
  XOR U36656 ( .A(x[77]), .B(y[77]), .Z(n26419) );
  XOR U36657 ( .A(x[76]), .B(y[76]), .Z(n26416) );
  XOR U36658 ( .A(x[75]), .B(y[75]), .Z(n26112) );
  XOR U36659 ( .A(x[74]), .B(y[74]), .Z(n26413) );
  XOR U36660 ( .A(x[73]), .B(y[73]), .Z(n26410) );
  XOR U36661 ( .A(x[72]), .B(y[72]), .Z(n26405) );
  XOR U36662 ( .A(x[71]), .B(y[71]), .Z(n26402) );
  XOR U36663 ( .A(x[70]), .B(y[70]), .Z(n26115) );
  XOR U36664 ( .A(x[69]), .B(y[69]), .Z(n26121) );
  XOR U36665 ( .A(x[68]), .B(y[68]), .Z(n26118) );
  XOR U36666 ( .A(x[67]), .B(y[67]), .Z(n26127) );
  XOR U36667 ( .A(x[66]), .B(y[66]), .Z(n26124) );
  XOR U36668 ( .A(x[65]), .B(y[65]), .Z(n26133) );
  XOR U36669 ( .A(x[64]), .B(y[64]), .Z(n26130) );
  XOR U36670 ( .A(x[63]), .B(y[63]), .Z(n26395) );
  XOR U36671 ( .A(x[62]), .B(y[62]), .Z(n26392) );
  XOR U36672 ( .A(x[61]), .B(y[61]), .Z(n26380) );
  XOR U36673 ( .A(x[60]), .B(y[60]), .Z(n26136) );
  XOR U36674 ( .A(x[59]), .B(y[59]), .Z(n26384) );
  XOR U36675 ( .A(x[58]), .B(y[58]), .Z(n26143) );
  XOR U36676 ( .A(x[57]), .B(y[57]), .Z(n26140) );
  XOR U36677 ( .A(x[56]), .B(y[56]), .Z(n26149) );
  XOR U36678 ( .A(x[55]), .B(y[55]), .Z(n26146) );
  XOR U36679 ( .A(x[54]), .B(y[54]), .Z(n26375) );
  XOR U36680 ( .A(x[53]), .B(y[53]), .Z(n26372) );
  XOR U36681 ( .A(x[52]), .B(y[52]), .Z(n26359) );
  XOR U36682 ( .A(x[51]), .B(y[51]), .Z(n26356) );
  XOR U36683 ( .A(x[50]), .B(y[50]), .Z(n26152) );
  XOR U36684 ( .A(x[49]), .B(y[49]), .Z(n26158) );
  XOR U36685 ( .A(x[48]), .B(y[48]), .Z(n26155) );
  XOR U36686 ( .A(x[47]), .B(y[47]), .Z(n26164) );
  XOR U36687 ( .A(x[46]), .B(y[46]), .Z(n26161) );
  XOR U36688 ( .A(x[45]), .B(y[45]), .Z(n26349) );
  XOR U36689 ( .A(x[44]), .B(y[44]), .Z(n26346) );
  XOR U36690 ( .A(x[43]), .B(y[43]), .Z(n26167) );
  XOR U36691 ( .A(x[42]), .B(y[42]), .Z(n26174) );
  XOR U36692 ( .A(x[41]), .B(y[41]), .Z(n26171) );
  XOR U36693 ( .A(x[40]), .B(y[40]), .Z(n26180) );
  XOR U36694 ( .A(x[39]), .B(y[39]), .Z(n26177) );
  XOR U36695 ( .A(x[38]), .B(y[38]), .Z(n26341) );
  XOR U36696 ( .A(x[37]), .B(y[37]), .Z(n26338) );
  XOR U36697 ( .A(x[36]), .B(y[36]), .Z(n26334) );
  XOR U36698 ( .A(x[35]), .B(y[35]), .Z(n26331) );
  XOR U36699 ( .A(x[34]), .B(y[34]), .Z(n26327) );
  XOR U36700 ( .A(x[33]), .B(y[33]), .Z(n26324) );
  XOR U36701 ( .A(x[32]), .B(y[32]), .Z(n26183) );
  XOR U36702 ( .A(x[31]), .B(y[31]), .Z(n26186) );
  XOR U36703 ( .A(x[30]), .B(y[30]), .Z(n26312) );
  XOR U36704 ( .A(x[29]), .B(y[29]), .Z(n26189) );
  XOR U36705 ( .A(x[28]), .B(y[28]), .Z(n26301) );
  XOR U36706 ( .A(x[27]), .B(y[27]), .Z(n26192) );
  XOR U36707 ( .A(x[26]), .B(y[26]), .Z(n26295) );
  XOR U36708 ( .A(x[25]), .B(y[25]), .Z(n26292) );
  XOR U36709 ( .A(x[24]), .B(y[24]), .Z(n26195) );
  XOR U36710 ( .A(x[23]), .B(y[23]), .Z(n26201) );
  XOR U36711 ( .A(x[22]), .B(y[22]), .Z(n26198) );
  XOR U36712 ( .A(x[21]), .B(y[21]), .Z(n26288) );
  XOR U36713 ( .A(x[20]), .B(y[20]), .Z(n26285) );
  XOR U36714 ( .A(x[19]), .B(y[19]), .Z(n26207) );
  XOR U36715 ( .A(x[18]), .B(y[18]), .Z(n26204) );
  XOR U36716 ( .A(x[17]), .B(y[17]), .Z(n26280) );
  XOR U36717 ( .A(x[16]), .B(y[16]), .Z(n26277) );
  XOR U36718 ( .A(x[15]), .B(y[15]), .Z(n26210) );
  XOR U36719 ( .A(x[14]), .B(y[14]), .Z(n26272) );
  XOR U36720 ( .A(x[13]), .B(y[13]), .Z(n26269) );
  XOR U36721 ( .A(x[12]), .B(y[12]), .Z(n26213) );
  XOR U36722 ( .A(x[11]), .B(y[11]), .Z(n26264) );
  XOR U36723 ( .A(x[10]), .B(y[10]), .Z(n26261) );
  XOR U36724 ( .A(x[9]), .B(y[9]), .Z(n26216) );
  XOR U36725 ( .A(x[8]), .B(y[8]), .Z(n26219) );
  XOR U36726 ( .A(x[7]), .B(y[7]), .Z(n26222) );
  XOR U36727 ( .A(x[6]), .B(y[6]), .Z(n26247) );
  XOR U36728 ( .A(x[5]), .B(y[5]), .Z(n26225) );
  XOR U36729 ( .A(x[4]), .B(y[4]), .Z(n26228) );
  XOR U36730 ( .A(x[3]), .B(y[3]), .Z(n26231) );
  XOR U36731 ( .A(x[2]), .B(y[2]), .Z(n26239) );
  IV U36732 ( .A(x[1]), .Z(n24501) );
  XOR U36733 ( .A(n24501), .B(y[1]), .Z(n26236) );
  XOR U36734 ( .A(x[0]), .B(y[0]), .Z(n26234) );
  XOR U36735 ( .A(n26236), .B(n26234), .Z(n26240) );
  XOR U36736 ( .A(n26239), .B(n26240), .Z(n26232) );
  XOR U36737 ( .A(n26231), .B(n26232), .Z(n26230) );
  XOR U36738 ( .A(n26228), .B(n26230), .Z(n26227) );
  XOR U36739 ( .A(n26225), .B(n26227), .Z(n26248) );
  XOR U36740 ( .A(n26247), .B(n26248), .Z(n26223) );
  XOR U36741 ( .A(n26222), .B(n26223), .Z(n26221) );
  XOR U36742 ( .A(n26219), .B(n26221), .Z(n26217) );
  XOR U36743 ( .A(n26216), .B(n26217), .Z(n26262) );
  XOR U36744 ( .A(n26261), .B(n26262), .Z(n26265) );
  XOR U36745 ( .A(n26264), .B(n26265), .Z(n26214) );
  XOR U36746 ( .A(n26213), .B(n26214), .Z(n26270) );
  XOR U36747 ( .A(n26269), .B(n26270), .Z(n26274) );
  XOR U36748 ( .A(n26272), .B(n26274), .Z(n26212) );
  XOR U36749 ( .A(n26210), .B(n26212), .Z(n26279) );
  XOR U36750 ( .A(n26277), .B(n26279), .Z(n26282) );
  XOR U36751 ( .A(n26280), .B(n26282), .Z(n26206) );
  XOR U36752 ( .A(n26204), .B(n26206), .Z(n26209) );
  XOR U36753 ( .A(n26207), .B(n26209), .Z(n26286) );
  XOR U36754 ( .A(n26285), .B(n26286), .Z(n26290) );
  XOR U36755 ( .A(n26288), .B(n26290), .Z(n26200) );
  XOR U36756 ( .A(n26198), .B(n26200), .Z(n26203) );
  XOR U36757 ( .A(n26201), .B(n26203), .Z(n26196) );
  XOR U36758 ( .A(n26195), .B(n26196), .Z(n26293) );
  XOR U36759 ( .A(n26292), .B(n26293), .Z(n26297) );
  XOR U36760 ( .A(n26295), .B(n26297), .Z(n26194) );
  XOR U36761 ( .A(n26192), .B(n26194), .Z(n26302) );
  XOR U36762 ( .A(n26301), .B(n26302), .Z(n26190) );
  XOR U36763 ( .A(n26189), .B(n26190), .Z(n26314) );
  XOR U36764 ( .A(n26312), .B(n26314), .Z(n26188) );
  XOR U36765 ( .A(n26186), .B(n26188), .Z(n26184) );
  XOR U36766 ( .A(n26183), .B(n26184), .Z(n26325) );
  XOR U36767 ( .A(n26324), .B(n26325), .Z(n26329) );
  XOR U36768 ( .A(n26327), .B(n26329), .Z(n26333) );
  XOR U36769 ( .A(n26331), .B(n26333), .Z(n26336) );
  XOR U36770 ( .A(n26334), .B(n26336), .Z(n26340) );
  XOR U36771 ( .A(n26338), .B(n26340), .Z(n26343) );
  XOR U36772 ( .A(n26341), .B(n26343), .Z(n26179) );
  XOR U36773 ( .A(n26177), .B(n26179), .Z(n26181) );
  XOR U36774 ( .A(n26180), .B(n26181), .Z(n26172) );
  XOR U36775 ( .A(n26171), .B(n26172), .Z(n26176) );
  XOR U36776 ( .A(n26174), .B(n26176), .Z(n26168) );
  XOR U36777 ( .A(n26167), .B(n26168), .Z(n26347) );
  XOR U36778 ( .A(n26346), .B(n26347), .Z(n26351) );
  XOR U36779 ( .A(n26349), .B(n26351), .Z(n26163) );
  XOR U36780 ( .A(n26161), .B(n26163), .Z(n26166) );
  XOR U36781 ( .A(n26164), .B(n26166), .Z(n26156) );
  XOR U36782 ( .A(n26155), .B(n26156), .Z(n26160) );
  XOR U36783 ( .A(n26158), .B(n26160), .Z(n26153) );
  XOR U36784 ( .A(n26152), .B(n26153), .Z(n26358) );
  XOR U36785 ( .A(n26356), .B(n26358), .Z(n26360) );
  XOR U36786 ( .A(n26359), .B(n26360), .Z(n26374) );
  XOR U36787 ( .A(n26372), .B(n26374), .Z(n26377) );
  XOR U36788 ( .A(n26375), .B(n26377), .Z(n26148) );
  XOR U36789 ( .A(n26146), .B(n26148), .Z(n26151) );
  XOR U36790 ( .A(n26149), .B(n26151), .Z(n26142) );
  XOR U36791 ( .A(n26140), .B(n26142), .Z(n26145) );
  XOR U36792 ( .A(n26143), .B(n26145), .Z(n26386) );
  XOR U36793 ( .A(n26384), .B(n26386), .Z(n26138) );
  XOR U36794 ( .A(n26136), .B(n26138), .Z(n26382) );
  XOR U36795 ( .A(n26380), .B(n26382), .Z(n26394) );
  XOR U36796 ( .A(n26392), .B(n26394), .Z(n26397) );
  XOR U36797 ( .A(n26395), .B(n26397), .Z(n26131) );
  XOR U36798 ( .A(n26130), .B(n26131), .Z(n26135) );
  XOR U36799 ( .A(n26133), .B(n26135), .Z(n26126) );
  XOR U36800 ( .A(n26124), .B(n26126), .Z(n26129) );
  XOR U36801 ( .A(n26127), .B(n26129), .Z(n26119) );
  XOR U36802 ( .A(n26118), .B(n26119), .Z(n26122) );
  XOR U36803 ( .A(n26121), .B(n26122), .Z(n26117) );
  XOR U36804 ( .A(n26115), .B(n26117), .Z(n26403) );
  XOR U36805 ( .A(n26402), .B(n26403), .Z(n26406) );
  XOR U36806 ( .A(n26405), .B(n26406), .Z(n26411) );
  XOR U36807 ( .A(n26410), .B(n26411), .Z(n26415) );
  XOR U36808 ( .A(n26413), .B(n26415), .Z(n26114) );
  XOR U36809 ( .A(n26112), .B(n26114), .Z(n26417) );
  XOR U36810 ( .A(n26416), .B(n26417), .Z(n26420) );
  XOR U36811 ( .A(n26419), .B(n26420), .Z(n26425) );
  XOR U36812 ( .A(n26423), .B(n26425), .Z(n26427) );
  XOR U36813 ( .A(n26426), .B(n26427), .Z(n26431) );
  XOR U36814 ( .A(n26430), .B(n26431), .Z(n26434) );
  XOR U36815 ( .A(n26433), .B(n26434), .Z(n26108) );
  XOR U36816 ( .A(n26106), .B(n26108), .Z(n26111) );
  XOR U36817 ( .A(n26109), .B(n26111), .Z(n26438) );
  XOR U36818 ( .A(n26437), .B(n26438), .Z(n26442) );
  XOR U36819 ( .A(n26440), .B(n26442), .Z(n26446) );
  XOR U36820 ( .A(n26444), .B(n26446), .Z(n26449) );
  XOR U36821 ( .A(n26447), .B(n26449), .Z(n26453) );
  XOR U36822 ( .A(n26451), .B(n26453), .Z(n26456) );
  XOR U36823 ( .A(n26454), .B(n26456), .Z(n26101) );
  XOR U36824 ( .A(n26100), .B(n26101), .Z(n26104) );
  XOR U36825 ( .A(n26103), .B(n26104), .Z(n26461) );
  XOR U36826 ( .A(n26459), .B(n26461), .Z(n26464) );
  XOR U36827 ( .A(n26462), .B(n26464), .Z(n26468) );
  XOR U36828 ( .A(n26466), .B(n26468), .Z(n26471) );
  XOR U36829 ( .A(n26469), .B(n26471), .Z(n26473) );
  XOR U36830 ( .A(n26472), .B(n26473), .Z(n26477) );
  XOR U36831 ( .A(n26475), .B(n26477), .Z(n26096) );
  XOR U36832 ( .A(n26094), .B(n26096), .Z(n26098) );
  XOR U36833 ( .A(n26097), .B(n26098), .Z(n26089) );
  XOR U36834 ( .A(n26088), .B(n26089), .Z(n26093) );
  XOR U36835 ( .A(n26091), .B(n26093), .Z(n26084) );
  XOR U36836 ( .A(n26082), .B(n26084), .Z(n26087) );
  XOR U36837 ( .A(n26085), .B(n26087), .Z(n26480) );
  XOR U36838 ( .A(n26479), .B(n26480), .Z(n26484) );
  XOR U36839 ( .A(n26482), .B(n26484), .Z(n26488) );
  XOR U36840 ( .A(n26486), .B(n26488), .Z(n26491) );
  XOR U36841 ( .A(n26489), .B(n26491), .Z(n26494) );
  XOR U36842 ( .A(n26493), .B(n26494), .Z(n26498) );
  XOR U36843 ( .A(n26496), .B(n26498), .Z(n26502) );
  XOR U36844 ( .A(n26500), .B(n26502), .Z(n26505) );
  XOR U36845 ( .A(n26503), .B(n26505), .Z(n26508) );
  XOR U36846 ( .A(n26507), .B(n26508), .Z(n26511) );
  XOR U36847 ( .A(n26510), .B(n26511), .Z(n26517) );
  XOR U36848 ( .A(n26515), .B(n26517), .Z(n26520) );
  XOR U36849 ( .A(n26518), .B(n26520), .Z(n26523) );
  XOR U36850 ( .A(n26521), .B(n26523), .Z(n26526) );
  XOR U36851 ( .A(n26524), .B(n26526), .Z(n26078) );
  XOR U36852 ( .A(n26076), .B(n26078), .Z(n26081) );
  XOR U36853 ( .A(n26079), .B(n26081), .Z(n26528) );
  XOR U36854 ( .A(n26527), .B(n26528), .Z(n26531) );
  XOR U36855 ( .A(n26530), .B(n26531), .Z(n26074) );
  XOR U36856 ( .A(n26073), .B(n26074), .Z(n26068) );
  XOR U36857 ( .A(n26067), .B(n26068), .Z(n26071) );
  XOR U36858 ( .A(n26070), .B(n26071), .Z(n26063) );
  XOR U36859 ( .A(n26061), .B(n26063), .Z(n26066) );
  XOR U36860 ( .A(n26064), .B(n26066), .Z(n26057) );
  XOR U36861 ( .A(n26055), .B(n26057), .Z(n26059) );
  XOR U36862 ( .A(n26058), .B(n26059), .Z(n26539) );
  XOR U36863 ( .A(n26537), .B(n26539), .Z(n26542) );
  XOR U36864 ( .A(n26540), .B(n26542), .Z(n26050) );
  XOR U36865 ( .A(n26049), .B(n26050), .Z(n26053) );
  XOR U36866 ( .A(n26052), .B(n26053), .Z(n26044) );
  XOR U36867 ( .A(n26043), .B(n26044), .Z(n26048) );
  XOR U36868 ( .A(n26046), .B(n26048), .Z(n26039) );
  XOR U36869 ( .A(n26037), .B(n26039), .Z(n26041) );
  XOR U36870 ( .A(n26040), .B(n26041), .Z(n26035) );
  XOR U36871 ( .A(n26034), .B(n26035), .Z(n26033) );
  XOR U36872 ( .A(n26031), .B(n26033), .Z(n26549) );
  XOR U36873 ( .A(n26547), .B(n26549), .Z(n26551) );
  XOR U36874 ( .A(n26550), .B(n26551), .Z(n26030) );
  XOR U36875 ( .A(n26028), .B(n26030), .Z(n26024) );
  XOR U36876 ( .A(n26022), .B(n26024), .Z(n26026) );
  XOR U36877 ( .A(n26025), .B(n26026), .Z(n26017) );
  XOR U36878 ( .A(n26016), .B(n26017), .Z(n26020) );
  XOR U36879 ( .A(n26019), .B(n26020), .Z(n26012) );
  XOR U36880 ( .A(n26010), .B(n26012), .Z(n26015) );
  XOR U36881 ( .A(n26013), .B(n26015), .Z(n26006) );
  XOR U36882 ( .A(n26004), .B(n26006), .Z(n26009) );
  XOR U36883 ( .A(n26007), .B(n26009), .Z(n26003) );
  XOR U36884 ( .A(n26001), .B(n26003), .Z(n25997) );
  XOR U36885 ( .A(n25995), .B(n25997), .Z(n25999) );
  XOR U36886 ( .A(n25998), .B(n25999), .Z(n25990) );
  XOR U36887 ( .A(n25988), .B(n25990), .Z(n25993) );
  XOR U36888 ( .A(n25991), .B(n25993), .Z(n25983) );
  XOR U36889 ( .A(n25982), .B(n25983), .Z(n25986) );
  XOR U36890 ( .A(n25985), .B(n25986), .Z(n26562) );
  XOR U36891 ( .A(n26560), .B(n26562), .Z(n26564) );
  XOR U36892 ( .A(n26563), .B(n26564), .Z(n25981) );
  XOR U36893 ( .A(n25979), .B(n25981), .Z(n25975) );
  XOR U36894 ( .A(n25973), .B(n25975), .Z(n25978) );
  XOR U36895 ( .A(n25976), .B(n25978), .Z(n25967) );
  XOR U36896 ( .A(n25966), .B(n25967), .Z(n25971) );
  XOR U36897 ( .A(n25969), .B(n25971), .Z(n25960) );
  XOR U36898 ( .A(n25959), .B(n25960), .Z(n25964) );
  XOR U36899 ( .A(n25962), .B(n25964), .Z(n25958) );
  XOR U36900 ( .A(n25956), .B(n25958), .Z(n26571) );
  XOR U36901 ( .A(n26570), .B(n26571), .Z(n26574) );
  XOR U36902 ( .A(n26573), .B(n26574), .Z(n26579) );
  XOR U36903 ( .A(n26577), .B(n26579), .Z(n26581) );
  XOR U36904 ( .A(n26580), .B(n26581), .Z(n25955) );
  XOR U36905 ( .A(n25953), .B(n25955), .Z(n26585) );
  XOR U36906 ( .A(n26584), .B(n26585), .Z(n26589) );
  XOR U36907 ( .A(n26587), .B(n26589), .Z(n26593) );
  XOR U36908 ( .A(n26591), .B(n26593), .Z(n26595) );
  XOR U36909 ( .A(n26594), .B(n26595), .Z(n26599) );
  XOR U36910 ( .A(n26598), .B(n26599), .Z(n26602) );
  XOR U36911 ( .A(n26601), .B(n26602), .Z(n25949) );
  XOR U36912 ( .A(n25947), .B(n25949), .Z(n25952) );
  XOR U36913 ( .A(n25950), .B(n25952), .Z(n25942) );
  XOR U36914 ( .A(n25941), .B(n25942), .Z(n25946) );
  XOR U36915 ( .A(n25944), .B(n25946), .Z(n25937) );
  XOR U36916 ( .A(n25935), .B(n25937), .Z(n25940) );
  XOR U36917 ( .A(n25938), .B(n25940), .Z(n26608) );
  XOR U36918 ( .A(n26607), .B(n26608), .Z(n26612) );
  XOR U36919 ( .A(n26610), .B(n26612), .Z(n26616) );
  XOR U36920 ( .A(n26615), .B(n26616), .Z(n26619) );
  XOR U36921 ( .A(n26618), .B(n26619), .Z(n26624) );
  XOR U36922 ( .A(n26622), .B(n26624), .Z(n26627) );
  XOR U36923 ( .A(n26625), .B(n26627), .Z(n25931) );
  XOR U36924 ( .A(n25929), .B(n25931), .Z(n25934) );
  XOR U36925 ( .A(n25932), .B(n25934), .Z(n25924) );
  XOR U36926 ( .A(n25923), .B(n25924), .Z(n25928) );
  XOR U36927 ( .A(n25926), .B(n25928), .Z(n25919) );
  XOR U36928 ( .A(n25917), .B(n25919), .Z(n25922) );
  XOR U36929 ( .A(n25920), .B(n25922), .Z(n26633) );
  XOR U36930 ( .A(n26631), .B(n26633), .Z(n26636) );
  XOR U36931 ( .A(n26634), .B(n26636), .Z(n25915) );
  XOR U36932 ( .A(n25914), .B(n25915), .Z(n25910) );
  XOR U36933 ( .A(n25908), .B(n25910), .Z(n25912) );
  XOR U36934 ( .A(n25911), .B(n25912), .Z(n25903) );
  XOR U36935 ( .A(n25902), .B(n25903), .Z(n25907) );
  XOR U36936 ( .A(n25905), .B(n25907), .Z(n25901) );
  XOR U36937 ( .A(n25899), .B(n25901), .Z(n25894) );
  XOR U36938 ( .A(n25893), .B(n25894), .Z(n25897) );
  XOR U36939 ( .A(n25896), .B(n25897), .Z(n25889) );
  XOR U36940 ( .A(n25887), .B(n25889), .Z(n25892) );
  XOR U36941 ( .A(n25890), .B(n25892), .Z(n25886) );
  XOR U36942 ( .A(n25884), .B(n25886), .Z(n26644) );
  XOR U36943 ( .A(n26642), .B(n26644), .Z(n25883) );
  XOR U36944 ( .A(n25881), .B(n25883), .Z(n26650) );
  XOR U36945 ( .A(n26648), .B(n26650), .Z(n26652) );
  XOR U36946 ( .A(n26651), .B(n26652), .Z(n26657) );
  XOR U36947 ( .A(n26655), .B(n26657), .Z(n26660) );
  XOR U36948 ( .A(n26658), .B(n26660), .Z(n25877) );
  XOR U36949 ( .A(n25875), .B(n25877), .Z(n25879) );
  XOR U36950 ( .A(n25878), .B(n25879), .Z(n25870) );
  XOR U36951 ( .A(n25869), .B(n25870), .Z(n25874) );
  XOR U36952 ( .A(n25872), .B(n25874), .Z(n25868) );
  XOR U36953 ( .A(n25866), .B(n25868), .Z(n26664) );
  XOR U36954 ( .A(n26663), .B(n26664), .Z(n26668) );
  XOR U36955 ( .A(n26666), .B(n26668), .Z(n26681) );
  XOR U36956 ( .A(n26679), .B(n26681), .Z(n26684) );
  XOR U36957 ( .A(n26682), .B(n26684), .Z(n26687) );
  XOR U36958 ( .A(n26686), .B(n26687), .Z(n26691) );
  XOR U36959 ( .A(n26689), .B(n26691), .Z(n26695) );
  XOR U36960 ( .A(n26693), .B(n26695), .Z(n26697) );
  XOR U36961 ( .A(n26696), .B(n26697), .Z(n26701) );
  XOR U36962 ( .A(n26700), .B(n26701), .Z(n26704) );
  XOR U36963 ( .A(n26703), .B(n26704), .Z(n26708) );
  XOR U36964 ( .A(n26706), .B(n26708), .Z(n26710) );
  XOR U36965 ( .A(n26709), .B(n26710), .Z(n25864) );
  XOR U36966 ( .A(n25863), .B(n25864), .Z(n25858) );
  XOR U36967 ( .A(n25857), .B(n25858), .Z(n25862) );
  XOR U36968 ( .A(n25860), .B(n25862), .Z(n25853) );
  XOR U36969 ( .A(n25851), .B(n25853), .Z(n25855) );
  XOR U36970 ( .A(n25854), .B(n25855), .Z(n25847) );
  XOR U36971 ( .A(n25845), .B(n25847), .Z(n25850) );
  XOR U36972 ( .A(n25848), .B(n25850), .Z(n26717) );
  XOR U36973 ( .A(n26716), .B(n26717), .Z(n26720) );
  XOR U36974 ( .A(n26719), .B(n26720), .Z(n26724) );
  XOR U36975 ( .A(n26723), .B(n26724), .Z(n26728) );
  XOR U36976 ( .A(n26726), .B(n26728), .Z(n46500) );
  XOR U36977 ( .A(n25843), .B(n46500), .Z(n26730) );
  XOR U36978 ( .A(n26729), .B(n26730), .Z(n26734) );
  XOR U36979 ( .A(n26732), .B(n26734), .Z(n26738) );
  XOR U36980 ( .A(n26736), .B(n26738), .Z(n26741) );
  XOR U36981 ( .A(n26739), .B(n26741), .Z(n26743) );
  XOR U36982 ( .A(n26742), .B(n26743), .Z(n26747) );
  XOR U36983 ( .A(n26745), .B(n26747), .Z(n25841) );
  XOR U36984 ( .A(n25839), .B(n25841), .Z(n26751) );
  XOR U36985 ( .A(n26749), .B(n26751), .Z(n26753) );
  XOR U36986 ( .A(n26752), .B(n26753), .Z(n25835) );
  XOR U36987 ( .A(n25833), .B(n25835), .Z(n25838) );
  XOR U36988 ( .A(n25836), .B(n25838), .Z(n25831) );
  XOR U36989 ( .A(n25829), .B(n25831), .Z(n26759) );
  XOR U36990 ( .A(n26758), .B(n26759), .Z(n25828) );
  XOR U36991 ( .A(n25826), .B(n25828), .Z(n26771) );
  XOR U36992 ( .A(n26769), .B(n26771), .Z(n26773) );
  XOR U36993 ( .A(n26772), .B(n26773), .Z(n25821) );
  XOR U36994 ( .A(n25820), .B(n25821), .Z(n25825) );
  XOR U36995 ( .A(n25823), .B(n25825), .Z(n26776) );
  XOR U36996 ( .A(n26775), .B(n26776), .Z(n26780) );
  XOR U36997 ( .A(n26778), .B(n26780), .Z(n25818) );
  XOR U36998 ( .A(n25817), .B(n25818), .Z(n25813) );
  XOR U36999 ( .A(n25811), .B(n25813), .Z(n25816) );
  XOR U37000 ( .A(n25814), .B(n25816), .Z(n25807) );
  XOR U37001 ( .A(n25805), .B(n25807), .Z(n25810) );
  XOR U37002 ( .A(n25808), .B(n25810), .Z(n25801) );
  XOR U37003 ( .A(n25799), .B(n25801), .Z(n25803) );
  XOR U37004 ( .A(n25802), .B(n25803), .Z(n25795) );
  XOR U37005 ( .A(n25793), .B(n25795), .Z(n25797) );
  XOR U37006 ( .A(n25796), .B(n25797), .Z(n25791) );
  XOR U37007 ( .A(n25790), .B(n25791), .Z(n26788) );
  XOR U37008 ( .A(n26786), .B(n26788), .Z(n25788) );
  XOR U37009 ( .A(n25787), .B(n25788), .Z(n26793) );
  XOR U37010 ( .A(n26792), .B(n26793), .Z(n26797) );
  XOR U37011 ( .A(n26795), .B(n26797), .Z(n26801) );
  XOR U37012 ( .A(n26799), .B(n26801), .Z(n26804) );
  XOR U37013 ( .A(n26802), .B(n26804), .Z(n26807) );
  XOR U37014 ( .A(n26806), .B(n26807), .Z(n26810) );
  XOR U37015 ( .A(n26809), .B(n26810), .Z(n25783) );
  XOR U37016 ( .A(n25781), .B(n25783), .Z(n25786) );
  XOR U37017 ( .A(n25784), .B(n25786), .Z(n25776) );
  XOR U37018 ( .A(n25775), .B(n25776), .Z(n25780) );
  XOR U37019 ( .A(n25778), .B(n25780), .Z(n26817) );
  XOR U37020 ( .A(n26816), .B(n26817), .Z(n25774) );
  XOR U37021 ( .A(n25772), .B(n25774), .Z(n25768) );
  XOR U37022 ( .A(n25766), .B(n25768), .Z(n25771) );
  XOR U37023 ( .A(n25769), .B(n25771), .Z(n25760) );
  XOR U37024 ( .A(n25759), .B(n25760), .Z(n25764) );
  XOR U37025 ( .A(n25762), .B(n25764), .Z(n25755) );
  XOR U37026 ( .A(n25753), .B(n25755), .Z(n25758) );
  XOR U37027 ( .A(n25756), .B(n25758), .Z(n26823) );
  XOR U37028 ( .A(n26821), .B(n26823), .Z(n26825) );
  XOR U37029 ( .A(n26824), .B(n26825), .Z(n25751) );
  XOR U37030 ( .A(n25750), .B(n25751), .Z(n26831) );
  XOR U37031 ( .A(n26830), .B(n26831), .Z(n25749) );
  XOR U37032 ( .A(n25747), .B(n25749), .Z(n26838) );
  XOR U37033 ( .A(n26836), .B(n26838), .Z(n26840) );
  XOR U37034 ( .A(n26839), .B(n26840), .Z(n26845) );
  XOR U37035 ( .A(n26843), .B(n26845), .Z(n26848) );
  XOR U37036 ( .A(n26846), .B(n26848), .Z(n26852) );
  XOR U37037 ( .A(n26850), .B(n26852), .Z(n26854) );
  XOR U37038 ( .A(n26853), .B(n26854), .Z(n26858) );
  XOR U37039 ( .A(n26857), .B(n26858), .Z(n26862) );
  XOR U37040 ( .A(n26860), .B(n26862), .Z(n26865) );
  XOR U37041 ( .A(n26863), .B(n26865), .Z(n26867) );
  XOR U37042 ( .A(n26866), .B(n26867), .Z(n25743) );
  XOR U37043 ( .A(n25741), .B(n25743), .Z(n25746) );
  XOR U37044 ( .A(n25744), .B(n25746), .Z(n25739) );
  XOR U37045 ( .A(n25738), .B(n25739), .Z(n26873) );
  XOR U37046 ( .A(n26872), .B(n26873), .Z(n26877) );
  XOR U37047 ( .A(n26875), .B(n26877), .Z(n26881) );
  XOR U37048 ( .A(n26879), .B(n26881), .Z(n26883) );
  XOR U37049 ( .A(n26882), .B(n26883), .Z(n26887) );
  XOR U37050 ( .A(n26886), .B(n26887), .Z(n26891) );
  XOR U37051 ( .A(n26889), .B(n26891), .Z(n25735) );
  XOR U37052 ( .A(n25734), .B(n25735), .Z(n25730) );
  XOR U37053 ( .A(n25728), .B(n25730), .Z(n25732) );
  XOR U37054 ( .A(n25731), .B(n25732), .Z(n25724) );
  XOR U37055 ( .A(n25722), .B(n25724), .Z(n25727) );
  XOR U37056 ( .A(n25725), .B(n25727), .Z(n25721) );
  XOR U37057 ( .A(n25719), .B(n25721), .Z(n26894) );
  XOR U37058 ( .A(n26893), .B(n26894), .Z(n26898) );
  XOR U37059 ( .A(n26896), .B(n26898), .Z(n25715) );
  XOR U37060 ( .A(n25713), .B(n25715), .Z(n25718) );
  XOR U37061 ( .A(n25716), .B(n25718), .Z(n25708) );
  XOR U37062 ( .A(n25707), .B(n25708), .Z(n25711) );
  XOR U37063 ( .A(n25710), .B(n25711), .Z(n25703) );
  XOR U37064 ( .A(n25701), .B(n25703), .Z(n25706) );
  XOR U37065 ( .A(n25704), .B(n25706), .Z(n25696) );
  XOR U37066 ( .A(n25695), .B(n25696), .Z(n25700) );
  XOR U37067 ( .A(n25698), .B(n25700), .Z(n26904) );
  XOR U37068 ( .A(n26902), .B(n26904), .Z(n26906) );
  XOR U37069 ( .A(n26905), .B(n26906), .Z(n25693) );
  XOR U37070 ( .A(n25692), .B(n25693), .Z(n25687) );
  XOR U37071 ( .A(n25686), .B(n25687), .Z(n25691) );
  XOR U37072 ( .A(n25689), .B(n25691), .Z(n25682) );
  XOR U37073 ( .A(n25680), .B(n25682), .Z(n25684) );
  XOR U37074 ( .A(n25683), .B(n25684), .Z(n25679) );
  XOR U37075 ( .A(n25677), .B(n25679), .Z(n26913) );
  XOR U37076 ( .A(n26912), .B(n26913), .Z(n25676) );
  XOR U37077 ( .A(n25674), .B(n25676), .Z(n26919) );
  XOR U37078 ( .A(n26918), .B(n26919), .Z(n26922) );
  XOR U37079 ( .A(n26921), .B(n26922), .Z(n26926) );
  XOR U37080 ( .A(n26925), .B(n26926), .Z(n26930) );
  XOR U37081 ( .A(n26928), .B(n26930), .Z(n26933) );
  XOR U37082 ( .A(n26932), .B(n26933), .Z(n26937) );
  XOR U37083 ( .A(n26935), .B(n26937), .Z(n25670) );
  XOR U37084 ( .A(n25668), .B(n25670), .Z(n25672) );
  XOR U37085 ( .A(n25671), .B(n25672), .Z(n25666) );
  XOR U37086 ( .A(n25665), .B(n25666), .Z(n26943) );
  XOR U37087 ( .A(n26941), .B(n26943), .Z(n26946) );
  XOR U37088 ( .A(n26944), .B(n26946), .Z(n26949) );
  XOR U37089 ( .A(n26948), .B(n26949), .Z(n26952) );
  XOR U37090 ( .A(n26951), .B(n26952), .Z(n25664) );
  XOR U37091 ( .A(n25662), .B(n25664), .Z(n26956) );
  XOR U37092 ( .A(n26954), .B(n26956), .Z(n26959) );
  XOR U37093 ( .A(n26957), .B(n26959), .Z(n26962) );
  XOR U37094 ( .A(n26961), .B(n26962), .Z(n26965) );
  XOR U37095 ( .A(n26964), .B(n26965), .Z(n25661) );
  XOR U37096 ( .A(n25659), .B(n25661), .Z(n26970) );
  XOR U37097 ( .A(n26968), .B(n26970), .Z(n26972) );
  XOR U37098 ( .A(n26971), .B(n26972), .Z(n26977) );
  XOR U37099 ( .A(n26975), .B(n26977), .Z(n26980) );
  XOR U37100 ( .A(n26978), .B(n26980), .Z(n26983) );
  XOR U37101 ( .A(n26982), .B(n26983), .Z(n26986) );
  XOR U37102 ( .A(n26985), .B(n26986), .Z(n26990) );
  XOR U37103 ( .A(n26989), .B(n26990), .Z(n26994) );
  XOR U37104 ( .A(n26992), .B(n26994), .Z(n26998) );
  XOR U37105 ( .A(n26996), .B(n26998), .Z(n27001) );
  XOR U37106 ( .A(n26999), .B(n27001), .Z(n25655) );
  XOR U37107 ( .A(n25653), .B(n25655), .Z(n25658) );
  XOR U37108 ( .A(n25656), .B(n25658), .Z(n25652) );
  XOR U37109 ( .A(n25650), .B(n25652), .Z(n25645) );
  XOR U37110 ( .A(n25644), .B(n25645), .Z(n25649) );
  XOR U37111 ( .A(n25647), .B(n25649), .Z(n27014) );
  XOR U37112 ( .A(n27012), .B(n27014), .Z(n27016) );
  XOR U37113 ( .A(n27015), .B(n27016), .Z(n27019) );
  XOR U37114 ( .A(n27018), .B(n27019), .Z(n27023) );
  XOR U37115 ( .A(n27021), .B(n27023), .Z(n25640) );
  XOR U37116 ( .A(n25638), .B(n25640), .Z(n25642) );
  XOR U37117 ( .A(n25641), .B(n25642), .Z(n27025) );
  XOR U37118 ( .A(n27024), .B(n27025), .Z(n27029) );
  XOR U37119 ( .A(n27027), .B(n27029), .Z(n25637) );
  XOR U37120 ( .A(n25635), .B(n25637), .Z(n27033) );
  XOR U37121 ( .A(n27032), .B(n27033), .Z(n25633) );
  XOR U37122 ( .A(n25632), .B(n25633), .Z(n27041) );
  XOR U37123 ( .A(n27040), .B(n27041), .Z(n27045) );
  XOR U37124 ( .A(n27043), .B(n27045), .Z(n25628) );
  XOR U37125 ( .A(n25626), .B(n25628), .Z(n25630) );
  XOR U37126 ( .A(n25629), .B(n25630), .Z(n25625) );
  XOR U37127 ( .A(n25623), .B(n25625), .Z(n27050) );
  XOR U37128 ( .A(n27048), .B(n27050), .Z(n28643) );
  XOR U37129 ( .A(n27051), .B(n28643), .Z(n27055) );
  XOR U37130 ( .A(n27054), .B(n27055), .Z(n27058) );
  XOR U37131 ( .A(n27057), .B(n27058), .Z(n27062) );
  XOR U37132 ( .A(n27061), .B(n27062), .Z(n27066) );
  XOR U37133 ( .A(n27064), .B(n27066), .Z(n25619) );
  XOR U37134 ( .A(n25617), .B(n25619), .Z(n25622) );
  XOR U37135 ( .A(n25620), .B(n25622), .Z(n25616) );
  XOR U37136 ( .A(n25614), .B(n25616), .Z(n27070) );
  XOR U37137 ( .A(n27068), .B(n27070), .Z(n27072) );
  XOR U37138 ( .A(n27071), .B(n27072), .Z(n27077) );
  XOR U37139 ( .A(n27075), .B(n27077), .Z(n27080) );
  XOR U37140 ( .A(n27078), .B(n27080), .Z(n27082) );
  XOR U37141 ( .A(n27081), .B(n27082), .Z(n27085) );
  XOR U37142 ( .A(n27084), .B(n27085), .Z(n27089) );
  XOR U37143 ( .A(n27088), .B(n27089), .Z(n27093) );
  XOR U37144 ( .A(n27091), .B(n27093), .Z(n25610) );
  XOR U37145 ( .A(n25608), .B(n25610), .Z(n25612) );
  XOR U37146 ( .A(n25611), .B(n25612), .Z(n25604) );
  XOR U37147 ( .A(n25602), .B(n25604), .Z(n25606) );
  XOR U37148 ( .A(n25605), .B(n25606), .Z(n27097) );
  XOR U37149 ( .A(n27096), .B(n27097), .Z(n27100) );
  XOR U37150 ( .A(n27099), .B(n27100), .Z(n25598) );
  XOR U37151 ( .A(n25596), .B(n25598), .Z(n25601) );
  XOR U37152 ( .A(n25599), .B(n25601), .Z(n25592) );
  XOR U37153 ( .A(n25590), .B(n25592), .Z(n25594) );
  XOR U37154 ( .A(n25593), .B(n25594), .Z(n25586) );
  XOR U37155 ( .A(n25584), .B(n25586), .Z(n25589) );
  XOR U37156 ( .A(n25587), .B(n25589), .Z(n27106) );
  XOR U37157 ( .A(n27105), .B(n27106), .Z(n27109) );
  XOR U37158 ( .A(n27108), .B(n27109), .Z(n25579) );
  XOR U37159 ( .A(n25578), .B(n25579), .Z(n25583) );
  XOR U37160 ( .A(n25581), .B(n25583), .Z(n27115) );
  XOR U37161 ( .A(n27113), .B(n27115), .Z(n27117) );
  XOR U37162 ( .A(n27116), .B(n27117), .Z(n25574) );
  XOR U37163 ( .A(n25572), .B(n25574), .Z(n25577) );
  XOR U37164 ( .A(n25575), .B(n25577), .Z(n27121) );
  XOR U37165 ( .A(n27120), .B(n27121), .Z(n27124) );
  XOR U37166 ( .A(n27123), .B(n27124), .Z(n25570) );
  XOR U37167 ( .A(n25569), .B(n25570), .Z(n27130) );
  XOR U37168 ( .A(n27128), .B(n27130), .Z(n25568) );
  XOR U37169 ( .A(n25566), .B(n25568), .Z(n25561) );
  XOR U37170 ( .A(n25560), .B(n25561), .Z(n25565) );
  XOR U37171 ( .A(n25563), .B(n25565), .Z(n27141) );
  XOR U37172 ( .A(n27139), .B(n27141), .Z(n27144) );
  XOR U37173 ( .A(n27142), .B(n27144), .Z(n25558) );
  XOR U37174 ( .A(n25557), .B(n25558), .Z(n25552) );
  XOR U37175 ( .A(n25551), .B(n25552), .Z(n25556) );
  XOR U37176 ( .A(n25554), .B(n25556), .Z(n25547) );
  XOR U37177 ( .A(n25545), .B(n25547), .Z(n25549) );
  XOR U37178 ( .A(n25548), .B(n25549), .Z(n25541) );
  XOR U37179 ( .A(n25539), .B(n25541), .Z(n25544) );
  XOR U37180 ( .A(n25542), .B(n25544), .Z(n27148) );
  XOR U37181 ( .A(n27147), .B(n27148), .Z(n27151) );
  XOR U37182 ( .A(n27150), .B(n27151), .Z(n27155) );
  XOR U37183 ( .A(n27154), .B(n27155), .Z(n27159) );
  XOR U37184 ( .A(n27157), .B(n27159), .Z(n27162) );
  XOR U37185 ( .A(n27160), .B(n27162), .Z(n27164) );
  XOR U37186 ( .A(n27163), .B(n27164), .Z(n25538) );
  XOR U37187 ( .A(n25536), .B(n25538), .Z(n27173) );
  XOR U37188 ( .A(n27171), .B(n27173), .Z(n25534) );
  XOR U37189 ( .A(n25532), .B(n25534), .Z(n27168) );
  XOR U37190 ( .A(n27167), .B(n27168), .Z(n25528) );
  XOR U37191 ( .A(n25526), .B(n25528), .Z(n25531) );
  XOR U37192 ( .A(n25529), .B(n25531), .Z(n25520) );
  XOR U37193 ( .A(n25519), .B(n25520), .Z(n25523) );
  XOR U37194 ( .A(n25522), .B(n25523), .Z(n27182) );
  XOR U37195 ( .A(n27180), .B(n27182), .Z(n27185) );
  XOR U37196 ( .A(n27183), .B(n27185), .Z(n25514) );
  XOR U37197 ( .A(n25513), .B(n25514), .Z(n25517) );
  XOR U37198 ( .A(n25516), .B(n25517), .Z(n25509) );
  XOR U37199 ( .A(n25507), .B(n25509), .Z(n25512) );
  XOR U37200 ( .A(n25510), .B(n25512), .Z(n25506) );
  XOR U37201 ( .A(n25504), .B(n25506), .Z(n25500) );
  XOR U37202 ( .A(n25498), .B(n25500), .Z(n25503) );
  XOR U37203 ( .A(n25501), .B(n25503), .Z(n27191) );
  XOR U37204 ( .A(n27189), .B(n27191), .Z(n27193) );
  XOR U37205 ( .A(n27192), .B(n27193), .Z(n25496) );
  XOR U37206 ( .A(n25495), .B(n25496), .Z(n25490) );
  XOR U37207 ( .A(n25489), .B(n25490), .Z(n25494) );
  XOR U37208 ( .A(n25492), .B(n25494), .Z(n25484) );
  XOR U37209 ( .A(n25483), .B(n25484), .Z(n25487) );
  XOR U37210 ( .A(n25486), .B(n25487), .Z(n27202) );
  XOR U37211 ( .A(n27200), .B(n27202), .Z(n25481) );
  XOR U37212 ( .A(n25479), .B(n25481), .Z(n27198) );
  XOR U37213 ( .A(n27196), .B(n27198), .Z(n25474) );
  XOR U37214 ( .A(n25473), .B(n25474), .Z(n25477) );
  XOR U37215 ( .A(n25476), .B(n25477), .Z(n25469) );
  XOR U37216 ( .A(n25467), .B(n25469), .Z(n25471) );
  XOR U37217 ( .A(n25470), .B(n25471), .Z(n25461) );
  XOR U37218 ( .A(n25460), .B(n25461), .Z(n25464) );
  XOR U37219 ( .A(n25463), .B(n25464), .Z(n25456) );
  XOR U37220 ( .A(n25454), .B(n25456), .Z(n25459) );
  XOR U37221 ( .A(n25457), .B(n25459), .Z(n25449) );
  XOR U37222 ( .A(n25448), .B(n25449), .Z(n25452) );
  XOR U37223 ( .A(n25451), .B(n25452), .Z(n27212) );
  XOR U37224 ( .A(n27210), .B(n27212), .Z(n27214) );
  XOR U37225 ( .A(n27213), .B(n27214), .Z(n27220) );
  XOR U37226 ( .A(n27219), .B(n27220), .Z(n25447) );
  XOR U37227 ( .A(n25445), .B(n25447), .Z(n25443) );
  XOR U37228 ( .A(n25441), .B(n25443), .Z(n25437) );
  XOR U37229 ( .A(n25435), .B(n25437), .Z(n25439) );
  XOR U37230 ( .A(n25438), .B(n25439), .Z(n25431) );
  XOR U37231 ( .A(n25429), .B(n25431), .Z(n25434) );
  XOR U37232 ( .A(n25432), .B(n25434), .Z(n25428) );
  XOR U37233 ( .A(n25426), .B(n25428), .Z(n25420) );
  XOR U37234 ( .A(n25419), .B(n25420), .Z(n25424) );
  XOR U37235 ( .A(n25422), .B(n25424), .Z(n25415) );
  XOR U37236 ( .A(n25413), .B(n25415), .Z(n25418) );
  XOR U37237 ( .A(n25416), .B(n25418), .Z(n25408) );
  XOR U37238 ( .A(n25407), .B(n25408), .Z(n25411) );
  XOR U37239 ( .A(n25410), .B(n25411), .Z(n25406) );
  XOR U37240 ( .A(n25404), .B(n25406), .Z(n25400) );
  XOR U37241 ( .A(n25398), .B(n25400), .Z(n25402) );
  XOR U37242 ( .A(n25401), .B(n25402), .Z(n25394) );
  XOR U37243 ( .A(n25392), .B(n25394), .Z(n25397) );
  XOR U37244 ( .A(n25395), .B(n25397), .Z(n25388) );
  XOR U37245 ( .A(n25386), .B(n25388), .Z(n25390) );
  XOR U37246 ( .A(n25389), .B(n25390), .Z(n25381) );
  XOR U37247 ( .A(n25380), .B(n25381), .Z(n25385) );
  XOR U37248 ( .A(n25383), .B(n25385), .Z(n25379) );
  XOR U37249 ( .A(n25377), .B(n25379), .Z(n27234) );
  XOR U37250 ( .A(n27233), .B(n27234), .Z(n27238) );
  XOR U37251 ( .A(n27236), .B(n27238), .Z(n27242) );
  XOR U37252 ( .A(n27240), .B(n27242), .Z(n27245) );
  XOR U37253 ( .A(n27243), .B(n27245), .Z(n25375) );
  XOR U37254 ( .A(n25374), .B(n25375), .Z(n25368) );
  XOR U37255 ( .A(n25367), .B(n25368), .Z(n25372) );
  XOR U37256 ( .A(n25370), .B(n25372), .Z(n25363) );
  XOR U37257 ( .A(n25361), .B(n25363), .Z(n25365) );
  XOR U37258 ( .A(n25364), .B(n25365), .Z(n27249) );
  XOR U37259 ( .A(n27247), .B(n27249), .Z(n27252) );
  XOR U37260 ( .A(n27250), .B(n27252), .Z(n25360) );
  XOR U37261 ( .A(n25358), .B(n25360), .Z(n27258) );
  XOR U37262 ( .A(n27257), .B(n27258), .Z(n25356) );
  XOR U37263 ( .A(n25355), .B(n25356), .Z(n25351) );
  XOR U37264 ( .A(n25349), .B(n25351), .Z(n25354) );
  XOR U37265 ( .A(n25352), .B(n25354), .Z(n27265) );
  XOR U37266 ( .A(n27264), .B(n27265), .Z(n27269) );
  XOR U37267 ( .A(n27267), .B(n27269), .Z(n25345) );
  XOR U37268 ( .A(n25343), .B(n25345), .Z(n25348) );
  XOR U37269 ( .A(n25346), .B(n25348), .Z(n27272) );
  XOR U37270 ( .A(n27271), .B(n27272), .Z(n27275) );
  XOR U37271 ( .A(n27274), .B(n27275), .Z(n25339) );
  XOR U37272 ( .A(n25337), .B(n25339), .Z(n25342) );
  XOR U37273 ( .A(n25340), .B(n25342), .Z(n27280) );
  XOR U37274 ( .A(n27279), .B(n27280), .Z(n27284) );
  XOR U37275 ( .A(n27282), .B(n27284), .Z(n27291) );
  XOR U37276 ( .A(n27289), .B(n27291), .Z(n25335) );
  XOR U37277 ( .A(n25333), .B(n25335), .Z(n27286) );
  XOR U37278 ( .A(n27285), .B(n27286), .Z(n25329) );
  XOR U37279 ( .A(n25327), .B(n25329), .Z(n25332) );
  XOR U37280 ( .A(n25330), .B(n25332), .Z(n25323) );
  XOR U37281 ( .A(n25321), .B(n25323), .Z(n25325) );
  XOR U37282 ( .A(n25324), .B(n25325), .Z(n25317) );
  XOR U37283 ( .A(n25315), .B(n25317), .Z(n25319) );
  XOR U37284 ( .A(n25318), .B(n25319), .Z(n25314) );
  XOR U37285 ( .A(n25312), .B(n25314), .Z(n25308) );
  XOR U37286 ( .A(n25306), .B(n25308), .Z(n25311) );
  XOR U37287 ( .A(n25309), .B(n25311), .Z(n25302) );
  XOR U37288 ( .A(n25300), .B(n25302), .Z(n25305) );
  XOR U37289 ( .A(n25303), .B(n25305), .Z(n25295) );
  XOR U37290 ( .A(n25294), .B(n25295), .Z(n25299) );
  XOR U37291 ( .A(n25297), .B(n25299), .Z(n25289) );
  XOR U37292 ( .A(n25288), .B(n25289), .Z(n25293) );
  XOR U37293 ( .A(n25291), .B(n25293), .Z(n27299) );
  XOR U37294 ( .A(n27298), .B(n27299), .Z(n27302) );
  XOR U37295 ( .A(n27301), .B(n27302), .Z(n27309) );
  XOR U37296 ( .A(n27307), .B(n27309), .Z(n25287) );
  XOR U37297 ( .A(n25285), .B(n25287), .Z(n25281) );
  XOR U37298 ( .A(n25279), .B(n25281), .Z(n25284) );
  XOR U37299 ( .A(n25282), .B(n25284), .Z(n25275) );
  XOR U37300 ( .A(n25273), .B(n25275), .Z(n25277) );
  XOR U37301 ( .A(n25276), .B(n25277), .Z(n25268) );
  XOR U37302 ( .A(n25267), .B(n25268), .Z(n25272) );
  XOR U37303 ( .A(n25270), .B(n25272), .Z(n27321) );
  XOR U37304 ( .A(n27319), .B(n27321), .Z(n27323) );
  XOR U37305 ( .A(n27322), .B(n27323), .Z(n25262) );
  XOR U37306 ( .A(n25261), .B(n25262), .Z(n25265) );
  XOR U37307 ( .A(n25264), .B(n25265), .Z(n27327) );
  XOR U37308 ( .A(n27326), .B(n27327), .Z(n27331) );
  XOR U37309 ( .A(n27329), .B(n27331), .Z(n27334) );
  XOR U37310 ( .A(n27333), .B(n27334), .Z(n27338) );
  XOR U37311 ( .A(n27336), .B(n27338), .Z(n27342) );
  XOR U37312 ( .A(n27340), .B(n27342), .Z(n27344) );
  XOR U37313 ( .A(n27343), .B(n27344), .Z(n25256) );
  XOR U37314 ( .A(n25255), .B(n25256), .Z(n25260) );
  XOR U37315 ( .A(n25258), .B(n25260), .Z(n27349) );
  XOR U37316 ( .A(n27347), .B(n27349), .Z(n27352) );
  XOR U37317 ( .A(n27350), .B(n27352), .Z(n25250) );
  XOR U37318 ( .A(n25249), .B(n25250), .Z(n25253) );
  XOR U37319 ( .A(n25252), .B(n25253), .Z(n27355) );
  XOR U37320 ( .A(n27353), .B(n27355), .Z(n27358) );
  XOR U37321 ( .A(n27356), .B(n27358), .Z(n27363) );
  XOR U37322 ( .A(n27362), .B(n27363), .Z(n25248) );
  XOR U37323 ( .A(n25246), .B(n25248), .Z(n27374) );
  XOR U37324 ( .A(n27372), .B(n27374), .Z(n27377) );
  XOR U37325 ( .A(n27375), .B(n27377), .Z(n27380) );
  XOR U37326 ( .A(n27379), .B(n27380), .Z(n27383) );
  XOR U37327 ( .A(n27382), .B(n27383), .Z(n27388) );
  XOR U37328 ( .A(n27386), .B(n27388), .Z(n27391) );
  XOR U37329 ( .A(n27389), .B(n27391), .Z(n25242) );
  XOR U37330 ( .A(n25240), .B(n25242), .Z(n25245) );
  XOR U37331 ( .A(n25243), .B(n25245), .Z(n25239) );
  XOR U37332 ( .A(n25237), .B(n25239), .Z(n27396) );
  XOR U37333 ( .A(n27394), .B(n27396), .Z(n27398) );
  XOR U37334 ( .A(n27397), .B(n27398), .Z(n27402) );
  XOR U37335 ( .A(n27401), .B(n27402), .Z(n27406) );
  XOR U37336 ( .A(n27404), .B(n27406), .Z(n27409) );
  XOR U37337 ( .A(n27407), .B(n27409), .Z(n27411) );
  XOR U37338 ( .A(n27410), .B(n27411), .Z(n25235) );
  XOR U37339 ( .A(n25233), .B(n25235), .Z(n27418) );
  XOR U37340 ( .A(n27416), .B(n27418), .Z(n25231) );
  XOR U37341 ( .A(n25230), .B(n25231), .Z(n25225) );
  XOR U37342 ( .A(n25224), .B(n25225), .Z(n25229) );
  XOR U37343 ( .A(n25227), .B(n25229), .Z(n25223) );
  XOR U37344 ( .A(n25221), .B(n25223), .Z(n27429) );
  XOR U37345 ( .A(n27427), .B(n27429), .Z(n27431) );
  XOR U37346 ( .A(n27430), .B(n27431), .Z(n25219) );
  XOR U37347 ( .A(n25218), .B(n25219), .Z(n25214) );
  XOR U37348 ( .A(n25212), .B(n25214), .Z(n25217) );
  XOR U37349 ( .A(n25215), .B(n25217), .Z(n25207) );
  XOR U37350 ( .A(n25206), .B(n25207), .Z(n25210) );
  XOR U37351 ( .A(n25209), .B(n25210), .Z(n25205) );
  XOR U37352 ( .A(n25203), .B(n25205), .Z(n25199) );
  XOR U37353 ( .A(n25197), .B(n25199), .Z(n25201) );
  XOR U37354 ( .A(n25200), .B(n25201), .Z(n25193) );
  XOR U37355 ( .A(n25191), .B(n25193), .Z(n25196) );
  XOR U37356 ( .A(n25194), .B(n25196), .Z(n25189) );
  XOR U37357 ( .A(n25188), .B(n25189), .Z(n27442) );
  XOR U37358 ( .A(n27441), .B(n27442), .Z(n25187) );
  XOR U37359 ( .A(n25185), .B(n25187), .Z(n25181) );
  XOR U37360 ( .A(n25179), .B(n25181), .Z(n25184) );
  XOR U37361 ( .A(n25182), .B(n25184), .Z(n25174) );
  XOR U37362 ( .A(n25173), .B(n25174), .Z(n25178) );
  XOR U37363 ( .A(n25176), .B(n25178), .Z(n25169) );
  XOR U37364 ( .A(n25167), .B(n25169), .Z(n25172) );
  XOR U37365 ( .A(n25170), .B(n25172), .Z(n27449) );
  XOR U37366 ( .A(n27448), .B(n27449), .Z(n27453) );
  XOR U37367 ( .A(n27451), .B(n27453), .Z(n27457) );
  XOR U37368 ( .A(n27455), .B(n27457), .Z(n27460) );
  XOR U37369 ( .A(n27458), .B(n27460), .Z(n27463) );
  XOR U37370 ( .A(n27461), .B(n27463), .Z(n27466) );
  XOR U37371 ( .A(n27464), .B(n27466), .Z(n25163) );
  XOR U37372 ( .A(n25161), .B(n25163), .Z(n25166) );
  XOR U37373 ( .A(n25164), .B(n25166), .Z(n27468) );
  XOR U37374 ( .A(n27467), .B(n27468), .Z(n27471) );
  XOR U37375 ( .A(n27470), .B(n27471), .Z(n25157) );
  XOR U37376 ( .A(n25155), .B(n25157), .Z(n25160) );
  XOR U37377 ( .A(n25158), .B(n25160), .Z(n25150) );
  XOR U37378 ( .A(n25149), .B(n25150), .Z(n25154) );
  XOR U37379 ( .A(n25152), .B(n25154), .Z(n25145) );
  XOR U37380 ( .A(n25143), .B(n25145), .Z(n25148) );
  XOR U37381 ( .A(n25146), .B(n25148), .Z(n27477) );
  XOR U37382 ( .A(n27475), .B(n27477), .Z(n27480) );
  XOR U37383 ( .A(n27478), .B(n27480), .Z(n25138) );
  XOR U37384 ( .A(n25137), .B(n25138), .Z(n25142) );
  XOR U37385 ( .A(n25140), .B(n25142), .Z(n25135) );
  XOR U37386 ( .A(n25133), .B(n25135), .Z(n25132) );
  XOR U37387 ( .A(n25130), .B(n25132), .Z(n27484) );
  XOR U37388 ( .A(n27482), .B(n27484), .Z(n27488) );
  XOR U37389 ( .A(n27486), .B(n27488), .Z(n27500) );
  XOR U37390 ( .A(n27498), .B(n27500), .Z(n27502) );
  XOR U37391 ( .A(n27501), .B(n27502), .Z(n25125) );
  XOR U37392 ( .A(n25124), .B(n25125), .Z(n25128) );
  XOR U37393 ( .A(n25127), .B(n25128), .Z(n25120) );
  XOR U37394 ( .A(n25118), .B(n25120), .Z(n25123) );
  XOR U37395 ( .A(n25121), .B(n25123), .Z(n25113) );
  XOR U37396 ( .A(n25112), .B(n25113), .Z(n25117) );
  XOR U37397 ( .A(n25115), .B(n25117), .Z(n25107) );
  XOR U37398 ( .A(n25106), .B(n25107), .Z(n25111) );
  XOR U37399 ( .A(n25109), .B(n25111), .Z(n25105) );
  XOR U37400 ( .A(n25103), .B(n25105), .Z(n25098) );
  XOR U37401 ( .A(n25097), .B(n25098), .Z(n25101) );
  XOR U37402 ( .A(n25100), .B(n25101), .Z(n25096) );
  XOR U37403 ( .A(n25094), .B(n25096), .Z(n27512) );
  XOR U37404 ( .A(n27510), .B(n27512), .Z(n27515) );
  XOR U37405 ( .A(n27513), .B(n27515), .Z(n25089) );
  XOR U37406 ( .A(n25088), .B(n25089), .Z(n25092) );
  XOR U37407 ( .A(n25091), .B(n25092), .Z(n25087) );
  XOR U37408 ( .A(n25085), .B(n25087), .Z(n27519) );
  XOR U37409 ( .A(n27518), .B(n27519), .Z(n27522) );
  XOR U37410 ( .A(n27521), .B(n27522), .Z(n25084) );
  XOR U37411 ( .A(n25082), .B(n25084), .Z(n25077) );
  XOR U37412 ( .A(n25076), .B(n25077), .Z(n25080) );
  XOR U37413 ( .A(n25079), .B(n25080), .Z(n25071) );
  XOR U37414 ( .A(n25070), .B(n25071), .Z(n25074) );
  XOR U37415 ( .A(n25073), .B(n25074), .Z(n25066) );
  XOR U37416 ( .A(n25064), .B(n25066), .Z(n25069) );
  XOR U37417 ( .A(n25067), .B(n25069), .Z(n25060) );
  XOR U37418 ( .A(n25058), .B(n25060), .Z(n25063) );
  XOR U37419 ( .A(n25061), .B(n25063), .Z(n25054) );
  XOR U37420 ( .A(n25052), .B(n25054), .Z(n25057) );
  XOR U37421 ( .A(n25055), .B(n25057), .Z(n25050) );
  XOR U37422 ( .A(n25049), .B(n25050), .Z(n27531) );
  XOR U37423 ( .A(n27530), .B(n27531), .Z(n27535) );
  XOR U37424 ( .A(n27533), .B(n27535), .Z(n27539) );
  XOR U37425 ( .A(n27538), .B(n27539), .Z(n27542) );
  XOR U37426 ( .A(n27541), .B(n27542), .Z(n25048) );
  XOR U37427 ( .A(n25046), .B(n25048), .Z(n27548) );
  XOR U37428 ( .A(n27547), .B(n27548), .Z(n25045) );
  XOR U37429 ( .A(n25043), .B(n25045), .Z(n27557) );
  XOR U37430 ( .A(n27556), .B(n27557), .Z(n25041) );
  XOR U37431 ( .A(n25040), .B(n25041), .Z(n27571) );
  XOR U37432 ( .A(n27570), .B(n27571), .Z(n27569) );
  XOR U37433 ( .A(n27567), .B(n27569), .Z(n25035) );
  XOR U37434 ( .A(n25034), .B(n25035), .Z(n25039) );
  XOR U37435 ( .A(n25037), .B(n25039), .Z(n25029) );
  XOR U37436 ( .A(n25027), .B(n25029), .Z(n25031) );
  XOR U37437 ( .A(n25030), .B(n25031), .Z(n25025) );
  XOR U37438 ( .A(n25024), .B(n25025), .Z(n25019) );
  XOR U37439 ( .A(n25018), .B(n25019), .Z(n25023) );
  XOR U37440 ( .A(n25021), .B(n25023), .Z(n25014) );
  XOR U37441 ( .A(n25012), .B(n25014), .Z(n25016) );
  XOR U37442 ( .A(n25015), .B(n25016), .Z(n25011) );
  XOR U37443 ( .A(n25009), .B(n25011), .Z(n27592) );
  XOR U37444 ( .A(n27590), .B(n27592), .Z(n25007) );
  XOR U37445 ( .A(n25005), .B(n25007), .Z(n27587) );
  XOR U37446 ( .A(n27586), .B(n27587), .Z(n25000) );
  XOR U37447 ( .A(n24999), .B(n25000), .Z(n25004) );
  XOR U37448 ( .A(n25002), .B(n25004), .Z(n24995) );
  XOR U37449 ( .A(n24993), .B(n24995), .Z(n24997) );
  XOR U37450 ( .A(n24996), .B(n24997), .Z(n24988) );
  XOR U37451 ( .A(n24987), .B(n24988), .Z(n24992) );
  XOR U37452 ( .A(n24990), .B(n24992), .Z(n24983) );
  XOR U37453 ( .A(n24981), .B(n24983), .Z(n24985) );
  XOR U37454 ( .A(n24984), .B(n24985), .Z(n27600) );
  XOR U37455 ( .A(n27599), .B(n27600), .Z(n27604) );
  XOR U37456 ( .A(n27602), .B(n27604), .Z(n24977) );
  XOR U37457 ( .A(n24975), .B(n24977), .Z(n24979) );
  XOR U37458 ( .A(n24978), .B(n24979), .Z(n27608) );
  XOR U37459 ( .A(n27606), .B(n27608), .Z(n27611) );
  XOR U37460 ( .A(n27609), .B(n27611), .Z(n24971) );
  XOR U37461 ( .A(n24969), .B(n24971), .Z(n24973) );
  XOR U37462 ( .A(n24972), .B(n24973), .Z(n27614) );
  XOR U37463 ( .A(n27613), .B(n27614), .Z(n27618) );
  XOR U37464 ( .A(n27616), .B(n27618), .Z(n24968) );
  XOR U37465 ( .A(n24966), .B(n24968), .Z(n24961) );
  XOR U37466 ( .A(n24960), .B(n24961), .Z(n24965) );
  XOR U37467 ( .A(n24963), .B(n24965), .Z(n24956) );
  XOR U37468 ( .A(n24954), .B(n24956), .Z(n24959) );
  XOR U37469 ( .A(n24957), .B(n24959), .Z(n27622) );
  XOR U37470 ( .A(n27621), .B(n27622), .Z(n27625) );
  XOR U37471 ( .A(n27624), .B(n27625), .Z(n24953) );
  XOR U37472 ( .A(n24951), .B(n24953), .Z(n24949) );
  XOR U37473 ( .A(n24947), .B(n24949), .Z(n24942) );
  XOR U37474 ( .A(n24941), .B(n24942), .Z(n24945) );
  XOR U37475 ( .A(n24944), .B(n24945), .Z(n24937) );
  XOR U37476 ( .A(n24935), .B(n24937), .Z(n24940) );
  XOR U37477 ( .A(n24938), .B(n24940), .Z(n24930) );
  XOR U37478 ( .A(n24929), .B(n24930), .Z(n24934) );
  XOR U37479 ( .A(n24932), .B(n24934), .Z(n27638) );
  XOR U37480 ( .A(n27636), .B(n27638), .Z(n27640) );
  XOR U37481 ( .A(n27639), .B(n27640), .Z(n27644) );
  XOR U37482 ( .A(n27643), .B(n27644), .Z(n27648) );
  XOR U37483 ( .A(n27646), .B(n27648), .Z(n24925) );
  XOR U37484 ( .A(n24923), .B(n24925), .Z(n24927) );
  XOR U37485 ( .A(n24926), .B(n24927), .Z(n24918) );
  XOR U37486 ( .A(n24917), .B(n24918), .Z(n24922) );
  XOR U37487 ( .A(n24920), .B(n24922), .Z(n24912) );
  XOR U37488 ( .A(n24911), .B(n24912), .Z(n24916) );
  XOR U37489 ( .A(n24914), .B(n24916), .Z(n24906) );
  XOR U37490 ( .A(n24905), .B(n24906), .Z(n24910) );
  XOR U37491 ( .A(n24908), .B(n24910), .Z(n27654) );
  XOR U37492 ( .A(n27652), .B(n27654), .Z(n27657) );
  XOR U37493 ( .A(n27655), .B(n27657), .Z(n27661) );
  XOR U37494 ( .A(n27659), .B(n27661), .Z(n27663) );
  XOR U37495 ( .A(n27662), .B(n27663), .Z(n24903) );
  XOR U37496 ( .A(n24902), .B(n24903), .Z(n24898) );
  XOR U37497 ( .A(n24896), .B(n24898), .Z(n24901) );
  XOR U37498 ( .A(n24899), .B(n24901), .Z(n27668) );
  XOR U37499 ( .A(n27666), .B(n27668), .Z(n27671) );
  XOR U37500 ( .A(n27669), .B(n27671), .Z(n24894) );
  XOR U37501 ( .A(n24893), .B(n24894), .Z(n27674) );
  XOR U37502 ( .A(n27673), .B(n27674), .Z(n27677) );
  XOR U37503 ( .A(n27676), .B(n27677), .Z(n24889) );
  XOR U37504 ( .A(n24887), .B(n24889), .Z(n24892) );
  XOR U37505 ( .A(n24890), .B(n24892), .Z(n24883) );
  XOR U37506 ( .A(n24881), .B(n24883), .Z(n24886) );
  XOR U37507 ( .A(n24884), .B(n24886), .Z(n24877) );
  XOR U37508 ( .A(n24875), .B(n24877), .Z(n24880) );
  XOR U37509 ( .A(n24878), .B(n24880), .Z(n24869) );
  XOR U37510 ( .A(n24868), .B(n24869), .Z(n24872) );
  XOR U37511 ( .A(n24871), .B(n24872), .Z(n24863) );
  XOR U37512 ( .A(n24861), .B(n24863), .Z(n24866) );
  XOR U37513 ( .A(n24864), .B(n24866), .Z(n24856) );
  XOR U37514 ( .A(n24855), .B(n24856), .Z(n24860) );
  XOR U37515 ( .A(n24858), .B(n24860), .Z(n24851) );
  XOR U37516 ( .A(n24849), .B(n24851), .Z(n24854) );
  XOR U37517 ( .A(n24852), .B(n24854), .Z(n27682) );
  XOR U37518 ( .A(n27681), .B(n27682), .Z(n27685) );
  XOR U37519 ( .A(n27684), .B(n27685), .Z(n24845) );
  XOR U37520 ( .A(n24843), .B(n24845), .Z(n24848) );
  XOR U37521 ( .A(n24846), .B(n24848), .Z(n27690) );
  XOR U37522 ( .A(n27689), .B(n27690), .Z(n27694) );
  XOR U37523 ( .A(n27692), .B(n27694), .Z(n27698) );
  XOR U37524 ( .A(n27696), .B(n27698), .Z(n27700) );
  XOR U37525 ( .A(n27699), .B(n27700), .Z(n27703) );
  XOR U37526 ( .A(n27702), .B(n27703), .Z(n27707) );
  XOR U37527 ( .A(n27705), .B(n27707), .Z(n24841) );
  XOR U37528 ( .A(n24840), .B(n24841), .Z(n24836) );
  XOR U37529 ( .A(n24834), .B(n24836), .Z(n24838) );
  XOR U37530 ( .A(n24837), .B(n24838), .Z(n24830) );
  XOR U37531 ( .A(n24828), .B(n24830), .Z(n24833) );
  XOR U37532 ( .A(n24831), .B(n24833), .Z(n24827) );
  XOR U37533 ( .A(n24825), .B(n24827), .Z(n27712) );
  XOR U37534 ( .A(n27711), .B(n27712), .Z(n24823) );
  XOR U37535 ( .A(n24822), .B(n24823), .Z(n24818) );
  XOR U37536 ( .A(n24816), .B(n24818), .Z(n24821) );
  XOR U37537 ( .A(n24819), .B(n24821), .Z(n24811) );
  XOR U37538 ( .A(n24810), .B(n24811), .Z(n24815) );
  XOR U37539 ( .A(n24813), .B(n24815), .Z(n24806) );
  XOR U37540 ( .A(n24804), .B(n24806), .Z(n24809) );
  XOR U37541 ( .A(n24807), .B(n24809), .Z(n24799) );
  XOR U37542 ( .A(n24798), .B(n24799), .Z(n24802) );
  XOR U37543 ( .A(n24801), .B(n24802), .Z(n24796) );
  XOR U37544 ( .A(n24794), .B(n24796), .Z(n24790) );
  XOR U37545 ( .A(n24788), .B(n24790), .Z(n24792) );
  XOR U37546 ( .A(n24791), .B(n24792), .Z(n24784) );
  XOR U37547 ( .A(n24782), .B(n24784), .Z(n24787) );
  XOR U37548 ( .A(n24785), .B(n24787), .Z(n24778) );
  XOR U37549 ( .A(n24776), .B(n24778), .Z(n24780) );
  XOR U37550 ( .A(n24779), .B(n24780), .Z(n24771) );
  XOR U37551 ( .A(n24770), .B(n24771), .Z(n24775) );
  XOR U37552 ( .A(n24773), .B(n24775), .Z(n24768) );
  XOR U37553 ( .A(n24767), .B(n24768), .Z(n24761) );
  XOR U37554 ( .A(n24760), .B(n24761), .Z(n24765) );
  XOR U37555 ( .A(n24763), .B(n24765), .Z(n27726) );
  XOR U37556 ( .A(n27724), .B(n27726), .Z(n27729) );
  XOR U37557 ( .A(n27727), .B(n27729), .Z(n24755) );
  XOR U37558 ( .A(n24754), .B(n24755), .Z(n24759) );
  XOR U37559 ( .A(n24757), .B(n24759), .Z(n24752) );
  XOR U37560 ( .A(n24751), .B(n24752), .Z(n27734) );
  XOR U37561 ( .A(n27733), .B(n27734), .Z(n27738) );
  XOR U37562 ( .A(n27736), .B(n27738), .Z(n27751) );
  XOR U37563 ( .A(n27749), .B(n27751), .Z(n27754) );
  XOR U37564 ( .A(n27752), .B(n27754), .Z(n24750) );
  XOR U37565 ( .A(n24748), .B(n24750), .Z(n24743) );
  XOR U37566 ( .A(n24742), .B(n24743), .Z(n24746) );
  XOR U37567 ( .A(n24745), .B(n24746), .Z(n24738) );
  XOR U37568 ( .A(n24736), .B(n24738), .Z(n24741) );
  XOR U37569 ( .A(n24739), .B(n24741), .Z(n24731) );
  XOR U37570 ( .A(n24730), .B(n24731), .Z(n24735) );
  XOR U37571 ( .A(n24733), .B(n24735), .Z(n24726) );
  XOR U37572 ( .A(n24724), .B(n24726), .Z(n24728) );
  XOR U37573 ( .A(n24727), .B(n24728), .Z(n27761) );
  XOR U37574 ( .A(n27760), .B(n27761), .Z(n27764) );
  XOR U37575 ( .A(n27763), .B(n27764), .Z(n24723) );
  XOR U37576 ( .A(n24721), .B(n24723), .Z(n27773) );
  XOR U37577 ( .A(n27772), .B(n27773), .Z(n27776) );
  XOR U37578 ( .A(n27775), .B(n27776), .Z(n24717) );
  XOR U37579 ( .A(n24715), .B(n24717), .Z(n24720) );
  XOR U37580 ( .A(n24718), .B(n24720), .Z(n24711) );
  XOR U37581 ( .A(n24709), .B(n24711), .Z(n24713) );
  XOR U37582 ( .A(n24712), .B(n24713), .Z(n24707) );
  XOR U37583 ( .A(n24706), .B(n24707), .Z(n24701) );
  XOR U37584 ( .A(n24699), .B(n24701), .Z(n24704) );
  XOR U37585 ( .A(n24702), .B(n24704), .Z(n24694) );
  XOR U37586 ( .A(n24693), .B(n24694), .Z(n24698) );
  XOR U37587 ( .A(n24696), .B(n24698), .Z(n24689) );
  XOR U37588 ( .A(n24687), .B(n24689), .Z(n24692) );
  XOR U37589 ( .A(n24690), .B(n24692), .Z(n24685) );
  XOR U37590 ( .A(n24684), .B(n24685), .Z(n27783) );
  XOR U37591 ( .A(n27782), .B(n27783), .Z(n27787) );
  XOR U37592 ( .A(n27785), .B(n27787), .Z(n27791) );
  XOR U37593 ( .A(n27789), .B(n27791), .Z(n27793) );
  XOR U37594 ( .A(n27792), .B(n27793), .Z(n24683) );
  XOR U37595 ( .A(n24681), .B(n24683), .Z(n27797) );
  XOR U37596 ( .A(n27795), .B(n27797), .Z(n27800) );
  XOR U37597 ( .A(n27798), .B(n27800), .Z(n27803) );
  XOR U37598 ( .A(n27802), .B(n27803), .Z(n27807) );
  XOR U37599 ( .A(n27805), .B(n27807), .Z(n24680) );
  XOR U37600 ( .A(n24678), .B(n24680), .Z(n27811) );
  XOR U37601 ( .A(n27809), .B(n27811), .Z(n27813) );
  XOR U37602 ( .A(n27812), .B(n27813), .Z(n27818) );
  XOR U37603 ( .A(n27816), .B(n27818), .Z(n27821) );
  XOR U37604 ( .A(n27819), .B(n27821), .Z(n27825) );
  XOR U37605 ( .A(n27823), .B(n27825), .Z(n27827) );
  XOR U37606 ( .A(n27826), .B(n27827), .Z(n24676) );
  XOR U37607 ( .A(n24674), .B(n24676), .Z(n24670) );
  XOR U37608 ( .A(n24668), .B(n24670), .Z(n24673) );
  XOR U37609 ( .A(n24671), .B(n24673), .Z(n24664) );
  XOR U37610 ( .A(n24662), .B(n24664), .Z(n24667) );
  XOR U37611 ( .A(n24665), .B(n24667), .Z(n24658) );
  XOR U37612 ( .A(n24656), .B(n24658), .Z(n24660) );
  XOR U37613 ( .A(n24659), .B(n24660), .Z(n24651) );
  XOR U37614 ( .A(n24650), .B(n24651), .Z(n24654) );
  XOR U37615 ( .A(n24653), .B(n24654), .Z(n24646) );
  XOR U37616 ( .A(n24644), .B(n24646), .Z(n24649) );
  XOR U37617 ( .A(n24647), .B(n24649), .Z(n27834) );
  XOR U37618 ( .A(n27833), .B(n27834), .Z(n27838) );
  XOR U37619 ( .A(n27836), .B(n27838), .Z(n24640) );
  XOR U37620 ( .A(n24638), .B(n24640), .Z(n24643) );
  XOR U37621 ( .A(n24641), .B(n24643), .Z(n24636) );
  XOR U37622 ( .A(n24635), .B(n24636), .Z(n27840) );
  XOR U37623 ( .A(n27839), .B(n27840), .Z(n27844) );
  XOR U37624 ( .A(n27842), .B(n27844), .Z(n24634) );
  XOR U37625 ( .A(n24632), .B(n24634), .Z(n24627) );
  XOR U37626 ( .A(n24626), .B(n24627), .Z(n24631) );
  XOR U37627 ( .A(n24629), .B(n24631), .Z(n24622) );
  XOR U37628 ( .A(n24620), .B(n24622), .Z(n24624) );
  XOR U37629 ( .A(n24623), .B(n24624), .Z(n24615) );
  XOR U37630 ( .A(n24614), .B(n24615), .Z(n24618) );
  XOR U37631 ( .A(n24617), .B(n24618), .Z(n27851) );
  XOR U37632 ( .A(n27849), .B(n27851), .Z(n27853) );
  XOR U37633 ( .A(n27852), .B(n27853), .Z(n24609) );
  XOR U37634 ( .A(n24608), .B(n24609), .Z(n24613) );
  XOR U37635 ( .A(n24611), .B(n24613), .Z(n24607) );
  XOR U37636 ( .A(n24605), .B(n24607), .Z(n27859) );
  XOR U37637 ( .A(n27857), .B(n27859), .Z(n27861) );
  XOR U37638 ( .A(n27860), .B(n27861), .Z(n27865) );
  XOR U37639 ( .A(n27864), .B(n27865), .Z(n27869) );
  XOR U37640 ( .A(n27867), .B(n27869), .Z(n24604) );
  XOR U37641 ( .A(n24602), .B(n24604), .Z(n27872) );
  XOR U37642 ( .A(n27871), .B(n27872), .Z(n27876) );
  XOR U37643 ( .A(n27874), .B(n27876), .Z(n27880) );
  XOR U37644 ( .A(n27878), .B(n27880), .Z(n27882) );
  XOR U37645 ( .A(n27881), .B(n27882), .Z(n27886) );
  XOR U37646 ( .A(n27885), .B(n27886), .Z(n27890) );
  XOR U37647 ( .A(n27888), .B(n27890), .Z(n24598) );
  XOR U37648 ( .A(n24596), .B(n24598), .Z(n24601) );
  XOR U37649 ( .A(n24599), .B(n24601), .Z(n27893) );
  XOR U37650 ( .A(n27892), .B(n27893), .Z(n27896) );
  XOR U37651 ( .A(n27895), .B(n27896), .Z(n24592) );
  XOR U37652 ( .A(n24590), .B(n24592), .Z(n24594) );
  XOR U37653 ( .A(n24593), .B(n24594), .Z(n27899) );
  XOR U37654 ( .A(n27898), .B(n27899), .Z(n27902) );
  XOR U37655 ( .A(n27901), .B(n27902), .Z(n24586) );
  XOR U37656 ( .A(n24584), .B(n24586), .Z(n24589) );
  XOR U37657 ( .A(n24587), .B(n24589), .Z(n27906) );
  XOR U37658 ( .A(n27905), .B(n27906), .Z(n27910) );
  XOR U37659 ( .A(n27908), .B(n27910), .Z(n27922) );
  XOR U37660 ( .A(n27920), .B(n27922), .Z(n27913) );
  XOR U37661 ( .A(n27912), .B(n27913), .Z(n27917) );
  XOR U37662 ( .A(n27916), .B(n27917), .Z(n24579) );
  XOR U37663 ( .A(n24578), .B(n24579), .Z(n24583) );
  XOR U37664 ( .A(n24581), .B(n24583), .Z(n24577) );
  XOR U37665 ( .A(n24575), .B(n24577), .Z(n27931) );
  XOR U37666 ( .A(n27929), .B(n27931), .Z(n27934) );
  XOR U37667 ( .A(n27932), .B(n27934), .Z(n27937) );
  XOR U37668 ( .A(n27936), .B(n27937), .Z(n27941) );
  XOR U37669 ( .A(n27939), .B(n27941), .Z(n24569) );
  XOR U37670 ( .A(n24568), .B(n24569), .Z(n24573) );
  XOR U37671 ( .A(n24571), .B(n24573), .Z(n24564) );
  XOR U37672 ( .A(n24562), .B(n24564), .Z(n24567) );
  XOR U37673 ( .A(n24565), .B(n24567), .Z(n24557) );
  XOR U37674 ( .A(n24556), .B(n24557), .Z(n24561) );
  XOR U37675 ( .A(n24559), .B(n24561), .Z(n24552) );
  XOR U37676 ( .A(n24550), .B(n24552), .Z(n24555) );
  XOR U37677 ( .A(n24553), .B(n24555), .Z(n27945) );
  XOR U37678 ( .A(n27944), .B(n27945), .Z(n27948) );
  XOR U37679 ( .A(n27947), .B(n27948), .Z(n27953) );
  XOR U37680 ( .A(n27951), .B(n27953), .Z(n27955) );
  XOR U37681 ( .A(n27954), .B(n27955), .Z(n27959) );
  XOR U37682 ( .A(n27958), .B(n27959), .Z(n27963) );
  XOR U37683 ( .A(n27961), .B(n27963), .Z(n27967) );
  XOR U37684 ( .A(n27965), .B(n27967), .Z(n27969) );
  XOR U37685 ( .A(n27968), .B(n27969), .Z(n27972) );
  XOR U37686 ( .A(n27971), .B(n27972), .Z(n27976) );
  XOR U37687 ( .A(n27974), .B(n27976), .Z(n27980) );
  XOR U37688 ( .A(n27978), .B(n27980), .Z(n27983) );
  XOR U37689 ( .A(n27981), .B(n27983), .Z(n24548) );
  XOR U37690 ( .A(n24547), .B(n24548), .Z(n27986) );
  XOR U37691 ( .A(n27985), .B(n27986), .Z(n27989) );
  XOR U37692 ( .A(n27988), .B(n27989), .Z(n24545) );
  XOR U37693 ( .A(n24544), .B(n24545), .Z(n27996) );
  XOR U37694 ( .A(n27995), .B(n27996), .Z(n24542) );
  XOR U37695 ( .A(n24541), .B(n24542), .Z(n28003) );
  XOR U37696 ( .A(n28001), .B(n28003), .Z(n28006) );
  XOR U37697 ( .A(n28004), .B(n28006), .Z(n28010) );
  XOR U37698 ( .A(n28008), .B(n28010), .Z(n28013) );
  XOR U37699 ( .A(n28011), .B(n28013), .Z(n28016) );
  XOR U37700 ( .A(n28014), .B(n28016), .Z(n28019) );
  XOR U37701 ( .A(n28017), .B(n28019), .Z(n24536) );
  XOR U37702 ( .A(n24535), .B(n24536), .Z(n24539) );
  XOR U37703 ( .A(n24538), .B(n24539), .Z(n24531) );
  XOR U37704 ( .A(n24529), .B(n24531), .Z(n24533) );
  XOR U37705 ( .A(n24532), .B(n24533), .Z(n24524) );
  XOR U37706 ( .A(n24523), .B(n24524), .Z(n24528) );
  XOR U37707 ( .A(n24526), .B(n24528), .Z(n28023) );
  XOR U37708 ( .A(n28021), .B(n28023), .Z(n28026) );
  XOR U37709 ( .A(n28024), .B(n28026), .Z(n24518) );
  XOR U37710 ( .A(n24517), .B(n24518), .Z(n24522) );
  XOR U37711 ( .A(n24520), .B(n24522), .Z(n24516) );
  XOR U37712 ( .A(n24514), .B(n24516), .Z(n28030) );
  XOR U37713 ( .A(n28029), .B(n28030), .Z(n28033) );
  XOR U37714 ( .A(n28032), .B(n28033), .Z(n24513) );
  XOR U37715 ( .A(n24511), .B(n24513), .Z(n24507) );
  XOR U37716 ( .A(n24505), .B(n24507), .Z(n24510) );
  XOR U37717 ( .A(n24508), .B(n24510), .Z(n28040) );
  XOR U37718 ( .A(n28039), .B(n28040), .Z(n24503) );
  XOR U37719 ( .A(n24502), .B(n24503), .Z(n28045) );
  XOR U37720 ( .A(n28044), .B(n28045), .Z(n28052) );
  XOR U37721 ( .A(n28053), .B(n28052), .Z(n28061) );
  XOR U37722 ( .A(n28062), .B(n28061), .Z(n37963) );
  XOR U37723 ( .A(n37962), .B(n37963), .Z(n28067) );
  XOR U37724 ( .A(n28066), .B(n28067), .Z(n28070) );
  XOR U37725 ( .A(n28069), .B(n28070), .Z(n31186) );
  XOR U37726 ( .A(n31185), .B(n31186), .Z(n34373) );
  XOR U37727 ( .A(n34372), .B(n34373), .Z(n34380) );
  XOR U37728 ( .A(n34379), .B(n34380), .Z(n34386) );
  XOR U37729 ( .A(n34385), .B(n34386), .Z(n37792) );
  XOR U37730 ( .A(n37791), .B(n37792), .Z(n37799) );
  XOR U37731 ( .A(n37798), .B(n37799), .Z(n37826) );
  XOR U37732 ( .A(n37824), .B(n37826), .Z(n37820) );
  XOR U37733 ( .A(n37819), .B(n37820), .Z(n37840) );
  XOR U37734 ( .A(n37839), .B(n37840), .Z(n37859) );
  XOR U37735 ( .A(n37858), .B(n37859), .Z(n37871) );
  XOR U37736 ( .A(n37870), .B(n37871), .Z(n37890) );
  XOR U37737 ( .A(n37889), .B(n37890), .Z(n37902) );
  XOR U37738 ( .A(n37901), .B(n37902), .Z(n37910) );
  XOR U37739 ( .A(n37909), .B(n37910), .Z(n37927) );
  XOR U37740 ( .A(n37926), .B(n37927), .Z(n37931) );
  XOR U37741 ( .A(n37930), .B(n37931), .Z(n37937) );
  XOR U37742 ( .A(n37936), .B(n37937), .Z(n44555) );
  XOR U37743 ( .A(n44554), .B(n44555), .Z(n44573) );
  XOR U37744 ( .A(n44572), .B(n44573), .Z(n44598) );
  XOR U37745 ( .A(n44597), .B(n44598), .Z(n44616) );
  XOR U37746 ( .A(n44615), .B(n44616), .Z(n44644) );
  XOR U37747 ( .A(n44643), .B(n44644), .Z(n44660) );
  XOR U37748 ( .A(n44659), .B(n44660), .Z(n44678) );
  XOR U37749 ( .A(n44677), .B(n44678), .Z(n48065) );
  XOR U37750 ( .A(n48064), .B(n48065), .Z(n48093) );
  XOR U37751 ( .A(n48092), .B(n48093), .Z(n54933) );
  XOR U37752 ( .A(n54932), .B(n54933), .Z(n54956) );
  XOR U37753 ( .A(n54955), .B(n54956), .Z(n54984) );
  XOR U37754 ( .A(n54983), .B(n54984), .Z(n55010) );
  XOR U37755 ( .A(n55009), .B(n55010), .Z(n55039) );
  XOR U37756 ( .A(n55038), .B(n55039), .Z(n55073) );
  XOR U37757 ( .A(n55074), .B(n55073), .Z(o[0]) );
  IV U37758 ( .A(n24502), .Z(n24504) );
  NOR U37759 ( .A(n24504), .B(n24503), .Z(n28048) );
  IV U37760 ( .A(n24505), .Z(n24506) );
  NOR U37761 ( .A(n24507), .B(n24506), .Z(n28087) );
  IV U37762 ( .A(n24508), .Z(n24509) );
  NOR U37763 ( .A(n24510), .B(n24509), .Z(n28082) );
  NOR U37764 ( .A(n28087), .B(n28082), .Z(n28037) );
  IV U37765 ( .A(n24511), .Z(n24512) );
  NOR U37766 ( .A(n24513), .B(n24512), .Z(n28085) );
  IV U37767 ( .A(n24514), .Z(n24515) );
  NOR U37768 ( .A(n24516), .B(n24515), .Z(n31164) );
  IV U37769 ( .A(n24517), .Z(n24519) );
  NOR U37770 ( .A(n24519), .B(n24518), .Z(n34342) );
  IV U37771 ( .A(n24520), .Z(n24521) );
  NOR U37772 ( .A(n24522), .B(n24521), .Z(n34348) );
  NOR U37773 ( .A(n34342), .B(n34348), .Z(n31163) );
  IV U37774 ( .A(n24523), .Z(n24525) );
  NOR U37775 ( .A(n24525), .B(n24524), .Z(n31211) );
  IV U37776 ( .A(n24526), .Z(n24527) );
  NOR U37777 ( .A(n24528), .B(n24527), .Z(n34335) );
  NOR U37778 ( .A(n31211), .B(n34335), .Z(n31157) );
  IV U37779 ( .A(n24529), .Z(n24530) );
  NOR U37780 ( .A(n24531), .B(n24530), .Z(n34317) );
  IV U37781 ( .A(n24532), .Z(n24534) );
  NOR U37782 ( .A(n24534), .B(n24533), .Z(n34327) );
  NOR U37783 ( .A(n34317), .B(n34327), .Z(n31151) );
  IV U37784 ( .A(n24535), .Z(n24537) );
  NOR U37785 ( .A(n24537), .B(n24536), .Z(n31147) );
  IV U37786 ( .A(n24538), .Z(n24540) );
  NOR U37787 ( .A(n24540), .B(n24539), .Z(n31152) );
  NOR U37788 ( .A(n31147), .B(n31152), .Z(n28020) );
  IV U37789 ( .A(n24541), .Z(n24543) );
  NOR U37790 ( .A(n24543), .B(n24542), .Z(n27999) );
  IV U37791 ( .A(n27999), .Z(n27994) );
  IV U37792 ( .A(n24544), .Z(n24546) );
  NOR U37793 ( .A(n24546), .B(n24545), .Z(n28093) );
  IV U37794 ( .A(n24547), .Z(n24549) );
  NOR U37795 ( .A(n24549), .B(n24548), .Z(n28098) );
  IV U37796 ( .A(n24550), .Z(n24551) );
  NOR U37797 ( .A(n24552), .B(n24551), .Z(n31247) );
  IV U37798 ( .A(n24553), .Z(n24554) );
  NOR U37799 ( .A(n24555), .B(n24554), .Z(n34248) );
  NOR U37800 ( .A(n31247), .B(n34248), .Z(n31103) );
  IV U37801 ( .A(n24556), .Z(n24558) );
  NOR U37802 ( .A(n24558), .B(n24557), .Z(n34464) );
  IV U37803 ( .A(n24559), .Z(n24560) );
  NOR U37804 ( .A(n24561), .B(n24560), .Z(n34457) );
  NOR U37805 ( .A(n34464), .B(n34457), .Z(n31101) );
  IV U37806 ( .A(n24562), .Z(n24563) );
  NOR U37807 ( .A(n24564), .B(n24563), .Z(n31086) );
  IV U37808 ( .A(n24565), .Z(n24566) );
  NOR U37809 ( .A(n24567), .B(n24566), .Z(n28117) );
  NOR U37810 ( .A(n31086), .B(n28117), .Z(n27943) );
  IV U37811 ( .A(n24568), .Z(n24570) );
  NOR U37812 ( .A(n24570), .B(n24569), .Z(n31261) );
  IV U37813 ( .A(n24571), .Z(n24572) );
  NOR U37814 ( .A(n24573), .B(n24572), .Z(n24574) );
  NOR U37815 ( .A(n31261), .B(n24574), .Z(n31091) );
  IV U37816 ( .A(n24575), .Z(n24576) );
  NOR U37817 ( .A(n24577), .B(n24576), .Z(n28127) );
  IV U37818 ( .A(n24578), .Z(n24580) );
  NOR U37819 ( .A(n24580), .B(n24579), .Z(n28136) );
  IV U37820 ( .A(n24581), .Z(n24582) );
  NOR U37821 ( .A(n24583), .B(n24582), .Z(n28132) );
  NOR U37822 ( .A(n28136), .B(n28132), .Z(n27928) );
  IV U37823 ( .A(n24584), .Z(n24585) );
  NOR U37824 ( .A(n24586), .B(n24585), .Z(n28141) );
  IV U37825 ( .A(n24587), .Z(n24588) );
  NOR U37826 ( .A(n24589), .B(n24588), .Z(n31055) );
  NOR U37827 ( .A(n28141), .B(n31055), .Z(n27904) );
  IV U37828 ( .A(n24590), .Z(n24591) );
  NOR U37829 ( .A(n24592), .B(n24591), .Z(n34209) );
  IV U37830 ( .A(n24593), .Z(n24595) );
  NOR U37831 ( .A(n24595), .B(n24594), .Z(n34204) );
  NOR U37832 ( .A(n34209), .B(n34204), .Z(n31049) );
  IV U37833 ( .A(n24596), .Z(n24597) );
  NOR U37834 ( .A(n24598), .B(n24597), .Z(n31292) );
  IV U37835 ( .A(n24599), .Z(n24600) );
  NOR U37836 ( .A(n24601), .B(n24600), .Z(n31288) );
  NOR U37837 ( .A(n31292), .B(n31288), .Z(n31043) );
  IV U37838 ( .A(n24602), .Z(n24603) );
  NOR U37839 ( .A(n24604), .B(n24603), .Z(n34504) );
  IV U37840 ( .A(n24605), .Z(n24606) );
  NOR U37841 ( .A(n24607), .B(n24606), .Z(n28154) );
  IV U37842 ( .A(n24608), .Z(n24610) );
  NOR U37843 ( .A(n24610), .B(n24609), .Z(n34180) );
  IV U37844 ( .A(n24611), .Z(n24612) );
  NOR U37845 ( .A(n24613), .B(n24612), .Z(n31314) );
  NOR U37846 ( .A(n34180), .B(n31314), .Z(n28153) );
  IV U37847 ( .A(n24614), .Z(n24616) );
  NOR U37848 ( .A(n24616), .B(n24615), .Z(n28164) );
  IV U37849 ( .A(n24617), .Z(n24619) );
  NOR U37850 ( .A(n24619), .B(n24618), .Z(n28166) );
  NOR U37851 ( .A(n28164), .B(n28166), .Z(n27848) );
  IV U37852 ( .A(n24620), .Z(n24621) );
  NOR U37853 ( .A(n24622), .B(n24621), .Z(n28175) );
  IV U37854 ( .A(n24623), .Z(n24625) );
  NOR U37855 ( .A(n24625), .B(n24624), .Z(n28173) );
  NOR U37856 ( .A(n28175), .B(n28173), .Z(n27847) );
  IV U37857 ( .A(n24626), .Z(n24628) );
  NOR U37858 ( .A(n24628), .B(n24627), .Z(n31005) );
  IV U37859 ( .A(n24629), .Z(n24630) );
  NOR U37860 ( .A(n24631), .B(n24630), .Z(n31010) );
  NOR U37861 ( .A(n31005), .B(n31010), .Z(n27846) );
  IV U37862 ( .A(n24632), .Z(n24633) );
  NOR U37863 ( .A(n24634), .B(n24633), .Z(n31004) );
  IV U37864 ( .A(n31004), .Z(n31001) );
  IV U37865 ( .A(n24635), .Z(n24637) );
  NOR U37866 ( .A(n24637), .B(n24636), .Z(n28181) );
  IV U37867 ( .A(n24638), .Z(n24639) );
  NOR U37868 ( .A(n24640), .B(n24639), .Z(n34158) );
  IV U37869 ( .A(n24641), .Z(n24642) );
  NOR U37870 ( .A(n24643), .B(n24642), .Z(n34153) );
  NOR U37871 ( .A(n34158), .B(n34153), .Z(n30996) );
  IV U37872 ( .A(n24644), .Z(n24645) );
  NOR U37873 ( .A(n24646), .B(n24645), .Z(n31335) );
  IV U37874 ( .A(n24647), .Z(n24648) );
  NOR U37875 ( .A(n24649), .B(n24648), .Z(n34141) );
  NOR U37876 ( .A(n31335), .B(n34141), .Z(n30978) );
  IV U37877 ( .A(n24650), .Z(n24652) );
  NOR U37878 ( .A(n24652), .B(n24651), .Z(n30953) );
  IV U37879 ( .A(n24653), .Z(n24655) );
  NOR U37880 ( .A(n24655), .B(n24654), .Z(n28183) );
  NOR U37881 ( .A(n30953), .B(n28183), .Z(n27832) );
  IV U37882 ( .A(n24656), .Z(n24657) );
  NOR U37883 ( .A(n24658), .B(n24657), .Z(n28187) );
  IV U37884 ( .A(n24659), .Z(n24661) );
  NOR U37885 ( .A(n24661), .B(n24660), .Z(n30958) );
  NOR U37886 ( .A(n28187), .B(n30958), .Z(n27830) );
  IV U37887 ( .A(n24662), .Z(n24663) );
  NOR U37888 ( .A(n24664), .B(n24663), .Z(n31348) );
  IV U37889 ( .A(n24665), .Z(n24666) );
  NOR U37890 ( .A(n24667), .B(n24666), .Z(n31341) );
  NOR U37891 ( .A(n31348), .B(n31341), .Z(n28186) );
  IV U37892 ( .A(n24668), .Z(n24669) );
  NOR U37893 ( .A(n24670), .B(n24669), .Z(n30938) );
  IV U37894 ( .A(n24671), .Z(n24672) );
  NOR U37895 ( .A(n24673), .B(n24672), .Z(n30949) );
  NOR U37896 ( .A(n30938), .B(n30949), .Z(n27829) );
  IV U37897 ( .A(n24674), .Z(n24675) );
  NOR U37898 ( .A(n24676), .B(n24675), .Z(n24677) );
  IV U37899 ( .A(n24677), .Z(n30943) );
  IV U37900 ( .A(n24678), .Z(n24679) );
  NOR U37901 ( .A(n24680), .B(n24679), .Z(n28196) );
  IV U37902 ( .A(n24681), .Z(n24682) );
  NOR U37903 ( .A(n24683), .B(n24682), .Z(n30919) );
  IV U37904 ( .A(n24684), .Z(n24686) );
  NOR U37905 ( .A(n24686), .B(n24685), .Z(n30900) );
  IV U37906 ( .A(n24687), .Z(n24688) );
  NOR U37907 ( .A(n24689), .B(n24688), .Z(n31379) );
  IV U37908 ( .A(n24690), .Z(n24691) );
  NOR U37909 ( .A(n24692), .B(n24691), .Z(n31375) );
  NOR U37910 ( .A(n31379), .B(n31375), .Z(n30881) );
  IV U37911 ( .A(n24693), .Z(n24695) );
  NOR U37912 ( .A(n24695), .B(n24694), .Z(n30882) );
  IV U37913 ( .A(n24696), .Z(n24697) );
  NOR U37914 ( .A(n24698), .B(n24697), .Z(n30884) );
  NOR U37915 ( .A(n30882), .B(n30884), .Z(n27781) );
  IV U37916 ( .A(n24699), .Z(n24700) );
  NOR U37917 ( .A(n24701), .B(n24700), .Z(n31384) );
  IV U37918 ( .A(n24702), .Z(n24703) );
  NOR U37919 ( .A(n24704), .B(n24703), .Z(n31389) );
  NOR U37920 ( .A(n31384), .B(n31389), .Z(n24705) );
  IV U37921 ( .A(n24705), .Z(n30876) );
  IV U37922 ( .A(n24706), .Z(n24708) );
  NOR U37923 ( .A(n24708), .B(n24707), .Z(n30875) );
  IV U37924 ( .A(n30875), .Z(n31398) );
  IV U37925 ( .A(n24709), .Z(n24710) );
  NOR U37926 ( .A(n24711), .B(n24710), .Z(n28206) );
  IV U37927 ( .A(n24712), .Z(n24714) );
  NOR U37928 ( .A(n24714), .B(n24713), .Z(n28204) );
  NOR U37929 ( .A(n28206), .B(n28204), .Z(n27780) );
  IV U37930 ( .A(n24715), .Z(n24716) );
  NOR U37931 ( .A(n24717), .B(n24716), .Z(n30868) );
  IV U37932 ( .A(n24718), .Z(n24719) );
  NOR U37933 ( .A(n24720), .B(n24719), .Z(n30865) );
  NOR U37934 ( .A(n30868), .B(n30865), .Z(n27778) );
  IV U37935 ( .A(n24721), .Z(n24722) );
  NOR U37936 ( .A(n24723), .B(n24722), .Z(n27768) );
  IV U37937 ( .A(n24724), .Z(n24725) );
  NOR U37938 ( .A(n24726), .B(n24725), .Z(n30819) );
  IV U37939 ( .A(n24727), .Z(n24729) );
  NOR U37940 ( .A(n24729), .B(n24728), .Z(n30837) );
  NOR U37941 ( .A(n30819), .B(n30837), .Z(n27759) );
  IV U37942 ( .A(n24730), .Z(n24732) );
  NOR U37943 ( .A(n24732), .B(n24731), .Z(n30822) );
  IV U37944 ( .A(n24733), .Z(n24734) );
  NOR U37945 ( .A(n24735), .B(n24734), .Z(n30829) );
  NOR U37946 ( .A(n30822), .B(n30829), .Z(n27758) );
  IV U37947 ( .A(n24736), .Z(n24737) );
  NOR U37948 ( .A(n24738), .B(n24737), .Z(n30807) );
  IV U37949 ( .A(n24739), .Z(n24740) );
  NOR U37950 ( .A(n24741), .B(n24740), .Z(n30814) );
  NOR U37951 ( .A(n30807), .B(n30814), .Z(n27757) );
  IV U37952 ( .A(n24742), .Z(n24744) );
  NOR U37953 ( .A(n24744), .B(n24743), .Z(n30803) );
  IV U37954 ( .A(n24745), .Z(n24747) );
  NOR U37955 ( .A(n24747), .B(n24746), .Z(n30809) );
  NOR U37956 ( .A(n30803), .B(n30809), .Z(n27756) );
  IV U37957 ( .A(n24748), .Z(n24749) );
  NOR U37958 ( .A(n24750), .B(n24749), .Z(n28211) );
  IV U37959 ( .A(n24751), .Z(n24753) );
  NOR U37960 ( .A(n24753), .B(n24752), .Z(n28220) );
  IV U37961 ( .A(n24754), .Z(n24756) );
  NOR U37962 ( .A(n24756), .B(n24755), .Z(n30798) );
  IV U37963 ( .A(n24757), .Z(n24758) );
  NOR U37964 ( .A(n24759), .B(n24758), .Z(n28223) );
  NOR U37965 ( .A(n30798), .B(n28223), .Z(n27731) );
  IV U37966 ( .A(n24760), .Z(n24762) );
  NOR U37967 ( .A(n24762), .B(n24761), .Z(n31425) );
  IV U37968 ( .A(n24763), .Z(n24764) );
  NOR U37969 ( .A(n24765), .B(n24764), .Z(n24766) );
  NOR U37970 ( .A(n31425), .B(n24766), .Z(n30790) );
  IV U37971 ( .A(n24767), .Z(n24769) );
  NOR U37972 ( .A(n24769), .B(n24768), .Z(n28227) );
  IV U37973 ( .A(n24770), .Z(n24772) );
  NOR U37974 ( .A(n24772), .B(n24771), .Z(n30767) );
  IV U37975 ( .A(n24773), .Z(n24774) );
  NOR U37976 ( .A(n24775), .B(n24774), .Z(n30785) );
  NOR U37977 ( .A(n30767), .B(n30785), .Z(n27723) );
  IV U37978 ( .A(n24776), .Z(n24777) );
  NOR U37979 ( .A(n24778), .B(n24777), .Z(n30770) );
  IV U37980 ( .A(n24779), .Z(n24781) );
  NOR U37981 ( .A(n24781), .B(n24780), .Z(n30777) );
  NOR U37982 ( .A(n30770), .B(n30777), .Z(n27722) );
  IV U37983 ( .A(n24782), .Z(n24783) );
  NOR U37984 ( .A(n24784), .B(n24783), .Z(n28234) );
  IV U37985 ( .A(n24785), .Z(n24786) );
  NOR U37986 ( .A(n24787), .B(n24786), .Z(n28231) );
  NOR U37987 ( .A(n28234), .B(n28231), .Z(n27721) );
  IV U37988 ( .A(n24788), .Z(n24789) );
  NOR U37989 ( .A(n24790), .B(n24789), .Z(n28240) );
  IV U37990 ( .A(n24791), .Z(n24793) );
  NOR U37991 ( .A(n24793), .B(n24792), .Z(n28237) );
  NOR U37992 ( .A(n28240), .B(n28237), .Z(n27720) );
  IV U37993 ( .A(n24794), .Z(n24795) );
  NOR U37994 ( .A(n24796), .B(n24795), .Z(n24797) );
  IV U37995 ( .A(n24797), .Z(n28245) );
  IV U37996 ( .A(n24798), .Z(n24800) );
  NOR U37997 ( .A(n24800), .B(n24799), .Z(n31442) );
  IV U37998 ( .A(n24801), .Z(n24803) );
  NOR U37999 ( .A(n24803), .B(n24802), .Z(n31437) );
  NOR U38000 ( .A(n31442), .B(n31437), .Z(n28243) );
  IV U38001 ( .A(n24804), .Z(n24805) );
  NOR U38002 ( .A(n24806), .B(n24805), .Z(n30761) );
  IV U38003 ( .A(n24807), .Z(n24808) );
  NOR U38004 ( .A(n24809), .B(n24808), .Z(n28247) );
  NOR U38005 ( .A(n30761), .B(n28247), .Z(n27719) );
  IV U38006 ( .A(n24810), .Z(n24812) );
  NOR U38007 ( .A(n24812), .B(n24811), .Z(n28252) );
  IV U38008 ( .A(n24813), .Z(n24814) );
  NOR U38009 ( .A(n24815), .B(n24814), .Z(n28250) );
  NOR U38010 ( .A(n28252), .B(n28250), .Z(n27718) );
  IV U38011 ( .A(n24816), .Z(n24817) );
  NOR U38012 ( .A(n24818), .B(n24817), .Z(n28255) );
  IV U38013 ( .A(n24819), .Z(n24820) );
  NOR U38014 ( .A(n24821), .B(n24820), .Z(n30747) );
  NOR U38015 ( .A(n28255), .B(n30747), .Z(n27717) );
  IV U38016 ( .A(n24822), .Z(n24824) );
  NOR U38017 ( .A(n24824), .B(n24823), .Z(n27715) );
  IV U38018 ( .A(n27715), .Z(n27710) );
  IV U38019 ( .A(n24825), .Z(n24826) );
  NOR U38020 ( .A(n24827), .B(n24826), .Z(n30731) );
  IV U38021 ( .A(n24828), .Z(n24829) );
  NOR U38022 ( .A(n24830), .B(n24829), .Z(n31463) );
  IV U38023 ( .A(n24831), .Z(n24832) );
  NOR U38024 ( .A(n24833), .B(n24832), .Z(n31456) );
  NOR U38025 ( .A(n31463), .B(n31456), .Z(n30730) );
  IV U38026 ( .A(n24834), .Z(n24835) );
  NOR U38027 ( .A(n24836), .B(n24835), .Z(n28264) );
  IV U38028 ( .A(n24837), .Z(n24839) );
  NOR U38029 ( .A(n24839), .B(n24838), .Z(n28261) );
  NOR U38030 ( .A(n28264), .B(n28261), .Z(n27708) );
  IV U38031 ( .A(n24840), .Z(n24842) );
  NOR U38032 ( .A(n24842), .B(n24841), .Z(n28266) );
  IV U38033 ( .A(n24843), .Z(n24844) );
  NOR U38034 ( .A(n24845), .B(n24844), .Z(n31495) );
  IV U38035 ( .A(n24846), .Z(n24847) );
  NOR U38036 ( .A(n24848), .B(n24847), .Z(n31490) );
  NOR U38037 ( .A(n31495), .B(n31490), .Z(n28272) );
  IV U38038 ( .A(n24849), .Z(n24850) );
  NOR U38039 ( .A(n24851), .B(n24850), .Z(n31501) );
  IV U38040 ( .A(n24852), .Z(n24853) );
  NOR U38041 ( .A(n24854), .B(n24853), .Z(n34014) );
  NOR U38042 ( .A(n31501), .B(n34014), .Z(n30716) );
  IV U38043 ( .A(n24855), .Z(n24857) );
  NOR U38044 ( .A(n24857), .B(n24856), .Z(n31516) );
  IV U38045 ( .A(n24858), .Z(n24859) );
  NOR U38046 ( .A(n24860), .B(n24859), .Z(n31505) );
  NOR U38047 ( .A(n31516), .B(n31505), .Z(n30714) );
  IV U38048 ( .A(n24861), .Z(n24862) );
  NOR U38049 ( .A(n24863), .B(n24862), .Z(n31519) );
  IV U38050 ( .A(n24864), .Z(n24865) );
  NOR U38051 ( .A(n24866), .B(n24865), .Z(n31511) );
  NOR U38052 ( .A(n31519), .B(n31511), .Z(n24867) );
  IV U38053 ( .A(n24867), .Z(n30710) );
  IV U38054 ( .A(n24868), .Z(n24870) );
  NOR U38055 ( .A(n24870), .B(n24869), .Z(n34004) );
  IV U38056 ( .A(n24871), .Z(n24873) );
  NOR U38057 ( .A(n24873), .B(n24872), .Z(n31522) );
  NOR U38058 ( .A(n34004), .B(n31522), .Z(n24874) );
  IV U38059 ( .A(n24874), .Z(n30708) );
  IV U38060 ( .A(n24875), .Z(n24876) );
  NOR U38061 ( .A(n24877), .B(n24876), .Z(n30698) );
  IV U38062 ( .A(n24878), .Z(n24879) );
  NOR U38063 ( .A(n24880), .B(n24879), .Z(n28279) );
  NOR U38064 ( .A(n30698), .B(n28279), .Z(n27680) );
  IV U38065 ( .A(n24881), .Z(n24882) );
  NOR U38066 ( .A(n24883), .B(n24882), .Z(n31532) );
  IV U38067 ( .A(n24884), .Z(n24885) );
  NOR U38068 ( .A(n24886), .B(n24885), .Z(n31527) );
  NOR U38069 ( .A(n31532), .B(n31527), .Z(n30702) );
  IV U38070 ( .A(n24887), .Z(n24888) );
  NOR U38071 ( .A(n24889), .B(n24888), .Z(n31540) );
  IV U38072 ( .A(n24890), .Z(n24891) );
  NOR U38073 ( .A(n24892), .B(n24891), .Z(n31535) );
  NOR U38074 ( .A(n31540), .B(n31535), .Z(n30692) );
  IV U38075 ( .A(n24893), .Z(n24895) );
  NOR U38076 ( .A(n24895), .B(n24894), .Z(n28285) );
  IV U38077 ( .A(n24896), .Z(n24897) );
  NOR U38078 ( .A(n24898), .B(n24897), .Z(n31562) );
  IV U38079 ( .A(n24899), .Z(n24900) );
  NOR U38080 ( .A(n24901), .B(n24900), .Z(n31550) );
  NOR U38081 ( .A(n31562), .B(n31550), .Z(n28295) );
  IV U38082 ( .A(n24902), .Z(n24904) );
  NOR U38083 ( .A(n24904), .B(n24903), .Z(n33992) );
  IV U38084 ( .A(n24905), .Z(n24907) );
  NOR U38085 ( .A(n24907), .B(n24906), .Z(n34755) );
  IV U38086 ( .A(n24908), .Z(n24909) );
  NOR U38087 ( .A(n24910), .B(n24909), .Z(n37371) );
  NOR U38088 ( .A(n34755), .B(n37371), .Z(n28316) );
  IV U38089 ( .A(n24911), .Z(n24913) );
  NOR U38090 ( .A(n24913), .B(n24912), .Z(n28317) );
  IV U38091 ( .A(n24914), .Z(n24915) );
  NOR U38092 ( .A(n24916), .B(n24915), .Z(n28314) );
  NOR U38093 ( .A(n28317), .B(n28314), .Z(n27651) );
  IV U38094 ( .A(n24917), .Z(n24919) );
  NOR U38095 ( .A(n24919), .B(n24918), .Z(n28324) );
  IV U38096 ( .A(n24920), .Z(n24921) );
  NOR U38097 ( .A(n24922), .B(n24921), .Z(n28320) );
  NOR U38098 ( .A(n28324), .B(n28320), .Z(n27650) );
  IV U38099 ( .A(n24923), .Z(n24924) );
  NOR U38100 ( .A(n24925), .B(n24924), .Z(n33971) );
  IV U38101 ( .A(n24926), .Z(n24928) );
  NOR U38102 ( .A(n24928), .B(n24927), .Z(n31573) );
  NOR U38103 ( .A(n33971), .B(n31573), .Z(n28323) );
  IV U38104 ( .A(n24929), .Z(n24931) );
  NOR U38105 ( .A(n24931), .B(n24930), .Z(n30659) );
  IV U38106 ( .A(n24932), .Z(n24933) );
  NOR U38107 ( .A(n24934), .B(n24933), .Z(n28331) );
  NOR U38108 ( .A(n30659), .B(n28331), .Z(n27635) );
  IV U38109 ( .A(n24935), .Z(n24936) );
  NOR U38110 ( .A(n24937), .B(n24936), .Z(n30651) );
  IV U38111 ( .A(n24938), .Z(n24939) );
  NOR U38112 ( .A(n24940), .B(n24939), .Z(n28334) );
  NOR U38113 ( .A(n30651), .B(n28334), .Z(n27634) );
  IV U38114 ( .A(n24941), .Z(n24943) );
  NOR U38115 ( .A(n24943), .B(n24942), .Z(n28339) );
  IV U38116 ( .A(n24944), .Z(n24946) );
  NOR U38117 ( .A(n24946), .B(n24945), .Z(n28336) );
  NOR U38118 ( .A(n28339), .B(n28336), .Z(n27633) );
  IV U38119 ( .A(n24947), .Z(n24948) );
  NOR U38120 ( .A(n24949), .B(n24948), .Z(n24950) );
  IV U38121 ( .A(n24950), .Z(n28343) );
  IV U38122 ( .A(n24951), .Z(n24952) );
  NOR U38123 ( .A(n24953), .B(n24952), .Z(n27629) );
  IV U38124 ( .A(n24954), .Z(n24955) );
  NOR U38125 ( .A(n24956), .B(n24955), .Z(n33929) );
  IV U38126 ( .A(n24957), .Z(n24958) );
  NOR U38127 ( .A(n24959), .B(n24958), .Z(n33935) );
  NOR U38128 ( .A(n33929), .B(n33935), .Z(n28350) );
  IV U38129 ( .A(n24960), .Z(n24962) );
  NOR U38130 ( .A(n24962), .B(n24961), .Z(n30640) );
  IV U38131 ( .A(n24963), .Z(n24964) );
  NOR U38132 ( .A(n24965), .B(n24964), .Z(n30645) );
  NOR U38133 ( .A(n30640), .B(n30645), .Z(n27620) );
  IV U38134 ( .A(n24966), .Z(n24967) );
  NOR U38135 ( .A(n24968), .B(n24967), .Z(n30638) );
  IV U38136 ( .A(n24969), .Z(n24970) );
  NOR U38137 ( .A(n24971), .B(n24970), .Z(n33906) );
  IV U38138 ( .A(n24972), .Z(n24974) );
  NOR U38139 ( .A(n24974), .B(n24973), .Z(n33911) );
  NOR U38140 ( .A(n33906), .B(n33911), .Z(n28357) );
  IV U38141 ( .A(n24975), .Z(n24976) );
  NOR U38142 ( .A(n24977), .B(n24976), .Z(n30631) );
  IV U38143 ( .A(n24978), .Z(n24980) );
  NOR U38144 ( .A(n24980), .B(n24979), .Z(n28364) );
  NOR U38145 ( .A(n30631), .B(n28364), .Z(n27605) );
  IV U38146 ( .A(n24981), .Z(n24982) );
  NOR U38147 ( .A(n24983), .B(n24982), .Z(n33901) );
  IV U38148 ( .A(n24984), .Z(n24986) );
  NOR U38149 ( .A(n24986), .B(n24985), .Z(n31603) );
  NOR U38150 ( .A(n33901), .B(n31603), .Z(n28368) );
  IV U38151 ( .A(n24987), .Z(n24989) );
  NOR U38152 ( .A(n24989), .B(n24988), .Z(n34826) );
  IV U38153 ( .A(n24990), .Z(n24991) );
  NOR U38154 ( .A(n24992), .B(n24991), .Z(n34819) );
  NOR U38155 ( .A(n34826), .B(n34819), .Z(n28367) );
  IV U38156 ( .A(n24993), .Z(n24994) );
  NOR U38157 ( .A(n24995), .B(n24994), .Z(n37296) );
  IV U38158 ( .A(n24996), .Z(n24998) );
  NOR U38159 ( .A(n24998), .B(n24997), .Z(n37302) );
  NOR U38160 ( .A(n37296), .B(n37302), .Z(n28370) );
  IV U38161 ( .A(n24999), .Z(n25001) );
  NOR U38162 ( .A(n25001), .B(n25000), .Z(n41635) );
  IV U38163 ( .A(n25002), .Z(n25003) );
  NOR U38164 ( .A(n25004), .B(n25003), .Z(n41625) );
  NOR U38165 ( .A(n41635), .B(n41625), .Z(n30626) );
  IV U38166 ( .A(n25005), .Z(n25006) );
  NOR U38167 ( .A(n25007), .B(n25006), .Z(n25008) );
  IV U38168 ( .A(n25008), .Z(n27594) );
  IV U38169 ( .A(n25009), .Z(n25010) );
  NOR U38170 ( .A(n25011), .B(n25010), .Z(n30606) );
  IV U38171 ( .A(n25012), .Z(n25013) );
  NOR U38172 ( .A(n25014), .B(n25013), .Z(n34840) );
  IV U38173 ( .A(n25015), .Z(n25017) );
  NOR U38174 ( .A(n25017), .B(n25016), .Z(n37284) );
  NOR U38175 ( .A(n34840), .B(n37284), .Z(n33882) );
  IV U38176 ( .A(n25018), .Z(n25020) );
  NOR U38177 ( .A(n25020), .B(n25019), .Z(n28371) );
  IV U38178 ( .A(n25021), .Z(n25022) );
  NOR U38179 ( .A(n25023), .B(n25022), .Z(n30602) );
  NOR U38180 ( .A(n28371), .B(n30602), .Z(n27584) );
  IV U38181 ( .A(n25024), .Z(n25026) );
  NOR U38182 ( .A(n25026), .B(n25025), .Z(n28373) );
  IV U38183 ( .A(n25027), .Z(n25028) );
  NOR U38184 ( .A(n25029), .B(n25028), .Z(n37282) );
  IV U38185 ( .A(n25030), .Z(n25032) );
  NOR U38186 ( .A(n25032), .B(n25031), .Z(n25033) );
  NOR U38187 ( .A(n37282), .B(n25033), .Z(n28377) );
  IV U38188 ( .A(n25034), .Z(n25036) );
  NOR U38189 ( .A(n25036), .B(n25035), .Z(n30585) );
  IV U38190 ( .A(n25037), .Z(n25038) );
  NOR U38191 ( .A(n25039), .B(n25038), .Z(n30583) );
  NOR U38192 ( .A(n30585), .B(n30583), .Z(n27583) );
  IV U38193 ( .A(n25040), .Z(n25042) );
  NOR U38194 ( .A(n25042), .B(n25041), .Z(n27565) );
  IV U38195 ( .A(n27565), .Z(n27555) );
  IV U38196 ( .A(n25043), .Z(n25044) );
  NOR U38197 ( .A(n25045), .B(n25044), .Z(n27552) );
  IV U38198 ( .A(n27552), .Z(n27545) );
  IV U38199 ( .A(n25046), .Z(n25047) );
  NOR U38200 ( .A(n25048), .B(n25047), .Z(n27550) );
  IV U38201 ( .A(n27550), .Z(n28385) );
  IV U38202 ( .A(n25049), .Z(n25051) );
  NOR U38203 ( .A(n25051), .B(n25050), .Z(n28396) );
  IV U38204 ( .A(n25052), .Z(n25053) );
  NOR U38205 ( .A(n25054), .B(n25053), .Z(n28404) );
  IV U38206 ( .A(n25055), .Z(n25056) );
  NOR U38207 ( .A(n25057), .B(n25056), .Z(n28399) );
  NOR U38208 ( .A(n28404), .B(n28399), .Z(n31640) );
  IV U38209 ( .A(n25058), .Z(n25059) );
  NOR U38210 ( .A(n25060), .B(n25059), .Z(n31648) );
  IV U38211 ( .A(n25061), .Z(n25062) );
  NOR U38212 ( .A(n25063), .B(n25062), .Z(n31643) );
  NOR U38213 ( .A(n31648), .B(n31643), .Z(n28403) );
  IV U38214 ( .A(n25064), .Z(n25065) );
  NOR U38215 ( .A(n25066), .B(n25065), .Z(n30569) );
  IV U38216 ( .A(n25067), .Z(n25068) );
  NOR U38217 ( .A(n25069), .B(n25068), .Z(n30575) );
  NOR U38218 ( .A(n30569), .B(n30575), .Z(n27528) );
  IV U38219 ( .A(n25070), .Z(n25072) );
  NOR U38220 ( .A(n25072), .B(n25071), .Z(n30563) );
  IV U38221 ( .A(n25073), .Z(n25075) );
  NOR U38222 ( .A(n25075), .B(n25074), .Z(n30571) );
  NOR U38223 ( .A(n30563), .B(n30571), .Z(n27527) );
  IV U38224 ( .A(n25076), .Z(n25078) );
  NOR U38225 ( .A(n25078), .B(n25077), .Z(n30558) );
  IV U38226 ( .A(n25079), .Z(n25081) );
  NOR U38227 ( .A(n25081), .B(n25080), .Z(n30565) );
  NOR U38228 ( .A(n30558), .B(n30565), .Z(n27526) );
  IV U38229 ( .A(n25082), .Z(n25083) );
  NOR U38230 ( .A(n25084), .B(n25083), .Z(n30556) );
  IV U38231 ( .A(n25085), .Z(n25086) );
  NOR U38232 ( .A(n25087), .B(n25086), .Z(n28411) );
  IV U38233 ( .A(n25088), .Z(n25090) );
  NOR U38234 ( .A(n25090), .B(n25089), .Z(n30545) );
  IV U38235 ( .A(n25091), .Z(n25093) );
  NOR U38236 ( .A(n25093), .B(n25092), .Z(n30552) );
  NOR U38237 ( .A(n30545), .B(n30552), .Z(n27517) );
  IV U38238 ( .A(n25094), .Z(n25095) );
  NOR U38239 ( .A(n25096), .B(n25095), .Z(n30537) );
  IV U38240 ( .A(n25097), .Z(n25099) );
  NOR U38241 ( .A(n25099), .B(n25098), .Z(n30520) );
  IV U38242 ( .A(n25100), .Z(n25102) );
  NOR U38243 ( .A(n25102), .B(n25101), .Z(n30530) );
  NOR U38244 ( .A(n30520), .B(n30530), .Z(n27508) );
  IV U38245 ( .A(n25103), .Z(n25104) );
  NOR U38246 ( .A(n25105), .B(n25104), .Z(n30522) );
  IV U38247 ( .A(n25106), .Z(n25108) );
  NOR U38248 ( .A(n25108), .B(n25107), .Z(n28417) );
  IV U38249 ( .A(n25109), .Z(n25110) );
  NOR U38250 ( .A(n25111), .B(n25110), .Z(n30525) );
  NOR U38251 ( .A(n28417), .B(n30525), .Z(n27507) );
  IV U38252 ( .A(n25112), .Z(n25114) );
  NOR U38253 ( .A(n25114), .B(n25113), .Z(n30512) );
  IV U38254 ( .A(n25115), .Z(n25116) );
  NOR U38255 ( .A(n25117), .B(n25116), .Z(n28419) );
  NOR U38256 ( .A(n30512), .B(n28419), .Z(n27506) );
  IV U38257 ( .A(n25118), .Z(n25119) );
  NOR U38258 ( .A(n25120), .B(n25119), .Z(n30491) );
  IV U38259 ( .A(n25121), .Z(n25122) );
  NOR U38260 ( .A(n25123), .B(n25122), .Z(n30509) );
  NOR U38261 ( .A(n30491), .B(n30509), .Z(n27505) );
  IV U38262 ( .A(n25124), .Z(n25126) );
  NOR U38263 ( .A(n25126), .B(n25125), .Z(n30493) );
  IV U38264 ( .A(n25127), .Z(n25129) );
  NOR U38265 ( .A(n25129), .B(n25128), .Z(n30488) );
  NOR U38266 ( .A(n30493), .B(n30488), .Z(n27504) );
  IV U38267 ( .A(n25130), .Z(n25131) );
  NOR U38268 ( .A(n25132), .B(n25131), .Z(n27490) );
  IV U38269 ( .A(n25133), .Z(n25134) );
  NOR U38270 ( .A(n25135), .B(n25134), .Z(n25136) );
  IV U38271 ( .A(n25136), .Z(n28425) );
  IV U38272 ( .A(n25137), .Z(n25139) );
  NOR U38273 ( .A(n25139), .B(n25138), .Z(n33777) );
  IV U38274 ( .A(n25140), .Z(n25141) );
  NOR U38275 ( .A(n25142), .B(n25141), .Z(n33781) );
  NOR U38276 ( .A(n33777), .B(n33781), .Z(n30482) );
  IV U38277 ( .A(n25143), .Z(n25144) );
  NOR U38278 ( .A(n25145), .B(n25144), .Z(n33767) );
  IV U38279 ( .A(n25146), .Z(n25147) );
  NOR U38280 ( .A(n25148), .B(n25147), .Z(n31681) );
  NOR U38281 ( .A(n33767), .B(n31681), .Z(n30477) );
  IV U38282 ( .A(n25149), .Z(n25151) );
  NOR U38283 ( .A(n25151), .B(n25150), .Z(n31685) );
  IV U38284 ( .A(n25152), .Z(n25153) );
  NOR U38285 ( .A(n25154), .B(n25153), .Z(n33764) );
  NOR U38286 ( .A(n31685), .B(n33764), .Z(n30475) );
  IV U38287 ( .A(n25155), .Z(n25156) );
  NOR U38288 ( .A(n25157), .B(n25156), .Z(n28426) );
  IV U38289 ( .A(n25158), .Z(n25159) );
  NOR U38290 ( .A(n25160), .B(n25159), .Z(n30471) );
  NOR U38291 ( .A(n28426), .B(n30471), .Z(n27474) );
  IV U38292 ( .A(n25161), .Z(n25162) );
  NOR U38293 ( .A(n25163), .B(n25162), .Z(n37185) );
  IV U38294 ( .A(n25164), .Z(n25165) );
  NOR U38295 ( .A(n25166), .B(n25165), .Z(n34980) );
  NOR U38296 ( .A(n37185), .B(n34980), .Z(n30452) );
  IV U38297 ( .A(n25167), .Z(n25168) );
  NOR U38298 ( .A(n25169), .B(n25168), .Z(n31708) );
  IV U38299 ( .A(n25170), .Z(n25171) );
  NOR U38300 ( .A(n25172), .B(n25171), .Z(n31703) );
  NOR U38301 ( .A(n31708), .B(n31703), .Z(n28432) );
  IV U38302 ( .A(n25173), .Z(n25175) );
  NOR U38303 ( .A(n25175), .B(n25174), .Z(n30425) );
  IV U38304 ( .A(n25176), .Z(n25177) );
  NOR U38305 ( .A(n25178), .B(n25177), .Z(n30419) );
  NOR U38306 ( .A(n30425), .B(n30419), .Z(n28433) );
  IV U38307 ( .A(n25179), .Z(n25180) );
  NOR U38308 ( .A(n25181), .B(n25180), .Z(n30411) );
  IV U38309 ( .A(n25182), .Z(n25183) );
  NOR U38310 ( .A(n25184), .B(n25183), .Z(n30406) );
  NOR U38311 ( .A(n30411), .B(n30406), .Z(n27447) );
  IV U38312 ( .A(n25185), .Z(n25186) );
  NOR U38313 ( .A(n25187), .B(n25186), .Z(n27445) );
  IV U38314 ( .A(n27445), .Z(n27440) );
  IV U38315 ( .A(n25188), .Z(n25190) );
  NOR U38316 ( .A(n25190), .B(n25189), .Z(n28434) );
  IV U38317 ( .A(n25191), .Z(n25192) );
  NOR U38318 ( .A(n25193), .B(n25192), .Z(n28440) );
  IV U38319 ( .A(n25194), .Z(n25195) );
  NOR U38320 ( .A(n25196), .B(n25195), .Z(n28445) );
  NOR U38321 ( .A(n28440), .B(n28445), .Z(n27438) );
  IV U38322 ( .A(n25197), .Z(n25198) );
  NOR U38323 ( .A(n25199), .B(n25198), .Z(n30400) );
  IV U38324 ( .A(n25200), .Z(n25202) );
  NOR U38325 ( .A(n25202), .B(n25201), .Z(n28442) );
  NOR U38326 ( .A(n30400), .B(n28442), .Z(n27437) );
  IV U38327 ( .A(n25203), .Z(n25204) );
  NOR U38328 ( .A(n25205), .B(n25204), .Z(n30394) );
  IV U38329 ( .A(n25206), .Z(n25208) );
  NOR U38330 ( .A(n25208), .B(n25207), .Z(n28449) );
  IV U38331 ( .A(n25209), .Z(n25211) );
  NOR U38332 ( .A(n25211), .B(n25210), .Z(n30396) );
  NOR U38333 ( .A(n28449), .B(n30396), .Z(n27436) );
  IV U38334 ( .A(n25212), .Z(n25213) );
  NOR U38335 ( .A(n25214), .B(n25213), .Z(n30382) );
  IV U38336 ( .A(n25215), .Z(n25216) );
  NOR U38337 ( .A(n25217), .B(n25216), .Z(n30376) );
  NOR U38338 ( .A(n30382), .B(n30376), .Z(n27435) );
  IV U38339 ( .A(n25218), .Z(n25220) );
  NOR U38340 ( .A(n25220), .B(n25219), .Z(n30380) );
  IV U38341 ( .A(n25221), .Z(n25222) );
  NOR U38342 ( .A(n25223), .B(n25222), .Z(n30370) );
  IV U38343 ( .A(n25224), .Z(n25226) );
  NOR U38344 ( .A(n25226), .B(n25225), .Z(n35026) );
  IV U38345 ( .A(n25227), .Z(n25228) );
  NOR U38346 ( .A(n25229), .B(n25228), .Z(n37123) );
  NOR U38347 ( .A(n35026), .B(n37123), .Z(n30369) );
  IV U38348 ( .A(n25230), .Z(n25232) );
  NOR U38349 ( .A(n25232), .B(n25231), .Z(n27421) );
  IV U38350 ( .A(n27421), .Z(n27414) );
  IV U38351 ( .A(n25233), .Z(n25234) );
  NOR U38352 ( .A(n25235), .B(n25234), .Z(n25236) );
  IV U38353 ( .A(n25236), .Z(n30361) );
  IV U38354 ( .A(n25237), .Z(n25238) );
  NOR U38355 ( .A(n25239), .B(n25238), .Z(n28457) );
  IV U38356 ( .A(n25240), .Z(n25241) );
  NOR U38357 ( .A(n25242), .B(n25241), .Z(n37106) );
  IV U38358 ( .A(n25243), .Z(n25244) );
  NOR U38359 ( .A(n25245), .B(n25244), .Z(n37115) );
  NOR U38360 ( .A(n37106), .B(n37115), .Z(n28462) );
  IV U38361 ( .A(n25246), .Z(n25247) );
  NOR U38362 ( .A(n25248), .B(n25247), .Z(n27370) );
  IV U38363 ( .A(n27370), .Z(n27361) );
  IV U38364 ( .A(n25249), .Z(n25251) );
  NOR U38365 ( .A(n25251), .B(n25250), .Z(n31742) );
  IV U38366 ( .A(n25252), .Z(n25254) );
  NOR U38367 ( .A(n25254), .B(n25253), .Z(n31738) );
  NOR U38368 ( .A(n31742), .B(n31738), .Z(n30309) );
  IV U38369 ( .A(n25255), .Z(n25257) );
  NOR U38370 ( .A(n25257), .B(n25256), .Z(n33675) );
  IV U38371 ( .A(n25258), .Z(n25259) );
  NOR U38372 ( .A(n25260), .B(n25259), .Z(n31747) );
  NOR U38373 ( .A(n33675), .B(n31747), .Z(n30303) );
  IV U38374 ( .A(n25261), .Z(n25263) );
  NOR U38375 ( .A(n25263), .B(n25262), .Z(n30292) );
  IV U38376 ( .A(n25264), .Z(n25266) );
  NOR U38377 ( .A(n25266), .B(n25265), .Z(n30286) );
  NOR U38378 ( .A(n30292), .B(n30286), .Z(n28486) );
  IV U38379 ( .A(n25267), .Z(n25269) );
  NOR U38380 ( .A(n25269), .B(n25268), .Z(n33643) );
  IV U38381 ( .A(n25270), .Z(n25271) );
  NOR U38382 ( .A(n25272), .B(n25271), .Z(n31755) );
  NOR U38383 ( .A(n33643), .B(n31755), .Z(n30277) );
  IV U38384 ( .A(n25273), .Z(n25274) );
  NOR U38385 ( .A(n25275), .B(n25274), .Z(n28487) );
  IV U38386 ( .A(n25276), .Z(n25278) );
  NOR U38387 ( .A(n25278), .B(n25277), .Z(n28489) );
  NOR U38388 ( .A(n28487), .B(n28489), .Z(n27318) );
  IV U38389 ( .A(n25279), .Z(n25280) );
  NOR U38390 ( .A(n25281), .B(n25280), .Z(n28496) );
  IV U38391 ( .A(n25282), .Z(n25283) );
  NOR U38392 ( .A(n25284), .B(n25283), .Z(n28492) );
  NOR U38393 ( .A(n28496), .B(n28492), .Z(n27317) );
  IV U38394 ( .A(n25285), .Z(n25286) );
  NOR U38395 ( .A(n25287), .B(n25286), .Z(n27315) );
  IV U38396 ( .A(n27315), .Z(n27306) );
  IV U38397 ( .A(n25288), .Z(n25290) );
  NOR U38398 ( .A(n25290), .B(n25289), .Z(n37037) );
  IV U38399 ( .A(n25291), .Z(n25292) );
  NOR U38400 ( .A(n25293), .B(n25292), .Z(n35123) );
  NOR U38401 ( .A(n37037), .B(n35123), .Z(n28504) );
  IV U38402 ( .A(n25294), .Z(n25296) );
  NOR U38403 ( .A(n25296), .B(n25295), .Z(n31778) );
  IV U38404 ( .A(n25297), .Z(n25298) );
  NOR U38405 ( .A(n25299), .B(n25298), .Z(n31773) );
  NOR U38406 ( .A(n31778), .B(n31773), .Z(n28510) );
  IV U38407 ( .A(n25300), .Z(n25301) );
  NOR U38408 ( .A(n25302), .B(n25301), .Z(n35134) );
  IV U38409 ( .A(n25303), .Z(n25304) );
  NOR U38410 ( .A(n25305), .B(n25304), .Z(n37026) );
  NOR U38411 ( .A(n35134), .B(n37026), .Z(n31784) );
  IV U38412 ( .A(n25306), .Z(n25307) );
  NOR U38413 ( .A(n25308), .B(n25307), .Z(n33595) );
  IV U38414 ( .A(n25309), .Z(n25310) );
  NOR U38415 ( .A(n25311), .B(n25310), .Z(n31785) );
  NOR U38416 ( .A(n33595), .B(n31785), .Z(n28516) );
  IV U38417 ( .A(n25312), .Z(n25313) );
  NOR U38418 ( .A(n25314), .B(n25313), .Z(n28513) );
  IV U38419 ( .A(n25315), .Z(n25316) );
  NOR U38420 ( .A(n25317), .B(n25316), .Z(n33589) );
  IV U38421 ( .A(n25318), .Z(n25320) );
  NOR U38422 ( .A(n25320), .B(n25319), .Z(n33582) );
  NOR U38423 ( .A(n33589), .B(n33582), .Z(n28520) );
  IV U38424 ( .A(n25321), .Z(n25322) );
  NOR U38425 ( .A(n25323), .B(n25322), .Z(n31795) );
  IV U38426 ( .A(n25324), .Z(n25326) );
  NOR U38427 ( .A(n25326), .B(n25325), .Z(n31789) );
  NOR U38428 ( .A(n31795), .B(n31789), .Z(n28518) );
  IV U38429 ( .A(n25327), .Z(n25328) );
  NOR U38430 ( .A(n25329), .B(n25328), .Z(n30260) );
  IV U38431 ( .A(n25330), .Z(n25331) );
  NOR U38432 ( .A(n25332), .B(n25331), .Z(n30254) );
  NOR U38433 ( .A(n30260), .B(n30254), .Z(n27297) );
  IV U38434 ( .A(n25333), .Z(n25334) );
  NOR U38435 ( .A(n25335), .B(n25334), .Z(n25336) );
  IV U38436 ( .A(n25336), .Z(n27292) );
  IV U38437 ( .A(n25337), .Z(n25338) );
  NOR U38438 ( .A(n25339), .B(n25338), .Z(n28526) );
  IV U38439 ( .A(n25340), .Z(n25341) );
  NOR U38440 ( .A(n25342), .B(n25341), .Z(n30231) );
  NOR U38441 ( .A(n28526), .B(n30231), .Z(n27278) );
  IV U38442 ( .A(n25343), .Z(n25344) );
  NOR U38443 ( .A(n25345), .B(n25344), .Z(n35163) );
  IV U38444 ( .A(n25346), .Z(n25347) );
  NOR U38445 ( .A(n25348), .B(n25347), .Z(n35153) );
  NOR U38446 ( .A(n35163), .B(n35153), .Z(n30207) );
  IV U38447 ( .A(n25349), .Z(n25350) );
  NOR U38448 ( .A(n25351), .B(n25350), .Z(n30194) );
  IV U38449 ( .A(n25352), .Z(n25353) );
  NOR U38450 ( .A(n25354), .B(n25353), .Z(n28531) );
  NOR U38451 ( .A(n30194), .B(n28531), .Z(n30189) );
  IV U38452 ( .A(n25355), .Z(n25357) );
  NOR U38453 ( .A(n25357), .B(n25356), .Z(n27261) );
  IV U38454 ( .A(n27261), .Z(n27256) );
  IV U38455 ( .A(n25358), .Z(n25359) );
  NOR U38456 ( .A(n25360), .B(n25359), .Z(n28535) );
  IV U38457 ( .A(n25361), .Z(n25362) );
  NOR U38458 ( .A(n25363), .B(n25362), .Z(n33545) );
  IV U38459 ( .A(n25364), .Z(n25366) );
  NOR U38460 ( .A(n25366), .B(n25365), .Z(n33550) );
  NOR U38461 ( .A(n33545), .B(n33550), .Z(n30179) );
  IV U38462 ( .A(n25367), .Z(n25369) );
  NOR U38463 ( .A(n25369), .B(n25368), .Z(n33543) );
  IV U38464 ( .A(n25370), .Z(n25371) );
  NOR U38465 ( .A(n25372), .B(n25371), .Z(n25373) );
  NOR U38466 ( .A(n33543), .B(n25373), .Z(n28540) );
  IV U38467 ( .A(n25374), .Z(n25376) );
  NOR U38468 ( .A(n25376), .B(n25375), .Z(n30175) );
  IV U38469 ( .A(n25377), .Z(n25378) );
  NOR U38470 ( .A(n25379), .B(n25378), .Z(n28547) );
  IV U38471 ( .A(n25380), .Z(n25382) );
  NOR U38472 ( .A(n25382), .B(n25381), .Z(n28553) );
  IV U38473 ( .A(n25383), .Z(n25384) );
  NOR U38474 ( .A(n25385), .B(n25384), .Z(n30165) );
  NOR U38475 ( .A(n28553), .B(n30165), .Z(n27232) );
  IV U38476 ( .A(n25386), .Z(n25387) );
  NOR U38477 ( .A(n25388), .B(n25387), .Z(n33529) );
  IV U38478 ( .A(n25389), .Z(n25391) );
  NOR U38479 ( .A(n25391), .B(n25390), .Z(n33520) );
  NOR U38480 ( .A(n33529), .B(n33520), .Z(n28552) );
  IV U38481 ( .A(n25392), .Z(n25393) );
  NOR U38482 ( .A(n25394), .B(n25393), .Z(n33506) );
  IV U38483 ( .A(n25395), .Z(n25396) );
  NOR U38484 ( .A(n25397), .B(n25396), .Z(n31833) );
  NOR U38485 ( .A(n33506), .B(n31833), .Z(n28557) );
  IV U38486 ( .A(n25398), .Z(n25399) );
  NOR U38487 ( .A(n25400), .B(n25399), .Z(n33498) );
  IV U38488 ( .A(n25401), .Z(n25403) );
  NOR U38489 ( .A(n25403), .B(n25402), .Z(n33509) );
  NOR U38490 ( .A(n33498), .B(n33509), .Z(n28560) );
  IV U38491 ( .A(n25404), .Z(n25405) );
  NOR U38492 ( .A(n25406), .B(n25405), .Z(n28558) );
  IV U38493 ( .A(n25407), .Z(n25409) );
  NOR U38494 ( .A(n25409), .B(n25408), .Z(n31845) );
  IV U38495 ( .A(n25410), .Z(n25412) );
  NOR U38496 ( .A(n25412), .B(n25411), .Z(n31841) );
  NOR U38497 ( .A(n31845), .B(n31841), .Z(n28564) );
  IV U38498 ( .A(n25413), .Z(n25414) );
  NOR U38499 ( .A(n25415), .B(n25414), .Z(n31852) );
  IV U38500 ( .A(n25416), .Z(n25417) );
  NOR U38501 ( .A(n25418), .B(n25417), .Z(n31848) );
  NOR U38502 ( .A(n31852), .B(n31848), .Z(n28562) );
  IV U38503 ( .A(n25419), .Z(n25421) );
  NOR U38504 ( .A(n25421), .B(n25420), .Z(n33490) );
  IV U38505 ( .A(n25422), .Z(n25423) );
  NOR U38506 ( .A(n25424), .B(n25423), .Z(n31855) );
  NOR U38507 ( .A(n33490), .B(n31855), .Z(n25425) );
  IV U38508 ( .A(n25425), .Z(n28567) );
  IV U38509 ( .A(n25426), .Z(n25427) );
  NOR U38510 ( .A(n25428), .B(n25427), .Z(n28566) );
  IV U38511 ( .A(n28566), .Z(n33484) );
  IV U38512 ( .A(n25429), .Z(n25430) );
  NOR U38513 ( .A(n25431), .B(n25430), .Z(n30152) );
  IV U38514 ( .A(n25432), .Z(n25433) );
  NOR U38515 ( .A(n25434), .B(n25433), .Z(n30158) );
  NOR U38516 ( .A(n30152), .B(n30158), .Z(n27231) );
  IV U38517 ( .A(n25435), .Z(n25436) );
  NOR U38518 ( .A(n25437), .B(n25436), .Z(n28570) );
  IV U38519 ( .A(n25438), .Z(n25440) );
  NOR U38520 ( .A(n25440), .B(n25439), .Z(n30154) );
  NOR U38521 ( .A(n28570), .B(n30154), .Z(n27229) );
  IV U38522 ( .A(n25441), .Z(n25442) );
  NOR U38523 ( .A(n25443), .B(n25442), .Z(n25444) );
  IV U38524 ( .A(n25444), .Z(n28574) );
  IV U38525 ( .A(n25445), .Z(n25446) );
  NOR U38526 ( .A(n25447), .B(n25446), .Z(n31871) );
  IV U38527 ( .A(n31871), .Z(n27218) );
  IV U38528 ( .A(n25448), .Z(n25450) );
  NOR U38529 ( .A(n25450), .B(n25449), .Z(n36874) );
  IV U38530 ( .A(n25451), .Z(n25453) );
  NOR U38531 ( .A(n25453), .B(n25452), .Z(n36881) );
  NOR U38532 ( .A(n36874), .B(n36881), .Z(n31879) );
  IV U38533 ( .A(n25454), .Z(n25455) );
  NOR U38534 ( .A(n25456), .B(n25455), .Z(n33459) );
  IV U38535 ( .A(n25457), .Z(n25458) );
  NOR U38536 ( .A(n25459), .B(n25458), .Z(n33466) );
  NOR U38537 ( .A(n33459), .B(n33466), .Z(n28581) );
  IV U38538 ( .A(n25460), .Z(n25462) );
  NOR U38539 ( .A(n25462), .B(n25461), .Z(n33458) );
  IV U38540 ( .A(n25463), .Z(n25465) );
  NOR U38541 ( .A(n25465), .B(n25464), .Z(n25466) );
  NOR U38542 ( .A(n33458), .B(n25466), .Z(n28586) );
  IV U38543 ( .A(n25467), .Z(n25468) );
  NOR U38544 ( .A(n25469), .B(n25468), .Z(n30129) );
  IV U38545 ( .A(n25470), .Z(n25472) );
  NOR U38546 ( .A(n25472), .B(n25471), .Z(n30143) );
  NOR U38547 ( .A(n30129), .B(n30143), .Z(n27209) );
  IV U38548 ( .A(n25473), .Z(n25475) );
  NOR U38549 ( .A(n25475), .B(n25474), .Z(n30136) );
  IV U38550 ( .A(n25476), .Z(n25478) );
  NOR U38551 ( .A(n25478), .B(n25477), .Z(n30132) );
  NOR U38552 ( .A(n30136), .B(n30132), .Z(n27208) );
  IV U38553 ( .A(n25479), .Z(n25480) );
  NOR U38554 ( .A(n25481), .B(n25480), .Z(n25482) );
  IV U38555 ( .A(n25482), .Z(n27203) );
  IV U38556 ( .A(n25483), .Z(n25485) );
  NOR U38557 ( .A(n25485), .B(n25484), .Z(n31893) );
  IV U38558 ( .A(n25486), .Z(n25488) );
  NOR U38559 ( .A(n25488), .B(n25487), .Z(n33431) );
  NOR U38560 ( .A(n31893), .B(n33431), .Z(n30122) );
  IV U38561 ( .A(n25489), .Z(n25491) );
  NOR U38562 ( .A(n25491), .B(n25490), .Z(n30105) );
  IV U38563 ( .A(n25492), .Z(n25493) );
  NOR U38564 ( .A(n25494), .B(n25493), .Z(n28589) );
  NOR U38565 ( .A(n30105), .B(n28589), .Z(n27195) );
  IV U38566 ( .A(n25495), .Z(n25497) );
  NOR U38567 ( .A(n25497), .B(n25496), .Z(n30110) );
  IV U38568 ( .A(n25498), .Z(n25499) );
  NOR U38569 ( .A(n25500), .B(n25499), .Z(n33418) );
  IV U38570 ( .A(n25501), .Z(n25502) );
  NOR U38571 ( .A(n25503), .B(n25502), .Z(n31903) );
  NOR U38572 ( .A(n33418), .B(n31903), .Z(n30096) );
  IV U38573 ( .A(n25504), .Z(n25505) );
  NOR U38574 ( .A(n25506), .B(n25505), .Z(n33420) );
  IV U38575 ( .A(n33420), .Z(n28595) );
  IV U38576 ( .A(n25507), .Z(n25508) );
  NOR U38577 ( .A(n25509), .B(n25508), .Z(n31913) );
  IV U38578 ( .A(n25510), .Z(n25511) );
  NOR U38579 ( .A(n25512), .B(n25511), .Z(n31909) );
  NOR U38580 ( .A(n31913), .B(n31909), .Z(n30090) );
  IV U38581 ( .A(n25513), .Z(n25515) );
  NOR U38582 ( .A(n25515), .B(n25514), .Z(n30079) );
  IV U38583 ( .A(n25516), .Z(n25518) );
  NOR U38584 ( .A(n25518), .B(n25517), .Z(n30086) );
  NOR U38585 ( .A(n30079), .B(n30086), .Z(n27187) );
  IV U38586 ( .A(n25519), .Z(n25521) );
  NOR U38587 ( .A(n25521), .B(n25520), .Z(n33400) );
  IV U38588 ( .A(n25522), .Z(n25524) );
  NOR U38589 ( .A(n25524), .B(n25523), .Z(n25525) );
  NOR U38590 ( .A(n33400), .B(n25525), .Z(n30069) );
  IV U38591 ( .A(n25526), .Z(n25527) );
  NOR U38592 ( .A(n25528), .B(n25527), .Z(n31923) );
  IV U38593 ( .A(n25529), .Z(n25530) );
  NOR U38594 ( .A(n25531), .B(n25530), .Z(n31919) );
  NOR U38595 ( .A(n31923), .B(n31919), .Z(n28598) );
  IV U38596 ( .A(n25532), .Z(n25533) );
  NOR U38597 ( .A(n25534), .B(n25533), .Z(n25535) );
  IV U38598 ( .A(n25535), .Z(n27175) );
  IV U38599 ( .A(n25536), .Z(n25537) );
  NOR U38600 ( .A(n25538), .B(n25537), .Z(n28604) );
  IV U38601 ( .A(n25539), .Z(n25540) );
  NOR U38602 ( .A(n25541), .B(n25540), .Z(n31946) );
  IV U38603 ( .A(n25542), .Z(n25543) );
  NOR U38604 ( .A(n25544), .B(n25543), .Z(n33380) );
  NOR U38605 ( .A(n31946), .B(n33380), .Z(n30058) );
  IV U38606 ( .A(n25545), .Z(n25546) );
  NOR U38607 ( .A(n25547), .B(n25546), .Z(n36775) );
  IV U38608 ( .A(n25548), .Z(n25550) );
  NOR U38609 ( .A(n25550), .B(n25549), .Z(n35294) );
  NOR U38610 ( .A(n36775), .B(n35294), .Z(n30057) );
  IV U38611 ( .A(n25551), .Z(n25553) );
  NOR U38612 ( .A(n25553), .B(n25552), .Z(n30042) );
  IV U38613 ( .A(n25554), .Z(n25555) );
  NOR U38614 ( .A(n25556), .B(n25555), .Z(n30053) );
  NOR U38615 ( .A(n30042), .B(n30053), .Z(n27146) );
  IV U38616 ( .A(n25557), .Z(n25559) );
  NOR U38617 ( .A(n25559), .B(n25558), .Z(n30047) );
  IV U38618 ( .A(n25560), .Z(n25562) );
  NOR U38619 ( .A(n25562), .B(n25561), .Z(n31962) );
  IV U38620 ( .A(n25563), .Z(n25564) );
  NOR U38621 ( .A(n25565), .B(n25564), .Z(n31958) );
  NOR U38622 ( .A(n31962), .B(n31958), .Z(n30036) );
  IV U38623 ( .A(n25566), .Z(n25567) );
  NOR U38624 ( .A(n25568), .B(n25567), .Z(n27134) );
  IV U38625 ( .A(n27134), .Z(n27127) );
  IV U38626 ( .A(n25569), .Z(n25571) );
  NOR U38627 ( .A(n25571), .B(n25570), .Z(n30026) );
  IV U38628 ( .A(n25572), .Z(n25573) );
  NOR U38629 ( .A(n25574), .B(n25573), .Z(n30022) );
  IV U38630 ( .A(n25575), .Z(n25576) );
  NOR U38631 ( .A(n25577), .B(n25576), .Z(n28614) );
  NOR U38632 ( .A(n30022), .B(n28614), .Z(n27119) );
  IV U38633 ( .A(n25578), .Z(n25580) );
  NOR U38634 ( .A(n25580), .B(n25579), .Z(n35330) );
  IV U38635 ( .A(n25581), .Z(n25582) );
  NOR U38636 ( .A(n25583), .B(n25582), .Z(n35325) );
  NOR U38637 ( .A(n35330), .B(n35325), .Z(n31978) );
  IV U38638 ( .A(n25584), .Z(n25585) );
  NOR U38639 ( .A(n25586), .B(n25585), .Z(n28616) );
  IV U38640 ( .A(n25587), .Z(n25588) );
  NOR U38641 ( .A(n25589), .B(n25588), .Z(n33349) );
  NOR U38642 ( .A(n28616), .B(n33349), .Z(n27104) );
  IV U38643 ( .A(n25590), .Z(n25591) );
  NOR U38644 ( .A(n25592), .B(n25591), .Z(n35343) );
  IV U38645 ( .A(n25593), .Z(n25595) );
  NOR U38646 ( .A(n25595), .B(n25594), .Z(n35335) );
  NOR U38647 ( .A(n35343), .B(n35335), .Z(n29992) );
  IV U38648 ( .A(n25596), .Z(n25597) );
  NOR U38649 ( .A(n25598), .B(n25597), .Z(n29978) );
  IV U38650 ( .A(n25599), .Z(n25600) );
  NOR U38651 ( .A(n25601), .B(n25600), .Z(n29987) );
  NOR U38652 ( .A(n29978), .B(n29987), .Z(n27103) );
  IV U38653 ( .A(n25602), .Z(n25603) );
  NOR U38654 ( .A(n25604), .B(n25603), .Z(n28623) );
  IV U38655 ( .A(n25605), .Z(n25607) );
  NOR U38656 ( .A(n25607), .B(n25606), .Z(n29972) );
  NOR U38657 ( .A(n28623), .B(n29972), .Z(n27095) );
  IV U38658 ( .A(n25608), .Z(n25609) );
  NOR U38659 ( .A(n25610), .B(n25609), .Z(n32002) );
  IV U38660 ( .A(n25611), .Z(n25613) );
  NOR U38661 ( .A(n25613), .B(n25612), .Z(n31998) );
  NOR U38662 ( .A(n32002), .B(n31998), .Z(n29967) );
  IV U38663 ( .A(n25614), .Z(n25615) );
  NOR U38664 ( .A(n25616), .B(n25615), .Z(n28634) );
  IV U38665 ( .A(n25617), .Z(n25618) );
  NOR U38666 ( .A(n25619), .B(n25618), .Z(n32012) );
  IV U38667 ( .A(n25620), .Z(n25621) );
  NOR U38668 ( .A(n25622), .B(n25621), .Z(n33313) );
  NOR U38669 ( .A(n32012), .B(n33313), .Z(n29937) );
  IV U38670 ( .A(n25623), .Z(n25624) );
  NOR U38671 ( .A(n25625), .B(n25624), .Z(n29916) );
  IV U38672 ( .A(n25626), .Z(n25627) );
  NOR U38673 ( .A(n25628), .B(n25627), .Z(n29905) );
  IV U38674 ( .A(n25629), .Z(n25631) );
  NOR U38675 ( .A(n25631), .B(n25630), .Z(n29913) );
  NOR U38676 ( .A(n29905), .B(n29913), .Z(n27046) );
  IV U38677 ( .A(n25632), .Z(n25634) );
  NOR U38678 ( .A(n25634), .B(n25633), .Z(n27038) );
  IV U38679 ( .A(n27038), .Z(n27031) );
  IV U38680 ( .A(n25635), .Z(n25636) );
  NOR U38681 ( .A(n25637), .B(n25636), .Z(n27035) );
  IV U38682 ( .A(n27035), .Z(n29899) );
  IV U38683 ( .A(n25638), .Z(n25639) );
  NOR U38684 ( .A(n25640), .B(n25639), .Z(n32044) );
  IV U38685 ( .A(n25641), .Z(n25643) );
  NOR U38686 ( .A(n25643), .B(n25642), .Z(n32037) );
  NOR U38687 ( .A(n32044), .B(n32037), .Z(n29890) );
  IV U38688 ( .A(n25644), .Z(n25646) );
  NOR U38689 ( .A(n25646), .B(n25645), .Z(n27006) );
  IV U38690 ( .A(n25647), .Z(n25648) );
  NOR U38691 ( .A(n25649), .B(n25648), .Z(n27008) );
  IV U38692 ( .A(n25650), .Z(n25651) );
  NOR U38693 ( .A(n25652), .B(n25651), .Z(n29855) );
  IV U38694 ( .A(n25653), .Z(n25654) );
  NOR U38695 ( .A(n25655), .B(n25654), .Z(n29864) );
  IV U38696 ( .A(n25656), .Z(n25657) );
  NOR U38697 ( .A(n25658), .B(n25657), .Z(n29876) );
  NOR U38698 ( .A(n29864), .B(n29876), .Z(n29861) );
  IV U38699 ( .A(n25659), .Z(n25660) );
  NOR U38700 ( .A(n25661), .B(n25660), .Z(n29823) );
  IV U38701 ( .A(n25662), .Z(n25663) );
  NOR U38702 ( .A(n25664), .B(n25663), .Z(n29806) );
  IV U38703 ( .A(n25665), .Z(n25667) );
  NOR U38704 ( .A(n25667), .B(n25666), .Z(n28654) );
  IV U38705 ( .A(n25668), .Z(n25669) );
  NOR U38706 ( .A(n25670), .B(n25669), .Z(n28663) );
  IV U38707 ( .A(n25671), .Z(n25673) );
  NOR U38708 ( .A(n25673), .B(n25672), .Z(n28660) );
  NOR U38709 ( .A(n28663), .B(n28660), .Z(n26939) );
  IV U38710 ( .A(n25674), .Z(n25675) );
  NOR U38711 ( .A(n25676), .B(n25675), .Z(n26916) );
  IV U38712 ( .A(n26916), .Z(n26911) );
  IV U38713 ( .A(n25677), .Z(n25678) );
  NOR U38714 ( .A(n25679), .B(n25678), .Z(n28675) );
  IV U38715 ( .A(n25680), .Z(n25681) );
  NOR U38716 ( .A(n25682), .B(n25681), .Z(n33208) );
  IV U38717 ( .A(n25683), .Z(n25685) );
  NOR U38718 ( .A(n25685), .B(n25684), .Z(n32127) );
  NOR U38719 ( .A(n33208), .B(n32127), .Z(n28679) );
  IV U38720 ( .A(n25686), .Z(n25688) );
  NOR U38721 ( .A(n25688), .B(n25687), .Z(n28686) );
  IV U38722 ( .A(n25689), .Z(n25690) );
  NOR U38723 ( .A(n25691), .B(n25690), .Z(n28683) );
  NOR U38724 ( .A(n28686), .B(n28683), .Z(n26909) );
  IV U38725 ( .A(n25692), .Z(n25694) );
  NOR U38726 ( .A(n25694), .B(n25693), .Z(n29781) );
  IV U38727 ( .A(n25695), .Z(n25697) );
  NOR U38728 ( .A(n25697), .B(n25696), .Z(n33182) );
  IV U38729 ( .A(n25698), .Z(n25699) );
  NOR U38730 ( .A(n25700), .B(n25699), .Z(n32133) );
  NOR U38731 ( .A(n33182), .B(n32133), .Z(n29773) );
  IV U38732 ( .A(n25701), .Z(n25702) );
  NOR U38733 ( .A(n25703), .B(n25702), .Z(n33177) );
  IV U38734 ( .A(n25704), .Z(n25705) );
  NOR U38735 ( .A(n25706), .B(n25705), .Z(n33185) );
  NOR U38736 ( .A(n33177), .B(n33185), .Z(n29763) );
  IV U38737 ( .A(n25707), .Z(n25709) );
  NOR U38738 ( .A(n25709), .B(n25708), .Z(n28691) );
  IV U38739 ( .A(n25710), .Z(n25712) );
  NOR U38740 ( .A(n25712), .B(n25711), .Z(n29764) );
  NOR U38741 ( .A(n28691), .B(n29764), .Z(n26901) );
  IV U38742 ( .A(n25713), .Z(n25714) );
  NOR U38743 ( .A(n25715), .B(n25714), .Z(n28693) );
  IV U38744 ( .A(n25716), .Z(n25717) );
  NOR U38745 ( .A(n25718), .B(n25717), .Z(n28689) );
  NOR U38746 ( .A(n28693), .B(n28689), .Z(n26900) );
  IV U38747 ( .A(n25719), .Z(n25720) );
  NOR U38748 ( .A(n25721), .B(n25720), .Z(n28701) );
  IV U38749 ( .A(n25722), .Z(n25723) );
  NOR U38750 ( .A(n25724), .B(n25723), .Z(n33156) );
  IV U38751 ( .A(n25725), .Z(n25726) );
  NOR U38752 ( .A(n25727), .B(n25726), .Z(n33172) );
  NOR U38753 ( .A(n33156), .B(n33172), .Z(n28700) );
  IV U38754 ( .A(n25728), .Z(n25729) );
  NOR U38755 ( .A(n25730), .B(n25729), .Z(n28711) );
  IV U38756 ( .A(n25731), .Z(n25733) );
  NOR U38757 ( .A(n25733), .B(n25732), .Z(n28708) );
  NOR U38758 ( .A(n28711), .B(n28708), .Z(n26892) );
  IV U38759 ( .A(n25734), .Z(n25736) );
  NOR U38760 ( .A(n25736), .B(n25735), .Z(n25737) );
  IV U38761 ( .A(n25737), .Z(n28716) );
  IV U38762 ( .A(n25738), .Z(n25740) );
  NOR U38763 ( .A(n25740), .B(n25739), .Z(n28723) );
  IV U38764 ( .A(n25741), .Z(n25742) );
  NOR U38765 ( .A(n25743), .B(n25742), .Z(n28730) );
  IV U38766 ( .A(n25744), .Z(n25745) );
  NOR U38767 ( .A(n25746), .B(n25745), .Z(n28725) );
  NOR U38768 ( .A(n28730), .B(n28725), .Z(n26870) );
  IV U38769 ( .A(n25747), .Z(n25748) );
  NOR U38770 ( .A(n25749), .B(n25748), .Z(n26834) );
  IV U38771 ( .A(n26834), .Z(n26829) );
  IV U38772 ( .A(n25750), .Z(n25752) );
  NOR U38773 ( .A(n25752), .B(n25751), .Z(n28748) );
  IV U38774 ( .A(n25753), .Z(n25754) );
  NOR U38775 ( .A(n25755), .B(n25754), .Z(n35503) );
  IV U38776 ( .A(n25756), .Z(n25757) );
  NOR U38777 ( .A(n25758), .B(n25757), .Z(n35498) );
  NOR U38778 ( .A(n35503), .B(n35498), .Z(n32198) );
  IV U38779 ( .A(n25759), .Z(n25761) );
  NOR U38780 ( .A(n25761), .B(n25760), .Z(n35513) );
  IV U38781 ( .A(n25762), .Z(n25763) );
  NOR U38782 ( .A(n25764), .B(n25763), .Z(n25765) );
  NOR U38783 ( .A(n35513), .B(n25765), .Z(n28755) );
  IV U38784 ( .A(n25766), .Z(n25767) );
  NOR U38785 ( .A(n25768), .B(n25767), .Z(n33092) );
  IV U38786 ( .A(n25769), .Z(n25770) );
  NOR U38787 ( .A(n25771), .B(n25770), .Z(n33097) );
  NOR U38788 ( .A(n33092), .B(n33097), .Z(n28757) );
  IV U38789 ( .A(n25772), .Z(n25773) );
  NOR U38790 ( .A(n25774), .B(n25773), .Z(n26820) );
  IV U38791 ( .A(n26820), .Z(n26815) );
  IV U38792 ( .A(n25775), .Z(n25777) );
  NOR U38793 ( .A(n25777), .B(n25776), .Z(n29698) );
  IV U38794 ( .A(n25778), .Z(n25779) );
  NOR U38795 ( .A(n25780), .B(n25779), .Z(n28765) );
  NOR U38796 ( .A(n29698), .B(n28765), .Z(n26814) );
  IV U38797 ( .A(n25781), .Z(n25782) );
  NOR U38798 ( .A(n25783), .B(n25782), .Z(n28767) );
  IV U38799 ( .A(n25784), .Z(n25785) );
  NOR U38800 ( .A(n25786), .B(n25785), .Z(n29694) );
  NOR U38801 ( .A(n28767), .B(n29694), .Z(n26813) );
  IV U38802 ( .A(n25787), .Z(n25789) );
  NOR U38803 ( .A(n25789), .B(n25788), .Z(n26790) );
  IV U38804 ( .A(n26790), .Z(n26785) );
  IV U38805 ( .A(n25790), .Z(n25792) );
  NOR U38806 ( .A(n25792), .B(n25791), .Z(n28782) );
  IV U38807 ( .A(n25793), .Z(n25794) );
  NOR U38808 ( .A(n25795), .B(n25794), .Z(n35552) );
  IV U38809 ( .A(n25796), .Z(n25798) );
  NOR U38810 ( .A(n25798), .B(n25797), .Z(n36467) );
  NOR U38811 ( .A(n35552), .B(n36467), .Z(n28785) );
  IV U38812 ( .A(n25799), .Z(n25800) );
  NOR U38813 ( .A(n25801), .B(n25800), .Z(n28790) );
  IV U38814 ( .A(n25802), .Z(n25804) );
  NOR U38815 ( .A(n25804), .B(n25803), .Z(n28786) );
  NOR U38816 ( .A(n28790), .B(n28786), .Z(n26783) );
  IV U38817 ( .A(n25805), .Z(n25806) );
  NOR U38818 ( .A(n25807), .B(n25806), .Z(n33048) );
  IV U38819 ( .A(n25808), .Z(n25809) );
  NOR U38820 ( .A(n25810), .B(n25809), .Z(n32219) );
  NOR U38821 ( .A(n33048), .B(n32219), .Z(n28789) );
  IV U38822 ( .A(n25811), .Z(n25812) );
  NOR U38823 ( .A(n25813), .B(n25812), .Z(n28797) );
  IV U38824 ( .A(n25814), .Z(n25815) );
  NOR U38825 ( .A(n25816), .B(n25815), .Z(n28794) );
  NOR U38826 ( .A(n28797), .B(n28794), .Z(n26782) );
  IV U38827 ( .A(n25817), .Z(n25819) );
  NOR U38828 ( .A(n25819), .B(n25818), .Z(n29663) );
  IV U38829 ( .A(n25820), .Z(n25822) );
  NOR U38830 ( .A(n25822), .B(n25821), .Z(n33018) );
  IV U38831 ( .A(n25823), .Z(n25824) );
  NOR U38832 ( .A(n25825), .B(n25824), .Z(n33034) );
  NOR U38833 ( .A(n33018), .B(n33034), .Z(n29658) );
  IV U38834 ( .A(n25826), .Z(n25827) );
  NOR U38835 ( .A(n25828), .B(n25827), .Z(n26764) );
  IV U38836 ( .A(n26764), .Z(n26757) );
  IV U38837 ( .A(n25829), .Z(n25830) );
  NOR U38838 ( .A(n25831), .B(n25830), .Z(n25832) );
  IV U38839 ( .A(n25832), .Z(n28801) );
  IV U38840 ( .A(n25833), .Z(n25834) );
  NOR U38841 ( .A(n25835), .B(n25834), .Z(n32223) );
  IV U38842 ( .A(n25836), .Z(n25837) );
  NOR U38843 ( .A(n25838), .B(n25837), .Z(n33000) );
  NOR U38844 ( .A(n32223), .B(n33000), .Z(n29648) );
  IV U38845 ( .A(n25839), .Z(n25840) );
  NOR U38846 ( .A(n25841), .B(n25840), .Z(n25842) );
  IV U38847 ( .A(n25842), .Z(n29640) );
  IV U38848 ( .A(n25843), .Z(n25844) );
  NOR U38849 ( .A(n46500), .B(n25844), .Z(n32976) );
  IV U38850 ( .A(n25845), .Z(n25846) );
  NOR U38851 ( .A(n25847), .B(n25846), .Z(n29616) );
  IV U38852 ( .A(n25848), .Z(n25849) );
  NOR U38853 ( .A(n25850), .B(n25849), .Z(n29612) );
  NOR U38854 ( .A(n29616), .B(n29612), .Z(n26714) );
  IV U38855 ( .A(n25851), .Z(n25852) );
  NOR U38856 ( .A(n25853), .B(n25852), .Z(n32261) );
  IV U38857 ( .A(n25854), .Z(n25856) );
  NOR U38858 ( .A(n25856), .B(n25855), .Z(n32257) );
  NOR U38859 ( .A(n32261), .B(n32257), .Z(n29608) );
  IV U38860 ( .A(n25857), .Z(n25859) );
  NOR U38861 ( .A(n25859), .B(n25858), .Z(n29600) );
  IV U38862 ( .A(n25860), .Z(n25861) );
  NOR U38863 ( .A(n25862), .B(n25861), .Z(n29604) );
  NOR U38864 ( .A(n29600), .B(n29604), .Z(n26713) );
  IV U38865 ( .A(n25863), .Z(n25865) );
  NOR U38866 ( .A(n25865), .B(n25864), .Z(n29581) );
  IV U38867 ( .A(n25866), .Z(n25867) );
  NOR U38868 ( .A(n25868), .B(n25867), .Z(n28819) );
  IV U38869 ( .A(n25869), .Z(n25871) );
  NOR U38870 ( .A(n25871), .B(n25870), .Z(n32940) );
  IV U38871 ( .A(n25872), .Z(n25873) );
  NOR U38872 ( .A(n25874), .B(n25873), .Z(n32947) );
  NOR U38873 ( .A(n32940), .B(n32947), .Z(n29547) );
  IV U38874 ( .A(n25875), .Z(n25876) );
  NOR U38875 ( .A(n25877), .B(n25876), .Z(n36336) );
  IV U38876 ( .A(n25878), .Z(n25880) );
  NOR U38877 ( .A(n25880), .B(n25879), .Z(n36343) );
  NOR U38878 ( .A(n36336), .B(n36343), .Z(n29550) );
  IV U38879 ( .A(n25881), .Z(n25882) );
  NOR U38880 ( .A(n25883), .B(n25882), .Z(n26646) );
  IV U38881 ( .A(n26646), .Z(n26641) );
  IV U38882 ( .A(n25884), .Z(n25885) );
  NOR U38883 ( .A(n25886), .B(n25885), .Z(n28840) );
  IV U38884 ( .A(n25887), .Z(n25888) );
  NOR U38885 ( .A(n25889), .B(n25888), .Z(n32916) );
  IV U38886 ( .A(n25890), .Z(n25891) );
  NOR U38887 ( .A(n25892), .B(n25891), .Z(n32922) );
  NOR U38888 ( .A(n32916), .B(n32922), .Z(n28839) );
  IV U38889 ( .A(n25893), .Z(n25895) );
  NOR U38890 ( .A(n25895), .B(n25894), .Z(n29541) );
  IV U38891 ( .A(n25896), .Z(n25898) );
  NOR U38892 ( .A(n25898), .B(n25897), .Z(n28844) );
  NOR U38893 ( .A(n29541), .B(n28844), .Z(n26639) );
  IV U38894 ( .A(n25899), .Z(n25900) );
  NOR U38895 ( .A(n25901), .B(n25900), .Z(n29539) );
  IV U38896 ( .A(n25902), .Z(n25904) );
  NOR U38897 ( .A(n25904), .B(n25903), .Z(n32285) );
  IV U38898 ( .A(n25905), .Z(n25906) );
  NOR U38899 ( .A(n25907), .B(n25906), .Z(n32907) );
  NOR U38900 ( .A(n32285), .B(n32907), .Z(n28848) );
  IV U38901 ( .A(n25908), .Z(n25909) );
  NOR U38902 ( .A(n25910), .B(n25909), .Z(n29530) );
  IV U38903 ( .A(n25911), .Z(n25913) );
  NOR U38904 ( .A(n25913), .B(n25912), .Z(n28849) );
  NOR U38905 ( .A(n29530), .B(n28849), .Z(n26638) );
  IV U38906 ( .A(n25914), .Z(n25916) );
  NOR U38907 ( .A(n25916), .B(n25915), .Z(n29523) );
  IV U38908 ( .A(n25917), .Z(n25918) );
  NOR U38909 ( .A(n25919), .B(n25918), .Z(n29518) );
  IV U38910 ( .A(n25920), .Z(n25921) );
  NOR U38911 ( .A(n25922), .B(n25921), .Z(n28860) );
  NOR U38912 ( .A(n29518), .B(n28860), .Z(n26630) );
  IV U38913 ( .A(n25923), .Z(n25925) );
  NOR U38914 ( .A(n25925), .B(n25924), .Z(n29506) );
  IV U38915 ( .A(n25926), .Z(n25927) );
  NOR U38916 ( .A(n25928), .B(n25927), .Z(n29502) );
  NOR U38917 ( .A(n29506), .B(n29502), .Z(n26629) );
  IV U38918 ( .A(n25929), .Z(n25930) );
  NOR U38919 ( .A(n25931), .B(n25930), .Z(n29497) );
  IV U38920 ( .A(n25932), .Z(n25933) );
  NOR U38921 ( .A(n25934), .B(n25933), .Z(n29491) );
  NOR U38922 ( .A(n29497), .B(n29491), .Z(n26628) );
  IV U38923 ( .A(n25935), .Z(n25936) );
  NOR U38924 ( .A(n25937), .B(n25936), .Z(n29480) );
  IV U38925 ( .A(n25938), .Z(n25939) );
  NOR U38926 ( .A(n25940), .B(n25939), .Z(n28866) );
  NOR U38927 ( .A(n29480), .B(n28866), .Z(n26606) );
  IV U38928 ( .A(n25941), .Z(n25943) );
  NOR U38929 ( .A(n25943), .B(n25942), .Z(n29458) );
  IV U38930 ( .A(n25944), .Z(n25945) );
  NOR U38931 ( .A(n25946), .B(n25945), .Z(n28868) );
  NOR U38932 ( .A(n29458), .B(n28868), .Z(n26605) );
  IV U38933 ( .A(n25947), .Z(n25948) );
  NOR U38934 ( .A(n25949), .B(n25948), .Z(n29452) );
  IV U38935 ( .A(n25950), .Z(n25951) );
  NOR U38936 ( .A(n25952), .B(n25951), .Z(n29462) );
  NOR U38937 ( .A(n29452), .B(n29462), .Z(n26604) );
  IV U38938 ( .A(n25953), .Z(n25954) );
  NOR U38939 ( .A(n25955), .B(n25954), .Z(n29435) );
  IV U38940 ( .A(n25956), .Z(n25957) );
  NOR U38941 ( .A(n25958), .B(n25957), .Z(n29419) );
  IV U38942 ( .A(n25959), .Z(n25961) );
  NOR U38943 ( .A(n25961), .B(n25960), .Z(n32858) );
  IV U38944 ( .A(n25962), .Z(n25963) );
  NOR U38945 ( .A(n25964), .B(n25963), .Z(n25965) );
  NOR U38946 ( .A(n32858), .B(n25965), .Z(n29415) );
  IV U38947 ( .A(n25966), .Z(n25968) );
  NOR U38948 ( .A(n25968), .B(n25967), .Z(n32350) );
  IV U38949 ( .A(n25969), .Z(n25970) );
  NOR U38950 ( .A(n25971), .B(n25970), .Z(n25972) );
  NOR U38951 ( .A(n32350), .B(n25972), .Z(n29414) );
  IV U38952 ( .A(n25973), .Z(n25974) );
  NOR U38953 ( .A(n25975), .B(n25974), .Z(n29404) );
  IV U38954 ( .A(n25976), .Z(n25977) );
  NOR U38955 ( .A(n25978), .B(n25977), .Z(n28876) );
  NOR U38956 ( .A(n29404), .B(n28876), .Z(n26568) );
  IV U38957 ( .A(n25979), .Z(n25980) );
  NOR U38958 ( .A(n25981), .B(n25980), .Z(n29406) );
  IV U38959 ( .A(n25982), .Z(n25984) );
  NOR U38960 ( .A(n25984), .B(n25983), .Z(n32365) );
  IV U38961 ( .A(n25985), .Z(n25987) );
  NOR U38962 ( .A(n25987), .B(n25986), .Z(n32361) );
  NOR U38963 ( .A(n32365), .B(n32361), .Z(n29397) );
  IV U38964 ( .A(n25988), .Z(n25989) );
  NOR U38965 ( .A(n25990), .B(n25989), .Z(n32375) );
  IV U38966 ( .A(n25991), .Z(n25992) );
  NOR U38967 ( .A(n25993), .B(n25992), .Z(n25994) );
  NOR U38968 ( .A(n32375), .B(n25994), .Z(n28879) );
  IV U38969 ( .A(n25995), .Z(n25996) );
  NOR U38970 ( .A(n25997), .B(n25996), .Z(n28880) );
  IV U38971 ( .A(n25998), .Z(n26000) );
  NOR U38972 ( .A(n26000), .B(n25999), .Z(n29392) );
  NOR U38973 ( .A(n28880), .B(n29392), .Z(n26558) );
  IV U38974 ( .A(n26001), .Z(n26002) );
  NOR U38975 ( .A(n26003), .B(n26002), .Z(n29370) );
  IV U38976 ( .A(n26004), .Z(n26005) );
  NOR U38977 ( .A(n26006), .B(n26005), .Z(n29378) );
  IV U38978 ( .A(n26007), .Z(n26008) );
  NOR U38979 ( .A(n26009), .B(n26008), .Z(n29382) );
  NOR U38980 ( .A(n29378), .B(n29382), .Z(n29375) );
  IV U38981 ( .A(n26010), .Z(n26011) );
  NOR U38982 ( .A(n26012), .B(n26011), .Z(n28884) );
  IV U38983 ( .A(n26013), .Z(n26014) );
  NOR U38984 ( .A(n26015), .B(n26014), .Z(n29364) );
  NOR U38985 ( .A(n28884), .B(n29364), .Z(n26557) );
  IV U38986 ( .A(n26016), .Z(n26018) );
  NOR U38987 ( .A(n26018), .B(n26017), .Z(n28885) );
  IV U38988 ( .A(n26019), .Z(n26021) );
  NOR U38989 ( .A(n26021), .B(n26020), .Z(n28882) );
  NOR U38990 ( .A(n28885), .B(n28882), .Z(n26556) );
  IV U38991 ( .A(n26022), .Z(n26023) );
  NOR U38992 ( .A(n26024), .B(n26023), .Z(n29348) );
  IV U38993 ( .A(n26025), .Z(n26027) );
  NOR U38994 ( .A(n26027), .B(n26026), .Z(n28892) );
  NOR U38995 ( .A(n29348), .B(n28892), .Z(n26555) );
  IV U38996 ( .A(n26028), .Z(n26029) );
  NOR U38997 ( .A(n26030), .B(n26029), .Z(n29351) );
  IV U38998 ( .A(n26031), .Z(n26032) );
  NOR U38999 ( .A(n26033), .B(n26032), .Z(n29341) );
  IV U39000 ( .A(n26034), .Z(n26036) );
  NOR U39001 ( .A(n26036), .B(n26035), .Z(n28895) );
  IV U39002 ( .A(n26037), .Z(n26038) );
  NOR U39003 ( .A(n26039), .B(n26038), .Z(n28898) );
  IV U39004 ( .A(n26040), .Z(n26042) );
  NOR U39005 ( .A(n26042), .B(n26041), .Z(n29335) );
  NOR U39006 ( .A(n28898), .B(n29335), .Z(n26545) );
  IV U39007 ( .A(n26043), .Z(n26045) );
  NOR U39008 ( .A(n26045), .B(n26044), .Z(n32401) );
  IV U39009 ( .A(n26046), .Z(n26047) );
  NOR U39010 ( .A(n26048), .B(n26047), .Z(n32395) );
  NOR U39011 ( .A(n32401), .B(n32395), .Z(n29331) );
  IV U39012 ( .A(n26049), .Z(n26051) );
  NOR U39013 ( .A(n26051), .B(n26050), .Z(n28900) );
  IV U39014 ( .A(n26052), .Z(n26054) );
  NOR U39015 ( .A(n26054), .B(n26053), .Z(n29327) );
  NOR U39016 ( .A(n28900), .B(n29327), .Z(n26544) );
  IV U39017 ( .A(n26055), .Z(n26056) );
  NOR U39018 ( .A(n26057), .B(n26056), .Z(n28913) );
  IV U39019 ( .A(n26058), .Z(n26060) );
  NOR U39020 ( .A(n26060), .B(n26059), .Z(n28905) );
  NOR U39021 ( .A(n28913), .B(n28905), .Z(n26536) );
  IV U39022 ( .A(n26061), .Z(n26062) );
  NOR U39023 ( .A(n26063), .B(n26062), .Z(n28916) );
  IV U39024 ( .A(n26064), .Z(n26065) );
  NOR U39025 ( .A(n26066), .B(n26065), .Z(n28911) );
  NOR U39026 ( .A(n28916), .B(n28911), .Z(n26535) );
  IV U39027 ( .A(n26067), .Z(n26069) );
  NOR U39028 ( .A(n26069), .B(n26068), .Z(n29317) );
  IV U39029 ( .A(n26070), .Z(n26072) );
  NOR U39030 ( .A(n26072), .B(n26071), .Z(n29323) );
  NOR U39031 ( .A(n29317), .B(n29323), .Z(n26534) );
  IV U39032 ( .A(n26073), .Z(n26075) );
  NOR U39033 ( .A(n26075), .B(n26074), .Z(n29316) );
  IV U39034 ( .A(n26076), .Z(n26077) );
  NOR U39035 ( .A(n26078), .B(n26077), .Z(n32425) );
  IV U39036 ( .A(n26079), .Z(n26080) );
  NOR U39037 ( .A(n26081), .B(n26080), .Z(n32420) );
  NOR U39038 ( .A(n32425), .B(n32420), .Z(n28920) );
  IV U39039 ( .A(n26082), .Z(n26083) );
  NOR U39040 ( .A(n26084), .B(n26083), .Z(n29254) );
  IV U39041 ( .A(n26085), .Z(n26086) );
  NOR U39042 ( .A(n26087), .B(n26086), .Z(n29251) );
  NOR U39043 ( .A(n29254), .B(n29251), .Z(n26478) );
  IV U39044 ( .A(n26088), .Z(n26090) );
  NOR U39045 ( .A(n26090), .B(n26089), .Z(n32455) );
  IV U39046 ( .A(n26091), .Z(n26092) );
  NOR U39047 ( .A(n26093), .B(n26092), .Z(n32450) );
  NOR U39048 ( .A(n32455), .B(n32450), .Z(n28932) );
  IV U39049 ( .A(n26094), .Z(n26095) );
  NOR U39050 ( .A(n26096), .B(n26095), .Z(n32743) );
  IV U39051 ( .A(n26097), .Z(n26099) );
  NOR U39052 ( .A(n26099), .B(n26098), .Z(n32458) );
  NOR U39053 ( .A(n32743), .B(n32458), .Z(n28931) );
  IV U39054 ( .A(n26100), .Z(n26102) );
  NOR U39055 ( .A(n26102), .B(n26101), .Z(n28940) );
  IV U39056 ( .A(n26103), .Z(n26105) );
  NOR U39057 ( .A(n26105), .B(n26104), .Z(n29232) );
  NOR U39058 ( .A(n28940), .B(n29232), .Z(n26458) );
  IV U39059 ( .A(n26106), .Z(n26107) );
  NOR U39060 ( .A(n26108), .B(n26107), .Z(n35879) );
  IV U39061 ( .A(n26109), .Z(n26110) );
  NOR U39062 ( .A(n26111), .B(n26110), .Z(n35871) );
  NOR U39063 ( .A(n35879), .B(n35871), .Z(n28951) );
  IV U39064 ( .A(n26112), .Z(n26113) );
  NOR U39065 ( .A(n26114), .B(n26113), .Z(n29192) );
  IV U39066 ( .A(n26115), .Z(n26116) );
  NOR U39067 ( .A(n26117), .B(n26116), .Z(n32505) );
  IV U39068 ( .A(n26118), .Z(n26120) );
  NOR U39069 ( .A(n26120), .B(n26119), .Z(n29183) );
  IV U39070 ( .A(n26121), .Z(n26123) );
  NOR U39071 ( .A(n26123), .B(n26122), .Z(n28962) );
  NOR U39072 ( .A(n29183), .B(n28962), .Z(n26400) );
  IV U39073 ( .A(n26124), .Z(n26125) );
  NOR U39074 ( .A(n26126), .B(n26125), .Z(n32512) );
  IV U39075 ( .A(n26127), .Z(n26128) );
  NOR U39076 ( .A(n26129), .B(n26128), .Z(n32516) );
  NOR U39077 ( .A(n32512), .B(n32516), .Z(n29187) );
  IV U39078 ( .A(n26130), .Z(n26132) );
  NOR U39079 ( .A(n26132), .B(n26131), .Z(n29159) );
  IV U39080 ( .A(n26133), .Z(n26134) );
  NOR U39081 ( .A(n26135), .B(n26134), .Z(n29179) );
  NOR U39082 ( .A(n29159), .B(n29179), .Z(n26399) );
  IV U39083 ( .A(n26136), .Z(n26137) );
  NOR U39084 ( .A(n26138), .B(n26137), .Z(n26139) );
  IV U39085 ( .A(n26139), .Z(n26387) );
  IV U39086 ( .A(n26140), .Z(n26141) );
  NOR U39087 ( .A(n26142), .B(n26141), .Z(n32535) );
  IV U39088 ( .A(n26143), .Z(n26144) );
  NOR U39089 ( .A(n26145), .B(n26144), .Z(n32530) );
  NOR U39090 ( .A(n32535), .B(n32530), .Z(n29153) );
  IV U39091 ( .A(n26146), .Z(n26147) );
  NOR U39092 ( .A(n26148), .B(n26147), .Z(n29127) );
  IV U39093 ( .A(n26149), .Z(n26150) );
  NOR U39094 ( .A(n26151), .B(n26150), .Z(n28967) );
  NOR U39095 ( .A(n29127), .B(n28967), .Z(n26379) );
  IV U39096 ( .A(n26152), .Z(n26154) );
  NOR U39097 ( .A(n26154), .B(n26153), .Z(n28969) );
  IV U39098 ( .A(n26155), .Z(n26157) );
  NOR U39099 ( .A(n26157), .B(n26156), .Z(n28974) );
  IV U39100 ( .A(n26158), .Z(n26159) );
  NOR U39101 ( .A(n26160), .B(n26159), .Z(n28972) );
  NOR U39102 ( .A(n28974), .B(n28972), .Z(n26354) );
  IV U39103 ( .A(n26161), .Z(n26162) );
  NOR U39104 ( .A(n26163), .B(n26162), .Z(n28980) );
  IV U39105 ( .A(n26164), .Z(n26165) );
  NOR U39106 ( .A(n26166), .B(n26165), .Z(n28978) );
  NOR U39107 ( .A(n28980), .B(n28978), .Z(n26353) );
  IV U39108 ( .A(n26167), .Z(n26169) );
  NOR U39109 ( .A(n26169), .B(n26168), .Z(n26170) );
  IV U39110 ( .A(n26170), .Z(n28990) );
  IV U39111 ( .A(n26171), .Z(n26173) );
  NOR U39112 ( .A(n26173), .B(n26172), .Z(n32652) );
  IV U39113 ( .A(n26174), .Z(n26175) );
  NOR U39114 ( .A(n26176), .B(n26175), .Z(n32551) );
  NOR U39115 ( .A(n32652), .B(n32551), .Z(n28991) );
  IV U39116 ( .A(n26177), .Z(n26178) );
  NOR U39117 ( .A(n26179), .B(n26178), .Z(n29109) );
  IV U39118 ( .A(n26180), .Z(n26182) );
  NOR U39119 ( .A(n26182), .B(n26181), .Z(n29103) );
  NOR U39120 ( .A(n29109), .B(n29103), .Z(n26345) );
  IV U39121 ( .A(n26183), .Z(n26185) );
  NOR U39122 ( .A(n26185), .B(n26184), .Z(n29008) );
  IV U39123 ( .A(n26186), .Z(n26187) );
  NOR U39124 ( .A(n26188), .B(n26187), .Z(n26321) );
  IV U39125 ( .A(n26321), .Z(n29095) );
  IV U39126 ( .A(n26189), .Z(n26191) );
  NOR U39127 ( .A(n26191), .B(n26190), .Z(n26309) );
  IV U39128 ( .A(n26309), .Z(n26300) );
  IV U39129 ( .A(n26192), .Z(n26193) );
  NOR U39130 ( .A(n26194), .B(n26193), .Z(n29012) );
  IV U39131 ( .A(n26195), .Z(n26197) );
  NOR U39132 ( .A(n26197), .B(n26196), .Z(n29025) );
  IV U39133 ( .A(n26198), .Z(n26199) );
  NOR U39134 ( .A(n26200), .B(n26199), .Z(n29029) );
  IV U39135 ( .A(n26201), .Z(n26202) );
  NOR U39136 ( .A(n26203), .B(n26202), .Z(n29022) );
  NOR U39137 ( .A(n29029), .B(n29022), .Z(n26291) );
  IV U39138 ( .A(n26204), .Z(n26205) );
  NOR U39139 ( .A(n26206), .B(n26205), .Z(n29038) );
  IV U39140 ( .A(n26207), .Z(n26208) );
  NOR U39141 ( .A(n26209), .B(n26208), .Z(n29033) );
  NOR U39142 ( .A(n29038), .B(n29033), .Z(n26284) );
  IV U39143 ( .A(n26210), .Z(n26211) );
  NOR U39144 ( .A(n26212), .B(n26211), .Z(n29041) );
  IV U39145 ( .A(n26213), .Z(n26215) );
  NOR U39146 ( .A(n26215), .B(n26214), .Z(n29051) );
  IV U39147 ( .A(n26216), .Z(n26218) );
  NOR U39148 ( .A(n26218), .B(n26217), .Z(n29076) );
  IV U39149 ( .A(n26219), .Z(n26220) );
  NOR U39150 ( .A(n26221), .B(n26220), .Z(n26255) );
  IV U39151 ( .A(n26222), .Z(n26224) );
  NOR U39152 ( .A(n26224), .B(n26223), .Z(n26252) );
  IV U39153 ( .A(n26252), .Z(n26246) );
  IV U39154 ( .A(n26225), .Z(n26226) );
  NOR U39155 ( .A(n26227), .B(n26226), .Z(n26251) );
  IV U39156 ( .A(n26228), .Z(n26229) );
  NOR U39157 ( .A(n26230), .B(n26229), .Z(n26238) );
  IV U39158 ( .A(n26231), .Z(n26233) );
  NOR U39159 ( .A(n26233), .B(n26232), .Z(n29055) );
  IV U39160 ( .A(n26234), .Z(n26235) );
  NOR U39161 ( .A(n26236), .B(n26235), .Z(n29059) );
  IV U39162 ( .A(n29059), .Z(n29057) );
  XOR U39163 ( .A(n29055), .B(n29057), .Z(n26237) );
  NOR U39164 ( .A(n26238), .B(n26237), .Z(n26244) );
  IV U39165 ( .A(n26238), .Z(n29060) );
  IV U39166 ( .A(n26239), .Z(n26241) );
  NOR U39167 ( .A(n26241), .B(n26240), .Z(n29058) );
  XOR U39168 ( .A(n29060), .B(n29058), .Z(n26242) );
  NOR U39169 ( .A(n29059), .B(n26242), .Z(n26243) );
  NOR U39170 ( .A(n26244), .B(n26243), .Z(n29064) );
  XOR U39171 ( .A(n26251), .B(n29064), .Z(n26245) );
  NOR U39172 ( .A(n26246), .B(n26245), .Z(n32611) );
  IV U39173 ( .A(n26247), .Z(n26249) );
  NOR U39174 ( .A(n26249), .B(n26248), .Z(n26250) );
  NOR U39175 ( .A(n26251), .B(n26250), .Z(n29065) );
  XOR U39176 ( .A(n29065), .B(n29064), .Z(n26256) );
  NOR U39177 ( .A(n26252), .B(n26256), .Z(n26253) );
  NOR U39178 ( .A(n32611), .B(n26253), .Z(n26254) );
  NOR U39179 ( .A(n26255), .B(n26254), .Z(n26259) );
  IV U39180 ( .A(n26255), .Z(n26258) );
  IV U39181 ( .A(n26256), .Z(n26257) );
  NOR U39182 ( .A(n26258), .B(n26257), .Z(n29080) );
  NOR U39183 ( .A(n26259), .B(n29080), .Z(n26260) );
  IV U39184 ( .A(n26260), .Z(n29077) );
  XOR U39185 ( .A(n29076), .B(n29077), .Z(n29071) );
  IV U39186 ( .A(n26261), .Z(n26263) );
  NOR U39187 ( .A(n26263), .B(n26262), .Z(n29073) );
  IV U39188 ( .A(n26264), .Z(n26266) );
  NOR U39189 ( .A(n26266), .B(n26265), .Z(n29070) );
  NOR U39190 ( .A(n29073), .B(n29070), .Z(n26267) );
  XOR U39191 ( .A(n29071), .B(n26267), .Z(n26268) );
  IV U39192 ( .A(n26268), .Z(n29053) );
  XOR U39193 ( .A(n29051), .B(n29053), .Z(n29049) );
  IV U39194 ( .A(n26269), .Z(n26271) );
  NOR U39195 ( .A(n26271), .B(n26270), .Z(n29050) );
  IV U39196 ( .A(n26272), .Z(n26273) );
  NOR U39197 ( .A(n26274), .B(n26273), .Z(n29047) );
  NOR U39198 ( .A(n29050), .B(n29047), .Z(n26275) );
  XOR U39199 ( .A(n29049), .B(n26275), .Z(n26276) );
  IV U39200 ( .A(n26276), .Z(n29042) );
  XOR U39201 ( .A(n29041), .B(n29042), .Z(n29045) );
  IV U39202 ( .A(n26277), .Z(n26278) );
  NOR U39203 ( .A(n26279), .B(n26278), .Z(n29044) );
  IV U39204 ( .A(n26280), .Z(n26281) );
  NOR U39205 ( .A(n26282), .B(n26281), .Z(n29036) );
  NOR U39206 ( .A(n29044), .B(n29036), .Z(n26283) );
  XOR U39207 ( .A(n29045), .B(n26283), .Z(n29034) );
  XOR U39208 ( .A(n26284), .B(n29034), .Z(n32622) );
  IV U39209 ( .A(n26285), .Z(n26287) );
  NOR U39210 ( .A(n26287), .B(n26286), .Z(n32587) );
  IV U39211 ( .A(n26288), .Z(n26289) );
  NOR U39212 ( .A(n26290), .B(n26289), .Z(n32621) );
  NOR U39213 ( .A(n32587), .B(n32621), .Z(n29028) );
  XOR U39214 ( .A(n32622), .B(n29028), .Z(n29023) );
  XOR U39215 ( .A(n26291), .B(n29023), .Z(n29026) );
  XOR U39216 ( .A(n29025), .B(n29026), .Z(n29018) );
  IV U39217 ( .A(n26292), .Z(n26294) );
  NOR U39218 ( .A(n26294), .B(n26293), .Z(n29020) );
  IV U39219 ( .A(n26295), .Z(n26296) );
  NOR U39220 ( .A(n26297), .B(n26296), .Z(n29017) );
  NOR U39221 ( .A(n29020), .B(n29017), .Z(n26298) );
  XOR U39222 ( .A(n29018), .B(n26298), .Z(n29011) );
  XOR U39223 ( .A(n29012), .B(n29011), .Z(n26306) );
  IV U39224 ( .A(n26306), .Z(n26299) );
  NOR U39225 ( .A(n26300), .B(n26299), .Z(n32578) );
  NOR U39226 ( .A(n29012), .B(n29011), .Z(n26305) );
  IV U39227 ( .A(n26301), .Z(n26303) );
  NOR U39228 ( .A(n26303), .B(n26302), .Z(n26307) );
  IV U39229 ( .A(n26307), .Z(n26304) );
  NOR U39230 ( .A(n26305), .B(n26304), .Z(n29010) );
  NOR U39231 ( .A(n26307), .B(n26306), .Z(n26308) );
  NOR U39232 ( .A(n29010), .B(n26308), .Z(n26315) );
  NOR U39233 ( .A(n26309), .B(n26315), .Z(n26310) );
  NOR U39234 ( .A(n32578), .B(n26310), .Z(n26318) );
  IV U39235 ( .A(n26318), .Z(n26311) );
  NOR U39236 ( .A(n29095), .B(n26311), .Z(n29089) );
  IV U39237 ( .A(n26312), .Z(n26313) );
  NOR U39238 ( .A(n26314), .B(n26313), .Z(n26319) );
  IV U39239 ( .A(n26319), .Z(n26317) );
  IV U39240 ( .A(n26315), .Z(n26316) );
  NOR U39241 ( .A(n26317), .B(n26316), .Z(n32575) );
  NOR U39242 ( .A(n26319), .B(n26318), .Z(n26320) );
  NOR U39243 ( .A(n32575), .B(n26320), .Z(n29009) );
  NOR U39244 ( .A(n26321), .B(n29009), .Z(n26322) );
  NOR U39245 ( .A(n29089), .B(n26322), .Z(n26323) );
  IV U39246 ( .A(n26323), .Z(n29092) );
  XOR U39247 ( .A(n29008), .B(n29092), .Z(n29003) );
  IV U39248 ( .A(n26324), .Z(n26326) );
  NOR U39249 ( .A(n26326), .B(n26325), .Z(n29005) );
  IV U39250 ( .A(n26327), .Z(n26328) );
  NOR U39251 ( .A(n26329), .B(n26328), .Z(n29002) );
  NOR U39252 ( .A(n29005), .B(n29002), .Z(n26330) );
  XOR U39253 ( .A(n29003), .B(n26330), .Z(n28996) );
  IV U39254 ( .A(n26331), .Z(n26332) );
  NOR U39255 ( .A(n26333), .B(n26332), .Z(n28999) );
  IV U39256 ( .A(n26334), .Z(n26335) );
  NOR U39257 ( .A(n26336), .B(n26335), .Z(n28997) );
  NOR U39258 ( .A(n28999), .B(n28997), .Z(n26337) );
  XOR U39259 ( .A(n28996), .B(n26337), .Z(n29114) );
  IV U39260 ( .A(n26338), .Z(n26339) );
  NOR U39261 ( .A(n26340), .B(n26339), .Z(n29110) );
  IV U39262 ( .A(n26341), .Z(n26342) );
  NOR U39263 ( .A(n26343), .B(n26342), .Z(n29113) );
  NOR U39264 ( .A(n29110), .B(n29113), .Z(n26344) );
  XOR U39265 ( .A(n29114), .B(n26344), .Z(n29104) );
  XOR U39266 ( .A(n26345), .B(n29104), .Z(n32553) );
  XOR U39267 ( .A(n28991), .B(n32553), .Z(n28987) );
  XOR U39268 ( .A(n28990), .B(n28987), .Z(n28984) );
  IV U39269 ( .A(n26346), .Z(n26348) );
  NOR U39270 ( .A(n26348), .B(n26347), .Z(n28986) );
  IV U39271 ( .A(n26349), .Z(n26350) );
  NOR U39272 ( .A(n26351), .B(n26350), .Z(n28983) );
  NOR U39273 ( .A(n28986), .B(n28983), .Z(n26352) );
  XOR U39274 ( .A(n28984), .B(n26352), .Z(n28977) );
  XOR U39275 ( .A(n26353), .B(n28977), .Z(n28975) );
  XOR U39276 ( .A(n26354), .B(n28975), .Z(n26355) );
  IV U39277 ( .A(n26355), .Z(n28971) );
  XOR U39278 ( .A(n28969), .B(n28971), .Z(n26366) );
  IV U39279 ( .A(n26366), .Z(n26364) );
  IV U39280 ( .A(n26356), .Z(n26357) );
  NOR U39281 ( .A(n26358), .B(n26357), .Z(n26368) );
  IV U39282 ( .A(n26359), .Z(n26361) );
  NOR U39283 ( .A(n26361), .B(n26360), .Z(n26365) );
  NOR U39284 ( .A(n26368), .B(n26365), .Z(n26362) );
  IV U39285 ( .A(n26362), .Z(n26363) );
  NOR U39286 ( .A(n26364), .B(n26363), .Z(n26371) );
  IV U39287 ( .A(n26365), .Z(n26367) );
  NOR U39288 ( .A(n26367), .B(n26366), .Z(n32673) );
  IV U39289 ( .A(n26368), .Z(n26369) );
  NOR U39290 ( .A(n28971), .B(n26369), .Z(n32665) );
  NOR U39291 ( .A(n32673), .B(n32665), .Z(n29126) );
  IV U39292 ( .A(n29126), .Z(n26370) );
  NOR U39293 ( .A(n26371), .B(n26370), .Z(n29132) );
  IV U39294 ( .A(n26372), .Z(n26373) );
  NOR U39295 ( .A(n26374), .B(n26373), .Z(n29134) );
  IV U39296 ( .A(n26375), .Z(n26376) );
  NOR U39297 ( .A(n26377), .B(n26376), .Z(n29131) );
  NOR U39298 ( .A(n29134), .B(n29131), .Z(n26378) );
  XOR U39299 ( .A(n29132), .B(n26378), .Z(n29128) );
  XOR U39300 ( .A(n26379), .B(n29128), .Z(n29152) );
  XOR U39301 ( .A(n29153), .B(n29152), .Z(n29155) );
  NOR U39302 ( .A(n26387), .B(n29155), .Z(n32684) );
  IV U39303 ( .A(n26380), .Z(n26381) );
  NOR U39304 ( .A(n26382), .B(n26381), .Z(n26383) );
  IV U39305 ( .A(n26383), .Z(n28965) );
  IV U39306 ( .A(n26384), .Z(n26385) );
  NOR U39307 ( .A(n26386), .B(n26385), .Z(n29154) );
  XOR U39308 ( .A(n29154), .B(n29155), .Z(n28964) );
  XOR U39309 ( .A(n28965), .B(n28964), .Z(n26390) );
  IV U39310 ( .A(n28964), .Z(n26388) );
  NOR U39311 ( .A(n26388), .B(n26387), .Z(n26389) );
  NOR U39312 ( .A(n26390), .B(n26389), .Z(n26391) );
  NOR U39313 ( .A(n32684), .B(n26391), .Z(n29165) );
  IV U39314 ( .A(n26392), .Z(n26393) );
  NOR U39315 ( .A(n26394), .B(n26393), .Z(n29160) );
  IV U39316 ( .A(n26395), .Z(n26396) );
  NOR U39317 ( .A(n26397), .B(n26396), .Z(n29172) );
  NOR U39318 ( .A(n29160), .B(n29172), .Z(n26398) );
  XOR U39319 ( .A(n29165), .B(n26398), .Z(n29180) );
  XOR U39320 ( .A(n26399), .B(n29180), .Z(n29186) );
  XOR U39321 ( .A(n29187), .B(n29186), .Z(n29184) );
  XOR U39322 ( .A(n26400), .B(n29184), .Z(n26401) );
  IV U39323 ( .A(n26401), .Z(n32506) );
  XOR U39324 ( .A(n32505), .B(n32506), .Z(n28957) );
  IV U39325 ( .A(n28957), .Z(n26409) );
  IV U39326 ( .A(n26402), .Z(n26404) );
  NOR U39327 ( .A(n26404), .B(n26403), .Z(n28960) );
  IV U39328 ( .A(n26405), .Z(n26407) );
  NOR U39329 ( .A(n26407), .B(n26406), .Z(n28956) );
  NOR U39330 ( .A(n28960), .B(n28956), .Z(n26408) );
  XOR U39331 ( .A(n26409), .B(n26408), .Z(n32493) );
  IV U39332 ( .A(n26410), .Z(n26412) );
  NOR U39333 ( .A(n26412), .B(n26411), .Z(n32699) );
  IV U39334 ( .A(n26413), .Z(n26414) );
  NOR U39335 ( .A(n26415), .B(n26414), .Z(n32492) );
  NOR U39336 ( .A(n32699), .B(n32492), .Z(n29191) );
  XOR U39337 ( .A(n32493), .B(n29191), .Z(n28952) );
  IV U39338 ( .A(n28952), .Z(n29193) );
  XOR U39339 ( .A(n29192), .B(n29193), .Z(n29198) );
  IV U39340 ( .A(n26416), .Z(n26418) );
  NOR U39341 ( .A(n26418), .B(n26417), .Z(n28953) );
  IV U39342 ( .A(n26419), .Z(n26421) );
  NOR U39343 ( .A(n26421), .B(n26420), .Z(n29197) );
  NOR U39344 ( .A(n28953), .B(n29197), .Z(n26422) );
  XOR U39345 ( .A(n29198), .B(n26422), .Z(n29200) );
  IV U39346 ( .A(n26423), .Z(n26424) );
  NOR U39347 ( .A(n26425), .B(n26424), .Z(n29201) );
  IV U39348 ( .A(n26426), .Z(n26428) );
  NOR U39349 ( .A(n26428), .B(n26427), .Z(n29203) );
  NOR U39350 ( .A(n29201), .B(n29203), .Z(n26429) );
  XOR U39351 ( .A(n29200), .B(n26429), .Z(n29212) );
  IV U39352 ( .A(n26430), .Z(n26432) );
  NOR U39353 ( .A(n26432), .B(n26431), .Z(n29211) );
  IV U39354 ( .A(n26433), .Z(n26435) );
  NOR U39355 ( .A(n26435), .B(n26434), .Z(n29208) );
  NOR U39356 ( .A(n29211), .B(n29208), .Z(n26436) );
  XOR U39357 ( .A(n29212), .B(n26436), .Z(n28950) );
  XOR U39358 ( .A(n28951), .B(n28950), .Z(n29228) );
  IV U39359 ( .A(n26437), .Z(n26439) );
  NOR U39360 ( .A(n26439), .B(n26438), .Z(n28948) );
  IV U39361 ( .A(n26440), .Z(n26441) );
  NOR U39362 ( .A(n26442), .B(n26441), .Z(n29227) );
  NOR U39363 ( .A(n28948), .B(n29227), .Z(n26443) );
  XOR U39364 ( .A(n29228), .B(n26443), .Z(n28945) );
  IV U39365 ( .A(n26444), .Z(n26445) );
  NOR U39366 ( .A(n26446), .B(n26445), .Z(n29224) );
  IV U39367 ( .A(n26447), .Z(n26448) );
  NOR U39368 ( .A(n26449), .B(n26448), .Z(n28946) );
  NOR U39369 ( .A(n29224), .B(n28946), .Z(n26450) );
  XOR U39370 ( .A(n28945), .B(n26450), .Z(n28943) );
  IV U39371 ( .A(n26451), .Z(n26452) );
  NOR U39372 ( .A(n26453), .B(n26452), .Z(n28942) );
  IV U39373 ( .A(n26454), .Z(n26455) );
  NOR U39374 ( .A(n26456), .B(n26455), .Z(n32727) );
  NOR U39375 ( .A(n28942), .B(n32727), .Z(n26457) );
  XOR U39376 ( .A(n28943), .B(n26457), .Z(n29236) );
  XOR U39377 ( .A(n26458), .B(n29236), .Z(n29242) );
  IV U39378 ( .A(n26459), .Z(n26460) );
  NOR U39379 ( .A(n26461), .B(n26460), .Z(n29235) );
  IV U39380 ( .A(n26462), .Z(n26463) );
  NOR U39381 ( .A(n26464), .B(n26463), .Z(n29241) );
  NOR U39382 ( .A(n29235), .B(n29241), .Z(n26465) );
  XOR U39383 ( .A(n29242), .B(n26465), .Z(n28934) );
  IV U39384 ( .A(n26466), .Z(n26467) );
  NOR U39385 ( .A(n26468), .B(n26467), .Z(n32733) );
  IV U39386 ( .A(n26469), .Z(n26470) );
  NOR U39387 ( .A(n26471), .B(n26470), .Z(n32740) );
  NOR U39388 ( .A(n32733), .B(n32740), .Z(n28935) );
  XOR U39389 ( .A(n28934), .B(n28935), .Z(n32465) );
  IV U39390 ( .A(n26472), .Z(n26474) );
  NOR U39391 ( .A(n26474), .B(n26473), .Z(n32463) );
  IV U39392 ( .A(n26475), .Z(n26476) );
  NOR U39393 ( .A(n26477), .B(n26476), .Z(n32747) );
  NOR U39394 ( .A(n32463), .B(n32747), .Z(n28936) );
  XOR U39395 ( .A(n32465), .B(n28936), .Z(n28930) );
  XOR U39396 ( .A(n28931), .B(n28930), .Z(n32451) );
  XOR U39397 ( .A(n28932), .B(n32451), .Z(n29252) );
  XOR U39398 ( .A(n26478), .B(n29252), .Z(n29269) );
  IV U39399 ( .A(n26479), .Z(n26481) );
  NOR U39400 ( .A(n26481), .B(n26480), .Z(n29247) );
  IV U39401 ( .A(n26482), .Z(n26483) );
  NOR U39402 ( .A(n26484), .B(n26483), .Z(n29268) );
  NOR U39403 ( .A(n29247), .B(n29268), .Z(n26485) );
  XOR U39404 ( .A(n29269), .B(n26485), .Z(n28929) );
  IV U39405 ( .A(n26486), .Z(n26487) );
  NOR U39406 ( .A(n26488), .B(n26487), .Z(n35846) );
  IV U39407 ( .A(n26489), .Z(n26490) );
  NOR U39408 ( .A(n26491), .B(n26490), .Z(n26492) );
  NOR U39409 ( .A(n35846), .B(n26492), .Z(n29266) );
  XOR U39410 ( .A(n28929), .B(n29266), .Z(n29284) );
  IV U39411 ( .A(n26493), .Z(n26495) );
  NOR U39412 ( .A(n26495), .B(n26494), .Z(n29275) );
  IV U39413 ( .A(n26496), .Z(n26497) );
  NOR U39414 ( .A(n26498), .B(n26497), .Z(n29283) );
  NOR U39415 ( .A(n29275), .B(n29283), .Z(n26499) );
  XOR U39416 ( .A(n29284), .B(n26499), .Z(n28926) );
  IV U39417 ( .A(n26500), .Z(n26501) );
  NOR U39418 ( .A(n26502), .B(n26501), .Z(n28927) );
  IV U39419 ( .A(n26503), .Z(n26504) );
  NOR U39420 ( .A(n26505), .B(n26504), .Z(n29290) );
  NOR U39421 ( .A(n28927), .B(n29290), .Z(n26506) );
  XOR U39422 ( .A(n28926), .B(n26506), .Z(n28924) );
  IV U39423 ( .A(n28924), .Z(n26514) );
  IV U39424 ( .A(n26507), .Z(n26509) );
  NOR U39425 ( .A(n26509), .B(n26508), .Z(n28923) );
  IV U39426 ( .A(n26510), .Z(n26512) );
  NOR U39427 ( .A(n26512), .B(n26511), .Z(n28921) );
  NOR U39428 ( .A(n28923), .B(n28921), .Z(n26513) );
  XOR U39429 ( .A(n26514), .B(n26513), .Z(n32437) );
  IV U39430 ( .A(n26515), .Z(n26516) );
  NOR U39431 ( .A(n26517), .B(n26516), .Z(n32440) );
  IV U39432 ( .A(n26518), .Z(n26519) );
  NOR U39433 ( .A(n26520), .B(n26519), .Z(n32436) );
  NOR U39434 ( .A(n32440), .B(n32436), .Z(n29294) );
  XOR U39435 ( .A(n32437), .B(n29294), .Z(n29295) );
  IV U39436 ( .A(n26521), .Z(n26522) );
  NOR U39437 ( .A(n26523), .B(n26522), .Z(n32433) );
  IV U39438 ( .A(n26524), .Z(n26525) );
  NOR U39439 ( .A(n26526), .B(n26525), .Z(n32428) );
  NOR U39440 ( .A(n32433), .B(n32428), .Z(n29296) );
  XOR U39441 ( .A(n29295), .B(n29296), .Z(n32421) );
  XOR U39442 ( .A(n28920), .B(n32421), .Z(n29305) );
  IV U39443 ( .A(n26527), .Z(n26529) );
  NOR U39444 ( .A(n26529), .B(n26528), .Z(n29302) );
  IV U39445 ( .A(n26530), .Z(n26532) );
  NOR U39446 ( .A(n26532), .B(n26531), .Z(n28919) );
  NOR U39447 ( .A(n29302), .B(n28919), .Z(n26533) );
  XOR U39448 ( .A(n29305), .B(n26533), .Z(n29318) );
  XOR U39449 ( .A(n29316), .B(n29318), .Z(n29324) );
  XOR U39450 ( .A(n26534), .B(n29324), .Z(n28910) );
  XOR U39451 ( .A(n26535), .B(n28910), .Z(n28914) );
  XOR U39452 ( .A(n26536), .B(n28914), .Z(n28902) );
  IV U39453 ( .A(n26537), .Z(n26538) );
  NOR U39454 ( .A(n26539), .B(n26538), .Z(n28907) );
  IV U39455 ( .A(n26540), .Z(n26541) );
  NOR U39456 ( .A(n26542), .B(n26541), .Z(n32808) );
  NOR U39457 ( .A(n28907), .B(n32808), .Z(n26543) );
  XOR U39458 ( .A(n28902), .B(n26543), .Z(n29328) );
  XOR U39459 ( .A(n26544), .B(n29328), .Z(n29330) );
  XOR U39460 ( .A(n29331), .B(n29330), .Z(n29336) );
  XOR U39461 ( .A(n26545), .B(n29336), .Z(n26546) );
  IV U39462 ( .A(n26546), .Z(n28896) );
  XOR U39463 ( .A(n28895), .B(n28896), .Z(n29344) );
  XOR U39464 ( .A(n29341), .B(n29344), .Z(n29356) );
  IV U39465 ( .A(n29356), .Z(n26554) );
  IV U39466 ( .A(n26547), .Z(n26548) );
  NOR U39467 ( .A(n26549), .B(n26548), .Z(n29343) );
  IV U39468 ( .A(n26550), .Z(n26552) );
  NOR U39469 ( .A(n26552), .B(n26551), .Z(n29355) );
  NOR U39470 ( .A(n29343), .B(n29355), .Z(n26553) );
  XOR U39471 ( .A(n26554), .B(n26553), .Z(n29353) );
  XOR U39472 ( .A(n29351), .B(n29353), .Z(n28893) );
  XOR U39473 ( .A(n26555), .B(n28893), .Z(n28886) );
  XOR U39474 ( .A(n26556), .B(n28886), .Z(n29365) );
  XOR U39475 ( .A(n26557), .B(n29365), .Z(n29374) );
  XOR U39476 ( .A(n29375), .B(n29374), .Z(n29371) );
  XOR U39477 ( .A(n29370), .B(n29371), .Z(n29393) );
  XOR U39478 ( .A(n26558), .B(n29393), .Z(n26559) );
  IV U39479 ( .A(n26559), .Z(n32377) );
  XOR U39480 ( .A(n28879), .B(n32377), .Z(n29399) );
  XOR U39481 ( .A(n29397), .B(n29399), .Z(n32358) );
  IV U39482 ( .A(n32358), .Z(n26567) );
  IV U39483 ( .A(n26560), .Z(n26561) );
  NOR U39484 ( .A(n26562), .B(n26561), .Z(n29396) );
  IV U39485 ( .A(n26563), .Z(n26565) );
  NOR U39486 ( .A(n26565), .B(n26564), .Z(n29409) );
  NOR U39487 ( .A(n29396), .B(n29409), .Z(n26566) );
  XOR U39488 ( .A(n26567), .B(n26566), .Z(n29408) );
  XOR U39489 ( .A(n29406), .B(n29408), .Z(n28877) );
  XOR U39490 ( .A(n26568), .B(n28877), .Z(n29413) );
  XOR U39491 ( .A(n29414), .B(n29413), .Z(n32342) );
  XOR U39492 ( .A(n29415), .B(n32342), .Z(n26569) );
  IV U39493 ( .A(n26569), .Z(n29422) );
  XOR U39494 ( .A(n29419), .B(n29422), .Z(n28874) );
  IV U39495 ( .A(n26570), .Z(n26572) );
  NOR U39496 ( .A(n26572), .B(n26571), .Z(n29421) );
  IV U39497 ( .A(n26573), .Z(n26575) );
  NOR U39498 ( .A(n26575), .B(n26574), .Z(n28873) );
  NOR U39499 ( .A(n29421), .B(n28873), .Z(n26576) );
  XOR U39500 ( .A(n28874), .B(n26576), .Z(n28870) );
  IV U39501 ( .A(n26577), .Z(n26578) );
  NOR U39502 ( .A(n26579), .B(n26578), .Z(n28871) );
  IV U39503 ( .A(n26580), .Z(n26582) );
  NOR U39504 ( .A(n26582), .B(n26581), .Z(n29432) );
  NOR U39505 ( .A(n28871), .B(n29432), .Z(n26583) );
  XOR U39506 ( .A(n28870), .B(n26583), .Z(n29438) );
  XOR U39507 ( .A(n29435), .B(n29438), .Z(n29445) );
  IV U39508 ( .A(n26584), .Z(n26586) );
  NOR U39509 ( .A(n26586), .B(n26585), .Z(n29437) );
  IV U39510 ( .A(n26587), .Z(n26588) );
  NOR U39511 ( .A(n26589), .B(n26588), .Z(n29444) );
  NOR U39512 ( .A(n29437), .B(n29444), .Z(n26590) );
  XOR U39513 ( .A(n29445), .B(n26590), .Z(n29441) );
  IV U39514 ( .A(n26591), .Z(n26592) );
  NOR U39515 ( .A(n26593), .B(n26592), .Z(n29442) );
  IV U39516 ( .A(n26594), .Z(n26596) );
  NOR U39517 ( .A(n26596), .B(n26595), .Z(n29448) );
  NOR U39518 ( .A(n29442), .B(n29448), .Z(n26597) );
  XOR U39519 ( .A(n29441), .B(n26597), .Z(n32878) );
  IV U39520 ( .A(n26598), .Z(n26600) );
  NOR U39521 ( .A(n26600), .B(n26599), .Z(n32329) );
  IV U39522 ( .A(n26601), .Z(n26603) );
  NOR U39523 ( .A(n26603), .B(n26602), .Z(n32877) );
  NOR U39524 ( .A(n32329), .B(n32877), .Z(n29455) );
  XOR U39525 ( .A(n32878), .B(n29455), .Z(n29453) );
  XOR U39526 ( .A(n26604), .B(n29453), .Z(n29460) );
  XOR U39527 ( .A(n26605), .B(n29460), .Z(n28864) );
  XOR U39528 ( .A(n26606), .B(n28864), .Z(n29484) );
  IV U39529 ( .A(n26607), .Z(n26609) );
  NOR U39530 ( .A(n26609), .B(n26608), .Z(n29478) );
  IV U39531 ( .A(n26610), .Z(n26611) );
  NOR U39532 ( .A(n26612), .B(n26611), .Z(n29483) );
  NOR U39533 ( .A(n29478), .B(n29483), .Z(n26613) );
  XOR U39534 ( .A(n29484), .B(n26613), .Z(n26614) );
  IV U39535 ( .A(n26614), .Z(n29476) );
  IV U39536 ( .A(n26615), .Z(n26617) );
  NOR U39537 ( .A(n26617), .B(n26616), .Z(n29474) );
  IV U39538 ( .A(n26618), .Z(n26620) );
  NOR U39539 ( .A(n26620), .B(n26619), .Z(n28862) );
  NOR U39540 ( .A(n29474), .B(n28862), .Z(n26621) );
  XOR U39541 ( .A(n29476), .B(n26621), .Z(n29495) );
  IV U39542 ( .A(n29495), .Z(n32311) );
  IV U39543 ( .A(n26622), .Z(n26623) );
  NOR U39544 ( .A(n26624), .B(n26623), .Z(n32314) );
  IV U39545 ( .A(n26625), .Z(n26626) );
  NOR U39546 ( .A(n26627), .B(n26626), .Z(n32310) );
  NOR U39547 ( .A(n32314), .B(n32310), .Z(n29496) );
  IV U39548 ( .A(n29496), .Z(n29494) );
  XOR U39549 ( .A(n32311), .B(n29494), .Z(n29492) );
  XOR U39550 ( .A(n26628), .B(n29492), .Z(n29501) );
  XOR U39551 ( .A(n26629), .B(n29501), .Z(n29519) );
  XOR U39552 ( .A(n26630), .B(n29519), .Z(n28853) );
  IV U39553 ( .A(n26631), .Z(n26632) );
  NOR U39554 ( .A(n26633), .B(n26632), .Z(n28857) );
  IV U39555 ( .A(n26634), .Z(n26635) );
  NOR U39556 ( .A(n26636), .B(n26635), .Z(n28852) );
  NOR U39557 ( .A(n28857), .B(n28852), .Z(n26637) );
  XOR U39558 ( .A(n28853), .B(n26637), .Z(n29532) );
  XOR U39559 ( .A(n29523), .B(n29532), .Z(n28850) );
  XOR U39560 ( .A(n26638), .B(n28850), .Z(n28847) );
  XOR U39561 ( .A(n28848), .B(n28847), .Z(n29542) );
  XOR U39562 ( .A(n29539), .B(n29542), .Z(n28845) );
  XOR U39563 ( .A(n26639), .B(n28845), .Z(n28838) );
  XOR U39564 ( .A(n28839), .B(n28838), .Z(n28841) );
  XOR U39565 ( .A(n28840), .B(n28841), .Z(n26640) );
  NOR U39566 ( .A(n26641), .B(n26640), .Z(n35653) );
  IV U39567 ( .A(n26642), .Z(n26643) );
  NOR U39568 ( .A(n26644), .B(n26643), .Z(n28835) );
  NOR U39569 ( .A(n28840), .B(n28835), .Z(n26645) );
  XOR U39570 ( .A(n26645), .B(n28841), .Z(n28832) );
  NOR U39571 ( .A(n26646), .B(n28832), .Z(n26647) );
  NOR U39572 ( .A(n35653), .B(n26647), .Z(n28828) );
  IV U39573 ( .A(n26648), .Z(n26649) );
  NOR U39574 ( .A(n26650), .B(n26649), .Z(n28831) );
  IV U39575 ( .A(n26651), .Z(n26653) );
  NOR U39576 ( .A(n26653), .B(n26652), .Z(n28827) );
  NOR U39577 ( .A(n28831), .B(n28827), .Z(n26654) );
  XOR U39578 ( .A(n28828), .B(n26654), .Z(n28826) );
  IV U39579 ( .A(n26655), .Z(n26656) );
  NOR U39580 ( .A(n26657), .B(n26656), .Z(n28824) );
  IV U39581 ( .A(n26658), .Z(n26659) );
  NOR U39582 ( .A(n26660), .B(n26659), .Z(n28822) );
  NOR U39583 ( .A(n28824), .B(n28822), .Z(n26661) );
  XOR U39584 ( .A(n28826), .B(n26661), .Z(n29549) );
  XOR U39585 ( .A(n29550), .B(n29549), .Z(n32942) );
  XOR U39586 ( .A(n29547), .B(n32942), .Z(n26662) );
  IV U39587 ( .A(n26662), .Z(n28820) );
  XOR U39588 ( .A(n28819), .B(n28820), .Z(n26675) );
  IV U39589 ( .A(n26675), .Z(n26671) );
  IV U39590 ( .A(n26663), .Z(n26665) );
  NOR U39591 ( .A(n26665), .B(n26664), .Z(n26672) );
  IV U39592 ( .A(n26666), .Z(n26667) );
  NOR U39593 ( .A(n26668), .B(n26667), .Z(n26674) );
  NOR U39594 ( .A(n26672), .B(n26674), .Z(n26669) );
  IV U39595 ( .A(n26669), .Z(n26670) );
  NOR U39596 ( .A(n26671), .B(n26670), .Z(n26678) );
  IV U39597 ( .A(n26672), .Z(n26673) );
  NOR U39598 ( .A(n26673), .B(n28820), .Z(n32278) );
  IV U39599 ( .A(n26674), .Z(n26676) );
  NOR U39600 ( .A(n26676), .B(n26675), .Z(n32273) );
  NOR U39601 ( .A(n32278), .B(n32273), .Z(n26677) );
  IV U39602 ( .A(n26677), .Z(n28818) );
  NOR U39603 ( .A(n26678), .B(n28818), .Z(n28816) );
  IV U39604 ( .A(n26679), .Z(n26680) );
  NOR U39605 ( .A(n26681), .B(n26680), .Z(n28815) );
  IV U39606 ( .A(n26682), .Z(n26683) );
  NOR U39607 ( .A(n26684), .B(n26683), .Z(n29566) );
  NOR U39608 ( .A(n28815), .B(n29566), .Z(n26685) );
  XOR U39609 ( .A(n28816), .B(n26685), .Z(n29564) );
  IV U39610 ( .A(n26686), .Z(n26688) );
  NOR U39611 ( .A(n26688), .B(n26687), .Z(n28813) );
  IV U39612 ( .A(n26689), .Z(n26690) );
  NOR U39613 ( .A(n26691), .B(n26690), .Z(n29562) );
  NOR U39614 ( .A(n28813), .B(n29562), .Z(n26692) );
  XOR U39615 ( .A(n29564), .B(n26692), .Z(n28807) );
  IV U39616 ( .A(n26693), .Z(n26694) );
  NOR U39617 ( .A(n26695), .B(n26694), .Z(n28809) );
  IV U39618 ( .A(n26696), .Z(n26698) );
  NOR U39619 ( .A(n26698), .B(n26697), .Z(n28806) );
  NOR U39620 ( .A(n28809), .B(n28806), .Z(n26699) );
  XOR U39621 ( .A(n28807), .B(n26699), .Z(n35618) );
  IV U39622 ( .A(n26700), .Z(n26702) );
  NOR U39623 ( .A(n26702), .B(n26701), .Z(n35624) );
  IV U39624 ( .A(n26703), .Z(n26705) );
  NOR U39625 ( .A(n26705), .B(n26704), .Z(n35613) );
  NOR U39626 ( .A(n35624), .B(n35613), .Z(n29584) );
  XOR U39627 ( .A(n35618), .B(n29584), .Z(n29578) );
  IV U39628 ( .A(n26706), .Z(n26707) );
  NOR U39629 ( .A(n26708), .B(n26707), .Z(n29587) );
  IV U39630 ( .A(n26709), .Z(n26711) );
  NOR U39631 ( .A(n26711), .B(n26710), .Z(n29577) );
  NOR U39632 ( .A(n29587), .B(n29577), .Z(n26712) );
  XOR U39633 ( .A(n29578), .B(n26712), .Z(n29602) );
  XOR U39634 ( .A(n29581), .B(n29602), .Z(n29605) );
  XOR U39635 ( .A(n26713), .B(n29605), .Z(n29607) );
  XOR U39636 ( .A(n29608), .B(n29607), .Z(n29615) );
  XOR U39637 ( .A(n26714), .B(n29615), .Z(n26715) );
  IV U39638 ( .A(n26715), .Z(n29621) );
  IV U39639 ( .A(n26716), .Z(n26718) );
  NOR U39640 ( .A(n26718), .B(n26717), .Z(n29614) );
  IV U39641 ( .A(n26719), .Z(n26721) );
  NOR U39642 ( .A(n26721), .B(n26720), .Z(n29620) );
  NOR U39643 ( .A(n29614), .B(n29620), .Z(n26722) );
  XOR U39644 ( .A(n29621), .B(n26722), .Z(n29624) );
  IV U39645 ( .A(n29624), .Z(n32245) );
  IV U39646 ( .A(n26723), .Z(n26725) );
  NOR U39647 ( .A(n26725), .B(n26724), .Z(n32243) );
  IV U39648 ( .A(n26726), .Z(n26727) );
  NOR U39649 ( .A(n26728), .B(n26727), .Z(n32972) );
  NOR U39650 ( .A(n32243), .B(n32972), .Z(n29625) );
  IV U39651 ( .A(n29625), .Z(n29623) );
  XOR U39652 ( .A(n32245), .B(n29623), .Z(n32978) );
  XOR U39653 ( .A(n32976), .B(n32978), .Z(n28804) );
  IV U39654 ( .A(n26729), .Z(n26731) );
  NOR U39655 ( .A(n26731), .B(n26730), .Z(n32983) );
  IV U39656 ( .A(n26732), .Z(n26733) );
  NOR U39657 ( .A(n26734), .B(n26733), .Z(n28803) );
  NOR U39658 ( .A(n32983), .B(n28803), .Z(n26735) );
  XOR U39659 ( .A(n28804), .B(n26735), .Z(n29632) );
  IV U39660 ( .A(n26736), .Z(n26737) );
  NOR U39661 ( .A(n26738), .B(n26737), .Z(n39699) );
  IV U39662 ( .A(n26739), .Z(n26740) );
  NOR U39663 ( .A(n26741), .B(n26740), .Z(n39705) );
  NOR U39664 ( .A(n39699), .B(n39705), .Z(n32992) );
  XOR U39665 ( .A(n29632), .B(n32992), .Z(n29637) );
  IV U39666 ( .A(n26742), .Z(n26744) );
  NOR U39667 ( .A(n26744), .B(n26743), .Z(n29633) );
  IV U39668 ( .A(n26745), .Z(n26746) );
  NOR U39669 ( .A(n26747), .B(n26746), .Z(n29636) );
  NOR U39670 ( .A(n29633), .B(n29636), .Z(n26748) );
  XOR U39671 ( .A(n29637), .B(n26748), .Z(n29639) );
  XOR U39672 ( .A(n29640), .B(n29639), .Z(n29650) );
  IV U39673 ( .A(n26749), .Z(n26750) );
  NOR U39674 ( .A(n26751), .B(n26750), .Z(n29641) );
  IV U39675 ( .A(n26752), .Z(n26754) );
  NOR U39676 ( .A(n26754), .B(n26753), .Z(n29649) );
  NOR U39677 ( .A(n29641), .B(n29649), .Z(n26755) );
  XOR U39678 ( .A(n29650), .B(n26755), .Z(n29647) );
  XOR U39679 ( .A(n29648), .B(n29647), .Z(n28800) );
  XOR U39680 ( .A(n28801), .B(n28800), .Z(n26767) );
  IV U39681 ( .A(n26767), .Z(n26756) );
  NOR U39682 ( .A(n26757), .B(n26756), .Z(n33010) );
  IV U39683 ( .A(n26758), .Z(n26760) );
  NOR U39684 ( .A(n26760), .B(n26759), .Z(n26763) );
  IV U39685 ( .A(n26763), .Z(n26761) );
  NOR U39686 ( .A(n26761), .B(n28800), .Z(n33005) );
  NOR U39687 ( .A(n33010), .B(n33005), .Z(n26762) );
  IV U39688 ( .A(n26762), .Z(n33020) );
  NOR U39689 ( .A(n26764), .B(n26763), .Z(n26765) );
  IV U39690 ( .A(n26765), .Z(n26766) );
  NOR U39691 ( .A(n26767), .B(n26766), .Z(n26768) );
  NOR U39692 ( .A(n33020), .B(n26768), .Z(n29654) );
  IV U39693 ( .A(n26769), .Z(n26770) );
  NOR U39694 ( .A(n26771), .B(n26770), .Z(n33026) );
  IV U39695 ( .A(n26772), .Z(n26774) );
  NOR U39696 ( .A(n26774), .B(n26773), .Z(n33013) );
  NOR U39697 ( .A(n33026), .B(n33013), .Z(n29655) );
  XOR U39698 ( .A(n29654), .B(n29655), .Z(n33021) );
  XOR U39699 ( .A(n29658), .B(n33021), .Z(n29660) );
  IV U39700 ( .A(n26775), .Z(n26777) );
  NOR U39701 ( .A(n26777), .B(n26776), .Z(n29659) );
  IV U39702 ( .A(n26778), .Z(n26779) );
  NOR U39703 ( .A(n26780), .B(n26779), .Z(n29668) );
  NOR U39704 ( .A(n29659), .B(n29668), .Z(n26781) );
  XOR U39705 ( .A(n29660), .B(n26781), .Z(n29664) );
  XOR U39706 ( .A(n29663), .B(n29664), .Z(n28795) );
  XOR U39707 ( .A(n26782), .B(n28795), .Z(n28788) );
  XOR U39708 ( .A(n28789), .B(n28788), .Z(n28791) );
  XOR U39709 ( .A(n26783), .B(n28791), .Z(n28784) );
  XOR U39710 ( .A(n28785), .B(n28784), .Z(n29682) );
  XOR U39711 ( .A(n28782), .B(n29682), .Z(n26784) );
  NOR U39712 ( .A(n26785), .B(n26784), .Z(n33070) );
  IV U39713 ( .A(n26786), .Z(n26787) );
  NOR U39714 ( .A(n26788), .B(n26787), .Z(n29681) );
  NOR U39715 ( .A(n28782), .B(n29681), .Z(n26789) );
  XOR U39716 ( .A(n26789), .B(n29682), .Z(n29685) );
  NOR U39717 ( .A(n26790), .B(n29685), .Z(n26791) );
  NOR U39718 ( .A(n33070), .B(n26791), .Z(n29691) );
  IV U39719 ( .A(n26792), .Z(n26794) );
  NOR U39720 ( .A(n26794), .B(n26793), .Z(n29684) );
  IV U39721 ( .A(n26795), .Z(n26796) );
  NOR U39722 ( .A(n26797), .B(n26796), .Z(n29690) );
  NOR U39723 ( .A(n29684), .B(n29690), .Z(n26798) );
  XOR U39724 ( .A(n29691), .B(n26798), .Z(n28781) );
  IV U39725 ( .A(n26799), .Z(n26800) );
  NOR U39726 ( .A(n26801), .B(n26800), .Z(n28779) );
  IV U39727 ( .A(n26802), .Z(n26803) );
  NOR U39728 ( .A(n26804), .B(n26803), .Z(n28777) );
  NOR U39729 ( .A(n28779), .B(n28777), .Z(n26805) );
  XOR U39730 ( .A(n28781), .B(n26805), .Z(n28772) );
  IV U39731 ( .A(n26806), .Z(n26808) );
  NOR U39732 ( .A(n26808), .B(n26807), .Z(n28768) );
  IV U39733 ( .A(n26809), .Z(n26811) );
  NOR U39734 ( .A(n26811), .B(n26810), .Z(n28771) );
  NOR U39735 ( .A(n28768), .B(n28771), .Z(n26812) );
  XOR U39736 ( .A(n28772), .B(n26812), .Z(n29695) );
  XOR U39737 ( .A(n26813), .B(n29695), .Z(n28764) );
  XOR U39738 ( .A(n26814), .B(n28764), .Z(n28762) );
  NOR U39739 ( .A(n26815), .B(n28762), .Z(n32201) );
  IV U39740 ( .A(n26816), .Z(n26818) );
  NOR U39741 ( .A(n26818), .B(n26817), .Z(n28761) );
  XOR U39742 ( .A(n28761), .B(n28762), .Z(n33093) );
  IV U39743 ( .A(n33093), .Z(n26819) );
  NOR U39744 ( .A(n26820), .B(n26819), .Z(n28760) );
  NOR U39745 ( .A(n32201), .B(n28760), .Z(n28756) );
  XOR U39746 ( .A(n28757), .B(n28756), .Z(n35515) );
  XOR U39747 ( .A(n28755), .B(n35515), .Z(n32197) );
  XOR U39748 ( .A(n32198), .B(n32197), .Z(n32190) );
  IV U39749 ( .A(n26821), .Z(n26822) );
  NOR U39750 ( .A(n26823), .B(n26822), .Z(n32193) );
  IV U39751 ( .A(n26824), .Z(n26826) );
  NOR U39752 ( .A(n26826), .B(n26825), .Z(n32188) );
  NOR U39753 ( .A(n32193), .B(n32188), .Z(n26827) );
  IV U39754 ( .A(n26827), .Z(n28752) );
  XOR U39755 ( .A(n32190), .B(n28752), .Z(n29719) );
  XOR U39756 ( .A(n28748), .B(n29719), .Z(n26828) );
  NOR U39757 ( .A(n26829), .B(n26828), .Z(n32181) );
  IV U39758 ( .A(n26830), .Z(n26832) );
  NOR U39759 ( .A(n26832), .B(n26831), .Z(n29717) );
  NOR U39760 ( .A(n28748), .B(n29717), .Z(n26833) );
  XOR U39761 ( .A(n29719), .B(n26833), .Z(n29721) );
  NOR U39762 ( .A(n26834), .B(n29721), .Z(n26835) );
  NOR U39763 ( .A(n32181), .B(n26835), .Z(n28745) );
  IV U39764 ( .A(n26836), .Z(n26837) );
  NOR U39765 ( .A(n26838), .B(n26837), .Z(n29720) );
  IV U39766 ( .A(n26839), .Z(n26841) );
  NOR U39767 ( .A(n26841), .B(n26840), .Z(n28744) );
  NOR U39768 ( .A(n29720), .B(n28744), .Z(n26842) );
  XOR U39769 ( .A(n28745), .B(n26842), .Z(n29731) );
  IV U39770 ( .A(n26843), .Z(n26844) );
  NOR U39771 ( .A(n26845), .B(n26844), .Z(n29727) );
  IV U39772 ( .A(n26846), .Z(n26847) );
  NOR U39773 ( .A(n26848), .B(n26847), .Z(n29729) );
  NOR U39774 ( .A(n29727), .B(n29729), .Z(n26849) );
  XOR U39775 ( .A(n29731), .B(n26849), .Z(n28737) );
  IV U39776 ( .A(n26850), .Z(n26851) );
  NOR U39777 ( .A(n26852), .B(n26851), .Z(n28741) );
  IV U39778 ( .A(n26853), .Z(n26855) );
  NOR U39779 ( .A(n26855), .B(n26854), .Z(n28736) );
  NOR U39780 ( .A(n28741), .B(n28736), .Z(n26856) );
  XOR U39781 ( .A(n28737), .B(n26856), .Z(n29737) );
  IV U39782 ( .A(n26857), .Z(n26859) );
  NOR U39783 ( .A(n26859), .B(n26858), .Z(n33120) );
  IV U39784 ( .A(n26860), .Z(n26861) );
  NOR U39785 ( .A(n26862), .B(n26861), .Z(n32176) );
  NOR U39786 ( .A(n33120), .B(n32176), .Z(n29739) );
  XOR U39787 ( .A(n29737), .B(n29739), .Z(n28728) );
  IV U39788 ( .A(n26863), .Z(n26864) );
  NOR U39789 ( .A(n26865), .B(n26864), .Z(n28733) );
  IV U39790 ( .A(n26866), .Z(n26868) );
  NOR U39791 ( .A(n26868), .B(n26867), .Z(n28727) );
  NOR U39792 ( .A(n28733), .B(n28727), .Z(n26869) );
  XOR U39793 ( .A(n28728), .B(n26869), .Z(n28731) );
  XOR U39794 ( .A(n26870), .B(n28731), .Z(n26871) );
  IV U39795 ( .A(n26871), .Z(n29748) );
  XOR U39796 ( .A(n28723), .B(n29748), .Z(n29753) );
  IV U39797 ( .A(n26872), .Z(n26874) );
  NOR U39798 ( .A(n26874), .B(n26873), .Z(n29746) );
  IV U39799 ( .A(n26875), .Z(n26876) );
  NOR U39800 ( .A(n26877), .B(n26876), .Z(n29752) );
  NOR U39801 ( .A(n29746), .B(n29752), .Z(n26878) );
  XOR U39802 ( .A(n29753), .B(n26878), .Z(n28719) );
  IV U39803 ( .A(n26879), .Z(n26880) );
  NOR U39804 ( .A(n26881), .B(n26880), .Z(n29749) );
  IV U39805 ( .A(n26882), .Z(n26884) );
  NOR U39806 ( .A(n26884), .B(n26883), .Z(n28720) );
  NOR U39807 ( .A(n29749), .B(n28720), .Z(n26885) );
  XOR U39808 ( .A(n28719), .B(n26885), .Z(n32161) );
  IV U39809 ( .A(n26886), .Z(n26888) );
  NOR U39810 ( .A(n26888), .B(n26887), .Z(n32159) );
  IV U39811 ( .A(n26889), .Z(n26890) );
  NOR U39812 ( .A(n26891), .B(n26890), .Z(n33151) );
  NOR U39813 ( .A(n32159), .B(n33151), .Z(n28718) );
  XOR U39814 ( .A(n32161), .B(n28718), .Z(n28712) );
  XOR U39815 ( .A(n28716), .B(n28712), .Z(n28709) );
  XOR U39816 ( .A(n26892), .B(n28709), .Z(n28699) );
  XOR U39817 ( .A(n28700), .B(n28699), .Z(n28705) );
  XOR U39818 ( .A(n28701), .B(n28705), .Z(n28697) );
  IV U39819 ( .A(n26893), .Z(n26895) );
  NOR U39820 ( .A(n26895), .B(n26894), .Z(n28704) );
  IV U39821 ( .A(n26896), .Z(n26897) );
  NOR U39822 ( .A(n26898), .B(n26897), .Z(n28696) );
  NOR U39823 ( .A(n28704), .B(n28696), .Z(n26899) );
  XOR U39824 ( .A(n28697), .B(n26899), .Z(n28688) );
  XOR U39825 ( .A(n26900), .B(n28688), .Z(n29765) );
  XOR U39826 ( .A(n26901), .B(n29765), .Z(n29762) );
  XOR U39827 ( .A(n29763), .B(n29762), .Z(n32134) );
  XOR U39828 ( .A(n29773), .B(n32134), .Z(n29770) );
  IV U39829 ( .A(n26902), .Z(n26903) );
  NOR U39830 ( .A(n26904), .B(n26903), .Z(n29769) );
  IV U39831 ( .A(n26905), .Z(n26907) );
  NOR U39832 ( .A(n26907), .B(n26906), .Z(n29778) );
  NOR U39833 ( .A(n29769), .B(n29778), .Z(n26908) );
  XOR U39834 ( .A(n29770), .B(n26908), .Z(n29782) );
  XOR U39835 ( .A(n29781), .B(n29782), .Z(n28684) );
  XOR U39836 ( .A(n26909), .B(n28684), .Z(n28678) );
  XOR U39837 ( .A(n28679), .B(n28678), .Z(n28676) );
  XOR U39838 ( .A(n28675), .B(n28676), .Z(n26910) );
  NOR U39839 ( .A(n26911), .B(n26910), .Z(n32119) );
  IV U39840 ( .A(n26912), .Z(n26914) );
  NOR U39841 ( .A(n26914), .B(n26913), .Z(n28673) );
  NOR U39842 ( .A(n28675), .B(n28673), .Z(n26915) );
  XOR U39843 ( .A(n26915), .B(n28676), .Z(n28670) );
  NOR U39844 ( .A(n26916), .B(n28670), .Z(n26917) );
  NOR U39845 ( .A(n32119), .B(n26917), .Z(n29787) );
  IV U39846 ( .A(n26918), .Z(n26920) );
  NOR U39847 ( .A(n26920), .B(n26919), .Z(n28669) );
  IV U39848 ( .A(n26921), .Z(n26923) );
  NOR U39849 ( .A(n26923), .B(n26922), .Z(n29786) );
  NOR U39850 ( .A(n28669), .B(n29786), .Z(n26924) );
  XOR U39851 ( .A(n29787), .B(n26924), .Z(n29797) );
  IV U39852 ( .A(n26925), .Z(n26927) );
  NOR U39853 ( .A(n26927), .B(n26926), .Z(n29790) );
  IV U39854 ( .A(n26928), .Z(n26929) );
  NOR U39855 ( .A(n26930), .B(n26929), .Z(n29795) );
  NOR U39856 ( .A(n29790), .B(n29795), .Z(n26931) );
  XOR U39857 ( .A(n29797), .B(n26931), .Z(n28667) );
  IV U39858 ( .A(n26932), .Z(n26934) );
  NOR U39859 ( .A(n26934), .B(n26933), .Z(n29792) );
  IV U39860 ( .A(n26935), .Z(n26936) );
  NOR U39861 ( .A(n26937), .B(n26936), .Z(n28666) );
  NOR U39862 ( .A(n29792), .B(n28666), .Z(n26938) );
  XOR U39863 ( .A(n28667), .B(n26938), .Z(n28664) );
  XOR U39864 ( .A(n26939), .B(n28664), .Z(n26940) );
  IV U39865 ( .A(n26940), .Z(n28657) );
  XOR U39866 ( .A(n28654), .B(n28657), .Z(n28652) );
  IV U39867 ( .A(n26941), .Z(n26942) );
  NOR U39868 ( .A(n26943), .B(n26942), .Z(n28656) );
  IV U39869 ( .A(n26944), .Z(n26945) );
  NOR U39870 ( .A(n26946), .B(n26945), .Z(n28651) );
  NOR U39871 ( .A(n28656), .B(n28651), .Z(n26947) );
  XOR U39872 ( .A(n28652), .B(n26947), .Z(n29804) );
  IV U39873 ( .A(n26948), .Z(n26950) );
  NOR U39874 ( .A(n26950), .B(n26949), .Z(n32098) );
  IV U39875 ( .A(n26951), .Z(n26953) );
  NOR U39876 ( .A(n26953), .B(n26952), .Z(n32091) );
  NOR U39877 ( .A(n32098), .B(n32091), .Z(n29805) );
  XOR U39878 ( .A(n29804), .B(n29805), .Z(n29807) );
  XOR U39879 ( .A(n29806), .B(n29807), .Z(n29817) );
  IV U39880 ( .A(n26954), .Z(n26955) );
  NOR U39881 ( .A(n26956), .B(n26955), .Z(n29802) );
  IV U39882 ( .A(n26957), .Z(n26958) );
  NOR U39883 ( .A(n26959), .B(n26958), .Z(n29816) );
  NOR U39884 ( .A(n29802), .B(n29816), .Z(n26960) );
  XOR U39885 ( .A(n29817), .B(n26960), .Z(n29813) );
  IV U39886 ( .A(n26961), .Z(n26963) );
  NOR U39887 ( .A(n26963), .B(n26962), .Z(n29814) );
  IV U39888 ( .A(n26964), .Z(n26966) );
  NOR U39889 ( .A(n26966), .B(n26965), .Z(n29820) );
  NOR U39890 ( .A(n29814), .B(n29820), .Z(n26967) );
  XOR U39891 ( .A(n29813), .B(n26967), .Z(n29824) );
  XOR U39892 ( .A(n29823), .B(n29824), .Z(n28647) );
  IV U39893 ( .A(n26968), .Z(n26969) );
  NOR U39894 ( .A(n26970), .B(n26969), .Z(n28649) );
  IV U39895 ( .A(n26971), .Z(n26973) );
  NOR U39896 ( .A(n26973), .B(n26972), .Z(n28646) );
  NOR U39897 ( .A(n28649), .B(n28646), .Z(n26974) );
  XOR U39898 ( .A(n28647), .B(n26974), .Z(n29837) );
  IV U39899 ( .A(n26975), .Z(n26976) );
  NOR U39900 ( .A(n26977), .B(n26976), .Z(n29831) );
  IV U39901 ( .A(n26978), .Z(n26979) );
  NOR U39902 ( .A(n26980), .B(n26979), .Z(n29833) );
  NOR U39903 ( .A(n29831), .B(n29833), .Z(n26981) );
  XOR U39904 ( .A(n29837), .B(n26981), .Z(n29844) );
  IV U39905 ( .A(n26982), .Z(n26984) );
  NOR U39906 ( .A(n26984), .B(n26983), .Z(n29836) );
  IV U39907 ( .A(n26985), .Z(n26987) );
  NOR U39908 ( .A(n26987), .B(n26986), .Z(n29843) );
  NOR U39909 ( .A(n29836), .B(n29843), .Z(n26988) );
  XOR U39910 ( .A(n29844), .B(n26988), .Z(n29847) );
  IV U39911 ( .A(n26989), .Z(n26991) );
  NOR U39912 ( .A(n26991), .B(n26990), .Z(n29848) );
  IV U39913 ( .A(n26992), .Z(n26993) );
  NOR U39914 ( .A(n26994), .B(n26993), .Z(n29850) );
  NOR U39915 ( .A(n29848), .B(n29850), .Z(n26995) );
  XOR U39916 ( .A(n29847), .B(n26995), .Z(n32065) );
  IV U39917 ( .A(n26996), .Z(n26997) );
  NOR U39918 ( .A(n26998), .B(n26997), .Z(n32064) );
  IV U39919 ( .A(n26999), .Z(n27000) );
  NOR U39920 ( .A(n27001), .B(n27000), .Z(n33246) );
  NOR U39921 ( .A(n32064), .B(n33246), .Z(n29846) );
  IV U39922 ( .A(n29846), .Z(n29865) );
  XOR U39923 ( .A(n32065), .B(n29865), .Z(n29860) );
  XOR U39924 ( .A(n29861), .B(n29860), .Z(n27002) );
  IV U39925 ( .A(n27002), .Z(n29856) );
  XOR U39926 ( .A(n29855), .B(n29856), .Z(n27009) );
  IV U39927 ( .A(n27009), .Z(n27003) );
  NOR U39928 ( .A(n27008), .B(n27003), .Z(n27004) );
  IV U39929 ( .A(n27004), .Z(n27005) );
  NOR U39930 ( .A(n27006), .B(n27005), .Z(n33276) );
  IV U39931 ( .A(n27006), .Z(n27007) );
  NOR U39932 ( .A(n27007), .B(n29856), .Z(n33257) );
  IV U39933 ( .A(n27008), .Z(n27010) );
  NOR U39934 ( .A(n27010), .B(n27009), .Z(n33261) );
  NOR U39935 ( .A(n33257), .B(n33261), .Z(n27011) );
  IV U39936 ( .A(n27011), .Z(n33269) );
  NOR U39937 ( .A(n33276), .B(n33269), .Z(n29884) );
  IV U39938 ( .A(n27012), .Z(n27013) );
  NOR U39939 ( .A(n27014), .B(n27013), .Z(n33267) );
  IV U39940 ( .A(n27015), .Z(n27017) );
  NOR U39941 ( .A(n27017), .B(n27016), .Z(n33279) );
  NOR U39942 ( .A(n33267), .B(n33279), .Z(n29886) );
  XOR U39943 ( .A(n29884), .B(n29886), .Z(n32052) );
  IV U39944 ( .A(n27018), .Z(n27020) );
  NOR U39945 ( .A(n27020), .B(n27019), .Z(n32056) );
  IV U39946 ( .A(n27021), .Z(n27022) );
  NOR U39947 ( .A(n27023), .B(n27022), .Z(n32050) );
  NOR U39948 ( .A(n32056), .B(n32050), .Z(n29888) );
  XOR U39949 ( .A(n32052), .B(n29888), .Z(n29889) );
  XOR U39950 ( .A(n29890), .B(n29889), .Z(n32034) );
  IV U39951 ( .A(n27024), .Z(n27026) );
  NOR U39952 ( .A(n27026), .B(n27025), .Z(n32041) );
  IV U39953 ( .A(n27027), .Z(n27028) );
  NOR U39954 ( .A(n27029), .B(n27028), .Z(n32032) );
  NOR U39955 ( .A(n32041), .B(n32032), .Z(n29894) );
  XOR U39956 ( .A(n32034), .B(n29894), .Z(n29896) );
  XOR U39957 ( .A(n29899), .B(n29896), .Z(n27030) );
  NOR U39958 ( .A(n27031), .B(n27030), .Z(n33289) );
  IV U39959 ( .A(n27032), .Z(n27034) );
  NOR U39960 ( .A(n27034), .B(n27033), .Z(n29895) );
  NOR U39961 ( .A(n27035), .B(n29895), .Z(n27036) );
  XOR U39962 ( .A(n27036), .B(n29896), .Z(n33293) );
  IV U39963 ( .A(n33293), .Z(n27037) );
  NOR U39964 ( .A(n27038), .B(n27037), .Z(n27039) );
  NOR U39965 ( .A(n33289), .B(n27039), .Z(n29903) );
  IV U39966 ( .A(n27040), .Z(n27042) );
  NOR U39967 ( .A(n27042), .B(n27041), .Z(n33291) );
  IV U39968 ( .A(n27043), .Z(n27044) );
  NOR U39969 ( .A(n27045), .B(n27044), .Z(n33298) );
  NOR U39970 ( .A(n33291), .B(n33298), .Z(n29904) );
  XOR U39971 ( .A(n29903), .B(n29904), .Z(n29914) );
  XOR U39972 ( .A(n27046), .B(n29914), .Z(n27047) );
  IV U39973 ( .A(n27047), .Z(n29917) );
  XOR U39974 ( .A(n29916), .B(n29917), .Z(n28642) );
  IV U39975 ( .A(n27048), .Z(n27049) );
  NOR U39976 ( .A(n27050), .B(n27049), .Z(n29910) );
  IV U39977 ( .A(n27051), .Z(n28645) );
  NOR U39978 ( .A(n28645), .B(n28643), .Z(n27052) );
  NOR U39979 ( .A(n29910), .B(n27052), .Z(n27053) );
  XOR U39980 ( .A(n28642), .B(n27053), .Z(n28639) );
  IV U39981 ( .A(n27054), .Z(n27056) );
  NOR U39982 ( .A(n27056), .B(n27055), .Z(n28640) );
  IV U39983 ( .A(n27057), .Z(n27059) );
  NOR U39984 ( .A(n27059), .B(n27058), .Z(n29927) );
  NOR U39985 ( .A(n28640), .B(n29927), .Z(n27060) );
  XOR U39986 ( .A(n28639), .B(n27060), .Z(n29934) );
  IV U39987 ( .A(n27061), .Z(n27063) );
  NOR U39988 ( .A(n27063), .B(n27062), .Z(n29933) );
  IV U39989 ( .A(n27064), .Z(n27065) );
  NOR U39990 ( .A(n27066), .B(n27065), .Z(n29924) );
  NOR U39991 ( .A(n29933), .B(n29924), .Z(n27067) );
  XOR U39992 ( .A(n29934), .B(n27067), .Z(n29936) );
  XOR U39993 ( .A(n29937), .B(n29936), .Z(n28637) );
  XOR U39994 ( .A(n28634), .B(n28637), .Z(n29946) );
  IV U39995 ( .A(n27068), .Z(n27069) );
  NOR U39996 ( .A(n27070), .B(n27069), .Z(n28636) );
  IV U39997 ( .A(n27071), .Z(n27073) );
  NOR U39998 ( .A(n27073), .B(n27072), .Z(n29945) );
  NOR U39999 ( .A(n28636), .B(n29945), .Z(n27074) );
  XOR U40000 ( .A(n29946), .B(n27074), .Z(n28632) );
  IV U40001 ( .A(n27075), .Z(n27076) );
  NOR U40002 ( .A(n27077), .B(n27076), .Z(n36699) );
  IV U40003 ( .A(n27078), .Z(n27079) );
  NOR U40004 ( .A(n27080), .B(n27079), .Z(n36709) );
  NOR U40005 ( .A(n36699), .B(n36709), .Z(n28633) );
  XOR U40006 ( .A(n28632), .B(n28633), .Z(n29957) );
  IV U40007 ( .A(n27081), .Z(n27083) );
  NOR U40008 ( .A(n27083), .B(n27082), .Z(n29956) );
  IV U40009 ( .A(n27084), .Z(n27086) );
  NOR U40010 ( .A(n27086), .B(n27085), .Z(n29953) );
  NOR U40011 ( .A(n29956), .B(n29953), .Z(n27087) );
  XOR U40012 ( .A(n29957), .B(n27087), .Z(n28626) );
  IV U40013 ( .A(n27088), .Z(n27090) );
  NOR U40014 ( .A(n27090), .B(n27089), .Z(n28629) );
  IV U40015 ( .A(n27091), .Z(n27092) );
  NOR U40016 ( .A(n27093), .B(n27092), .Z(n28627) );
  NOR U40017 ( .A(n28629), .B(n28627), .Z(n27094) );
  XOR U40018 ( .A(n28626), .B(n27094), .Z(n31999) );
  XOR U40019 ( .A(n29967), .B(n31999), .Z(n28624) );
  XOR U40020 ( .A(n27095), .B(n28624), .Z(n29979) );
  IV U40021 ( .A(n27096), .Z(n27098) );
  NOR U40022 ( .A(n27098), .B(n27097), .Z(n29980) );
  IV U40023 ( .A(n27099), .Z(n27101) );
  NOR U40024 ( .A(n27101), .B(n27100), .Z(n28620) );
  NOR U40025 ( .A(n29980), .B(n28620), .Z(n27102) );
  XOR U40026 ( .A(n29979), .B(n27102), .Z(n29988) );
  XOR U40027 ( .A(n27103), .B(n29988), .Z(n35340) );
  XOR U40028 ( .A(n29992), .B(n35340), .Z(n28617) );
  XOR U40029 ( .A(n27104), .B(n28617), .Z(n30009) );
  IV U40030 ( .A(n30009), .Z(n27112) );
  IV U40031 ( .A(n27105), .Z(n27107) );
  NOR U40032 ( .A(n27107), .B(n27106), .Z(n30005) );
  IV U40033 ( .A(n27108), .Z(n27110) );
  NOR U40034 ( .A(n27110), .B(n27109), .Z(n30008) );
  NOR U40035 ( .A(n30005), .B(n30008), .Z(n27111) );
  XOR U40036 ( .A(n27112), .B(n27111), .Z(n31976) );
  XOR U40037 ( .A(n31978), .B(n31976), .Z(n30014) );
  IV U40038 ( .A(n27113), .Z(n27114) );
  NOR U40039 ( .A(n27115), .B(n27114), .Z(n36737) );
  IV U40040 ( .A(n27116), .Z(n27118) );
  NOR U40041 ( .A(n27118), .B(n27117), .Z(n35317) );
  NOR U40042 ( .A(n36737), .B(n35317), .Z(n30015) );
  XOR U40043 ( .A(n30014), .B(n30015), .Z(n30021) );
  XOR U40044 ( .A(n27119), .B(n30021), .Z(n30030) );
  IV U40045 ( .A(n27120), .Z(n27122) );
  NOR U40046 ( .A(n27122), .B(n27121), .Z(n30020) );
  IV U40047 ( .A(n27123), .Z(n27125) );
  NOR U40048 ( .A(n27125), .B(n27124), .Z(n30029) );
  NOR U40049 ( .A(n30020), .B(n30029), .Z(n27126) );
  XOR U40050 ( .A(n30030), .B(n27126), .Z(n30028) );
  XOR U40051 ( .A(n30026), .B(n30028), .Z(n27133) );
  NOR U40052 ( .A(n27127), .B(n27133), .Z(n31965) );
  IV U40053 ( .A(n27128), .Z(n27129) );
  NOR U40054 ( .A(n27130), .B(n27129), .Z(n27135) );
  IV U40055 ( .A(n27135), .Z(n27131) );
  NOR U40056 ( .A(n30028), .B(n27131), .Z(n31968) );
  NOR U40057 ( .A(n31965), .B(n31968), .Z(n27132) );
  IV U40058 ( .A(n27132), .Z(n30035) );
  NOR U40059 ( .A(n30035), .B(n27133), .Z(n27138) );
  NOR U40060 ( .A(n27135), .B(n27134), .Z(n27136) );
  NOR U40061 ( .A(n27136), .B(n30035), .Z(n27137) );
  NOR U40062 ( .A(n27138), .B(n27137), .Z(n31959) );
  XOR U40063 ( .A(n30036), .B(n31959), .Z(n30038) );
  IV U40064 ( .A(n27139), .Z(n27140) );
  NOR U40065 ( .A(n27141), .B(n27140), .Z(n30037) );
  IV U40066 ( .A(n27142), .Z(n27143) );
  NOR U40067 ( .A(n27144), .B(n27143), .Z(n30044) );
  NOR U40068 ( .A(n30037), .B(n30044), .Z(n27145) );
  XOR U40069 ( .A(n30038), .B(n27145), .Z(n30048) );
  XOR U40070 ( .A(n30047), .B(n30048), .Z(n30054) );
  XOR U40071 ( .A(n27146), .B(n30054), .Z(n30056) );
  XOR U40072 ( .A(n30057), .B(n30056), .Z(n31948) );
  XOR U40073 ( .A(n30058), .B(n31948), .Z(n28612) );
  IV U40074 ( .A(n27147), .Z(n27149) );
  NOR U40075 ( .A(n27149), .B(n27148), .Z(n30062) );
  IV U40076 ( .A(n27150), .Z(n27152) );
  NOR U40077 ( .A(n27152), .B(n27151), .Z(n28611) );
  NOR U40078 ( .A(n30062), .B(n28611), .Z(n27153) );
  XOR U40079 ( .A(n28612), .B(n27153), .Z(n35288) );
  IV U40080 ( .A(n27154), .Z(n27156) );
  NOR U40081 ( .A(n27156), .B(n27155), .Z(n35291) );
  IV U40082 ( .A(n27157), .Z(n27158) );
  NOR U40083 ( .A(n27159), .B(n27158), .Z(n35283) );
  NOR U40084 ( .A(n35291), .B(n35283), .Z(n28608) );
  XOR U40085 ( .A(n35288), .B(n28608), .Z(n28609) );
  IV U40086 ( .A(n27160), .Z(n27161) );
  NOR U40087 ( .A(n27162), .B(n27161), .Z(n35278) );
  IV U40088 ( .A(n27163), .Z(n27165) );
  NOR U40089 ( .A(n27165), .B(n27164), .Z(n36797) );
  NOR U40090 ( .A(n35278), .B(n36797), .Z(n31940) );
  XOR U40091 ( .A(n28609), .B(n31940), .Z(n28605) );
  XOR U40092 ( .A(n28604), .B(n28605), .Z(n27166) );
  NOR U40093 ( .A(n27175), .B(n27166), .Z(n31930) );
  IV U40094 ( .A(n27167), .Z(n27169) );
  NOR U40095 ( .A(n27169), .B(n27168), .Z(n27170) );
  IV U40096 ( .A(n27170), .Z(n28600) );
  IV U40097 ( .A(n27171), .Z(n27172) );
  NOR U40098 ( .A(n27173), .B(n27172), .Z(n28601) );
  NOR U40099 ( .A(n28604), .B(n28601), .Z(n27174) );
  XOR U40100 ( .A(n27174), .B(n28605), .Z(n27176) );
  IV U40101 ( .A(n27176), .Z(n28599) );
  XOR U40102 ( .A(n28600), .B(n28599), .Z(n27178) );
  NOR U40103 ( .A(n27176), .B(n27175), .Z(n27177) );
  NOR U40104 ( .A(n27178), .B(n27177), .Z(n27179) );
  NOR U40105 ( .A(n31930), .B(n27179), .Z(n28597) );
  XOR U40106 ( .A(n28598), .B(n28597), .Z(n33394) );
  XOR U40107 ( .A(n30069), .B(n33394), .Z(n30080) );
  IV U40108 ( .A(n27180), .Z(n27181) );
  NOR U40109 ( .A(n27182), .B(n27181), .Z(n28596) );
  IV U40110 ( .A(n27183), .Z(n27184) );
  NOR U40111 ( .A(n27185), .B(n27184), .Z(n30076) );
  NOR U40112 ( .A(n28596), .B(n30076), .Z(n27186) );
  XOR U40113 ( .A(n30080), .B(n27186), .Z(n30087) );
  XOR U40114 ( .A(n27187), .B(n30087), .Z(n27188) );
  IV U40115 ( .A(n27188), .Z(n31910) );
  XOR U40116 ( .A(n30090), .B(n31910), .Z(n33419) );
  XOR U40117 ( .A(n28595), .B(n33419), .Z(n31905) );
  XOR U40118 ( .A(n30096), .B(n31905), .Z(n28592) );
  IV U40119 ( .A(n27189), .Z(n27190) );
  NOR U40120 ( .A(n27191), .B(n27190), .Z(n36824) );
  IV U40121 ( .A(n27192), .Z(n27194) );
  NOR U40122 ( .A(n27194), .B(n27193), .Z(n36831) );
  NOR U40123 ( .A(n36824), .B(n36831), .Z(n28593) );
  XOR U40124 ( .A(n28592), .B(n28593), .Z(n30111) );
  XOR U40125 ( .A(n30110), .B(n30111), .Z(n28590) );
  XOR U40126 ( .A(n27195), .B(n28590), .Z(n30121) );
  XOR U40127 ( .A(n30122), .B(n30121), .Z(n30124) );
  NOR U40128 ( .A(n27203), .B(n30124), .Z(n31889) );
  IV U40129 ( .A(n27196), .Z(n27197) );
  NOR U40130 ( .A(n27198), .B(n27197), .Z(n27199) );
  IV U40131 ( .A(n27199), .Z(n28588) );
  IV U40132 ( .A(n27200), .Z(n27201) );
  NOR U40133 ( .A(n27202), .B(n27201), .Z(n30123) );
  XOR U40134 ( .A(n30123), .B(n30124), .Z(n28587) );
  XOR U40135 ( .A(n28588), .B(n28587), .Z(n27206) );
  IV U40136 ( .A(n28587), .Z(n27204) );
  NOR U40137 ( .A(n27204), .B(n27203), .Z(n27205) );
  NOR U40138 ( .A(n27206), .B(n27205), .Z(n27207) );
  NOR U40139 ( .A(n31889), .B(n27207), .Z(n30133) );
  XOR U40140 ( .A(n27208), .B(n30133), .Z(n30145) );
  XOR U40141 ( .A(n27209), .B(n30145), .Z(n28585) );
  XOR U40142 ( .A(n28586), .B(n28585), .Z(n33461) );
  XOR U40143 ( .A(n28581), .B(n33461), .Z(n28582) );
  XOR U40144 ( .A(n31879), .B(n28582), .Z(n28579) );
  IV U40145 ( .A(n27210), .Z(n27211) );
  NOR U40146 ( .A(n27212), .B(n27211), .Z(n28578) );
  IV U40147 ( .A(n27213), .Z(n27215) );
  NOR U40148 ( .A(n27215), .B(n27214), .Z(n28576) );
  NOR U40149 ( .A(n28578), .B(n28576), .Z(n27216) );
  XOR U40150 ( .A(n28579), .B(n27216), .Z(n27224) );
  IV U40151 ( .A(n27224), .Z(n27217) );
  NOR U40152 ( .A(n27218), .B(n27217), .Z(n33474) );
  IV U40153 ( .A(n27219), .Z(n27221) );
  NOR U40154 ( .A(n27221), .B(n27220), .Z(n27225) );
  IV U40155 ( .A(n27225), .Z(n27223) );
  XOR U40156 ( .A(n28578), .B(n28579), .Z(n27222) );
  NOR U40157 ( .A(n27223), .B(n27222), .Z(n33471) );
  NOR U40158 ( .A(n27225), .B(n27224), .Z(n27226) );
  NOR U40159 ( .A(n33471), .B(n27226), .Z(n27227) );
  NOR U40160 ( .A(n31871), .B(n27227), .Z(n27228) );
  NOR U40161 ( .A(n33474), .B(n27228), .Z(n28571) );
  XOR U40162 ( .A(n28574), .B(n28571), .Z(n30155) );
  XOR U40163 ( .A(n27229), .B(n30155), .Z(n27230) );
  IV U40164 ( .A(n27230), .Z(n30160) );
  XOR U40165 ( .A(n27231), .B(n30160), .Z(n33483) );
  XOR U40166 ( .A(n33484), .B(n33483), .Z(n31857) );
  XOR U40167 ( .A(n28567), .B(n31857), .Z(n31849) );
  XOR U40168 ( .A(n28562), .B(n31849), .Z(n28563) );
  XOR U40169 ( .A(n28564), .B(n28563), .Z(n33502) );
  XOR U40170 ( .A(n28558), .B(n33502), .Z(n33510) );
  XOR U40171 ( .A(n28560), .B(n33510), .Z(n28556) );
  XOR U40172 ( .A(n28557), .B(n28556), .Z(n33526) );
  XOR U40173 ( .A(n28552), .B(n33526), .Z(n28554) );
  XOR U40174 ( .A(n27232), .B(n28554), .Z(n28551) );
  XOR U40175 ( .A(n28547), .B(n28551), .Z(n28545) );
  IV U40176 ( .A(n27233), .Z(n27235) );
  NOR U40177 ( .A(n27235), .B(n27234), .Z(n28549) );
  IV U40178 ( .A(n27236), .Z(n27237) );
  NOR U40179 ( .A(n27238), .B(n27237), .Z(n28544) );
  NOR U40180 ( .A(n28549), .B(n28544), .Z(n27239) );
  XOR U40181 ( .A(n28545), .B(n27239), .Z(n28541) );
  IV U40182 ( .A(n27240), .Z(n27241) );
  NOR U40183 ( .A(n27242), .B(n27241), .Z(n28542) );
  IV U40184 ( .A(n27243), .Z(n27244) );
  NOR U40185 ( .A(n27245), .B(n27244), .Z(n30172) );
  NOR U40186 ( .A(n28542), .B(n30172), .Z(n27246) );
  XOR U40187 ( .A(n28541), .B(n27246), .Z(n31813) );
  XOR U40188 ( .A(n30175), .B(n31813), .Z(n28539) );
  XOR U40189 ( .A(n28540), .B(n28539), .Z(n30178) );
  XOR U40190 ( .A(n30179), .B(n30178), .Z(n30181) );
  IV U40191 ( .A(n27247), .Z(n27248) );
  NOR U40192 ( .A(n27249), .B(n27248), .Z(n30180) );
  IV U40193 ( .A(n27250), .Z(n27251) );
  NOR U40194 ( .A(n27252), .B(n27251), .Z(n33563) );
  NOR U40195 ( .A(n30180), .B(n33563), .Z(n27253) );
  XOR U40196 ( .A(n30181), .B(n27253), .Z(n27254) );
  IV U40197 ( .A(n27254), .Z(n28536) );
  XOR U40198 ( .A(n28535), .B(n28536), .Z(n27255) );
  NOR U40199 ( .A(n27256), .B(n27255), .Z(n30190) );
  IV U40200 ( .A(n27257), .Z(n27259) );
  NOR U40201 ( .A(n27259), .B(n27258), .Z(n28532) );
  NOR U40202 ( .A(n28535), .B(n28532), .Z(n27260) );
  XOR U40203 ( .A(n27260), .B(n28536), .Z(n30195) );
  NOR U40204 ( .A(n27261), .B(n30195), .Z(n27262) );
  NOR U40205 ( .A(n30190), .B(n27262), .Z(n27263) );
  IV U40206 ( .A(n27263), .Z(n30188) );
  XOR U40207 ( .A(n30189), .B(n30188), .Z(n28529) );
  IV U40208 ( .A(n27264), .Z(n27266) );
  NOR U40209 ( .A(n27266), .B(n27265), .Z(n28528) );
  IV U40210 ( .A(n27267), .Z(n27268) );
  NOR U40211 ( .A(n27269), .B(n27268), .Z(n30208) );
  NOR U40212 ( .A(n28528), .B(n30208), .Z(n27270) );
  XOR U40213 ( .A(n28529), .B(n27270), .Z(n35158) );
  XOR U40214 ( .A(n30207), .B(n35158), .Z(n30214) );
  IV U40215 ( .A(n27271), .Z(n27273) );
  NOR U40216 ( .A(n27273), .B(n27272), .Z(n30217) );
  IV U40217 ( .A(n27274), .Z(n27276) );
  NOR U40218 ( .A(n27276), .B(n27275), .Z(n30213) );
  NOR U40219 ( .A(n30217), .B(n30213), .Z(n27277) );
  XOR U40220 ( .A(n30214), .B(n27277), .Z(n30232) );
  XOR U40221 ( .A(n27278), .B(n30232), .Z(n30236) );
  IV U40222 ( .A(n27279), .Z(n27281) );
  NOR U40223 ( .A(n27281), .B(n27280), .Z(n30240) );
  IV U40224 ( .A(n27282), .Z(n27283) );
  NOR U40225 ( .A(n27284), .B(n27283), .Z(n30245) );
  NOR U40226 ( .A(n30240), .B(n30245), .Z(n30237) );
  XOR U40227 ( .A(n30236), .B(n30237), .Z(n28524) );
  NOR U40228 ( .A(n27292), .B(n28524), .Z(n30263) );
  IV U40229 ( .A(n27285), .Z(n27287) );
  NOR U40230 ( .A(n27287), .B(n27286), .Z(n27288) );
  IV U40231 ( .A(n27288), .Z(n30259) );
  IV U40232 ( .A(n27289), .Z(n27290) );
  NOR U40233 ( .A(n27291), .B(n27290), .Z(n28523) );
  XOR U40234 ( .A(n28523), .B(n28524), .Z(n30258) );
  XOR U40235 ( .A(n30259), .B(n30258), .Z(n27295) );
  IV U40236 ( .A(n30258), .Z(n27293) );
  NOR U40237 ( .A(n27293), .B(n27292), .Z(n27294) );
  NOR U40238 ( .A(n27295), .B(n27294), .Z(n27296) );
  NOR U40239 ( .A(n30263), .B(n27296), .Z(n30255) );
  XOR U40240 ( .A(n27297), .B(n30255), .Z(n31792) );
  XOR U40241 ( .A(n28518), .B(n31792), .Z(n28519) );
  XOR U40242 ( .A(n28520), .B(n28519), .Z(n28514) );
  XOR U40243 ( .A(n28513), .B(n28514), .Z(n31786) );
  XOR U40244 ( .A(n28516), .B(n31786), .Z(n28509) );
  XOR U40245 ( .A(n31784), .B(n28509), .Z(n31775) );
  XOR U40246 ( .A(n28510), .B(n31775), .Z(n28503) );
  XOR U40247 ( .A(n28504), .B(n28503), .Z(n28506) );
  IV U40248 ( .A(n27298), .Z(n27300) );
  NOR U40249 ( .A(n27300), .B(n27299), .Z(n28505) );
  IV U40250 ( .A(n27301), .Z(n27303) );
  NOR U40251 ( .A(n27303), .B(n27302), .Z(n28500) );
  NOR U40252 ( .A(n28505), .B(n28500), .Z(n27304) );
  XOR U40253 ( .A(n28506), .B(n27304), .Z(n27312) );
  IV U40254 ( .A(n27312), .Z(n27305) );
  NOR U40255 ( .A(n27306), .B(n27305), .Z(n31765) );
  IV U40256 ( .A(n27307), .Z(n27308) );
  NOR U40257 ( .A(n27309), .B(n27308), .Z(n27313) );
  IV U40258 ( .A(n27313), .Z(n27311) );
  XOR U40259 ( .A(n28505), .B(n28506), .Z(n27310) );
  NOR U40260 ( .A(n27311), .B(n27310), .Z(n33617) );
  NOR U40261 ( .A(n27313), .B(n27312), .Z(n27314) );
  NOR U40262 ( .A(n33617), .B(n27314), .Z(n28497) );
  NOR U40263 ( .A(n27315), .B(n28497), .Z(n27316) );
  NOR U40264 ( .A(n31765), .B(n27316), .Z(n28493) );
  XOR U40265 ( .A(n27317), .B(n28493), .Z(n28491) );
  XOR U40266 ( .A(n27318), .B(n28491), .Z(n30276) );
  XOR U40267 ( .A(n30277), .B(n30276), .Z(n30279) );
  IV U40268 ( .A(n27319), .Z(n27320) );
  NOR U40269 ( .A(n27321), .B(n27320), .Z(n30278) );
  IV U40270 ( .A(n27322), .Z(n27324) );
  NOR U40271 ( .A(n27324), .B(n27323), .Z(n30273) );
  NOR U40272 ( .A(n30278), .B(n30273), .Z(n27325) );
  XOR U40273 ( .A(n30279), .B(n27325), .Z(n28485) );
  XOR U40274 ( .A(n28486), .B(n28485), .Z(n28481) );
  IV U40275 ( .A(n27326), .Z(n27328) );
  NOR U40276 ( .A(n27328), .B(n27327), .Z(n28480) );
  IV U40277 ( .A(n27329), .Z(n27330) );
  NOR U40278 ( .A(n27331), .B(n27330), .Z(n28477) );
  NOR U40279 ( .A(n28480), .B(n28477), .Z(n27332) );
  XOR U40280 ( .A(n28481), .B(n27332), .Z(n28475) );
  IV U40281 ( .A(n27333), .Z(n27335) );
  NOR U40282 ( .A(n27335), .B(n27334), .Z(n33664) );
  IV U40283 ( .A(n27336), .Z(n27337) );
  NOR U40284 ( .A(n27338), .B(n27337), .Z(n27339) );
  NOR U40285 ( .A(n33664), .B(n27339), .Z(n28476) );
  XOR U40286 ( .A(n28475), .B(n28476), .Z(n30300) );
  IV U40287 ( .A(n27340), .Z(n27341) );
  NOR U40288 ( .A(n27342), .B(n27341), .Z(n28473) );
  IV U40289 ( .A(n27343), .Z(n27345) );
  NOR U40290 ( .A(n27345), .B(n27344), .Z(n30299) );
  NOR U40291 ( .A(n28473), .B(n30299), .Z(n27346) );
  XOR U40292 ( .A(n30300), .B(n27346), .Z(n30302) );
  XOR U40293 ( .A(n30303), .B(n30302), .Z(n37076) );
  IV U40294 ( .A(n27347), .Z(n27348) );
  NOR U40295 ( .A(n27349), .B(n27348), .Z(n37071) );
  IV U40296 ( .A(n27350), .Z(n27351) );
  NOR U40297 ( .A(n27352), .B(n27351), .Z(n37080) );
  NOR U40298 ( .A(n37071), .B(n37080), .Z(n28472) );
  XOR U40299 ( .A(n37076), .B(n28472), .Z(n30308) );
  XOR U40300 ( .A(n30309), .B(n30308), .Z(n28470) );
  IV U40301 ( .A(n27353), .Z(n27354) );
  NOR U40302 ( .A(n27355), .B(n27354), .Z(n28469) );
  IV U40303 ( .A(n27356), .Z(n27357) );
  NOR U40304 ( .A(n27358), .B(n27357), .Z(n28467) );
  NOR U40305 ( .A(n28469), .B(n28467), .Z(n27359) );
  XOR U40306 ( .A(n28470), .B(n27359), .Z(n27367) );
  IV U40307 ( .A(n27367), .Z(n27360) );
  NOR U40308 ( .A(n27361), .B(n27360), .Z(n31733) );
  IV U40309 ( .A(n27362), .Z(n27364) );
  NOR U40310 ( .A(n27364), .B(n27363), .Z(n27368) );
  IV U40311 ( .A(n27368), .Z(n27366) );
  XOR U40312 ( .A(n28469), .B(n28470), .Z(n27365) );
  NOR U40313 ( .A(n27366), .B(n27365), .Z(n31730) );
  NOR U40314 ( .A(n27368), .B(n27367), .Z(n27369) );
  NOR U40315 ( .A(n31730), .B(n27369), .Z(n30327) );
  NOR U40316 ( .A(n27370), .B(n30327), .Z(n27371) );
  NOR U40317 ( .A(n31733), .B(n27371), .Z(n30319) );
  IV U40318 ( .A(n27372), .Z(n27373) );
  NOR U40319 ( .A(n27374), .B(n27373), .Z(n30326) );
  IV U40320 ( .A(n27375), .Z(n27376) );
  NOR U40321 ( .A(n27377), .B(n27376), .Z(n30318) );
  NOR U40322 ( .A(n30326), .B(n30318), .Z(n27378) );
  XOR U40323 ( .A(n30319), .B(n27378), .Z(n30339) );
  IV U40324 ( .A(n27379), .Z(n27381) );
  NOR U40325 ( .A(n27381), .B(n27380), .Z(n30323) );
  IV U40326 ( .A(n27382), .Z(n27384) );
  NOR U40327 ( .A(n27384), .B(n27383), .Z(n30337) );
  NOR U40328 ( .A(n30323), .B(n30337), .Z(n27385) );
  XOR U40329 ( .A(n30339), .B(n27385), .Z(n28465) );
  IV U40330 ( .A(n27386), .Z(n27387) );
  NOR U40331 ( .A(n27388), .B(n27387), .Z(n28464) );
  IV U40332 ( .A(n27389), .Z(n27390) );
  NOR U40333 ( .A(n27391), .B(n27390), .Z(n30344) );
  NOR U40334 ( .A(n28464), .B(n30344), .Z(n27392) );
  XOR U40335 ( .A(n28465), .B(n27392), .Z(n37111) );
  XOR U40336 ( .A(n28462), .B(n37111), .Z(n27393) );
  IV U40337 ( .A(n27393), .Z(n28460) );
  XOR U40338 ( .A(n28457), .B(n28460), .Z(n28455) );
  IV U40339 ( .A(n27394), .Z(n27395) );
  NOR U40340 ( .A(n27396), .B(n27395), .Z(n28459) );
  IV U40341 ( .A(n27397), .Z(n27399) );
  NOR U40342 ( .A(n27399), .B(n27398), .Z(n28454) );
  NOR U40343 ( .A(n28459), .B(n28454), .Z(n27400) );
  XOR U40344 ( .A(n28455), .B(n27400), .Z(n30349) );
  IV U40345 ( .A(n27401), .Z(n27403) );
  NOR U40346 ( .A(n27403), .B(n27402), .Z(n33702) );
  IV U40347 ( .A(n27404), .Z(n27405) );
  NOR U40348 ( .A(n27406), .B(n27405), .Z(n33709) );
  NOR U40349 ( .A(n33702), .B(n33709), .Z(n30350) );
  XOR U40350 ( .A(n30349), .B(n30350), .Z(n30357) );
  IV U40351 ( .A(n27407), .Z(n27408) );
  NOR U40352 ( .A(n27409), .B(n27408), .Z(n30351) );
  IV U40353 ( .A(n27410), .Z(n27412) );
  NOR U40354 ( .A(n27412), .B(n27411), .Z(n30356) );
  NOR U40355 ( .A(n30351), .B(n30356), .Z(n27413) );
  XOR U40356 ( .A(n30357), .B(n27413), .Z(n27415) );
  XOR U40357 ( .A(n30361), .B(n27415), .Z(n27420) );
  NOR U40358 ( .A(n27414), .B(n27420), .Z(n37120) );
  IV U40359 ( .A(n27415), .Z(n30362) );
  IV U40360 ( .A(n27416), .Z(n27417) );
  NOR U40361 ( .A(n27418), .B(n27417), .Z(n27422) );
  IV U40362 ( .A(n27422), .Z(n27419) );
  NOR U40363 ( .A(n30362), .B(n27419), .Z(n35036) );
  NOR U40364 ( .A(n37120), .B(n35036), .Z(n30360) );
  IV U40365 ( .A(n30360), .Z(n30367) );
  NOR U40366 ( .A(n30367), .B(n27420), .Z(n27425) );
  NOR U40367 ( .A(n27422), .B(n27421), .Z(n27423) );
  NOR U40368 ( .A(n27423), .B(n30367), .Z(n27424) );
  NOR U40369 ( .A(n27425), .B(n27424), .Z(n35033) );
  XOR U40370 ( .A(n30369), .B(n35033), .Z(n27426) );
  IV U40371 ( .A(n27426), .Z(n30374) );
  XOR U40372 ( .A(n30370), .B(n30374), .Z(n28452) );
  IV U40373 ( .A(n28452), .Z(n27434) );
  IV U40374 ( .A(n27427), .Z(n27428) );
  NOR U40375 ( .A(n27429), .B(n27428), .Z(n30373) );
  IV U40376 ( .A(n27430), .Z(n27432) );
  NOR U40377 ( .A(n27432), .B(n27431), .Z(n28451) );
  NOR U40378 ( .A(n30373), .B(n28451), .Z(n27433) );
  XOR U40379 ( .A(n27434), .B(n27433), .Z(n30384) );
  XOR U40380 ( .A(n30380), .B(n30384), .Z(n30377) );
  XOR U40381 ( .A(n27435), .B(n30377), .Z(n28448) );
  XOR U40382 ( .A(n27436), .B(n28448), .Z(n30401) );
  XOR U40383 ( .A(n30394), .B(n30401), .Z(n28443) );
  XOR U40384 ( .A(n27437), .B(n28443), .Z(n28439) );
  XOR U40385 ( .A(n27438), .B(n28439), .Z(n28437) );
  XOR U40386 ( .A(n28434), .B(n28437), .Z(n27439) );
  NOR U40387 ( .A(n27440), .B(n27439), .Z(n33748) );
  IV U40388 ( .A(n27441), .Z(n27443) );
  NOR U40389 ( .A(n27443), .B(n27442), .Z(n28436) );
  NOR U40390 ( .A(n28434), .B(n28436), .Z(n27444) );
  XOR U40391 ( .A(n27444), .B(n28437), .Z(n30412) );
  NOR U40392 ( .A(n27445), .B(n30412), .Z(n27446) );
  NOR U40393 ( .A(n33748), .B(n27446), .Z(n30407) );
  XOR U40394 ( .A(n27447), .B(n30407), .Z(n30428) );
  XOR U40395 ( .A(n28433), .B(n30428), .Z(n28431) );
  XOR U40396 ( .A(n28432), .B(n28431), .Z(n30438) );
  IV U40397 ( .A(n27448), .Z(n27450) );
  NOR U40398 ( .A(n27450), .B(n27449), .Z(n30437) );
  IV U40399 ( .A(n27451), .Z(n27452) );
  NOR U40400 ( .A(n27453), .B(n27452), .Z(n30435) );
  NOR U40401 ( .A(n30437), .B(n30435), .Z(n27454) );
  XOR U40402 ( .A(n30438), .B(n27454), .Z(n28429) );
  IV U40403 ( .A(n27455), .Z(n27456) );
  NOR U40404 ( .A(n27457), .B(n27456), .Z(n34988) );
  IV U40405 ( .A(n27458), .Z(n27459) );
  NOR U40406 ( .A(n27460), .B(n27459), .Z(n37178) );
  NOR U40407 ( .A(n34988), .B(n37178), .Z(n28430) );
  XOR U40408 ( .A(n28429), .B(n28430), .Z(n31694) );
  IV U40409 ( .A(n27461), .Z(n27462) );
  NOR U40410 ( .A(n27463), .B(n27462), .Z(n31697) );
  IV U40411 ( .A(n27464), .Z(n27465) );
  NOR U40412 ( .A(n27466), .B(n27465), .Z(n31692) );
  NOR U40413 ( .A(n31697), .B(n31692), .Z(n30450) );
  XOR U40414 ( .A(n31694), .B(n30450), .Z(n30451) );
  XOR U40415 ( .A(n30452), .B(n30451), .Z(n30459) );
  IV U40416 ( .A(n27467), .Z(n27469) );
  NOR U40417 ( .A(n27469), .B(n27468), .Z(n30458) );
  IV U40418 ( .A(n27470), .Z(n27472) );
  NOR U40419 ( .A(n27472), .B(n27471), .Z(n30455) );
  NOR U40420 ( .A(n30458), .B(n30455), .Z(n27473) );
  XOR U40421 ( .A(n30459), .B(n27473), .Z(n28427) );
  XOR U40422 ( .A(n27474), .B(n28427), .Z(n33766) );
  XOR U40423 ( .A(n30475), .B(n33766), .Z(n30476) );
  XOR U40424 ( .A(n30477), .B(n30476), .Z(n33773) );
  IV U40425 ( .A(n27475), .Z(n27476) );
  NOR U40426 ( .A(n27477), .B(n27476), .Z(n37194) );
  IV U40427 ( .A(n27478), .Z(n27479) );
  NOR U40428 ( .A(n27480), .B(n27479), .Z(n34954) );
  NOR U40429 ( .A(n37194), .B(n34954), .Z(n33775) );
  XOR U40430 ( .A(n33773), .B(n33775), .Z(n30481) );
  XOR U40431 ( .A(n30482), .B(n30481), .Z(n28424) );
  XOR U40432 ( .A(n28425), .B(n28424), .Z(n27481) );
  NOR U40433 ( .A(n27490), .B(n27481), .Z(n27492) );
  IV U40434 ( .A(n27482), .Z(n27483) );
  NOR U40435 ( .A(n27484), .B(n27483), .Z(n27485) );
  IV U40436 ( .A(n27485), .Z(n27493) );
  NOR U40437 ( .A(n27492), .B(n27493), .Z(n31677) );
  IV U40438 ( .A(n27486), .Z(n27487) );
  NOR U40439 ( .A(n27488), .B(n27487), .Z(n27489) );
  IV U40440 ( .A(n27489), .Z(n28423) );
  IV U40441 ( .A(n27490), .Z(n27491) );
  NOR U40442 ( .A(n27491), .B(n28424), .Z(n33790) );
  NOR U40443 ( .A(n27492), .B(n33790), .Z(n27494) );
  IV U40444 ( .A(n27494), .Z(n28422) );
  XOR U40445 ( .A(n28423), .B(n28422), .Z(n27496) );
  NOR U40446 ( .A(n27494), .B(n27493), .Z(n27495) );
  NOR U40447 ( .A(n27496), .B(n27495), .Z(n27497) );
  NOR U40448 ( .A(n31677), .B(n27497), .Z(n30496) );
  IV U40449 ( .A(n27498), .Z(n27499) );
  NOR U40450 ( .A(n27500), .B(n27499), .Z(n34940) );
  IV U40451 ( .A(n27501), .Z(n27503) );
  NOR U40452 ( .A(n27503), .B(n27502), .Z(n34932) );
  NOR U40453 ( .A(n34940), .B(n34932), .Z(n30497) );
  XOR U40454 ( .A(n30496), .B(n30497), .Z(n30494) );
  XOR U40455 ( .A(n27504), .B(n30494), .Z(n30513) );
  XOR U40456 ( .A(n27505), .B(n30513), .Z(n28420) );
  XOR U40457 ( .A(n27506), .B(n28420), .Z(n28416) );
  XOR U40458 ( .A(n27507), .B(n28416), .Z(n30523) );
  XOR U40459 ( .A(n30522), .B(n30523), .Z(n30531) );
  XOR U40460 ( .A(n27508), .B(n30531), .Z(n27509) );
  IV U40461 ( .A(n27509), .Z(n30542) );
  XOR U40462 ( .A(n30537), .B(n30542), .Z(n30548) );
  IV U40463 ( .A(n27510), .Z(n27511) );
  NOR U40464 ( .A(n27512), .B(n27511), .Z(n30540) );
  IV U40465 ( .A(n27513), .Z(n27514) );
  NOR U40466 ( .A(n27515), .B(n27514), .Z(n30547) );
  NOR U40467 ( .A(n30540), .B(n30547), .Z(n27516) );
  XOR U40468 ( .A(n30548), .B(n27516), .Z(n30544) );
  XOR U40469 ( .A(n27517), .B(n30544), .Z(n28414) );
  XOR U40470 ( .A(n28411), .B(n28414), .Z(n28409) );
  IV U40471 ( .A(n28409), .Z(n27525) );
  IV U40472 ( .A(n27518), .Z(n27520) );
  NOR U40473 ( .A(n27520), .B(n27519), .Z(n28413) );
  IV U40474 ( .A(n27521), .Z(n27523) );
  NOR U40475 ( .A(n27523), .B(n27522), .Z(n28408) );
  NOR U40476 ( .A(n28413), .B(n28408), .Z(n27524) );
  XOR U40477 ( .A(n27525), .B(n27524), .Z(n30560) );
  XOR U40478 ( .A(n30556), .B(n30560), .Z(n30566) );
  XOR U40479 ( .A(n27526), .B(n30566), .Z(n30562) );
  XOR U40480 ( .A(n27527), .B(n30562), .Z(n30576) );
  XOR U40481 ( .A(n27528), .B(n30576), .Z(n28402) );
  XOR U40482 ( .A(n28403), .B(n28402), .Z(n31639) );
  XOR U40483 ( .A(n31640), .B(n31639), .Z(n27529) );
  IV U40484 ( .A(n27529), .Z(n28397) );
  XOR U40485 ( .A(n28396), .B(n28397), .Z(n28391) );
  IV U40486 ( .A(n28391), .Z(n27537) );
  IV U40487 ( .A(n27530), .Z(n27532) );
  NOR U40488 ( .A(n27532), .B(n27531), .Z(n28393) );
  IV U40489 ( .A(n27533), .Z(n27534) );
  NOR U40490 ( .A(n27535), .B(n27534), .Z(n28390) );
  NOR U40491 ( .A(n28393), .B(n28390), .Z(n27536) );
  XOR U40492 ( .A(n27537), .B(n27536), .Z(n31628) );
  IV U40493 ( .A(n27538), .Z(n27540) );
  NOR U40494 ( .A(n27540), .B(n27539), .Z(n33852) );
  IV U40495 ( .A(n27541), .Z(n27543) );
  NOR U40496 ( .A(n27543), .B(n27542), .Z(n31627) );
  NOR U40497 ( .A(n33852), .B(n31627), .Z(n28387) );
  XOR U40498 ( .A(n31628), .B(n28387), .Z(n27546) );
  XOR U40499 ( .A(n28385), .B(n27546), .Z(n27544) );
  NOR U40500 ( .A(n27545), .B(n27544), .Z(n31619) );
  IV U40501 ( .A(n27546), .Z(n28384) );
  IV U40502 ( .A(n27547), .Z(n27549) );
  NOR U40503 ( .A(n27549), .B(n27548), .Z(n28382) );
  NOR U40504 ( .A(n27550), .B(n28382), .Z(n27551) );
  XOR U40505 ( .A(n28384), .B(n27551), .Z(n27559) );
  NOR U40506 ( .A(n27552), .B(n27559), .Z(n27553) );
  NOR U40507 ( .A(n31619), .B(n27553), .Z(n27562) );
  IV U40508 ( .A(n27562), .Z(n27554) );
  NOR U40509 ( .A(n27555), .B(n27554), .Z(n33862) );
  IV U40510 ( .A(n27556), .Z(n27558) );
  NOR U40511 ( .A(n27558), .B(n27557), .Z(n27563) );
  IV U40512 ( .A(n27563), .Z(n27561) );
  IV U40513 ( .A(n27559), .Z(n27560) );
  NOR U40514 ( .A(n27561), .B(n27560), .Z(n31617) );
  NOR U40515 ( .A(n27563), .B(n27562), .Z(n27564) );
  NOR U40516 ( .A(n31617), .B(n27564), .Z(n27573) );
  NOR U40517 ( .A(n27565), .B(n27573), .Z(n27566) );
  NOR U40518 ( .A(n33862), .B(n27566), .Z(n28378) );
  IV U40519 ( .A(n27567), .Z(n27568) );
  NOR U40520 ( .A(n27569), .B(n27568), .Z(n27580) );
  IV U40521 ( .A(n27580), .Z(n28380) );
  NOR U40522 ( .A(n28378), .B(n28380), .Z(n27582) );
  IV U40523 ( .A(n27570), .Z(n27572) );
  NOR U40524 ( .A(n27572), .B(n27571), .Z(n27576) );
  IV U40525 ( .A(n27576), .Z(n27575) );
  IV U40526 ( .A(n27573), .Z(n27574) );
  NOR U40527 ( .A(n27575), .B(n27574), .Z(n33865) );
  NOR U40528 ( .A(n28378), .B(n27576), .Z(n27577) );
  NOR U40529 ( .A(n33865), .B(n27577), .Z(n27578) );
  IV U40530 ( .A(n27578), .Z(n27579) );
  NOR U40531 ( .A(n27580), .B(n27579), .Z(n27581) );
  NOR U40532 ( .A(n27582), .B(n27581), .Z(n30586) );
  XOR U40533 ( .A(n27583), .B(n30586), .Z(n28376) );
  XOR U40534 ( .A(n28377), .B(n28376), .Z(n28374) );
  XOR U40535 ( .A(n28373), .B(n28374), .Z(n30603) );
  XOR U40536 ( .A(n27584), .B(n30603), .Z(n30605) );
  XOR U40537 ( .A(n33882), .B(n30605), .Z(n30611) );
  XOR U40538 ( .A(n30606), .B(n30611), .Z(n27585) );
  NOR U40539 ( .A(n27594), .B(n27585), .Z(n30621) );
  IV U40540 ( .A(n27586), .Z(n27588) );
  NOR U40541 ( .A(n27588), .B(n27587), .Z(n27589) );
  IV U40542 ( .A(n27589), .Z(n30624) );
  IV U40543 ( .A(n27590), .Z(n27591) );
  NOR U40544 ( .A(n27592), .B(n27591), .Z(n30610) );
  NOR U40545 ( .A(n30606), .B(n30610), .Z(n27593) );
  XOR U40546 ( .A(n27593), .B(n30611), .Z(n27595) );
  IV U40547 ( .A(n27595), .Z(n30623) );
  XOR U40548 ( .A(n30624), .B(n30623), .Z(n27597) );
  NOR U40549 ( .A(n27595), .B(n27594), .Z(n27596) );
  NOR U40550 ( .A(n27597), .B(n27596), .Z(n27598) );
  NOR U40551 ( .A(n30621), .B(n27598), .Z(n30625) );
  XOR U40552 ( .A(n30626), .B(n30625), .Z(n37298) );
  XOR U40553 ( .A(n28370), .B(n37298), .Z(n28366) );
  XOR U40554 ( .A(n28367), .B(n28366), .Z(n31605) );
  XOR U40555 ( .A(n28368), .B(n31605), .Z(n30629) );
  IV U40556 ( .A(n27599), .Z(n27601) );
  NOR U40557 ( .A(n27601), .B(n27600), .Z(n31600) );
  IV U40558 ( .A(n27602), .Z(n27603) );
  NOR U40559 ( .A(n27604), .B(n27603), .Z(n31595) );
  NOR U40560 ( .A(n31600), .B(n31595), .Z(n30630) );
  XOR U40561 ( .A(n30629), .B(n30630), .Z(n30632) );
  XOR U40562 ( .A(n27605), .B(n30632), .Z(n28362) );
  IV U40563 ( .A(n27606), .Z(n27607) );
  NOR U40564 ( .A(n27608), .B(n27607), .Z(n31587) );
  IV U40565 ( .A(n27609), .Z(n27610) );
  NOR U40566 ( .A(n27611), .B(n27610), .Z(n27612) );
  NOR U40567 ( .A(n31587), .B(n27612), .Z(n28363) );
  XOR U40568 ( .A(n28362), .B(n28363), .Z(n33908) );
  XOR U40569 ( .A(n28357), .B(n33908), .Z(n28355) );
  IV U40570 ( .A(n27613), .Z(n27615) );
  NOR U40571 ( .A(n27615), .B(n27614), .Z(n28358) );
  IV U40572 ( .A(n27616), .Z(n27617) );
  NOR U40573 ( .A(n27618), .B(n27617), .Z(n28354) );
  NOR U40574 ( .A(n28358), .B(n28354), .Z(n27619) );
  XOR U40575 ( .A(n28355), .B(n27619), .Z(n30642) );
  XOR U40576 ( .A(n30638), .B(n30642), .Z(n30646) );
  XOR U40577 ( .A(n27620), .B(n30646), .Z(n28349) );
  XOR U40578 ( .A(n28350), .B(n28349), .Z(n28347) );
  IV U40579 ( .A(n27621), .Z(n27623) );
  NOR U40580 ( .A(n27623), .B(n27622), .Z(n28344) );
  IV U40581 ( .A(n27624), .Z(n27626) );
  NOR U40582 ( .A(n27626), .B(n27625), .Z(n28346) );
  NOR U40583 ( .A(n28344), .B(n28346), .Z(n27627) );
  XOR U40584 ( .A(n28347), .B(n27627), .Z(n27628) );
  NOR U40585 ( .A(n27629), .B(n27628), .Z(n27632) );
  IV U40586 ( .A(n27629), .Z(n27631) );
  XOR U40587 ( .A(n28344), .B(n28347), .Z(n27630) );
  NOR U40588 ( .A(n27631), .B(n27630), .Z(n38348) );
  NOR U40589 ( .A(n27632), .B(n38348), .Z(n28340) );
  XOR U40590 ( .A(n28343), .B(n28340), .Z(n28337) );
  XOR U40591 ( .A(n27633), .B(n28337), .Z(n28333) );
  XOR U40592 ( .A(n27634), .B(n28333), .Z(n30660) );
  XOR U40593 ( .A(n27635), .B(n30660), .Z(n28329) );
  IV U40594 ( .A(n27636), .Z(n27637) );
  NOR U40595 ( .A(n27638), .B(n27637), .Z(n28328) );
  IV U40596 ( .A(n27639), .Z(n27641) );
  NOR U40597 ( .A(n27641), .B(n27640), .Z(n30675) );
  NOR U40598 ( .A(n28328), .B(n30675), .Z(n27642) );
  XOR U40599 ( .A(n28329), .B(n27642), .Z(n30683) );
  IV U40600 ( .A(n27643), .Z(n27645) );
  NOR U40601 ( .A(n27645), .B(n27644), .Z(n30678) );
  IV U40602 ( .A(n27646), .Z(n27647) );
  NOR U40603 ( .A(n27648), .B(n27647), .Z(n30681) );
  NOR U40604 ( .A(n30678), .B(n30681), .Z(n27649) );
  XOR U40605 ( .A(n30683), .B(n27649), .Z(n28322) );
  XOR U40606 ( .A(n28323), .B(n28322), .Z(n28325) );
  XOR U40607 ( .A(n27650), .B(n28325), .Z(n28313) );
  XOR U40608 ( .A(n27651), .B(n28313), .Z(n34760) );
  XOR U40609 ( .A(n28316), .B(n34760), .Z(n28305) );
  IV U40610 ( .A(n27652), .Z(n27653) );
  NOR U40611 ( .A(n27654), .B(n27653), .Z(n28304) );
  IV U40612 ( .A(n27655), .Z(n27656) );
  NOR U40613 ( .A(n27657), .B(n27656), .Z(n28308) );
  NOR U40614 ( .A(n28304), .B(n28308), .Z(n27658) );
  XOR U40615 ( .A(n28305), .B(n27658), .Z(n28303) );
  IV U40616 ( .A(n27659), .Z(n27660) );
  NOR U40617 ( .A(n27661), .B(n27660), .Z(n28301) );
  IV U40618 ( .A(n27662), .Z(n27664) );
  NOR U40619 ( .A(n27664), .B(n27663), .Z(n28299) );
  NOR U40620 ( .A(n28301), .B(n28299), .Z(n27665) );
  XOR U40621 ( .A(n28303), .B(n27665), .Z(n28294) );
  IV U40622 ( .A(n28294), .Z(n33993) );
  XOR U40623 ( .A(n33992), .B(n33993), .Z(n31551) );
  XOR U40624 ( .A(n28295), .B(n31551), .Z(n28288) );
  IV U40625 ( .A(n27666), .Z(n27667) );
  NOR U40626 ( .A(n27668), .B(n27667), .Z(n28291) );
  IV U40627 ( .A(n27669), .Z(n27670) );
  NOR U40628 ( .A(n27671), .B(n27670), .Z(n28289) );
  NOR U40629 ( .A(n28291), .B(n28289), .Z(n27672) );
  XOR U40630 ( .A(n28288), .B(n27672), .Z(n28286) );
  XOR U40631 ( .A(n28285), .B(n28286), .Z(n30694) );
  IV U40632 ( .A(n27673), .Z(n27675) );
  NOR U40633 ( .A(n27675), .B(n27674), .Z(n28282) );
  IV U40634 ( .A(n27676), .Z(n27678) );
  NOR U40635 ( .A(n27678), .B(n27677), .Z(n30693) );
  NOR U40636 ( .A(n28282), .B(n30693), .Z(n27679) );
  XOR U40637 ( .A(n30694), .B(n27679), .Z(n30691) );
  XOR U40638 ( .A(n30692), .B(n30691), .Z(n31528) );
  XOR U40639 ( .A(n30702), .B(n31528), .Z(n28280) );
  XOR U40640 ( .A(n27680), .B(n28280), .Z(n31523) );
  XOR U40641 ( .A(n30708), .B(n31523), .Z(n31513) );
  XOR U40642 ( .A(n30710), .B(n31513), .Z(n31507) );
  XOR U40643 ( .A(n30714), .B(n31507), .Z(n30715) );
  XOR U40644 ( .A(n30716), .B(n30715), .Z(n34009) );
  IV U40645 ( .A(n34009), .Z(n27688) );
  IV U40646 ( .A(n27681), .Z(n27683) );
  NOR U40647 ( .A(n27683), .B(n27682), .Z(n34008) );
  IV U40648 ( .A(n27684), .Z(n27686) );
  NOR U40649 ( .A(n27686), .B(n27685), .Z(n27687) );
  NOR U40650 ( .A(n34008), .B(n27687), .Z(n28277) );
  XOR U40651 ( .A(n27688), .B(n28277), .Z(n31492) );
  XOR U40652 ( .A(n28272), .B(n31492), .Z(n28270) );
  IV U40653 ( .A(n27689), .Z(n27691) );
  NOR U40654 ( .A(n27691), .B(n27690), .Z(n28273) );
  IV U40655 ( .A(n27692), .Z(n27693) );
  NOR U40656 ( .A(n27694), .B(n27693), .Z(n28269) );
  NOR U40657 ( .A(n28273), .B(n28269), .Z(n27695) );
  XOR U40658 ( .A(n28270), .B(n27695), .Z(n31478) );
  IV U40659 ( .A(n27696), .Z(n27697) );
  NOR U40660 ( .A(n27698), .B(n27697), .Z(n31484) );
  IV U40661 ( .A(n27699), .Z(n27701) );
  NOR U40662 ( .A(n27701), .B(n27700), .Z(n31477) );
  NOR U40663 ( .A(n31484), .B(n31477), .Z(n30722) );
  XOR U40664 ( .A(n31478), .B(n30722), .Z(n30723) );
  IV U40665 ( .A(n27702), .Z(n27704) );
  NOR U40666 ( .A(n27704), .B(n27703), .Z(n37458) );
  IV U40667 ( .A(n27705), .Z(n27706) );
  NOR U40668 ( .A(n27707), .B(n27706), .Z(n37467) );
  NOR U40669 ( .A(n37458), .B(n37467), .Z(n30724) );
  XOR U40670 ( .A(n30723), .B(n30724), .Z(n28267) );
  XOR U40671 ( .A(n28266), .B(n28267), .Z(n28262) );
  XOR U40672 ( .A(n27708), .B(n28262), .Z(n30729) );
  XOR U40673 ( .A(n30730), .B(n30729), .Z(n30732) );
  XOR U40674 ( .A(n30731), .B(n30732), .Z(n27709) );
  NOR U40675 ( .A(n27710), .B(n27709), .Z(n30739) );
  IV U40676 ( .A(n27711), .Z(n27713) );
  NOR U40677 ( .A(n27713), .B(n27712), .Z(n28259) );
  NOR U40678 ( .A(n30731), .B(n28259), .Z(n27714) );
  XOR U40679 ( .A(n27714), .B(n30732), .Z(n28256) );
  NOR U40680 ( .A(n27715), .B(n28256), .Z(n27716) );
  NOR U40681 ( .A(n30739), .B(n27716), .Z(n30748) );
  XOR U40682 ( .A(n27717), .B(n30748), .Z(n28254) );
  XOR U40683 ( .A(n27718), .B(n28254), .Z(n28248) );
  XOR U40684 ( .A(n27719), .B(n28248), .Z(n31438) );
  XOR U40685 ( .A(n28243), .B(n31438), .Z(n28241) );
  XOR U40686 ( .A(n28245), .B(n28241), .Z(n28238) );
  XOR U40687 ( .A(n27720), .B(n28238), .Z(n28230) );
  XOR U40688 ( .A(n27721), .B(n28230), .Z(n30778) );
  XOR U40689 ( .A(n27722), .B(n30778), .Z(n30766) );
  XOR U40690 ( .A(n27723), .B(n30766), .Z(n31426) );
  XOR U40691 ( .A(n28227), .B(n31426), .Z(n30789) );
  XOR U40692 ( .A(n30790), .B(n30789), .Z(n28225) );
  IV U40693 ( .A(n27724), .Z(n27725) );
  NOR U40694 ( .A(n27726), .B(n27725), .Z(n37538) );
  IV U40695 ( .A(n27727), .Z(n27728) );
  NOR U40696 ( .A(n27729), .B(n27728), .Z(n27730) );
  NOR U40697 ( .A(n37538), .B(n27730), .Z(n28226) );
  XOR U40698 ( .A(n28225), .B(n28226), .Z(n30799) );
  XOR U40699 ( .A(n27731), .B(n30799), .Z(n27732) );
  IV U40700 ( .A(n27732), .Z(n28222) );
  XOR U40701 ( .A(n28220), .B(n28222), .Z(n27743) );
  IV U40702 ( .A(n27743), .Z(n27741) );
  IV U40703 ( .A(n27733), .Z(n27735) );
  NOR U40704 ( .A(n27735), .B(n27734), .Z(n27745) );
  IV U40705 ( .A(n27736), .Z(n27737) );
  NOR U40706 ( .A(n27738), .B(n27737), .Z(n27742) );
  NOR U40707 ( .A(n27745), .B(n27742), .Z(n27739) );
  IV U40708 ( .A(n27739), .Z(n27740) );
  NOR U40709 ( .A(n27741), .B(n27740), .Z(n27748) );
  IV U40710 ( .A(n27742), .Z(n27744) );
  NOR U40711 ( .A(n27744), .B(n27743), .Z(n34065) );
  IV U40712 ( .A(n27745), .Z(n27746) );
  NOR U40713 ( .A(n28222), .B(n27746), .Z(n34060) );
  NOR U40714 ( .A(n34065), .B(n34060), .Z(n27747) );
  IV U40715 ( .A(n27747), .Z(n28219) );
  NOR U40716 ( .A(n27748), .B(n28219), .Z(n28214) );
  IV U40717 ( .A(n27749), .Z(n27750) );
  NOR U40718 ( .A(n27751), .B(n27750), .Z(n28216) );
  IV U40719 ( .A(n27752), .Z(n27753) );
  NOR U40720 ( .A(n27754), .B(n27753), .Z(n28213) );
  NOR U40721 ( .A(n28216), .B(n28213), .Z(n27755) );
  XOR U40722 ( .A(n28214), .B(n27755), .Z(n30805) );
  XOR U40723 ( .A(n28211), .B(n30805), .Z(n30810) );
  XOR U40724 ( .A(n27756), .B(n30810), .Z(n30806) );
  XOR U40725 ( .A(n27757), .B(n30806), .Z(n30830) );
  XOR U40726 ( .A(n27758), .B(n30830), .Z(n30818) );
  XOR U40727 ( .A(n27759), .B(n30818), .Z(n30841) );
  IV U40728 ( .A(n27760), .Z(n27762) );
  NOR U40729 ( .A(n27762), .B(n27761), .Z(n30840) );
  IV U40730 ( .A(n27763), .Z(n27765) );
  NOR U40731 ( .A(n27765), .B(n27764), .Z(n28209) );
  NOR U40732 ( .A(n30840), .B(n28209), .Z(n27766) );
  XOR U40733 ( .A(n30841), .B(n27766), .Z(n27767) );
  NOR U40734 ( .A(n27768), .B(n27767), .Z(n27771) );
  IV U40735 ( .A(n27768), .Z(n27770) );
  XOR U40736 ( .A(n30840), .B(n30841), .Z(n27769) );
  NOR U40737 ( .A(n27770), .B(n27769), .Z(n30857) );
  NOR U40738 ( .A(n27771), .B(n30857), .Z(n30852) );
  IV U40739 ( .A(n27772), .Z(n27774) );
  NOR U40740 ( .A(n27774), .B(n27773), .Z(n31414) );
  IV U40741 ( .A(n27775), .Z(n27777) );
  NOR U40742 ( .A(n27777), .B(n27776), .Z(n31408) );
  NOR U40743 ( .A(n31414), .B(n31408), .Z(n30853) );
  XOR U40744 ( .A(n30852), .B(n30853), .Z(n30869) );
  XOR U40745 ( .A(n27778), .B(n30869), .Z(n27779) );
  IV U40746 ( .A(n27779), .Z(n28208) );
  XOR U40747 ( .A(n27780), .B(n28208), .Z(n31385) );
  XOR U40748 ( .A(n31398), .B(n31385), .Z(n31391) );
  XOR U40749 ( .A(n30876), .B(n31391), .Z(n30886) );
  XOR U40750 ( .A(n27781), .B(n30886), .Z(n30880) );
  XOR U40751 ( .A(n30881), .B(n30880), .Z(n30903) );
  XOR U40752 ( .A(n30900), .B(n30903), .Z(n30892) );
  IV U40753 ( .A(n27782), .Z(n27784) );
  NOR U40754 ( .A(n27784), .B(n27783), .Z(n30902) );
  IV U40755 ( .A(n27785), .Z(n27786) );
  NOR U40756 ( .A(n27787), .B(n27786), .Z(n30891) );
  NOR U40757 ( .A(n30902), .B(n30891), .Z(n27788) );
  XOR U40758 ( .A(n30892), .B(n27788), .Z(n28201) );
  IV U40759 ( .A(n27789), .Z(n27790) );
  NOR U40760 ( .A(n27791), .B(n27790), .Z(n30895) );
  IV U40761 ( .A(n27792), .Z(n27794) );
  NOR U40762 ( .A(n27794), .B(n27793), .Z(n28202) );
  NOR U40763 ( .A(n30895), .B(n28202), .Z(n31366) );
  XOR U40764 ( .A(n28201), .B(n31366), .Z(n30922) );
  XOR U40765 ( .A(n30919), .B(n30922), .Z(n30929) );
  IV U40766 ( .A(n27795), .Z(n27796) );
  NOR U40767 ( .A(n27797), .B(n27796), .Z(n30921) );
  IV U40768 ( .A(n27798), .Z(n27799) );
  NOR U40769 ( .A(n27800), .B(n27799), .Z(n30928) );
  NOR U40770 ( .A(n30921), .B(n30928), .Z(n27801) );
  XOR U40771 ( .A(n30929), .B(n27801), .Z(n28198) );
  IV U40772 ( .A(n27802), .Z(n27804) );
  NOR U40773 ( .A(n27804), .B(n27803), .Z(n30925) );
  IV U40774 ( .A(n27805), .Z(n27806) );
  NOR U40775 ( .A(n27807), .B(n27806), .Z(n28199) );
  NOR U40776 ( .A(n30925), .B(n28199), .Z(n27808) );
  XOR U40777 ( .A(n28198), .B(n27808), .Z(n30932) );
  XOR U40778 ( .A(n28196), .B(n30932), .Z(n28194) );
  IV U40779 ( .A(n27809), .Z(n27810) );
  NOR U40780 ( .A(n27811), .B(n27810), .Z(n30931) );
  IV U40781 ( .A(n27812), .Z(n27814) );
  NOR U40782 ( .A(n27814), .B(n27813), .Z(n28193) );
  NOR U40783 ( .A(n30931), .B(n28193), .Z(n27815) );
  XOR U40784 ( .A(n28194), .B(n27815), .Z(n28190) );
  IV U40785 ( .A(n27816), .Z(n27817) );
  NOR U40786 ( .A(n27818), .B(n27817), .Z(n28191) );
  IV U40787 ( .A(n27819), .Z(n27820) );
  NOR U40788 ( .A(n27821), .B(n27820), .Z(n30935) );
  NOR U40789 ( .A(n28191), .B(n30935), .Z(n27822) );
  XOR U40790 ( .A(n28190), .B(n27822), .Z(n31357) );
  IV U40791 ( .A(n27823), .Z(n27824) );
  NOR U40792 ( .A(n27825), .B(n27824), .Z(n34129) );
  IV U40793 ( .A(n27826), .Z(n27828) );
  NOR U40794 ( .A(n27828), .B(n27827), .Z(n31356) );
  NOR U40795 ( .A(n34129), .B(n31356), .Z(n30941) );
  XOR U40796 ( .A(n31357), .B(n30941), .Z(n30939) );
  XOR U40797 ( .A(n30943), .B(n30939), .Z(n30950) );
  XOR U40798 ( .A(n27829), .B(n30950), .Z(n28185) );
  XOR U40799 ( .A(n28186), .B(n28185), .Z(n30959) );
  XOR U40800 ( .A(n27830), .B(n30959), .Z(n27831) );
  IV U40801 ( .A(n27831), .Z(n30955) );
  XOR U40802 ( .A(n27832), .B(n30955), .Z(n30980) );
  XOR U40803 ( .A(n30978), .B(n30980), .Z(n30973) );
  IV U40804 ( .A(n27833), .Z(n27835) );
  NOR U40805 ( .A(n27835), .B(n27834), .Z(n30977) );
  IV U40806 ( .A(n27836), .Z(n27837) );
  NOR U40807 ( .A(n27838), .B(n27837), .Z(n30988) );
  NOR U40808 ( .A(n30977), .B(n30988), .Z(n30974) );
  XOR U40809 ( .A(n30973), .B(n30974), .Z(n30995) );
  XOR U40810 ( .A(n30996), .B(n30995), .Z(n30999) );
  XOR U40811 ( .A(n28181), .B(n30999), .Z(n28179) );
  IV U40812 ( .A(n27839), .Z(n27841) );
  NOR U40813 ( .A(n27841), .B(n27840), .Z(n30998) );
  IV U40814 ( .A(n27842), .Z(n27843) );
  NOR U40815 ( .A(n27844), .B(n27843), .Z(n28178) );
  NOR U40816 ( .A(n30998), .B(n28178), .Z(n27845) );
  XOR U40817 ( .A(n28179), .B(n27845), .Z(n31003) );
  XOR U40818 ( .A(n31001), .B(n31003), .Z(n31011) );
  XOR U40819 ( .A(n27846), .B(n31011), .Z(n28172) );
  XOR U40820 ( .A(n27847), .B(n28172), .Z(n28167) );
  XOR U40821 ( .A(n27848), .B(n28167), .Z(n28159) );
  IV U40822 ( .A(n27849), .Z(n27850) );
  NOR U40823 ( .A(n27851), .B(n27850), .Z(n28161) );
  IV U40824 ( .A(n27852), .Z(n27854) );
  NOR U40825 ( .A(n27854), .B(n27853), .Z(n28158) );
  NOR U40826 ( .A(n28161), .B(n28158), .Z(n27855) );
  XOR U40827 ( .A(n28159), .B(n27855), .Z(n31315) );
  XOR U40828 ( .A(n28153), .B(n31315), .Z(n27856) );
  IV U40829 ( .A(n27856), .Z(n28155) );
  XOR U40830 ( .A(n28154), .B(n28155), .Z(n31020) );
  IV U40831 ( .A(n27857), .Z(n27858) );
  NOR U40832 ( .A(n27859), .B(n27858), .Z(n28151) );
  IV U40833 ( .A(n27860), .Z(n27862) );
  NOR U40834 ( .A(n27862), .B(n27861), .Z(n31019) );
  NOR U40835 ( .A(n28151), .B(n31019), .Z(n27863) );
  XOR U40836 ( .A(n31020), .B(n27863), .Z(n31016) );
  IV U40837 ( .A(n27864), .Z(n27866) );
  NOR U40838 ( .A(n27866), .B(n27865), .Z(n31017) );
  IV U40839 ( .A(n27867), .Z(n27868) );
  NOR U40840 ( .A(n27869), .B(n27868), .Z(n31023) );
  NOR U40841 ( .A(n31017), .B(n31023), .Z(n27870) );
  XOR U40842 ( .A(n31016), .B(n27870), .Z(n34505) );
  XOR U40843 ( .A(n34504), .B(n34505), .Z(n31031) );
  IV U40844 ( .A(n27871), .Z(n27873) );
  NOR U40845 ( .A(n27873), .B(n27872), .Z(n31026) );
  IV U40846 ( .A(n27874), .Z(n27875) );
  NOR U40847 ( .A(n27876), .B(n27875), .Z(n31030) );
  NOR U40848 ( .A(n31026), .B(n31030), .Z(n27877) );
  XOR U40849 ( .A(n31031), .B(n27877), .Z(n28145) );
  IV U40850 ( .A(n27878), .Z(n27879) );
  NOR U40851 ( .A(n27880), .B(n27879), .Z(n28148) );
  IV U40852 ( .A(n27881), .Z(n27883) );
  NOR U40853 ( .A(n27883), .B(n27882), .Z(n28146) );
  NOR U40854 ( .A(n28148), .B(n28146), .Z(n27884) );
  XOR U40855 ( .A(n28145), .B(n27884), .Z(n34196) );
  IV U40856 ( .A(n27885), .Z(n27887) );
  NOR U40857 ( .A(n27887), .B(n27886), .Z(n34194) );
  IV U40858 ( .A(n27888), .Z(n27889) );
  NOR U40859 ( .A(n27890), .B(n27889), .Z(n34201) );
  NOR U40860 ( .A(n34194), .B(n34201), .Z(n28144) );
  XOR U40861 ( .A(n34196), .B(n28144), .Z(n27891) );
  IV U40862 ( .A(n27891), .Z(n31289) );
  XOR U40863 ( .A(n31043), .B(n31289), .Z(n31044) );
  IV U40864 ( .A(n27892), .Z(n27894) );
  NOR U40865 ( .A(n27894), .B(n27893), .Z(n31285) );
  IV U40866 ( .A(n27895), .Z(n27897) );
  NOR U40867 ( .A(n27897), .B(n27896), .Z(n31280) );
  NOR U40868 ( .A(n31285), .B(n31280), .Z(n31045) );
  XOR U40869 ( .A(n31044), .B(n31045), .Z(n34205) );
  XOR U40870 ( .A(n31049), .B(n34205), .Z(n31050) );
  IV U40871 ( .A(n27898), .Z(n27900) );
  NOR U40872 ( .A(n27900), .B(n27899), .Z(n34215) );
  IV U40873 ( .A(n27901), .Z(n27903) );
  NOR U40874 ( .A(n27903), .B(n27902), .Z(n31275) );
  NOR U40875 ( .A(n34215), .B(n31275), .Z(n31051) );
  XOR U40876 ( .A(n31050), .B(n31051), .Z(n31056) );
  XOR U40877 ( .A(n27904), .B(n31056), .Z(n31059) );
  IV U40878 ( .A(n27905), .Z(n27907) );
  NOR U40879 ( .A(n27907), .B(n27906), .Z(n31058) );
  IV U40880 ( .A(n27908), .Z(n27909) );
  NOR U40881 ( .A(n27910), .B(n27909), .Z(n31063) );
  NOR U40882 ( .A(n31058), .B(n31063), .Z(n27911) );
  XOR U40883 ( .A(n31059), .B(n27911), .Z(n31071) );
  IV U40884 ( .A(n27912), .Z(n27914) );
  NOR U40885 ( .A(n27914), .B(n27913), .Z(n27915) );
  IV U40886 ( .A(n27915), .Z(n27923) );
  NOR U40887 ( .A(n31071), .B(n27923), .Z(n31077) );
  IV U40888 ( .A(n27916), .Z(n27918) );
  NOR U40889 ( .A(n27918), .B(n27917), .Z(n27919) );
  IV U40890 ( .A(n27919), .Z(n28140) );
  IV U40891 ( .A(n27920), .Z(n27921) );
  NOR U40892 ( .A(n27922), .B(n27921), .Z(n31069) );
  XOR U40893 ( .A(n31069), .B(n31071), .Z(n28139) );
  XOR U40894 ( .A(n28140), .B(n28139), .Z(n27926) );
  IV U40895 ( .A(n28139), .Z(n27924) );
  NOR U40896 ( .A(n27924), .B(n27923), .Z(n27925) );
  NOR U40897 ( .A(n27926), .B(n27925), .Z(n27927) );
  NOR U40898 ( .A(n31077), .B(n27927), .Z(n28133) );
  XOR U40899 ( .A(n27928), .B(n28133), .Z(n28131) );
  XOR U40900 ( .A(n28127), .B(n28131), .Z(n31083) );
  IV U40901 ( .A(n27929), .Z(n27930) );
  NOR U40902 ( .A(n27931), .B(n27930), .Z(n28129) );
  IV U40903 ( .A(n27932), .Z(n27933) );
  NOR U40904 ( .A(n27934), .B(n27933), .Z(n31082) );
  NOR U40905 ( .A(n28129), .B(n31082), .Z(n27935) );
  XOR U40906 ( .A(n31083), .B(n27935), .Z(n28120) );
  IV U40907 ( .A(n27936), .Z(n27938) );
  NOR U40908 ( .A(n27938), .B(n27937), .Z(n28124) );
  IV U40909 ( .A(n27939), .Z(n27940) );
  NOR U40910 ( .A(n27941), .B(n27940), .Z(n28121) );
  NOR U40911 ( .A(n28124), .B(n28121), .Z(n27942) );
  XOR U40912 ( .A(n28120), .B(n27942), .Z(n31262) );
  XOR U40913 ( .A(n31091), .B(n31262), .Z(n28118) );
  XOR U40914 ( .A(n27943), .B(n28118), .Z(n34461) );
  XOR U40915 ( .A(n31101), .B(n34461), .Z(n31102) );
  XOR U40916 ( .A(n31103), .B(n31102), .Z(n31107) );
  IV U40917 ( .A(n27944), .Z(n27946) );
  NOR U40918 ( .A(n27946), .B(n27945), .Z(n31106) );
  IV U40919 ( .A(n27947), .Z(n27949) );
  NOR U40920 ( .A(n27949), .B(n27948), .Z(n31246) );
  NOR U40921 ( .A(n31106), .B(n31246), .Z(n27950) );
  XOR U40922 ( .A(n31107), .B(n27950), .Z(n28110) );
  IV U40923 ( .A(n27951), .Z(n27952) );
  NOR U40924 ( .A(n27953), .B(n27952), .Z(n28107) );
  IV U40925 ( .A(n27954), .Z(n27956) );
  NOR U40926 ( .A(n27956), .B(n27955), .Z(n28111) );
  NOR U40927 ( .A(n28107), .B(n28111), .Z(n27957) );
  XOR U40928 ( .A(n28110), .B(n27957), .Z(n28104) );
  IV U40929 ( .A(n27958), .Z(n27960) );
  NOR U40930 ( .A(n27960), .B(n27959), .Z(n28106) );
  IV U40931 ( .A(n27961), .Z(n27962) );
  NOR U40932 ( .A(n27963), .B(n27962), .Z(n28103) );
  NOR U40933 ( .A(n28106), .B(n28103), .Z(n27964) );
  XOR U40934 ( .A(n28104), .B(n27964), .Z(n31110) );
  IV U40935 ( .A(n27965), .Z(n27966) );
  NOR U40936 ( .A(n27967), .B(n27966), .Z(n34272) );
  IV U40937 ( .A(n27968), .Z(n27970) );
  NOR U40938 ( .A(n27970), .B(n27969), .Z(n34268) );
  NOR U40939 ( .A(n34272), .B(n34268), .Z(n31111) );
  XOR U40940 ( .A(n31110), .B(n31111), .Z(n31120) );
  IV U40941 ( .A(n27971), .Z(n27973) );
  NOR U40942 ( .A(n27973), .B(n27972), .Z(n31112) );
  IV U40943 ( .A(n27974), .Z(n27975) );
  NOR U40944 ( .A(n27976), .B(n27975), .Z(n31119) );
  NOR U40945 ( .A(n31112), .B(n31119), .Z(n27977) );
  XOR U40946 ( .A(n31120), .B(n27977), .Z(n31116) );
  IV U40947 ( .A(n27978), .Z(n27979) );
  NOR U40948 ( .A(n27980), .B(n27979), .Z(n31117) );
  IV U40949 ( .A(n27981), .Z(n27982) );
  NOR U40950 ( .A(n27983), .B(n27982), .Z(n31123) );
  NOR U40951 ( .A(n31117), .B(n31123), .Z(n27984) );
  XOR U40952 ( .A(n31116), .B(n27984), .Z(n28101) );
  XOR U40953 ( .A(n28098), .B(n28101), .Z(n31130) );
  IV U40954 ( .A(n31130), .Z(n27992) );
  IV U40955 ( .A(n27985), .Z(n27987) );
  NOR U40956 ( .A(n27987), .B(n27986), .Z(n28100) );
  IV U40957 ( .A(n27988), .Z(n27990) );
  NOR U40958 ( .A(n27990), .B(n27989), .Z(n31129) );
  NOR U40959 ( .A(n28100), .B(n31129), .Z(n27991) );
  XOR U40960 ( .A(n27992), .B(n27991), .Z(n28097) );
  XOR U40961 ( .A(n28093), .B(n28097), .Z(n27993) );
  NOR U40962 ( .A(n27994), .B(n27993), .Z(n34306) );
  IV U40963 ( .A(n27995), .Z(n27997) );
  NOR U40964 ( .A(n27997), .B(n27996), .Z(n28095) );
  NOR U40965 ( .A(n28093), .B(n28095), .Z(n27998) );
  XOR U40966 ( .A(n28097), .B(n27998), .Z(n31135) );
  NOR U40967 ( .A(n27999), .B(n31135), .Z(n28000) );
  NOR U40968 ( .A(n34306), .B(n28000), .Z(n31140) );
  IV U40969 ( .A(n28001), .Z(n28002) );
  NOR U40970 ( .A(n28003), .B(n28002), .Z(n31134) );
  IV U40971 ( .A(n28004), .Z(n28005) );
  NOR U40972 ( .A(n28006), .B(n28005), .Z(n31139) );
  NOR U40973 ( .A(n31134), .B(n31139), .Z(n28007) );
  XOR U40974 ( .A(n31140), .B(n28007), .Z(n31223) );
  IV U40975 ( .A(n28008), .Z(n28009) );
  NOR U40976 ( .A(n28010), .B(n28009), .Z(n31226) );
  IV U40977 ( .A(n28011), .Z(n28012) );
  NOR U40978 ( .A(n28013), .B(n28012), .Z(n31222) );
  NOR U40979 ( .A(n31226), .B(n31222), .Z(n31138) );
  XOR U40980 ( .A(n31223), .B(n31138), .Z(n31145) );
  IV U40981 ( .A(n28014), .Z(n28015) );
  NOR U40982 ( .A(n28016), .B(n28015), .Z(n37721) );
  IV U40983 ( .A(n28017), .Z(n28018) );
  NOR U40984 ( .A(n28019), .B(n28018), .Z(n37730) );
  NOR U40985 ( .A(n37721), .B(n37730), .Z(n31146) );
  XOR U40986 ( .A(n31145), .B(n31146), .Z(n31153) );
  XOR U40987 ( .A(n28020), .B(n31153), .Z(n31150) );
  XOR U40988 ( .A(n31151), .B(n31150), .Z(n31213) );
  XOR U40989 ( .A(n31157), .B(n31213), .Z(n28091) );
  IV U40990 ( .A(n28021), .Z(n28022) );
  NOR U40991 ( .A(n28023), .B(n28022), .Z(n31158) );
  IV U40992 ( .A(n28024), .Z(n28025) );
  NOR U40993 ( .A(n28026), .B(n28025), .Z(n28090) );
  NOR U40994 ( .A(n31158), .B(n28090), .Z(n28027) );
  XOR U40995 ( .A(n28091), .B(n28027), .Z(n34344) );
  XOR U40996 ( .A(n31163), .B(n34344), .Z(n28028) );
  IV U40997 ( .A(n28028), .Z(n31167) );
  XOR U40998 ( .A(n31164), .B(n31167), .Z(n31173) );
  IV U40999 ( .A(n31173), .Z(n28036) );
  IV U41000 ( .A(n28029), .Z(n28031) );
  NOR U41001 ( .A(n28031), .B(n28030), .Z(n31166) );
  IV U41002 ( .A(n28032), .Z(n28034) );
  NOR U41003 ( .A(n28034), .B(n28033), .Z(n31172) );
  NOR U41004 ( .A(n31166), .B(n31172), .Z(n28035) );
  XOR U41005 ( .A(n28036), .B(n28035), .Z(n28089) );
  XOR U41006 ( .A(n28085), .B(n28089), .Z(n28083) );
  XOR U41007 ( .A(n28037), .B(n28083), .Z(n28038) );
  IV U41008 ( .A(n28038), .Z(n31179) );
  IV U41009 ( .A(n28039), .Z(n28041) );
  NOR U41010 ( .A(n28041), .B(n28040), .Z(n28042) );
  IV U41011 ( .A(n28042), .Z(n31178) );
  XOR U41012 ( .A(n31179), .B(n31178), .Z(n28043) );
  NOR U41013 ( .A(n28048), .B(n28043), .Z(n28050) );
  IV U41014 ( .A(n28044), .Z(n28046) );
  NOR U41015 ( .A(n28046), .B(n28045), .Z(n28047) );
  IV U41016 ( .A(n28047), .Z(n28054) );
  NOR U41017 ( .A(n28050), .B(n28054), .Z(n31192) );
  IV U41018 ( .A(n28048), .Z(n28049) );
  NOR U41019 ( .A(n31179), .B(n28049), .Z(n31197) );
  NOR U41020 ( .A(n28050), .B(n31197), .Z(n28051) );
  IV U41021 ( .A(n28051), .Z(n28081) );
  NOR U41022 ( .A(n28053), .B(n28052), .Z(n28055) );
  IV U41023 ( .A(n28055), .Z(n28080) );
  XOR U41024 ( .A(n28081), .B(n28080), .Z(n28057) );
  NOR U41025 ( .A(n28055), .B(n28054), .Z(n28056) );
  NOR U41026 ( .A(n28057), .B(n28056), .Z(n28058) );
  NOR U41027 ( .A(n31192), .B(n28058), .Z(n28059) );
  IV U41028 ( .A(n28059), .Z(n37970) );
  NOR U41029 ( .A(n28061), .B(n28060), .Z(n28065) );
  IV U41030 ( .A(n28061), .Z(n28063) );
  NOR U41031 ( .A(n28063), .B(n28062), .Z(n37973) );
  NOR U41032 ( .A(n37973), .B(n37962), .Z(n28064) );
  NOR U41033 ( .A(n28065), .B(n28064), .Z(n28075) );
  XOR U41034 ( .A(n37970), .B(n28075), .Z(n28079) );
  IV U41035 ( .A(n28066), .Z(n28068) );
  NOR U41036 ( .A(n28068), .B(n28067), .Z(n28077) );
  IV U41037 ( .A(n28069), .Z(n28071) );
  NOR U41038 ( .A(n28071), .B(n28070), .Z(n28073) );
  NOR U41039 ( .A(n28077), .B(n28073), .Z(n28072) );
  XOR U41040 ( .A(n28079), .B(n28072), .Z(n34378) );
  IV U41041 ( .A(n34378), .Z(n34376) );
  IV U41042 ( .A(n28073), .Z(n28074) );
  NOR U41043 ( .A(n28079), .B(n28074), .Z(n31189) );
  IV U41044 ( .A(n28075), .Z(n28076) );
  NOR U41045 ( .A(n37970), .B(n28076), .Z(n34367) );
  IV U41046 ( .A(n28077), .Z(n28078) );
  NOR U41047 ( .A(n28079), .B(n28078), .Z(n34369) );
  NOR U41048 ( .A(n34367), .B(n34369), .Z(n31182) );
  NOR U41049 ( .A(n28081), .B(n28080), .Z(n31194) );
  IV U41050 ( .A(n28082), .Z(n28084) );
  NOR U41051 ( .A(n28084), .B(n28083), .Z(n34357) );
  IV U41052 ( .A(n28085), .Z(n28086) );
  NOR U41053 ( .A(n28089), .B(n28086), .Z(n31205) );
  IV U41054 ( .A(n28087), .Z(n28088) );
  NOR U41055 ( .A(n28089), .B(n28088), .Z(n31199) );
  NOR U41056 ( .A(n31205), .B(n31199), .Z(n31176) );
  IV U41057 ( .A(n28090), .Z(n28092) );
  IV U41058 ( .A(n28091), .Z(n31159) );
  NOR U41059 ( .A(n28092), .B(n31159), .Z(n34340) );
  IV U41060 ( .A(n28093), .Z(n28094) );
  NOR U41061 ( .A(n28097), .B(n28094), .Z(n31237) );
  IV U41062 ( .A(n28095), .Z(n28096) );
  NOR U41063 ( .A(n28097), .B(n28096), .Z(n31232) );
  NOR U41064 ( .A(n31237), .B(n31232), .Z(n31132) );
  IV U41065 ( .A(n28098), .Z(n28099) );
  NOR U41066 ( .A(n28099), .B(n28101), .Z(n34291) );
  IV U41067 ( .A(n28100), .Z(n28102) );
  NOR U41068 ( .A(n28102), .B(n28101), .Z(n34302) );
  NOR U41069 ( .A(n34291), .B(n34302), .Z(n31128) );
  IV U41070 ( .A(n28103), .Z(n28105) );
  NOR U41071 ( .A(n28105), .B(n28104), .Z(n31240) );
  IV U41072 ( .A(n28106), .Z(n28109) );
  IV U41073 ( .A(n28107), .Z(n28113) );
  XOR U41074 ( .A(n28113), .B(n28110), .Z(n28108) );
  NOR U41075 ( .A(n28109), .B(n28108), .Z(n34259) );
  IV U41076 ( .A(n28110), .Z(n28114) );
  IV U41077 ( .A(n28111), .Z(n28112) );
  NOR U41078 ( .A(n28114), .B(n28112), .Z(n34256) );
  NOR U41079 ( .A(n28114), .B(n28113), .Z(n28116) );
  IV U41080 ( .A(n31246), .Z(n28115) );
  NOR U41081 ( .A(n28115), .B(n31107), .Z(n34253) );
  NOR U41082 ( .A(n28116), .B(n34253), .Z(n31243) );
  IV U41083 ( .A(n28117), .Z(n28119) );
  IV U41084 ( .A(n28118), .Z(n31087) );
  NOR U41085 ( .A(n28119), .B(n31087), .Z(n31099) );
  IV U41086 ( .A(n31099), .Z(n31085) );
  IV U41087 ( .A(n28120), .Z(n28126) );
  IV U41088 ( .A(n28121), .Z(n28122) );
  NOR U41089 ( .A(n28126), .B(n28122), .Z(n28123) );
  IV U41090 ( .A(n28123), .Z(n31259) );
  IV U41091 ( .A(n28124), .Z(n28125) );
  NOR U41092 ( .A(n28126), .B(n28125), .Z(n31266) );
  IV U41093 ( .A(n28127), .Z(n28128) );
  NOR U41094 ( .A(n28131), .B(n28128), .Z(n31269) );
  IV U41095 ( .A(n28129), .Z(n28130) );
  NOR U41096 ( .A(n28131), .B(n28130), .Z(n34236) );
  NOR U41097 ( .A(n31269), .B(n34236), .Z(n31081) );
  IV U41098 ( .A(n28132), .Z(n28134) );
  IV U41099 ( .A(n28133), .Z(n28137) );
  NOR U41100 ( .A(n28134), .B(n28137), .Z(n28135) );
  IV U41101 ( .A(n28135), .Z(n34232) );
  IV U41102 ( .A(n28136), .Z(n28138) );
  NOR U41103 ( .A(n28138), .B(n28137), .Z(n34229) );
  NOR U41104 ( .A(n28140), .B(n28139), .Z(n34225) );
  IV U41105 ( .A(n31077), .Z(n31068) );
  IV U41106 ( .A(n28141), .Z(n28142) );
  NOR U41107 ( .A(n28142), .B(n31056), .Z(n28143) );
  IV U41108 ( .A(n28143), .Z(n34219) );
  NOR U41109 ( .A(n28144), .B(n34196), .Z(n31042) );
  IV U41110 ( .A(n28145), .Z(n28150) );
  IV U41111 ( .A(n28146), .Z(n28147) );
  NOR U41112 ( .A(n28150), .B(n28147), .Z(n31037) );
  IV U41113 ( .A(n28148), .Z(n28149) );
  NOR U41114 ( .A(n28150), .B(n28149), .Z(n31034) );
  IV U41115 ( .A(n31034), .Z(n31029) );
  IV U41116 ( .A(n28151), .Z(n28152) );
  NOR U41117 ( .A(n28152), .B(n28155), .Z(n31308) );
  NOR U41118 ( .A(n28153), .B(n31315), .Z(n28157) );
  IV U41119 ( .A(n28154), .Z(n28156) );
  NOR U41120 ( .A(n28156), .B(n28155), .Z(n31311) );
  NOR U41121 ( .A(n28157), .B(n31311), .Z(n31014) );
  IV U41122 ( .A(n28158), .Z(n28160) );
  IV U41123 ( .A(n28159), .Z(n28162) );
  NOR U41124 ( .A(n28160), .B(n28162), .Z(n34185) );
  IV U41125 ( .A(n28161), .Z(n28163) );
  NOR U41126 ( .A(n28163), .B(n28162), .Z(n31319) );
  IV U41127 ( .A(n28164), .Z(n28165) );
  NOR U41128 ( .A(n28165), .B(n28167), .Z(n31321) );
  IV U41129 ( .A(n31321), .Z(n34178) );
  IV U41130 ( .A(n28166), .Z(n28168) );
  NOR U41131 ( .A(n28168), .B(n28167), .Z(n28169) );
  IV U41132 ( .A(n28169), .Z(n31323) );
  XOR U41133 ( .A(n34178), .B(n31323), .Z(n28170) );
  NOR U41134 ( .A(n31319), .B(n28170), .Z(n28171) );
  IV U41135 ( .A(n28171), .Z(n31013) );
  IV U41136 ( .A(n28172), .Z(n28177) );
  IV U41137 ( .A(n28173), .Z(n28174) );
  NOR U41138 ( .A(n28177), .B(n28174), .Z(n34174) );
  IV U41139 ( .A(n28175), .Z(n28176) );
  NOR U41140 ( .A(n28177), .B(n28176), .Z(n31327) );
  IV U41141 ( .A(n28178), .Z(n28180) );
  NOR U41142 ( .A(n28180), .B(n28179), .Z(n34167) );
  IV U41143 ( .A(n28181), .Z(n28182) );
  NOR U41144 ( .A(n28182), .B(n30999), .Z(n31332) );
  IV U41145 ( .A(n30980), .Z(n31337) );
  NOR U41146 ( .A(n30978), .B(n31337), .Z(n30982) );
  IV U41147 ( .A(n28183), .Z(n28184) );
  NOR U41148 ( .A(n30955), .B(n28184), .Z(n30968) );
  IV U41149 ( .A(n28185), .Z(n31342) );
  NOR U41150 ( .A(n31342), .B(n28186), .Z(n28189) );
  IV U41151 ( .A(n28187), .Z(n28188) );
  NOR U41152 ( .A(n28188), .B(n30959), .Z(n34134) );
  NOR U41153 ( .A(n28189), .B(n34134), .Z(n30952) );
  IV U41154 ( .A(n28190), .Z(n30937) );
  IV U41155 ( .A(n28191), .Z(n28192) );
  NOR U41156 ( .A(n30937), .B(n28192), .Z(n34124) );
  IV U41157 ( .A(n28193), .Z(n28195) );
  NOR U41158 ( .A(n28195), .B(n28194), .Z(n34121) );
  IV U41159 ( .A(n28196), .Z(n28197) );
  NOR U41160 ( .A(n28197), .B(n30932), .Z(n34583) );
  IV U41161 ( .A(n28198), .Z(n30927) );
  IV U41162 ( .A(n28199), .Z(n28200) );
  NOR U41163 ( .A(n30927), .B(n28200), .Z(n34588) );
  NOR U41164 ( .A(n34583), .B(n34588), .Z(n34116) );
  IV U41165 ( .A(n28201), .Z(n31367) );
  IV U41166 ( .A(n28202), .Z(n28203) );
  NOR U41167 ( .A(n31367), .B(n28203), .Z(n34598) );
  IV U41168 ( .A(n28204), .Z(n28205) );
  NOR U41169 ( .A(n28208), .B(n28205), .Z(n31395) );
  IV U41170 ( .A(n28206), .Z(n28207) );
  NOR U41171 ( .A(n28208), .B(n28207), .Z(n30872) );
  IV U41172 ( .A(n30872), .Z(n30864) );
  IV U41173 ( .A(n28209), .Z(n28210) );
  NOR U41174 ( .A(n28210), .B(n30841), .Z(n30848) );
  IV U41175 ( .A(n28211), .Z(n28212) );
  NOR U41176 ( .A(n30805), .B(n28212), .Z(n34074) );
  IV U41177 ( .A(n28213), .Z(n28215) );
  IV U41178 ( .A(n28214), .Z(n28217) );
  NOR U41179 ( .A(n28215), .B(n28217), .Z(n34071) );
  IV U41180 ( .A(n28216), .Z(n28218) );
  NOR U41181 ( .A(n28218), .B(n28217), .Z(n34067) );
  NOR U41182 ( .A(n28219), .B(n34067), .Z(n30802) );
  IV U41183 ( .A(n28220), .Z(n28221) );
  NOR U41184 ( .A(n28222), .B(n28221), .Z(n37545) );
  IV U41185 ( .A(n28223), .Z(n28224) );
  NOR U41186 ( .A(n28224), .B(n30799), .Z(n37540) );
  NOR U41187 ( .A(n37545), .B(n37540), .Z(n34059) );
  IV U41188 ( .A(n28225), .Z(n37527) );
  NOR U41189 ( .A(n28226), .B(n37527), .Z(n30796) );
  IV U41190 ( .A(n30796), .Z(n30788) );
  IV U41191 ( .A(n28227), .Z(n28228) );
  NOR U41192 ( .A(n28228), .B(n31426), .Z(n28229) );
  IV U41193 ( .A(n28229), .Z(n31433) );
  IV U41194 ( .A(n28230), .Z(n28236) );
  IV U41195 ( .A(n28231), .Z(n28232) );
  NOR U41196 ( .A(n28236), .B(n28232), .Z(n28233) );
  IV U41197 ( .A(n28233), .Z(n34690) );
  IV U41198 ( .A(n28234), .Z(n28235) );
  NOR U41199 ( .A(n28236), .B(n28235), .Z(n31435) );
  IV U41200 ( .A(n28237), .Z(n28239) );
  NOR U41201 ( .A(n28239), .B(n28238), .Z(n34039) );
  IV U41202 ( .A(n28240), .Z(n28242) );
  IV U41203 ( .A(n28241), .Z(n28244) );
  NOR U41204 ( .A(n28242), .B(n28244), .Z(n34033) );
  NOR U41205 ( .A(n34039), .B(n34033), .Z(n30765) );
  NOR U41206 ( .A(n31438), .B(n28243), .Z(n28246) );
  NOR U41207 ( .A(n28245), .B(n28244), .Z(n34034) );
  NOR U41208 ( .A(n28246), .B(n34034), .Z(n30764) );
  IV U41209 ( .A(n28247), .Z(n28249) );
  IV U41210 ( .A(n28248), .Z(n30762) );
  NOR U41211 ( .A(n28249), .B(n30762), .Z(n31448) );
  IV U41212 ( .A(n28250), .Z(n28251) );
  NOR U41213 ( .A(n28254), .B(n28251), .Z(n30757) );
  IV U41214 ( .A(n28252), .Z(n28253) );
  NOR U41215 ( .A(n28254), .B(n28253), .Z(n30755) );
  IV U41216 ( .A(n30755), .Z(n30746) );
  IV U41217 ( .A(n28255), .Z(n28258) );
  IV U41218 ( .A(n28256), .Z(n28257) );
  NOR U41219 ( .A(n28258), .B(n28257), .Z(n30742) );
  IV U41220 ( .A(n28259), .Z(n28260) );
  NOR U41221 ( .A(n28260), .B(n30732), .Z(n30736) );
  IV U41222 ( .A(n30736), .Z(n30728) );
  IV U41223 ( .A(n28261), .Z(n28263) );
  NOR U41224 ( .A(n28263), .B(n28262), .Z(n31460) );
  IV U41225 ( .A(n28264), .Z(n28265) );
  NOR U41226 ( .A(n28265), .B(n28267), .Z(n31471) );
  IV U41227 ( .A(n28266), .Z(n28268) );
  NOR U41228 ( .A(n28268), .B(n28267), .Z(n31468) );
  IV U41229 ( .A(n28269), .Z(n28271) );
  IV U41230 ( .A(n28270), .Z(n28274) );
  NOR U41231 ( .A(n28271), .B(n28274), .Z(n31481) );
  NOR U41232 ( .A(n28272), .B(n31492), .Z(n28276) );
  IV U41233 ( .A(n28273), .Z(n28275) );
  NOR U41234 ( .A(n28275), .B(n28274), .Z(n31487) );
  NOR U41235 ( .A(n28276), .B(n31487), .Z(n30720) );
  NOR U41236 ( .A(n28277), .B(n34009), .Z(n28278) );
  IV U41237 ( .A(n28278), .Z(n31498) );
  IV U41238 ( .A(n28279), .Z(n28281) );
  IV U41239 ( .A(n28280), .Z(n30699) );
  NOR U41240 ( .A(n28281), .B(n30699), .Z(n34000) );
  IV U41241 ( .A(n28282), .Z(n28283) );
  NOR U41242 ( .A(n28283), .B(n28286), .Z(n28284) );
  IV U41243 ( .A(n28284), .Z(n31546) );
  IV U41244 ( .A(n28285), .Z(n28287) );
  NOR U41245 ( .A(n28287), .B(n28286), .Z(n31548) );
  IV U41246 ( .A(n28288), .Z(n28293) );
  IV U41247 ( .A(n28289), .Z(n28290) );
  NOR U41248 ( .A(n28293), .B(n28290), .Z(n31554) );
  NOR U41249 ( .A(n31548), .B(n31554), .Z(n30689) );
  IV U41250 ( .A(n28291), .Z(n28292) );
  NOR U41251 ( .A(n28293), .B(n28292), .Z(n31557) );
  NOR U41252 ( .A(n33992), .B(n28294), .Z(n28298) );
  IV U41253 ( .A(n28295), .Z(n28296) );
  NOR U41254 ( .A(n28296), .B(n31551), .Z(n28297) );
  NOR U41255 ( .A(n28298), .B(n28297), .Z(n30688) );
  IV U41256 ( .A(n28299), .Z(n28300) );
  NOR U41257 ( .A(n28303), .B(n28300), .Z(n33989) );
  IV U41258 ( .A(n28301), .Z(n28302) );
  NOR U41259 ( .A(n28303), .B(n28302), .Z(n33987) );
  IV U41260 ( .A(n28304), .Z(n28306) );
  IV U41261 ( .A(n28305), .Z(n28309) );
  NOR U41262 ( .A(n28306), .B(n28309), .Z(n28307) );
  IV U41263 ( .A(n28307), .Z(n33979) );
  IV U41264 ( .A(n28308), .Z(n28310) );
  NOR U41265 ( .A(n28310), .B(n28309), .Z(n28311) );
  IV U41266 ( .A(n28311), .Z(n31566) );
  XOR U41267 ( .A(n33979), .B(n31566), .Z(n28312) );
  NOR U41268 ( .A(n33987), .B(n28312), .Z(n30687) );
  IV U41269 ( .A(n28313), .Z(n28319) );
  IV U41270 ( .A(n28314), .Z(n28315) );
  NOR U41271 ( .A(n28319), .B(n28315), .Z(n34763) );
  NOR U41272 ( .A(n28316), .B(n34760), .Z(n33981) );
  NOR U41273 ( .A(n34763), .B(n33981), .Z(n30686) );
  IV U41274 ( .A(n28317), .Z(n28318) );
  NOR U41275 ( .A(n28319), .B(n28318), .Z(n34769) );
  IV U41276 ( .A(n28320), .Z(n28321) );
  NOR U41277 ( .A(n28321), .B(n28325), .Z(n31571) );
  NOR U41278 ( .A(n34769), .B(n31571), .Z(n30685) );
  IV U41279 ( .A(n28322), .Z(n31574) );
  NOR U41280 ( .A(n28323), .B(n31574), .Z(n28327) );
  IV U41281 ( .A(n28324), .Z(n28326) );
  NOR U41282 ( .A(n28326), .B(n28325), .Z(n31567) );
  NOR U41283 ( .A(n28327), .B(n31567), .Z(n30684) );
  IV U41284 ( .A(n28328), .Z(n28330) );
  IV U41285 ( .A(n28329), .Z(n30676) );
  NOR U41286 ( .A(n28330), .B(n30676), .Z(n30670) );
  IV U41287 ( .A(n28331), .Z(n28332) );
  NOR U41288 ( .A(n28332), .B(n30660), .Z(n30668) );
  IV U41289 ( .A(n30668), .Z(n30658) );
  IV U41290 ( .A(n28333), .Z(n30653) );
  IV U41291 ( .A(n28334), .Z(n28335) );
  NOR U41292 ( .A(n30653), .B(n28335), .Z(n30655) );
  IV U41293 ( .A(n30655), .Z(n30650) );
  IV U41294 ( .A(n28336), .Z(n28338) );
  NOR U41295 ( .A(n28338), .B(n28337), .Z(n33950) );
  IV U41296 ( .A(n28339), .Z(n28341) );
  IV U41297 ( .A(n28340), .Z(n28342) );
  NOR U41298 ( .A(n28341), .B(n28342), .Z(n33947) );
  NOR U41299 ( .A(n28343), .B(n28342), .Z(n38343) );
  NOR U41300 ( .A(n38348), .B(n38343), .Z(n34792) );
  IV U41301 ( .A(n28344), .Z(n28345) );
  NOR U41302 ( .A(n28345), .B(n28347), .Z(n33938) );
  IV U41303 ( .A(n28346), .Z(n28348) );
  NOR U41304 ( .A(n28348), .B(n28347), .Z(n33942) );
  IV U41305 ( .A(n28349), .Z(n33931) );
  NOR U41306 ( .A(n28350), .B(n33931), .Z(n28351) );
  NOR U41307 ( .A(n33942), .B(n28351), .Z(n28352) );
  IV U41308 ( .A(n28352), .Z(n28353) );
  NOR U41309 ( .A(n33938), .B(n28353), .Z(n30648) );
  IV U41310 ( .A(n28354), .Z(n28356) );
  IV U41311 ( .A(n28355), .Z(n28359) );
  NOR U41312 ( .A(n28356), .B(n28359), .Z(n33919) );
  NOR U41313 ( .A(n28357), .B(n33908), .Z(n28361) );
  IV U41314 ( .A(n28358), .Z(n28360) );
  NOR U41315 ( .A(n28360), .B(n28359), .Z(n33914) );
  NOR U41316 ( .A(n28361), .B(n33914), .Z(n30636) );
  IV U41317 ( .A(n28362), .Z(n31588) );
  NOR U41318 ( .A(n28363), .B(n31588), .Z(n31580) );
  IV U41319 ( .A(n28364), .Z(n28365) );
  NOR U41320 ( .A(n28365), .B(n30632), .Z(n31584) );
  IV U41321 ( .A(n28366), .Z(n34823) );
  NOR U41322 ( .A(n28367), .B(n34823), .Z(n33897) );
  NOR U41323 ( .A(n28368), .B(n31605), .Z(n28369) );
  NOR U41324 ( .A(n33897), .B(n28369), .Z(n30628) );
  NOR U41325 ( .A(n28370), .B(n37298), .Z(n33898) );
  IV U41326 ( .A(n28371), .Z(n28372) );
  NOR U41327 ( .A(n28372), .B(n28374), .Z(n33872) );
  IV U41328 ( .A(n28373), .Z(n28375) );
  NOR U41329 ( .A(n28375), .B(n28374), .Z(n30597) );
  IV U41330 ( .A(n28376), .Z(n34855) );
  NOR U41331 ( .A(n28377), .B(n34855), .Z(n30594) );
  IV U41332 ( .A(n30594), .Z(n30582) );
  IV U41333 ( .A(n28378), .Z(n28379) );
  NOR U41334 ( .A(n28380), .B(n28379), .Z(n28381) );
  IV U41335 ( .A(n28381), .Z(n33870) );
  NOR U41336 ( .A(n31617), .B(n31619), .Z(n30581) );
  IV U41337 ( .A(n28382), .Z(n28383) );
  NOR U41338 ( .A(n28383), .B(n28384), .Z(n31622) );
  NOR U41339 ( .A(n28385), .B(n28384), .Z(n31624) );
  NOR U41340 ( .A(n31622), .B(n31624), .Z(n28386) );
  IV U41341 ( .A(n28386), .Z(n28389) );
  NOR U41342 ( .A(n31628), .B(n28387), .Z(n28388) );
  NOR U41343 ( .A(n28389), .B(n28388), .Z(n30580) );
  IV U41344 ( .A(n28390), .Z(n28392) );
  NOR U41345 ( .A(n28392), .B(n28391), .Z(n31632) );
  IV U41346 ( .A(n28393), .Z(n28394) );
  NOR U41347 ( .A(n28394), .B(n28397), .Z(n28395) );
  IV U41348 ( .A(n28395), .Z(n33850) );
  IV U41349 ( .A(n28396), .Z(n28398) );
  NOR U41350 ( .A(n28398), .B(n28397), .Z(n31636) );
  IV U41351 ( .A(n28399), .Z(n28400) );
  NOR U41352 ( .A(n28400), .B(n31639), .Z(n28401) );
  NOR U41353 ( .A(n31636), .B(n28401), .Z(n30579) );
  IV U41354 ( .A(n28402), .Z(n31645) );
  NOR U41355 ( .A(n31645), .B(n28403), .Z(n28406) );
  IV U41356 ( .A(n28404), .Z(n28405) );
  NOR U41357 ( .A(n28405), .B(n31639), .Z(n34872) );
  NOR U41358 ( .A(n28406), .B(n34872), .Z(n28407) );
  IV U41359 ( .A(n28407), .Z(n37245) );
  IV U41360 ( .A(n28408), .Z(n28410) );
  NOR U41361 ( .A(n28410), .B(n28409), .Z(n31654) );
  IV U41362 ( .A(n28411), .Z(n28412) );
  NOR U41363 ( .A(n28412), .B(n28414), .Z(n33823) );
  IV U41364 ( .A(n28413), .Z(n28415) );
  NOR U41365 ( .A(n28415), .B(n28414), .Z(n33827) );
  NOR U41366 ( .A(n33823), .B(n33827), .Z(n31659) );
  IV U41367 ( .A(n28416), .Z(n30527) );
  IV U41368 ( .A(n28417), .Z(n28418) );
  NOR U41369 ( .A(n30527), .B(n28418), .Z(n31666) );
  IV U41370 ( .A(n28419), .Z(n28421) );
  NOR U41371 ( .A(n28421), .B(n28420), .Z(n31672) );
  NOR U41372 ( .A(n31666), .B(n31672), .Z(n30518) );
  NOR U41373 ( .A(n28423), .B(n28422), .Z(n31679) );
  NOR U41374 ( .A(n28425), .B(n28424), .Z(n33787) );
  IV U41375 ( .A(n28426), .Z(n28428) );
  IV U41376 ( .A(n28427), .Z(n30472) );
  NOR U41377 ( .A(n28428), .B(n30472), .Z(n30469) );
  IV U41378 ( .A(n30469), .Z(n30454) );
  IV U41379 ( .A(n28429), .Z(n34993) );
  NOR U41380 ( .A(n34993), .B(n28430), .Z(n30447) );
  IV U41381 ( .A(n30447), .Z(n30434) );
  IV U41382 ( .A(n28431), .Z(n31705) );
  NOR U41383 ( .A(n28432), .B(n31705), .Z(n30433) );
  NOR U41384 ( .A(n30428), .B(n28433), .Z(n30418) );
  IV U41385 ( .A(n28434), .Z(n28435) );
  NOR U41386 ( .A(n28435), .B(n28437), .Z(n31712) );
  IV U41387 ( .A(n28436), .Z(n28438) );
  NOR U41388 ( .A(n28438), .B(n28437), .Z(n33745) );
  NOR U41389 ( .A(n31712), .B(n33745), .Z(n30405) );
  IV U41390 ( .A(n28439), .Z(n28447) );
  IV U41391 ( .A(n28440), .Z(n28441) );
  NOR U41392 ( .A(n28447), .B(n28441), .Z(n33742) );
  IV U41393 ( .A(n28442), .Z(n28444) );
  NOR U41394 ( .A(n28444), .B(n28443), .Z(n31719) );
  NOR U41395 ( .A(n33742), .B(n31719), .Z(n30404) );
  IV U41396 ( .A(n28445), .Z(n28446) );
  NOR U41397 ( .A(n28447), .B(n28446), .Z(n31717) );
  IV U41398 ( .A(n28448), .Z(n30398) );
  IV U41399 ( .A(n28449), .Z(n28450) );
  NOR U41400 ( .A(n30398), .B(n28450), .Z(n30390) );
  IV U41401 ( .A(n28451), .Z(n28453) );
  NOR U41402 ( .A(n28453), .B(n28452), .Z(n33731) );
  IV U41403 ( .A(n28454), .Z(n28456) );
  NOR U41404 ( .A(n28456), .B(n28455), .Z(n33700) );
  IV U41405 ( .A(n28457), .Z(n28458) );
  NOR U41406 ( .A(n28458), .B(n28460), .Z(n35062) );
  IV U41407 ( .A(n28459), .Z(n28461) );
  NOR U41408 ( .A(n28461), .B(n28460), .Z(n35057) );
  NOR U41409 ( .A(n35062), .B(n35057), .Z(n33698) );
  IV U41410 ( .A(n33698), .Z(n28463) );
  NOR U41411 ( .A(n28462), .B(n37111), .Z(n33695) );
  NOR U41412 ( .A(n28463), .B(n33695), .Z(n30347) );
  IV U41413 ( .A(n28464), .Z(n28466) );
  IV U41414 ( .A(n28465), .Z(n30345) );
  NOR U41415 ( .A(n28466), .B(n30345), .Z(n30341) );
  IV U41416 ( .A(n30341), .Z(n30336) );
  IV U41417 ( .A(n28467), .Z(n28468) );
  NOR U41418 ( .A(n28468), .B(n28470), .Z(n30314) );
  IV U41419 ( .A(n28469), .Z(n28471) );
  NOR U41420 ( .A(n28471), .B(n28470), .Z(n30312) );
  IV U41421 ( .A(n30312), .Z(n30307) );
  NOR U41422 ( .A(n28472), .B(n37076), .Z(n31745) );
  IV U41423 ( .A(n28473), .Z(n28474) );
  NOR U41424 ( .A(n28474), .B(n30300), .Z(n33665) );
  IV U41425 ( .A(n28475), .Z(n33654) );
  NOR U41426 ( .A(n33654), .B(n28476), .Z(n33659) );
  IV U41427 ( .A(n28477), .Z(n28478) );
  NOR U41428 ( .A(n28478), .B(n28481), .Z(n28479) );
  IV U41429 ( .A(n28479), .Z(n31752) );
  IV U41430 ( .A(n28480), .Z(n28482) );
  NOR U41431 ( .A(n28482), .B(n28481), .Z(n28483) );
  IV U41432 ( .A(n28483), .Z(n33649) );
  XOR U41433 ( .A(n31752), .B(n33649), .Z(n28484) );
  NOR U41434 ( .A(n33659), .B(n28484), .Z(n30298) );
  IV U41435 ( .A(n28485), .Z(n30289) );
  NOR U41436 ( .A(n28486), .B(n30289), .Z(n30285) );
  IV U41437 ( .A(n28487), .Z(n28488) );
  NOR U41438 ( .A(n28491), .B(n28488), .Z(n31760) );
  IV U41439 ( .A(n28489), .Z(n28490) );
  NOR U41440 ( .A(n28491), .B(n28490), .Z(n31759) );
  NOR U41441 ( .A(n31760), .B(n31759), .Z(n30271) );
  IV U41442 ( .A(n28492), .Z(n28495) );
  IV U41443 ( .A(n28493), .Z(n28494) );
  NOR U41444 ( .A(n28495), .B(n28494), .Z(n31763) );
  IV U41445 ( .A(n28496), .Z(n28499) );
  IV U41446 ( .A(n28497), .Z(n28498) );
  NOR U41447 ( .A(n28499), .B(n28498), .Z(n33614) );
  IV U41448 ( .A(n28500), .Z(n28501) );
  NOR U41449 ( .A(n28501), .B(n28506), .Z(n28502) );
  IV U41450 ( .A(n28502), .Z(n31772) );
  IV U41451 ( .A(n28503), .Z(n35124) );
  NOR U41452 ( .A(n28504), .B(n35124), .Z(n28508) );
  IV U41453 ( .A(n28505), .Z(n28507) );
  NOR U41454 ( .A(n28507), .B(n28506), .Z(n35117) );
  NOR U41455 ( .A(n28508), .B(n35117), .Z(n31769) );
  IV U41456 ( .A(n28509), .Z(n31782) );
  NOR U41457 ( .A(n31784), .B(n31782), .Z(n28512) );
  NOR U41458 ( .A(n28510), .B(n31775), .Z(n28511) );
  NOR U41459 ( .A(n28512), .B(n28511), .Z(n30270) );
  IV U41460 ( .A(n28513), .Z(n28515) );
  NOR U41461 ( .A(n28515), .B(n28514), .Z(n33599) );
  NOR U41462 ( .A(n28516), .B(n31786), .Z(n28517) );
  NOR U41463 ( .A(n33599), .B(n28517), .Z(n30269) );
  NOR U41464 ( .A(n28518), .B(n31792), .Z(n28522) );
  IV U41465 ( .A(n28519), .Z(n33585) );
  NOR U41466 ( .A(n28520), .B(n33585), .Z(n28521) );
  NOR U41467 ( .A(n28522), .B(n28521), .Z(n30268) );
  IV U41468 ( .A(n28523), .Z(n28525) );
  NOR U41469 ( .A(n28525), .B(n28524), .Z(n30252) );
  IV U41470 ( .A(n30252), .Z(n30235) );
  IV U41471 ( .A(n28526), .Z(n28527) );
  NOR U41472 ( .A(n28527), .B(n30232), .Z(n30229) );
  IV U41473 ( .A(n30229), .Z(n30212) );
  IV U41474 ( .A(n28528), .Z(n28530) );
  IV U41475 ( .A(n28529), .Z(n30209) );
  NOR U41476 ( .A(n28530), .B(n30209), .Z(n30201) );
  IV U41477 ( .A(n28531), .Z(n30187) );
  IV U41478 ( .A(n28532), .Z(n28533) );
  NOR U41479 ( .A(n28533), .B(n28536), .Z(n33556) );
  IV U41480 ( .A(n33563), .Z(n28534) );
  NOR U41481 ( .A(n28534), .B(n30181), .Z(n31808) );
  IV U41482 ( .A(n28535), .Z(n28537) );
  NOR U41483 ( .A(n28537), .B(n28536), .Z(n28538) );
  NOR U41484 ( .A(n31808), .B(n28538), .Z(n33559) );
  NOR U41485 ( .A(n28540), .B(n28539), .Z(n33539) );
  IV U41486 ( .A(n28541), .Z(n30174) );
  IV U41487 ( .A(n28542), .Z(n28543) );
  NOR U41488 ( .A(n30174), .B(n28543), .Z(n31820) );
  IV U41489 ( .A(n28544), .Z(n28546) );
  NOR U41490 ( .A(n28546), .B(n28545), .Z(n31822) );
  NOR U41491 ( .A(n31820), .B(n31822), .Z(n30171) );
  IV U41492 ( .A(n28547), .Z(n28548) );
  NOR U41493 ( .A(n28551), .B(n28548), .Z(n31828) );
  IV U41494 ( .A(n28549), .Z(n28550) );
  NOR U41495 ( .A(n28551), .B(n28550), .Z(n31826) );
  NOR U41496 ( .A(n31828), .B(n31826), .Z(n30170) );
  NOR U41497 ( .A(n28552), .B(n33526), .Z(n33517) );
  IV U41498 ( .A(n28553), .Z(n28555) );
  IV U41499 ( .A(n28554), .Z(n30166) );
  NOR U41500 ( .A(n28555), .B(n30166), .Z(n33536) );
  NOR U41501 ( .A(n33517), .B(n33536), .Z(n30169) );
  IV U41502 ( .A(n28556), .Z(n31834) );
  NOR U41503 ( .A(n28557), .B(n31834), .Z(n30164) );
  IV U41504 ( .A(n28558), .Z(n28559) );
  NOR U41505 ( .A(n28559), .B(n33502), .Z(n31839) );
  NOR U41506 ( .A(n28560), .B(n33510), .Z(n28561) );
  NOR U41507 ( .A(n31839), .B(n28561), .Z(n30163) );
  NOR U41508 ( .A(n28562), .B(n31849), .Z(n33500) );
  IV U41509 ( .A(n28563), .Z(n31842) );
  NOR U41510 ( .A(n28564), .B(n31842), .Z(n28565) );
  NOR U41511 ( .A(n33500), .B(n28565), .Z(n30162) );
  NOR U41512 ( .A(n28566), .B(n33483), .Z(n28569) );
  NOR U41513 ( .A(n31857), .B(n28567), .Z(n28568) );
  NOR U41514 ( .A(n28569), .B(n28568), .Z(n30161) );
  IV U41515 ( .A(n28570), .Z(n28572) );
  IV U41516 ( .A(n28571), .Z(n28573) );
  NOR U41517 ( .A(n28572), .B(n28573), .Z(n30148) );
  NOR U41518 ( .A(n28574), .B(n28573), .Z(n28575) );
  NOR U41519 ( .A(n33474), .B(n28575), .Z(n31868) );
  IV U41520 ( .A(n28576), .Z(n28577) );
  NOR U41521 ( .A(n28577), .B(n28579), .Z(n31873) );
  IV U41522 ( .A(n28578), .Z(n28580) );
  NOR U41523 ( .A(n28580), .B(n28579), .Z(n31872) );
  NOR U41524 ( .A(n31873), .B(n31872), .Z(n30147) );
  NOR U41525 ( .A(n28581), .B(n33461), .Z(n28584) );
  IV U41526 ( .A(n28582), .Z(n31877) );
  NOR U41527 ( .A(n31879), .B(n31877), .Z(n28583) );
  NOR U41528 ( .A(n28584), .B(n28583), .Z(n30146) );
  IV U41529 ( .A(n28585), .Z(n31880) );
  NOR U41530 ( .A(n28586), .B(n31880), .Z(n33454) );
  NOR U41531 ( .A(n28588), .B(n28587), .Z(n33442) );
  IV U41532 ( .A(n28589), .Z(n28591) );
  NOR U41533 ( .A(n28591), .B(n28590), .Z(n31899) );
  IV U41534 ( .A(n28592), .Z(n36828) );
  NOR U41535 ( .A(n28593), .B(n36828), .Z(n30102) );
  IV U41536 ( .A(n33419), .Z(n28594) );
  NOR U41537 ( .A(n28595), .B(n28594), .Z(n30094) );
  IV U41538 ( .A(n30094), .Z(n30089) );
  IV U41539 ( .A(n28596), .Z(n30081) );
  IV U41540 ( .A(n30080), .Z(n30077) );
  NOR U41541 ( .A(n30081), .B(n30077), .Z(n30074) );
  IV U41542 ( .A(n30074), .Z(n30068) );
  IV U41543 ( .A(n28597), .Z(n31920) );
  NOR U41544 ( .A(n28598), .B(n31920), .Z(n30067) );
  NOR U41545 ( .A(n28600), .B(n28599), .Z(n31926) );
  IV U41546 ( .A(n28601), .Z(n28602) );
  NOR U41547 ( .A(n28602), .B(n28605), .Z(n31932) );
  NOR U41548 ( .A(n31932), .B(n31930), .Z(n28603) );
  IV U41549 ( .A(n28603), .Z(n28607) );
  IV U41550 ( .A(n28604), .Z(n28606) );
  NOR U41551 ( .A(n28606), .B(n28605), .Z(n31934) );
  NOR U41552 ( .A(n28607), .B(n31934), .Z(n30066) );
  NOR U41553 ( .A(n35288), .B(n28608), .Z(n31941) );
  IV U41554 ( .A(n28609), .Z(n31938) );
  NOR U41555 ( .A(n31940), .B(n31938), .Z(n28610) );
  NOR U41556 ( .A(n31941), .B(n28610), .Z(n30065) );
  IV U41557 ( .A(n28611), .Z(n28613) );
  IV U41558 ( .A(n28612), .Z(n30063) );
  NOR U41559 ( .A(n28613), .B(n30063), .Z(n33376) );
  IV U41560 ( .A(n28614), .Z(n28615) );
  NOR U41561 ( .A(n28615), .B(n30021), .Z(n30018) );
  IV U41562 ( .A(n30018), .Z(n30013) );
  IV U41563 ( .A(n28616), .Z(n28618) );
  IV U41564 ( .A(n28617), .Z(n30003) );
  NOR U41565 ( .A(n28618), .B(n30003), .Z(n28619) );
  IV U41566 ( .A(n28619), .Z(n29999) );
  IV U41567 ( .A(n28620), .Z(n28621) );
  NOR U41568 ( .A(n28621), .B(n29979), .Z(n28622) );
  IV U41569 ( .A(n28622), .Z(n31989) );
  IV U41570 ( .A(n28623), .Z(n28625) );
  IV U41571 ( .A(n28624), .Z(n29973) );
  NOR U41572 ( .A(n28625), .B(n29973), .Z(n29970) );
  IV U41573 ( .A(n29970), .Z(n29966) );
  IV U41574 ( .A(n28626), .Z(n28631) );
  IV U41575 ( .A(n28627), .Z(n28628) );
  NOR U41576 ( .A(n28631), .B(n28628), .Z(n32005) );
  IV U41577 ( .A(n28629), .Z(n28630) );
  NOR U41578 ( .A(n28631), .B(n28630), .Z(n29963) );
  IV U41579 ( .A(n29963), .Z(n29952) );
  IV U41580 ( .A(n28632), .Z(n36704) );
  NOR U41581 ( .A(n36704), .B(n28633), .Z(n29959) );
  IV U41582 ( .A(n29959), .Z(n32010) );
  IV U41583 ( .A(n28634), .Z(n28635) );
  NOR U41584 ( .A(n28635), .B(n28637), .Z(n33316) );
  IV U41585 ( .A(n28636), .Z(n28638) );
  NOR U41586 ( .A(n28638), .B(n28637), .Z(n33311) );
  NOR U41587 ( .A(n33316), .B(n33311), .Z(n29950) );
  IV U41588 ( .A(n28639), .Z(n29929) );
  IV U41589 ( .A(n28640), .Z(n28641) );
  NOR U41590 ( .A(n29929), .B(n28641), .Z(n32023) );
  NOR U41591 ( .A(n28643), .B(n28642), .Z(n28644) );
  IV U41592 ( .A(n28644), .Z(n36666) );
  NOR U41593 ( .A(n28645), .B(n36666), .Z(n33305) );
  NOR U41594 ( .A(n32023), .B(n33305), .Z(n29923) );
  IV U41595 ( .A(n28646), .Z(n28648) );
  NOR U41596 ( .A(n28648), .B(n28647), .Z(n29830) );
  IV U41597 ( .A(n29830), .Z(n29828) );
  IV U41598 ( .A(n28649), .Z(n28650) );
  NOR U41599 ( .A(n28650), .B(n29824), .Z(n32081) );
  IV U41600 ( .A(n28651), .Z(n28653) );
  NOR U41601 ( .A(n28653), .B(n28652), .Z(n32095) );
  IV U41602 ( .A(n28654), .Z(n28655) );
  NOR U41603 ( .A(n28655), .B(n28657), .Z(n32101) );
  IV U41604 ( .A(n28656), .Z(n28658) );
  NOR U41605 ( .A(n28658), .B(n28657), .Z(n32103) );
  NOR U41606 ( .A(n32101), .B(n32103), .Z(n28659) );
  IV U41607 ( .A(n28659), .Z(n28662) );
  IV U41608 ( .A(n28660), .Z(n28661) );
  NOR U41609 ( .A(n28661), .B(n28664), .Z(n36583) );
  NOR U41610 ( .A(n28662), .B(n36583), .Z(n29800) );
  IV U41611 ( .A(n28663), .Z(n28665) );
  NOR U41612 ( .A(n28665), .B(n28664), .Z(n36576) );
  IV U41613 ( .A(n28666), .Z(n28668) );
  IV U41614 ( .A(n28667), .Z(n29793) );
  NOR U41615 ( .A(n28668), .B(n29793), .Z(n32109) );
  IV U41616 ( .A(n32109), .Z(n32107) );
  IV U41617 ( .A(n28669), .Z(n28672) );
  IV U41618 ( .A(n28670), .Z(n28671) );
  NOR U41619 ( .A(n28672), .B(n28671), .Z(n32116) );
  IV U41620 ( .A(n28673), .Z(n28674) );
  NOR U41621 ( .A(n28674), .B(n28676), .Z(n32122) );
  IV U41622 ( .A(n28675), .Z(n28677) );
  NOR U41623 ( .A(n28677), .B(n28676), .Z(n32124) );
  IV U41624 ( .A(n28678), .Z(n32128) );
  NOR U41625 ( .A(n32128), .B(n28679), .Z(n28680) );
  NOR U41626 ( .A(n32124), .B(n28680), .Z(n28681) );
  IV U41627 ( .A(n28681), .Z(n28682) );
  NOR U41628 ( .A(n32122), .B(n28682), .Z(n29784) );
  IV U41629 ( .A(n28683), .Z(n28685) );
  NOR U41630 ( .A(n28685), .B(n28684), .Z(n33204) );
  IV U41631 ( .A(n28686), .Z(n28687) );
  NOR U41632 ( .A(n28687), .B(n29782), .Z(n33201) );
  IV U41633 ( .A(n28688), .Z(n28695) );
  IV U41634 ( .A(n28689), .Z(n28690) );
  NOR U41635 ( .A(n28695), .B(n28690), .Z(n32143) );
  IV U41636 ( .A(n28691), .Z(n28692) );
  NOR U41637 ( .A(n28692), .B(n29765), .Z(n32141) );
  NOR U41638 ( .A(n32143), .B(n32141), .Z(n29761) );
  IV U41639 ( .A(n28693), .Z(n28694) );
  NOR U41640 ( .A(n28695), .B(n28694), .Z(n32146) );
  IV U41641 ( .A(n28696), .Z(n28698) );
  NOR U41642 ( .A(n28698), .B(n28697), .Z(n32149) );
  NOR U41643 ( .A(n32146), .B(n32149), .Z(n29760) );
  IV U41644 ( .A(n28699), .Z(n33158) );
  NOR U41645 ( .A(n33158), .B(n28700), .Z(n28703) );
  IV U41646 ( .A(n28701), .Z(n28702) );
  NOR U41647 ( .A(n28702), .B(n28705), .Z(n32153) );
  NOR U41648 ( .A(n28703), .B(n32153), .Z(n29759) );
  IV U41649 ( .A(n28704), .Z(n28706) );
  NOR U41650 ( .A(n28706), .B(n28705), .Z(n28707) );
  IV U41651 ( .A(n28707), .Z(n32152) );
  IV U41652 ( .A(n28708), .Z(n28710) );
  NOR U41653 ( .A(n28710), .B(n28709), .Z(n33162) );
  IV U41654 ( .A(n28711), .Z(n28713) );
  IV U41655 ( .A(n28712), .Z(n28715) );
  NOR U41656 ( .A(n28713), .B(n28715), .Z(n28714) );
  IV U41657 ( .A(n28714), .Z(n32157) );
  NOR U41658 ( .A(n28716), .B(n28715), .Z(n32155) );
  IV U41659 ( .A(n32155), .Z(n33150) );
  XOR U41660 ( .A(n32157), .B(n33150), .Z(n28717) );
  NOR U41661 ( .A(n33162), .B(n28717), .Z(n29757) );
  NOR U41662 ( .A(n28718), .B(n32161), .Z(n28722) );
  IV U41663 ( .A(n28719), .Z(n29751) );
  IV U41664 ( .A(n28720), .Z(n28721) );
  NOR U41665 ( .A(n29751), .B(n28721), .Z(n32166) );
  NOR U41666 ( .A(n28722), .B(n32166), .Z(n29756) );
  IV U41667 ( .A(n28723), .Z(n28724) );
  NOR U41668 ( .A(n29748), .B(n28724), .Z(n33141) );
  IV U41669 ( .A(n28725), .Z(n28726) );
  NOR U41670 ( .A(n28726), .B(n28731), .Z(n33131) );
  IV U41671 ( .A(n28727), .Z(n28729) );
  IV U41672 ( .A(n28728), .Z(n28734) );
  NOR U41673 ( .A(n28729), .B(n28734), .Z(n32173) );
  IV U41674 ( .A(n28730), .Z(n28732) );
  NOR U41675 ( .A(n28732), .B(n28731), .Z(n33134) );
  NOR U41676 ( .A(n32173), .B(n33134), .Z(n29745) );
  IV U41677 ( .A(n28733), .Z(n28735) );
  NOR U41678 ( .A(n28735), .B(n28734), .Z(n29743) );
  IV U41679 ( .A(n29743), .Z(n29734) );
  IV U41680 ( .A(n28736), .Z(n28739) );
  IV U41681 ( .A(n28737), .Z(n28738) );
  NOR U41682 ( .A(n28739), .B(n28738), .Z(n28740) );
  IV U41683 ( .A(n28740), .Z(n32179) );
  IV U41684 ( .A(n28741), .Z(n28743) );
  XOR U41685 ( .A(n29727), .B(n29731), .Z(n28742) );
  NOR U41686 ( .A(n28743), .B(n28742), .Z(n33115) );
  IV U41687 ( .A(n28744), .Z(n28747) );
  IV U41688 ( .A(n28745), .Z(n28746) );
  NOR U41689 ( .A(n28747), .B(n28746), .Z(n33106) );
  IV U41690 ( .A(n28748), .Z(n28749) );
  NOR U41691 ( .A(n29719), .B(n28749), .Z(n28750) );
  IV U41692 ( .A(n28750), .Z(n32184) );
  IV U41693 ( .A(n32198), .Z(n28751) );
  NOR U41694 ( .A(n32197), .B(n28751), .Z(n28754) );
  NOR U41695 ( .A(n32190), .B(n28752), .Z(n28753) );
  NOR U41696 ( .A(n28754), .B(n28753), .Z(n29716) );
  NOR U41697 ( .A(n35515), .B(n28755), .Z(n32196) );
  IV U41698 ( .A(n28756), .Z(n33099) );
  IV U41699 ( .A(n28757), .Z(n28758) );
  NOR U41700 ( .A(n33099), .B(n28758), .Z(n28759) );
  NOR U41701 ( .A(n28760), .B(n28759), .Z(n29715) );
  IV U41702 ( .A(n28761), .Z(n28763) );
  NOR U41703 ( .A(n28763), .B(n28762), .Z(n29709) );
  IV U41704 ( .A(n28764), .Z(n29700) );
  IV U41705 ( .A(n28765), .Z(n28766) );
  NOR U41706 ( .A(n29700), .B(n28766), .Z(n29706) );
  IV U41707 ( .A(n29706), .Z(n29697) );
  IV U41708 ( .A(n28767), .Z(n28770) );
  IV U41709 ( .A(n28768), .Z(n28775) );
  XOR U41710 ( .A(n28775), .B(n28772), .Z(n28769) );
  NOR U41711 ( .A(n28770), .B(n28769), .Z(n33084) );
  IV U41712 ( .A(n28771), .Z(n28773) );
  IV U41713 ( .A(n28772), .Z(n28774) );
  NOR U41714 ( .A(n28773), .B(n28774), .Z(n35536) );
  NOR U41715 ( .A(n28775), .B(n28774), .Z(n35540) );
  NOR U41716 ( .A(n35536), .B(n35540), .Z(n28776) );
  IV U41717 ( .A(n28776), .Z(n33081) );
  IV U41718 ( .A(n28777), .Z(n28778) );
  NOR U41719 ( .A(n28781), .B(n28778), .Z(n35543) );
  IV U41720 ( .A(n28779), .Z(n28780) );
  NOR U41721 ( .A(n28781), .B(n28780), .Z(n32207) );
  IV U41722 ( .A(n28782), .Z(n28783) );
  NOR U41723 ( .A(n28783), .B(n29682), .Z(n33056) );
  IV U41724 ( .A(n28784), .Z(n35557) );
  NOR U41725 ( .A(n28785), .B(n35557), .Z(n33059) );
  IV U41726 ( .A(n28786), .Z(n28787) );
  NOR U41727 ( .A(n28787), .B(n28791), .Z(n32214) );
  NOR U41728 ( .A(n33059), .B(n32214), .Z(n29680) );
  IV U41729 ( .A(n28788), .Z(n33050) );
  NOR U41730 ( .A(n33050), .B(n28789), .Z(n28793) );
  IV U41731 ( .A(n28790), .Z(n28792) );
  NOR U41732 ( .A(n28792), .B(n28791), .Z(n32217) );
  NOR U41733 ( .A(n28793), .B(n32217), .Z(n29679) );
  IV U41734 ( .A(n28794), .Z(n28796) );
  NOR U41735 ( .A(n28796), .B(n28795), .Z(n33043) );
  IV U41736 ( .A(n28797), .Z(n28798) );
  NOR U41737 ( .A(n28798), .B(n29664), .Z(n28799) );
  IV U41738 ( .A(n28799), .Z(n33042) );
  NOR U41739 ( .A(n28801), .B(n28800), .Z(n28802) );
  IV U41740 ( .A(n28802), .Z(n33004) );
  IV U41741 ( .A(n28803), .Z(n28805) );
  NOR U41742 ( .A(n28805), .B(n28804), .Z(n32981) );
  IV U41743 ( .A(n28806), .Z(n28808) );
  IV U41744 ( .A(n28807), .Z(n28810) );
  NOR U41745 ( .A(n28808), .B(n28810), .Z(n32270) );
  IV U41746 ( .A(n28809), .Z(n28811) );
  NOR U41747 ( .A(n28811), .B(n28810), .Z(n28812) );
  IV U41748 ( .A(n28812), .Z(n32269) );
  IV U41749 ( .A(n28813), .Z(n28814) );
  NOR U41750 ( .A(n29564), .B(n28814), .Z(n29573) );
  IV U41751 ( .A(n28815), .Z(n28817) );
  IV U41752 ( .A(n28816), .Z(n29567) );
  NOR U41753 ( .A(n28817), .B(n29567), .Z(n32956) );
  NOR U41754 ( .A(n28818), .B(n32956), .Z(n29560) );
  IV U41755 ( .A(n28819), .Z(n28821) );
  NOR U41756 ( .A(n28821), .B(n28820), .Z(n32275) );
  IV U41757 ( .A(n28822), .Z(n28823) );
  NOR U41758 ( .A(n28826), .B(n28823), .Z(n32936) );
  IV U41759 ( .A(n28824), .Z(n28825) );
  NOR U41760 ( .A(n28826), .B(n28825), .Z(n32934) );
  IV U41761 ( .A(n28827), .Z(n28830) );
  IV U41762 ( .A(n28828), .Z(n28829) );
  NOR U41763 ( .A(n28830), .B(n28829), .Z(n32929) );
  IV U41764 ( .A(n28831), .Z(n28834) );
  IV U41765 ( .A(n28832), .Z(n28833) );
  NOR U41766 ( .A(n28834), .B(n28833), .Z(n35647) );
  NOR U41767 ( .A(n35653), .B(n35647), .Z(n32928) );
  IV U41768 ( .A(n32928), .Z(n28837) );
  IV U41769 ( .A(n28835), .Z(n28836) );
  NOR U41770 ( .A(n28836), .B(n28841), .Z(n32280) );
  NOR U41771 ( .A(n28837), .B(n32280), .Z(n29546) );
  IV U41772 ( .A(n28838), .Z(n32918) );
  NOR U41773 ( .A(n32918), .B(n28839), .Z(n28843) );
  IV U41774 ( .A(n28840), .Z(n28842) );
  NOR U41775 ( .A(n28842), .B(n28841), .Z(n32925) );
  NOR U41776 ( .A(n28843), .B(n32925), .Z(n29545) );
  IV U41777 ( .A(n28844), .Z(n28846) );
  NOR U41778 ( .A(n28846), .B(n28845), .Z(n32281) );
  IV U41779 ( .A(n28847), .Z(n32286) );
  NOR U41780 ( .A(n32286), .B(n28848), .Z(n29538) );
  IV U41781 ( .A(n28849), .Z(n28851) );
  NOR U41782 ( .A(n28851), .B(n28850), .Z(n29535) );
  IV U41783 ( .A(n29535), .Z(n29522) );
  IV U41784 ( .A(n28852), .Z(n28855) );
  IV U41785 ( .A(n28853), .Z(n28854) );
  NOR U41786 ( .A(n28855), .B(n28854), .Z(n28856) );
  IV U41787 ( .A(n28856), .Z(n32294) );
  IV U41788 ( .A(n28857), .Z(n28859) );
  XOR U41789 ( .A(n29518), .B(n29519), .Z(n28858) );
  NOR U41790 ( .A(n28859), .B(n28858), .Z(n32291) );
  IV U41791 ( .A(n28860), .Z(n28861) );
  NOR U41792 ( .A(n28861), .B(n29519), .Z(n32296) );
  IV U41793 ( .A(n28862), .Z(n28863) );
  NOR U41794 ( .A(n29476), .B(n28863), .Z(n32899) );
  IV U41795 ( .A(n29480), .Z(n28865) );
  IV U41796 ( .A(n28864), .Z(n29479) );
  NOR U41797 ( .A(n28865), .B(n29479), .Z(n32895) );
  IV U41798 ( .A(n28866), .Z(n28867) );
  NOR U41799 ( .A(n28867), .B(n29479), .Z(n32322) );
  NOR U41800 ( .A(n32895), .B(n32322), .Z(n29470) );
  IV U41801 ( .A(n29470), .Z(n29469) );
  IV U41802 ( .A(n28868), .Z(n28869) );
  NOR U41803 ( .A(n29460), .B(n28869), .Z(n32891) );
  IV U41804 ( .A(n28870), .Z(n29434) );
  IV U41805 ( .A(n28871), .Z(n28872) );
  NOR U41806 ( .A(n29434), .B(n28872), .Z(n32861) );
  IV U41807 ( .A(n28873), .Z(n28875) );
  NOR U41808 ( .A(n28875), .B(n28874), .Z(n29429) );
  IV U41809 ( .A(n29429), .Z(n29418) );
  IV U41810 ( .A(n28876), .Z(n28878) );
  NOR U41811 ( .A(n28878), .B(n28877), .Z(n32848) );
  NOR U41812 ( .A(n32377), .B(n28879), .Z(n32368) );
  IV U41813 ( .A(n28880), .Z(n28881) );
  NOR U41814 ( .A(n28881), .B(n29371), .Z(n29390) );
  IV U41815 ( .A(n29390), .Z(n29369) );
  IV U41816 ( .A(n28886), .Z(n28890) );
  IV U41817 ( .A(n28882), .Z(n28883) );
  NOR U41818 ( .A(n28890), .B(n28883), .Z(n32828) );
  IV U41819 ( .A(n28884), .Z(n28888) );
  IV U41820 ( .A(n28885), .Z(n28889) );
  XOR U41821 ( .A(n28889), .B(n28886), .Z(n28887) );
  NOR U41822 ( .A(n28888), .B(n28887), .Z(n32387) );
  NOR U41823 ( .A(n32828), .B(n32387), .Z(n29363) );
  NOR U41824 ( .A(n28890), .B(n28889), .Z(n28891) );
  IV U41825 ( .A(n28891), .Z(n32827) );
  IV U41826 ( .A(n28892), .Z(n28894) );
  NOR U41827 ( .A(n28894), .B(n28893), .Z(n32823) );
  IV U41828 ( .A(n28895), .Z(n28897) );
  NOR U41829 ( .A(n28897), .B(n28896), .Z(n29339) );
  IV U41830 ( .A(n29339), .Z(n29334) );
  IV U41831 ( .A(n28898), .Z(n28899) );
  NOR U41832 ( .A(n28899), .B(n29336), .Z(n32809) );
  IV U41833 ( .A(n28900), .Z(n28901) );
  NOR U41834 ( .A(n28901), .B(n29328), .Z(n28904) );
  IV U41835 ( .A(n28902), .Z(n28909) );
  IV U41836 ( .A(n32808), .Z(n28903) );
  NOR U41837 ( .A(n28909), .B(n28903), .Z(n32799) );
  NOR U41838 ( .A(n28904), .B(n32799), .Z(n32805) );
  IV U41839 ( .A(n28905), .Z(n28906) );
  NOR U41840 ( .A(n28906), .B(n28914), .Z(n36200) );
  IV U41841 ( .A(n28907), .Z(n28908) );
  NOR U41842 ( .A(n28909), .B(n28908), .Z(n35805) );
  NOR U41843 ( .A(n36200), .B(n35805), .Z(n32798) );
  IV U41844 ( .A(n28910), .Z(n28918) );
  IV U41845 ( .A(n28911), .Z(n28912) );
  NOR U41846 ( .A(n28918), .B(n28912), .Z(n32407) );
  IV U41847 ( .A(n28913), .Z(n28915) );
  NOR U41848 ( .A(n28915), .B(n28914), .Z(n32794) );
  NOR U41849 ( .A(n32407), .B(n32794), .Z(n29326) );
  IV U41850 ( .A(n28916), .Z(n28917) );
  NOR U41851 ( .A(n28918), .B(n28917), .Z(n32412) );
  IV U41852 ( .A(n28919), .Z(n29306) );
  NOR U41853 ( .A(n28920), .B(n32421), .Z(n29301) );
  IV U41854 ( .A(n28921), .Z(n28922) );
  NOR U41855 ( .A(n28922), .B(n28924), .Z(n32443) );
  IV U41856 ( .A(n28923), .Z(n28925) );
  NOR U41857 ( .A(n28925), .B(n28924), .Z(n32773) );
  IV U41858 ( .A(n28926), .Z(n29292) );
  IV U41859 ( .A(n28927), .Z(n28928) );
  NOR U41860 ( .A(n29292), .B(n28928), .Z(n29288) );
  IV U41861 ( .A(n29288), .Z(n29274) );
  IV U41862 ( .A(n28929), .Z(n29267) );
  IV U41863 ( .A(n28930), .Z(n32459) );
  NOR U41864 ( .A(n28931), .B(n32459), .Z(n29258) );
  NOR U41865 ( .A(n28932), .B(n32451), .Z(n28933) );
  NOR U41866 ( .A(n29258), .B(n28933), .Z(n29246) );
  IV U41867 ( .A(n28934), .Z(n32735) );
  NOR U41868 ( .A(n32735), .B(n28935), .Z(n28938) );
  NOR U41869 ( .A(n28936), .B(n32465), .Z(n28937) );
  NOR U41870 ( .A(n28938), .B(n28937), .Z(n29244) );
  IV U41871 ( .A(n32727), .Z(n28939) );
  NOR U41872 ( .A(n28939), .B(n28943), .Z(n36113) );
  IV U41873 ( .A(n28940), .Z(n29237) );
  IV U41874 ( .A(n29236), .Z(n29233) );
  NOR U41875 ( .A(n29237), .B(n29233), .Z(n28941) );
  NOR U41876 ( .A(n36113), .B(n28941), .Z(n32724) );
  IV U41877 ( .A(n28942), .Z(n28944) );
  NOR U41878 ( .A(n28944), .B(n28943), .Z(n35868) );
  IV U41879 ( .A(n28945), .Z(n29226) );
  IV U41880 ( .A(n28946), .Z(n28947) );
  NOR U41881 ( .A(n29226), .B(n28947), .Z(n32472) );
  IV U41882 ( .A(n28948), .Z(n28949) );
  NOR U41883 ( .A(n28949), .B(n29228), .Z(n32710) );
  IV U41884 ( .A(n28950), .Z(n35876) );
  NOR U41885 ( .A(n28951), .B(n35876), .Z(n29221) );
  IV U41886 ( .A(n29221), .Z(n29207) );
  NOR U41887 ( .A(n29192), .B(n28952), .Z(n28955) );
  IV U41888 ( .A(n28953), .Z(n28954) );
  NOR U41889 ( .A(n28955), .B(n28954), .Z(n32482) );
  IV U41890 ( .A(n28956), .Z(n28958) );
  NOR U41891 ( .A(n28958), .B(n28957), .Z(n28959) );
  IV U41892 ( .A(n28959), .Z(n32698) );
  NOR U41893 ( .A(n32505), .B(n28960), .Z(n28961) );
  NOR U41894 ( .A(n28961), .B(n32506), .Z(n32496) );
  IV U41895 ( .A(n28962), .Z(n28963) );
  NOR U41896 ( .A(n28963), .B(n29184), .Z(n32501) );
  NOR U41897 ( .A(n28965), .B(n28964), .Z(n28966) );
  IV U41898 ( .A(n28966), .Z(n32688) );
  IV U41899 ( .A(n28967), .Z(n28968) );
  NOR U41900 ( .A(n28968), .B(n29128), .Z(n29148) );
  IV U41901 ( .A(n28969), .Z(n28970) );
  NOR U41902 ( .A(n28971), .B(n28970), .Z(n32663) );
  IV U41903 ( .A(n28972), .Z(n28973) );
  NOR U41904 ( .A(n28973), .B(n28975), .Z(n32539) );
  NOR U41905 ( .A(n32663), .B(n32539), .Z(n29125) );
  IV U41906 ( .A(n28974), .Z(n28976) );
  NOR U41907 ( .A(n28976), .B(n28975), .Z(n32660) );
  IV U41908 ( .A(n28977), .Z(n28982) );
  IV U41909 ( .A(n28978), .Z(n28979) );
  NOR U41910 ( .A(n28982), .B(n28979), .Z(n32657) );
  NOR U41911 ( .A(n32660), .B(n32657), .Z(n29124) );
  IV U41912 ( .A(n28980), .Z(n28981) );
  NOR U41913 ( .A(n28982), .B(n28981), .Z(n32541) );
  IV U41914 ( .A(n28983), .Z(n28985) );
  NOR U41915 ( .A(n28985), .B(n28984), .Z(n32543) );
  NOR U41916 ( .A(n32541), .B(n32543), .Z(n29123) );
  IV U41917 ( .A(n28986), .Z(n28988) );
  IV U41918 ( .A(n28987), .Z(n28989) );
  NOR U41919 ( .A(n28988), .B(n28989), .Z(n32547) );
  NOR U41920 ( .A(n28990), .B(n28989), .Z(n32549) );
  NOR U41921 ( .A(n32553), .B(n28991), .Z(n28992) );
  NOR U41922 ( .A(n32549), .B(n28992), .Z(n28993) );
  IV U41923 ( .A(n28993), .Z(n28994) );
  NOR U41924 ( .A(n32547), .B(n28994), .Z(n29122) );
  IV U41925 ( .A(n29110), .Z(n28995) );
  NOR U41926 ( .A(n28995), .B(n29114), .Z(n32563) );
  IV U41927 ( .A(n28996), .Z(n29001) );
  IV U41928 ( .A(n28997), .Z(n28998) );
  NOR U41929 ( .A(n29001), .B(n28998), .Z(n32560) );
  IV U41930 ( .A(n28999), .Z(n29000) );
  NOR U41931 ( .A(n29001), .B(n29000), .Z(n32569) );
  IV U41932 ( .A(n29002), .Z(n29004) );
  NOR U41933 ( .A(n29004), .B(n29003), .Z(n32566) );
  IV U41934 ( .A(n29005), .Z(n29006) );
  NOR U41935 ( .A(n29006), .B(n29092), .Z(n29007) );
  IV U41936 ( .A(n29007), .Z(n32574) );
  IV U41937 ( .A(n29008), .Z(n29093) );
  IV U41938 ( .A(n29009), .Z(n29088) );
  IV U41939 ( .A(n29010), .Z(n32582) );
  IV U41940 ( .A(n29011), .Z(n29014) );
  IV U41941 ( .A(n29012), .Z(n29013) );
  NOR U41942 ( .A(n29014), .B(n29013), .Z(n32580) );
  IV U41943 ( .A(n32580), .Z(n32638) );
  XOR U41944 ( .A(n32582), .B(n32638), .Z(n29015) );
  NOR U41945 ( .A(n32578), .B(n29015), .Z(n29016) );
  IV U41946 ( .A(n29016), .Z(n29087) );
  IV U41947 ( .A(n29017), .Z(n29019) );
  NOR U41948 ( .A(n29019), .B(n29018), .Z(n32583) );
  IV U41949 ( .A(n29020), .Z(n29021) );
  NOR U41950 ( .A(n29021), .B(n29026), .Z(n32640) );
  IV U41951 ( .A(n29022), .Z(n29024) );
  IV U41952 ( .A(n29023), .Z(n29030) );
  NOR U41953 ( .A(n29024), .B(n29030), .Z(n32628) );
  IV U41954 ( .A(n29025), .Z(n29027) );
  NOR U41955 ( .A(n29027), .B(n29026), .Z(n32634) );
  NOR U41956 ( .A(n32628), .B(n32634), .Z(n29086) );
  NOR U41957 ( .A(n29028), .B(n32622), .Z(n29032) );
  IV U41958 ( .A(n29029), .Z(n29031) );
  NOR U41959 ( .A(n29031), .B(n29030), .Z(n32630) );
  NOR U41960 ( .A(n29032), .B(n32630), .Z(n29085) );
  IV U41961 ( .A(n29033), .Z(n29035) );
  IV U41962 ( .A(n29034), .Z(n29039) );
  NOR U41963 ( .A(n29035), .B(n29039), .Z(n32591) );
  IV U41964 ( .A(n29036), .Z(n29037) );
  NOR U41965 ( .A(n29037), .B(n29045), .Z(n32597) );
  IV U41966 ( .A(n29038), .Z(n29040) );
  NOR U41967 ( .A(n29040), .B(n29039), .Z(n32595) );
  NOR U41968 ( .A(n32597), .B(n32595), .Z(n29084) );
  IV U41969 ( .A(n29041), .Z(n29043) );
  NOR U41970 ( .A(n29043), .B(n29042), .Z(n32603) );
  IV U41971 ( .A(n29044), .Z(n29046) );
  NOR U41972 ( .A(n29046), .B(n29045), .Z(n32616) );
  NOR U41973 ( .A(n32603), .B(n32616), .Z(n29083) );
  IV U41974 ( .A(n29047), .Z(n29048) );
  NOR U41975 ( .A(n29049), .B(n29048), .Z(n32601) );
  IV U41976 ( .A(n32601), .Z(n32600) );
  NOR U41977 ( .A(n29051), .B(n29050), .Z(n29052) );
  NOR U41978 ( .A(n29053), .B(n29052), .Z(n29054) );
  IV U41979 ( .A(n29054), .Z(n32607) );
  IV U41980 ( .A(n29055), .Z(n29056) );
  NOR U41981 ( .A(n29057), .B(n29056), .Z(n32610) );
  NOR U41982 ( .A(n29059), .B(n29058), .Z(n29061) );
  NOR U41983 ( .A(n29061), .B(n29060), .Z(n29062) );
  NOR U41984 ( .A(n32611), .B(n29062), .Z(n29063) );
  NOR U41985 ( .A(n32610), .B(n29063), .Z(n29069) );
  NOR U41986 ( .A(n29065), .B(n29064), .Z(n29066) );
  NOR U41987 ( .A(n32610), .B(n29066), .Z(n29067) );
  NOR U41988 ( .A(n32611), .B(n29067), .Z(n29068) );
  NOR U41989 ( .A(n29069), .B(n29068), .Z(n32612) );
  IV U41990 ( .A(n32612), .Z(n32613) );
  IV U41991 ( .A(n29070), .Z(n29072) );
  NOR U41992 ( .A(n29072), .B(n29071), .Z(n32604) );
  IV U41993 ( .A(n29073), .Z(n29074) );
  NOR U41994 ( .A(n29074), .B(n29077), .Z(n29075) );
  IV U41995 ( .A(n29075), .Z(n32615) );
  IV U41996 ( .A(n29076), .Z(n29078) );
  NOR U41997 ( .A(n29078), .B(n29077), .Z(n29079) );
  NOR U41998 ( .A(n29080), .B(n29079), .Z(n32614) );
  XOR U41999 ( .A(n32615), .B(n32614), .Z(n29081) );
  NOR U42000 ( .A(n32604), .B(n29081), .Z(n29082) );
  XOR U42001 ( .A(n32613), .B(n29082), .Z(n32606) );
  XOR U42002 ( .A(n32607), .B(n32606), .Z(n32602) );
  XOR U42003 ( .A(n32600), .B(n32602), .Z(n32617) );
  XOR U42004 ( .A(n29083), .B(n32617), .Z(n32594) );
  XOR U42005 ( .A(n29084), .B(n32594), .Z(n32592) );
  XOR U42006 ( .A(n32591), .B(n32592), .Z(n32631) );
  XOR U42007 ( .A(n29085), .B(n32631), .Z(n32627) );
  XOR U42008 ( .A(n29086), .B(n32627), .Z(n32642) );
  XOR U42009 ( .A(n32640), .B(n32642), .Z(n32585) );
  XOR U42010 ( .A(n32583), .B(n32585), .Z(n32637) );
  XOR U42011 ( .A(n29087), .B(n32637), .Z(n32576) );
  NOR U42012 ( .A(n29088), .B(n32576), .Z(n29090) );
  IV U42013 ( .A(n29090), .Z(n29094) );
  NOR U42014 ( .A(n29093), .B(n29094), .Z(n35942) );
  IV U42015 ( .A(n29089), .Z(n29091) );
  NOR U42016 ( .A(n29091), .B(n29090), .Z(n29101) );
  NOR U42017 ( .A(n29093), .B(n29092), .Z(n29098) );
  NOR U42018 ( .A(n29095), .B(n29094), .Z(n36004) );
  XOR U42019 ( .A(n32576), .B(n32575), .Z(n29096) );
  NOR U42020 ( .A(n36004), .B(n29096), .Z(n29097) );
  NOR U42021 ( .A(n29098), .B(n29097), .Z(n29099) );
  IV U42022 ( .A(n29099), .Z(n29100) );
  NOR U42023 ( .A(n29101), .B(n29100), .Z(n29102) );
  NOR U42024 ( .A(n35942), .B(n29102), .Z(n32572) );
  XOR U42025 ( .A(n32574), .B(n32572), .Z(n32567) );
  XOR U42026 ( .A(n32566), .B(n32567), .Z(n32571) );
  XOR U42027 ( .A(n32569), .B(n32571), .Z(n32562) );
  XOR U42028 ( .A(n32560), .B(n32562), .Z(n32564) );
  XOR U42029 ( .A(n32563), .B(n32564), .Z(n29108) );
  IV U42030 ( .A(n29103), .Z(n29106) );
  IV U42031 ( .A(n29104), .Z(n29105) );
  NOR U42032 ( .A(n29106), .B(n29105), .Z(n29120) );
  IV U42033 ( .A(n29120), .Z(n29107) );
  NOR U42034 ( .A(n29108), .B(n29107), .Z(n35928) );
  IV U42035 ( .A(n29109), .Z(n29112) );
  XOR U42036 ( .A(n29110), .B(n29114), .Z(n29111) );
  NOR U42037 ( .A(n29112), .B(n29111), .Z(n32556) );
  IV U42038 ( .A(n29113), .Z(n29115) );
  NOR U42039 ( .A(n29115), .B(n29114), .Z(n32558) );
  NOR U42040 ( .A(n32563), .B(n32558), .Z(n29116) );
  IV U42041 ( .A(n29116), .Z(n29117) );
  NOR U42042 ( .A(n32556), .B(n29117), .Z(n29118) );
  XOR U42043 ( .A(n29118), .B(n32564), .Z(n29119) );
  NOR U42044 ( .A(n29120), .B(n29119), .Z(n29121) );
  NOR U42045 ( .A(n35928), .B(n29121), .Z(n32546) );
  XOR U42046 ( .A(n29122), .B(n32546), .Z(n32545) );
  XOR U42047 ( .A(n29123), .B(n32545), .Z(n32658) );
  XOR U42048 ( .A(n29124), .B(n32658), .Z(n32667) );
  XOR U42049 ( .A(n29125), .B(n32667), .Z(n29137) );
  XOR U42050 ( .A(n29126), .B(n29137), .Z(n29139) );
  IV U42051 ( .A(n29127), .Z(n29129) );
  NOR U42052 ( .A(n29129), .B(n29128), .Z(n29145) );
  IV U42053 ( .A(n29145), .Z(n29130) );
  NOR U42054 ( .A(n29139), .B(n29130), .Z(n35917) );
  IV U42055 ( .A(n29131), .Z(n29133) );
  IV U42056 ( .A(n29132), .Z(n29135) );
  NOR U42057 ( .A(n29133), .B(n29135), .Z(n32669) );
  IV U42058 ( .A(n29134), .Z(n29136) );
  NOR U42059 ( .A(n29136), .B(n29135), .Z(n29141) );
  IV U42060 ( .A(n29141), .Z(n29138) );
  IV U42061 ( .A(n29137), .Z(n32674) );
  NOR U42062 ( .A(n29138), .B(n32674), .Z(n32538) );
  IV U42063 ( .A(n29139), .Z(n29140) );
  NOR U42064 ( .A(n29141), .B(n29140), .Z(n29142) );
  NOR U42065 ( .A(n32538), .B(n29142), .Z(n29143) );
  IV U42066 ( .A(n29143), .Z(n32670) );
  XOR U42067 ( .A(n32669), .B(n32670), .Z(n29149) );
  IV U42068 ( .A(n29149), .Z(n29144) );
  NOR U42069 ( .A(n29145), .B(n29144), .Z(n29146) );
  NOR U42070 ( .A(n35917), .B(n29146), .Z(n29147) );
  NOR U42071 ( .A(n29148), .B(n29147), .Z(n29151) );
  IV U42072 ( .A(n29148), .Z(n29150) );
  NOR U42073 ( .A(n29150), .B(n29149), .Z(n36061) );
  NOR U42074 ( .A(n29151), .B(n36061), .Z(n32528) );
  IV U42075 ( .A(n29152), .Z(n32532) );
  NOR U42076 ( .A(n32532), .B(n29153), .Z(n29157) );
  IV U42077 ( .A(n29154), .Z(n29156) );
  NOR U42078 ( .A(n29156), .B(n29155), .Z(n32527) );
  NOR U42079 ( .A(n29157), .B(n32527), .Z(n29158) );
  XOR U42080 ( .A(n32528), .B(n29158), .Z(n32686) );
  XOR U42081 ( .A(n32684), .B(n32686), .Z(n32687) );
  XOR U42082 ( .A(n32688), .B(n32687), .Z(n29168) );
  IV U42083 ( .A(n29168), .Z(n29164) );
  IV U42084 ( .A(n29159), .Z(n29162) );
  IV U42085 ( .A(n29160), .Z(n29166) );
  XOR U42086 ( .A(n29166), .B(n29165), .Z(n29161) );
  NOR U42087 ( .A(n29162), .B(n29161), .Z(n29177) );
  IV U42088 ( .A(n29177), .Z(n29163) );
  NOR U42089 ( .A(n29164), .B(n29163), .Z(n36079) );
  IV U42090 ( .A(n29165), .Z(n29173) );
  NOR U42091 ( .A(n29166), .B(n29173), .Z(n29169) );
  IV U42092 ( .A(n29169), .Z(n29167) );
  NOR U42093 ( .A(n32686), .B(n29167), .Z(n36074) );
  NOR U42094 ( .A(n29169), .B(n29168), .Z(n29170) );
  NOR U42095 ( .A(n36074), .B(n29170), .Z(n29171) );
  IV U42096 ( .A(n29171), .Z(n32692) );
  IV U42097 ( .A(n29172), .Z(n29174) );
  NOR U42098 ( .A(n29174), .B(n29173), .Z(n29175) );
  IV U42099 ( .A(n29175), .Z(n32693) );
  XOR U42100 ( .A(n32692), .B(n32693), .Z(n29176) );
  NOR U42101 ( .A(n29177), .B(n29176), .Z(n29178) );
  NOR U42102 ( .A(n36079), .B(n29178), .Z(n32522) );
  IV U42103 ( .A(n29179), .Z(n29181) );
  NOR U42104 ( .A(n29181), .B(n29180), .Z(n29182) );
  IV U42105 ( .A(n29182), .Z(n32523) );
  XOR U42106 ( .A(n32522), .B(n32523), .Z(n32520) );
  IV U42107 ( .A(n32520), .Z(n29190) );
  IV U42108 ( .A(n29183), .Z(n29185) );
  NOR U42109 ( .A(n29185), .B(n29184), .Z(n32503) );
  IV U42110 ( .A(n29186), .Z(n32518) );
  NOR U42111 ( .A(n32518), .B(n29187), .Z(n29188) );
  NOR U42112 ( .A(n32503), .B(n29188), .Z(n29189) );
  XOR U42113 ( .A(n29190), .B(n29189), .Z(n32510) );
  XOR U42114 ( .A(n32501), .B(n32510), .Z(n32497) );
  XOR U42115 ( .A(n32496), .B(n32497), .Z(n32697) );
  XOR U42116 ( .A(n32698), .B(n32697), .Z(n32489) );
  NOR U42117 ( .A(n32493), .B(n29191), .Z(n29195) );
  IV U42118 ( .A(n29192), .Z(n29194) );
  NOR U42119 ( .A(n29194), .B(n29193), .Z(n32488) );
  NOR U42120 ( .A(n29195), .B(n32488), .Z(n29196) );
  XOR U42121 ( .A(n32489), .B(n29196), .Z(n32484) );
  XOR U42122 ( .A(n32482), .B(n32484), .Z(n32487) );
  IV U42123 ( .A(n29197), .Z(n29199) );
  NOR U42124 ( .A(n29199), .B(n29198), .Z(n32485) );
  XOR U42125 ( .A(n32487), .B(n32485), .Z(n32481) );
  IV U42126 ( .A(n29200), .Z(n29205) );
  IV U42127 ( .A(n29201), .Z(n29202) );
  NOR U42128 ( .A(n29205), .B(n29202), .Z(n32479) );
  IV U42129 ( .A(n29203), .Z(n29204) );
  NOR U42130 ( .A(n29205), .B(n29204), .Z(n32477) );
  NOR U42131 ( .A(n32479), .B(n32477), .Z(n29206) );
  XOR U42132 ( .A(n32481), .B(n29206), .Z(n29216) );
  IV U42133 ( .A(n29216), .Z(n35872) );
  NOR U42134 ( .A(n29207), .B(n35872), .Z(n32714) );
  IV U42135 ( .A(n29208), .Z(n29209) );
  NOR U42136 ( .A(n29209), .B(n29212), .Z(n29210) );
  IV U42137 ( .A(n29210), .Z(n32707) );
  IV U42138 ( .A(n29211), .Z(n29213) );
  NOR U42139 ( .A(n29213), .B(n29212), .Z(n29217) );
  IV U42140 ( .A(n29217), .Z(n29215) );
  XOR U42141 ( .A(n32479), .B(n32481), .Z(n29214) );
  NOR U42142 ( .A(n29215), .B(n29214), .Z(n36101) );
  NOR U42143 ( .A(n29217), .B(n29216), .Z(n29218) );
  NOR U42144 ( .A(n36101), .B(n29218), .Z(n29219) );
  IV U42145 ( .A(n29219), .Z(n32706) );
  XOR U42146 ( .A(n32707), .B(n32706), .Z(n29220) );
  NOR U42147 ( .A(n29221), .B(n29220), .Z(n29222) );
  NOR U42148 ( .A(n32714), .B(n29222), .Z(n29223) );
  IV U42149 ( .A(n29223), .Z(n32711) );
  XOR U42150 ( .A(n32710), .B(n32711), .Z(n32717) );
  IV U42151 ( .A(n32717), .Z(n29231) );
  IV U42152 ( .A(n29224), .Z(n29225) );
  NOR U42153 ( .A(n29226), .B(n29225), .Z(n32475) );
  IV U42154 ( .A(n29227), .Z(n29229) );
  NOR U42155 ( .A(n29229), .B(n29228), .Z(n32715) );
  NOR U42156 ( .A(n32475), .B(n32715), .Z(n29230) );
  XOR U42157 ( .A(n29231), .B(n29230), .Z(n32474) );
  XOR U42158 ( .A(n32472), .B(n32474), .Z(n36110) );
  XOR U42159 ( .A(n35868), .B(n36110), .Z(n32723) );
  XOR U42160 ( .A(n32724), .B(n32723), .Z(n32469) );
  IV U42161 ( .A(n29232), .Z(n29234) );
  NOR U42162 ( .A(n29234), .B(n29233), .Z(n32468) );
  IV U42163 ( .A(n29235), .Z(n29239) );
  XOR U42164 ( .A(n29237), .B(n29236), .Z(n29238) );
  NOR U42165 ( .A(n29239), .B(n29238), .Z(n32728) );
  NOR U42166 ( .A(n32468), .B(n32728), .Z(n29240) );
  XOR U42167 ( .A(n32469), .B(n29240), .Z(n32734) );
  IV U42168 ( .A(n29241), .Z(n29243) );
  NOR U42169 ( .A(n29243), .B(n29242), .Z(n32731) );
  XOR U42170 ( .A(n32734), .B(n32731), .Z(n32464) );
  XOR U42171 ( .A(n29244), .B(n32464), .Z(n29245) );
  IV U42172 ( .A(n29245), .Z(n32460) );
  XOR U42173 ( .A(n29246), .B(n32460), .Z(n29257) );
  IV U42174 ( .A(n29257), .Z(n29250) );
  IV U42175 ( .A(n29247), .Z(n29248) );
  NOR U42176 ( .A(n29248), .B(n29269), .Z(n29262) );
  IV U42177 ( .A(n29262), .Z(n29249) );
  NOR U42178 ( .A(n29250), .B(n29249), .Z(n39119) );
  IV U42179 ( .A(n29251), .Z(n29253) );
  IV U42180 ( .A(n29252), .Z(n29255) );
  NOR U42181 ( .A(n29253), .B(n29255), .Z(n32449) );
  IV U42182 ( .A(n32449), .Z(n39126) );
  IV U42183 ( .A(n29254), .Z(n29256) );
  NOR U42184 ( .A(n29256), .B(n29255), .Z(n32448) );
  NOR U42185 ( .A(n32448), .B(n29257), .Z(n29259) );
  XOR U42186 ( .A(n29258), .B(n32460), .Z(n32756) );
  IV U42187 ( .A(n32448), .Z(n39131) );
  NOR U42188 ( .A(n32756), .B(n39131), .Z(n32760) );
  NOR U42189 ( .A(n29259), .B(n32760), .Z(n29260) );
  IV U42190 ( .A(n29260), .Z(n32759) );
  XOR U42191 ( .A(n39126), .B(n32759), .Z(n29261) );
  NOR U42192 ( .A(n29262), .B(n29261), .Z(n29263) );
  NOR U42193 ( .A(n39119), .B(n29263), .Z(n29264) );
  IV U42194 ( .A(n29264), .Z(n32767) );
  NOR U42195 ( .A(n29267), .B(n32767), .Z(n29265) );
  IV U42196 ( .A(n29265), .Z(n35847) );
  NOR U42197 ( .A(n29266), .B(n35847), .Z(n32769) );
  NOR U42198 ( .A(n29267), .B(n29266), .Z(n29272) );
  IV U42199 ( .A(n29268), .Z(n29270) );
  NOR U42200 ( .A(n29270), .B(n29269), .Z(n32766) );
  XOR U42201 ( .A(n32766), .B(n32767), .Z(n29277) );
  IV U42202 ( .A(n29277), .Z(n29271) );
  NOR U42203 ( .A(n29272), .B(n29271), .Z(n29273) );
  NOR U42204 ( .A(n32769), .B(n29273), .Z(n29279) );
  IV U42205 ( .A(n29279), .Z(n36175) );
  NOR U42206 ( .A(n29274), .B(n36175), .Z(n36169) );
  IV U42207 ( .A(n29275), .Z(n29276) );
  NOR U42208 ( .A(n29276), .B(n29284), .Z(n29280) );
  IV U42209 ( .A(n29280), .Z(n29278) );
  NOR U42210 ( .A(n29278), .B(n29277), .Z(n35845) );
  NOR U42211 ( .A(n29280), .B(n29279), .Z(n29281) );
  NOR U42212 ( .A(n35845), .B(n29281), .Z(n29282) );
  IV U42213 ( .A(n29282), .Z(n32447) );
  IV U42214 ( .A(n29283), .Z(n29285) );
  NOR U42215 ( .A(n29285), .B(n29284), .Z(n29286) );
  IV U42216 ( .A(n29286), .Z(n32446) );
  XOR U42217 ( .A(n32447), .B(n32446), .Z(n29287) );
  NOR U42218 ( .A(n29288), .B(n29287), .Z(n29289) );
  NOR U42219 ( .A(n36169), .B(n29289), .Z(n32771) );
  IV U42220 ( .A(n29290), .Z(n29291) );
  NOR U42221 ( .A(n29292), .B(n29291), .Z(n29293) );
  IV U42222 ( .A(n29293), .Z(n36172) );
  XOR U42223 ( .A(n32771), .B(n36172), .Z(n32774) );
  XOR U42224 ( .A(n32773), .B(n32774), .Z(n32444) );
  XOR U42225 ( .A(n32443), .B(n32444), .Z(n32429) );
  IV U42226 ( .A(n32429), .Z(n29300) );
  NOR U42227 ( .A(n32437), .B(n29294), .Z(n29298) );
  IV U42228 ( .A(n29295), .Z(n32430) );
  NOR U42229 ( .A(n29296), .B(n32430), .Z(n29297) );
  NOR U42230 ( .A(n29298), .B(n29297), .Z(n29299) );
  XOR U42231 ( .A(n29300), .B(n29299), .Z(n32422) );
  XOR U42232 ( .A(n29301), .B(n32422), .Z(n29310) );
  IV U42233 ( .A(n29302), .Z(n29308) );
  XOR U42234 ( .A(n29308), .B(n29305), .Z(n29303) );
  NOR U42235 ( .A(n29310), .B(n29303), .Z(n29304) );
  IV U42236 ( .A(n29304), .Z(n32790) );
  NOR U42237 ( .A(n29306), .B(n32790), .Z(n32419) );
  IV U42238 ( .A(n29305), .Z(n29307) );
  NOR U42239 ( .A(n29306), .B(n29307), .Z(n29314) );
  NOR U42240 ( .A(n29308), .B(n29307), .Z(n29312) );
  IV U42241 ( .A(n29312), .Z(n29309) );
  NOR U42242 ( .A(n32422), .B(n29309), .Z(n32783) );
  IV U42243 ( .A(n29310), .Z(n29311) );
  NOR U42244 ( .A(n29312), .B(n29311), .Z(n29313) );
  NOR U42245 ( .A(n32783), .B(n29313), .Z(n32415) );
  NOR U42246 ( .A(n29314), .B(n32415), .Z(n29315) );
  NOR U42247 ( .A(n32419), .B(n29315), .Z(n29322) );
  IV U42248 ( .A(n29316), .Z(n32791) );
  NOR U42249 ( .A(n32791), .B(n29318), .Z(n29320) );
  IV U42250 ( .A(n29317), .Z(n29319) );
  NOR U42251 ( .A(n29319), .B(n29318), .Z(n32416) );
  NOR U42252 ( .A(n29320), .B(n32416), .Z(n29321) );
  XOR U42253 ( .A(n29322), .B(n29321), .Z(n32411) );
  IV U42254 ( .A(n29323), .Z(n29325) );
  NOR U42255 ( .A(n29325), .B(n29324), .Z(n32409) );
  XOR U42256 ( .A(n32411), .B(n32409), .Z(n32413) );
  XOR U42257 ( .A(n32412), .B(n32413), .Z(n32796) );
  XOR U42258 ( .A(n29326), .B(n32796), .Z(n32797) );
  XOR U42259 ( .A(n32798), .B(n32797), .Z(n32804) );
  XOR U42260 ( .A(n32805), .B(n32804), .Z(n32396) );
  IV U42261 ( .A(n29327), .Z(n29329) );
  NOR U42262 ( .A(n29329), .B(n29328), .Z(n32404) );
  IV U42263 ( .A(n29330), .Z(n32397) );
  NOR U42264 ( .A(n29331), .B(n32397), .Z(n29332) );
  NOR U42265 ( .A(n32404), .B(n29332), .Z(n29333) );
  XOR U42266 ( .A(n32396), .B(n29333), .Z(n32811) );
  XOR U42267 ( .A(n32809), .B(n32811), .Z(n32813) );
  NOR U42268 ( .A(n29334), .B(n32813), .Z(n35788) );
  IV U42269 ( .A(n29335), .Z(n29337) );
  NOR U42270 ( .A(n29337), .B(n29336), .Z(n32812) );
  XOR U42271 ( .A(n32812), .B(n32813), .Z(n32393) );
  IV U42272 ( .A(n32393), .Z(n29338) );
  NOR U42273 ( .A(n29339), .B(n29338), .Z(n29340) );
  NOR U42274 ( .A(n35788), .B(n29340), .Z(n29347) );
  IV U42275 ( .A(n29341), .Z(n29342) );
  NOR U42276 ( .A(n29342), .B(n29344), .Z(n32392) );
  IV U42277 ( .A(n29343), .Z(n29345) );
  NOR U42278 ( .A(n29345), .B(n29344), .Z(n32390) );
  NOR U42279 ( .A(n32392), .B(n32390), .Z(n29346) );
  XOR U42280 ( .A(n29347), .B(n29346), .Z(n32819) );
  IV U42281 ( .A(n29348), .Z(n29349) );
  NOR U42282 ( .A(n29353), .B(n29349), .Z(n29359) );
  IV U42283 ( .A(n29359), .Z(n29350) );
  NOR U42284 ( .A(n32819), .B(n29350), .Z(n36212) );
  IV U42285 ( .A(n29351), .Z(n29352) );
  NOR U42286 ( .A(n29353), .B(n29352), .Z(n29354) );
  IV U42287 ( .A(n29354), .Z(n32821) );
  IV U42288 ( .A(n29355), .Z(n29357) );
  NOR U42289 ( .A(n29357), .B(n29356), .Z(n32817) );
  XOR U42290 ( .A(n32817), .B(n32819), .Z(n32820) );
  XOR U42291 ( .A(n32821), .B(n32820), .Z(n29358) );
  NOR U42292 ( .A(n29359), .B(n29358), .Z(n29360) );
  NOR U42293 ( .A(n36212), .B(n29360), .Z(n29361) );
  IV U42294 ( .A(n29361), .Z(n32824) );
  XOR U42295 ( .A(n32823), .B(n32824), .Z(n32829) );
  XOR U42296 ( .A(n32827), .B(n32829), .Z(n29362) );
  XOR U42297 ( .A(n29363), .B(n29362), .Z(n32385) );
  IV U42298 ( .A(n29364), .Z(n29366) );
  NOR U42299 ( .A(n29366), .B(n29365), .Z(n29367) );
  IV U42300 ( .A(n29367), .Z(n32384) );
  XOR U42301 ( .A(n32385), .B(n32384), .Z(n29376) );
  IV U42302 ( .A(n29376), .Z(n29368) );
  NOR U42303 ( .A(n29369), .B(n29368), .Z(n32381) );
  IV U42304 ( .A(n29370), .Z(n29372) );
  NOR U42305 ( .A(n29372), .B(n29371), .Z(n29373) );
  IV U42306 ( .A(n29373), .Z(n32383) );
  IV U42307 ( .A(n29374), .Z(n29379) );
  NOR U42308 ( .A(n29379), .B(n29375), .Z(n29377) );
  NOR U42309 ( .A(n29377), .B(n29376), .Z(n29387) );
  IV U42310 ( .A(n29378), .Z(n29381) );
  NOR U42311 ( .A(n29379), .B(n32385), .Z(n29380) );
  IV U42312 ( .A(n29380), .Z(n29383) );
  NOR U42313 ( .A(n29381), .B(n29383), .Z(n32836) );
  IV U42314 ( .A(n29382), .Z(n29384) );
  NOR U42315 ( .A(n29384), .B(n29383), .Z(n32833) );
  NOR U42316 ( .A(n32836), .B(n32833), .Z(n29385) );
  IV U42317 ( .A(n29385), .Z(n29386) );
  NOR U42318 ( .A(n29387), .B(n29386), .Z(n29388) );
  IV U42319 ( .A(n29388), .Z(n32382) );
  XOR U42320 ( .A(n32383), .B(n32382), .Z(n29389) );
  NOR U42321 ( .A(n29390), .B(n29389), .Z(n29391) );
  NOR U42322 ( .A(n32381), .B(n29391), .Z(n32372) );
  IV U42323 ( .A(n29392), .Z(n29394) );
  NOR U42324 ( .A(n29394), .B(n29393), .Z(n29395) );
  IV U42325 ( .A(n29395), .Z(n32373) );
  XOR U42326 ( .A(n32372), .B(n32373), .Z(n32376) );
  XOR U42327 ( .A(n32368), .B(n32376), .Z(n32357) );
  IV U42328 ( .A(n29399), .Z(n32362) );
  NOR U42329 ( .A(n29397), .B(n32362), .Z(n29402) );
  IV U42330 ( .A(n29396), .Z(n32360) );
  IV U42331 ( .A(n29397), .Z(n29398) );
  NOR U42332 ( .A(n29399), .B(n29398), .Z(n29400) );
  NOR U42333 ( .A(n32360), .B(n29400), .Z(n29401) );
  NOR U42334 ( .A(n29402), .B(n29401), .Z(n29403) );
  XOR U42335 ( .A(n32357), .B(n29403), .Z(n32355) );
  IV U42336 ( .A(n29404), .Z(n29405) );
  NOR U42337 ( .A(n29408), .B(n29405), .Z(n32846) );
  IV U42338 ( .A(n29406), .Z(n29407) );
  NOR U42339 ( .A(n29408), .B(n29407), .Z(n35751) );
  IV U42340 ( .A(n29409), .Z(n35763) );
  NOR U42341 ( .A(n32358), .B(n35763), .Z(n29410) );
  NOR U42342 ( .A(n35751), .B(n29410), .Z(n32356) );
  IV U42343 ( .A(n32356), .Z(n29411) );
  NOR U42344 ( .A(n32846), .B(n29411), .Z(n29412) );
  XOR U42345 ( .A(n32355), .B(n29412), .Z(n32849) );
  XOR U42346 ( .A(n32848), .B(n32849), .Z(n32854) );
  IV U42347 ( .A(n29413), .Z(n32351) );
  NOR U42348 ( .A(n32351), .B(n29414), .Z(n32346) );
  NOR U42349 ( .A(n29415), .B(n32342), .Z(n32853) );
  NOR U42350 ( .A(n32346), .B(n32853), .Z(n29416) );
  XOR U42351 ( .A(n32854), .B(n29416), .Z(n29426) );
  IV U42352 ( .A(n29426), .Z(n29417) );
  NOR U42353 ( .A(n29418), .B(n29417), .Z(n35727) );
  IV U42354 ( .A(n29419), .Z(n29420) );
  NOR U42355 ( .A(n29420), .B(n29422), .Z(n36246) );
  IV U42356 ( .A(n29421), .Z(n29423) );
  NOR U42357 ( .A(n29423), .B(n29422), .Z(n35732) );
  NOR U42358 ( .A(n36246), .B(n35732), .Z(n29424) );
  XOR U42359 ( .A(n32346), .B(n32854), .Z(n35734) );
  NOR U42360 ( .A(n29424), .B(n35734), .Z(n32860) );
  IV U42361 ( .A(n29424), .Z(n29425) );
  NOR U42362 ( .A(n29426), .B(n29425), .Z(n29427) );
  NOR U42363 ( .A(n32860), .B(n29427), .Z(n29428) );
  NOR U42364 ( .A(n29429), .B(n29428), .Z(n29430) );
  NOR U42365 ( .A(n35727), .B(n29430), .Z(n29431) );
  IV U42366 ( .A(n29431), .Z(n32862) );
  XOR U42367 ( .A(n32861), .B(n32862), .Z(n32866) );
  IV U42368 ( .A(n29432), .Z(n29433) );
  NOR U42369 ( .A(n29434), .B(n29433), .Z(n32864) );
  XOR U42370 ( .A(n32866), .B(n32864), .Z(n32870) );
  IV U42371 ( .A(n29435), .Z(n29436) );
  NOR U42372 ( .A(n29436), .B(n29438), .Z(n32869) );
  IV U42373 ( .A(n29437), .Z(n29439) );
  NOR U42374 ( .A(n29439), .B(n29438), .Z(n32340) );
  NOR U42375 ( .A(n32869), .B(n32340), .Z(n29440) );
  XOR U42376 ( .A(n32870), .B(n29440), .Z(n32334) );
  IV U42377 ( .A(n29441), .Z(n29450) );
  IV U42378 ( .A(n29442), .Z(n29443) );
  NOR U42379 ( .A(n29450), .B(n29443), .Z(n32335) );
  IV U42380 ( .A(n29444), .Z(n29446) );
  NOR U42381 ( .A(n29446), .B(n29445), .Z(n32337) );
  NOR U42382 ( .A(n32335), .B(n32337), .Z(n29447) );
  XOR U42383 ( .A(n32334), .B(n29447), .Z(n32328) );
  IV U42384 ( .A(n29448), .Z(n29449) );
  NOR U42385 ( .A(n29450), .B(n29449), .Z(n29451) );
  IV U42386 ( .A(n29451), .Z(n32327) );
  XOR U42387 ( .A(n32328), .B(n32327), .Z(n32332) );
  IV U42388 ( .A(n29452), .Z(n29454) );
  IV U42389 ( .A(n29453), .Z(n29463) );
  NOR U42390 ( .A(n29454), .B(n29463), .Z(n32874) );
  NOR U42391 ( .A(n29455), .B(n32878), .Z(n29456) );
  NOR U42392 ( .A(n32874), .B(n29456), .Z(n29457) );
  XOR U42393 ( .A(n32332), .B(n29457), .Z(n32326) );
  IV U42394 ( .A(n29458), .Z(n29459) );
  NOR U42395 ( .A(n29460), .B(n29459), .Z(n29465) );
  IV U42396 ( .A(n29465), .Z(n29461) );
  NOR U42397 ( .A(n32326), .B(n29461), .Z(n35718) );
  IV U42398 ( .A(n29462), .Z(n29464) );
  NOR U42399 ( .A(n29464), .B(n29463), .Z(n32324) );
  XOR U42400 ( .A(n32324), .B(n32326), .Z(n32896) );
  IV U42401 ( .A(n32896), .Z(n29471) );
  NOR U42402 ( .A(n29471), .B(n29465), .Z(n29466) );
  NOR U42403 ( .A(n35718), .B(n29466), .Z(n29467) );
  IV U42404 ( .A(n29467), .Z(n32892) );
  XOR U42405 ( .A(n32891), .B(n32892), .Z(n29468) );
  NOR U42406 ( .A(n29469), .B(n29468), .Z(n29473) );
  NOR U42407 ( .A(n29471), .B(n29470), .Z(n29472) );
  NOR U42408 ( .A(n29473), .B(n29472), .Z(n32319) );
  IV U42409 ( .A(n29474), .Z(n29475) );
  NOR U42410 ( .A(n29476), .B(n29475), .Z(n29488) );
  IV U42411 ( .A(n29488), .Z(n29477) );
  NOR U42412 ( .A(n32319), .B(n29477), .Z(n35699) );
  IV U42413 ( .A(n29478), .Z(n29482) );
  XOR U42414 ( .A(n29480), .B(n29479), .Z(n29481) );
  NOR U42415 ( .A(n29482), .B(n29481), .Z(n32317) );
  XOR U42416 ( .A(n32317), .B(n32319), .Z(n32321) );
  IV U42417 ( .A(n29483), .Z(n29485) );
  NOR U42418 ( .A(n29485), .B(n29484), .Z(n29486) );
  IV U42419 ( .A(n29486), .Z(n32320) );
  XOR U42420 ( .A(n32321), .B(n32320), .Z(n29487) );
  NOR U42421 ( .A(n29488), .B(n29487), .Z(n29489) );
  NOR U42422 ( .A(n35699), .B(n29489), .Z(n29490) );
  IV U42423 ( .A(n29490), .Z(n32900) );
  XOR U42424 ( .A(n32899), .B(n32900), .Z(n32306) );
  IV U42425 ( .A(n29491), .Z(n29493) );
  NOR U42426 ( .A(n29493), .B(n29492), .Z(n32302) );
  NOR U42427 ( .A(n29495), .B(n29494), .Z(n29499) );
  NOR U42428 ( .A(n29496), .B(n32311), .Z(n32309) );
  NOR U42429 ( .A(n29497), .B(n32309), .Z(n29498) );
  NOR U42430 ( .A(n29499), .B(n29498), .Z(n32304) );
  NOR U42431 ( .A(n32302), .B(n32304), .Z(n29500) );
  XOR U42432 ( .A(n32306), .B(n29500), .Z(n29512) );
  IV U42433 ( .A(n29512), .Z(n29505) );
  IV U42434 ( .A(n29501), .Z(n29508) );
  IV U42435 ( .A(n29502), .Z(n29503) );
  NOR U42436 ( .A(n29508), .B(n29503), .Z(n29515) );
  IV U42437 ( .A(n29515), .Z(n29504) );
  NOR U42438 ( .A(n29505), .B(n29504), .Z(n35686) );
  XOR U42439 ( .A(n32304), .B(n32306), .Z(n29510) );
  IV U42440 ( .A(n29506), .Z(n29507) );
  NOR U42441 ( .A(n29508), .B(n29507), .Z(n29511) );
  IV U42442 ( .A(n29511), .Z(n29509) );
  NOR U42443 ( .A(n29510), .B(n29509), .Z(n35688) );
  NOR U42444 ( .A(n29512), .B(n29511), .Z(n29513) );
  NOR U42445 ( .A(n35688), .B(n29513), .Z(n29514) );
  NOR U42446 ( .A(n29515), .B(n29514), .Z(n29516) );
  NOR U42447 ( .A(n35686), .B(n29516), .Z(n29517) );
  IV U42448 ( .A(n29517), .Z(n32300) );
  IV U42449 ( .A(n29518), .Z(n29520) );
  NOR U42450 ( .A(n29520), .B(n29519), .Z(n32299) );
  XOR U42451 ( .A(n32300), .B(n32299), .Z(n32297) );
  XOR U42452 ( .A(n32296), .B(n32297), .Z(n32292) );
  XOR U42453 ( .A(n32291), .B(n32292), .Z(n32295) );
  XOR U42454 ( .A(n32294), .B(n32295), .Z(n29526) );
  IV U42455 ( .A(n29526), .Z(n29521) );
  NOR U42456 ( .A(n29522), .B(n29521), .Z(n42457) );
  IV U42457 ( .A(n29523), .Z(n29524) );
  NOR U42458 ( .A(n29532), .B(n29524), .Z(n29527) );
  IV U42459 ( .A(n29527), .Z(n29525) );
  NOR U42460 ( .A(n29525), .B(n32295), .Z(n35677) );
  NOR U42461 ( .A(n29527), .B(n29526), .Z(n29528) );
  NOR U42462 ( .A(n35677), .B(n29528), .Z(n29529) );
  IV U42463 ( .A(n29529), .Z(n32290) );
  IV U42464 ( .A(n29530), .Z(n29531) );
  NOR U42465 ( .A(n29532), .B(n29531), .Z(n29533) );
  IV U42466 ( .A(n29533), .Z(n32289) );
  XOR U42467 ( .A(n32290), .B(n32289), .Z(n29534) );
  NOR U42468 ( .A(n29535), .B(n29534), .Z(n29536) );
  NOR U42469 ( .A(n42457), .B(n29536), .Z(n29537) );
  IV U42470 ( .A(n29537), .Z(n36329) );
  XOR U42471 ( .A(n29538), .B(n36329), .Z(n32283) );
  IV U42472 ( .A(n32283), .Z(n29544) );
  IV U42473 ( .A(n29539), .Z(n29540) );
  NOR U42474 ( .A(n29540), .B(n29542), .Z(n36313) );
  IV U42475 ( .A(n29541), .Z(n29543) );
  NOR U42476 ( .A(n29543), .B(n29542), .Z(n36324) );
  NOR U42477 ( .A(n36313), .B(n36324), .Z(n32284) );
  XOR U42478 ( .A(n29544), .B(n32284), .Z(n32917) );
  XOR U42479 ( .A(n32281), .B(n32917), .Z(n32926) );
  XOR U42480 ( .A(n29545), .B(n32926), .Z(n35654) );
  XOR U42481 ( .A(n29546), .B(n35654), .Z(n32930) );
  XOR U42482 ( .A(n32929), .B(n32930), .Z(n36337) );
  XOR U42483 ( .A(n32934), .B(n36337), .Z(n32937) );
  XOR U42484 ( .A(n32936), .B(n32937), .Z(n32941) );
  IV U42485 ( .A(n32941), .Z(n29553) );
  NOR U42486 ( .A(n29547), .B(n32942), .Z(n29557) );
  IV U42487 ( .A(n29557), .Z(n29548) );
  NOR U42488 ( .A(n29553), .B(n29548), .Z(n29559) );
  IV U42489 ( .A(n29549), .Z(n36340) );
  NOR U42490 ( .A(n29550), .B(n36340), .Z(n29552) );
  IV U42491 ( .A(n29552), .Z(n29551) );
  NOR U42492 ( .A(n29551), .B(n36337), .Z(n32945) );
  NOR U42493 ( .A(n29553), .B(n29552), .Z(n29554) );
  NOR U42494 ( .A(n32945), .B(n29554), .Z(n29555) );
  IV U42495 ( .A(n29555), .Z(n29556) );
  NOR U42496 ( .A(n29557), .B(n29556), .Z(n29558) );
  NOR U42497 ( .A(n29559), .B(n29558), .Z(n32276) );
  XOR U42498 ( .A(n32275), .B(n32276), .Z(n32958) );
  XOR U42499 ( .A(n29560), .B(n32958), .Z(n29561) );
  IV U42500 ( .A(n29561), .Z(n32955) );
  IV U42501 ( .A(n29562), .Z(n29563) );
  NOR U42502 ( .A(n29564), .B(n29563), .Z(n29570) );
  IV U42503 ( .A(n29570), .Z(n29565) );
  NOR U42504 ( .A(n32955), .B(n29565), .Z(n35633) );
  IV U42505 ( .A(n29566), .Z(n29568) );
  NOR U42506 ( .A(n29568), .B(n29567), .Z(n32953) );
  XOR U42507 ( .A(n32953), .B(n32955), .Z(n29574) );
  IV U42508 ( .A(n29574), .Z(n29569) );
  NOR U42509 ( .A(n29570), .B(n29569), .Z(n29571) );
  NOR U42510 ( .A(n35633), .B(n29571), .Z(n29572) );
  NOR U42511 ( .A(n29573), .B(n29572), .Z(n29576) );
  IV U42512 ( .A(n29573), .Z(n29575) );
  NOR U42513 ( .A(n29575), .B(n29574), .Z(n35630) );
  NOR U42514 ( .A(n29576), .B(n35630), .Z(n29586) );
  XOR U42515 ( .A(n32269), .B(n29586), .Z(n32272) );
  XOR U42516 ( .A(n32270), .B(n32272), .Z(n32268) );
  IV U42517 ( .A(n29577), .Z(n29579) );
  IV U42518 ( .A(n29578), .Z(n29588) );
  NOR U42519 ( .A(n29579), .B(n29588), .Z(n29580) );
  IV U42520 ( .A(n29580), .Z(n29595) );
  NOR U42521 ( .A(n32268), .B(n29595), .Z(n36374) );
  IV U42522 ( .A(n29581), .Z(n29582) );
  NOR U42523 ( .A(n29602), .B(n29582), .Z(n29583) );
  IV U42524 ( .A(n29583), .Z(n32965) );
  NOR U42525 ( .A(n35618), .B(n29584), .Z(n29585) );
  IV U42526 ( .A(n29585), .Z(n29590) );
  IV U42527 ( .A(n29586), .Z(n35614) );
  NOR U42528 ( .A(n29590), .B(n35614), .Z(n32963) );
  IV U42529 ( .A(n29587), .Z(n29589) );
  NOR U42530 ( .A(n29589), .B(n29588), .Z(n29591) );
  IV U42531 ( .A(n29591), .Z(n32267) );
  XOR U42532 ( .A(n32268), .B(n32267), .Z(n29593) );
  NOR U42533 ( .A(n29591), .B(n29590), .Z(n29592) );
  NOR U42534 ( .A(n29593), .B(n29592), .Z(n29594) );
  NOR U42535 ( .A(n32963), .B(n29594), .Z(n29596) );
  IV U42536 ( .A(n29596), .Z(n32964) );
  XOR U42537 ( .A(n32965), .B(n32964), .Z(n29598) );
  NOR U42538 ( .A(n29596), .B(n29595), .Z(n29597) );
  NOR U42539 ( .A(n29598), .B(n29597), .Z(n29599) );
  NOR U42540 ( .A(n36374), .B(n29599), .Z(n32966) );
  IV U42541 ( .A(n29600), .Z(n29601) );
  NOR U42542 ( .A(n29602), .B(n29601), .Z(n29603) );
  IV U42543 ( .A(n29603), .Z(n32967) );
  XOR U42544 ( .A(n32966), .B(n32967), .Z(n32266) );
  IV U42545 ( .A(n29604), .Z(n29606) );
  NOR U42546 ( .A(n29606), .B(n29605), .Z(n32264) );
  XOR U42547 ( .A(n32266), .B(n32264), .Z(n32255) );
  IV U42548 ( .A(n29607), .Z(n32258) );
  NOR U42549 ( .A(n32258), .B(n29608), .Z(n29610) );
  IV U42550 ( .A(n29616), .Z(n29609) );
  NOR U42551 ( .A(n29609), .B(n29615), .Z(n32254) );
  NOR U42552 ( .A(n29610), .B(n32254), .Z(n29611) );
  XOR U42553 ( .A(n32255), .B(n29611), .Z(n32248) );
  IV U42554 ( .A(n29612), .Z(n29613) );
  NOR U42555 ( .A(n29613), .B(n29615), .Z(n32251) );
  IV U42556 ( .A(n29614), .Z(n29618) );
  XOR U42557 ( .A(n29616), .B(n29615), .Z(n29617) );
  NOR U42558 ( .A(n29618), .B(n29617), .Z(n32249) );
  NOR U42559 ( .A(n32251), .B(n32249), .Z(n29619) );
  XOR U42560 ( .A(n32248), .B(n29619), .Z(n32244) );
  IV U42561 ( .A(n29620), .Z(n29622) );
  NOR U42562 ( .A(n29622), .B(n29621), .Z(n32241) );
  XOR U42563 ( .A(n32244), .B(n32241), .Z(n32977) );
  NOR U42564 ( .A(n29624), .B(n29623), .Z(n29630) );
  NOR U42565 ( .A(n32245), .B(n29625), .Z(n29628) );
  NOR U42566 ( .A(n32976), .B(n32983), .Z(n29626) );
  IV U42567 ( .A(n29626), .Z(n29627) );
  NOR U42568 ( .A(n29628), .B(n29627), .Z(n29629) );
  NOR U42569 ( .A(n29630), .B(n29629), .Z(n29631) );
  XOR U42570 ( .A(n32977), .B(n29631), .Z(n32986) );
  XOR U42571 ( .A(n32981), .B(n32986), .Z(n32994) );
  IV U42572 ( .A(n29632), .Z(n32990) );
  NOR U42573 ( .A(n32990), .B(n32992), .Z(n32993) );
  IV U42574 ( .A(n29633), .Z(n29634) );
  NOR U42575 ( .A(n29634), .B(n29637), .Z(n32238) );
  NOR U42576 ( .A(n32993), .B(n32238), .Z(n29635) );
  XOR U42577 ( .A(n32994), .B(n29635), .Z(n32230) );
  IV U42578 ( .A(n29636), .Z(n29638) );
  NOR U42579 ( .A(n29638), .B(n29637), .Z(n32236) );
  IV U42580 ( .A(n29639), .Z(n29643) );
  NOR U42581 ( .A(n29643), .B(n29640), .Z(n32233) );
  IV U42582 ( .A(n29641), .Z(n29642) );
  NOR U42583 ( .A(n29643), .B(n29642), .Z(n32231) );
  NOR U42584 ( .A(n32233), .B(n32231), .Z(n29644) );
  IV U42585 ( .A(n29644), .Z(n29645) );
  NOR U42586 ( .A(n32236), .B(n29645), .Z(n29646) );
  XOR U42587 ( .A(n32230), .B(n29646), .Z(n32228) );
  IV U42588 ( .A(n29647), .Z(n32224) );
  NOR U42589 ( .A(n32224), .B(n29648), .Z(n29652) );
  IV U42590 ( .A(n29649), .Z(n29651) );
  NOR U42591 ( .A(n29651), .B(n29650), .Z(n32227) );
  NOR U42592 ( .A(n29652), .B(n32227), .Z(n29653) );
  XOR U42593 ( .A(n32228), .B(n29653), .Z(n33003) );
  XOR U42594 ( .A(n33004), .B(n33003), .Z(n33019) );
  IV U42595 ( .A(n29654), .Z(n33014) );
  NOR U42596 ( .A(n29655), .B(n33014), .Z(n29656) );
  NOR U42597 ( .A(n29656), .B(n33020), .Z(n29657) );
  XOR U42598 ( .A(n33019), .B(n29657), .Z(n29674) );
  NOR U42599 ( .A(n29658), .B(n33021), .Z(n29671) );
  IV U42600 ( .A(n29659), .Z(n29661) );
  IV U42601 ( .A(n29660), .Z(n29669) );
  NOR U42602 ( .A(n29661), .B(n29669), .Z(n35577) );
  NOR U42603 ( .A(n29671), .B(n35577), .Z(n29662) );
  XOR U42604 ( .A(n29674), .B(n29662), .Z(n29667) );
  IV U42605 ( .A(n29663), .Z(n29665) );
  NOR U42606 ( .A(n29665), .B(n29664), .Z(n29677) );
  IV U42607 ( .A(n29677), .Z(n29666) );
  NOR U42608 ( .A(n29667), .B(n29666), .Z(n35564) );
  IV U42609 ( .A(n29668), .Z(n29670) );
  NOR U42610 ( .A(n29670), .B(n29669), .Z(n35569) );
  NOR U42611 ( .A(n35569), .B(n29671), .Z(n29672) );
  IV U42612 ( .A(n29672), .Z(n29673) );
  NOR U42613 ( .A(n35577), .B(n29673), .Z(n29675) );
  IV U42614 ( .A(n29674), .Z(n35571) );
  XOR U42615 ( .A(n29675), .B(n35571), .Z(n29676) );
  NOR U42616 ( .A(n29677), .B(n29676), .Z(n29678) );
  NOR U42617 ( .A(n35564), .B(n29678), .Z(n33040) );
  XOR U42618 ( .A(n33042), .B(n33040), .Z(n33044) );
  XOR U42619 ( .A(n33043), .B(n33044), .Z(n33052) );
  XOR U42620 ( .A(n29679), .B(n33052), .Z(n32213) );
  XOR U42621 ( .A(n29680), .B(n32213), .Z(n33057) );
  XOR U42622 ( .A(n33056), .B(n33057), .Z(n33066) );
  IV U42623 ( .A(n33066), .Z(n33071) );
  IV U42624 ( .A(n29681), .Z(n29683) );
  NOR U42625 ( .A(n29683), .B(n29682), .Z(n32211) );
  IV U42626 ( .A(n29684), .Z(n29687) );
  IV U42627 ( .A(n29685), .Z(n29686) );
  NOR U42628 ( .A(n29687), .B(n29686), .Z(n33065) );
  NOR U42629 ( .A(n33070), .B(n33065), .Z(n32210) );
  IV U42630 ( .A(n32210), .Z(n29688) );
  NOR U42631 ( .A(n32211), .B(n29688), .Z(n29689) );
  XOR U42632 ( .A(n33071), .B(n29689), .Z(n32206) );
  IV U42633 ( .A(n29690), .Z(n29693) );
  IV U42634 ( .A(n29691), .Z(n29692) );
  NOR U42635 ( .A(n29693), .B(n29692), .Z(n32204) );
  XOR U42636 ( .A(n32206), .B(n32204), .Z(n32208) );
  XOR U42637 ( .A(n32207), .B(n32208), .Z(n35544) );
  XOR U42638 ( .A(n35543), .B(n35544), .Z(n35537) );
  XOR U42639 ( .A(n33081), .B(n35537), .Z(n33086) );
  XOR U42640 ( .A(n33084), .B(n33086), .Z(n33089) );
  IV U42641 ( .A(n29694), .Z(n29696) );
  NOR U42642 ( .A(n29696), .B(n29695), .Z(n33087) );
  XOR U42643 ( .A(n33089), .B(n33087), .Z(n29702) );
  NOR U42644 ( .A(n29697), .B(n29702), .Z(n35528) );
  IV U42645 ( .A(n29698), .Z(n29699) );
  NOR U42646 ( .A(n29700), .B(n29699), .Z(n29704) );
  IV U42647 ( .A(n29704), .Z(n29701) );
  NOR U42648 ( .A(n29701), .B(n33089), .Z(n32203) );
  IV U42649 ( .A(n29702), .Z(n29703) );
  NOR U42650 ( .A(n29704), .B(n29703), .Z(n29705) );
  NOR U42651 ( .A(n32203), .B(n29705), .Z(n29710) );
  NOR U42652 ( .A(n29706), .B(n29710), .Z(n29707) );
  NOR U42653 ( .A(n35528), .B(n29707), .Z(n29708) );
  NOR U42654 ( .A(n29709), .B(n29708), .Z(n29713) );
  IV U42655 ( .A(n29709), .Z(n29712) );
  IV U42656 ( .A(n29710), .Z(n29711) );
  NOR U42657 ( .A(n29712), .B(n29711), .Z(n35531) );
  NOR U42658 ( .A(n29713), .B(n35531), .Z(n29714) );
  IV U42659 ( .A(n29714), .Z(n33098) );
  XOR U42660 ( .A(n29715), .B(n33098), .Z(n35506) );
  XOR U42661 ( .A(n32196), .B(n35506), .Z(n32189) );
  XOR U42662 ( .A(n29716), .B(n32189), .Z(n32183) );
  XOR U42663 ( .A(n32184), .B(n32183), .Z(n32186) );
  IV U42664 ( .A(n29717), .Z(n29718) );
  NOR U42665 ( .A(n29719), .B(n29718), .Z(n32185) );
  IV U42666 ( .A(n29720), .Z(n29723) );
  IV U42667 ( .A(n29721), .Z(n29722) );
  NOR U42668 ( .A(n29723), .B(n29722), .Z(n33109) );
  NOR U42669 ( .A(n32181), .B(n33109), .Z(n29724) );
  IV U42670 ( .A(n29724), .Z(n29725) );
  NOR U42671 ( .A(n32185), .B(n29725), .Z(n29726) );
  XOR U42672 ( .A(n32186), .B(n29726), .Z(n33108) );
  XOR U42673 ( .A(n33106), .B(n33108), .Z(n39800) );
  IV U42674 ( .A(n39800), .Z(n29732) );
  IV U42675 ( .A(n29727), .Z(n29728) );
  NOR U42676 ( .A(n29731), .B(n29728), .Z(n39795) );
  IV U42677 ( .A(n29729), .Z(n29730) );
  NOR U42678 ( .A(n29731), .B(n29730), .Z(n39803) );
  NOR U42679 ( .A(n39795), .B(n39803), .Z(n33114) );
  XOR U42680 ( .A(n29732), .B(n33114), .Z(n33116) );
  XOR U42681 ( .A(n33115), .B(n33116), .Z(n32180) );
  XOR U42682 ( .A(n32179), .B(n32180), .Z(n29735) );
  IV U42683 ( .A(n29735), .Z(n29733) );
  NOR U42684 ( .A(n29734), .B(n29733), .Z(n35487) );
  NOR U42685 ( .A(n29737), .B(n29739), .Z(n29736) );
  NOR U42686 ( .A(n29736), .B(n29735), .Z(n29741) );
  NOR U42687 ( .A(n29737), .B(n32180), .Z(n29738) );
  IV U42688 ( .A(n29738), .Z(n33121) );
  NOR U42689 ( .A(n33121), .B(n29739), .Z(n29740) );
  NOR U42690 ( .A(n29741), .B(n29740), .Z(n29742) );
  NOR U42691 ( .A(n29743), .B(n29742), .Z(n29744) );
  NOR U42692 ( .A(n35487), .B(n29744), .Z(n32174) );
  XOR U42693 ( .A(n29745), .B(n32174), .Z(n33133) );
  XOR U42694 ( .A(n33131), .B(n33133), .Z(n33142) );
  XOR U42695 ( .A(n33141), .B(n33142), .Z(n32171) );
  IV U42696 ( .A(n29746), .Z(n29747) );
  NOR U42697 ( .A(n29748), .B(n29747), .Z(n32169) );
  XOR U42698 ( .A(n32171), .B(n32169), .Z(n33139) );
  IV U42699 ( .A(n29749), .Z(n29750) );
  NOR U42700 ( .A(n29751), .B(n29750), .Z(n32164) );
  IV U42701 ( .A(n29752), .Z(n29754) );
  NOR U42702 ( .A(n29754), .B(n29753), .Z(n33137) );
  NOR U42703 ( .A(n32164), .B(n33137), .Z(n29755) );
  XOR U42704 ( .A(n33139), .B(n29755), .Z(n32160) );
  XOR U42705 ( .A(n29756), .B(n32160), .Z(n33164) );
  XOR U42706 ( .A(n29757), .B(n33164), .Z(n32151) );
  XOR U42707 ( .A(n32152), .B(n32151), .Z(n29758) );
  XOR U42708 ( .A(n29759), .B(n29758), .Z(n32145) );
  XOR U42709 ( .A(n29760), .B(n32145), .Z(n32144) );
  XOR U42710 ( .A(n29761), .B(n32144), .Z(n32139) );
  IV U42711 ( .A(n29762), .Z(n33179) );
  NOR U42712 ( .A(n33179), .B(n29763), .Z(n29767) );
  IV U42713 ( .A(n29764), .Z(n29766) );
  NOR U42714 ( .A(n29766), .B(n29765), .Z(n32138) );
  NOR U42715 ( .A(n29767), .B(n32138), .Z(n29768) );
  XOR U42716 ( .A(n32139), .B(n29768), .Z(n32135) );
  IV U42717 ( .A(n29769), .Z(n29771) );
  IV U42718 ( .A(n29770), .Z(n29779) );
  NOR U42719 ( .A(n29771), .B(n29779), .Z(n29776) );
  IV U42720 ( .A(n29776), .Z(n29772) );
  NOR U42721 ( .A(n32135), .B(n29772), .Z(n36563) );
  NOR U42722 ( .A(n29773), .B(n32134), .Z(n29774) );
  XOR U42723 ( .A(n29774), .B(n32135), .Z(n50097) );
  IV U42724 ( .A(n50097), .Z(n29775) );
  NOR U42725 ( .A(n29776), .B(n29775), .Z(n29777) );
  NOR U42726 ( .A(n36563), .B(n29777), .Z(n32131) );
  IV U42727 ( .A(n29778), .Z(n29780) );
  NOR U42728 ( .A(n29780), .B(n29779), .Z(n33196) );
  IV U42729 ( .A(n29781), .Z(n29783) );
  NOR U42730 ( .A(n29783), .B(n29782), .Z(n33192) );
  NOR U42731 ( .A(n33196), .B(n33192), .Z(n32132) );
  XOR U42732 ( .A(n32131), .B(n32132), .Z(n33202) );
  XOR U42733 ( .A(n33201), .B(n33202), .Z(n33206) );
  XOR U42734 ( .A(n33204), .B(n33206), .Z(n32125) );
  XOR U42735 ( .A(n29784), .B(n32125), .Z(n29785) );
  IV U42736 ( .A(n29785), .Z(n32121) );
  XOR U42737 ( .A(n32119), .B(n32121), .Z(n32117) );
  XOR U42738 ( .A(n32116), .B(n32117), .Z(n33215) );
  IV U42739 ( .A(n29786), .Z(n29789) );
  IV U42740 ( .A(n29787), .Z(n29788) );
  NOR U42741 ( .A(n29789), .B(n29788), .Z(n33213) );
  XOR U42742 ( .A(n33215), .B(n33213), .Z(n35416) );
  IV U42743 ( .A(n29790), .Z(n29791) );
  NOR U42744 ( .A(n29797), .B(n29791), .Z(n32114) );
  IV U42745 ( .A(n29792), .Z(n29794) );
  NOR U42746 ( .A(n29794), .B(n29793), .Z(n35414) );
  IV U42747 ( .A(n29795), .Z(n29796) );
  NOR U42748 ( .A(n29797), .B(n29796), .Z(n35419) );
  NOR U42749 ( .A(n35414), .B(n35419), .Z(n32113) );
  IV U42750 ( .A(n32113), .Z(n29798) );
  NOR U42751 ( .A(n32114), .B(n29798), .Z(n29799) );
  XOR U42752 ( .A(n35416), .B(n29799), .Z(n32108) );
  XOR U42753 ( .A(n32107), .B(n32108), .Z(n36585) );
  XOR U42754 ( .A(n36576), .B(n36585), .Z(n32105) );
  XOR U42755 ( .A(n29800), .B(n32105), .Z(n29801) );
  IV U42756 ( .A(n29801), .Z(n32097) );
  XOR U42757 ( .A(n32095), .B(n32097), .Z(n33230) );
  IV U42758 ( .A(n29802), .Z(n29803) );
  NOR U42759 ( .A(n29803), .B(n29807), .Z(n32089) );
  IV U42760 ( .A(n29804), .Z(n32092) );
  NOR U42761 ( .A(n32092), .B(n29805), .Z(n29809) );
  IV U42762 ( .A(n29806), .Z(n29808) );
  NOR U42763 ( .A(n29808), .B(n29807), .Z(n33229) );
  NOR U42764 ( .A(n29809), .B(n33229), .Z(n29810) );
  IV U42765 ( .A(n29810), .Z(n29811) );
  NOR U42766 ( .A(n32089), .B(n29811), .Z(n29812) );
  XOR U42767 ( .A(n33230), .B(n29812), .Z(n32086) );
  IV U42768 ( .A(n29813), .Z(n29822) );
  IV U42769 ( .A(n29814), .Z(n29815) );
  NOR U42770 ( .A(n29822), .B(n29815), .Z(n33235) );
  IV U42771 ( .A(n29816), .Z(n29818) );
  NOR U42772 ( .A(n29818), .B(n29817), .Z(n32087) );
  NOR U42773 ( .A(n33235), .B(n32087), .Z(n29819) );
  XOR U42774 ( .A(n32086), .B(n29819), .Z(n33233) );
  IV U42775 ( .A(n29820), .Z(n29821) );
  NOR U42776 ( .A(n29822), .B(n29821), .Z(n33232) );
  IV U42777 ( .A(n29823), .Z(n29825) );
  NOR U42778 ( .A(n29825), .B(n29824), .Z(n32084) );
  NOR U42779 ( .A(n33232), .B(n32084), .Z(n29826) );
  XOR U42780 ( .A(n33233), .B(n29826), .Z(n32080) );
  XOR U42781 ( .A(n32081), .B(n32080), .Z(n29829) );
  IV U42782 ( .A(n29829), .Z(n29827) );
  NOR U42783 ( .A(n29828), .B(n29827), .Z(n35394) );
  NOR U42784 ( .A(n29830), .B(n29829), .Z(n33241) );
  IV U42785 ( .A(n29837), .Z(n29835) );
  IV U42786 ( .A(n29831), .Z(n29838) );
  NOR U42787 ( .A(n29835), .B(n29838), .Z(n33239) );
  XOR U42788 ( .A(n33241), .B(n33239), .Z(n29832) );
  NOR U42789 ( .A(n35394), .B(n29832), .Z(n29842) );
  IV U42790 ( .A(n29833), .Z(n29834) );
  NOR U42791 ( .A(n29835), .B(n29834), .Z(n32076) );
  IV U42792 ( .A(n29836), .Z(n29840) );
  XOR U42793 ( .A(n29838), .B(n29837), .Z(n29839) );
  NOR U42794 ( .A(n29840), .B(n29839), .Z(n32073) );
  NOR U42795 ( .A(n32076), .B(n32073), .Z(n29841) );
  XOR U42796 ( .A(n29842), .B(n29841), .Z(n32070) );
  IV U42797 ( .A(n29843), .Z(n29845) );
  NOR U42798 ( .A(n29845), .B(n29844), .Z(n32068) );
  XOR U42799 ( .A(n32070), .B(n32068), .Z(n32071) );
  NOR U42800 ( .A(n29846), .B(n32065), .Z(n29870) );
  IV U42801 ( .A(n29847), .Z(n29852) );
  IV U42802 ( .A(n29848), .Z(n29849) );
  NOR U42803 ( .A(n29852), .B(n29849), .Z(n29867) );
  IV U42804 ( .A(n29867), .Z(n32072) );
  IV U42805 ( .A(n29850), .Z(n29851) );
  NOR U42806 ( .A(n29852), .B(n29851), .Z(n29868) );
  IV U42807 ( .A(n29868), .Z(n32063) );
  XOR U42808 ( .A(n32072), .B(n32063), .Z(n29853) );
  NOR U42809 ( .A(n29870), .B(n29853), .Z(n29854) );
  XOR U42810 ( .A(n32071), .B(n29854), .Z(n29863) );
  IV U42811 ( .A(n29863), .Z(n29859) );
  IV U42812 ( .A(n29855), .Z(n29857) );
  NOR U42813 ( .A(n29857), .B(n29856), .Z(n29882) );
  IV U42814 ( .A(n29882), .Z(n29858) );
  NOR U42815 ( .A(n29859), .B(n29858), .Z(n35385) );
  NOR U42816 ( .A(n29861), .B(n29860), .Z(n29862) );
  NOR U42817 ( .A(n29863), .B(n29862), .Z(n29881) );
  IV U42818 ( .A(n29864), .Z(n29875) );
  IV U42819 ( .A(n32065), .Z(n29866) );
  NOR U42820 ( .A(n29866), .B(n29865), .Z(n29873) );
  XOR U42821 ( .A(n29867), .B(n32071), .Z(n32062) );
  XOR U42822 ( .A(n29868), .B(n32062), .Z(n29869) );
  NOR U42823 ( .A(n29870), .B(n29869), .Z(n29871) );
  IV U42824 ( .A(n29871), .Z(n29872) );
  NOR U42825 ( .A(n29873), .B(n29872), .Z(n29874) );
  IV U42826 ( .A(n29874), .Z(n29877) );
  NOR U42827 ( .A(n29875), .B(n29877), .Z(n33254) );
  IV U42828 ( .A(n29876), .Z(n29878) );
  NOR U42829 ( .A(n29878), .B(n29877), .Z(n35389) );
  NOR U42830 ( .A(n33254), .B(n35389), .Z(n29879) );
  IV U42831 ( .A(n29879), .Z(n29880) );
  NOR U42832 ( .A(n29881), .B(n29880), .Z(n33262) );
  NOR U42833 ( .A(n29882), .B(n33262), .Z(n29883) );
  NOR U42834 ( .A(n35385), .B(n29883), .Z(n32051) );
  IV U42835 ( .A(n29884), .Z(n29885) );
  NOR U42836 ( .A(n29886), .B(n29885), .Z(n32060) );
  NOR U42837 ( .A(n32060), .B(n33269), .Z(n29887) );
  XOR U42838 ( .A(n32051), .B(n29887), .Z(n32048) );
  NOR U42839 ( .A(n29888), .B(n32052), .Z(n29892) );
  IV U42840 ( .A(n29889), .Z(n32045) );
  NOR U42841 ( .A(n29890), .B(n32045), .Z(n29891) );
  NOR U42842 ( .A(n29892), .B(n29891), .Z(n29893) );
  XOR U42843 ( .A(n32048), .B(n29893), .Z(n32033) );
  NOR U42844 ( .A(n29894), .B(n32034), .Z(n29901) );
  IV U42845 ( .A(n29895), .Z(n29897) );
  IV U42846 ( .A(n29896), .Z(n29898) );
  NOR U42847 ( .A(n29897), .B(n29898), .Z(n35370) );
  NOR U42848 ( .A(n29899), .B(n29898), .Z(n36639) );
  NOR U42849 ( .A(n35370), .B(n36639), .Z(n33287) );
  IV U42850 ( .A(n33287), .Z(n29900) );
  NOR U42851 ( .A(n29901), .B(n29900), .Z(n29902) );
  XOR U42852 ( .A(n32033), .B(n29902), .Z(n33299) );
  XOR U42853 ( .A(n33289), .B(n33299), .Z(n33292) );
  IV U42854 ( .A(n29903), .Z(n33300) );
  NOR U42855 ( .A(n29904), .B(n33300), .Z(n29907) );
  IV U42856 ( .A(n29905), .Z(n29906) );
  NOR U42857 ( .A(n29906), .B(n29914), .Z(n32030) );
  NOR U42858 ( .A(n29907), .B(n32030), .Z(n29908) );
  XOR U42859 ( .A(n33292), .B(n29908), .Z(n29909) );
  IV U42860 ( .A(n29909), .Z(n32029) );
  IV U42861 ( .A(n29910), .Z(n29911) );
  NOR U42862 ( .A(n29911), .B(n29917), .Z(n29912) );
  IV U42863 ( .A(n29912), .Z(n29920) );
  NOR U42864 ( .A(n32029), .B(n29920), .Z(n36653) );
  IV U42865 ( .A(n29913), .Z(n29915) );
  NOR U42866 ( .A(n29915), .B(n29914), .Z(n32027) );
  IV U42867 ( .A(n29916), .Z(n29918) );
  NOR U42868 ( .A(n29918), .B(n29917), .Z(n32025) );
  NOR U42869 ( .A(n32027), .B(n32025), .Z(n29919) );
  XOR U42870 ( .A(n32029), .B(n29919), .Z(n29922) );
  NOR U42871 ( .A(n32025), .B(n29920), .Z(n29921) );
  NOR U42872 ( .A(n29922), .B(n29921), .Z(n33307) );
  NOR U42873 ( .A(n36653), .B(n33307), .Z(n32022) );
  XOR U42874 ( .A(n29923), .B(n32022), .Z(n32021) );
  IV U42875 ( .A(n29924), .Z(n29925) );
  NOR U42876 ( .A(n29925), .B(n29934), .Z(n29931) );
  IV U42877 ( .A(n29931), .Z(n29926) );
  NOR U42878 ( .A(n32021), .B(n29926), .Z(n35362) );
  IV U42879 ( .A(n29927), .Z(n29928) );
  NOR U42880 ( .A(n29929), .B(n29928), .Z(n32019) );
  XOR U42881 ( .A(n32019), .B(n32021), .Z(n32017) );
  IV U42882 ( .A(n32017), .Z(n29930) );
  NOR U42883 ( .A(n29931), .B(n29930), .Z(n29932) );
  NOR U42884 ( .A(n35362), .B(n29932), .Z(n29940) );
  IV U42885 ( .A(n29933), .Z(n29935) );
  NOR U42886 ( .A(n29935), .B(n29934), .Z(n32016) );
  IV U42887 ( .A(n29936), .Z(n32013) );
  NOR U42888 ( .A(n29937), .B(n32013), .Z(n29938) );
  NOR U42889 ( .A(n32016), .B(n29938), .Z(n29941) );
  IV U42890 ( .A(n29941), .Z(n29939) );
  NOR U42891 ( .A(n29940), .B(n29939), .Z(n29943) );
  NOR U42892 ( .A(n29941), .B(n32017), .Z(n29942) );
  NOR U42893 ( .A(n29943), .B(n29942), .Z(n29944) );
  IV U42894 ( .A(n29944), .Z(n33317) );
  IV U42895 ( .A(n29945), .Z(n29947) );
  NOR U42896 ( .A(n29947), .B(n29946), .Z(n29948) );
  IV U42897 ( .A(n29948), .Z(n32011) );
  XOR U42898 ( .A(n33317), .B(n32011), .Z(n29949) );
  XOR U42899 ( .A(n29950), .B(n29949), .Z(n36701) );
  IV U42900 ( .A(n36701), .Z(n29961) );
  XOR U42901 ( .A(n32010), .B(n29961), .Z(n29951) );
  NOR U42902 ( .A(n29952), .B(n29951), .Z(n36712) );
  IV U42903 ( .A(n29953), .Z(n29954) );
  NOR U42904 ( .A(n29954), .B(n29957), .Z(n29955) );
  IV U42905 ( .A(n29955), .Z(n32009) );
  IV U42906 ( .A(n29956), .Z(n29958) );
  NOR U42907 ( .A(n29958), .B(n29957), .Z(n33323) );
  NOR U42908 ( .A(n29959), .B(n33323), .Z(n29960) );
  XOR U42909 ( .A(n29961), .B(n29960), .Z(n32008) );
  XOR U42910 ( .A(n32009), .B(n32008), .Z(n29962) );
  NOR U42911 ( .A(n29963), .B(n29962), .Z(n29964) );
  NOR U42912 ( .A(n36712), .B(n29964), .Z(n29965) );
  IV U42913 ( .A(n29965), .Z(n32007) );
  XOR U42914 ( .A(n32005), .B(n32007), .Z(n31995) );
  NOR U42915 ( .A(n29966), .B(n31995), .Z(n33331) );
  NOR U42916 ( .A(n29967), .B(n31999), .Z(n29968) );
  XOR U42917 ( .A(n29968), .B(n31995), .Z(n31992) );
  IV U42918 ( .A(n31992), .Z(n29969) );
  NOR U42919 ( .A(n29970), .B(n29969), .Z(n29971) );
  NOR U42920 ( .A(n33331), .B(n29971), .Z(n29977) );
  IV U42921 ( .A(n29972), .Z(n29974) );
  NOR U42922 ( .A(n29974), .B(n29973), .Z(n31994) );
  IV U42923 ( .A(n29980), .Z(n29975) );
  NOR U42924 ( .A(n29975), .B(n29979), .Z(n31991) );
  NOR U42925 ( .A(n31994), .B(n31991), .Z(n29976) );
  XOR U42926 ( .A(n29977), .B(n29976), .Z(n31990) );
  XOR U42927 ( .A(n31989), .B(n31990), .Z(n29986) );
  IV U42928 ( .A(n29986), .Z(n29984) );
  IV U42929 ( .A(n29978), .Z(n29982) );
  XOR U42930 ( .A(n29980), .B(n29979), .Z(n29981) );
  NOR U42931 ( .A(n29982), .B(n29981), .Z(n29985) );
  IV U42932 ( .A(n29985), .Z(n29983) );
  NOR U42933 ( .A(n29984), .B(n29983), .Z(n35349) );
  NOR U42934 ( .A(n29986), .B(n29985), .Z(n31988) );
  IV U42935 ( .A(n29987), .Z(n29990) );
  IV U42936 ( .A(n29988), .Z(n29989) );
  NOR U42937 ( .A(n29990), .B(n29989), .Z(n31986) );
  XOR U42938 ( .A(n31988), .B(n31986), .Z(n29991) );
  NOR U42939 ( .A(n35349), .B(n29991), .Z(n30000) );
  IV U42940 ( .A(n30000), .Z(n33343) );
  NOR U42941 ( .A(n29999), .B(n33343), .Z(n36730) );
  NOR U42942 ( .A(n35340), .B(n29992), .Z(n29997) );
  IV U42943 ( .A(n29997), .Z(n29994) );
  NOR U42944 ( .A(n31988), .B(n35349), .Z(n29993) );
  IV U42945 ( .A(n29993), .Z(n35336) );
  NOR U42946 ( .A(n29994), .B(n35336), .Z(n29995) );
  NOR U42947 ( .A(n36730), .B(n29995), .Z(n29996) );
  IV U42948 ( .A(n29996), .Z(n33340) );
  NOR U42949 ( .A(n29997), .B(n30000), .Z(n29998) );
  NOR U42950 ( .A(n33340), .B(n29998), .Z(n30002) );
  NOR U42951 ( .A(n30000), .B(n29999), .Z(n30001) );
  NOR U42952 ( .A(n30002), .B(n30001), .Z(n33346) );
  IV U42953 ( .A(n33349), .Z(n30004) );
  NOR U42954 ( .A(n30004), .B(n30003), .Z(n33342) );
  IV U42955 ( .A(n30005), .Z(n30006) );
  NOR U42956 ( .A(n30006), .B(n30009), .Z(n30007) );
  NOR U42957 ( .A(n33342), .B(n30007), .Z(n33345) );
  XOR U42958 ( .A(n33346), .B(n33345), .Z(n31975) );
  IV U42959 ( .A(n30008), .Z(n30010) );
  NOR U42960 ( .A(n30010), .B(n30009), .Z(n31983) );
  NOR U42961 ( .A(n31978), .B(n31976), .Z(n30011) );
  NOR U42962 ( .A(n31983), .B(n30011), .Z(n30012) );
  XOR U42963 ( .A(n31975), .B(n30012), .Z(n35319) );
  NOR U42964 ( .A(n30013), .B(n35319), .Z(n36743) );
  IV U42965 ( .A(n30014), .Z(n35322) );
  NOR U42966 ( .A(n30015), .B(n35322), .Z(n31979) );
  IV U42967 ( .A(n30022), .Z(n30016) );
  NOR U42968 ( .A(n30016), .B(n30021), .Z(n31973) );
  NOR U42969 ( .A(n31979), .B(n31973), .Z(n30017) );
  XOR U42970 ( .A(n30017), .B(n35319), .Z(n33360) );
  NOR U42971 ( .A(n30018), .B(n33360), .Z(n30019) );
  NOR U42972 ( .A(n36743), .B(n30019), .Z(n33355) );
  IV U42973 ( .A(n30020), .Z(n30024) );
  XOR U42974 ( .A(n30022), .B(n30021), .Z(n30023) );
  NOR U42975 ( .A(n30024), .B(n30023), .Z(n30025) );
  IV U42976 ( .A(n30025), .Z(n33356) );
  XOR U42977 ( .A(n33355), .B(n33356), .Z(n31971) );
  IV U42978 ( .A(n31971), .Z(n30034) );
  IV U42979 ( .A(n30026), .Z(n30027) );
  NOR U42980 ( .A(n30028), .B(n30027), .Z(n31970) );
  IV U42981 ( .A(n30029), .Z(n30032) );
  IV U42982 ( .A(n30030), .Z(n30031) );
  NOR U42983 ( .A(n30032), .B(n30031), .Z(n33361) );
  NOR U42984 ( .A(n31970), .B(n33361), .Z(n30033) );
  XOR U42985 ( .A(n30034), .B(n30033), .Z(n31967) );
  XOR U42986 ( .A(n30035), .B(n31967), .Z(n33367) );
  NOR U42987 ( .A(n30036), .B(n31959), .Z(n30040) );
  IV U42988 ( .A(n30037), .Z(n30039) );
  IV U42989 ( .A(n30038), .Z(n30045) );
  NOR U42990 ( .A(n30039), .B(n30045), .Z(n33366) );
  NOR U42991 ( .A(n30040), .B(n33366), .Z(n30041) );
  XOR U42992 ( .A(n33367), .B(n30041), .Z(n31955) );
  IV U42993 ( .A(n30042), .Z(n30043) );
  NOR U42994 ( .A(n30043), .B(n30048), .Z(n33369) );
  IV U42995 ( .A(n30044), .Z(n30046) );
  NOR U42996 ( .A(n30046), .B(n30045), .Z(n31956) );
  IV U42997 ( .A(n30047), .Z(n30049) );
  NOR U42998 ( .A(n30049), .B(n30048), .Z(n33371) );
  NOR U42999 ( .A(n31956), .B(n33371), .Z(n30050) );
  IV U43000 ( .A(n30050), .Z(n30051) );
  NOR U43001 ( .A(n33369), .B(n30051), .Z(n30052) );
  XOR U43002 ( .A(n31955), .B(n30052), .Z(n35296) );
  IV U43003 ( .A(n30053), .Z(n30055) );
  NOR U43004 ( .A(n30055), .B(n30054), .Z(n31953) );
  XOR U43005 ( .A(n35296), .B(n31953), .Z(n31947) );
  IV U43006 ( .A(n31947), .Z(n30061) );
  IV U43007 ( .A(n30056), .Z(n35299) );
  NOR U43008 ( .A(n35299), .B(n30057), .Z(n31951) );
  NOR U43009 ( .A(n30058), .B(n31948), .Z(n30059) );
  NOR U43010 ( .A(n31951), .B(n30059), .Z(n30060) );
  XOR U43011 ( .A(n30061), .B(n30060), .Z(n35285) );
  IV U43012 ( .A(n30062), .Z(n30064) );
  NOR U43013 ( .A(n30064), .B(n30063), .Z(n31943) );
  XOR U43014 ( .A(n35285), .B(n31943), .Z(n33377) );
  XOR U43015 ( .A(n33376), .B(n33377), .Z(n31937) );
  XOR U43016 ( .A(n30065), .B(n31937), .Z(n31929) );
  XOR U43017 ( .A(n30066), .B(n31929), .Z(n31927) );
  XOR U43018 ( .A(n31926), .B(n31927), .Z(n33393) );
  XOR U43019 ( .A(n30067), .B(n33393), .Z(n33402) );
  NOR U43020 ( .A(n30068), .B(n33402), .Z(n35266) );
  NOR U43021 ( .A(n30069), .B(n33394), .Z(n30072) );
  IV U43022 ( .A(n30072), .Z(n30070) );
  NOR U43023 ( .A(n30070), .B(n33393), .Z(n33398) );
  IV U43024 ( .A(n33402), .Z(n30071) );
  NOR U43025 ( .A(n30072), .B(n30071), .Z(n30073) );
  NOR U43026 ( .A(n33398), .B(n30073), .Z(n33405) );
  NOR U43027 ( .A(n30074), .B(n33405), .Z(n30075) );
  NOR U43028 ( .A(n35266), .B(n30075), .Z(n30085) );
  IV U43029 ( .A(n30076), .Z(n30078) );
  NOR U43030 ( .A(n30078), .B(n30077), .Z(n33401) );
  IV U43031 ( .A(n30079), .Z(n30083) );
  XOR U43032 ( .A(n30081), .B(n30080), .Z(n30082) );
  NOR U43033 ( .A(n30083), .B(n30082), .Z(n33406) );
  NOR U43034 ( .A(n33401), .B(n33406), .Z(n30084) );
  XOR U43035 ( .A(n30085), .B(n30084), .Z(n31918) );
  IV U43036 ( .A(n30086), .Z(n30088) );
  NOR U43037 ( .A(n30088), .B(n30087), .Z(n31916) );
  XOR U43038 ( .A(n31918), .B(n31916), .Z(n30091) );
  NOR U43039 ( .A(n30089), .B(n30091), .Z(n43580) );
  NOR U43040 ( .A(n31910), .B(n30090), .Z(n30092) );
  XOR U43041 ( .A(n30092), .B(n30091), .Z(n31904) );
  IV U43042 ( .A(n31904), .Z(n30093) );
  NOR U43043 ( .A(n30094), .B(n30093), .Z(n30095) );
  NOR U43044 ( .A(n43580), .B(n30095), .Z(n30101) );
  NOR U43045 ( .A(n30096), .B(n31905), .Z(n30097) );
  NOR U43046 ( .A(n30101), .B(n30097), .Z(n30100) );
  IV U43047 ( .A(n30097), .Z(n30098) );
  NOR U43048 ( .A(n30098), .B(n31904), .Z(n30099) );
  NOR U43049 ( .A(n30100), .B(n30099), .Z(n30109) );
  NOR U43050 ( .A(n30102), .B(n30109), .Z(n31898) );
  IV U43051 ( .A(n30101), .Z(n36825) );
  IV U43052 ( .A(n30102), .Z(n30103) );
  NOR U43053 ( .A(n36825), .B(n30103), .Z(n30104) );
  NOR U43054 ( .A(n31898), .B(n30104), .Z(n30115) );
  IV U43055 ( .A(n30115), .Z(n30108) );
  IV U43056 ( .A(n30105), .Z(n30106) );
  NOR U43057 ( .A(n30106), .B(n30111), .Z(n30118) );
  IV U43058 ( .A(n30118), .Z(n30107) );
  NOR U43059 ( .A(n30108), .B(n30107), .Z(n35250) );
  IV U43060 ( .A(n30109), .Z(n30114) );
  IV U43061 ( .A(n30110), .Z(n30112) );
  NOR U43062 ( .A(n30112), .B(n30111), .Z(n30116) );
  IV U43063 ( .A(n30116), .Z(n30113) );
  NOR U43064 ( .A(n30114), .B(n30113), .Z(n35252) );
  NOR U43065 ( .A(n30116), .B(n30115), .Z(n30117) );
  NOR U43066 ( .A(n35252), .B(n30117), .Z(n30119) );
  NOR U43067 ( .A(n30119), .B(n30118), .Z(n30120) );
  NOR U43068 ( .A(n35250), .B(n30120), .Z(n31897) );
  IV U43069 ( .A(n31897), .Z(n31900) );
  XOR U43070 ( .A(n31899), .B(n31900), .Z(n33429) );
  IV U43071 ( .A(n33429), .Z(n30128) );
  IV U43072 ( .A(n30121), .Z(n31894) );
  NOR U43073 ( .A(n31894), .B(n30122), .Z(n30126) );
  IV U43074 ( .A(n30123), .Z(n30125) );
  NOR U43075 ( .A(n30125), .B(n30124), .Z(n33428) );
  NOR U43076 ( .A(n30126), .B(n33428), .Z(n30127) );
  XOR U43077 ( .A(n30128), .B(n30127), .Z(n31891) );
  XOR U43078 ( .A(n31889), .B(n31891), .Z(n33443) );
  XOR U43079 ( .A(n33442), .B(n33443), .Z(n33440) );
  IV U43080 ( .A(n30129), .Z(n30130) );
  NOR U43081 ( .A(n30145), .B(n30130), .Z(n30140) );
  IV U43082 ( .A(n30140), .Z(n30131) );
  NOR U43083 ( .A(n33440), .B(n30131), .Z(n35240) );
  IV U43084 ( .A(n30132), .Z(n30134) );
  IV U43085 ( .A(n30133), .Z(n30137) );
  NOR U43086 ( .A(n30134), .B(n30137), .Z(n30135) );
  IV U43087 ( .A(n30135), .Z(n31888) );
  IV U43088 ( .A(n30136), .Z(n30138) );
  NOR U43089 ( .A(n30138), .B(n30137), .Z(n33438) );
  XOR U43090 ( .A(n33440), .B(n33438), .Z(n31887) );
  XOR U43091 ( .A(n31888), .B(n31887), .Z(n30139) );
  NOR U43092 ( .A(n30140), .B(n30139), .Z(n30141) );
  NOR U43093 ( .A(n35240), .B(n30141), .Z(n30142) );
  IV U43094 ( .A(n30142), .Z(n31886) );
  IV U43095 ( .A(n30143), .Z(n30144) );
  NOR U43096 ( .A(n30145), .B(n30144), .Z(n31884) );
  XOR U43097 ( .A(n31886), .B(n31884), .Z(n33460) );
  XOR U43098 ( .A(n33454), .B(n33460), .Z(n31876) );
  XOR U43099 ( .A(n30146), .B(n31876), .Z(n33475) );
  XOR U43100 ( .A(n30147), .B(n33475), .Z(n33472) );
  XOR U43101 ( .A(n33471), .B(n33472), .Z(n31867) );
  XOR U43102 ( .A(n31868), .B(n31867), .Z(n30149) );
  NOR U43103 ( .A(n30148), .B(n30149), .Z(n31866) );
  IV U43104 ( .A(n30148), .Z(n30151) );
  IV U43105 ( .A(n30149), .Z(n30150) );
  NOR U43106 ( .A(n30151), .B(n30150), .Z(n36890) );
  NOR U43107 ( .A(n31866), .B(n36890), .Z(n31861) );
  IV U43108 ( .A(n30152), .Z(n30153) );
  NOR U43109 ( .A(n30160), .B(n30153), .Z(n31862) );
  IV U43110 ( .A(n30154), .Z(n30156) );
  NOR U43111 ( .A(n30156), .B(n30155), .Z(n31864) );
  NOR U43112 ( .A(n31862), .B(n31864), .Z(n30157) );
  XOR U43113 ( .A(n31861), .B(n30157), .Z(n33492) );
  IV U43114 ( .A(n30158), .Z(n30159) );
  NOR U43115 ( .A(n30160), .B(n30159), .Z(n33482) );
  XOR U43116 ( .A(n33492), .B(n33482), .Z(n31856) );
  XOR U43117 ( .A(n30161), .B(n31856), .Z(n33499) );
  XOR U43118 ( .A(n30162), .B(n33499), .Z(n31838) );
  XOR U43119 ( .A(n30163), .B(n31838), .Z(n33523) );
  XOR U43120 ( .A(n30164), .B(n33523), .Z(n33537) );
  IV U43121 ( .A(n30165), .Z(n30167) );
  NOR U43122 ( .A(n30167), .B(n30166), .Z(n31831) );
  XOR U43123 ( .A(n33537), .B(n31831), .Z(n30168) );
  XOR U43124 ( .A(n30169), .B(n30168), .Z(n31825) );
  XOR U43125 ( .A(n30170), .B(n31825), .Z(n31824) );
  XOR U43126 ( .A(n30171), .B(n31824), .Z(n31811) );
  IV U43127 ( .A(n30172), .Z(n30173) );
  NOR U43128 ( .A(n30174), .B(n30173), .Z(n31817) );
  IV U43129 ( .A(n30175), .Z(n30176) );
  NOR U43130 ( .A(n30176), .B(n31813), .Z(n31810) );
  NOR U43131 ( .A(n31817), .B(n31810), .Z(n30177) );
  XOR U43132 ( .A(n31811), .B(n30177), .Z(n33547) );
  XOR U43133 ( .A(n33539), .B(n33547), .Z(n33554) );
  IV U43134 ( .A(n30178), .Z(n33546) );
  NOR U43135 ( .A(n30179), .B(n33546), .Z(n30183) );
  IV U43136 ( .A(n30180), .Z(n30182) );
  NOR U43137 ( .A(n30182), .B(n30181), .Z(n33553) );
  NOR U43138 ( .A(n30183), .B(n33553), .Z(n30184) );
  XOR U43139 ( .A(n33554), .B(n30184), .Z(n31807) );
  XOR U43140 ( .A(n33559), .B(n31807), .Z(n33557) );
  XOR U43141 ( .A(n33556), .B(n33557), .Z(n31805) );
  NOR U43142 ( .A(n30188), .B(n31805), .Z(n30185) );
  IV U43143 ( .A(n30185), .Z(n30186) );
  NOR U43144 ( .A(n30187), .B(n30186), .Z(n35166) );
  NOR U43145 ( .A(n30189), .B(n30188), .Z(n30191) );
  IV U43146 ( .A(n30190), .Z(n31806) );
  XOR U43147 ( .A(n31806), .B(n31805), .Z(n30196) );
  NOR U43148 ( .A(n30191), .B(n30196), .Z(n30192) );
  NOR U43149 ( .A(n35166), .B(n30192), .Z(n30193) );
  NOR U43150 ( .A(n30201), .B(n30193), .Z(n30206) );
  IV U43151 ( .A(n30194), .Z(n30200) );
  IV U43152 ( .A(n30195), .Z(n30197) );
  IV U43153 ( .A(n30196), .Z(n30203) );
  NOR U43154 ( .A(n30197), .B(n30203), .Z(n30198) );
  IV U43155 ( .A(n30198), .Z(n30199) );
  NOR U43156 ( .A(n30200), .B(n30199), .Z(n35175) );
  IV U43157 ( .A(n30201), .Z(n30202) );
  NOR U43158 ( .A(n30203), .B(n30202), .Z(n35169) );
  NOR U43159 ( .A(n35175), .B(n35169), .Z(n30204) );
  IV U43160 ( .A(n30204), .Z(n30205) );
  NOR U43161 ( .A(n30206), .B(n30205), .Z(n30221) );
  IV U43162 ( .A(n30221), .Z(n35155) );
  NOR U43163 ( .A(n30207), .B(n35158), .Z(n31802) );
  IV U43164 ( .A(n30208), .Z(n30210) );
  NOR U43165 ( .A(n30210), .B(n30209), .Z(n30220) );
  NOR U43166 ( .A(n31802), .B(n30220), .Z(n30211) );
  XOR U43167 ( .A(n35155), .B(n30211), .Z(n30224) );
  IV U43168 ( .A(n30224), .Z(n36993) );
  NOR U43169 ( .A(n30212), .B(n36993), .Z(n36991) );
  IV U43170 ( .A(n30213), .Z(n30215) );
  IV U43171 ( .A(n30214), .Z(n30218) );
  NOR U43172 ( .A(n30215), .B(n30218), .Z(n30216) );
  IV U43173 ( .A(n30216), .Z(n31801) );
  IV U43174 ( .A(n30217), .Z(n30219) );
  NOR U43175 ( .A(n30219), .B(n30218), .Z(n30225) );
  IV U43176 ( .A(n30225), .Z(n30223) );
  IV U43177 ( .A(n30220), .Z(n31804) );
  XOR U43178 ( .A(n31804), .B(n30221), .Z(n30222) );
  NOR U43179 ( .A(n30223), .B(n30222), .Z(n36984) );
  NOR U43180 ( .A(n30225), .B(n30224), .Z(n30226) );
  NOR U43181 ( .A(n36984), .B(n30226), .Z(n30227) );
  IV U43182 ( .A(n30227), .Z(n31800) );
  XOR U43183 ( .A(n31801), .B(n31800), .Z(n30228) );
  NOR U43184 ( .A(n30229), .B(n30228), .Z(n30230) );
  NOR U43185 ( .A(n36991), .B(n30230), .Z(n30241) );
  IV U43186 ( .A(n30231), .Z(n30233) );
  NOR U43187 ( .A(n30233), .B(n30232), .Z(n33570) );
  XOR U43188 ( .A(n30241), .B(n33570), .Z(n30238) );
  IV U43189 ( .A(n30238), .Z(n30234) );
  NOR U43190 ( .A(n30235), .B(n30234), .Z(n35148) );
  IV U43191 ( .A(n30236), .Z(n30242) );
  NOR U43192 ( .A(n30237), .B(n30242), .Z(n30239) );
  NOR U43193 ( .A(n30239), .B(n30238), .Z(n30250) );
  IV U43194 ( .A(n30240), .Z(n30244) );
  IV U43195 ( .A(n30241), .Z(n33571) );
  NOR U43196 ( .A(n30242), .B(n33571), .Z(n30243) );
  IV U43197 ( .A(n30243), .Z(n30246) );
  NOR U43198 ( .A(n30244), .B(n30246), .Z(n35150) );
  IV U43199 ( .A(n30245), .Z(n30247) );
  NOR U43200 ( .A(n30247), .B(n30246), .Z(n35145) );
  NOR U43201 ( .A(n35150), .B(n35145), .Z(n30248) );
  IV U43202 ( .A(n30248), .Z(n30249) );
  NOR U43203 ( .A(n30250), .B(n30249), .Z(n30251) );
  NOR U43204 ( .A(n30252), .B(n30251), .Z(n30253) );
  NOR U43205 ( .A(n35148), .B(n30253), .Z(n30264) );
  IV U43206 ( .A(n30264), .Z(n33575) );
  IV U43207 ( .A(n30254), .Z(n30256) );
  IV U43208 ( .A(n30255), .Z(n30261) );
  NOR U43209 ( .A(n30256), .B(n30261), .Z(n30266) );
  IV U43210 ( .A(n30266), .Z(n30257) );
  NOR U43211 ( .A(n33575), .B(n30257), .Z(n37016) );
  NOR U43212 ( .A(n30259), .B(n30258), .Z(n33579) );
  IV U43213 ( .A(n30260), .Z(n30262) );
  NOR U43214 ( .A(n30262), .B(n30261), .Z(n31798) );
  NOR U43215 ( .A(n33579), .B(n31798), .Z(n30265) );
  IV U43216 ( .A(n30263), .Z(n33576) );
  XOR U43217 ( .A(n33576), .B(n30264), .Z(n33580) );
  XOR U43218 ( .A(n30265), .B(n33580), .Z(n31790) );
  NOR U43219 ( .A(n30266), .B(n31790), .Z(n30267) );
  NOR U43220 ( .A(n37016), .B(n30267), .Z(n33583) );
  XOR U43221 ( .A(n30268), .B(n33583), .Z(n33601) );
  XOR U43222 ( .A(n30269), .B(n33601), .Z(n31774) );
  XOR U43223 ( .A(n30270), .B(n31774), .Z(n35125) );
  XOR U43224 ( .A(n31769), .B(n35125), .Z(n31770) );
  XOR U43225 ( .A(n31772), .B(n31770), .Z(n33618) );
  XOR U43226 ( .A(n33617), .B(n33618), .Z(n31766) );
  XOR U43227 ( .A(n31765), .B(n31766), .Z(n33616) );
  XOR U43228 ( .A(n33614), .B(n33616), .Z(n33634) );
  XOR U43229 ( .A(n31763), .B(n33634), .Z(n33637) );
  XOR U43230 ( .A(n30271), .B(n33637), .Z(n30272) );
  IV U43231 ( .A(n30272), .Z(n35106) );
  IV U43232 ( .A(n30273), .Z(n30274) );
  NOR U43233 ( .A(n30274), .B(n30279), .Z(n31753) );
  IV U43234 ( .A(n31753), .Z(n30275) );
  NOR U43235 ( .A(n35106), .B(n30275), .Z(n37050) );
  IV U43236 ( .A(n30276), .Z(n31756) );
  NOR U43237 ( .A(n30277), .B(n31756), .Z(n30281) );
  IV U43238 ( .A(n30278), .Z(n30280) );
  NOR U43239 ( .A(n30280), .B(n30279), .Z(n35105) );
  NOR U43240 ( .A(n30281), .B(n35105), .Z(n30282) );
  XOR U43241 ( .A(n30282), .B(n35106), .Z(n30287) );
  NOR U43242 ( .A(n31753), .B(n30287), .Z(n30283) );
  NOR U43243 ( .A(n37050), .B(n30283), .Z(n30284) );
  NOR U43244 ( .A(n30285), .B(n30284), .Z(n30297) );
  IV U43245 ( .A(n30286), .Z(n30291) );
  IV U43246 ( .A(n30287), .Z(n30288) );
  NOR U43247 ( .A(n30289), .B(n30288), .Z(n30290) );
  IV U43248 ( .A(n30290), .Z(n30293) );
  NOR U43249 ( .A(n30291), .B(n30293), .Z(n37054) );
  IV U43250 ( .A(n30292), .Z(n30294) );
  NOR U43251 ( .A(n30294), .B(n30293), .Z(n37047) );
  NOR U43252 ( .A(n37054), .B(n37047), .Z(n30295) );
  IV U43253 ( .A(n30295), .Z(n30296) );
  NOR U43254 ( .A(n30297), .B(n30296), .Z(n33648) );
  XOR U43255 ( .A(n30298), .B(n33648), .Z(n33666) );
  XOR U43256 ( .A(n33665), .B(n33666), .Z(n33669) );
  IV U43257 ( .A(n33669), .Z(n30306) );
  IV U43258 ( .A(n30299), .Z(n30301) );
  NOR U43259 ( .A(n30301), .B(n30300), .Z(n33668) );
  IV U43260 ( .A(n30302), .Z(n31748) );
  NOR U43261 ( .A(n30303), .B(n31748), .Z(n30304) );
  NOR U43262 ( .A(n33668), .B(n30304), .Z(n30305) );
  XOR U43263 ( .A(n30306), .B(n30305), .Z(n37073) );
  XOR U43264 ( .A(n31745), .B(n37073), .Z(n35073) );
  NOR U43265 ( .A(n30307), .B(n35073), .Z(n35077) );
  NOR U43266 ( .A(n30314), .B(n35077), .Z(n31736) );
  IV U43267 ( .A(n31736), .Z(n30313) );
  IV U43268 ( .A(n30308), .Z(n31739) );
  NOR U43269 ( .A(n30309), .B(n31739), .Z(n30310) );
  NOR U43270 ( .A(n31745), .B(n30310), .Z(n30311) );
  XOR U43271 ( .A(n37073), .B(n30311), .Z(n30315) );
  NOR U43272 ( .A(n30312), .B(n30315), .Z(n31737) );
  NOR U43273 ( .A(n30313), .B(n31737), .Z(n30317) );
  IV U43274 ( .A(n30314), .Z(n35076) );
  NOR U43275 ( .A(n35076), .B(n30315), .Z(n30316) );
  NOR U43276 ( .A(n30317), .B(n30316), .Z(n31732) );
  XOR U43277 ( .A(n31730), .B(n31732), .Z(n31734) );
  IV U43278 ( .A(n30318), .Z(n30321) );
  IV U43279 ( .A(n30319), .Z(n30320) );
  NOR U43280 ( .A(n30321), .B(n30320), .Z(n30322) );
  IV U43281 ( .A(n30322), .Z(n30330) );
  NOR U43282 ( .A(n31734), .B(n30330), .Z(n37086) );
  IV U43283 ( .A(n30323), .Z(n30324) );
  NOR U43284 ( .A(n30339), .B(n30324), .Z(n30325) );
  IV U43285 ( .A(n30325), .Z(n33686) );
  IV U43286 ( .A(n30326), .Z(n30329) );
  IV U43287 ( .A(n30327), .Z(n30328) );
  NOR U43288 ( .A(n30329), .B(n30328), .Z(n33681) );
  XOR U43289 ( .A(n31733), .B(n31734), .Z(n33682) );
  XOR U43290 ( .A(n33681), .B(n33682), .Z(n33685) );
  XOR U43291 ( .A(n33686), .B(n33685), .Z(n30333) );
  IV U43292 ( .A(n33685), .Z(n30331) );
  NOR U43293 ( .A(n30331), .B(n30330), .Z(n30332) );
  NOR U43294 ( .A(n30333), .B(n30332), .Z(n30334) );
  NOR U43295 ( .A(n37086), .B(n30334), .Z(n30335) );
  IV U43296 ( .A(n30335), .Z(n33688) );
  NOR U43297 ( .A(n30336), .B(n33688), .Z(n35065) );
  IV U43298 ( .A(n30337), .Z(n30338) );
  NOR U43299 ( .A(n30339), .B(n30338), .Z(n33687) );
  XOR U43300 ( .A(n33687), .B(n33688), .Z(n37107) );
  IV U43301 ( .A(n37107), .Z(n30340) );
  NOR U43302 ( .A(n30341), .B(n30340), .Z(n30342) );
  NOR U43303 ( .A(n35065), .B(n30342), .Z(n30343) );
  IV U43304 ( .A(n30343), .Z(n33692) );
  IV U43305 ( .A(n30344), .Z(n30346) );
  NOR U43306 ( .A(n30346), .B(n30345), .Z(n33691) );
  XOR U43307 ( .A(n33692), .B(n33691), .Z(n35058) );
  XOR U43308 ( .A(n30347), .B(n35058), .Z(n30348) );
  IV U43309 ( .A(n30348), .Z(n33703) );
  XOR U43310 ( .A(n33700), .B(n33703), .Z(n33716) );
  IV U43311 ( .A(n30349), .Z(n33704) );
  NOR U43312 ( .A(n33704), .B(n30350), .Z(n30353) );
  IV U43313 ( .A(n30351), .Z(n30352) );
  NOR U43314 ( .A(n30352), .B(n30357), .Z(n33714) );
  NOR U43315 ( .A(n30353), .B(n33714), .Z(n30354) );
  XOR U43316 ( .A(n33716), .B(n30354), .Z(n30355) );
  IV U43317 ( .A(n30355), .Z(n33713) );
  IV U43318 ( .A(n30356), .Z(n30358) );
  NOR U43319 ( .A(n30358), .B(n30357), .Z(n30359) );
  IV U43320 ( .A(n30359), .Z(n33712) );
  XOR U43321 ( .A(n33713), .B(n33712), .Z(n30364) );
  IV U43322 ( .A(n30364), .Z(n35038) );
  NOR U43323 ( .A(n30360), .B(n35038), .Z(n35027) );
  NOR U43324 ( .A(n30362), .B(n30361), .Z(n30365) );
  IV U43325 ( .A(n30365), .Z(n30363) );
  NOR U43326 ( .A(n33713), .B(n30363), .Z(n35041) );
  NOR U43327 ( .A(n30365), .B(n30364), .Z(n30366) );
  NOR U43328 ( .A(n35041), .B(n30366), .Z(n33719) );
  NOR U43329 ( .A(n33719), .B(n30367), .Z(n30368) );
  NOR U43330 ( .A(n35027), .B(n30368), .Z(n33727) );
  NOR U43331 ( .A(n30369), .B(n35033), .Z(n33720) );
  IV U43332 ( .A(n30370), .Z(n30371) );
  NOR U43333 ( .A(n30371), .B(n30374), .Z(n33726) );
  NOR U43334 ( .A(n33720), .B(n33726), .Z(n30372) );
  XOR U43335 ( .A(n33727), .B(n30372), .Z(n33725) );
  IV U43336 ( .A(n30373), .Z(n30375) );
  NOR U43337 ( .A(n30375), .B(n30374), .Z(n33723) );
  XOR U43338 ( .A(n33725), .B(n33723), .Z(n33732) );
  XOR U43339 ( .A(n33731), .B(n33732), .Z(n33739) );
  IV U43340 ( .A(n30376), .Z(n30378) );
  NOR U43341 ( .A(n30378), .B(n30377), .Z(n30386) );
  IV U43342 ( .A(n30386), .Z(n30379) );
  NOR U43343 ( .A(n33739), .B(n30379), .Z(n37136) );
  IV U43344 ( .A(n30380), .Z(n30381) );
  NOR U43345 ( .A(n30384), .B(n30381), .Z(n33734) );
  IV U43346 ( .A(n30382), .Z(n30383) );
  NOR U43347 ( .A(n30384), .B(n30383), .Z(n33737) );
  NOR U43348 ( .A(n33734), .B(n33737), .Z(n30385) );
  XOR U43349 ( .A(n30385), .B(n33739), .Z(n30389) );
  NOR U43350 ( .A(n30386), .B(n30389), .Z(n30387) );
  NOR U43351 ( .A(n37136), .B(n30387), .Z(n30388) );
  NOR U43352 ( .A(n30390), .B(n30388), .Z(n30393) );
  IV U43353 ( .A(n30389), .Z(n30392) );
  IV U43354 ( .A(n30390), .Z(n30391) );
  NOR U43355 ( .A(n30392), .B(n30391), .Z(n37139) );
  NOR U43356 ( .A(n30393), .B(n37139), .Z(n31725) );
  IV U43357 ( .A(n30394), .Z(n30395) );
  NOR U43358 ( .A(n30395), .B(n30401), .Z(n31724) );
  IV U43359 ( .A(n30396), .Z(n30397) );
  NOR U43360 ( .A(n30398), .B(n30397), .Z(n31727) );
  NOR U43361 ( .A(n31724), .B(n31727), .Z(n30399) );
  XOR U43362 ( .A(n31725), .B(n30399), .Z(n31723) );
  IV U43363 ( .A(n30400), .Z(n30402) );
  NOR U43364 ( .A(n30402), .B(n30401), .Z(n31721) );
  XOR U43365 ( .A(n31723), .B(n31721), .Z(n33743) );
  XOR U43366 ( .A(n31717), .B(n33743), .Z(n30403) );
  XOR U43367 ( .A(n30404), .B(n30403), .Z(n31715) );
  XOR U43368 ( .A(n30405), .B(n31715), .Z(n33749) );
  IV U43369 ( .A(n30406), .Z(n30409) );
  IV U43370 ( .A(n30407), .Z(n30408) );
  NOR U43371 ( .A(n30409), .B(n30408), .Z(n30416) );
  IV U43372 ( .A(n30416), .Z(n30410) );
  NOR U43373 ( .A(n33749), .B(n30410), .Z(n37160) );
  IV U43374 ( .A(n30411), .Z(n30414) );
  IV U43375 ( .A(n30412), .Z(n30413) );
  NOR U43376 ( .A(n30414), .B(n30413), .Z(n31711) );
  NOR U43377 ( .A(n33748), .B(n31711), .Z(n30415) );
  XOR U43378 ( .A(n30415), .B(n33749), .Z(n30426) );
  NOR U43379 ( .A(n30416), .B(n30426), .Z(n30417) );
  NOR U43380 ( .A(n37160), .B(n30417), .Z(n30420) );
  NOR U43381 ( .A(n30418), .B(n30420), .Z(n30432) );
  IV U43382 ( .A(n30419), .Z(n30424) );
  IV U43383 ( .A(n30420), .Z(n30421) );
  NOR U43384 ( .A(n30428), .B(n30421), .Z(n30422) );
  IV U43385 ( .A(n30422), .Z(n30423) );
  NOR U43386 ( .A(n30424), .B(n30423), .Z(n38487) );
  IV U43387 ( .A(n30425), .Z(n30431) );
  IV U43388 ( .A(n30426), .Z(n30427) );
  NOR U43389 ( .A(n30428), .B(n30427), .Z(n30429) );
  IV U43390 ( .A(n30429), .Z(n30430) );
  NOR U43391 ( .A(n30431), .B(n30430), .Z(n40422) );
  NOR U43392 ( .A(n38487), .B(n40422), .Z(n37159) );
  IV U43393 ( .A(n37159), .Z(n33753) );
  NOR U43394 ( .A(n30432), .B(n33753), .Z(n30442) );
  XOR U43395 ( .A(n30433), .B(n30442), .Z(n30440) );
  IV U43396 ( .A(n30440), .Z(n34989) );
  NOR U43397 ( .A(n30434), .B(n34989), .Z(n33756) );
  IV U43398 ( .A(n30435), .Z(n30436) );
  NOR U43399 ( .A(n30436), .B(n30438), .Z(n31700) );
  IV U43400 ( .A(n30437), .Z(n30439) );
  NOR U43401 ( .A(n30439), .B(n30438), .Z(n30441) );
  NOR U43402 ( .A(n30441), .B(n30440), .Z(n30444) );
  IV U43403 ( .A(n30441), .Z(n30443) );
  IV U43404 ( .A(n30442), .Z(n31704) );
  NOR U43405 ( .A(n30443), .B(n31704), .Z(n34996) );
  NOR U43406 ( .A(n30444), .B(n34996), .Z(n30445) );
  IV U43407 ( .A(n30445), .Z(n31701) );
  XOR U43408 ( .A(n31700), .B(n31701), .Z(n31693) );
  IV U43409 ( .A(n31693), .Z(n30446) );
  NOR U43410 ( .A(n30447), .B(n30446), .Z(n30448) );
  NOR U43411 ( .A(n33756), .B(n30448), .Z(n30449) );
  IV U43412 ( .A(n30449), .Z(n34982) );
  NOR U43413 ( .A(n30450), .B(n31694), .Z(n30461) );
  IV U43414 ( .A(n30451), .Z(n34985) );
  NOR U43415 ( .A(n30452), .B(n34985), .Z(n31690) );
  NOR U43416 ( .A(n30461), .B(n31690), .Z(n30453) );
  XOR U43417 ( .A(n34982), .B(n30453), .Z(n30464) );
  IV U43418 ( .A(n30464), .Z(n34974) );
  NOR U43419 ( .A(n30454), .B(n34974), .Z(n34975) );
  IV U43420 ( .A(n30455), .Z(n30456) );
  NOR U43421 ( .A(n30456), .B(n30459), .Z(n30457) );
  IV U43422 ( .A(n30457), .Z(n33759) );
  IV U43423 ( .A(n30458), .Z(n30460) );
  NOR U43424 ( .A(n30460), .B(n30459), .Z(n30465) );
  IV U43425 ( .A(n30465), .Z(n30463) );
  XOR U43426 ( .A(n30461), .B(n34982), .Z(n30462) );
  NOR U43427 ( .A(n30463), .B(n30462), .Z(n37188) );
  NOR U43428 ( .A(n30465), .B(n30464), .Z(n30466) );
  NOR U43429 ( .A(n37188), .B(n30466), .Z(n30467) );
  IV U43430 ( .A(n30467), .Z(n33758) );
  XOR U43431 ( .A(n33759), .B(n33758), .Z(n30468) );
  NOR U43432 ( .A(n30469), .B(n30468), .Z(n30470) );
  NOR U43433 ( .A(n34975), .B(n30470), .Z(n31686) );
  IV U43434 ( .A(n30471), .Z(n30473) );
  NOR U43435 ( .A(n30473), .B(n30472), .Z(n30474) );
  IV U43436 ( .A(n30474), .Z(n34971) );
  XOR U43437 ( .A(n31686), .B(n34971), .Z(n34964) );
  NOR U43438 ( .A(n33766), .B(n30475), .Z(n30479) );
  IV U43439 ( .A(n30476), .Z(n33768) );
  NOR U43440 ( .A(n30477), .B(n33768), .Z(n30478) );
  NOR U43441 ( .A(n30479), .B(n30478), .Z(n30480) );
  XOR U43442 ( .A(n34964), .B(n30480), .Z(n33772) );
  NOR U43443 ( .A(n33775), .B(n33773), .Z(n30484) );
  IV U43444 ( .A(n30481), .Z(n33782) );
  NOR U43445 ( .A(n30482), .B(n33782), .Z(n30483) );
  NOR U43446 ( .A(n30484), .B(n30483), .Z(n30485) );
  XOR U43447 ( .A(n33772), .B(n30485), .Z(n33788) );
  XOR U43448 ( .A(n33787), .B(n33788), .Z(n33791) );
  IV U43449 ( .A(n33791), .Z(n30487) );
  NOR U43450 ( .A(n33790), .B(n31677), .Z(n30486) );
  XOR U43451 ( .A(n30487), .B(n30486), .Z(n34933) );
  XOR U43452 ( .A(n31679), .B(n34933), .Z(n30501) );
  IV U43453 ( .A(n30488), .Z(n30489) );
  NOR U43454 ( .A(n30489), .B(n30494), .Z(n30490) );
  IV U43455 ( .A(n30490), .Z(n30504) );
  NOR U43456 ( .A(n30501), .B(n30504), .Z(n34929) );
  IV U43457 ( .A(n30513), .Z(n30511) );
  IV U43458 ( .A(n30491), .Z(n30514) );
  NOR U43459 ( .A(n30511), .B(n30514), .Z(n30492) );
  IV U43460 ( .A(n30492), .Z(n33797) );
  IV U43461 ( .A(n30493), .Z(n30495) );
  NOR U43462 ( .A(n30495), .B(n30494), .Z(n30500) );
  IV U43463 ( .A(n30496), .Z(n34937) );
  NOR U43464 ( .A(n30497), .B(n34937), .Z(n31675) );
  NOR U43465 ( .A(n31679), .B(n31675), .Z(n30498) );
  XOR U43466 ( .A(n34933), .B(n30498), .Z(n30499) );
  NOR U43467 ( .A(n30500), .B(n30499), .Z(n30503) );
  IV U43468 ( .A(n30500), .Z(n30502) );
  NOR U43469 ( .A(n30502), .B(n30501), .Z(n34926) );
  NOR U43470 ( .A(n30503), .B(n34926), .Z(n30505) );
  IV U43471 ( .A(n30505), .Z(n33796) );
  XOR U43472 ( .A(n33797), .B(n33796), .Z(n30507) );
  NOR U43473 ( .A(n30505), .B(n30504), .Z(n30506) );
  NOR U43474 ( .A(n30507), .B(n30506), .Z(n30508) );
  NOR U43475 ( .A(n34929), .B(n30508), .Z(n31669) );
  IV U43476 ( .A(n30509), .Z(n30510) );
  NOR U43477 ( .A(n30511), .B(n30510), .Z(n33798) );
  IV U43478 ( .A(n30512), .Z(n30516) );
  XOR U43479 ( .A(n30514), .B(n30513), .Z(n30515) );
  NOR U43480 ( .A(n30516), .B(n30515), .Z(n31670) );
  NOR U43481 ( .A(n33798), .B(n31670), .Z(n30517) );
  XOR U43482 ( .A(n31669), .B(n30517), .Z(n31674) );
  XOR U43483 ( .A(n30518), .B(n31674), .Z(n30519) );
  IV U43484 ( .A(n30519), .Z(n34912) );
  IV U43485 ( .A(n30520), .Z(n30521) );
  NOR U43486 ( .A(n30521), .B(n30523), .Z(n33806) );
  IV U43487 ( .A(n30522), .Z(n30524) );
  NOR U43488 ( .A(n30524), .B(n30523), .Z(n34911) );
  IV U43489 ( .A(n30525), .Z(n30526) );
  NOR U43490 ( .A(n30527), .B(n30526), .Z(n34916) );
  NOR U43491 ( .A(n34911), .B(n34916), .Z(n33803) );
  IV U43492 ( .A(n33803), .Z(n30528) );
  NOR U43493 ( .A(n33806), .B(n30528), .Z(n30529) );
  XOR U43494 ( .A(n34912), .B(n30529), .Z(n30535) );
  IV U43495 ( .A(n30535), .Z(n30534) );
  IV U43496 ( .A(n30530), .Z(n30532) );
  NOR U43497 ( .A(n30532), .B(n30531), .Z(n30536) );
  IV U43498 ( .A(n30536), .Z(n30533) );
  NOR U43499 ( .A(n30534), .B(n30533), .Z(n34908) );
  NOR U43500 ( .A(n30536), .B(n30535), .Z(n33816) );
  IV U43501 ( .A(n30537), .Z(n30538) );
  NOR U43502 ( .A(n30542), .B(n30538), .Z(n33814) );
  XOR U43503 ( .A(n33816), .B(n33814), .Z(n30539) );
  NOR U43504 ( .A(n34908), .B(n30539), .Z(n33809) );
  IV U43505 ( .A(n30540), .Z(n30541) );
  NOR U43506 ( .A(n30542), .B(n30541), .Z(n30543) );
  IV U43507 ( .A(n30543), .Z(n33812) );
  XOR U43508 ( .A(n33809), .B(n33812), .Z(n31665) );
  IV U43509 ( .A(n31665), .Z(n30551) );
  IV U43510 ( .A(n30544), .Z(n30554) );
  IV U43511 ( .A(n30545), .Z(n30546) );
  NOR U43512 ( .A(n30554), .B(n30546), .Z(n31663) );
  IV U43513 ( .A(n30547), .Z(n30549) );
  NOR U43514 ( .A(n30549), .B(n30548), .Z(n33810) );
  NOR U43515 ( .A(n31663), .B(n33810), .Z(n30550) );
  XOR U43516 ( .A(n30551), .B(n30550), .Z(n31662) );
  IV U43517 ( .A(n30552), .Z(n30553) );
  NOR U43518 ( .A(n30554), .B(n30553), .Z(n31660) );
  XOR U43519 ( .A(n31662), .B(n31660), .Z(n33824) );
  XOR U43520 ( .A(n31659), .B(n33824), .Z(n30555) );
  IV U43521 ( .A(n30555), .Z(n31655) );
  XOR U43522 ( .A(n31654), .B(n31655), .Z(n33840) );
  IV U43523 ( .A(n30556), .Z(n30557) );
  NOR U43524 ( .A(n30560), .B(n30557), .Z(n31657) );
  IV U43525 ( .A(n30558), .Z(n30559) );
  NOR U43526 ( .A(n30560), .B(n30559), .Z(n33838) );
  NOR U43527 ( .A(n31657), .B(n33838), .Z(n30561) );
  XOR U43528 ( .A(n33840), .B(n30561), .Z(n31651) );
  IV U43529 ( .A(n30562), .Z(n30573) );
  IV U43530 ( .A(n30563), .Z(n30564) );
  NOR U43531 ( .A(n30573), .B(n30564), .Z(n31652) );
  IV U43532 ( .A(n30565), .Z(n30567) );
  NOR U43533 ( .A(n30567), .B(n30566), .Z(n33835) );
  NOR U43534 ( .A(n31652), .B(n33835), .Z(n30568) );
  XOR U43535 ( .A(n31651), .B(n30568), .Z(n33846) );
  IV U43536 ( .A(n30569), .Z(n30570) );
  NOR U43537 ( .A(n30570), .B(n30576), .Z(n33845) );
  IV U43538 ( .A(n30571), .Z(n30572) );
  NOR U43539 ( .A(n30573), .B(n30572), .Z(n33841) );
  NOR U43540 ( .A(n33845), .B(n33841), .Z(n30574) );
  XOR U43541 ( .A(n33846), .B(n30574), .Z(n31644) );
  IV U43542 ( .A(n30575), .Z(n30577) );
  NOR U43543 ( .A(n30577), .B(n30576), .Z(n30578) );
  IV U43544 ( .A(n30578), .Z(n33843) );
  XOR U43545 ( .A(n31644), .B(n33843), .Z(n34876) );
  XOR U43546 ( .A(n37245), .B(n34876), .Z(n31638) );
  XOR U43547 ( .A(n30579), .B(n31638), .Z(n33849) );
  XOR U43548 ( .A(n33850), .B(n33849), .Z(n31633) );
  XOR U43549 ( .A(n31632), .B(n31633), .Z(n31625) );
  XOR U43550 ( .A(n30580), .B(n31625), .Z(n31616) );
  XOR U43551 ( .A(n30581), .B(n31616), .Z(n33863) );
  XOR U43552 ( .A(n33862), .B(n33863), .Z(n33866) );
  XOR U43553 ( .A(n33865), .B(n33866), .Z(n33869) );
  XOR U43554 ( .A(n33870), .B(n33869), .Z(n30589) );
  IV U43555 ( .A(n30589), .Z(n34856) );
  NOR U43556 ( .A(n30582), .B(n34856), .Z(n37277) );
  IV U43557 ( .A(n30583), .Z(n30584) );
  NOR U43558 ( .A(n30584), .B(n30586), .Z(n31613) );
  IV U43559 ( .A(n30585), .Z(n30587) );
  NOR U43560 ( .A(n30587), .B(n30586), .Z(n30590) );
  IV U43561 ( .A(n30590), .Z(n30588) );
  NOR U43562 ( .A(n30588), .B(n33869), .Z(n37270) );
  NOR U43563 ( .A(n30590), .B(n30589), .Z(n30591) );
  NOR U43564 ( .A(n37270), .B(n30591), .Z(n30592) );
  IV U43565 ( .A(n30592), .Z(n31614) );
  XOR U43566 ( .A(n31613), .B(n31614), .Z(n30598) );
  IV U43567 ( .A(n30598), .Z(n30593) );
  NOR U43568 ( .A(n30594), .B(n30593), .Z(n30595) );
  NOR U43569 ( .A(n37277), .B(n30595), .Z(n30596) );
  NOR U43570 ( .A(n30597), .B(n30596), .Z(n30600) );
  IV U43571 ( .A(n30597), .Z(n30599) );
  NOR U43572 ( .A(n30599), .B(n30598), .Z(n37274) );
  NOR U43573 ( .A(n30600), .B(n37274), .Z(n30601) );
  IV U43574 ( .A(n30601), .Z(n33873) );
  XOR U43575 ( .A(n33872), .B(n33873), .Z(n33879) );
  IV U43576 ( .A(n30602), .Z(n30604) );
  NOR U43577 ( .A(n30604), .B(n30603), .Z(n33875) );
  XOR U43578 ( .A(n33879), .B(n33875), .Z(n31611) );
  IV U43579 ( .A(n30605), .Z(n33880) );
  NOR U43580 ( .A(n33880), .B(n33882), .Z(n30608) );
  IV U43581 ( .A(n30606), .Z(n30607) );
  NOR U43582 ( .A(n30607), .B(n30611), .Z(n31610) );
  NOR U43583 ( .A(n30608), .B(n31610), .Z(n30613) );
  XOR U43584 ( .A(n31611), .B(n30613), .Z(n30618) );
  IV U43585 ( .A(n30618), .Z(n30609) );
  IV U43586 ( .A(n30621), .Z(n34835) );
  NOR U43587 ( .A(n30609), .B(n34835), .Z(n33891) );
  IV U43588 ( .A(n30610), .Z(n30612) );
  NOR U43589 ( .A(n30612), .B(n30611), .Z(n30619) );
  IV U43590 ( .A(n30619), .Z(n30617) );
  IV U43591 ( .A(n30613), .Z(n30614) );
  NOR U43592 ( .A(n31611), .B(n30614), .Z(n30615) );
  IV U43593 ( .A(n30615), .Z(n30616) );
  NOR U43594 ( .A(n30617), .B(n30616), .Z(n34832) );
  NOR U43595 ( .A(n30619), .B(n30618), .Z(n30620) );
  NOR U43596 ( .A(n34832), .B(n30620), .Z(n31609) );
  NOR U43597 ( .A(n30621), .B(n31609), .Z(n30622) );
  NOR U43598 ( .A(n33891), .B(n30622), .Z(n33886) );
  NOR U43599 ( .A(n30624), .B(n30623), .Z(n33888) );
  IV U43600 ( .A(n30625), .Z(n41626) );
  NOR U43601 ( .A(n30626), .B(n41626), .Z(n31608) );
  NOR U43602 ( .A(n33888), .B(n31608), .Z(n30627) );
  XOR U43603 ( .A(n33886), .B(n30627), .Z(n34821) );
  XOR U43604 ( .A(n33898), .B(n34821), .Z(n31604) );
  XOR U43605 ( .A(n30628), .B(n31604), .Z(n31592) );
  IV U43606 ( .A(n30629), .Z(n31596) );
  NOR U43607 ( .A(n30630), .B(n31596), .Z(n30634) );
  IV U43608 ( .A(n30631), .Z(n30633) );
  NOR U43609 ( .A(n30633), .B(n30632), .Z(n31593) );
  NOR U43610 ( .A(n30634), .B(n31593), .Z(n30635) );
  XOR U43611 ( .A(n31592), .B(n30635), .Z(n31585) );
  XOR U43612 ( .A(n31584), .B(n31585), .Z(n33907) );
  XOR U43613 ( .A(n31580), .B(n33907), .Z(n33915) );
  XOR U43614 ( .A(n30636), .B(n33915), .Z(n30637) );
  IV U43615 ( .A(n30637), .Z(n33921) );
  XOR U43616 ( .A(n33919), .B(n33921), .Z(n33923) );
  IV U43617 ( .A(n33923), .Z(n30644) );
  IV U43618 ( .A(n30638), .Z(n30639) );
  NOR U43619 ( .A(n30642), .B(n30639), .Z(n33922) );
  IV U43620 ( .A(n30640), .Z(n30641) );
  NOR U43621 ( .A(n30642), .B(n30641), .Z(n33917) );
  NOR U43622 ( .A(n33922), .B(n33917), .Z(n30643) );
  XOR U43623 ( .A(n30644), .B(n30643), .Z(n33930) );
  IV U43624 ( .A(n30645), .Z(n30647) );
  NOR U43625 ( .A(n30647), .B(n30646), .Z(n33927) );
  XOR U43626 ( .A(n33930), .B(n33927), .Z(n33943) );
  XOR U43627 ( .A(n30648), .B(n33943), .Z(n33941) );
  XOR U43628 ( .A(n34792), .B(n33941), .Z(n33948) );
  XOR U43629 ( .A(n33947), .B(n33948), .Z(n33954) );
  XOR U43630 ( .A(n33950), .B(n33954), .Z(n30649) );
  NOR U43631 ( .A(n30650), .B(n30649), .Z(n37355) );
  IV U43632 ( .A(n30651), .Z(n30652) );
  NOR U43633 ( .A(n30653), .B(n30652), .Z(n33953) );
  NOR U43634 ( .A(n33953), .B(n33950), .Z(n30654) );
  XOR U43635 ( .A(n30654), .B(n33954), .Z(n30662) );
  NOR U43636 ( .A(n30655), .B(n30662), .Z(n30656) );
  NOR U43637 ( .A(n37355), .B(n30656), .Z(n30665) );
  IV U43638 ( .A(n30665), .Z(n30657) );
  NOR U43639 ( .A(n30658), .B(n30657), .Z(n34779) );
  IV U43640 ( .A(n30659), .Z(n30661) );
  NOR U43641 ( .A(n30661), .B(n30660), .Z(n30666) );
  IV U43642 ( .A(n30666), .Z(n30664) );
  IV U43643 ( .A(n30662), .Z(n30663) );
  NOR U43644 ( .A(n30664), .B(n30663), .Z(n34781) );
  NOR U43645 ( .A(n30666), .B(n30665), .Z(n30667) );
  NOR U43646 ( .A(n34781), .B(n30667), .Z(n30671) );
  NOR U43647 ( .A(n30668), .B(n30671), .Z(n30669) );
  NOR U43648 ( .A(n34779), .B(n30669), .Z(n33959) );
  NOR U43649 ( .A(n30670), .B(n33959), .Z(n30674) );
  IV U43650 ( .A(n30670), .Z(n30673) );
  IV U43651 ( .A(n30671), .Z(n30672) );
  NOR U43652 ( .A(n30673), .B(n30672), .Z(n37358) );
  NOR U43653 ( .A(n30674), .B(n37358), .Z(n33966) );
  IV U43654 ( .A(n30675), .Z(n30677) );
  NOR U43655 ( .A(n30677), .B(n30676), .Z(n33960) );
  IV U43656 ( .A(n30678), .Z(n30679) );
  NOR U43657 ( .A(n30683), .B(n30679), .Z(n33967) );
  NOR U43658 ( .A(n33960), .B(n33967), .Z(n30680) );
  XOR U43659 ( .A(n33966), .B(n30680), .Z(n31579) );
  IV U43660 ( .A(n30681), .Z(n30682) );
  NOR U43661 ( .A(n30683), .B(n30682), .Z(n31577) );
  XOR U43662 ( .A(n31579), .B(n31577), .Z(n31569) );
  XOR U43663 ( .A(n30684), .B(n31569), .Z(n31570) );
  XOR U43664 ( .A(n30685), .B(n31570), .Z(n34757) );
  XOR U43665 ( .A(n30686), .B(n34757), .Z(n33978) );
  XOR U43666 ( .A(n30687), .B(n33978), .Z(n37385) );
  XOR U43667 ( .A(n33989), .B(n37385), .Z(n33996) );
  XOR U43668 ( .A(n30688), .B(n33996), .Z(n31559) );
  XOR U43669 ( .A(n31557), .B(n31559), .Z(n31556) );
  XOR U43670 ( .A(n30689), .B(n31556), .Z(n30690) );
  IV U43671 ( .A(n30690), .Z(n31547) );
  XOR U43672 ( .A(n31546), .B(n31547), .Z(n31536) );
  IV U43673 ( .A(n30691), .Z(n31537) );
  NOR U43674 ( .A(n30692), .B(n31537), .Z(n30696) );
  IV U43675 ( .A(n30693), .Z(n30695) );
  NOR U43676 ( .A(n30695), .B(n30694), .Z(n31543) );
  NOR U43677 ( .A(n30696), .B(n31543), .Z(n30697) );
  XOR U43678 ( .A(n31536), .B(n30697), .Z(n31529) );
  IV U43679 ( .A(n30698), .Z(n30700) );
  NOR U43680 ( .A(n30700), .B(n30699), .Z(n30705) );
  IV U43681 ( .A(n30705), .Z(n30701) );
  NOR U43682 ( .A(n31529), .B(n30701), .Z(n34731) );
  NOR U43683 ( .A(n30702), .B(n31528), .Z(n30703) );
  XOR U43684 ( .A(n30703), .B(n31529), .Z(n31524) );
  IV U43685 ( .A(n31524), .Z(n30704) );
  NOR U43686 ( .A(n30705), .B(n30704), .Z(n30706) );
  NOR U43687 ( .A(n34731), .B(n30706), .Z(n30707) );
  IV U43688 ( .A(n30707), .Z(n34001) );
  XOR U43689 ( .A(n34000), .B(n34001), .Z(n31512) );
  IV U43690 ( .A(n31523), .Z(n30709) );
  NOR U43691 ( .A(n30709), .B(n30708), .Z(n30712) );
  NOR U43692 ( .A(n31513), .B(n30710), .Z(n30711) );
  NOR U43693 ( .A(n30712), .B(n30711), .Z(n30713) );
  XOR U43694 ( .A(n31512), .B(n30713), .Z(n31506) );
  NOR U43695 ( .A(n31507), .B(n30714), .Z(n30718) );
  IV U43696 ( .A(n30715), .Z(n31502) );
  NOR U43697 ( .A(n30716), .B(n31502), .Z(n30717) );
  NOR U43698 ( .A(n30718), .B(n30717), .Z(n30719) );
  XOR U43699 ( .A(n31506), .B(n30719), .Z(n31491) );
  XOR U43700 ( .A(n31498), .B(n31491), .Z(n31488) );
  XOR U43701 ( .A(n30720), .B(n31488), .Z(n30721) );
  IV U43702 ( .A(n30721), .Z(n31483) );
  XOR U43703 ( .A(n31481), .B(n31483), .Z(n37460) );
  IV U43704 ( .A(n37460), .Z(n30727) );
  NOR U43705 ( .A(n31478), .B(n30722), .Z(n30725) );
  IV U43706 ( .A(n30723), .Z(n37464) );
  NOR U43707 ( .A(n30724), .B(n37464), .Z(n31466) );
  NOR U43708 ( .A(n30725), .B(n31466), .Z(n30726) );
  XOR U43709 ( .A(n30727), .B(n30726), .Z(n31470) );
  XOR U43710 ( .A(n31468), .B(n31470), .Z(n31473) );
  XOR U43711 ( .A(n31471), .B(n31473), .Z(n31461) );
  XOR U43712 ( .A(n31460), .B(n31461), .Z(n31454) );
  NOR U43713 ( .A(n30728), .B(n31454), .Z(n37480) );
  IV U43714 ( .A(n30729), .Z(n31457) );
  NOR U43715 ( .A(n31457), .B(n30730), .Z(n30734) );
  IV U43716 ( .A(n30731), .Z(n30733) );
  NOR U43717 ( .A(n30733), .B(n30732), .Z(n31453) );
  NOR U43718 ( .A(n30734), .B(n31453), .Z(n30735) );
  XOR U43719 ( .A(n30735), .B(n31454), .Z(n30741) );
  NOR U43720 ( .A(n30736), .B(n30741), .Z(n30737) );
  NOR U43721 ( .A(n37480), .B(n30737), .Z(n30738) );
  IV U43722 ( .A(n30738), .Z(n34026) );
  IV U43723 ( .A(n30739), .Z(n34027) );
  XOR U43724 ( .A(n34026), .B(n34027), .Z(n30740) );
  NOR U43725 ( .A(n30742), .B(n30740), .Z(n30745) );
  IV U43726 ( .A(n30741), .Z(n30744) );
  IV U43727 ( .A(n30742), .Z(n30743) );
  NOR U43728 ( .A(n30744), .B(n30743), .Z(n37486) );
  NOR U43729 ( .A(n30745), .B(n37486), .Z(n30753) );
  IV U43730 ( .A(n30753), .Z(n37500) );
  NOR U43731 ( .A(n30746), .B(n37500), .Z(n37489) );
  NOR U43732 ( .A(n30757), .B(n37489), .Z(n31451) );
  IV U43733 ( .A(n31451), .Z(n30756) );
  IV U43734 ( .A(n30747), .Z(n30750) );
  IV U43735 ( .A(n30748), .Z(n30749) );
  NOR U43736 ( .A(n30750), .B(n30749), .Z(n30752) );
  IV U43737 ( .A(n30752), .Z(n30751) );
  NOR U43738 ( .A(n34026), .B(n30751), .Z(n34706) );
  NOR U43739 ( .A(n30753), .B(n30752), .Z(n30754) );
  NOR U43740 ( .A(n34706), .B(n30754), .Z(n30758) );
  NOR U43741 ( .A(n30755), .B(n30758), .Z(n31452) );
  NOR U43742 ( .A(n30756), .B(n31452), .Z(n30760) );
  IV U43743 ( .A(n30757), .Z(n37497) );
  NOR U43744 ( .A(n30758), .B(n37497), .Z(n30759) );
  NOR U43745 ( .A(n30760), .B(n30759), .Z(n31447) );
  IV U43746 ( .A(n30761), .Z(n30763) );
  NOR U43747 ( .A(n30763), .B(n30762), .Z(n31445) );
  XOR U43748 ( .A(n31447), .B(n31445), .Z(n31450) );
  XOR U43749 ( .A(n31448), .B(n31450), .Z(n34035) );
  XOR U43750 ( .A(n30764), .B(n34035), .Z(n34687) );
  XOR U43751 ( .A(n30765), .B(n34687), .Z(n47688) );
  XOR U43752 ( .A(n31435), .B(n47688), .Z(n34045) );
  XOR U43753 ( .A(n34690), .B(n34045), .Z(n30773) );
  IV U43754 ( .A(n30773), .Z(n34682) );
  IV U43755 ( .A(n30766), .Z(n30787) );
  IV U43756 ( .A(n30767), .Z(n30768) );
  NOR U43757 ( .A(n30787), .B(n30768), .Z(n30782) );
  IV U43758 ( .A(n30782), .Z(n30769) );
  NOR U43759 ( .A(n34682), .B(n30769), .Z(n34678) );
  IV U43760 ( .A(n30770), .Z(n30771) );
  NOR U43761 ( .A(n30771), .B(n30778), .Z(n30774) );
  IV U43762 ( .A(n30774), .Z(n30772) );
  NOR U43763 ( .A(n47688), .B(n30772), .Z(n37517) );
  NOR U43764 ( .A(n30774), .B(n30773), .Z(n30775) );
  NOR U43765 ( .A(n37517), .B(n30775), .Z(n30776) );
  IV U43766 ( .A(n30776), .Z(n44194) );
  IV U43767 ( .A(n30777), .Z(n30779) );
  NOR U43768 ( .A(n30779), .B(n30778), .Z(n30780) );
  IV U43769 ( .A(n30780), .Z(n44188) );
  XOR U43770 ( .A(n44194), .B(n44188), .Z(n30781) );
  NOR U43771 ( .A(n30782), .B(n30781), .Z(n30783) );
  NOR U43772 ( .A(n34678), .B(n30783), .Z(n30784) );
  IV U43773 ( .A(n30784), .Z(n31431) );
  IV U43774 ( .A(n30785), .Z(n30786) );
  NOR U43775 ( .A(n30787), .B(n30786), .Z(n31430) );
  XOR U43776 ( .A(n31431), .B(n31430), .Z(n31432) );
  XOR U43777 ( .A(n31433), .B(n31432), .Z(n30792) );
  IV U43778 ( .A(n30792), .Z(n37524) );
  NOR U43779 ( .A(n30788), .B(n37524), .Z(n37534) );
  NOR U43780 ( .A(n30790), .B(n30789), .Z(n30793) );
  IV U43781 ( .A(n30793), .Z(n30791) );
  NOR U43782 ( .A(n30791), .B(n31432), .Z(n31423) );
  NOR U43783 ( .A(n30793), .B(n30792), .Z(n30794) );
  NOR U43784 ( .A(n31423), .B(n30794), .Z(n30795) );
  NOR U43785 ( .A(n30796), .B(n30795), .Z(n30797) );
  NOR U43786 ( .A(n37534), .B(n30797), .Z(n34054) );
  IV U43787 ( .A(n30798), .Z(n30800) );
  NOR U43788 ( .A(n30800), .B(n30799), .Z(n30801) );
  IV U43789 ( .A(n30801), .Z(n34055) );
  XOR U43790 ( .A(n34054), .B(n34055), .Z(n37542) );
  XOR U43791 ( .A(n34059), .B(n37542), .Z(n34061) );
  XOR U43792 ( .A(n30802), .B(n34061), .Z(n34073) );
  XOR U43793 ( .A(n34071), .B(n34073), .Z(n34075) );
  XOR U43794 ( .A(n34074), .B(n34075), .Z(n34080) );
  IV U43795 ( .A(n30803), .Z(n30804) );
  NOR U43796 ( .A(n30805), .B(n30804), .Z(n34078) );
  XOR U43797 ( .A(n34080), .B(n34078), .Z(n34083) );
  IV U43798 ( .A(n30806), .Z(n30816) );
  IV U43799 ( .A(n30807), .Z(n30808) );
  NOR U43800 ( .A(n30816), .B(n30808), .Z(n31421) );
  IV U43801 ( .A(n30809), .Z(n30811) );
  NOR U43802 ( .A(n30811), .B(n30810), .Z(n34081) );
  NOR U43803 ( .A(n31421), .B(n34081), .Z(n30812) );
  XOR U43804 ( .A(n34083), .B(n30812), .Z(n30813) );
  IV U43805 ( .A(n30813), .Z(n31420) );
  IV U43806 ( .A(n30814), .Z(n30815) );
  NOR U43807 ( .A(n30816), .B(n30815), .Z(n30817) );
  IV U43808 ( .A(n30817), .Z(n31419) );
  XOR U43809 ( .A(n31420), .B(n31419), .Z(n30826) );
  IV U43810 ( .A(n30826), .Z(n41471) );
  IV U43811 ( .A(n30818), .Z(n30839) );
  IV U43812 ( .A(n30819), .Z(n30820) );
  NOR U43813 ( .A(n30839), .B(n30820), .Z(n30834) );
  IV U43814 ( .A(n30834), .Z(n30821) );
  NOR U43815 ( .A(n41471), .B(n30821), .Z(n34643) );
  IV U43816 ( .A(n30822), .Z(n30823) );
  NOR U43817 ( .A(n30823), .B(n30830), .Z(n30825) );
  IV U43818 ( .A(n30825), .Z(n30824) );
  NOR U43819 ( .A(n31420), .B(n30824), .Z(n34649) );
  NOR U43820 ( .A(n30826), .B(n30825), .Z(n30827) );
  NOR U43821 ( .A(n34649), .B(n30827), .Z(n30828) );
  IV U43822 ( .A(n30828), .Z(n31418) );
  IV U43823 ( .A(n30829), .Z(n30831) );
  NOR U43824 ( .A(n30831), .B(n30830), .Z(n30832) );
  IV U43825 ( .A(n30832), .Z(n31417) );
  XOR U43826 ( .A(n31418), .B(n31417), .Z(n30833) );
  NOR U43827 ( .A(n30834), .B(n30833), .Z(n30835) );
  NOR U43828 ( .A(n34643), .B(n30835), .Z(n30836) );
  IV U43829 ( .A(n30836), .Z(n34087) );
  IV U43830 ( .A(n30837), .Z(n30838) );
  NOR U43831 ( .A(n30839), .B(n30838), .Z(n30844) );
  IV U43832 ( .A(n30844), .Z(n41483) );
  XOR U43833 ( .A(n34087), .B(n41483), .Z(n30846) );
  IV U43834 ( .A(n30840), .Z(n30842) );
  NOR U43835 ( .A(n30842), .B(n30841), .Z(n30843) );
  IV U43836 ( .A(n30843), .Z(n30850) );
  NOR U43837 ( .A(n30844), .B(n30850), .Z(n30845) );
  NOR U43838 ( .A(n30846), .B(n30845), .Z(n30855) );
  IV U43839 ( .A(n30855), .Z(n30847) );
  NOR U43840 ( .A(n30848), .B(n30847), .Z(n30851) );
  IV U43841 ( .A(n30848), .Z(n30849) );
  NOR U43842 ( .A(n30849), .B(n34087), .Z(n38191) );
  NOR U43843 ( .A(n30850), .B(n34087), .Z(n38198) );
  NOR U43844 ( .A(n38191), .B(n38198), .Z(n34640) );
  IV U43845 ( .A(n34640), .Z(n34090) );
  NOR U43846 ( .A(n30851), .B(n34090), .Z(n31409) );
  IV U43847 ( .A(n30852), .Z(n31411) );
  NOR U43848 ( .A(n30853), .B(n31411), .Z(n30861) );
  IV U43849 ( .A(n30861), .Z(n30854) );
  NOR U43850 ( .A(n31409), .B(n30854), .Z(n30863) );
  IV U43851 ( .A(n30857), .Z(n30856) );
  NOR U43852 ( .A(n30856), .B(n30855), .Z(n34632) );
  NOR U43853 ( .A(n31409), .B(n30857), .Z(n30858) );
  NOR U43854 ( .A(n34632), .B(n30858), .Z(n30859) );
  IV U43855 ( .A(n30859), .Z(n30860) );
  NOR U43856 ( .A(n30861), .B(n30860), .Z(n30862) );
  NOR U43857 ( .A(n30863), .B(n30862), .Z(n31407) );
  NOR U43858 ( .A(n30864), .B(n31407), .Z(n34624) );
  IV U43859 ( .A(n30865), .Z(n30866) );
  NOR U43860 ( .A(n30866), .B(n30869), .Z(n30867) );
  IV U43861 ( .A(n30867), .Z(n31403) );
  IV U43862 ( .A(n30868), .Z(n30870) );
  NOR U43863 ( .A(n30870), .B(n30869), .Z(n31405) );
  XOR U43864 ( .A(n31407), .B(n31405), .Z(n31402) );
  XOR U43865 ( .A(n31403), .B(n31402), .Z(n30871) );
  NOR U43866 ( .A(n30872), .B(n30871), .Z(n30873) );
  NOR U43867 ( .A(n34624), .B(n30873), .Z(n30874) );
  IV U43868 ( .A(n30874), .Z(n31400) );
  XOR U43869 ( .A(n31395), .B(n31400), .Z(n31390) );
  NOR U43870 ( .A(n30875), .B(n31385), .Z(n30878) );
  NOR U43871 ( .A(n30876), .B(n31391), .Z(n30877) );
  NOR U43872 ( .A(n30878), .B(n30877), .Z(n30879) );
  XOR U43873 ( .A(n31390), .B(n30879), .Z(n31382) );
  IV U43874 ( .A(n31382), .Z(n30890) );
  IV U43875 ( .A(n30880), .Z(n31376) );
  NOR U43876 ( .A(n30881), .B(n31376), .Z(n30888) );
  IV U43877 ( .A(n30882), .Z(n30883) );
  NOR U43878 ( .A(n30886), .B(n30883), .Z(n30898) );
  IV U43879 ( .A(n30898), .Z(n31383) );
  IV U43880 ( .A(n30884), .Z(n30885) );
  NOR U43881 ( .A(n30886), .B(n30885), .Z(n30899) );
  IV U43882 ( .A(n30899), .Z(n34096) );
  XOR U43883 ( .A(n31383), .B(n34096), .Z(n30887) );
  NOR U43884 ( .A(n30888), .B(n30887), .Z(n30889) );
  XOR U43885 ( .A(n30890), .B(n30889), .Z(n30908) );
  IV U43886 ( .A(n30891), .Z(n30893) );
  NOR U43887 ( .A(n30893), .B(n30892), .Z(n30911) );
  IV U43888 ( .A(n30911), .Z(n30894) );
  NOR U43889 ( .A(n30908), .B(n30894), .Z(n34604) );
  IV U43890 ( .A(n30895), .Z(n30896) );
  NOR U43891 ( .A(n31367), .B(n30896), .Z(n30914) );
  NOR U43892 ( .A(n34604), .B(n30914), .Z(n30897) );
  IV U43893 ( .A(n30897), .Z(n30913) );
  XOR U43894 ( .A(n30898), .B(n31382), .Z(n34095) );
  XOR U43895 ( .A(n30899), .B(n34095), .Z(n31373) );
  IV U43896 ( .A(n31373), .Z(n30905) );
  IV U43897 ( .A(n30900), .Z(n30901) );
  NOR U43898 ( .A(n30901), .B(n30903), .Z(n31372) );
  IV U43899 ( .A(n30902), .Z(n30904) );
  NOR U43900 ( .A(n30904), .B(n30903), .Z(n31370) );
  NOR U43901 ( .A(n31372), .B(n31370), .Z(n30906) );
  NOR U43902 ( .A(n30905), .B(n30906), .Z(n30910) );
  IV U43903 ( .A(n30906), .Z(n30907) );
  NOR U43904 ( .A(n30908), .B(n30907), .Z(n30909) );
  NOR U43905 ( .A(n30910), .B(n30909), .Z(n34599) );
  IV U43906 ( .A(n34599), .Z(n30915) );
  NOR U43907 ( .A(n30911), .B(n30915), .Z(n30912) );
  NOR U43908 ( .A(n30913), .B(n30912), .Z(n30917) );
  IV U43909 ( .A(n30914), .Z(n37570) );
  NOR U43910 ( .A(n30915), .B(n37570), .Z(n30916) );
  NOR U43911 ( .A(n30917), .B(n30916), .Z(n30918) );
  XOR U43912 ( .A(n34598), .B(n30918), .Z(n34113) );
  IV U43913 ( .A(n30919), .Z(n30920) );
  NOR U43914 ( .A(n30920), .B(n30922), .Z(n31364) );
  IV U43915 ( .A(n30921), .Z(n30923) );
  NOR U43916 ( .A(n30923), .B(n30922), .Z(n34111) );
  NOR U43917 ( .A(n31364), .B(n34111), .Z(n30924) );
  XOR U43918 ( .A(n34113), .B(n30924), .Z(n34109) );
  IV U43919 ( .A(n30925), .Z(n30926) );
  NOR U43920 ( .A(n30927), .B(n30926), .Z(n34591) );
  IV U43921 ( .A(n30928), .Z(n30930) );
  NOR U43922 ( .A(n30930), .B(n30929), .Z(n34595) );
  NOR U43923 ( .A(n34591), .B(n34595), .Z(n34110) );
  XOR U43924 ( .A(n34109), .B(n34110), .Z(n34584) );
  XOR U43925 ( .A(n34116), .B(n34584), .Z(n34117) );
  IV U43926 ( .A(n30931), .Z(n30933) );
  NOR U43927 ( .A(n30933), .B(n30932), .Z(n30934) );
  IV U43928 ( .A(n30934), .Z(n34579) );
  XOR U43929 ( .A(n34117), .B(n34579), .Z(n34122) );
  XOR U43930 ( .A(n34121), .B(n34122), .Z(n34125) );
  XOR U43931 ( .A(n34124), .B(n34125), .Z(n31362) );
  IV U43932 ( .A(n30935), .Z(n30936) );
  NOR U43933 ( .A(n30937), .B(n30936), .Z(n31360) );
  XOR U43934 ( .A(n31362), .B(n31360), .Z(n31354) );
  IV U43935 ( .A(n31354), .Z(n30948) );
  IV U43936 ( .A(n30938), .Z(n30940) );
  IV U43937 ( .A(n30939), .Z(n30942) );
  NOR U43938 ( .A(n30940), .B(n30942), .Z(n31351) );
  NOR U43939 ( .A(n30941), .B(n31357), .Z(n30944) );
  NOR U43940 ( .A(n30943), .B(n30942), .Z(n31353) );
  NOR U43941 ( .A(n30944), .B(n31353), .Z(n30945) );
  IV U43942 ( .A(n30945), .Z(n30946) );
  NOR U43943 ( .A(n31351), .B(n30946), .Z(n30947) );
  XOR U43944 ( .A(n30948), .B(n30947), .Z(n31347) );
  IV U43945 ( .A(n30949), .Z(n30951) );
  NOR U43946 ( .A(n30951), .B(n30950), .Z(n31345) );
  XOR U43947 ( .A(n31347), .B(n31345), .Z(n34136) );
  XOR U43948 ( .A(n30952), .B(n34136), .Z(n30962) );
  IV U43949 ( .A(n30962), .Z(n30957) );
  IV U43950 ( .A(n30953), .Z(n30954) );
  NOR U43951 ( .A(n30955), .B(n30954), .Z(n30965) );
  IV U43952 ( .A(n30965), .Z(n30956) );
  NOR U43953 ( .A(n30957), .B(n30956), .Z(n34552) );
  IV U43954 ( .A(n30958), .Z(n30960) );
  NOR U43955 ( .A(n30960), .B(n30959), .Z(n30963) );
  IV U43956 ( .A(n30963), .Z(n30961) );
  NOR U43957 ( .A(n34136), .B(n30961), .Z(n34555) );
  NOR U43958 ( .A(n30963), .B(n30962), .Z(n30964) );
  NOR U43959 ( .A(n34555), .B(n30964), .Z(n30969) );
  NOR U43960 ( .A(n30965), .B(n30969), .Z(n30966) );
  NOR U43961 ( .A(n34552), .B(n30966), .Z(n30967) );
  NOR U43962 ( .A(n30968), .B(n30967), .Z(n30972) );
  IV U43963 ( .A(n30968), .Z(n30971) );
  IV U43964 ( .A(n30969), .Z(n30970) );
  NOR U43965 ( .A(n30971), .B(n30970), .Z(n34547) );
  NOR U43966 ( .A(n30972), .B(n34547), .Z(n30981) );
  XOR U43967 ( .A(n30982), .B(n30981), .Z(n30976) );
  NOR U43968 ( .A(n30974), .B(n30973), .Z(n30975) );
  NOR U43969 ( .A(n30976), .B(n30975), .Z(n30993) );
  IV U43970 ( .A(n30977), .Z(n30987) );
  IV U43971 ( .A(n30978), .Z(n30979) );
  NOR U43972 ( .A(n30980), .B(n30979), .Z(n30985) );
  IV U43973 ( .A(n30981), .Z(n31336) );
  NOR U43974 ( .A(n30982), .B(n31336), .Z(n30983) );
  IV U43975 ( .A(n30983), .Z(n30984) );
  NOR U43976 ( .A(n30985), .B(n30984), .Z(n30986) );
  IV U43977 ( .A(n30986), .Z(n30989) );
  NOR U43978 ( .A(n30987), .B(n30989), .Z(n34149) );
  IV U43979 ( .A(n30988), .Z(n30990) );
  NOR U43980 ( .A(n30990), .B(n30989), .Z(n37593) );
  NOR U43981 ( .A(n34149), .B(n37593), .Z(n30991) );
  IV U43982 ( .A(n30991), .Z(n30992) );
  NOR U43983 ( .A(n30993), .B(n30992), .Z(n30994) );
  IV U43984 ( .A(n30994), .Z(n34154) );
  IV U43985 ( .A(n30995), .Z(n34155) );
  NOR U43986 ( .A(n30996), .B(n34155), .Z(n30997) );
  XOR U43987 ( .A(n34154), .B(n30997), .Z(n31333) );
  XOR U43988 ( .A(n31332), .B(n31333), .Z(n34166) );
  IV U43989 ( .A(n30998), .Z(n31000) );
  NOR U43990 ( .A(n31000), .B(n30999), .Z(n34164) );
  XOR U43991 ( .A(n34166), .B(n34164), .Z(n34168) );
  XOR U43992 ( .A(n34167), .B(n34168), .Z(n34172) );
  IV U43993 ( .A(n34172), .Z(n31009) );
  IV U43994 ( .A(n31003), .Z(n31002) );
  NOR U43995 ( .A(n31002), .B(n31001), .Z(n34171) );
  NOR U43996 ( .A(n31004), .B(n31003), .Z(n31007) );
  IV U43997 ( .A(n31005), .Z(n31006) );
  NOR U43998 ( .A(n31007), .B(n31006), .Z(n31330) );
  NOR U43999 ( .A(n34171), .B(n31330), .Z(n31008) );
  XOR U44000 ( .A(n31009), .B(n31008), .Z(n31326) );
  IV U44001 ( .A(n31010), .Z(n31012) );
  NOR U44002 ( .A(n31012), .B(n31011), .Z(n31324) );
  XOR U44003 ( .A(n31326), .B(n31324), .Z(n31329) );
  XOR U44004 ( .A(n31327), .B(n31329), .Z(n34175) );
  XOR U44005 ( .A(n34174), .B(n34175), .Z(n34177) );
  XOR U44006 ( .A(n31013), .B(n34177), .Z(n34186) );
  XOR U44007 ( .A(n34185), .B(n34186), .Z(n31312) );
  XOR U44008 ( .A(n31014), .B(n31312), .Z(n31015) );
  IV U44009 ( .A(n31015), .Z(n31310) );
  XOR U44010 ( .A(n31308), .B(n31310), .Z(n31305) );
  IV U44011 ( .A(n31016), .Z(n31025) );
  IV U44012 ( .A(n31017), .Z(n31018) );
  NOR U44013 ( .A(n31025), .B(n31018), .Z(n31303) );
  IV U44014 ( .A(n31019), .Z(n31021) );
  NOR U44015 ( .A(n31021), .B(n31020), .Z(n31306) );
  NOR U44016 ( .A(n31303), .B(n31306), .Z(n31022) );
  XOR U44017 ( .A(n31305), .B(n31022), .Z(n31298) );
  IV U44018 ( .A(n31023), .Z(n31024) );
  NOR U44019 ( .A(n31025), .B(n31024), .Z(n31301) );
  NOR U44020 ( .A(n34504), .B(n31026), .Z(n31027) );
  NOR U44021 ( .A(n31027), .B(n34505), .Z(n31299) );
  NOR U44022 ( .A(n31301), .B(n31299), .Z(n31028) );
  XOR U44023 ( .A(n31298), .B(n31028), .Z(n31297) );
  NOR U44024 ( .A(n31029), .B(n31297), .Z(n37625) );
  IV U44025 ( .A(n31030), .Z(n31032) );
  NOR U44026 ( .A(n31032), .B(n31031), .Z(n31295) );
  XOR U44027 ( .A(n31297), .B(n31295), .Z(n31038) );
  IV U44028 ( .A(n31038), .Z(n31033) );
  NOR U44029 ( .A(n31034), .B(n31033), .Z(n31035) );
  NOR U44030 ( .A(n37625), .B(n31035), .Z(n31036) );
  NOR U44031 ( .A(n31037), .B(n31036), .Z(n31040) );
  IV U44032 ( .A(n31037), .Z(n31039) );
  NOR U44033 ( .A(n31039), .B(n31038), .Z(n37628) );
  NOR U44034 ( .A(n31040), .B(n37628), .Z(n31041) );
  IV U44035 ( .A(n31041), .Z(n34195) );
  XOR U44036 ( .A(n31042), .B(n34195), .Z(n31281) );
  NOR U44037 ( .A(n31043), .B(n31289), .Z(n31047) );
  IV U44038 ( .A(n31044), .Z(n31282) );
  NOR U44039 ( .A(n31045), .B(n31282), .Z(n31046) );
  NOR U44040 ( .A(n31047), .B(n31046), .Z(n31048) );
  XOR U44041 ( .A(n31281), .B(n31048), .Z(n31276) );
  NOR U44042 ( .A(n31049), .B(n34205), .Z(n31053) );
  IV U44043 ( .A(n31050), .Z(n31277) );
  NOR U44044 ( .A(n31051), .B(n31277), .Z(n31052) );
  NOR U44045 ( .A(n31053), .B(n31052), .Z(n31054) );
  XOR U44046 ( .A(n31276), .B(n31054), .Z(n34221) );
  XOR U44047 ( .A(n34219), .B(n34221), .Z(n31062) );
  IV U44048 ( .A(n31055), .Z(n31057) );
  NOR U44049 ( .A(n31057), .B(n31056), .Z(n34220) );
  IV U44050 ( .A(n31058), .Z(n31060) );
  IV U44051 ( .A(n31059), .Z(n31064) );
  NOR U44052 ( .A(n31060), .B(n31064), .Z(n31273) );
  NOR U44053 ( .A(n34220), .B(n31273), .Z(n31061) );
  XOR U44054 ( .A(n31062), .B(n31061), .Z(n31272) );
  IV U44055 ( .A(n31063), .Z(n31065) );
  NOR U44056 ( .A(n31065), .B(n31064), .Z(n31066) );
  IV U44057 ( .A(n31066), .Z(n31271) );
  XOR U44058 ( .A(n31272), .B(n31271), .Z(n31073) );
  IV U44059 ( .A(n31073), .Z(n31067) );
  NOR U44060 ( .A(n31068), .B(n31067), .Z(n37664) );
  IV U44061 ( .A(n31069), .Z(n31070) );
  NOR U44062 ( .A(n31071), .B(n31070), .Z(n31074) );
  IV U44063 ( .A(n31074), .Z(n31072) );
  NOR U44064 ( .A(n31272), .B(n31072), .Z(n37661) );
  NOR U44065 ( .A(n31074), .B(n31073), .Z(n31075) );
  NOR U44066 ( .A(n37661), .B(n31075), .Z(n31076) );
  NOR U44067 ( .A(n31077), .B(n31076), .Z(n31078) );
  NOR U44068 ( .A(n37664), .B(n31078), .Z(n31079) );
  IV U44069 ( .A(n31079), .Z(n34226) );
  XOR U44070 ( .A(n34225), .B(n34226), .Z(n34238) );
  XOR U44071 ( .A(n34229), .B(n34238), .Z(n34231) );
  XOR U44072 ( .A(n34232), .B(n34231), .Z(n31080) );
  XOR U44073 ( .A(n31081), .B(n31080), .Z(n34235) );
  IV U44074 ( .A(n31082), .Z(n31084) );
  NOR U44075 ( .A(n31084), .B(n31083), .Z(n34233) );
  XOR U44076 ( .A(n34235), .B(n34233), .Z(n31267) );
  XOR U44077 ( .A(n31266), .B(n31267), .Z(n31260) );
  XOR U44078 ( .A(n31259), .B(n31260), .Z(n31093) );
  IV U44079 ( .A(n31093), .Z(n31090) );
  NOR U44080 ( .A(n31085), .B(n31090), .Z(n34467) );
  IV U44081 ( .A(n31086), .Z(n31088) );
  NOR U44082 ( .A(n31088), .B(n31087), .Z(n31097) );
  IV U44083 ( .A(n31097), .Z(n31089) );
  NOR U44084 ( .A(n31090), .B(n31089), .Z(n34471) );
  NOR U44085 ( .A(n31091), .B(n31262), .Z(n31094) );
  IV U44086 ( .A(n31094), .Z(n31092) );
  NOR U44087 ( .A(n31092), .B(n31267), .Z(n31257) );
  NOR U44088 ( .A(n31094), .B(n31093), .Z(n31095) );
  NOR U44089 ( .A(n31257), .B(n31095), .Z(n31096) );
  NOR U44090 ( .A(n31097), .B(n31096), .Z(n31098) );
  NOR U44091 ( .A(n34471), .B(n31098), .Z(n31253) );
  NOR U44092 ( .A(n31099), .B(n31253), .Z(n31100) );
  NOR U44093 ( .A(n34467), .B(n31100), .Z(n31248) );
  NOR U44094 ( .A(n34461), .B(n31101), .Z(n31252) );
  IV U44095 ( .A(n31102), .Z(n31249) );
  NOR U44096 ( .A(n31103), .B(n31249), .Z(n31104) );
  NOR U44097 ( .A(n31252), .B(n31104), .Z(n31105) );
  XOR U44098 ( .A(n31248), .B(n31105), .Z(n34247) );
  IV U44099 ( .A(n31106), .Z(n31108) );
  NOR U44100 ( .A(n31108), .B(n31107), .Z(n34245) );
  XOR U44101 ( .A(n34247), .B(n34245), .Z(n34255) );
  XOR U44102 ( .A(n31243), .B(n34255), .Z(n31109) );
  IV U44103 ( .A(n31109), .Z(n34257) );
  XOR U44104 ( .A(n34256), .B(n34257), .Z(n34260) );
  XOR U44105 ( .A(n34259), .B(n34260), .Z(n31241) );
  XOR U44106 ( .A(n31240), .B(n31241), .Z(n34285) );
  IV U44107 ( .A(n31110), .Z(n34269) );
  NOR U44108 ( .A(n34269), .B(n31111), .Z(n31114) );
  IV U44109 ( .A(n31112), .Z(n31113) );
  NOR U44110 ( .A(n31113), .B(n31120), .Z(n34283) );
  NOR U44111 ( .A(n31114), .B(n34283), .Z(n31115) );
  XOR U44112 ( .A(n34285), .B(n31115), .Z(n34280) );
  IV U44113 ( .A(n31116), .Z(n31125) );
  IV U44114 ( .A(n31117), .Z(n31118) );
  NOR U44115 ( .A(n31125), .B(n31118), .Z(n34287) );
  IV U44116 ( .A(n31119), .Z(n31121) );
  NOR U44117 ( .A(n31121), .B(n31120), .Z(n34281) );
  NOR U44118 ( .A(n34287), .B(n34281), .Z(n31122) );
  XOR U44119 ( .A(n34280), .B(n31122), .Z(n34304) );
  IV U44120 ( .A(n31123), .Z(n31124) );
  NOR U44121 ( .A(n31125), .B(n31124), .Z(n31126) );
  IV U44122 ( .A(n31126), .Z(n34294) );
  XOR U44123 ( .A(n34304), .B(n34294), .Z(n31127) );
  XOR U44124 ( .A(n31128), .B(n31127), .Z(n31236) );
  IV U44125 ( .A(n31129), .Z(n31131) );
  NOR U44126 ( .A(n31131), .B(n31130), .Z(n31234) );
  XOR U44127 ( .A(n31236), .B(n31234), .Z(n31238) );
  XOR U44128 ( .A(n31132), .B(n31238), .Z(n31133) );
  IV U44129 ( .A(n31133), .Z(n34307) );
  XOR U44130 ( .A(n34306), .B(n34307), .Z(n34311) );
  IV U44131 ( .A(n31134), .Z(n31137) );
  IV U44132 ( .A(n31135), .Z(n31136) );
  NOR U44133 ( .A(n31137), .B(n31136), .Z(n34309) );
  XOR U44134 ( .A(n34311), .B(n34309), .Z(n31231) );
  NOR U44135 ( .A(n31223), .B(n31138), .Z(n31143) );
  IV U44136 ( .A(n31139), .Z(n31142) );
  IV U44137 ( .A(n31140), .Z(n31141) );
  NOR U44138 ( .A(n31142), .B(n31141), .Z(n31229) );
  NOR U44139 ( .A(n31143), .B(n31229), .Z(n31144) );
  XOR U44140 ( .A(n31231), .B(n31144), .Z(n31220) );
  IV U44141 ( .A(n31145), .Z(n37726) );
  NOR U44142 ( .A(n31146), .B(n37726), .Z(n31219) );
  IV U44143 ( .A(n31147), .Z(n31148) );
  NOR U44144 ( .A(n31148), .B(n31153), .Z(n34315) );
  NOR U44145 ( .A(n31219), .B(n34315), .Z(n31149) );
  XOR U44146 ( .A(n31220), .B(n31149), .Z(n34318) );
  IV U44147 ( .A(n31150), .Z(n34319) );
  NOR U44148 ( .A(n34319), .B(n31151), .Z(n31155) );
  IV U44149 ( .A(n31152), .Z(n31154) );
  NOR U44150 ( .A(n31154), .B(n31153), .Z(n31216) );
  NOR U44151 ( .A(n31155), .B(n31216), .Z(n31156) );
  XOR U44152 ( .A(n34318), .B(n31156), .Z(n34331) );
  NOR U44153 ( .A(n31157), .B(n31213), .Z(n31161) );
  IV U44154 ( .A(n31158), .Z(n31160) );
  NOR U44155 ( .A(n31160), .B(n31159), .Z(n34332) );
  NOR U44156 ( .A(n31161), .B(n34332), .Z(n31162) );
  XOR U44157 ( .A(n34331), .B(n31162), .Z(n34343) );
  XOR U44158 ( .A(n34340), .B(n34343), .Z(n37745) );
  NOR U44159 ( .A(n31163), .B(n34344), .Z(n31170) );
  IV U44160 ( .A(n31164), .Z(n31165) );
  NOR U44161 ( .A(n31165), .B(n31167), .Z(n37743) );
  IV U44162 ( .A(n31166), .Z(n31168) );
  NOR U44163 ( .A(n31168), .B(n31167), .Z(n37750) );
  NOR U44164 ( .A(n37743), .B(n37750), .Z(n31208) );
  IV U44165 ( .A(n31208), .Z(n31169) );
  NOR U44166 ( .A(n31170), .B(n31169), .Z(n31171) );
  XOR U44167 ( .A(n37745), .B(n31171), .Z(n31203) );
  IV U44168 ( .A(n31172), .Z(n31174) );
  NOR U44169 ( .A(n31174), .B(n31173), .Z(n31204) );
  IV U44170 ( .A(n31204), .Z(n31201) );
  XOR U44171 ( .A(n31203), .B(n31201), .Z(n31175) );
  XOR U44172 ( .A(n31176), .B(n31175), .Z(n31177) );
  IV U44173 ( .A(n31177), .Z(n34359) );
  XOR U44174 ( .A(n34357), .B(n34359), .Z(n34361) );
  IV U44175 ( .A(n34361), .Z(n31181) );
  NOR U44176 ( .A(n31179), .B(n31178), .Z(n34360) );
  NOR U44177 ( .A(n34360), .B(n31197), .Z(n31180) );
  XOR U44178 ( .A(n31181), .B(n31180), .Z(n37771) );
  XOR U44179 ( .A(n31192), .B(n37771), .Z(n31195) );
  XOR U44180 ( .A(n31194), .B(n31195), .Z(n34370) );
  XOR U44181 ( .A(n31182), .B(n34370), .Z(n31183) );
  IV U44182 ( .A(n31183), .Z(n31191) );
  XOR U44183 ( .A(n31189), .B(n31191), .Z(n34398) );
  NOR U44184 ( .A(n34376), .B(n34398), .Z(n31184) );
  IV U44185 ( .A(n31184), .Z(n34392) );
  IV U44186 ( .A(n31185), .Z(n31187) );
  NOR U44187 ( .A(n31187), .B(n31186), .Z(n34375) );
  IV U44188 ( .A(n34375), .Z(n31188) );
  NOR U44189 ( .A(n34392), .B(n31188), .Z(n34403) );
  IV U44190 ( .A(n31189), .Z(n31190) );
  NOR U44191 ( .A(n31191), .B(n31190), .Z(n34400) );
  IV U44192 ( .A(n31192), .Z(n31193) );
  NOR U44193 ( .A(n37771), .B(n31193), .Z(n34409) );
  IV U44194 ( .A(n31194), .Z(n31196) );
  NOR U44195 ( .A(n31196), .B(n31195), .Z(n34406) );
  NOR U44196 ( .A(n34409), .B(n34406), .Z(n34365) );
  IV U44197 ( .A(n31197), .Z(n31198) );
  NOR U44198 ( .A(n31198), .B(n34361), .Z(n37755) );
  IV U44199 ( .A(n31203), .Z(n31202) );
  IV U44200 ( .A(n31199), .Z(n31200) );
  NOR U44201 ( .A(n31202), .B(n31200), .Z(n34412) );
  NOR U44202 ( .A(n31202), .B(n31201), .Z(n34420) );
  NOR U44203 ( .A(n31204), .B(n31203), .Z(n31207) );
  IV U44204 ( .A(n31205), .Z(n31206) );
  NOR U44205 ( .A(n31207), .B(n31206), .Z(n34417) );
  NOR U44206 ( .A(n34420), .B(n34417), .Z(n31210) );
  NOR U44207 ( .A(n37745), .B(n31208), .Z(n31209) );
  XOR U44208 ( .A(n31210), .B(n31209), .Z(n34356) );
  IV U44209 ( .A(n31211), .Z(n31215) );
  XOR U44210 ( .A(n31216), .B(n34318), .Z(n31212) );
  NOR U44211 ( .A(n31213), .B(n31212), .Z(n31214) );
  IV U44212 ( .A(n31214), .Z(n34336) );
  NOR U44213 ( .A(n31215), .B(n34336), .Z(n34427) );
  IV U44214 ( .A(n31216), .Z(n31217) );
  NOR U44215 ( .A(n31217), .B(n34318), .Z(n31218) );
  IV U44216 ( .A(n31218), .Z(n34322) );
  IV U44217 ( .A(n31219), .Z(n31221) );
  IV U44218 ( .A(n31220), .Z(n37723) );
  NOR U44219 ( .A(n31221), .B(n37723), .Z(n34314) );
  IV U44220 ( .A(n31222), .Z(n31225) );
  NOR U44221 ( .A(n31223), .B(n31231), .Z(n31224) );
  IV U44222 ( .A(n31224), .Z(n31227) );
  NOR U44223 ( .A(n31225), .B(n31227), .Z(n37718) );
  IV U44224 ( .A(n31226), .Z(n31228) );
  NOR U44225 ( .A(n31228), .B(n31227), .Z(n37714) );
  IV U44226 ( .A(n31229), .Z(n31230) );
  NOR U44227 ( .A(n31231), .B(n31230), .Z(n37711) );
  IV U44228 ( .A(n31232), .Z(n31233) );
  NOR U44229 ( .A(n31233), .B(n31238), .Z(n34436) );
  IV U44230 ( .A(n31234), .Z(n31235) );
  NOR U44231 ( .A(n31236), .B(n31235), .Z(n41068) );
  IV U44232 ( .A(n31237), .Z(n31239) );
  NOR U44233 ( .A(n31239), .B(n31238), .Z(n38016) );
  NOR U44234 ( .A(n41068), .B(n38016), .Z(n34442) );
  IV U44235 ( .A(n31240), .Z(n31242) );
  NOR U44236 ( .A(n31242), .B(n31241), .Z(n34264) );
  NOR U44237 ( .A(n31243), .B(n34255), .Z(n31244) );
  IV U44238 ( .A(n31244), .Z(n31245) );
  NOR U44239 ( .A(n31246), .B(n31245), .Z(n37687) );
  IV U44240 ( .A(n31247), .Z(n31251) );
  IV U44241 ( .A(n31248), .Z(n34458) );
  NOR U44242 ( .A(n31249), .B(n34458), .Z(n31250) );
  IV U44243 ( .A(n31250), .Z(n34249) );
  NOR U44244 ( .A(n31251), .B(n34249), .Z(n34454) );
  IV U44245 ( .A(n31252), .Z(n31255) );
  IV U44246 ( .A(n31253), .Z(n31254) );
  NOR U44247 ( .A(n31255), .B(n31254), .Z(n31256) );
  NOR U44248 ( .A(n34467), .B(n31256), .Z(n34243) );
  IV U44249 ( .A(n31257), .Z(n31258) );
  NOR U44250 ( .A(n31261), .B(n31258), .Z(n34473) );
  NOR U44251 ( .A(n34471), .B(n34473), .Z(n34242) );
  NOR U44252 ( .A(n31260), .B(n31259), .Z(n41306) );
  IV U44253 ( .A(n31261), .Z(n31265) );
  NOR U44254 ( .A(n31262), .B(n31267), .Z(n31263) );
  IV U44255 ( .A(n31263), .Z(n31264) );
  NOR U44256 ( .A(n31265), .B(n31264), .Z(n34476) );
  NOR U44257 ( .A(n41306), .B(n34476), .Z(n34241) );
  IV U44258 ( .A(n31266), .Z(n31268) );
  NOR U44259 ( .A(n31268), .B(n31267), .Z(n44415) );
  IV U44260 ( .A(n31269), .Z(n31270) );
  NOR U44261 ( .A(n31270), .B(n34238), .Z(n37674) );
  NOR U44262 ( .A(n31272), .B(n31271), .Z(n34481) );
  IV U44263 ( .A(n31273), .Z(n31274) );
  NOR U44264 ( .A(n34221), .B(n31274), .Z(n34484) );
  NOR U44265 ( .A(n34481), .B(n34484), .Z(n34224) );
  IV U44266 ( .A(n31275), .Z(n31279) );
  IV U44267 ( .A(n31276), .Z(n34206) );
  NOR U44268 ( .A(n34206), .B(n31277), .Z(n31278) );
  IV U44269 ( .A(n31278), .Z(n34216) );
  NOR U44270 ( .A(n31279), .B(n34216), .Z(n37653) );
  IV U44271 ( .A(n31280), .Z(n31284) );
  NOR U44272 ( .A(n31282), .B(n31281), .Z(n31283) );
  IV U44273 ( .A(n31283), .Z(n31286) );
  NOR U44274 ( .A(n31284), .B(n31286), .Z(n37642) );
  IV U44275 ( .A(n31285), .Z(n31287) );
  NOR U44276 ( .A(n31287), .B(n31286), .Z(n34490) );
  IV U44277 ( .A(n31288), .Z(n31291) );
  NOR U44278 ( .A(n31289), .B(n34195), .Z(n31290) );
  IV U44279 ( .A(n31290), .Z(n31293) );
  NOR U44280 ( .A(n31291), .B(n31293), .Z(n37638) );
  IV U44281 ( .A(n31292), .Z(n31294) );
  NOR U44282 ( .A(n31294), .B(n31293), .Z(n37635) );
  IV U44283 ( .A(n31295), .Z(n31296) );
  NOR U44284 ( .A(n31297), .B(n31296), .Z(n34497) );
  IV U44285 ( .A(n31298), .Z(n34509) );
  IV U44286 ( .A(n31299), .Z(n31300) );
  NOR U44287 ( .A(n34509), .B(n31300), .Z(n34500) );
  IV U44288 ( .A(n31301), .Z(n31302) );
  NOR U44289 ( .A(n34509), .B(n31302), .Z(n34513) );
  IV U44290 ( .A(n31303), .Z(n31304) );
  NOR U44291 ( .A(n31305), .B(n31304), .Z(n34515) );
  NOR U44292 ( .A(n34513), .B(n34515), .Z(n34192) );
  IV U44293 ( .A(n31306), .Z(n31307) );
  NOR U44294 ( .A(n31310), .B(n31307), .Z(n37620) );
  IV U44295 ( .A(n31308), .Z(n31309) );
  NOR U44296 ( .A(n31310), .B(n31309), .Z(n37617) );
  IV U44297 ( .A(n31311), .Z(n31313) );
  NOR U44298 ( .A(n31313), .B(n31312), .Z(n37613) );
  IV U44299 ( .A(n31314), .Z(n31317) );
  NOR U44300 ( .A(n31315), .B(n34186), .Z(n31316) );
  IV U44301 ( .A(n31316), .Z(n34181) );
  NOR U44302 ( .A(n31317), .B(n34181), .Z(n31318) );
  IV U44303 ( .A(n31318), .Z(n37612) );
  IV U44304 ( .A(n31319), .Z(n31320) );
  NOR U44305 ( .A(n31320), .B(n34177), .Z(n34521) );
  XOR U44306 ( .A(n31321), .B(n34177), .Z(n31322) );
  NOR U44307 ( .A(n31323), .B(n31322), .Z(n34518) );
  IV U44308 ( .A(n31324), .Z(n31325) );
  NOR U44309 ( .A(n31326), .B(n31325), .Z(n40936) );
  IV U44310 ( .A(n31327), .Z(n31328) );
  NOR U44311 ( .A(n31329), .B(n31328), .Z(n40941) );
  NOR U44312 ( .A(n40936), .B(n40941), .Z(n34526) );
  IV U44313 ( .A(n31330), .Z(n31331) );
  NOR U44314 ( .A(n34172), .B(n31331), .Z(n34534) );
  IV U44315 ( .A(n31332), .Z(n31334) );
  NOR U44316 ( .A(n31334), .B(n31333), .Z(n34162) );
  IV U44317 ( .A(n34162), .Z(n34152) );
  IV U44318 ( .A(n34149), .Z(n34140) );
  IV U44319 ( .A(n31335), .Z(n31339) );
  NOR U44320 ( .A(n31337), .B(n31336), .Z(n31338) );
  IV U44321 ( .A(n31338), .Z(n34142) );
  NOR U44322 ( .A(n31339), .B(n34142), .Z(n31340) );
  IV U44323 ( .A(n31340), .Z(n34546) );
  IV U44324 ( .A(n31341), .Z(n31344) );
  NOR U44325 ( .A(n31342), .B(n31347), .Z(n31343) );
  IV U44326 ( .A(n31343), .Z(n31349) );
  NOR U44327 ( .A(n31344), .B(n31349), .Z(n34557) );
  IV U44328 ( .A(n31345), .Z(n31346) );
  NOR U44329 ( .A(n31347), .B(n31346), .Z(n37587) );
  IV U44330 ( .A(n31348), .Z(n31350) );
  NOR U44331 ( .A(n31350), .B(n31349), .Z(n34563) );
  NOR U44332 ( .A(n37587), .B(n34563), .Z(n34132) );
  IV U44333 ( .A(n31351), .Z(n31352) );
  NOR U44334 ( .A(n31354), .B(n31352), .Z(n37583) );
  IV U44335 ( .A(n31353), .Z(n31355) );
  NOR U44336 ( .A(n31355), .B(n31354), .Z(n37580) );
  IV U44337 ( .A(n31356), .Z(n31359) );
  NOR U44338 ( .A(n31357), .B(n34125), .Z(n31358) );
  IV U44339 ( .A(n31358), .Z(n34130) );
  NOR U44340 ( .A(n31359), .B(n34130), .Z(n34568) );
  IV U44341 ( .A(n31360), .Z(n31361) );
  NOR U44342 ( .A(n31362), .B(n31361), .Z(n31363) );
  IV U44343 ( .A(n31363), .Z(n34571) );
  IV U44344 ( .A(n31364), .Z(n31365) );
  NOR U44345 ( .A(n34113), .B(n31365), .Z(n37572) );
  NOR U44346 ( .A(n31367), .B(n31366), .Z(n31368) );
  IV U44347 ( .A(n31368), .Z(n31369) );
  NOR U44348 ( .A(n31369), .B(n34599), .Z(n34108) );
  IV U44349 ( .A(n31370), .Z(n31371) );
  NOR U44350 ( .A(n31373), .B(n31371), .Z(n34606) );
  NOR U44351 ( .A(n34606), .B(n34604), .Z(n34106) );
  IV U44352 ( .A(n31372), .Z(n31374) );
  NOR U44353 ( .A(n31374), .B(n31373), .Z(n37565) );
  IV U44354 ( .A(n31375), .Z(n31378) );
  NOR U44355 ( .A(n31376), .B(n31382), .Z(n31377) );
  IV U44356 ( .A(n31377), .Z(n31380) );
  NOR U44357 ( .A(n31378), .B(n31380), .Z(n37562) );
  IV U44358 ( .A(n31379), .Z(n31381) );
  NOR U44359 ( .A(n31381), .B(n31380), .Z(n34100) );
  IV U44360 ( .A(n34100), .Z(n34094) );
  NOR U44361 ( .A(n31383), .B(n31382), .Z(n34609) );
  IV U44362 ( .A(n31384), .Z(n31388) );
  IV U44363 ( .A(n31385), .Z(n31397) );
  NOR U44364 ( .A(n31397), .B(n31400), .Z(n31386) );
  IV U44365 ( .A(n31386), .Z(n31387) );
  NOR U44366 ( .A(n31388), .B(n31387), .Z(n34617) );
  IV U44367 ( .A(n31389), .Z(n31394) );
  NOR U44368 ( .A(n31391), .B(n31390), .Z(n31392) );
  IV U44369 ( .A(n31392), .Z(n31393) );
  NOR U44370 ( .A(n31394), .B(n31393), .Z(n34615) );
  NOR U44371 ( .A(n34617), .B(n34615), .Z(n34093) );
  IV U44372 ( .A(n31395), .Z(n31396) );
  NOR U44373 ( .A(n31396), .B(n31400), .Z(n34622) );
  NOR U44374 ( .A(n31398), .B(n31397), .Z(n31399) );
  IV U44375 ( .A(n31399), .Z(n31401) );
  NOR U44376 ( .A(n31401), .B(n31400), .Z(n34620) );
  NOR U44377 ( .A(n34622), .B(n34620), .Z(n34092) );
  NOR U44378 ( .A(n31403), .B(n31402), .Z(n31404) );
  IV U44379 ( .A(n31404), .Z(n34630) );
  IV U44380 ( .A(n31405), .Z(n31406) );
  NOR U44381 ( .A(n31407), .B(n31406), .Z(n38181) );
  IV U44382 ( .A(n31408), .Z(n31413) );
  IV U44383 ( .A(n31409), .Z(n31410) );
  NOR U44384 ( .A(n31411), .B(n31410), .Z(n31412) );
  IV U44385 ( .A(n31412), .Z(n31415) );
  NOR U44386 ( .A(n31413), .B(n31415), .Z(n38186) );
  NOR U44387 ( .A(n38181), .B(n38186), .Z(n34627) );
  IV U44388 ( .A(n31414), .Z(n31416) );
  NOR U44389 ( .A(n31416), .B(n31415), .Z(n34635) );
  NOR U44390 ( .A(n31418), .B(n31417), .Z(n34646) );
  NOR U44391 ( .A(n31420), .B(n31419), .Z(n34651) );
  NOR U44392 ( .A(n34651), .B(n34649), .Z(n34085) );
  IV U44393 ( .A(n31421), .Z(n31422) );
  NOR U44394 ( .A(n34083), .B(n31422), .Z(n34657) );
  IV U44395 ( .A(n31423), .Z(n31424) );
  NOR U44396 ( .A(n31425), .B(n31424), .Z(n37521) );
  IV U44397 ( .A(n31425), .Z(n31429) );
  NOR U44398 ( .A(n31426), .B(n37524), .Z(n31427) );
  IV U44399 ( .A(n31427), .Z(n31428) );
  NOR U44400 ( .A(n31429), .B(n31428), .Z(n34673) );
  IV U44401 ( .A(n31430), .Z(n34685) );
  NOR U44402 ( .A(n34685), .B(n31431), .Z(n31434) );
  NOR U44403 ( .A(n31433), .B(n31432), .Z(n34676) );
  NOR U44404 ( .A(n31434), .B(n34676), .Z(n34052) );
  NOR U44405 ( .A(n44188), .B(n44194), .Z(n37515) );
  NOR U44406 ( .A(n37517), .B(n37515), .Z(n34051) );
  IV U44407 ( .A(n31435), .Z(n31436) );
  NOR U44408 ( .A(n47688), .B(n31436), .Z(n34043) );
  IV U44409 ( .A(n34043), .Z(n34038) );
  IV U44410 ( .A(n31437), .Z(n31440) );
  NOR U44411 ( .A(n31438), .B(n31447), .Z(n31439) );
  IV U44412 ( .A(n31439), .Z(n31443) );
  NOR U44413 ( .A(n31440), .B(n31443), .Z(n31441) );
  IV U44414 ( .A(n31441), .Z(n37509) );
  IV U44415 ( .A(n31442), .Z(n31444) );
  NOR U44416 ( .A(n31444), .B(n31443), .Z(n37505) );
  IV U44417 ( .A(n31445), .Z(n31446) );
  NOR U44418 ( .A(n31447), .B(n31446), .Z(n37502) );
  IV U44419 ( .A(n31448), .Z(n31449) );
  NOR U44420 ( .A(n31450), .B(n31449), .Z(n34704) );
  NOR U44421 ( .A(n37502), .B(n34704), .Z(n34031) );
  NOR U44422 ( .A(n31452), .B(n31451), .Z(n34030) );
  IV U44423 ( .A(n31453), .Z(n31455) );
  NOR U44424 ( .A(n31455), .B(n31454), .Z(n37477) );
  IV U44425 ( .A(n31456), .Z(n31459) );
  NOR U44426 ( .A(n31457), .B(n31461), .Z(n31458) );
  IV U44427 ( .A(n31458), .Z(n31464) );
  NOR U44428 ( .A(n31459), .B(n31464), .Z(n37473) );
  NOR U44429 ( .A(n37477), .B(n37473), .Z(n34025) );
  IV U44430 ( .A(n31460), .Z(n31462) );
  NOR U44431 ( .A(n31462), .B(n31461), .Z(n34712) );
  IV U44432 ( .A(n31463), .Z(n31465) );
  NOR U44433 ( .A(n31465), .B(n31464), .Z(n34710) );
  NOR U44434 ( .A(n34712), .B(n34710), .Z(n34024) );
  IV U44435 ( .A(n31466), .Z(n31467) );
  NOR U44436 ( .A(n37460), .B(n31467), .Z(n31476) );
  IV U44437 ( .A(n31468), .Z(n31469) );
  NOR U44438 ( .A(n31470), .B(n31469), .Z(n34715) );
  IV U44439 ( .A(n31471), .Z(n31472) );
  NOR U44440 ( .A(n31473), .B(n31472), .Z(n37470) );
  NOR U44441 ( .A(n34715), .B(n37470), .Z(n31474) );
  IV U44442 ( .A(n31474), .Z(n31475) );
  NOR U44443 ( .A(n31476), .B(n31475), .Z(n34023) );
  IV U44444 ( .A(n31477), .Z(n31480) );
  NOR U44445 ( .A(n31478), .B(n31483), .Z(n31479) );
  IV U44446 ( .A(n31479), .Z(n31485) );
  NOR U44447 ( .A(n31480), .B(n31485), .Z(n34020) );
  IV U44448 ( .A(n31481), .Z(n31482) );
  NOR U44449 ( .A(n31483), .B(n31482), .Z(n37453) );
  IV U44450 ( .A(n31484), .Z(n31486) );
  NOR U44451 ( .A(n31486), .B(n31485), .Z(n37455) );
  NOR U44452 ( .A(n37453), .B(n37455), .Z(n34019) );
  IV U44453 ( .A(n31487), .Z(n31489) );
  NOR U44454 ( .A(n31489), .B(n31488), .Z(n37448) );
  IV U44455 ( .A(n31490), .Z(n31494) );
  IV U44456 ( .A(n31491), .Z(n34010) );
  NOR U44457 ( .A(n34010), .B(n31492), .Z(n31493) );
  IV U44458 ( .A(n31493), .Z(n31496) );
  NOR U44459 ( .A(n31494), .B(n31496), .Z(n37445) );
  IV U44460 ( .A(n31495), .Z(n31497) );
  NOR U44461 ( .A(n31497), .B(n31496), .Z(n37441) );
  NOR U44462 ( .A(n34010), .B(n31498), .Z(n31499) );
  IV U44463 ( .A(n31499), .Z(n31500) );
  NOR U44464 ( .A(n34008), .B(n31500), .Z(n37438) );
  IV U44465 ( .A(n31501), .Z(n31504) );
  NOR U44466 ( .A(n31502), .B(n31506), .Z(n31503) );
  IV U44467 ( .A(n31503), .Z(n34015) );
  NOR U44468 ( .A(n31504), .B(n34015), .Z(n37428) );
  IV U44469 ( .A(n31505), .Z(n31509) );
  NOR U44470 ( .A(n31507), .B(n31506), .Z(n31508) );
  IV U44471 ( .A(n31508), .Z(n31517) );
  NOR U44472 ( .A(n31509), .B(n31517), .Z(n31510) );
  IV U44473 ( .A(n31510), .Z(n34721) );
  IV U44474 ( .A(n31511), .Z(n31515) );
  NOR U44475 ( .A(n31513), .B(n31512), .Z(n31514) );
  IV U44476 ( .A(n31514), .Z(n31520) );
  NOR U44477 ( .A(n31515), .B(n31520), .Z(n34726) );
  IV U44478 ( .A(n31516), .Z(n31518) );
  NOR U44479 ( .A(n31518), .B(n31517), .Z(n37425) );
  NOR U44480 ( .A(n34726), .B(n37425), .Z(n34007) );
  IV U44481 ( .A(n31519), .Z(n31521) );
  NOR U44482 ( .A(n31521), .B(n31520), .Z(n34723) );
  IV U44483 ( .A(n31522), .Z(n31526) );
  NOR U44484 ( .A(n31524), .B(n31523), .Z(n31525) );
  IV U44485 ( .A(n31525), .Z(n34005) );
  NOR U44486 ( .A(n31526), .B(n34005), .Z(n37421) );
  IV U44487 ( .A(n31527), .Z(n31531) );
  NOR U44488 ( .A(n31529), .B(n31528), .Z(n31530) );
  IV U44489 ( .A(n31530), .Z(n31533) );
  NOR U44490 ( .A(n31531), .B(n31533), .Z(n34735) );
  IV U44491 ( .A(n31532), .Z(n31534) );
  NOR U44492 ( .A(n31534), .B(n31533), .Z(n34737) );
  NOR U44493 ( .A(n34735), .B(n34737), .Z(n33999) );
  IV U44494 ( .A(n31535), .Z(n31539) );
  IV U44495 ( .A(n31536), .Z(n31545) );
  NOR U44496 ( .A(n31537), .B(n31545), .Z(n31538) );
  IV U44497 ( .A(n31538), .Z(n31541) );
  NOR U44498 ( .A(n31539), .B(n31541), .Z(n34742) );
  IV U44499 ( .A(n31540), .Z(n31542) );
  NOR U44500 ( .A(n31542), .B(n31541), .Z(n34745) );
  IV U44501 ( .A(n31543), .Z(n31544) );
  NOR U44502 ( .A(n31545), .B(n31544), .Z(n37400) );
  NOR U44503 ( .A(n31547), .B(n31546), .Z(n38291) );
  IV U44504 ( .A(n31548), .Z(n31549) );
  NOR U44505 ( .A(n31549), .B(n31559), .Z(n38295) );
  NOR U44506 ( .A(n38291), .B(n38295), .Z(n34749) );
  IV U44507 ( .A(n31550), .Z(n31553) );
  NOR U44508 ( .A(n31551), .B(n33996), .Z(n31552) );
  IV U44509 ( .A(n31552), .Z(n31563) );
  NOR U44510 ( .A(n31553), .B(n31563), .Z(n37392) );
  IV U44511 ( .A(n31554), .Z(n31555) );
  NOR U44512 ( .A(n31556), .B(n31555), .Z(n34750) );
  IV U44513 ( .A(n31557), .Z(n31558) );
  NOR U44514 ( .A(n31559), .B(n31558), .Z(n37395) );
  NOR U44515 ( .A(n34750), .B(n37395), .Z(n31560) );
  IV U44516 ( .A(n31560), .Z(n31561) );
  NOR U44517 ( .A(n37392), .B(n31561), .Z(n33998) );
  IV U44518 ( .A(n31562), .Z(n31564) );
  NOR U44519 ( .A(n31564), .B(n31563), .Z(n37389) );
  XOR U44520 ( .A(n33978), .B(n33979), .Z(n31565) );
  NOR U44521 ( .A(n31566), .B(n31565), .Z(n33985) );
  IV U44522 ( .A(n33985), .Z(n33977) );
  IV U44523 ( .A(n31567), .Z(n31568) );
  NOR U44524 ( .A(n31569), .B(n31568), .Z(n38323) );
  IV U44525 ( .A(n31570), .Z(n34765) );
  IV U44526 ( .A(n31571), .Z(n31572) );
  NOR U44527 ( .A(n34765), .B(n31572), .Z(n38318) );
  NOR U44528 ( .A(n38323), .B(n38318), .Z(n34768) );
  IV U44529 ( .A(n34768), .Z(n33974) );
  IV U44530 ( .A(n31573), .Z(n31576) );
  NOR U44531 ( .A(n31579), .B(n31574), .Z(n31575) );
  IV U44532 ( .A(n31575), .Z(n33972) );
  NOR U44533 ( .A(n31576), .B(n33972), .Z(n37366) );
  IV U44534 ( .A(n31577), .Z(n31578) );
  NOR U44535 ( .A(n31579), .B(n31578), .Z(n34776) );
  NOR U44536 ( .A(n34781), .B(n34779), .Z(n33957) );
  IV U44537 ( .A(n31580), .Z(n31581) );
  NOR U44538 ( .A(n31581), .B(n33907), .Z(n31582) );
  IV U44539 ( .A(n31582), .Z(n31583) );
  NOR U44540 ( .A(n31587), .B(n31583), .Z(n37323) );
  IV U44541 ( .A(n31584), .Z(n31586) );
  NOR U44542 ( .A(n31586), .B(n31585), .Z(n34814) );
  IV U44543 ( .A(n31587), .Z(n31591) );
  NOR U44544 ( .A(n31588), .B(n33907), .Z(n31589) );
  IV U44545 ( .A(n31589), .Z(n31590) );
  NOR U44546 ( .A(n31591), .B(n31590), .Z(n37320) );
  NOR U44547 ( .A(n34814), .B(n37320), .Z(n33904) );
  IV U44548 ( .A(n31592), .Z(n31597) );
  IV U44549 ( .A(n31593), .Z(n31594) );
  NOR U44550 ( .A(n31597), .B(n31594), .Z(n37315) );
  IV U44551 ( .A(n31595), .Z(n31599) );
  NOR U44552 ( .A(n31597), .B(n31596), .Z(n31598) );
  IV U44553 ( .A(n31598), .Z(n31601) );
  NOR U44554 ( .A(n31599), .B(n31601), .Z(n37312) );
  IV U44555 ( .A(n31600), .Z(n31602) );
  NOR U44556 ( .A(n31602), .B(n31601), .Z(n37308) );
  IV U44557 ( .A(n31603), .Z(n31607) );
  NOR U44558 ( .A(n31605), .B(n31604), .Z(n31606) );
  IV U44559 ( .A(n31606), .Z(n33902) );
  NOR U44560 ( .A(n31607), .B(n33902), .Z(n37305) );
  IV U44561 ( .A(n31608), .Z(n33887) );
  IV U44562 ( .A(n31609), .Z(n33884) );
  IV U44563 ( .A(n31610), .Z(n31612) );
  NOR U44564 ( .A(n31612), .B(n31611), .Z(n34836) );
  IV U44565 ( .A(n31613), .Z(n31615) );
  NOR U44566 ( .A(n31615), .B(n31614), .Z(n34850) );
  IV U44567 ( .A(n31616), .Z(n31621) );
  IV U44568 ( .A(n31617), .Z(n31618) );
  NOR U44569 ( .A(n31621), .B(n31618), .Z(n34860) );
  IV U44570 ( .A(n31619), .Z(n31620) );
  NOR U44571 ( .A(n31621), .B(n31620), .Z(n37260) );
  IV U44572 ( .A(n31622), .Z(n31623) );
  NOR U44573 ( .A(n31623), .B(n31625), .Z(n37257) );
  NOR U44574 ( .A(n37260), .B(n37257), .Z(n33860) );
  IV U44575 ( .A(n31624), .Z(n31626) );
  NOR U44576 ( .A(n31626), .B(n31625), .Z(n37254) );
  IV U44577 ( .A(n31627), .Z(n31630) );
  NOR U44578 ( .A(n31628), .B(n31633), .Z(n31629) );
  IV U44579 ( .A(n31629), .Z(n33853) );
  NOR U44580 ( .A(n31630), .B(n33853), .Z(n31631) );
  IV U44581 ( .A(n31631), .Z(n37252) );
  IV U44582 ( .A(n31632), .Z(n31634) );
  NOR U44583 ( .A(n31634), .B(n31633), .Z(n31635) );
  IV U44584 ( .A(n31635), .Z(n33855) );
  IV U44585 ( .A(n31636), .Z(n31637) );
  NOR U44586 ( .A(n31638), .B(n31637), .Z(n34868) );
  NOR U44587 ( .A(n31640), .B(n31639), .Z(n31641) );
  IV U44588 ( .A(n31641), .Z(n31642) );
  NOR U44589 ( .A(n31642), .B(n34876), .Z(n37240) );
  IV U44590 ( .A(n31643), .Z(n31647) );
  IV U44591 ( .A(n31644), .Z(n33844) );
  NOR U44592 ( .A(n31645), .B(n33844), .Z(n31646) );
  IV U44593 ( .A(n31646), .Z(n31649) );
  NOR U44594 ( .A(n31647), .B(n31649), .Z(n34880) );
  IV U44595 ( .A(n31648), .Z(n31650) );
  NOR U44596 ( .A(n31650), .B(n31649), .Z(n34877) );
  IV U44597 ( .A(n31651), .Z(n33837) );
  IV U44598 ( .A(n31652), .Z(n31653) );
  NOR U44599 ( .A(n33837), .B(n31653), .Z(n34884) );
  IV U44600 ( .A(n31654), .Z(n31656) );
  NOR U44601 ( .A(n31656), .B(n31655), .Z(n37224) );
  IV U44602 ( .A(n31657), .Z(n31658) );
  NOR U44603 ( .A(n31658), .B(n33840), .Z(n37230) );
  NOR U44604 ( .A(n37224), .B(n37230), .Z(n33834) );
  NOR U44605 ( .A(n31659), .B(n33824), .Z(n33822) );
  IV U44606 ( .A(n31660), .Z(n31661) );
  NOR U44607 ( .A(n31662), .B(n31661), .Z(n34893) );
  IV U44608 ( .A(n31663), .Z(n31664) );
  NOR U44609 ( .A(n31665), .B(n31664), .Z(n34890) );
  IV U44610 ( .A(n31666), .Z(n31667) );
  NOR U44611 ( .A(n31667), .B(n31674), .Z(n31668) );
  IV U44612 ( .A(n31668), .Z(n34919) );
  IV U44613 ( .A(n31669), .Z(n33799) );
  IV U44614 ( .A(n31670), .Z(n31671) );
  NOR U44615 ( .A(n33799), .B(n31671), .Z(n37206) );
  IV U44616 ( .A(n31672), .Z(n31673) );
  NOR U44617 ( .A(n31674), .B(n31673), .Z(n37210) );
  NOR U44618 ( .A(n37206), .B(n37210), .Z(n33802) );
  IV U44619 ( .A(n31675), .Z(n31676) );
  NOR U44620 ( .A(n31676), .B(n34933), .Z(n33795) );
  IV U44621 ( .A(n31677), .Z(n31678) );
  NOR U44622 ( .A(n31678), .B(n33791), .Z(n34947) );
  IV U44623 ( .A(n31679), .Z(n31680) );
  NOR U44624 ( .A(n31680), .B(n34933), .Z(n34943) );
  NOR U44625 ( .A(n34947), .B(n34943), .Z(n33794) );
  IV U44626 ( .A(n31681), .Z(n31684) );
  NOR U44627 ( .A(n33768), .B(n34964), .Z(n31682) );
  IV U44628 ( .A(n31682), .Z(n31683) );
  NOR U44629 ( .A(n31684), .B(n31683), .Z(n34959) );
  IV U44630 ( .A(n31685), .Z(n31689) );
  IV U44631 ( .A(n31686), .Z(n33761) );
  NOR U44632 ( .A(n33766), .B(n33761), .Z(n31687) );
  IV U44633 ( .A(n31687), .Z(n31688) );
  NOR U44634 ( .A(n31689), .B(n31688), .Z(n34967) );
  IV U44635 ( .A(n31690), .Z(n31691) );
  NOR U44636 ( .A(n31691), .B(n34982), .Z(n33757) );
  IV U44637 ( .A(n31692), .Z(n31696) );
  NOR U44638 ( .A(n31694), .B(n31693), .Z(n31695) );
  IV U44639 ( .A(n31695), .Z(n31698) );
  NOR U44640 ( .A(n31696), .B(n31698), .Z(n37182) );
  IV U44641 ( .A(n31697), .Z(n31699) );
  NOR U44642 ( .A(n31699), .B(n31698), .Z(n37175) );
  IV U44643 ( .A(n31700), .Z(n31702) );
  NOR U44644 ( .A(n31702), .B(n31701), .Z(n37167) );
  NOR U44645 ( .A(n34996), .B(n37167), .Z(n33754) );
  IV U44646 ( .A(n31703), .Z(n31707) );
  NOR U44647 ( .A(n31705), .B(n31704), .Z(n31706) );
  IV U44648 ( .A(n31706), .Z(n31709) );
  NOR U44649 ( .A(n31707), .B(n31709), .Z(n35001) );
  IV U44650 ( .A(n31708), .Z(n31710) );
  NOR U44651 ( .A(n31710), .B(n31709), .Z(n34998) );
  IV U44652 ( .A(n31711), .Z(n31714) );
  IV U44653 ( .A(n31712), .Z(n31716) );
  XOR U44654 ( .A(n31716), .B(n31715), .Z(n31713) );
  NOR U44655 ( .A(n31714), .B(n31713), .Z(n35006) );
  NOR U44656 ( .A(n37160), .B(n35006), .Z(n33752) );
  IV U44657 ( .A(n31715), .Z(n33747) );
  NOR U44658 ( .A(n33747), .B(n31716), .Z(n37152) );
  IV U44659 ( .A(n31717), .Z(n31718) );
  NOR U44660 ( .A(n31718), .B(n33743), .Z(n35012) );
  IV U44661 ( .A(n31719), .Z(n31720) );
  NOR U44662 ( .A(n31720), .B(n33743), .Z(n35015) );
  IV U44663 ( .A(n31721), .Z(n31722) );
  NOR U44664 ( .A(n31723), .B(n31722), .Z(n37146) );
  IV U44665 ( .A(n31724), .Z(n31726) );
  IV U44666 ( .A(n31725), .Z(n31729) );
  NOR U44667 ( .A(n31726), .B(n31729), .Z(n37143) );
  IV U44668 ( .A(n31727), .Z(n31728) );
  NOR U44669 ( .A(n31729), .B(n31728), .Z(n35018) );
  NOR U44670 ( .A(n37139), .B(n35018), .Z(n33740) );
  IV U44671 ( .A(n31730), .Z(n31731) );
  NOR U44672 ( .A(n31732), .B(n31731), .Z(n35070) );
  IV U44673 ( .A(n31733), .Z(n31735) );
  NOR U44674 ( .A(n31735), .B(n31734), .Z(n35068) );
  NOR U44675 ( .A(n35070), .B(n35068), .Z(n33680) );
  NOR U44676 ( .A(n31737), .B(n31736), .Z(n33679) );
  IV U44677 ( .A(n31738), .Z(n31741) );
  NOR U44678 ( .A(n37073), .B(n31739), .Z(n31740) );
  IV U44679 ( .A(n31740), .Z(n31743) );
  NOR U44680 ( .A(n31741), .B(n31743), .Z(n35083) );
  IV U44681 ( .A(n31742), .Z(n31744) );
  NOR U44682 ( .A(n31744), .B(n31743), .Z(n35080) );
  IV U44683 ( .A(n31745), .Z(n31746) );
  NOR U44684 ( .A(n37073), .B(n31746), .Z(n33678) );
  IV U44685 ( .A(n31747), .Z(n31750) );
  NOR U44686 ( .A(n31748), .B(n33666), .Z(n31749) );
  IV U44687 ( .A(n31749), .Z(n33676) );
  NOR U44688 ( .A(n31750), .B(n33676), .Z(n37068) );
  XOR U44689 ( .A(n33649), .B(n33648), .Z(n31751) );
  NOR U44690 ( .A(n31752), .B(n31751), .Z(n33652) );
  IV U44691 ( .A(n33652), .Z(n33647) );
  NOR U44692 ( .A(n31753), .B(n35105), .Z(n31754) );
  NOR U44693 ( .A(n31754), .B(n35106), .Z(n33646) );
  IV U44694 ( .A(n31755), .Z(n31758) );
  NOR U44695 ( .A(n31756), .B(n33637), .Z(n31757) );
  IV U44696 ( .A(n31757), .Z(n33644) );
  NOR U44697 ( .A(n31758), .B(n33644), .Z(n35102) );
  IV U44698 ( .A(n31759), .Z(n33638) );
  IV U44699 ( .A(n31760), .Z(n31761) );
  NOR U44700 ( .A(n31761), .B(n33634), .Z(n31762) );
  IV U44701 ( .A(n31762), .Z(n35114) );
  IV U44702 ( .A(n31763), .Z(n31764) );
  NOR U44703 ( .A(n31764), .B(n33634), .Z(n35110) );
  IV U44704 ( .A(n31765), .Z(n31767) );
  NOR U44705 ( .A(n31767), .B(n31766), .Z(n31768) );
  IV U44706 ( .A(n31768), .Z(n33627) );
  NOR U44707 ( .A(n35125), .B(n31769), .Z(n35118) );
  IV U44708 ( .A(n31770), .Z(n31771) );
  NOR U44709 ( .A(n31772), .B(n31771), .Z(n35115) );
  NOR U44710 ( .A(n35118), .B(n35115), .Z(n33612) );
  IV U44711 ( .A(n31773), .Z(n31777) );
  IV U44712 ( .A(n31774), .Z(n31781) );
  NOR U44713 ( .A(n31775), .B(n31781), .Z(n31776) );
  IV U44714 ( .A(n31776), .Z(n31779) );
  NOR U44715 ( .A(n31777), .B(n31779), .Z(n37032) );
  IV U44716 ( .A(n31778), .Z(n31780) );
  NOR U44717 ( .A(n31780), .B(n31779), .Z(n37029) );
  NOR U44718 ( .A(n31782), .B(n31781), .Z(n31783) );
  IV U44719 ( .A(n31783), .Z(n35135) );
  NOR U44720 ( .A(n35135), .B(n31784), .Z(n33611) );
  IV U44721 ( .A(n31785), .Z(n31788) );
  NOR U44722 ( .A(n33601), .B(n31786), .Z(n31787) );
  IV U44723 ( .A(n31787), .Z(n33596) );
  NOR U44724 ( .A(n31788), .B(n33596), .Z(n35131) );
  IV U44725 ( .A(n31789), .Z(n31794) );
  IV U44726 ( .A(n31790), .Z(n31791) );
  NOR U44727 ( .A(n31792), .B(n31791), .Z(n31793) );
  IV U44728 ( .A(n31793), .Z(n31796) );
  NOR U44729 ( .A(n31794), .B(n31796), .Z(n37012) );
  IV U44730 ( .A(n31795), .Z(n31797) );
  NOR U44731 ( .A(n31797), .B(n31796), .Z(n37008) );
  IV U44732 ( .A(n31798), .Z(n31799) );
  NOR U44733 ( .A(n33575), .B(n31799), .Z(n37004) );
  NOR U44734 ( .A(n31801), .B(n31800), .Z(n36986) );
  NOR U44735 ( .A(n36984), .B(n36986), .Z(n33569) );
  IV U44736 ( .A(n31802), .Z(n31803) );
  NOR U44737 ( .A(n31803), .B(n35155), .Z(n33567) );
  NOR U44738 ( .A(n35155), .B(n31804), .Z(n35161) );
  NOR U44739 ( .A(n35169), .B(n35161), .Z(n33566) );
  NOR U44740 ( .A(n31806), .B(n31805), .Z(n35172) );
  IV U44741 ( .A(n31807), .Z(n33560) );
  IV U44742 ( .A(n31808), .Z(n31809) );
  NOR U44743 ( .A(n33560), .B(n31809), .Z(n36974) );
  IV U44744 ( .A(n31810), .Z(n31812) );
  IV U44745 ( .A(n31811), .Z(n31818) );
  NOR U44746 ( .A(n31812), .B(n31818), .Z(n41950) );
  IV U44747 ( .A(n33543), .Z(n31816) );
  NOR U44748 ( .A(n33547), .B(n31813), .Z(n31814) );
  IV U44749 ( .A(n31814), .Z(n31815) );
  NOR U44750 ( .A(n31816), .B(n31815), .Z(n41942) );
  NOR U44751 ( .A(n41950), .B(n41942), .Z(n35183) );
  IV U44752 ( .A(n31817), .Z(n31819) );
  NOR U44753 ( .A(n31819), .B(n31818), .Z(n35190) );
  IV U44754 ( .A(n31820), .Z(n31821) );
  NOR U44755 ( .A(n31821), .B(n31824), .Z(n35187) );
  IV U44756 ( .A(n31822), .Z(n31823) );
  NOR U44757 ( .A(n31824), .B(n31823), .Z(n36952) );
  IV U44758 ( .A(n31825), .Z(n31830) );
  IV U44759 ( .A(n31826), .Z(n31827) );
  NOR U44760 ( .A(n31830), .B(n31827), .Z(n36935) );
  IV U44761 ( .A(n31828), .Z(n31829) );
  NOR U44762 ( .A(n31830), .B(n31829), .Z(n35193) );
  IV U44763 ( .A(n31831), .Z(n31832) );
  NOR U44764 ( .A(n33537), .B(n31832), .Z(n36939) );
  IV U44765 ( .A(n31833), .Z(n31836) );
  NOR U44766 ( .A(n31834), .B(n33523), .Z(n31835) );
  IV U44767 ( .A(n31835), .Z(n33507) );
  NOR U44768 ( .A(n31836), .B(n33507), .Z(n31837) );
  IV U44769 ( .A(n31837), .Z(n35201) );
  IV U44770 ( .A(n31838), .Z(n33511) );
  IV U44771 ( .A(n31839), .Z(n31840) );
  NOR U44772 ( .A(n33511), .B(n31840), .Z(n36914) );
  IV U44773 ( .A(n31841), .Z(n31844) );
  NOR U44774 ( .A(n31842), .B(n33499), .Z(n31843) );
  IV U44775 ( .A(n31843), .Z(n31846) );
  NOR U44776 ( .A(n31844), .B(n31846), .Z(n35208) );
  IV U44777 ( .A(n31845), .Z(n31847) );
  NOR U44778 ( .A(n31847), .B(n31846), .Z(n35211) );
  IV U44779 ( .A(n31848), .Z(n31851) );
  NOR U44780 ( .A(n31849), .B(n33499), .Z(n31850) );
  IV U44781 ( .A(n31850), .Z(n31853) );
  NOR U44782 ( .A(n31851), .B(n31853), .Z(n36910) );
  NOR U44783 ( .A(n35211), .B(n36910), .Z(n33496) );
  IV U44784 ( .A(n31852), .Z(n31854) );
  NOR U44785 ( .A(n31854), .B(n31853), .Z(n36906) );
  IV U44786 ( .A(n31855), .Z(n31860) );
  NOR U44787 ( .A(n31857), .B(n31856), .Z(n31858) );
  IV U44788 ( .A(n31858), .Z(n31859) );
  NOR U44789 ( .A(n31860), .B(n31859), .Z(n36903) );
  IV U44790 ( .A(n31861), .Z(n35220) );
  IV U44791 ( .A(n31862), .Z(n31863) );
  NOR U44792 ( .A(n35220), .B(n31863), .Z(n36893) );
  IV U44793 ( .A(n31864), .Z(n31865) );
  NOR U44794 ( .A(n31866), .B(n31865), .Z(n36896) );
  NOR U44795 ( .A(n36890), .B(n36896), .Z(n33480) );
  NOR U44796 ( .A(n31868), .B(n31867), .Z(n31869) );
  IV U44797 ( .A(n31869), .Z(n31870) );
  NOR U44798 ( .A(n31871), .B(n31870), .Z(n36887) );
  IV U44799 ( .A(n33475), .Z(n31875) );
  IV U44800 ( .A(n31872), .Z(n33476) );
  NOR U44801 ( .A(n31875), .B(n33476), .Z(n35229) );
  IV U44802 ( .A(n31873), .Z(n31874) );
  NOR U44803 ( .A(n31875), .B(n31874), .Z(n35224) );
  NOR U44804 ( .A(n35229), .B(n35224), .Z(n33470) );
  NOR U44805 ( .A(n31877), .B(n31876), .Z(n31878) );
  IV U44806 ( .A(n31878), .Z(n36875) );
  NOR U44807 ( .A(n36875), .B(n31879), .Z(n33469) );
  IV U44808 ( .A(n33458), .Z(n31883) );
  NOR U44809 ( .A(n31880), .B(n33460), .Z(n31881) );
  IV U44810 ( .A(n31881), .Z(n31882) );
  NOR U44811 ( .A(n31883), .B(n31882), .Z(n35237) );
  IV U44812 ( .A(n31884), .Z(n31885) );
  NOR U44813 ( .A(n31886), .B(n31885), .Z(n36859) );
  NOR U44814 ( .A(n35240), .B(n36859), .Z(n33453) );
  NOR U44815 ( .A(n31888), .B(n31887), .Z(n33451) );
  IV U44816 ( .A(n33451), .Z(n33437) );
  IV U44817 ( .A(n31889), .Z(n31890) );
  NOR U44818 ( .A(n31891), .B(n31890), .Z(n31892) );
  IV U44819 ( .A(n31892), .Z(n36850) );
  IV U44820 ( .A(n31893), .Z(n31896) );
  NOR U44821 ( .A(n31894), .B(n31900), .Z(n31895) );
  IV U44822 ( .A(n31895), .Z(n33432) );
  NOR U44823 ( .A(n31896), .B(n33432), .Z(n35246) );
  NOR U44824 ( .A(n31898), .B(n31897), .Z(n31902) );
  IV U44825 ( .A(n31899), .Z(n31901) );
  NOR U44826 ( .A(n31901), .B(n31900), .Z(n36835) );
  NOR U44827 ( .A(n31902), .B(n36835), .Z(n33426) );
  IV U44828 ( .A(n31903), .Z(n31908) );
  NOR U44829 ( .A(n31905), .B(n31904), .Z(n31906) );
  IV U44830 ( .A(n31906), .Z(n31907) );
  NOR U44831 ( .A(n31908), .B(n31907), .Z(n35256) );
  IV U44832 ( .A(n31909), .Z(n31912) );
  NOR U44833 ( .A(n31910), .B(n31918), .Z(n31911) );
  IV U44834 ( .A(n31911), .Z(n31914) );
  NOR U44835 ( .A(n31912), .B(n31914), .Z(n36820) );
  IV U44836 ( .A(n31913), .Z(n31915) );
  NOR U44837 ( .A(n31915), .B(n31914), .Z(n33413) );
  IV U44838 ( .A(n31916), .Z(n31917) );
  NOR U44839 ( .A(n31918), .B(n31917), .Z(n33410) );
  IV U44840 ( .A(n33410), .Z(n33404) );
  IV U44841 ( .A(n31919), .Z(n31922) );
  NOR U44842 ( .A(n31920), .B(n31927), .Z(n31921) );
  IV U44843 ( .A(n31921), .Z(n31924) );
  NOR U44844 ( .A(n31922), .B(n31924), .Z(n36811) );
  IV U44845 ( .A(n31923), .Z(n31925) );
  NOR U44846 ( .A(n31925), .B(n31924), .Z(n35272) );
  IV U44847 ( .A(n31926), .Z(n31928) );
  NOR U44848 ( .A(n31928), .B(n31927), .Z(n35275) );
  IV U44849 ( .A(n31929), .Z(n31936) );
  IV U44850 ( .A(n31930), .Z(n31931) );
  NOR U44851 ( .A(n31936), .B(n31931), .Z(n36807) );
  NOR U44852 ( .A(n35275), .B(n36807), .Z(n33391) );
  IV U44853 ( .A(n31932), .Z(n31933) );
  NOR U44854 ( .A(n31936), .B(n31933), .Z(n36802) );
  IV U44855 ( .A(n31934), .Z(n31935) );
  NOR U44856 ( .A(n31936), .B(n31935), .Z(n36800) );
  NOR U44857 ( .A(n31938), .B(n31937), .Z(n31939) );
  IV U44858 ( .A(n31939), .Z(n35280) );
  NOR U44859 ( .A(n35280), .B(n31940), .Z(n33390) );
  IV U44860 ( .A(n31941), .Z(n31942) );
  NOR U44861 ( .A(n31942), .B(n35285), .Z(n33389) );
  IV U44862 ( .A(n31943), .Z(n31944) );
  NOR U44863 ( .A(n35285), .B(n31944), .Z(n31945) );
  IV U44864 ( .A(n31945), .Z(n33383) );
  IV U44865 ( .A(n31946), .Z(n31950) );
  NOR U44866 ( .A(n31948), .B(n31947), .Z(n31949) );
  IV U44867 ( .A(n31949), .Z(n33381) );
  NOR U44868 ( .A(n31950), .B(n33381), .Z(n36783) );
  IV U44869 ( .A(n31951), .Z(n31952) );
  NOR U44870 ( .A(n31952), .B(n35296), .Z(n33375) );
  IV U44871 ( .A(n31953), .Z(n31954) );
  NOR U44872 ( .A(n35296), .B(n31954), .Z(n35303) );
  IV U44873 ( .A(n31955), .Z(n33373) );
  IV U44874 ( .A(n31956), .Z(n31957) );
  NOR U44875 ( .A(n33373), .B(n31957), .Z(n36760) );
  IV U44876 ( .A(n31958), .Z(n31961) );
  NOR U44877 ( .A(n31967), .B(n31959), .Z(n31960) );
  IV U44878 ( .A(n31960), .Z(n31963) );
  NOR U44879 ( .A(n31961), .B(n31963), .Z(n36764) );
  IV U44880 ( .A(n31962), .Z(n31964) );
  NOR U44881 ( .A(n31964), .B(n31963), .Z(n35311) );
  IV U44882 ( .A(n31965), .Z(n31966) );
  NOR U44883 ( .A(n31967), .B(n31966), .Z(n35313) );
  NOR U44884 ( .A(n35311), .B(n35313), .Z(n33364) );
  IV U44885 ( .A(n31968), .Z(n31969) );
  NOR U44886 ( .A(n31969), .B(n31971), .Z(n36756) );
  IV U44887 ( .A(n31970), .Z(n31972) );
  NOR U44888 ( .A(n31972), .B(n31971), .Z(n36753) );
  IV U44889 ( .A(n31973), .Z(n31974) );
  NOR U44890 ( .A(n31974), .B(n35319), .Z(n36740) );
  IV U44891 ( .A(n31975), .Z(n31984) );
  NOR U44892 ( .A(n31976), .B(n31984), .Z(n31977) );
  IV U44893 ( .A(n31977), .Z(n35327) );
  NOR U44894 ( .A(n31978), .B(n35327), .Z(n31982) );
  IV U44895 ( .A(n31979), .Z(n31980) );
  NOR U44896 ( .A(n31980), .B(n35319), .Z(n31981) );
  NOR U44897 ( .A(n31982), .B(n31981), .Z(n33354) );
  IV U44898 ( .A(n31983), .Z(n31985) );
  NOR U44899 ( .A(n31985), .B(n31984), .Z(n33352) );
  IV U44900 ( .A(n33352), .Z(n33341) );
  IV U44901 ( .A(n31986), .Z(n31987) );
  NOR U44902 ( .A(n31988), .B(n31987), .Z(n35346) );
  NOR U44903 ( .A(n35349), .B(n35346), .Z(n33339) );
  NOR U44904 ( .A(n31990), .B(n31989), .Z(n35352) );
  IV U44905 ( .A(n31991), .Z(n31993) );
  NOR U44906 ( .A(n31993), .B(n31992), .Z(n35354) );
  NOR U44907 ( .A(n35352), .B(n35354), .Z(n33338) );
  IV U44908 ( .A(n31994), .Z(n31996) );
  NOR U44909 ( .A(n31996), .B(n31995), .Z(n31997) );
  IV U44910 ( .A(n31997), .Z(n33334) );
  IV U44911 ( .A(n31998), .Z(n32001) );
  NOR U44912 ( .A(n31999), .B(n32007), .Z(n32000) );
  IV U44913 ( .A(n32000), .Z(n32003) );
  NOR U44914 ( .A(n32001), .B(n32003), .Z(n36722) );
  IV U44915 ( .A(n32002), .Z(n32004) );
  NOR U44916 ( .A(n32004), .B(n32003), .Z(n36719) );
  IV U44917 ( .A(n32005), .Z(n32006) );
  NOR U44918 ( .A(n32007), .B(n32006), .Z(n36715) );
  NOR U44919 ( .A(n36712), .B(n36715), .Z(n33328) );
  NOR U44920 ( .A(n32009), .B(n32008), .Z(n33327) );
  IV U44921 ( .A(n33327), .Z(n33322) );
  NOR U44922 ( .A(n36701), .B(n32010), .Z(n33321) );
  NOR U44923 ( .A(n33317), .B(n32011), .Z(n36696) );
  IV U44924 ( .A(n32012), .Z(n32015) );
  NOR U44925 ( .A(n32013), .B(n32017), .Z(n32014) );
  IV U44926 ( .A(n32014), .Z(n33314) );
  NOR U44927 ( .A(n32015), .B(n33314), .Z(n35359) );
  IV U44928 ( .A(n32016), .Z(n32018) );
  NOR U44929 ( .A(n32018), .B(n32017), .Z(n36679) );
  IV U44930 ( .A(n32019), .Z(n32020) );
  NOR U44931 ( .A(n32021), .B(n32020), .Z(n36674) );
  IV U44932 ( .A(n32022), .Z(n36669) );
  IV U44933 ( .A(n32023), .Z(n32024) );
  NOR U44934 ( .A(n36669), .B(n32024), .Z(n35365) );
  NOR U44935 ( .A(n36674), .B(n35365), .Z(n33309) );
  IV U44936 ( .A(n32025), .Z(n32026) );
  NOR U44937 ( .A(n32029), .B(n32026), .Z(n38782) );
  IV U44938 ( .A(n32027), .Z(n32028) );
  NOR U44939 ( .A(n32029), .B(n32028), .Z(n39989) );
  NOR U44940 ( .A(n38782), .B(n39989), .Z(n35367) );
  IV U44941 ( .A(n32030), .Z(n32031) );
  NOR U44942 ( .A(n32031), .B(n33292), .Z(n36647) );
  IV U44943 ( .A(n32032), .Z(n32036) );
  IV U44944 ( .A(n32033), .Z(n35372) );
  NOR U44945 ( .A(n35372), .B(n32034), .Z(n32035) );
  IV U44946 ( .A(n32035), .Z(n32042) );
  NOR U44947 ( .A(n32036), .B(n32042), .Z(n36636) );
  IV U44948 ( .A(n32037), .Z(n32038) );
  NOR U44949 ( .A(n32038), .B(n32045), .Z(n32039) );
  IV U44950 ( .A(n32039), .Z(n32040) );
  NOR U44951 ( .A(n32040), .B(n32048), .Z(n35378) );
  IV U44952 ( .A(n32041), .Z(n32043) );
  NOR U44953 ( .A(n32043), .B(n32042), .Z(n36633) );
  NOR U44954 ( .A(n35378), .B(n36633), .Z(n33285) );
  IV U44955 ( .A(n32044), .Z(n32046) );
  NOR U44956 ( .A(n32046), .B(n32045), .Z(n32047) );
  IV U44957 ( .A(n32047), .Z(n32049) );
  NOR U44958 ( .A(n32049), .B(n32048), .Z(n36628) );
  IV U44959 ( .A(n32050), .Z(n32055) );
  IV U44960 ( .A(n32051), .Z(n33268) );
  XOR U44961 ( .A(n33269), .B(n33268), .Z(n32053) );
  NOR U44962 ( .A(n32053), .B(n32052), .Z(n32054) );
  IV U44963 ( .A(n32054), .Z(n32057) );
  NOR U44964 ( .A(n32055), .B(n32057), .Z(n36625) );
  IV U44965 ( .A(n32056), .Z(n32058) );
  NOR U44966 ( .A(n32058), .B(n32057), .Z(n32059) );
  IV U44967 ( .A(n32059), .Z(n35382) );
  IV U44968 ( .A(n32060), .Z(n32061) );
  NOR U44969 ( .A(n32061), .B(n33268), .Z(n33266) );
  IV U44970 ( .A(n33254), .Z(n33245) );
  NOR U44971 ( .A(n32063), .B(n32062), .Z(n38819) );
  IV U44972 ( .A(n32064), .Z(n32067) );
  NOR U44973 ( .A(n32065), .B(n32071), .Z(n32066) );
  IV U44974 ( .A(n32066), .Z(n33247) );
  NOR U44975 ( .A(n32067), .B(n33247), .Z(n38813) );
  NOR U44976 ( .A(n38819), .B(n38813), .Z(n36617) );
  IV U44977 ( .A(n32068), .Z(n32069) );
  NOR U44978 ( .A(n32070), .B(n32069), .Z(n38826) );
  NOR U44979 ( .A(n32072), .B(n32071), .Z(n38822) );
  NOR U44980 ( .A(n38826), .B(n38822), .Z(n36616) );
  IV U44981 ( .A(n32073), .Z(n32075) );
  NOR U44982 ( .A(n33241), .B(n35394), .Z(n32074) );
  IV U44983 ( .A(n32074), .Z(n32077) );
  NOR U44984 ( .A(n32075), .B(n32077), .Z(n36612) );
  IV U44985 ( .A(n32076), .Z(n32078) );
  NOR U44986 ( .A(n32078), .B(n32077), .Z(n32079) );
  IV U44987 ( .A(n32079), .Z(n36611) );
  IV U44988 ( .A(n32080), .Z(n32083) );
  IV U44989 ( .A(n32081), .Z(n32082) );
  NOR U44990 ( .A(n32083), .B(n32082), .Z(n35397) );
  IV U44991 ( .A(n32084), .Z(n32085) );
  NOR U44992 ( .A(n32085), .B(n33233), .Z(n36607) );
  NOR U44993 ( .A(n35397), .B(n36607), .Z(n42229) );
  IV U44994 ( .A(n32086), .Z(n33237) );
  IV U44995 ( .A(n32087), .Z(n32088) );
  NOR U44996 ( .A(n33237), .B(n32088), .Z(n35405) );
  IV U44997 ( .A(n32089), .Z(n32090) );
  NOR U44998 ( .A(n33230), .B(n32090), .Z(n35402) );
  IV U44999 ( .A(n32091), .Z(n32094) );
  NOR U45000 ( .A(n32092), .B(n32097), .Z(n32093) );
  IV U45001 ( .A(n32093), .Z(n32099) );
  NOR U45002 ( .A(n32094), .B(n32099), .Z(n36596) );
  IV U45003 ( .A(n32095), .Z(n32096) );
  NOR U45004 ( .A(n32097), .B(n32096), .Z(n36590) );
  IV U45005 ( .A(n32098), .Z(n32100) );
  NOR U45006 ( .A(n32100), .B(n32099), .Z(n36599) );
  NOR U45007 ( .A(n36590), .B(n36599), .Z(n33227) );
  IV U45008 ( .A(n32101), .Z(n32102) );
  NOR U45009 ( .A(n32102), .B(n32105), .Z(n36581) );
  IV U45010 ( .A(n32103), .Z(n32104) );
  NOR U45011 ( .A(n32105), .B(n32104), .Z(n36592) );
  NOR U45012 ( .A(n36581), .B(n36592), .Z(n33226) );
  IV U45013 ( .A(n32108), .Z(n32106) );
  NOR U45014 ( .A(n32107), .B(n32106), .Z(n35412) );
  NOR U45015 ( .A(n36576), .B(n36583), .Z(n32111) );
  NOR U45016 ( .A(n32109), .B(n32108), .Z(n32110) );
  NOR U45017 ( .A(n32111), .B(n32110), .Z(n32112) );
  NOR U45018 ( .A(n35412), .B(n32112), .Z(n33225) );
  NOR U45019 ( .A(n32113), .B(n35416), .Z(n33224) );
  IV U45020 ( .A(n32114), .Z(n32115) );
  NOR U45021 ( .A(n35416), .B(n32115), .Z(n33219) );
  IV U45022 ( .A(n33219), .Z(n33212) );
  IV U45023 ( .A(n32116), .Z(n32118) );
  NOR U45024 ( .A(n32118), .B(n32117), .Z(n35425) );
  IV U45025 ( .A(n32119), .Z(n32120) );
  NOR U45026 ( .A(n32121), .B(n32120), .Z(n39900) );
  IV U45027 ( .A(n32122), .Z(n32123) );
  NOR U45028 ( .A(n32123), .B(n32125), .Z(n38852) );
  NOR U45029 ( .A(n39900), .B(n38852), .Z(n35424) );
  IV U45030 ( .A(n32124), .Z(n32126) );
  NOR U45031 ( .A(n32126), .B(n32125), .Z(n35429) );
  IV U45032 ( .A(n32127), .Z(n32130) );
  NOR U45033 ( .A(n32128), .B(n33206), .Z(n32129) );
  IV U45034 ( .A(n32129), .Z(n33209) );
  NOR U45035 ( .A(n32130), .B(n33209), .Z(n35434) );
  NOR U45036 ( .A(n35429), .B(n35434), .Z(n33211) );
  IV U45037 ( .A(n32131), .Z(n33193) );
  NOR U45038 ( .A(n32132), .B(n33193), .Z(n33191) );
  IV U45039 ( .A(n32133), .Z(n32137) );
  NOR U45040 ( .A(n32135), .B(n32134), .Z(n32136) );
  IV U45041 ( .A(n32136), .Z(n33183) );
  NOR U45042 ( .A(n32137), .B(n33183), .Z(n36560) );
  IV U45043 ( .A(n32138), .Z(n32140) );
  IV U45044 ( .A(n32139), .Z(n33178) );
  NOR U45045 ( .A(n32140), .B(n33178), .Z(n35448) );
  IV U45046 ( .A(n32141), .Z(n32142) );
  NOR U45047 ( .A(n32144), .B(n32142), .Z(n36551) );
  IV U45048 ( .A(n32143), .Z(n35455) );
  NOR U45049 ( .A(n35455), .B(n32144), .Z(n32148) );
  IV U45050 ( .A(n32145), .Z(n35452) );
  IV U45051 ( .A(n32146), .Z(n32147) );
  NOR U45052 ( .A(n35452), .B(n32147), .Z(n35459) );
  NOR U45053 ( .A(n32148), .B(n35459), .Z(n33175) );
  IV U45054 ( .A(n32149), .Z(n32150) );
  NOR U45055 ( .A(n35452), .B(n32150), .Z(n35456) );
  IV U45056 ( .A(n32151), .Z(n33157) );
  NOR U45057 ( .A(n32152), .B(n33157), .Z(n35465) );
  IV U45058 ( .A(n32153), .Z(n32154) );
  NOR U45059 ( .A(n32154), .B(n33157), .Z(n35462) );
  XOR U45060 ( .A(n32155), .B(n33164), .Z(n32156) );
  NOR U45061 ( .A(n32157), .B(n32156), .Z(n32158) );
  IV U45062 ( .A(n32158), .Z(n36539) );
  IV U45063 ( .A(n32159), .Z(n32163) );
  IV U45064 ( .A(n32160), .Z(n32167) );
  NOR U45065 ( .A(n32161), .B(n32167), .Z(n32162) );
  IV U45066 ( .A(n32162), .Z(n33152) );
  NOR U45067 ( .A(n32163), .B(n33152), .Z(n36519) );
  IV U45068 ( .A(n32164), .Z(n32165) );
  NOR U45069 ( .A(n32165), .B(n33139), .Z(n35477) );
  IV U45070 ( .A(n32166), .Z(n32168) );
  NOR U45071 ( .A(n32168), .B(n32167), .Z(n36523) );
  NOR U45072 ( .A(n35477), .B(n36523), .Z(n33149) );
  IV U45073 ( .A(n32169), .Z(n32170) );
  NOR U45074 ( .A(n32171), .B(n32170), .Z(n32172) );
  IV U45075 ( .A(n32172), .Z(n33144) );
  IV U45076 ( .A(n32173), .Z(n32175) );
  IV U45077 ( .A(n32174), .Z(n33136) );
  NOR U45078 ( .A(n32175), .B(n33136), .Z(n35482) );
  NOR U45079 ( .A(n35487), .B(n35482), .Z(n33130) );
  IV U45080 ( .A(n32176), .Z(n32177) );
  NOR U45081 ( .A(n32177), .B(n33121), .Z(n32178) );
  IV U45082 ( .A(n32178), .Z(n35486) );
  NOR U45083 ( .A(n32180), .B(n32179), .Z(n33124) );
  IV U45084 ( .A(n32181), .Z(n32182) );
  NOR U45085 ( .A(n32182), .B(n32183), .Z(n36501) );
  NOR U45086 ( .A(n32184), .B(n32183), .Z(n38903) );
  IV U45087 ( .A(n32185), .Z(n32187) );
  IV U45088 ( .A(n32186), .Z(n33111) );
  NOR U45089 ( .A(n32187), .B(n33111), .Z(n38897) );
  NOR U45090 ( .A(n38903), .B(n38897), .Z(n36499) );
  IV U45091 ( .A(n32188), .Z(n32192) );
  NOR U45092 ( .A(n32190), .B(n32189), .Z(n32191) );
  IV U45093 ( .A(n32191), .Z(n32194) );
  NOR U45094 ( .A(n32192), .B(n32194), .Z(n35495) );
  IV U45095 ( .A(n32193), .Z(n32195) );
  NOR U45096 ( .A(n32195), .B(n32194), .Z(n35492) );
  IV U45097 ( .A(n32196), .Z(n35507) );
  IV U45098 ( .A(n32197), .Z(n35500) );
  NOR U45099 ( .A(n32198), .B(n35500), .Z(n32199) );
  XOR U45100 ( .A(n35507), .B(n32199), .Z(n32200) );
  NOR U45101 ( .A(n32200), .B(n35506), .Z(n33104) );
  IV U45102 ( .A(n32201), .Z(n32202) );
  NOR U45103 ( .A(n32202), .B(n33098), .Z(n35526) );
  NOR U45104 ( .A(n35531), .B(n35526), .Z(n33091) );
  IV U45105 ( .A(n32203), .Z(n36489) );
  IV U45106 ( .A(n32204), .Z(n32205) );
  NOR U45107 ( .A(n32206), .B(n32205), .Z(n36484) );
  IV U45108 ( .A(n32207), .Z(n32209) );
  NOR U45109 ( .A(n32209), .B(n32208), .Z(n35549) );
  NOR U45110 ( .A(n36484), .B(n35549), .Z(n33080) );
  NOR U45111 ( .A(n32210), .B(n33066), .Z(n33064) );
  IV U45112 ( .A(n32211), .Z(n33072) );
  NOR U45113 ( .A(n33072), .B(n33066), .Z(n32212) );
  IV U45114 ( .A(n32212), .Z(n36475) );
  IV U45115 ( .A(n32213), .Z(n35554) );
  IV U45116 ( .A(n32214), .Z(n32215) );
  NOR U45117 ( .A(n35554), .B(n32215), .Z(n32216) );
  IV U45118 ( .A(n32216), .Z(n35560) );
  IV U45119 ( .A(n32217), .Z(n32218) );
  NOR U45120 ( .A(n33052), .B(n32218), .Z(n35562) );
  IV U45121 ( .A(n32219), .Z(n32220) );
  NOR U45122 ( .A(n33050), .B(n32220), .Z(n32221) );
  IV U45123 ( .A(n32221), .Z(n32222) );
  NOR U45124 ( .A(n32222), .B(n33052), .Z(n36460) );
  NOR U45125 ( .A(n35562), .B(n36460), .Z(n33054) );
  IV U45126 ( .A(n32223), .Z(n32226) );
  NOR U45127 ( .A(n32224), .B(n32228), .Z(n32225) );
  IV U45128 ( .A(n32225), .Z(n33001) );
  NOR U45129 ( .A(n32226), .B(n33001), .Z(n36438) );
  IV U45130 ( .A(n32227), .Z(n32229) );
  NOR U45131 ( .A(n32229), .B(n32228), .Z(n36426) );
  NOR U45132 ( .A(n36438), .B(n36426), .Z(n32999) );
  IV U45133 ( .A(n32230), .Z(n32235) );
  IV U45134 ( .A(n32231), .Z(n32232) );
  NOR U45135 ( .A(n32235), .B(n32232), .Z(n36422) );
  IV U45136 ( .A(n32233), .Z(n32234) );
  NOR U45137 ( .A(n32235), .B(n32234), .Z(n36429) );
  IV U45138 ( .A(n32236), .Z(n32237) );
  NOR U45139 ( .A(n32237), .B(n32994), .Z(n36417) );
  IV U45140 ( .A(n32238), .Z(n32239) );
  NOR U45141 ( .A(n32994), .B(n32239), .Z(n32240) );
  IV U45142 ( .A(n32240), .Z(n36416) );
  IV U45143 ( .A(n32241), .Z(n32242) );
  NOR U45144 ( .A(n32244), .B(n32242), .Z(n36394) );
  IV U45145 ( .A(n32243), .Z(n32247) );
  NOR U45146 ( .A(n32245), .B(n32244), .Z(n32246) );
  IV U45147 ( .A(n32246), .Z(n32973) );
  NOR U45148 ( .A(n32247), .B(n32973), .Z(n36405) );
  NOR U45149 ( .A(n36394), .B(n36405), .Z(n32971) );
  IV U45150 ( .A(n32248), .Z(n32253) );
  IV U45151 ( .A(n32249), .Z(n32250) );
  NOR U45152 ( .A(n32253), .B(n32250), .Z(n35598) );
  IV U45153 ( .A(n32251), .Z(n32252) );
  NOR U45154 ( .A(n32253), .B(n32252), .Z(n36397) );
  IV U45155 ( .A(n32254), .Z(n32256) );
  NOR U45156 ( .A(n32256), .B(n32255), .Z(n36382) );
  IV U45157 ( .A(n32257), .Z(n32260) );
  NOR U45158 ( .A(n32258), .B(n32266), .Z(n32259) );
  IV U45159 ( .A(n32259), .Z(n32262) );
  NOR U45160 ( .A(n32260), .B(n32262), .Z(n35601) );
  IV U45161 ( .A(n32261), .Z(n32263) );
  NOR U45162 ( .A(n32263), .B(n32262), .Z(n36385) );
  IV U45163 ( .A(n32264), .Z(n32265) );
  NOR U45164 ( .A(n32266), .B(n32265), .Z(n35605) );
  NOR U45165 ( .A(n32268), .B(n32267), .Z(n35610) );
  NOR U45166 ( .A(n35614), .B(n32269), .Z(n35627) );
  IV U45167 ( .A(n32270), .Z(n32271) );
  NOR U45168 ( .A(n32272), .B(n32271), .Z(n35622) );
  NOR U45169 ( .A(n35627), .B(n35622), .Z(n32961) );
  IV U45170 ( .A(n32273), .Z(n32274) );
  NOR U45171 ( .A(n32274), .B(n32276), .Z(n36356) );
  IV U45172 ( .A(n32275), .Z(n32277) );
  NOR U45173 ( .A(n32277), .B(n32276), .Z(n36353) );
  IV U45174 ( .A(n32278), .Z(n32279) );
  NOR U45175 ( .A(n32279), .B(n32958), .Z(n36364) );
  NOR U45176 ( .A(n36353), .B(n36364), .Z(n32951) );
  IV U45177 ( .A(n35654), .Z(n35649) );
  IV U45178 ( .A(n32280), .Z(n35655) );
  NOR U45179 ( .A(n35649), .B(n35655), .Z(n35660) );
  IV U45180 ( .A(n32281), .Z(n32282) );
  NOR U45181 ( .A(n32282), .B(n32917), .Z(n32913) );
  NOR U45182 ( .A(n32284), .B(n32283), .Z(n32911) );
  IV U45183 ( .A(n32285), .Z(n32288) );
  NOR U45184 ( .A(n32286), .B(n36329), .Z(n32287) );
  IV U45185 ( .A(n32287), .Z(n32908) );
  NOR U45186 ( .A(n32288), .B(n32908), .Z(n42450) );
  NOR U45187 ( .A(n42457), .B(n42450), .Z(n36307) );
  NOR U45188 ( .A(n32290), .B(n32289), .Z(n35674) );
  NOR U45189 ( .A(n35677), .B(n35674), .Z(n32906) );
  IV U45190 ( .A(n32291), .Z(n32293) );
  NOR U45191 ( .A(n32293), .B(n32292), .Z(n36303) );
  NOR U45192 ( .A(n32295), .B(n32294), .Z(n35680) );
  NOR U45193 ( .A(n36303), .B(n35680), .Z(n32905) );
  IV U45194 ( .A(n32296), .Z(n32298) );
  NOR U45195 ( .A(n32298), .B(n32297), .Z(n35683) );
  IV U45196 ( .A(n32299), .Z(n32301) );
  NOR U45197 ( .A(n32301), .B(n32300), .Z(n36295) );
  NOR U45198 ( .A(n35686), .B(n36295), .Z(n32904) );
  IV U45199 ( .A(n32302), .Z(n32303) );
  NOR U45200 ( .A(n32303), .B(n32306), .Z(n35691) );
  NOR U45201 ( .A(n35691), .B(n35688), .Z(n32903) );
  IV U45202 ( .A(n32304), .Z(n32305) );
  NOR U45203 ( .A(n32306), .B(n32305), .Z(n32307) );
  IV U45204 ( .A(n32307), .Z(n32308) );
  NOR U45205 ( .A(n32309), .B(n32308), .Z(n35696) );
  IV U45206 ( .A(n32310), .Z(n32313) );
  NOR U45207 ( .A(n32311), .B(n32900), .Z(n32312) );
  IV U45208 ( .A(n32312), .Z(n32315) );
  NOR U45209 ( .A(n32313), .B(n32315), .Z(n35693) );
  IV U45210 ( .A(n32314), .Z(n32316) );
  NOR U45211 ( .A(n32316), .B(n32315), .Z(n35706) );
  IV U45212 ( .A(n32317), .Z(n32318) );
  NOR U45213 ( .A(n32319), .B(n32318), .Z(n35712) );
  NOR U45214 ( .A(n32321), .B(n32320), .Z(n35710) );
  NOR U45215 ( .A(n35712), .B(n35710), .Z(n32898) );
  IV U45216 ( .A(n32322), .Z(n32323) );
  NOR U45217 ( .A(n32323), .B(n32896), .Z(n36287) );
  IV U45218 ( .A(n32324), .Z(n32325) );
  NOR U45219 ( .A(n32326), .B(n32325), .Z(n32887) );
  NOR U45220 ( .A(n32328), .B(n32327), .Z(n36271) );
  IV U45221 ( .A(n32329), .Z(n32330) );
  NOR U45222 ( .A(n32330), .B(n32878), .Z(n32331) );
  IV U45223 ( .A(n32331), .Z(n32333) );
  IV U45224 ( .A(n32332), .Z(n32881) );
  NOR U45225 ( .A(n32333), .B(n32881), .Z(n36278) );
  NOR U45226 ( .A(n36271), .B(n36278), .Z(n32872) );
  IV U45227 ( .A(n32334), .Z(n32339) );
  IV U45228 ( .A(n32335), .Z(n32336) );
  NOR U45229 ( .A(n32339), .B(n32336), .Z(n35721) );
  IV U45230 ( .A(n32337), .Z(n32338) );
  NOR U45231 ( .A(n32339), .B(n32338), .Z(n36261) );
  IV U45232 ( .A(n32340), .Z(n32341) );
  NOR U45233 ( .A(n32862), .B(n32341), .Z(n35723) );
  IV U45234 ( .A(n32858), .Z(n32345) );
  NOR U45235 ( .A(n32342), .B(n32854), .Z(n32343) );
  IV U45236 ( .A(n32343), .Z(n32344) );
  NOR U45237 ( .A(n32345), .B(n32344), .Z(n35737) );
  IV U45238 ( .A(n32346), .Z(n32347) );
  NOR U45239 ( .A(n32347), .B(n32854), .Z(n32348) );
  IV U45240 ( .A(n32348), .Z(n32349) );
  NOR U45241 ( .A(n32350), .B(n32349), .Z(n35742) );
  NOR U45242 ( .A(n35737), .B(n35742), .Z(n32852) );
  IV U45243 ( .A(n32350), .Z(n32354) );
  NOR U45244 ( .A(n32351), .B(n32854), .Z(n32352) );
  IV U45245 ( .A(n32352), .Z(n32353) );
  NOR U45246 ( .A(n32354), .B(n32353), .Z(n35739) );
  IV U45247 ( .A(n32355), .Z(n35753) );
  NOR U45248 ( .A(n35753), .B(n32356), .Z(n32845) );
  NOR U45249 ( .A(n32358), .B(n32357), .Z(n32359) );
  IV U45250 ( .A(n32359), .Z(n35760) );
  NOR U45251 ( .A(n32360), .B(n35760), .Z(n35757) );
  IV U45252 ( .A(n32361), .Z(n32364) );
  NOR U45253 ( .A(n32362), .B(n32376), .Z(n32363) );
  IV U45254 ( .A(n32363), .Z(n32366) );
  NOR U45255 ( .A(n32364), .B(n32366), .Z(n35764) );
  NOR U45256 ( .A(n35757), .B(n35764), .Z(n32844) );
  IV U45257 ( .A(n32365), .Z(n32367) );
  NOR U45258 ( .A(n32367), .B(n32366), .Z(n35768) );
  IV U45259 ( .A(n32368), .Z(n32369) );
  NOR U45260 ( .A(n32369), .B(n32376), .Z(n32370) );
  IV U45261 ( .A(n32370), .Z(n32371) );
  NOR U45262 ( .A(n32375), .B(n32371), .Z(n35770) );
  NOR U45263 ( .A(n35768), .B(n35770), .Z(n32843) );
  IV U45264 ( .A(n32372), .Z(n32374) );
  NOR U45265 ( .A(n32374), .B(n32373), .Z(n36228) );
  IV U45266 ( .A(n32375), .Z(n32380) );
  NOR U45267 ( .A(n32377), .B(n32376), .Z(n32378) );
  IV U45268 ( .A(n32378), .Z(n32379) );
  NOR U45269 ( .A(n32380), .B(n32379), .Z(n36236) );
  NOR U45270 ( .A(n36228), .B(n36236), .Z(n32842) );
  IV U45271 ( .A(n32381), .Z(n36232) );
  NOR U45272 ( .A(n32383), .B(n32382), .Z(n32840) );
  IV U45273 ( .A(n32840), .Z(n32832) );
  NOR U45274 ( .A(n32385), .B(n32384), .Z(n32386) );
  IV U45275 ( .A(n32386), .Z(n36225) );
  IV U45276 ( .A(n32387), .Z(n32388) );
  NOR U45277 ( .A(n32829), .B(n32388), .Z(n32389) );
  IV U45278 ( .A(n32389), .Z(n36222) );
  IV U45279 ( .A(n32390), .Z(n32391) );
  NOR U45280 ( .A(n32393), .B(n32391), .Z(n35785) );
  IV U45281 ( .A(n32392), .Z(n32394) );
  NOR U45282 ( .A(n32394), .B(n32393), .Z(n35782) );
  IV U45283 ( .A(n32395), .Z(n32399) );
  IV U45284 ( .A(n32396), .Z(n32405) );
  NOR U45285 ( .A(n32397), .B(n32405), .Z(n32398) );
  IV U45286 ( .A(n32398), .Z(n32402) );
  NOR U45287 ( .A(n32399), .B(n32402), .Z(n32400) );
  IV U45288 ( .A(n32400), .Z(n36205) );
  IV U45289 ( .A(n32401), .Z(n32403) );
  NOR U45290 ( .A(n32403), .B(n32402), .Z(n35793) );
  IV U45291 ( .A(n32404), .Z(n32406) );
  NOR U45292 ( .A(n32406), .B(n32405), .Z(n35799) );
  IV U45293 ( .A(n32407), .Z(n32408) );
  NOR U45294 ( .A(n32408), .B(n32796), .Z(n35809) );
  IV U45295 ( .A(n32409), .Z(n32410) );
  NOR U45296 ( .A(n32411), .B(n32410), .Z(n35814) );
  IV U45297 ( .A(n32412), .Z(n32414) );
  NOR U45298 ( .A(n32414), .B(n32413), .Z(n35812) );
  NOR U45299 ( .A(n35814), .B(n35812), .Z(n32792) );
  IV U45300 ( .A(n32415), .Z(n32418) );
  IV U45301 ( .A(n32416), .Z(n32417) );
  NOR U45302 ( .A(n32418), .B(n32417), .Z(n35821) );
  IV U45303 ( .A(n32419), .Z(n32786) );
  IV U45304 ( .A(n32420), .Z(n32424) );
  NOR U45305 ( .A(n32422), .B(n32421), .Z(n32423) );
  IV U45306 ( .A(n32423), .Z(n32426) );
  NOR U45307 ( .A(n32424), .B(n32426), .Z(n35826) );
  IV U45308 ( .A(n32425), .Z(n32427) );
  NOR U45309 ( .A(n32427), .B(n32426), .Z(n35824) );
  NOR U45310 ( .A(n35826), .B(n35824), .Z(n32779) );
  IV U45311 ( .A(n32428), .Z(n32432) );
  NOR U45312 ( .A(n32430), .B(n32429), .Z(n32431) );
  IV U45313 ( .A(n32431), .Z(n32434) );
  NOR U45314 ( .A(n32432), .B(n32434), .Z(n35832) );
  IV U45315 ( .A(n32433), .Z(n32435) );
  NOR U45316 ( .A(n32435), .B(n32434), .Z(n35829) );
  IV U45317 ( .A(n32436), .Z(n32439) );
  NOR U45318 ( .A(n32437), .B(n32774), .Z(n32438) );
  IV U45319 ( .A(n32438), .Z(n32441) );
  NOR U45320 ( .A(n32439), .B(n32441), .Z(n35835) );
  IV U45321 ( .A(n32440), .Z(n32442) );
  NOR U45322 ( .A(n32442), .B(n32441), .Z(n36183) );
  IV U45323 ( .A(n32443), .Z(n32445) );
  NOR U45324 ( .A(n32445), .B(n32444), .Z(n35838) );
  NOR U45325 ( .A(n32447), .B(n32446), .Z(n35842) );
  NOR U45326 ( .A(n35845), .B(n35842), .Z(n32770) );
  NOR U45327 ( .A(n32449), .B(n32448), .Z(n32758) );
  IV U45328 ( .A(n32450), .Z(n32453) );
  NOR U45329 ( .A(n32460), .B(n32451), .Z(n32452) );
  IV U45330 ( .A(n32452), .Z(n32456) );
  NOR U45331 ( .A(n32453), .B(n32456), .Z(n32454) );
  IV U45332 ( .A(n32454), .Z(n35859) );
  IV U45333 ( .A(n32455), .Z(n32457) );
  NOR U45334 ( .A(n32457), .B(n32456), .Z(n39132) );
  IV U45335 ( .A(n32458), .Z(n32462) );
  NOR U45336 ( .A(n32460), .B(n32459), .Z(n32461) );
  IV U45337 ( .A(n32461), .Z(n32744) );
  NOR U45338 ( .A(n32462), .B(n32744), .Z(n39420) );
  NOR U45339 ( .A(n39132), .B(n39420), .Z(n36162) );
  IV U45340 ( .A(n32463), .Z(n32467) );
  NOR U45341 ( .A(n32465), .B(n32464), .Z(n32466) );
  IV U45342 ( .A(n32466), .Z(n32748) );
  NOR U45343 ( .A(n32467), .B(n32748), .Z(n36147) );
  IV U45344 ( .A(n32468), .Z(n32470) );
  IV U45345 ( .A(n32469), .Z(n32730) );
  NOR U45346 ( .A(n32470), .B(n32730), .Z(n36128) );
  NOR U45347 ( .A(n35868), .B(n36113), .Z(n32471) );
  NOR U45348 ( .A(n32471), .B(n36110), .Z(n36116) );
  IV U45349 ( .A(n32472), .Z(n32473) );
  NOR U45350 ( .A(n32474), .B(n32473), .Z(n39143) );
  IV U45351 ( .A(n32475), .Z(n32476) );
  NOR U45352 ( .A(n32476), .B(n32717), .Z(n39147) );
  NOR U45353 ( .A(n39143), .B(n39147), .Z(n36120) );
  IV U45354 ( .A(n32477), .Z(n32478) );
  NOR U45355 ( .A(n32481), .B(n32478), .Z(n36099) );
  IV U45356 ( .A(n32479), .Z(n32480) );
  NOR U45357 ( .A(n32481), .B(n32480), .Z(n35882) );
  IV U45358 ( .A(n32482), .Z(n32483) );
  NOR U45359 ( .A(n32484), .B(n32483), .Z(n36094) );
  IV U45360 ( .A(n32485), .Z(n32486) );
  NOR U45361 ( .A(n32487), .B(n32486), .Z(n35885) );
  NOR U45362 ( .A(n36094), .B(n35885), .Z(n32704) );
  IV U45363 ( .A(n32488), .Z(n32491) );
  IV U45364 ( .A(n32489), .Z(n32490) );
  NOR U45365 ( .A(n32491), .B(n32490), .Z(n36092) );
  IV U45366 ( .A(n32492), .Z(n32495) );
  NOR U45367 ( .A(n32493), .B(n32697), .Z(n32494) );
  IV U45368 ( .A(n32494), .Z(n32700) );
  NOR U45369 ( .A(n32495), .B(n32700), .Z(n35890) );
  IV U45370 ( .A(n32496), .Z(n32498) );
  NOR U45371 ( .A(n32498), .B(n32497), .Z(n32499) );
  IV U45372 ( .A(n32499), .Z(n32500) );
  NOR U45373 ( .A(n32505), .B(n32500), .Z(n35896) );
  IV U45374 ( .A(n32501), .Z(n32502) );
  NOR U45375 ( .A(n32510), .B(n32502), .Z(n39171) );
  IV U45376 ( .A(n32503), .Z(n32504) );
  NOR U45377 ( .A(n32504), .B(n32520), .Z(n39175) );
  NOR U45378 ( .A(n39171), .B(n39175), .Z(n35902) );
  IV U45379 ( .A(n35902), .Z(n32511) );
  IV U45380 ( .A(n32505), .Z(n32507) );
  NOR U45381 ( .A(n32507), .B(n32506), .Z(n32508) );
  IV U45382 ( .A(n32508), .Z(n32509) );
  NOR U45383 ( .A(n32510), .B(n32509), .Z(n35899) );
  NOR U45384 ( .A(n32511), .B(n35899), .Z(n32696) );
  IV U45385 ( .A(n32512), .Z(n32513) );
  NOR U45386 ( .A(n32518), .B(n32513), .Z(n32514) );
  IV U45387 ( .A(n32514), .Z(n32515) );
  NOR U45388 ( .A(n32515), .B(n32520), .Z(n35906) );
  IV U45389 ( .A(n32516), .Z(n32517) );
  NOR U45390 ( .A(n32518), .B(n32517), .Z(n32519) );
  IV U45391 ( .A(n32519), .Z(n32521) );
  NOR U45392 ( .A(n32521), .B(n32520), .Z(n35903) );
  IV U45393 ( .A(n32522), .Z(n32524) );
  NOR U45394 ( .A(n32524), .B(n32523), .Z(n36086) );
  NOR U45395 ( .A(n35903), .B(n36086), .Z(n32525) );
  IV U45396 ( .A(n32525), .Z(n32526) );
  NOR U45397 ( .A(n35906), .B(n32526), .Z(n32695) );
  IV U45398 ( .A(n32527), .Z(n32529) );
  IV U45399 ( .A(n32528), .Z(n32531) );
  NOR U45400 ( .A(n32529), .B(n32531), .Z(n35910) );
  IV U45401 ( .A(n32530), .Z(n32534) );
  NOR U45402 ( .A(n32532), .B(n32531), .Z(n32533) );
  IV U45403 ( .A(n32533), .Z(n32536) );
  NOR U45404 ( .A(n32534), .B(n32536), .Z(n36070) );
  IV U45405 ( .A(n32535), .Z(n32537) );
  NOR U45406 ( .A(n32537), .B(n32536), .Z(n36067) );
  NOR U45407 ( .A(n35917), .B(n36061), .Z(n32683) );
  IV U45408 ( .A(n32538), .Z(n32678) );
  IV U45409 ( .A(n32539), .Z(n32540) );
  NOR U45410 ( .A(n32667), .B(n32540), .Z(n35923) );
  IV U45411 ( .A(n32541), .Z(n32542) );
  NOR U45412 ( .A(n32545), .B(n32542), .Z(n36039) );
  IV U45413 ( .A(n32543), .Z(n32544) );
  NOR U45414 ( .A(n32545), .B(n32544), .Z(n36036) );
  IV U45415 ( .A(n32546), .Z(n32552) );
  IV U45416 ( .A(n32547), .Z(n32548) );
  NOR U45417 ( .A(n32552), .B(n32548), .Z(n36025) );
  IV U45418 ( .A(n32549), .Z(n32550) );
  NOR U45419 ( .A(n32550), .B(n32552), .Z(n36028) );
  IV U45420 ( .A(n32551), .Z(n32555) );
  NOR U45421 ( .A(n32553), .B(n32552), .Z(n32554) );
  IV U45422 ( .A(n32554), .Z(n32653) );
  NOR U45423 ( .A(n32555), .B(n32653), .Z(n36022) );
  NOR U45424 ( .A(n36028), .B(n36022), .Z(n32656) );
  IV U45425 ( .A(n32556), .Z(n32557) );
  NOR U45426 ( .A(n32564), .B(n32557), .Z(n36008) );
  IV U45427 ( .A(n32558), .Z(n32559) );
  NOR U45428 ( .A(n32559), .B(n32564), .Z(n35930) );
  IV U45429 ( .A(n32560), .Z(n32561) );
  NOR U45430 ( .A(n32562), .B(n32561), .Z(n39279) );
  IV U45431 ( .A(n32563), .Z(n32565) );
  NOR U45432 ( .A(n32565), .B(n32564), .Z(n39284) );
  NOR U45433 ( .A(n39279), .B(n39284), .Z(n36013) );
  IV U45434 ( .A(n32566), .Z(n32568) );
  NOR U45435 ( .A(n32568), .B(n32567), .Z(n35936) );
  IV U45436 ( .A(n32569), .Z(n32570) );
  NOR U45437 ( .A(n32571), .B(n32570), .Z(n35934) );
  NOR U45438 ( .A(n35936), .B(n35934), .Z(n32651) );
  IV U45439 ( .A(n32572), .Z(n32573) );
  NOR U45440 ( .A(n32574), .B(n32573), .Z(n35939) );
  NOR U45441 ( .A(n35942), .B(n35939), .Z(n32650) );
  IV U45442 ( .A(n32575), .Z(n32577) );
  NOR U45443 ( .A(n32577), .B(n32576), .Z(n36002) );
  NOR U45444 ( .A(n36004), .B(n36002), .Z(n32649) );
  IV U45445 ( .A(n32578), .Z(n32579) );
  NOR U45446 ( .A(n32579), .B(n32637), .Z(n35945) );
  XOR U45447 ( .A(n32580), .B(n32637), .Z(n32581) );
  NOR U45448 ( .A(n32582), .B(n32581), .Z(n35950) );
  NOR U45449 ( .A(n35945), .B(n35950), .Z(n32648) );
  IV U45450 ( .A(n32583), .Z(n32584) );
  NOR U45451 ( .A(n32585), .B(n32584), .Z(n32586) );
  IV U45452 ( .A(n32586), .Z(n32643) );
  IV U45453 ( .A(n32587), .Z(n32588) );
  NOR U45454 ( .A(n32588), .B(n32622), .Z(n32589) );
  IV U45455 ( .A(n32589), .Z(n32590) );
  NOR U45456 ( .A(n32590), .B(n32631), .Z(n35959) );
  IV U45457 ( .A(n32591), .Z(n32593) );
  NOR U45458 ( .A(n32593), .B(n32592), .Z(n35964) );
  IV U45459 ( .A(n32594), .Z(n32599) );
  IV U45460 ( .A(n32595), .Z(n32596) );
  NOR U45461 ( .A(n32599), .B(n32596), .Z(n35987) );
  NOR U45462 ( .A(n35964), .B(n35987), .Z(n32619) );
  IV U45463 ( .A(n32597), .Z(n32598) );
  NOR U45464 ( .A(n32599), .B(n32598), .Z(n35967) );
  IV U45465 ( .A(n32604), .Z(n32605) );
  NOR U45466 ( .A(n32605), .B(n32612), .Z(n32609) );
  NOR U45467 ( .A(n32607), .B(n32606), .Z(n32608) );
  NOR U45468 ( .A(n32609), .B(n32608), .Z(n35970) );
  XOR U45469 ( .A(n35970), .B(n35971), .Z(n35973) );
  XOR U45470 ( .A(n35974), .B(n35973), .Z(n35981) );
  IV U45471 ( .A(n32616), .Z(n32618) );
  NOR U45472 ( .A(n32618), .B(n32617), .Z(n35979) );
  XOR U45473 ( .A(n35981), .B(n35979), .Z(n35969) );
  XOR U45474 ( .A(n35967), .B(n35969), .Z(n35989) );
  XOR U45475 ( .A(n32619), .B(n35989), .Z(n32620) );
  IV U45476 ( .A(n32620), .Z(n35960) );
  XOR U45477 ( .A(n35959), .B(n35960), .Z(n35963) );
  IV U45478 ( .A(n32621), .Z(n32623) );
  NOR U45479 ( .A(n32623), .B(n32622), .Z(n32624) );
  IV U45480 ( .A(n32624), .Z(n32625) );
  NOR U45481 ( .A(n32625), .B(n32631), .Z(n32626) );
  IV U45482 ( .A(n32626), .Z(n35962) );
  XOR U45483 ( .A(n35963), .B(n35962), .Z(n35953) );
  IV U45484 ( .A(n32627), .Z(n32636) );
  IV U45485 ( .A(n32628), .Z(n32629) );
  NOR U45486 ( .A(n32636), .B(n32629), .Z(n35954) );
  IV U45487 ( .A(n32630), .Z(n32632) );
  NOR U45488 ( .A(n32632), .B(n32631), .Z(n35956) );
  NOR U45489 ( .A(n35954), .B(n35956), .Z(n32633) );
  XOR U45490 ( .A(n35953), .B(n32633), .Z(n35995) );
  IV U45491 ( .A(n32634), .Z(n32635) );
  NOR U45492 ( .A(n32636), .B(n32635), .Z(n35993) );
  XOR U45493 ( .A(n35995), .B(n35993), .Z(n35997) );
  NOR U45494 ( .A(n32643), .B(n35997), .Z(n39261) );
  NOR U45495 ( .A(n32638), .B(n32637), .Z(n32639) );
  IV U45496 ( .A(n32639), .Z(n35949) );
  IV U45497 ( .A(n32640), .Z(n32641) );
  NOR U45498 ( .A(n32642), .B(n32641), .Z(n35996) );
  XOR U45499 ( .A(n35996), .B(n35997), .Z(n35948) );
  XOR U45500 ( .A(n35949), .B(n35948), .Z(n32646) );
  IV U45501 ( .A(n35948), .Z(n32644) );
  NOR U45502 ( .A(n32644), .B(n32643), .Z(n32645) );
  NOR U45503 ( .A(n32646), .B(n32645), .Z(n32647) );
  NOR U45504 ( .A(n39261), .B(n32647), .Z(n35946) );
  XOR U45505 ( .A(n32648), .B(n35946), .Z(n36006) );
  XOR U45506 ( .A(n32649), .B(n36006), .Z(n35940) );
  XOR U45507 ( .A(n32650), .B(n35940), .Z(n35938) );
  XOR U45508 ( .A(n32651), .B(n35938), .Z(n36012) );
  XOR U45509 ( .A(n36013), .B(n36012), .Z(n35931) );
  XOR U45510 ( .A(n35930), .B(n35931), .Z(n36009) );
  XOR U45511 ( .A(n36008), .B(n36009), .Z(n36023) );
  IV U45512 ( .A(n32652), .Z(n32654) );
  NOR U45513 ( .A(n32654), .B(n32653), .Z(n35926) );
  NOR U45514 ( .A(n35928), .B(n35926), .Z(n32655) );
  XOR U45515 ( .A(n36023), .B(n32655), .Z(n36029) );
  XOR U45516 ( .A(n32656), .B(n36029), .Z(n36027) );
  XOR U45517 ( .A(n36025), .B(n36027), .Z(n36037) );
  XOR U45518 ( .A(n36036), .B(n36037), .Z(n36040) );
  XOR U45519 ( .A(n36039), .B(n36040), .Z(n36035) );
  IV U45520 ( .A(n32657), .Z(n32659) );
  IV U45521 ( .A(n32658), .Z(n32661) );
  NOR U45522 ( .A(n32659), .B(n32661), .Z(n36033) );
  XOR U45523 ( .A(n36035), .B(n36033), .Z(n36047) );
  IV U45524 ( .A(n32660), .Z(n32662) );
  NOR U45525 ( .A(n32662), .B(n32661), .Z(n36045) );
  XOR U45526 ( .A(n36047), .B(n36045), .Z(n35924) );
  XOR U45527 ( .A(n35923), .B(n35924), .Z(n36059) );
  IV U45528 ( .A(n32663), .Z(n32664) );
  NOR U45529 ( .A(n32667), .B(n32664), .Z(n35921) );
  IV U45530 ( .A(n32665), .Z(n32666) );
  NOR U45531 ( .A(n32667), .B(n32666), .Z(n36057) );
  NOR U45532 ( .A(n35921), .B(n36057), .Z(n32668) );
  XOR U45533 ( .A(n36059), .B(n32668), .Z(n32677) );
  IV U45534 ( .A(n32677), .Z(n35920) );
  NOR U45535 ( .A(n32678), .B(n35920), .Z(n39318) );
  IV U45536 ( .A(n32669), .Z(n32671) );
  NOR U45537 ( .A(n32671), .B(n32670), .Z(n32672) );
  IV U45538 ( .A(n32672), .Z(n35916) );
  IV U45539 ( .A(n32673), .Z(n32675) );
  NOR U45540 ( .A(n32675), .B(n32674), .Z(n32676) );
  IV U45541 ( .A(n32676), .Z(n35919) );
  XOR U45542 ( .A(n32677), .B(n35919), .Z(n35915) );
  XOR U45543 ( .A(n35916), .B(n35915), .Z(n32681) );
  IV U45544 ( .A(n35915), .Z(n32679) );
  NOR U45545 ( .A(n32679), .B(n32678), .Z(n32680) );
  NOR U45546 ( .A(n32681), .B(n32680), .Z(n32682) );
  NOR U45547 ( .A(n39318), .B(n32682), .Z(n36062) );
  XOR U45548 ( .A(n32683), .B(n36062), .Z(n36069) );
  XOR U45549 ( .A(n36067), .B(n36069), .Z(n36071) );
  XOR U45550 ( .A(n36070), .B(n36071), .Z(n35911) );
  XOR U45551 ( .A(n35910), .B(n35911), .Z(n36075) );
  IV U45552 ( .A(n32684), .Z(n32685) );
  NOR U45553 ( .A(n32686), .B(n32685), .Z(n35913) );
  NOR U45554 ( .A(n32688), .B(n32687), .Z(n35908) );
  NOR U45555 ( .A(n35913), .B(n35908), .Z(n32689) );
  IV U45556 ( .A(n32689), .Z(n32690) );
  NOR U45557 ( .A(n36074), .B(n32690), .Z(n32691) );
  XOR U45558 ( .A(n36075), .B(n32691), .Z(n36080) );
  NOR U45559 ( .A(n32693), .B(n32692), .Z(n36077) );
  NOR U45560 ( .A(n36077), .B(n36079), .Z(n32694) );
  XOR U45561 ( .A(n36080), .B(n32694), .Z(n36088) );
  XOR U45562 ( .A(n32695), .B(n36088), .Z(n35900) );
  XOR U45563 ( .A(n32696), .B(n35900), .Z(n35898) );
  XOR U45564 ( .A(n35896), .B(n35898), .Z(n35894) );
  IV U45565 ( .A(n35894), .Z(n32703) );
  NOR U45566 ( .A(n32698), .B(n32697), .Z(n35893) );
  IV U45567 ( .A(n32699), .Z(n32701) );
  NOR U45568 ( .A(n32701), .B(n32700), .Z(n35888) );
  NOR U45569 ( .A(n35893), .B(n35888), .Z(n32702) );
  XOR U45570 ( .A(n32703), .B(n32702), .Z(n35892) );
  XOR U45571 ( .A(n35890), .B(n35892), .Z(n36095) );
  XOR U45572 ( .A(n36092), .B(n36095), .Z(n35886) );
  XOR U45573 ( .A(n32704), .B(n35886), .Z(n32705) );
  IV U45574 ( .A(n32705), .Z(n35884) );
  XOR U45575 ( .A(n35882), .B(n35884), .Z(n36106) );
  XOR U45576 ( .A(n36099), .B(n36106), .Z(n36102) );
  NOR U45577 ( .A(n32707), .B(n32706), .Z(n36105) );
  NOR U45578 ( .A(n36101), .B(n36105), .Z(n32708) );
  XOR U45579 ( .A(n36102), .B(n32708), .Z(n32709) );
  IV U45580 ( .A(n32709), .Z(n35873) );
  IV U45581 ( .A(n32710), .Z(n32712) );
  NOR U45582 ( .A(n32712), .B(n32711), .Z(n32713) );
  IV U45583 ( .A(n32713), .Z(n32718) );
  NOR U45584 ( .A(n35873), .B(n32718), .Z(n39150) );
  XOR U45585 ( .A(n32714), .B(n35873), .Z(n35870) );
  IV U45586 ( .A(n32715), .Z(n32716) );
  NOR U45587 ( .A(n32717), .B(n32716), .Z(n32719) );
  IV U45588 ( .A(n32719), .Z(n35869) );
  XOR U45589 ( .A(n35870), .B(n35869), .Z(n32721) );
  NOR U45590 ( .A(n32719), .B(n32718), .Z(n32720) );
  NOR U45591 ( .A(n32721), .B(n32720), .Z(n32722) );
  NOR U45592 ( .A(n39150), .B(n32722), .Z(n36119) );
  XOR U45593 ( .A(n36120), .B(n36119), .Z(n36117) );
  XOR U45594 ( .A(n36116), .B(n36117), .Z(n36133) );
  NOR U45595 ( .A(n32724), .B(n32723), .Z(n32725) );
  IV U45596 ( .A(n32725), .Z(n32726) );
  NOR U45597 ( .A(n32727), .B(n32726), .Z(n36131) );
  XOR U45598 ( .A(n36133), .B(n36131), .Z(n36129) );
  XOR U45599 ( .A(n36128), .B(n36129), .Z(n35865) );
  IV U45600 ( .A(n32728), .Z(n32729) );
  NOR U45601 ( .A(n32730), .B(n32729), .Z(n35863) );
  XOR U45602 ( .A(n35865), .B(n35863), .Z(n36145) );
  IV U45603 ( .A(n36145), .Z(n32739) );
  IV U45604 ( .A(n32731), .Z(n32732) );
  NOR U45605 ( .A(n32734), .B(n32732), .Z(n35866) );
  IV U45606 ( .A(n32733), .Z(n32737) );
  NOR U45607 ( .A(n32735), .B(n32734), .Z(n32736) );
  IV U45608 ( .A(n32736), .Z(n32741) );
  NOR U45609 ( .A(n32737), .B(n32741), .Z(n36143) );
  NOR U45610 ( .A(n35866), .B(n36143), .Z(n32738) );
  XOR U45611 ( .A(n32739), .B(n32738), .Z(n35862) );
  IV U45612 ( .A(n32740), .Z(n32742) );
  NOR U45613 ( .A(n32742), .B(n32741), .Z(n35860) );
  XOR U45614 ( .A(n35862), .B(n35860), .Z(n36149) );
  XOR U45615 ( .A(n36147), .B(n36149), .Z(n36151) );
  IV U45616 ( .A(n32743), .Z(n32745) );
  NOR U45617 ( .A(n32745), .B(n32744), .Z(n32746) );
  IV U45618 ( .A(n32746), .Z(n32750) );
  NOR U45619 ( .A(n36151), .B(n32750), .Z(n39415) );
  IV U45620 ( .A(n32747), .Z(n32749) );
  NOR U45621 ( .A(n32749), .B(n32748), .Z(n32751) );
  IV U45622 ( .A(n32751), .Z(n36150) );
  XOR U45623 ( .A(n36151), .B(n36150), .Z(n32753) );
  NOR U45624 ( .A(n32751), .B(n32750), .Z(n32752) );
  NOR U45625 ( .A(n32753), .B(n32752), .Z(n36163) );
  NOR U45626 ( .A(n39415), .B(n36163), .Z(n35858) );
  XOR U45627 ( .A(n36162), .B(n35858), .Z(n32754) );
  XOR U45628 ( .A(n35859), .B(n32754), .Z(n32761) );
  IV U45629 ( .A(n32761), .Z(n32755) );
  NOR U45630 ( .A(n32756), .B(n32755), .Z(n32757) );
  IV U45631 ( .A(n32757), .Z(n39124) );
  NOR U45632 ( .A(n32758), .B(n39124), .Z(n36166) );
  NOR U45633 ( .A(n39126), .B(n32759), .Z(n32764) );
  NOR U45634 ( .A(n32761), .B(n32760), .Z(n32762) );
  IV U45635 ( .A(n32762), .Z(n32763) );
  NOR U45636 ( .A(n32764), .B(n32763), .Z(n32765) );
  NOR U45637 ( .A(n36166), .B(n32765), .Z(n35852) );
  IV U45638 ( .A(n32766), .Z(n32768) );
  NOR U45639 ( .A(n32768), .B(n32767), .Z(n39426) );
  NOR U45640 ( .A(n39119), .B(n39426), .Z(n35853) );
  XOR U45641 ( .A(n35852), .B(n35853), .Z(n35856) );
  XOR U45642 ( .A(n32769), .B(n35856), .Z(n35843) );
  IV U45643 ( .A(n35843), .Z(n35851) );
  XOR U45644 ( .A(n32770), .B(n35851), .Z(n36171) );
  XOR U45645 ( .A(n36169), .B(n36171), .Z(n36179) );
  IV U45646 ( .A(n36179), .Z(n32778) );
  IV U45647 ( .A(n32771), .Z(n32772) );
  NOR U45648 ( .A(n32772), .B(n36172), .Z(n32776) );
  IV U45649 ( .A(n32773), .Z(n32775) );
  NOR U45650 ( .A(n32775), .B(n32774), .Z(n36178) );
  NOR U45651 ( .A(n32776), .B(n36178), .Z(n32777) );
  XOR U45652 ( .A(n32778), .B(n32777), .Z(n35840) );
  XOR U45653 ( .A(n35838), .B(n35840), .Z(n36185) );
  XOR U45654 ( .A(n36183), .B(n36185), .Z(n35836) );
  XOR U45655 ( .A(n35835), .B(n35836), .Z(n35830) );
  XOR U45656 ( .A(n35829), .B(n35830), .Z(n35833) );
  XOR U45657 ( .A(n35832), .B(n35833), .Z(n35827) );
  XOR U45658 ( .A(n32779), .B(n35827), .Z(n32787) );
  IV U45659 ( .A(n32787), .Z(n32780) );
  NOR U45660 ( .A(n32786), .B(n32780), .Z(n39470) );
  IV U45661 ( .A(n32783), .Z(n32782) );
  XOR U45662 ( .A(n35824), .B(n35827), .Z(n32781) );
  NOR U45663 ( .A(n32782), .B(n32781), .Z(n39116) );
  NOR U45664 ( .A(n39470), .B(n39116), .Z(n36195) );
  IV U45665 ( .A(n36195), .Z(n32785) );
  NOR U45666 ( .A(n32783), .B(n32787), .Z(n32784) );
  NOR U45667 ( .A(n32785), .B(n32784), .Z(n32789) );
  NOR U45668 ( .A(n32787), .B(n32786), .Z(n32788) );
  NOR U45669 ( .A(n32789), .B(n32788), .Z(n35820) );
  NOR U45670 ( .A(n32791), .B(n32790), .Z(n35818) );
  XOR U45671 ( .A(n35820), .B(n35818), .Z(n35823) );
  XOR U45672 ( .A(n35821), .B(n35823), .Z(n35815) );
  XOR U45673 ( .A(n32792), .B(n35815), .Z(n32793) );
  IV U45674 ( .A(n32793), .Z(n35811) );
  XOR U45675 ( .A(n35809), .B(n35811), .Z(n36199) );
  IV U45676 ( .A(n32794), .Z(n32795) );
  NOR U45677 ( .A(n32796), .B(n32795), .Z(n36197) );
  XOR U45678 ( .A(n36199), .B(n36197), .Z(n35804) );
  IV U45679 ( .A(n35804), .Z(n32803) );
  IV U45680 ( .A(n32797), .Z(n35806) );
  NOR U45681 ( .A(n35806), .B(n32798), .Z(n32801) );
  IV U45682 ( .A(n32799), .Z(n32800) );
  NOR U45683 ( .A(n32804), .B(n32800), .Z(n35802) );
  NOR U45684 ( .A(n32801), .B(n35802), .Z(n32802) );
  XOR U45685 ( .A(n32803), .B(n32802), .Z(n35798) );
  NOR U45686 ( .A(n32805), .B(n32804), .Z(n32806) );
  IV U45687 ( .A(n32806), .Z(n32807) );
  NOR U45688 ( .A(n32808), .B(n32807), .Z(n35796) );
  XOR U45689 ( .A(n35798), .B(n35796), .Z(n35801) );
  XOR U45690 ( .A(n35799), .B(n35801), .Z(n35795) );
  XOR U45691 ( .A(n35793), .B(n35795), .Z(n36204) );
  XOR U45692 ( .A(n36205), .B(n36204), .Z(n35789) );
  IV U45693 ( .A(n32809), .Z(n32810) );
  NOR U45694 ( .A(n32811), .B(n32810), .Z(n36206) );
  IV U45695 ( .A(n32812), .Z(n32814) );
  NOR U45696 ( .A(n32814), .B(n32813), .Z(n35791) );
  NOR U45697 ( .A(n35788), .B(n35791), .Z(n32815) );
  XOR U45698 ( .A(n36206), .B(n32815), .Z(n32816) );
  XOR U45699 ( .A(n35789), .B(n32816), .Z(n35784) );
  XOR U45700 ( .A(n35782), .B(n35784), .Z(n35786) );
  XOR U45701 ( .A(n35785), .B(n35786), .Z(n36216) );
  IV U45702 ( .A(n32817), .Z(n32818) );
  NOR U45703 ( .A(n32819), .B(n32818), .Z(n35780) );
  NOR U45704 ( .A(n32821), .B(n32820), .Z(n36215) );
  NOR U45705 ( .A(n35780), .B(n36215), .Z(n32822) );
  XOR U45706 ( .A(n36216), .B(n32822), .Z(n35775) );
  IV U45707 ( .A(n32823), .Z(n32825) );
  NOR U45708 ( .A(n32825), .B(n32824), .Z(n35776) );
  NOR U45709 ( .A(n36212), .B(n35776), .Z(n32826) );
  XOR U45710 ( .A(n35775), .B(n32826), .Z(n39106) );
  NOR U45711 ( .A(n32827), .B(n32829), .Z(n39521) );
  IV U45712 ( .A(n32828), .Z(n32830) );
  NOR U45713 ( .A(n32830), .B(n32829), .Z(n39105) );
  NOR U45714 ( .A(n39521), .B(n39105), .Z(n35778) );
  XOR U45715 ( .A(n39106), .B(n35778), .Z(n36221) );
  XOR U45716 ( .A(n36222), .B(n36221), .Z(n36224) );
  XOR U45717 ( .A(n36225), .B(n36224), .Z(n32835) );
  IV U45718 ( .A(n32835), .Z(n32831) );
  NOR U45719 ( .A(n32832), .B(n32831), .Z(n39091) );
  IV U45720 ( .A(n32833), .Z(n35774) );
  IV U45721 ( .A(n32836), .Z(n32834) );
  NOR U45722 ( .A(n32834), .B(n36224), .Z(n39096) );
  NOR U45723 ( .A(n32836), .B(n32835), .Z(n32837) );
  NOR U45724 ( .A(n39096), .B(n32837), .Z(n32838) );
  IV U45725 ( .A(n32838), .Z(n35773) );
  XOR U45726 ( .A(n35774), .B(n35773), .Z(n32839) );
  NOR U45727 ( .A(n32840), .B(n32839), .Z(n32841) );
  NOR U45728 ( .A(n39091), .B(n32841), .Z(n36229) );
  XOR U45729 ( .A(n36232), .B(n36229), .Z(n36237) );
  XOR U45730 ( .A(n32842), .B(n36237), .Z(n35767) );
  XOR U45731 ( .A(n32843), .B(n35767), .Z(n35766) );
  XOR U45732 ( .A(n32844), .B(n35766), .Z(n35752) );
  XOR U45733 ( .A(n32845), .B(n35752), .Z(n35746) );
  IV U45734 ( .A(n32846), .Z(n32847) );
  NOR U45735 ( .A(n35753), .B(n32847), .Z(n35748) );
  IV U45736 ( .A(n32848), .Z(n32850) );
  NOR U45737 ( .A(n32850), .B(n32849), .Z(n35745) );
  NOR U45738 ( .A(n35748), .B(n35745), .Z(n32851) );
  XOR U45739 ( .A(n35746), .B(n32851), .Z(n35741) );
  XOR U45740 ( .A(n35739), .B(n35741), .Z(n35744) );
  XOR U45741 ( .A(n32852), .B(n35744), .Z(n36243) );
  IV U45742 ( .A(n32853), .Z(n32855) );
  NOR U45743 ( .A(n32855), .B(n32854), .Z(n32856) );
  IV U45744 ( .A(n32856), .Z(n32857) );
  NOR U45745 ( .A(n32858), .B(n32857), .Z(n32859) );
  IV U45746 ( .A(n32859), .Z(n36244) );
  XOR U45747 ( .A(n36243), .B(n36244), .Z(n35733) );
  XOR U45748 ( .A(n35733), .B(n32860), .Z(n35730) );
  XOR U45749 ( .A(n35727), .B(n35730), .Z(n36256) );
  IV U45750 ( .A(n36256), .Z(n32868) );
  IV U45751 ( .A(n32861), .Z(n32863) );
  NOR U45752 ( .A(n32863), .B(n32862), .Z(n35729) );
  IV U45753 ( .A(n32864), .Z(n32865) );
  NOR U45754 ( .A(n32866), .B(n32865), .Z(n36255) );
  NOR U45755 ( .A(n35729), .B(n36255), .Z(n32867) );
  XOR U45756 ( .A(n32868), .B(n32867), .Z(n36254) );
  IV U45757 ( .A(n32869), .Z(n32871) );
  NOR U45758 ( .A(n32871), .B(n32870), .Z(n36252) );
  XOR U45759 ( .A(n36254), .B(n36252), .Z(n35724) );
  XOR U45760 ( .A(n35723), .B(n35724), .Z(n36263) );
  XOR U45761 ( .A(n36261), .B(n36263), .Z(n36272) );
  XOR U45762 ( .A(n35721), .B(n36272), .Z(n36280) );
  XOR U45763 ( .A(n32872), .B(n36280), .Z(n32873) );
  IV U45764 ( .A(n32873), .Z(n36277) );
  IV U45765 ( .A(n32874), .Z(n32875) );
  NOR U45766 ( .A(n32881), .B(n32875), .Z(n32884) );
  IV U45767 ( .A(n32884), .Z(n32876) );
  NOR U45768 ( .A(n36277), .B(n32876), .Z(n39056) );
  IV U45769 ( .A(n32877), .Z(n32879) );
  NOR U45770 ( .A(n32879), .B(n32878), .Z(n32880) );
  IV U45771 ( .A(n32880), .Z(n32882) );
  NOR U45772 ( .A(n32882), .B(n32881), .Z(n36275) );
  XOR U45773 ( .A(n36275), .B(n36277), .Z(n32888) );
  IV U45774 ( .A(n32888), .Z(n32883) );
  NOR U45775 ( .A(n32884), .B(n32883), .Z(n32885) );
  NOR U45776 ( .A(n39056), .B(n32885), .Z(n32886) );
  NOR U45777 ( .A(n32887), .B(n32886), .Z(n32890) );
  IV U45778 ( .A(n32887), .Z(n32889) );
  NOR U45779 ( .A(n32889), .B(n32888), .Z(n39572) );
  NOR U45780 ( .A(n32890), .B(n39572), .Z(n35716) );
  IV U45781 ( .A(n32891), .Z(n32893) );
  NOR U45782 ( .A(n32893), .B(n32892), .Z(n35715) );
  NOR U45783 ( .A(n35718), .B(n35715), .Z(n32894) );
  XOR U45784 ( .A(n35716), .B(n32894), .Z(n36286) );
  IV U45785 ( .A(n32895), .Z(n32897) );
  NOR U45786 ( .A(n32897), .B(n32896), .Z(n36284) );
  XOR U45787 ( .A(n36286), .B(n36284), .Z(n36289) );
  XOR U45788 ( .A(n36287), .B(n36289), .Z(n35713) );
  XOR U45789 ( .A(n32898), .B(n35713), .Z(n35700) );
  IV U45790 ( .A(n32899), .Z(n32901) );
  NOR U45791 ( .A(n32901), .B(n32900), .Z(n35702) );
  NOR U45792 ( .A(n35699), .B(n35702), .Z(n32902) );
  XOR U45793 ( .A(n35700), .B(n32902), .Z(n35708) );
  XOR U45794 ( .A(n35706), .B(n35708), .Z(n35695) );
  XOR U45795 ( .A(n35693), .B(n35695), .Z(n35698) );
  XOR U45796 ( .A(n35696), .B(n35698), .Z(n35689) );
  XOR U45797 ( .A(n32903), .B(n35689), .Z(n35685) );
  XOR U45798 ( .A(n32904), .B(n35685), .Z(n36304) );
  XOR U45799 ( .A(n35683), .B(n36304), .Z(n35681) );
  XOR U45800 ( .A(n32905), .B(n35681), .Z(n35673) );
  XOR U45801 ( .A(n32906), .B(n35673), .Z(n42454) );
  XOR U45802 ( .A(n36307), .B(n42454), .Z(n35669) );
  IV U45803 ( .A(n32907), .Z(n32909) );
  NOR U45804 ( .A(n32909), .B(n32908), .Z(n32910) );
  IV U45805 ( .A(n32910), .Z(n35670) );
  XOR U45806 ( .A(n35669), .B(n35670), .Z(n36314) );
  XOR U45807 ( .A(n32911), .B(n36314), .Z(n32912) );
  IV U45808 ( .A(n32912), .Z(n36326) );
  NOR U45809 ( .A(n32913), .B(n36326), .Z(n32915) );
  IV U45810 ( .A(n32913), .Z(n32914) );
  NOR U45811 ( .A(n32914), .B(n36314), .Z(n39620) );
  NOR U45812 ( .A(n32915), .B(n39620), .Z(n36330) );
  IV U45813 ( .A(n32916), .Z(n32920) );
  NOR U45814 ( .A(n32918), .B(n32917), .Z(n32919) );
  IV U45815 ( .A(n32919), .Z(n32923) );
  NOR U45816 ( .A(n32920), .B(n32923), .Z(n32921) );
  IV U45817 ( .A(n32921), .Z(n36331) );
  XOR U45818 ( .A(n36330), .B(n36331), .Z(n35665) );
  IV U45819 ( .A(n32922), .Z(n32924) );
  NOR U45820 ( .A(n32924), .B(n32923), .Z(n35663) );
  XOR U45821 ( .A(n35665), .B(n35663), .Z(n35668) );
  IV U45822 ( .A(n32925), .Z(n32927) );
  NOR U45823 ( .A(n32927), .B(n32926), .Z(n35666) );
  XOR U45824 ( .A(n35668), .B(n35666), .Z(n35661) );
  XOR U45825 ( .A(n35660), .B(n35661), .Z(n35648) );
  NOR U45826 ( .A(n32928), .B(n35649), .Z(n32932) );
  IV U45827 ( .A(n32929), .Z(n32931) );
  NOR U45828 ( .A(n32931), .B(n32930), .Z(n35645) );
  NOR U45829 ( .A(n32932), .B(n35645), .Z(n32933) );
  XOR U45830 ( .A(n35648), .B(n32933), .Z(n35639) );
  IV U45831 ( .A(n32934), .Z(n32935) );
  NOR U45832 ( .A(n32935), .B(n36337), .Z(n35642) );
  IV U45833 ( .A(n32936), .Z(n32938) );
  NOR U45834 ( .A(n32938), .B(n32937), .Z(n35640) );
  NOR U45835 ( .A(n35642), .B(n35640), .Z(n32939) );
  XOR U45836 ( .A(n35639), .B(n32939), .Z(n36347) );
  IV U45837 ( .A(n32940), .Z(n32944) );
  NOR U45838 ( .A(n32942), .B(n32941), .Z(n32943) );
  IV U45839 ( .A(n32943), .Z(n32948) );
  NOR U45840 ( .A(n32944), .B(n32948), .Z(n36346) );
  NOR U45841 ( .A(n32945), .B(n36346), .Z(n32946) );
  XOR U45842 ( .A(n36347), .B(n32946), .Z(n36350) );
  IV U45843 ( .A(n32947), .Z(n32949) );
  NOR U45844 ( .A(n32949), .B(n32948), .Z(n32950) );
  IV U45845 ( .A(n32950), .Z(n36351) );
  XOR U45846 ( .A(n36350), .B(n36351), .Z(n36366) );
  XOR U45847 ( .A(n32951), .B(n36366), .Z(n32952) );
  IV U45848 ( .A(n32952), .Z(n36358) );
  XOR U45849 ( .A(n36356), .B(n36358), .Z(n36362) );
  IV U45850 ( .A(n36362), .Z(n32960) );
  IV U45851 ( .A(n32953), .Z(n32954) );
  NOR U45852 ( .A(n32955), .B(n32954), .Z(n35636) );
  IV U45853 ( .A(n32956), .Z(n32957) );
  NOR U45854 ( .A(n32958), .B(n32957), .Z(n36360) );
  NOR U45855 ( .A(n35636), .B(n36360), .Z(n32959) );
  XOR U45856 ( .A(n32960), .B(n32959), .Z(n35631) );
  XOR U45857 ( .A(n35630), .B(n35631), .Z(n35634) );
  XOR U45858 ( .A(n35633), .B(n35634), .Z(n35628) );
  XOR U45859 ( .A(n32961), .B(n35628), .Z(n32962) );
  IV U45860 ( .A(n32962), .Z(n35615) );
  XOR U45861 ( .A(n32963), .B(n35615), .Z(n35612) );
  XOR U45862 ( .A(n35610), .B(n35612), .Z(n36375) );
  XOR U45863 ( .A(n36374), .B(n36375), .Z(n36378) );
  IV U45864 ( .A(n36378), .Z(n32970) );
  NOR U45865 ( .A(n32965), .B(n32964), .Z(n36377) );
  IV U45866 ( .A(n32966), .Z(n32968) );
  NOR U45867 ( .A(n32968), .B(n32967), .Z(n35608) );
  NOR U45868 ( .A(n36377), .B(n35608), .Z(n32969) );
  XOR U45869 ( .A(n32970), .B(n32969), .Z(n35607) );
  XOR U45870 ( .A(n35605), .B(n35607), .Z(n36386) );
  XOR U45871 ( .A(n36385), .B(n36386), .Z(n35603) );
  XOR U45872 ( .A(n35601), .B(n35603), .Z(n49190) );
  XOR U45873 ( .A(n36382), .B(n49190), .Z(n36398) );
  XOR U45874 ( .A(n36397), .B(n36398), .Z(n35599) );
  XOR U45875 ( .A(n35598), .B(n35599), .Z(n36407) );
  XOR U45876 ( .A(n32971), .B(n36407), .Z(n36408) );
  IV U45877 ( .A(n32972), .Z(n32974) );
  NOR U45878 ( .A(n32974), .B(n32973), .Z(n32975) );
  IV U45879 ( .A(n32975), .Z(n36409) );
  XOR U45880 ( .A(n36408), .B(n36409), .Z(n35591) );
  IV U45881 ( .A(n32976), .Z(n35594) );
  NOR U45882 ( .A(n32978), .B(n32977), .Z(n32979) );
  IV U45883 ( .A(n32979), .Z(n35592) );
  NOR U45884 ( .A(n35594), .B(n35592), .Z(n32980) );
  XOR U45885 ( .A(n35591), .B(n32980), .Z(n35597) );
  IV U45886 ( .A(n32981), .Z(n32982) );
  NOR U45887 ( .A(n32982), .B(n32986), .Z(n35589) );
  IV U45888 ( .A(n32983), .Z(n32984) );
  NOR U45889 ( .A(n32984), .B(n35592), .Z(n35595) );
  NOR U45890 ( .A(n35589), .B(n35595), .Z(n32985) );
  XOR U45891 ( .A(n35597), .B(n32985), .Z(n32997) );
  IV U45892 ( .A(n32997), .Z(n32987) );
  NOR U45893 ( .A(n32987), .B(n32986), .Z(n32988) );
  IV U45894 ( .A(n32988), .Z(n32989) );
  NOR U45895 ( .A(n32990), .B(n32989), .Z(n32991) );
  IV U45896 ( .A(n32991), .Z(n39700) );
  NOR U45897 ( .A(n32992), .B(n39700), .Z(n36413) );
  IV U45898 ( .A(n32993), .Z(n32995) );
  NOR U45899 ( .A(n32995), .B(n32994), .Z(n32996) );
  NOR U45900 ( .A(n32997), .B(n32996), .Z(n32998) );
  NOR U45901 ( .A(n36413), .B(n32998), .Z(n36414) );
  XOR U45902 ( .A(n36416), .B(n36414), .Z(n36419) );
  XOR U45903 ( .A(n36417), .B(n36419), .Z(n36431) );
  XOR U45904 ( .A(n36429), .B(n36431), .Z(n36423) );
  XOR U45905 ( .A(n36422), .B(n36423), .Z(n36439) );
  XOR U45906 ( .A(n32999), .B(n36439), .Z(n35581) );
  IV U45907 ( .A(n33000), .Z(n33002) );
  NOR U45908 ( .A(n33002), .B(n33001), .Z(n35586) );
  IV U45909 ( .A(n33003), .Z(n33012) );
  NOR U45910 ( .A(n33012), .B(n33004), .Z(n35584) );
  IV U45911 ( .A(n33005), .Z(n33006) );
  NOR U45912 ( .A(n33006), .B(n33019), .Z(n35580) );
  NOR U45913 ( .A(n35584), .B(n35580), .Z(n33007) );
  IV U45914 ( .A(n33007), .Z(n33008) );
  NOR U45915 ( .A(n35586), .B(n33008), .Z(n33009) );
  XOR U45916 ( .A(n35581), .B(n33009), .Z(n36443) );
  IV U45917 ( .A(n33010), .Z(n33011) );
  NOR U45918 ( .A(n33012), .B(n33011), .Z(n36441) );
  XOR U45919 ( .A(n36443), .B(n36441), .Z(n36446) );
  IV U45920 ( .A(n33013), .Z(n33016) );
  NOR U45921 ( .A(n33014), .B(n33019), .Z(n33015) );
  IV U45922 ( .A(n33015), .Z(n33027) );
  NOR U45923 ( .A(n33016), .B(n33027), .Z(n33017) );
  IV U45924 ( .A(n33017), .Z(n33029) );
  NOR U45925 ( .A(n36446), .B(n33029), .Z(n36448) );
  IV U45926 ( .A(n33018), .Z(n33024) );
  XOR U45927 ( .A(n33020), .B(n33019), .Z(n33022) );
  NOR U45928 ( .A(n33022), .B(n33021), .Z(n33023) );
  IV U45929 ( .A(n33023), .Z(n33035) );
  NOR U45930 ( .A(n33024), .B(n33035), .Z(n33025) );
  IV U45931 ( .A(n33025), .Z(n36450) );
  IV U45932 ( .A(n33026), .Z(n33028) );
  NOR U45933 ( .A(n33028), .B(n33027), .Z(n36444) );
  XOR U45934 ( .A(n36446), .B(n36444), .Z(n36449) );
  XOR U45935 ( .A(n36450), .B(n36449), .Z(n33032) );
  IV U45936 ( .A(n36449), .Z(n33030) );
  NOR U45937 ( .A(n33030), .B(n33029), .Z(n33031) );
  NOR U45938 ( .A(n33032), .B(n33031), .Z(n33033) );
  NOR U45939 ( .A(n36448), .B(n33033), .Z(n35574) );
  IV U45940 ( .A(n33034), .Z(n33036) );
  NOR U45941 ( .A(n33036), .B(n33035), .Z(n33037) );
  IV U45942 ( .A(n33037), .Z(n35575) );
  XOR U45943 ( .A(n35574), .B(n35575), .Z(n35570) );
  NOR U45944 ( .A(n35569), .B(n35577), .Z(n33038) );
  NOR U45945 ( .A(n33038), .B(n35571), .Z(n33039) );
  XOR U45946 ( .A(n35570), .B(n33039), .Z(n35567) );
  XOR U45947 ( .A(n35564), .B(n35567), .Z(n36457) );
  IV U45948 ( .A(n36457), .Z(n33047) );
  IV U45949 ( .A(n33040), .Z(n33041) );
  NOR U45950 ( .A(n33042), .B(n33041), .Z(n35566) );
  IV U45951 ( .A(n33043), .Z(n33045) );
  NOR U45952 ( .A(n33045), .B(n33044), .Z(n36456) );
  NOR U45953 ( .A(n35566), .B(n36456), .Z(n33046) );
  XOR U45954 ( .A(n33047), .B(n33046), .Z(n36455) );
  IV U45955 ( .A(n33048), .Z(n33049) );
  NOR U45956 ( .A(n33050), .B(n33049), .Z(n33051) );
  IV U45957 ( .A(n33051), .Z(n33053) );
  NOR U45958 ( .A(n33053), .B(n33052), .Z(n36453) );
  XOR U45959 ( .A(n36455), .B(n36453), .Z(n36462) );
  XOR U45960 ( .A(n33054), .B(n36462), .Z(n33055) );
  IV U45961 ( .A(n33055), .Z(n35561) );
  XOR U45962 ( .A(n35560), .B(n35561), .Z(n35553) );
  IV U45963 ( .A(n33056), .Z(n33058) );
  NOR U45964 ( .A(n33058), .B(n33057), .Z(n36463) );
  IV U45965 ( .A(n33059), .Z(n33060) );
  NOR U45966 ( .A(n33060), .B(n35554), .Z(n33061) );
  NOR U45967 ( .A(n36463), .B(n33061), .Z(n33062) );
  XOR U45968 ( .A(n35553), .B(n33062), .Z(n36476) );
  XOR U45969 ( .A(n36475), .B(n36476), .Z(n33063) );
  NOR U45970 ( .A(n33064), .B(n33063), .Z(n33079) );
  IV U45971 ( .A(n33065), .Z(n33069) );
  NOR U45972 ( .A(n36476), .B(n33066), .Z(n33067) );
  IV U45973 ( .A(n33067), .Z(n33068) );
  NOR U45974 ( .A(n33069), .B(n33068), .Z(n38947) );
  IV U45975 ( .A(n33070), .Z(n33076) );
  XOR U45976 ( .A(n33072), .B(n33071), .Z(n33073) );
  NOR U45977 ( .A(n36476), .B(n33073), .Z(n33074) );
  IV U45978 ( .A(n33074), .Z(n33075) );
  NOR U45979 ( .A(n33076), .B(n33075), .Z(n36482) );
  NOR U45980 ( .A(n38947), .B(n36482), .Z(n33077) );
  IV U45981 ( .A(n33077), .Z(n33078) );
  NOR U45982 ( .A(n33079), .B(n33078), .Z(n35550) );
  XOR U45983 ( .A(n33080), .B(n35550), .Z(n35547) );
  NOR U45984 ( .A(n33081), .B(n35537), .Z(n33082) );
  NOR U45985 ( .A(n33082), .B(n35544), .Z(n33083) );
  XOR U45986 ( .A(n35547), .B(n33083), .Z(n36492) );
  IV U45987 ( .A(n33084), .Z(n33085) );
  NOR U45988 ( .A(n33086), .B(n33085), .Z(n35534) );
  IV U45989 ( .A(n33087), .Z(n33088) );
  NOR U45990 ( .A(n33089), .B(n33088), .Z(n36491) );
  NOR U45991 ( .A(n35534), .B(n36491), .Z(n33090) );
  XOR U45992 ( .A(n36492), .B(n33090), .Z(n36488) );
  XOR U45993 ( .A(n36489), .B(n36488), .Z(n35529) );
  XOR U45994 ( .A(n35528), .B(n35529), .Z(n35532) );
  XOR U45995 ( .A(n33091), .B(n35532), .Z(n35520) );
  IV U45996 ( .A(n33092), .Z(n33096) );
  NOR U45997 ( .A(n33093), .B(n33098), .Z(n33094) );
  IV U45998 ( .A(n33094), .Z(n33095) );
  NOR U45999 ( .A(n33096), .B(n33095), .Z(n35521) );
  IV U46000 ( .A(n33097), .Z(n33102) );
  NOR U46001 ( .A(n33099), .B(n33098), .Z(n33100) );
  IV U46002 ( .A(n33100), .Z(n33101) );
  NOR U46003 ( .A(n33102), .B(n33101), .Z(n35523) );
  NOR U46004 ( .A(n35521), .B(n35523), .Z(n33103) );
  XOR U46005 ( .A(n35520), .B(n33103), .Z(n35509) );
  XOR U46006 ( .A(n33104), .B(n35509), .Z(n35493) );
  XOR U46007 ( .A(n35492), .B(n35493), .Z(n35496) );
  XOR U46008 ( .A(n35495), .B(n35496), .Z(n38898) );
  XOR U46009 ( .A(n36499), .B(n38898), .Z(n33105) );
  IV U46010 ( .A(n33105), .Z(n36502) );
  XOR U46011 ( .A(n36501), .B(n36502), .Z(n36508) );
  IV U46012 ( .A(n36508), .Z(n33113) );
  IV U46013 ( .A(n33106), .Z(n33107) );
  NOR U46014 ( .A(n33108), .B(n33107), .Z(n36507) );
  IV U46015 ( .A(n33109), .Z(n33110) );
  NOR U46016 ( .A(n33111), .B(n33110), .Z(n36504) );
  NOR U46017 ( .A(n36507), .B(n36504), .Z(n33112) );
  XOR U46018 ( .A(n33113), .B(n33112), .Z(n39797) );
  NOR U46019 ( .A(n33114), .B(n39800), .Z(n36510) );
  IV U46020 ( .A(n33115), .Z(n33117) );
  NOR U46021 ( .A(n33117), .B(n33116), .Z(n35490) );
  NOR U46022 ( .A(n36510), .B(n35490), .Z(n33118) );
  XOR U46023 ( .A(n39797), .B(n33118), .Z(n33119) );
  NOR U46024 ( .A(n33124), .B(n33119), .Z(n33127) );
  IV U46025 ( .A(n33120), .Z(n33122) );
  NOR U46026 ( .A(n33122), .B(n33121), .Z(n33128) );
  IV U46027 ( .A(n33128), .Z(n33123) );
  NOR U46028 ( .A(n33127), .B(n33123), .Z(n36514) );
  IV U46029 ( .A(n33124), .Z(n33126) );
  XOR U46030 ( .A(n36510), .B(n39797), .Z(n33125) );
  NOR U46031 ( .A(n33126), .B(n33125), .Z(n39809) );
  NOR U46032 ( .A(n39809), .B(n33127), .Z(n38886) );
  NOR U46033 ( .A(n33128), .B(n38886), .Z(n33129) );
  NOR U46034 ( .A(n36514), .B(n33129), .Z(n35484) );
  XOR U46035 ( .A(n35486), .B(n35484), .Z(n35488) );
  XOR U46036 ( .A(n33130), .B(n35488), .Z(n35480) );
  IV U46037 ( .A(n33131), .Z(n33132) );
  NOR U46038 ( .A(n33133), .B(n33132), .Z(n42300) );
  IV U46039 ( .A(n33134), .Z(n33135) );
  NOR U46040 ( .A(n33136), .B(n33135), .Z(n43268) );
  NOR U46041 ( .A(n42300), .B(n43268), .Z(n35481) );
  XOR U46042 ( .A(n35480), .B(n35481), .Z(n36516) );
  NOR U46043 ( .A(n33144), .B(n36516), .Z(n42292) );
  IV U46044 ( .A(n33137), .Z(n33138) );
  NOR U46045 ( .A(n33139), .B(n33138), .Z(n33140) );
  IV U46046 ( .A(n33140), .Z(n35476) );
  IV U46047 ( .A(n33141), .Z(n33143) );
  NOR U46048 ( .A(n33143), .B(n33142), .Z(n36515) );
  XOR U46049 ( .A(n36515), .B(n36516), .Z(n35475) );
  XOR U46050 ( .A(n35476), .B(n35475), .Z(n33147) );
  IV U46051 ( .A(n35475), .Z(n33145) );
  NOR U46052 ( .A(n33145), .B(n33144), .Z(n33146) );
  NOR U46053 ( .A(n33147), .B(n33146), .Z(n33148) );
  NOR U46054 ( .A(n42292), .B(n33148), .Z(n35478) );
  XOR U46055 ( .A(n33149), .B(n35478), .Z(n36521) );
  XOR U46056 ( .A(n36519), .B(n36521), .Z(n36535) );
  IV U46057 ( .A(n36535), .Z(n33155) );
  NOR U46058 ( .A(n33164), .B(n33150), .Z(n36534) );
  IV U46059 ( .A(n33151), .Z(n33153) );
  NOR U46060 ( .A(n33153), .B(n33152), .Z(n35473) );
  NOR U46061 ( .A(n36534), .B(n35473), .Z(n33154) );
  XOR U46062 ( .A(n33155), .B(n33154), .Z(n36540) );
  XOR U46063 ( .A(n36539), .B(n36540), .Z(n33165) );
  IV U46064 ( .A(n33165), .Z(n49073) );
  IV U46065 ( .A(n33156), .Z(n33160) );
  NOR U46066 ( .A(n33158), .B(n33157), .Z(n33159) );
  IV U46067 ( .A(n33159), .Z(n33173) );
  NOR U46068 ( .A(n33160), .B(n33173), .Z(n33169) );
  IV U46069 ( .A(n33169), .Z(n33161) );
  NOR U46070 ( .A(n49073), .B(n33161), .Z(n35472) );
  IV U46071 ( .A(n33162), .Z(n33163) );
  NOR U46072 ( .A(n33164), .B(n33163), .Z(n33166) );
  IV U46073 ( .A(n33166), .Z(n49063) );
  NOR U46074 ( .A(n36540), .B(n49063), .Z(n36538) );
  NOR U46075 ( .A(n33166), .B(n33165), .Z(n33167) );
  NOR U46076 ( .A(n36538), .B(n33167), .Z(n33168) );
  NOR U46077 ( .A(n33169), .B(n33168), .Z(n33170) );
  NOR U46078 ( .A(n35472), .B(n33170), .Z(n33171) );
  IV U46079 ( .A(n33171), .Z(n35470) );
  IV U46080 ( .A(n33172), .Z(n33174) );
  NOR U46081 ( .A(n33174), .B(n33173), .Z(n35468) );
  XOR U46082 ( .A(n35470), .B(n35468), .Z(n35463) );
  XOR U46083 ( .A(n35462), .B(n35463), .Z(n35466) );
  XOR U46084 ( .A(n35465), .B(n35466), .Z(n35457) );
  XOR U46085 ( .A(n35456), .B(n35457), .Z(n35461) );
  XOR U46086 ( .A(n33175), .B(n35461), .Z(n33176) );
  IV U46087 ( .A(n33176), .Z(n36553) );
  XOR U46088 ( .A(n36551), .B(n36553), .Z(n35449) );
  XOR U46089 ( .A(n35448), .B(n35449), .Z(n36549) );
  IV U46090 ( .A(n33177), .Z(n33181) );
  NOR U46091 ( .A(n33179), .B(n33178), .Z(n33180) );
  IV U46092 ( .A(n33180), .Z(n33186) );
  NOR U46093 ( .A(n33181), .B(n33186), .Z(n36547) );
  XOR U46094 ( .A(n36549), .B(n36547), .Z(n35447) );
  IV U46095 ( .A(n33182), .Z(n33184) );
  NOR U46096 ( .A(n33184), .B(n33183), .Z(n35443) );
  IV U46097 ( .A(n33185), .Z(n33187) );
  NOR U46098 ( .A(n33187), .B(n33186), .Z(n35445) );
  NOR U46099 ( .A(n35443), .B(n35445), .Z(n33188) );
  XOR U46100 ( .A(n35447), .B(n33188), .Z(n33189) );
  IV U46101 ( .A(n33189), .Z(n36562) );
  XOR U46102 ( .A(n36560), .B(n36562), .Z(n36564) );
  XOR U46103 ( .A(n36563), .B(n36564), .Z(n50105) );
  IV U46104 ( .A(n50105), .Z(n33190) );
  NOR U46105 ( .A(n33191), .B(n33190), .Z(n33200) );
  IV U46106 ( .A(n33192), .Z(n33195) );
  NOR U46107 ( .A(n33193), .B(n36564), .Z(n33194) );
  IV U46108 ( .A(n33194), .Z(n33197) );
  NOR U46109 ( .A(n33195), .B(n33197), .Z(n39875) );
  IV U46110 ( .A(n33196), .Z(n50099) );
  NOR U46111 ( .A(n50099), .B(n33197), .Z(n39874) );
  NOR U46112 ( .A(n39875), .B(n39874), .Z(n33198) );
  IV U46113 ( .A(n33198), .Z(n33199) );
  NOR U46114 ( .A(n33200), .B(n33199), .Z(n35438) );
  IV U46115 ( .A(n33201), .Z(n33203) );
  NOR U46116 ( .A(n33203), .B(n33202), .Z(n35441) );
  IV U46117 ( .A(n33204), .Z(n33205) );
  NOR U46118 ( .A(n33206), .B(n33205), .Z(n35437) );
  NOR U46119 ( .A(n35441), .B(n35437), .Z(n33207) );
  XOR U46120 ( .A(n35438), .B(n33207), .Z(n35436) );
  IV U46121 ( .A(n33208), .Z(n33210) );
  NOR U46122 ( .A(n33210), .B(n33209), .Z(n35432) );
  XOR U46123 ( .A(n35436), .B(n35432), .Z(n35431) );
  XOR U46124 ( .A(n33211), .B(n35431), .Z(n35423) );
  XOR U46125 ( .A(n35424), .B(n35423), .Z(n35426) );
  XOR U46126 ( .A(n35425), .B(n35426), .Z(n33218) );
  NOR U46127 ( .A(n33212), .B(n33218), .Z(n39913) );
  IV U46128 ( .A(n33213), .Z(n33214) );
  NOR U46129 ( .A(n33215), .B(n33214), .Z(n33220) );
  IV U46130 ( .A(n33220), .Z(n33216) );
  NOR U46131 ( .A(n33216), .B(n35426), .Z(n39909) );
  NOR U46132 ( .A(n39913), .B(n39909), .Z(n33217) );
  IV U46133 ( .A(n33217), .Z(n35422) );
  NOR U46134 ( .A(n35422), .B(n33218), .Z(n33223) );
  NOR U46135 ( .A(n33220), .B(n33219), .Z(n33221) );
  NOR U46136 ( .A(n33221), .B(n35422), .Z(n33222) );
  NOR U46137 ( .A(n33223), .B(n33222), .Z(n35415) );
  XOR U46138 ( .A(n33224), .B(n35415), .Z(n36584) );
  XOR U46139 ( .A(n33225), .B(n36584), .Z(n36580) );
  XOR U46140 ( .A(n33226), .B(n36580), .Z(n36600) );
  XOR U46141 ( .A(n33227), .B(n36600), .Z(n33228) );
  IV U46142 ( .A(n33228), .Z(n36598) );
  XOR U46143 ( .A(n36596), .B(n36598), .Z(n35410) );
  IV U46144 ( .A(n33229), .Z(n33231) );
  NOR U46145 ( .A(n33231), .B(n33230), .Z(n35408) );
  XOR U46146 ( .A(n35410), .B(n35408), .Z(n35403) );
  XOR U46147 ( .A(n35402), .B(n35403), .Z(n35406) );
  XOR U46148 ( .A(n35405), .B(n35406), .Z(n36606) );
  IV U46149 ( .A(n33232), .Z(n33234) );
  NOR U46150 ( .A(n33234), .B(n33233), .Z(n36604) );
  IV U46151 ( .A(n33235), .Z(n33236) );
  NOR U46152 ( .A(n33237), .B(n33236), .Z(n35400) );
  NOR U46153 ( .A(n36604), .B(n35400), .Z(n33238) );
  XOR U46154 ( .A(n36606), .B(n33238), .Z(n35398) );
  XOR U46155 ( .A(n42229), .B(n35398), .Z(n35395) );
  IV U46156 ( .A(n33239), .Z(n33240) );
  NOR U46157 ( .A(n33241), .B(n33240), .Z(n35392) );
  NOR U46158 ( .A(n35394), .B(n35392), .Z(n33242) );
  XOR U46159 ( .A(n35395), .B(n33242), .Z(n36609) );
  XOR U46160 ( .A(n36611), .B(n36609), .Z(n36614) );
  XOR U46161 ( .A(n36612), .B(n36614), .Z(n38823) );
  XOR U46162 ( .A(n36616), .B(n38823), .Z(n33243) );
  IV U46163 ( .A(n33243), .Z(n38816) );
  XOR U46164 ( .A(n36617), .B(n38816), .Z(n33251) );
  IV U46165 ( .A(n33251), .Z(n33244) );
  NOR U46166 ( .A(n33245), .B(n33244), .Z(n42207) );
  IV U46167 ( .A(n33246), .Z(n33248) );
  NOR U46168 ( .A(n33248), .B(n33247), .Z(n33250) );
  IV U46169 ( .A(n33250), .Z(n33249) );
  NOR U46170 ( .A(n38816), .B(n33249), .Z(n38810) );
  NOR U46171 ( .A(n33251), .B(n33250), .Z(n33252) );
  NOR U46172 ( .A(n38810), .B(n33252), .Z(n33253) );
  NOR U46173 ( .A(n33254), .B(n33253), .Z(n33255) );
  NOR U46174 ( .A(n42207), .B(n33255), .Z(n33256) );
  IV U46175 ( .A(n33256), .Z(n35390) );
  XOR U46176 ( .A(n35389), .B(n35390), .Z(n35386) );
  IV U46177 ( .A(n33257), .Z(n33258) );
  NOR U46178 ( .A(n33258), .B(n33268), .Z(n35383) );
  NOR U46179 ( .A(n35385), .B(n35383), .Z(n33259) );
  XOR U46180 ( .A(n35386), .B(n33259), .Z(n33260) );
  IV U46181 ( .A(n33260), .Z(n36622) );
  IV U46182 ( .A(n33261), .Z(n33264) );
  IV U46183 ( .A(n33262), .Z(n33263) );
  NOR U46184 ( .A(n33264), .B(n33263), .Z(n33265) );
  IV U46185 ( .A(n33265), .Z(n36621) );
  XOR U46186 ( .A(n36622), .B(n36621), .Z(n33271) );
  NOR U46187 ( .A(n33266), .B(n33271), .Z(n33284) );
  IV U46188 ( .A(n33267), .Z(n33278) );
  NOR U46189 ( .A(n33269), .B(n33268), .Z(n33270) );
  IV U46190 ( .A(n33270), .Z(n33273) );
  IV U46191 ( .A(n33271), .Z(n33272) );
  NOR U46192 ( .A(n33273), .B(n33272), .Z(n33274) );
  IV U46193 ( .A(n33274), .Z(n33275) );
  NOR U46194 ( .A(n33276), .B(n33275), .Z(n33277) );
  IV U46195 ( .A(n33277), .Z(n33280) );
  NOR U46196 ( .A(n33278), .B(n33280), .Z(n38804) );
  IV U46197 ( .A(n33279), .Z(n33281) );
  NOR U46198 ( .A(n33281), .B(n33280), .Z(n38801) );
  NOR U46199 ( .A(n38804), .B(n38801), .Z(n33282) );
  IV U46200 ( .A(n33282), .Z(n33283) );
  NOR U46201 ( .A(n33284), .B(n33283), .Z(n35380) );
  XOR U46202 ( .A(n35382), .B(n35380), .Z(n36626) );
  XOR U46203 ( .A(n36625), .B(n36626), .Z(n36629) );
  XOR U46204 ( .A(n36628), .B(n36629), .Z(n36635) );
  XOR U46205 ( .A(n33285), .B(n36635), .Z(n33286) );
  IV U46206 ( .A(n33286), .Z(n36638) );
  XOR U46207 ( .A(n36636), .B(n36638), .Z(n35371) );
  NOR U46208 ( .A(n33287), .B(n35372), .Z(n33288) );
  XOR U46209 ( .A(n35371), .B(n33288), .Z(n35376) );
  IV U46210 ( .A(n33289), .Z(n33290) );
  NOR U46211 ( .A(n33290), .B(n33299), .Z(n35375) );
  IV U46212 ( .A(n33291), .Z(n33296) );
  NOR U46213 ( .A(n33293), .B(n33292), .Z(n33294) );
  IV U46214 ( .A(n33294), .Z(n33295) );
  NOR U46215 ( .A(n33296), .B(n33295), .Z(n35368) );
  NOR U46216 ( .A(n35375), .B(n35368), .Z(n33297) );
  XOR U46217 ( .A(n35376), .B(n33297), .Z(n36644) );
  IV U46218 ( .A(n33298), .Z(n33303) );
  NOR U46219 ( .A(n33300), .B(n33299), .Z(n33301) );
  IV U46220 ( .A(n33301), .Z(n33302) );
  NOR U46221 ( .A(n33303), .B(n33302), .Z(n33304) );
  IV U46222 ( .A(n33304), .Z(n36645) );
  XOR U46223 ( .A(n36644), .B(n36645), .Z(n36649) );
  XOR U46224 ( .A(n36647), .B(n36649), .Z(n38784) );
  XOR U46225 ( .A(n35367), .B(n38784), .Z(n36654) );
  IV U46226 ( .A(n33305), .Z(n33306) );
  NOR U46227 ( .A(n33307), .B(n33306), .Z(n33308) );
  NOR U46228 ( .A(n36653), .B(n33308), .Z(n36663) );
  XOR U46229 ( .A(n36654), .B(n36663), .Z(n36675) );
  XOR U46230 ( .A(n33309), .B(n36675), .Z(n33310) );
  IV U46231 ( .A(n33310), .Z(n36681) );
  XOR U46232 ( .A(n36679), .B(n36681), .Z(n35363) );
  XOR U46233 ( .A(n35362), .B(n35363), .Z(n35360) );
  XOR U46234 ( .A(n35359), .B(n35360), .Z(n38773) );
  IV U46235 ( .A(n38773), .Z(n33320) );
  IV U46236 ( .A(n33311), .Z(n33312) );
  NOR U46237 ( .A(n33312), .B(n33317), .Z(n36691) );
  IV U46238 ( .A(n33313), .Z(n33315) );
  NOR U46239 ( .A(n33315), .B(n33314), .Z(n40006) );
  IV U46240 ( .A(n33316), .Z(n33318) );
  NOR U46241 ( .A(n33318), .B(n33317), .Z(n38770) );
  NOR U46242 ( .A(n40006), .B(n38770), .Z(n36689) );
  IV U46243 ( .A(n36689), .Z(n36690) );
  NOR U46244 ( .A(n36691), .B(n36690), .Z(n33319) );
  XOR U46245 ( .A(n33320), .B(n33319), .Z(n36697) );
  XOR U46246 ( .A(n36696), .B(n36697), .Z(n36700) );
  XOR U46247 ( .A(n33321), .B(n36700), .Z(n35357) );
  NOR U46248 ( .A(n33322), .B(n35357), .Z(n43468) );
  IV U46249 ( .A(n33323), .Z(n33324) );
  NOR U46250 ( .A(n36701), .B(n33324), .Z(n33325) );
  IV U46251 ( .A(n33325), .Z(n35358) );
  XOR U46252 ( .A(n35358), .B(n35357), .Z(n33326) );
  NOR U46253 ( .A(n33327), .B(n33326), .Z(n36714) );
  NOR U46254 ( .A(n43468), .B(n36714), .Z(n36716) );
  XOR U46255 ( .A(n33328), .B(n36716), .Z(n36721) );
  XOR U46256 ( .A(n36719), .B(n36721), .Z(n36723) );
  XOR U46257 ( .A(n36722), .B(n36723), .Z(n33330) );
  NOR U46258 ( .A(n33334), .B(n33330), .Z(n38756) );
  IV U46259 ( .A(n33331), .Z(n33329) );
  NOR U46260 ( .A(n33329), .B(n36723), .Z(n38761) );
  NOR U46261 ( .A(n38756), .B(n38761), .Z(n36726) );
  IV U46262 ( .A(n36726), .Z(n33333) );
  IV U46263 ( .A(n33330), .Z(n33335) );
  NOR U46264 ( .A(n33331), .B(n33335), .Z(n33332) );
  NOR U46265 ( .A(n33333), .B(n33332), .Z(n33337) );
  NOR U46266 ( .A(n33335), .B(n33334), .Z(n33336) );
  NOR U46267 ( .A(n33337), .B(n33336), .Z(n35356) );
  XOR U46268 ( .A(n33338), .B(n35356), .Z(n35347) );
  XOR U46269 ( .A(n33339), .B(n35347), .Z(n35337) );
  XOR U46270 ( .A(n33340), .B(n35337), .Z(n36729) );
  NOR U46271 ( .A(n33341), .B(n36729), .Z(n38739) );
  IV U46272 ( .A(n33342), .Z(n33344) );
  NOR U46273 ( .A(n33344), .B(n33343), .Z(n36727) );
  XOR U46274 ( .A(n36729), .B(n36727), .Z(n35334) );
  NOR U46275 ( .A(n33346), .B(n33345), .Z(n33347) );
  IV U46276 ( .A(n33347), .Z(n33348) );
  NOR U46277 ( .A(n33349), .B(n33348), .Z(n33350) );
  IV U46278 ( .A(n33350), .Z(n35333) );
  XOR U46279 ( .A(n35334), .B(n35333), .Z(n33351) );
  NOR U46280 ( .A(n33352), .B(n33351), .Z(n33353) );
  NOR U46281 ( .A(n38739), .B(n33353), .Z(n35318) );
  XOR U46282 ( .A(n33354), .B(n35318), .Z(n36742) );
  XOR U46283 ( .A(n36740), .B(n36742), .Z(n36750) );
  IV U46284 ( .A(n36750), .Z(n33359) );
  IV U46285 ( .A(n33355), .Z(n33357) );
  NOR U46286 ( .A(n33357), .B(n33356), .Z(n36749) );
  NOR U46287 ( .A(n36743), .B(n36749), .Z(n33358) );
  XOR U46288 ( .A(n33359), .B(n33358), .Z(n36748) );
  IV U46289 ( .A(n33360), .Z(n33363) );
  IV U46290 ( .A(n33361), .Z(n33362) );
  NOR U46291 ( .A(n33363), .B(n33362), .Z(n36746) );
  XOR U46292 ( .A(n36748), .B(n36746), .Z(n36755) );
  XOR U46293 ( .A(n36753), .B(n36755), .Z(n36757) );
  XOR U46294 ( .A(n36756), .B(n36757), .Z(n35315) );
  XOR U46295 ( .A(n33364), .B(n35315), .Z(n33365) );
  IV U46296 ( .A(n33365), .Z(n36766) );
  XOR U46297 ( .A(n36764), .B(n36766), .Z(n35309) );
  IV U46298 ( .A(n33366), .Z(n33368) );
  NOR U46299 ( .A(n33368), .B(n33367), .Z(n35307) );
  XOR U46300 ( .A(n35309), .B(n35307), .Z(n36761) );
  XOR U46301 ( .A(n36760), .B(n36761), .Z(n38706) );
  IV U46302 ( .A(n38706), .Z(n33374) );
  IV U46303 ( .A(n33369), .Z(n33370) );
  NOR U46304 ( .A(n33373), .B(n33370), .Z(n38704) );
  IV U46305 ( .A(n33371), .Z(n33372) );
  NOR U46306 ( .A(n33373), .B(n33372), .Z(n38711) );
  NOR U46307 ( .A(n38704), .B(n38711), .Z(n36773) );
  XOR U46308 ( .A(n33374), .B(n36773), .Z(n35304) );
  XOR U46309 ( .A(n35303), .B(n35304), .Z(n35295) );
  XOR U46310 ( .A(n33375), .B(n35295), .Z(n36784) );
  XOR U46311 ( .A(n36783), .B(n36784), .Z(n36787) );
  NOR U46312 ( .A(n33383), .B(n36787), .Z(n36790) );
  IV U46313 ( .A(n33376), .Z(n33378) );
  NOR U46314 ( .A(n33378), .B(n33377), .Z(n33379) );
  IV U46315 ( .A(n33379), .Z(n36794) );
  IV U46316 ( .A(n33380), .Z(n33382) );
  NOR U46317 ( .A(n33382), .B(n33381), .Z(n36786) );
  XOR U46318 ( .A(n36786), .B(n36787), .Z(n36793) );
  XOR U46319 ( .A(n36794), .B(n36793), .Z(n33386) );
  IV U46320 ( .A(n36793), .Z(n33384) );
  NOR U46321 ( .A(n33384), .B(n33383), .Z(n33385) );
  NOR U46322 ( .A(n33386), .B(n33385), .Z(n33387) );
  NOR U46323 ( .A(n36790), .B(n33387), .Z(n33388) );
  IV U46324 ( .A(n33388), .Z(n35284) );
  XOR U46325 ( .A(n33389), .B(n35284), .Z(n35279) );
  XOR U46326 ( .A(n33390), .B(n35279), .Z(n36809) );
  XOR U46327 ( .A(n36800), .B(n36809), .Z(n36803) );
  XOR U46328 ( .A(n36802), .B(n36803), .Z(n35276) );
  XOR U46329 ( .A(n33391), .B(n35276), .Z(n33392) );
  IV U46330 ( .A(n33392), .Z(n35274) );
  XOR U46331 ( .A(n35272), .B(n35274), .Z(n36812) );
  XOR U46332 ( .A(n36811), .B(n36812), .Z(n36816) );
  IV U46333 ( .A(n33400), .Z(n33397) );
  NOR U46334 ( .A(n33394), .B(n33393), .Z(n33395) );
  IV U46335 ( .A(n33395), .Z(n33396) );
  NOR U46336 ( .A(n33397), .B(n33396), .Z(n36814) );
  XOR U46337 ( .A(n36816), .B(n36814), .Z(n35271) );
  IV U46338 ( .A(n33398), .Z(n33399) );
  NOR U46339 ( .A(n33400), .B(n33399), .Z(n35269) );
  XOR U46340 ( .A(n35271), .B(n35269), .Z(n35267) );
  XOR U46341 ( .A(n35266), .B(n35267), .Z(n35262) );
  IV U46342 ( .A(n33401), .Z(n33403) );
  NOR U46343 ( .A(n33403), .B(n33402), .Z(n35260) );
  XOR U46344 ( .A(n35262), .B(n35260), .Z(n35265) );
  NOR U46345 ( .A(n33404), .B(n35265), .Z(n38668) );
  IV U46346 ( .A(n33405), .Z(n33408) );
  IV U46347 ( .A(n33406), .Z(n33407) );
  NOR U46348 ( .A(n33408), .B(n33407), .Z(n35263) );
  XOR U46349 ( .A(n35265), .B(n35263), .Z(n33414) );
  IV U46350 ( .A(n33414), .Z(n33409) );
  NOR U46351 ( .A(n33410), .B(n33409), .Z(n33411) );
  NOR U46352 ( .A(n38668), .B(n33411), .Z(n33412) );
  NOR U46353 ( .A(n33413), .B(n33412), .Z(n33416) );
  IV U46354 ( .A(n33413), .Z(n33415) );
  NOR U46355 ( .A(n33415), .B(n33414), .Z(n38671) );
  NOR U46356 ( .A(n33416), .B(n38671), .Z(n33417) );
  IV U46357 ( .A(n33417), .Z(n36821) );
  XOR U46358 ( .A(n36820), .B(n36821), .Z(n42041) );
  IV U46359 ( .A(n42041), .Z(n33425) );
  IV U46360 ( .A(n33418), .Z(n33424) );
  NOR U46361 ( .A(n33420), .B(n33419), .Z(n33421) );
  NOR U46362 ( .A(n33421), .B(n36825), .Z(n33422) );
  IV U46363 ( .A(n33422), .Z(n33423) );
  NOR U46364 ( .A(n33424), .B(n33423), .Z(n42039) );
  NOR U46365 ( .A(n43580), .B(n42039), .Z(n35255) );
  XOR U46366 ( .A(n33425), .B(n35255), .Z(n35258) );
  XOR U46367 ( .A(n35256), .B(n35258), .Z(n36836) );
  XOR U46368 ( .A(n33426), .B(n36836), .Z(n33427) );
  IV U46369 ( .A(n33427), .Z(n35248) );
  XOR U46370 ( .A(n35246), .B(n35248), .Z(n36840) );
  IV U46371 ( .A(n36840), .Z(n33435) );
  IV U46372 ( .A(n33428), .Z(n33430) );
  NOR U46373 ( .A(n33430), .B(n33429), .Z(n35244) );
  IV U46374 ( .A(n33431), .Z(n33433) );
  NOR U46375 ( .A(n33433), .B(n33432), .Z(n36838) );
  NOR U46376 ( .A(n35244), .B(n36838), .Z(n33434) );
  XOR U46377 ( .A(n33435), .B(n33434), .Z(n36851) );
  XOR U46378 ( .A(n36850), .B(n36851), .Z(n33446) );
  IV U46379 ( .A(n33446), .Z(n33436) );
  NOR U46380 ( .A(n33437), .B(n33436), .Z(n40127) );
  IV U46381 ( .A(n33438), .Z(n33439) );
  NOR U46382 ( .A(n33440), .B(n33439), .Z(n33441) );
  IV U46383 ( .A(n33441), .Z(n36848) );
  IV U46384 ( .A(n33442), .Z(n33444) );
  NOR U46385 ( .A(n33444), .B(n33443), .Z(n33447) );
  IV U46386 ( .A(n33447), .Z(n33445) );
  NOR U46387 ( .A(n36851), .B(n33445), .Z(n35243) );
  NOR U46388 ( .A(n33447), .B(n33446), .Z(n33448) );
  NOR U46389 ( .A(n35243), .B(n33448), .Z(n33449) );
  IV U46390 ( .A(n33449), .Z(n36847) );
  XOR U46391 ( .A(n36848), .B(n36847), .Z(n33450) );
  NOR U46392 ( .A(n33451), .B(n33450), .Z(n33452) );
  NOR U46393 ( .A(n40127), .B(n33452), .Z(n35241) );
  XOR U46394 ( .A(n33453), .B(n35241), .Z(n35238) );
  XOR U46395 ( .A(n35237), .B(n35238), .Z(n35236) );
  IV U46396 ( .A(n35236), .Z(n33465) );
  IV U46397 ( .A(n33454), .Z(n33455) );
  NOR U46398 ( .A(n33455), .B(n33460), .Z(n33456) );
  IV U46399 ( .A(n33456), .Z(n33457) );
  NOR U46400 ( .A(n33458), .B(n33457), .Z(n35234) );
  IV U46401 ( .A(n33459), .Z(n33463) );
  NOR U46402 ( .A(n33461), .B(n33460), .Z(n33462) );
  IV U46403 ( .A(n33462), .Z(n33467) );
  NOR U46404 ( .A(n33463), .B(n33467), .Z(n35232) );
  NOR U46405 ( .A(n35234), .B(n35232), .Z(n33464) );
  XOR U46406 ( .A(n33465), .B(n33464), .Z(n36873) );
  IV U46407 ( .A(n33466), .Z(n33468) );
  NOR U46408 ( .A(n33468), .B(n33467), .Z(n36871) );
  XOR U46409 ( .A(n36873), .B(n36871), .Z(n36876) );
  XOR U46410 ( .A(n33469), .B(n36876), .Z(n35230) );
  XOR U46411 ( .A(n33470), .B(n35230), .Z(n35222) );
  IV U46412 ( .A(n33471), .Z(n33473) );
  NOR U46413 ( .A(n33473), .B(n33472), .Z(n35226) );
  IV U46414 ( .A(n33474), .Z(n33478) );
  XOR U46415 ( .A(n33476), .B(n33475), .Z(n33477) );
  NOR U46416 ( .A(n33478), .B(n33477), .Z(n35221) );
  NOR U46417 ( .A(n35226), .B(n35221), .Z(n33479) );
  XOR U46418 ( .A(n35222), .B(n33479), .Z(n36888) );
  XOR U46419 ( .A(n36887), .B(n36888), .Z(n36898) );
  XOR U46420 ( .A(n33480), .B(n36898), .Z(n33481) );
  IV U46421 ( .A(n33481), .Z(n36895) );
  XOR U46422 ( .A(n36893), .B(n36895), .Z(n36902) );
  IV U46423 ( .A(n36902), .Z(n33489) );
  IV U46424 ( .A(n33482), .Z(n35217) );
  NOR U46425 ( .A(n33492), .B(n35217), .Z(n33487) );
  IV U46426 ( .A(n33483), .Z(n33491) );
  NOR U46427 ( .A(n33484), .B(n33491), .Z(n33485) );
  IV U46428 ( .A(n33485), .Z(n33486) );
  NOR U46429 ( .A(n33492), .B(n33486), .Z(n36900) );
  NOR U46430 ( .A(n33487), .B(n36900), .Z(n33488) );
  XOR U46431 ( .A(n33489), .B(n33488), .Z(n35216) );
  IV U46432 ( .A(n33490), .Z(n33495) );
  NOR U46433 ( .A(n33492), .B(n33491), .Z(n33493) );
  IV U46434 ( .A(n33493), .Z(n33494) );
  NOR U46435 ( .A(n33495), .B(n33494), .Z(n35214) );
  XOR U46436 ( .A(n35216), .B(n35214), .Z(n36905) );
  XOR U46437 ( .A(n36903), .B(n36905), .Z(n36912) );
  XOR U46438 ( .A(n36906), .B(n36912), .Z(n35213) );
  XOR U46439 ( .A(n33496), .B(n35213), .Z(n33497) );
  IV U46440 ( .A(n33497), .Z(n35210) );
  XOR U46441 ( .A(n35208), .B(n35210), .Z(n36915) );
  XOR U46442 ( .A(n36914), .B(n36915), .Z(n35207) );
  IV U46443 ( .A(n33498), .Z(n33505) );
  XOR U46444 ( .A(n33500), .B(n33499), .Z(n33501) );
  NOR U46445 ( .A(n33502), .B(n33501), .Z(n33503) );
  IV U46446 ( .A(n33503), .Z(n33504) );
  NOR U46447 ( .A(n33505), .B(n33504), .Z(n35205) );
  XOR U46448 ( .A(n35207), .B(n35205), .Z(n36932) );
  IV U46449 ( .A(n36932), .Z(n33516) );
  IV U46450 ( .A(n33506), .Z(n33508) );
  NOR U46451 ( .A(n33508), .B(n33507), .Z(n36931) );
  IV U46452 ( .A(n33509), .Z(n33514) );
  NOR U46453 ( .A(n33511), .B(n33510), .Z(n33512) );
  IV U46454 ( .A(n33512), .Z(n33513) );
  NOR U46455 ( .A(n33514), .B(n33513), .Z(n35203) );
  NOR U46456 ( .A(n36931), .B(n35203), .Z(n33515) );
  XOR U46457 ( .A(n33516), .B(n33515), .Z(n35202) );
  XOR U46458 ( .A(n35201), .B(n35202), .Z(n33521) );
  IV U46459 ( .A(n33517), .Z(n33518) );
  NOR U46460 ( .A(n33518), .B(n33523), .Z(n33519) );
  NOR U46461 ( .A(n33521), .B(n33519), .Z(n33534) );
  IV U46462 ( .A(n33520), .Z(n33528) );
  IV U46463 ( .A(n33521), .Z(n33522) );
  NOR U46464 ( .A(n33523), .B(n33522), .Z(n33524) );
  IV U46465 ( .A(n33524), .Z(n33525) );
  NOR U46466 ( .A(n33526), .B(n33525), .Z(n33527) );
  IV U46467 ( .A(n33527), .Z(n33530) );
  NOR U46468 ( .A(n33528), .B(n33530), .Z(n40201) );
  IV U46469 ( .A(n33529), .Z(n33531) );
  NOR U46470 ( .A(n33531), .B(n33530), .Z(n40197) );
  NOR U46471 ( .A(n40201), .B(n40197), .Z(n33532) );
  IV U46472 ( .A(n33532), .Z(n33533) );
  NOR U46473 ( .A(n33534), .B(n33533), .Z(n33535) );
  IV U46474 ( .A(n33535), .Z(n35199) );
  IV U46475 ( .A(n33536), .Z(n33538) );
  NOR U46476 ( .A(n33538), .B(n33537), .Z(n35197) );
  XOR U46477 ( .A(n35199), .B(n35197), .Z(n36940) );
  XOR U46478 ( .A(n36939), .B(n36940), .Z(n35194) );
  XOR U46479 ( .A(n35193), .B(n35194), .Z(n36936) );
  XOR U46480 ( .A(n36935), .B(n36936), .Z(n36953) );
  XOR U46481 ( .A(n36952), .B(n36953), .Z(n35188) );
  XOR U46482 ( .A(n35187), .B(n35188), .Z(n35191) );
  XOR U46483 ( .A(n35190), .B(n35191), .Z(n41943) );
  XOR U46484 ( .A(n35183), .B(n41943), .Z(n35184) );
  IV U46485 ( .A(n33539), .Z(n33540) );
  NOR U46486 ( .A(n33547), .B(n33540), .Z(n33541) );
  IV U46487 ( .A(n33541), .Z(n33542) );
  NOR U46488 ( .A(n33543), .B(n33542), .Z(n33544) );
  IV U46489 ( .A(n33544), .Z(n35185) );
  XOR U46490 ( .A(n35184), .B(n35185), .Z(n36961) );
  IV U46491 ( .A(n33545), .Z(n33549) );
  NOR U46492 ( .A(n33547), .B(n33546), .Z(n33548) );
  IV U46493 ( .A(n33548), .Z(n33551) );
  NOR U46494 ( .A(n33549), .B(n33551), .Z(n36959) );
  XOR U46495 ( .A(n36961), .B(n36959), .Z(n35182) );
  IV U46496 ( .A(n33550), .Z(n33552) );
  NOR U46497 ( .A(n33552), .B(n33551), .Z(n35180) );
  XOR U46498 ( .A(n35182), .B(n35180), .Z(n36973) );
  IV U46499 ( .A(n33553), .Z(n33555) );
  NOR U46500 ( .A(n33555), .B(n33554), .Z(n36971) );
  XOR U46501 ( .A(n36973), .B(n36971), .Z(n36975) );
  XOR U46502 ( .A(n36974), .B(n36975), .Z(n36980) );
  IV U46503 ( .A(n36980), .Z(n33565) );
  IV U46504 ( .A(n33556), .Z(n33558) );
  NOR U46505 ( .A(n33558), .B(n33557), .Z(n35178) );
  NOR U46506 ( .A(n33560), .B(n33559), .Z(n33561) );
  IV U46507 ( .A(n33561), .Z(n33562) );
  NOR U46508 ( .A(n33563), .B(n33562), .Z(n36978) );
  NOR U46509 ( .A(n35178), .B(n36978), .Z(n33564) );
  XOR U46510 ( .A(n33565), .B(n33564), .Z(n35174) );
  XOR U46511 ( .A(n35172), .B(n35174), .Z(n35176) );
  XOR U46512 ( .A(n35175), .B(n35176), .Z(n35167) );
  XOR U46513 ( .A(n35166), .B(n35167), .Z(n35170) );
  XOR U46514 ( .A(n33566), .B(n35170), .Z(n35154) );
  XOR U46515 ( .A(n33567), .B(n35154), .Z(n33568) );
  XOR U46516 ( .A(n33569), .B(n33568), .Z(n36990) );
  IV U46517 ( .A(n36990), .Z(n33574) );
  IV U46518 ( .A(n33570), .Z(n36996) );
  NOR U46519 ( .A(n36996), .B(n33571), .Z(n33572) );
  NOR U46520 ( .A(n36991), .B(n33572), .Z(n33573) );
  XOR U46521 ( .A(n33574), .B(n33573), .Z(n35152) );
  XOR U46522 ( .A(n35150), .B(n35152), .Z(n35146) );
  XOR U46523 ( .A(n35145), .B(n35146), .Z(n36999) );
  IV U46524 ( .A(n36999), .Z(n33578) );
  NOR U46525 ( .A(n33576), .B(n33575), .Z(n36998) );
  NOR U46526 ( .A(n35148), .B(n36998), .Z(n33577) );
  XOR U46527 ( .A(n33578), .B(n33577), .Z(n37003) );
  IV U46528 ( .A(n33579), .Z(n33581) );
  NOR U46529 ( .A(n33581), .B(n33580), .Z(n37001) );
  XOR U46530 ( .A(n37003), .B(n37001), .Z(n37006) );
  XOR U46531 ( .A(n37004), .B(n37006), .Z(n37017) );
  XOR U46532 ( .A(n37016), .B(n37017), .Z(n37009) );
  XOR U46533 ( .A(n37008), .B(n37009), .Z(n37013) );
  XOR U46534 ( .A(n37012), .B(n37013), .Z(n35144) );
  IV U46535 ( .A(n33582), .Z(n33587) );
  IV U46536 ( .A(n33583), .Z(n33584) );
  NOR U46537 ( .A(n33585), .B(n33584), .Z(n33586) );
  IV U46538 ( .A(n33586), .Z(n33590) );
  NOR U46539 ( .A(n33587), .B(n33590), .Z(n33593) );
  IV U46540 ( .A(n33593), .Z(n33588) );
  NOR U46541 ( .A(n35144), .B(n33588), .Z(n38572) );
  IV U46542 ( .A(n33589), .Z(n33591) );
  NOR U46543 ( .A(n33591), .B(n33590), .Z(n33592) );
  IV U46544 ( .A(n33592), .Z(n35143) );
  XOR U46545 ( .A(n35143), .B(n35144), .Z(n33598) );
  NOR U46546 ( .A(n33593), .B(n33598), .Z(n33594) );
  NOR U46547 ( .A(n38572), .B(n33594), .Z(n35139) );
  IV U46548 ( .A(n33595), .Z(n33597) );
  NOR U46549 ( .A(n33597), .B(n33596), .Z(n33608) );
  IV U46550 ( .A(n33608), .Z(n35140) );
  NOR U46551 ( .A(n35139), .B(n35140), .Z(n33610) );
  IV U46552 ( .A(n33598), .Z(n33603) );
  IV U46553 ( .A(n33599), .Z(n33600) );
  NOR U46554 ( .A(n33601), .B(n33600), .Z(n33604) );
  IV U46555 ( .A(n33604), .Z(n33602) );
  NOR U46556 ( .A(n33603), .B(n33602), .Z(n43723) );
  NOR U46557 ( .A(n35139), .B(n33604), .Z(n33605) );
  NOR U46558 ( .A(n43723), .B(n33605), .Z(n33606) );
  IV U46559 ( .A(n33606), .Z(n33607) );
  NOR U46560 ( .A(n33608), .B(n33607), .Z(n33609) );
  NOR U46561 ( .A(n33610), .B(n33609), .Z(n35132) );
  XOR U46562 ( .A(n35131), .B(n35132), .Z(n35136) );
  XOR U46563 ( .A(n33611), .B(n35136), .Z(n37030) );
  XOR U46564 ( .A(n37029), .B(n37030), .Z(n37034) );
  XOR U46565 ( .A(n37032), .B(n37034), .Z(n35128) );
  XOR U46566 ( .A(n33612), .B(n35128), .Z(n33622) );
  IV U46567 ( .A(n33622), .Z(n33613) );
  NOR U46568 ( .A(n33627), .B(n33613), .Z(n43743) );
  IV U46569 ( .A(n33614), .Z(n33615) );
  NOR U46570 ( .A(n33616), .B(n33615), .Z(n33629) );
  IV U46571 ( .A(n33629), .Z(n33626) );
  IV U46572 ( .A(n33617), .Z(n33619) );
  NOR U46573 ( .A(n33619), .B(n33618), .Z(n33623) );
  IV U46574 ( .A(n33623), .Z(n33621) );
  XOR U46575 ( .A(n35118), .B(n35128), .Z(n33620) );
  NOR U46576 ( .A(n33621), .B(n33620), .Z(n40305) );
  NOR U46577 ( .A(n33623), .B(n33622), .Z(n33624) );
  NOR U46578 ( .A(n40305), .B(n33624), .Z(n33628) );
  IV U46579 ( .A(n33628), .Z(n33625) );
  NOR U46580 ( .A(n33626), .B(n33625), .Z(n43749) );
  NOR U46581 ( .A(n43743), .B(n43749), .Z(n38571) );
  IV U46582 ( .A(n38571), .Z(n37042) );
  NOR U46583 ( .A(n37042), .B(n33627), .Z(n33632) );
  NOR U46584 ( .A(n33629), .B(n33628), .Z(n33630) );
  NOR U46585 ( .A(n33630), .B(n37042), .Z(n33631) );
  NOR U46586 ( .A(n33632), .B(n33631), .Z(n35111) );
  XOR U46587 ( .A(n35110), .B(n35111), .Z(n35113) );
  XOR U46588 ( .A(n35114), .B(n35113), .Z(n33640) );
  IV U46589 ( .A(n33640), .Z(n33633) );
  NOR U46590 ( .A(n33634), .B(n33633), .Z(n33635) );
  IV U46591 ( .A(n33635), .Z(n33636) );
  NOR U46592 ( .A(n33638), .B(n33636), .Z(n40314) );
  NOR U46593 ( .A(n33638), .B(n33637), .Z(n33639) );
  NOR U46594 ( .A(n33640), .B(n33639), .Z(n33641) );
  NOR U46595 ( .A(n40314), .B(n33641), .Z(n33642) );
  IV U46596 ( .A(n33642), .Z(n37045) );
  IV U46597 ( .A(n33643), .Z(n33645) );
  NOR U46598 ( .A(n33645), .B(n33644), .Z(n37043) );
  XOR U46599 ( .A(n37045), .B(n37043), .Z(n35103) );
  XOR U46600 ( .A(n35102), .B(n35103), .Z(n37051) );
  XOR U46601 ( .A(n33646), .B(n37051), .Z(n37048) );
  NOR U46602 ( .A(n33647), .B(n37048), .Z(n41846) );
  XOR U46603 ( .A(n37047), .B(n37048), .Z(n37055) );
  IV U46604 ( .A(n33648), .Z(n33660) );
  NOR U46605 ( .A(n33660), .B(n33649), .Z(n35100) );
  NOR U46606 ( .A(n37054), .B(n35100), .Z(n33650) );
  XOR U46607 ( .A(n37055), .B(n33650), .Z(n33651) );
  NOR U46608 ( .A(n33652), .B(n33651), .Z(n33653) );
  NOR U46609 ( .A(n41846), .B(n33653), .Z(n35094) );
  IV U46610 ( .A(n33664), .Z(n33657) );
  NOR U46611 ( .A(n33654), .B(n33660), .Z(n33655) );
  IV U46612 ( .A(n33655), .Z(n33656) );
  NOR U46613 ( .A(n33657), .B(n33656), .Z(n33658) );
  IV U46614 ( .A(n33658), .Z(n35095) );
  XOR U46615 ( .A(n35094), .B(n35095), .Z(n35092) );
  IV U46616 ( .A(n35092), .Z(n33674) );
  IV U46617 ( .A(n33659), .Z(n33661) );
  NOR U46618 ( .A(n33661), .B(n33660), .Z(n33662) );
  IV U46619 ( .A(n33662), .Z(n33663) );
  NOR U46620 ( .A(n33664), .B(n33663), .Z(n35096) );
  IV U46621 ( .A(n33665), .Z(n33667) );
  NOR U46622 ( .A(n33667), .B(n33666), .Z(n35091) );
  IV U46623 ( .A(n33668), .Z(n33670) );
  NOR U46624 ( .A(n33670), .B(n33669), .Z(n35089) );
  NOR U46625 ( .A(n35091), .B(n35089), .Z(n33671) );
  IV U46626 ( .A(n33671), .Z(n33672) );
  NOR U46627 ( .A(n35096), .B(n33672), .Z(n33673) );
  XOR U46628 ( .A(n33674), .B(n33673), .Z(n35088) );
  IV U46629 ( .A(n33675), .Z(n33677) );
  NOR U46630 ( .A(n33677), .B(n33676), .Z(n35086) );
  XOR U46631 ( .A(n35088), .B(n35086), .Z(n37069) );
  XOR U46632 ( .A(n37068), .B(n37069), .Z(n37072) );
  XOR U46633 ( .A(n33678), .B(n37072), .Z(n35082) );
  XOR U46634 ( .A(n35080), .B(n35082), .Z(n35084) );
  XOR U46635 ( .A(n35083), .B(n35084), .Z(n35078) );
  XOR U46636 ( .A(n33679), .B(n35078), .Z(n35071) );
  XOR U46637 ( .A(n33680), .B(n35071), .Z(n37087) );
  IV U46638 ( .A(n33681), .Z(n33683) );
  NOR U46639 ( .A(n33683), .B(n33682), .Z(n37084) );
  NOR U46640 ( .A(n37084), .B(n37086), .Z(n33684) );
  XOR U46641 ( .A(n37087), .B(n33684), .Z(n37096) );
  NOR U46642 ( .A(n33686), .B(n33685), .Z(n37094) );
  IV U46643 ( .A(n33687), .Z(n33689) );
  NOR U46644 ( .A(n33689), .B(n33688), .Z(n37092) );
  NOR U46645 ( .A(n37094), .B(n37092), .Z(n33690) );
  XOR U46646 ( .A(n37096), .B(n33690), .Z(n35066) );
  IV U46647 ( .A(n33691), .Z(n33693) );
  NOR U46648 ( .A(n33693), .B(n33692), .Z(n37103) );
  NOR U46649 ( .A(n35065), .B(n37103), .Z(n33694) );
  XOR U46650 ( .A(n35066), .B(n33694), .Z(n37108) );
  IV U46651 ( .A(n33695), .Z(n33696) );
  NOR U46652 ( .A(n37107), .B(n33696), .Z(n33697) );
  XOR U46653 ( .A(n37108), .B(n33697), .Z(n35059) );
  NOR U46654 ( .A(n33698), .B(n35058), .Z(n33699) );
  XOR U46655 ( .A(n35059), .B(n33699), .Z(n35056) );
  IV U46656 ( .A(n33700), .Z(n33701) );
  NOR U46657 ( .A(n33703), .B(n33701), .Z(n35054) );
  IV U46658 ( .A(n33702), .Z(n33706) );
  NOR U46659 ( .A(n33704), .B(n33703), .Z(n33705) );
  IV U46660 ( .A(n33705), .Z(n33710) );
  NOR U46661 ( .A(n33706), .B(n33710), .Z(n35052) );
  NOR U46662 ( .A(n35054), .B(n35052), .Z(n33707) );
  XOR U46663 ( .A(n35056), .B(n33707), .Z(n33708) );
  IV U46664 ( .A(n33708), .Z(n35048) );
  IV U46665 ( .A(n33709), .Z(n33711) );
  NOR U46666 ( .A(n33711), .B(n33710), .Z(n35046) );
  XOR U46667 ( .A(n35048), .B(n35046), .Z(n35051) );
  IV U46668 ( .A(n35051), .Z(n33718) );
  NOR U46669 ( .A(n33713), .B(n33712), .Z(n35044) );
  IV U46670 ( .A(n33714), .Z(n33715) );
  NOR U46671 ( .A(n33716), .B(n33715), .Z(n35049) );
  NOR U46672 ( .A(n35044), .B(n35049), .Z(n33717) );
  XOR U46673 ( .A(n33718), .B(n33717), .Z(n35043) );
  XOR U46674 ( .A(n35041), .B(n35043), .Z(n35037) );
  XOR U46675 ( .A(n35027), .B(n35037), .Z(n35025) );
  IV U46676 ( .A(n33719), .Z(n35030) );
  IV U46677 ( .A(n33720), .Z(n33721) );
  NOR U46678 ( .A(n35030), .B(n33721), .Z(n33722) );
  XOR U46679 ( .A(n35025), .B(n33722), .Z(n37128) );
  IV U46680 ( .A(n33723), .Z(n33724) );
  NOR U46681 ( .A(n33725), .B(n33724), .Z(n35023) );
  IV U46682 ( .A(n33726), .Z(n33729) );
  IV U46683 ( .A(n33727), .Z(n33728) );
  NOR U46684 ( .A(n33729), .B(n33728), .Z(n37126) );
  NOR U46685 ( .A(n35023), .B(n37126), .Z(n33730) );
  XOR U46686 ( .A(n37128), .B(n33730), .Z(n35021) );
  IV U46687 ( .A(n33731), .Z(n33733) );
  NOR U46688 ( .A(n33733), .B(n33732), .Z(n35020) );
  IV U46689 ( .A(n33734), .Z(n33735) );
  NOR U46690 ( .A(n33735), .B(n33739), .Z(n37132) );
  NOR U46691 ( .A(n35020), .B(n37132), .Z(n33736) );
  XOR U46692 ( .A(n35021), .B(n33736), .Z(n37131) );
  IV U46693 ( .A(n33737), .Z(n33738) );
  NOR U46694 ( .A(n33739), .B(n33738), .Z(n37129) );
  XOR U46695 ( .A(n37131), .B(n37129), .Z(n37137) );
  XOR U46696 ( .A(n37136), .B(n37137), .Z(n37140) );
  XOR U46697 ( .A(n33740), .B(n37140), .Z(n33741) );
  IV U46698 ( .A(n33741), .Z(n37145) );
  XOR U46699 ( .A(n37143), .B(n37145), .Z(n37147) );
  XOR U46700 ( .A(n37146), .B(n37147), .Z(n35016) );
  XOR U46701 ( .A(n35015), .B(n35016), .Z(n35011) );
  IV U46702 ( .A(n33742), .Z(n33744) );
  NOR U46703 ( .A(n33744), .B(n33743), .Z(n35009) );
  XOR U46704 ( .A(n35011), .B(n35009), .Z(n35013) );
  XOR U46705 ( .A(n35012), .B(n35013), .Z(n37153) );
  XOR U46706 ( .A(n37152), .B(n37153), .Z(n37156) );
  IV U46707 ( .A(n33745), .Z(n33746) );
  NOR U46708 ( .A(n33747), .B(n33746), .Z(n37155) );
  IV U46709 ( .A(n33748), .Z(n33750) );
  NOR U46710 ( .A(n33750), .B(n33749), .Z(n35004) );
  NOR U46711 ( .A(n37155), .B(n35004), .Z(n33751) );
  XOR U46712 ( .A(n37156), .B(n33751), .Z(n35007) );
  XOR U46713 ( .A(n33752), .B(n35007), .Z(n38488) );
  XOR U46714 ( .A(n33753), .B(n38488), .Z(n34999) );
  XOR U46715 ( .A(n34998), .B(n34999), .Z(n35002) );
  XOR U46716 ( .A(n35001), .B(n35002), .Z(n37168) );
  XOR U46717 ( .A(n33754), .B(n37168), .Z(n33755) );
  IV U46718 ( .A(n33755), .Z(n34990) );
  XOR U46719 ( .A(n33756), .B(n34990), .Z(n37177) );
  XOR U46720 ( .A(n37175), .B(n37177), .Z(n37183) );
  XOR U46721 ( .A(n37182), .B(n37183), .Z(n34981) );
  XOR U46722 ( .A(n33757), .B(n34981), .Z(n37189) );
  NOR U46723 ( .A(n33759), .B(n33758), .Z(n34978) );
  NOR U46724 ( .A(n37188), .B(n34978), .Z(n33760) );
  XOR U46725 ( .A(n37189), .B(n33760), .Z(n34970) );
  NOR U46726 ( .A(n33761), .B(n34971), .Z(n33762) );
  NOR U46727 ( .A(n34975), .B(n33762), .Z(n33763) );
  XOR U46728 ( .A(n34970), .B(n33763), .Z(n34968) );
  XOR U46729 ( .A(n34967), .B(n34968), .Z(n34963) );
  IV U46730 ( .A(n33764), .Z(n33765) );
  NOR U46731 ( .A(n33766), .B(n33765), .Z(n34962) );
  IV U46732 ( .A(n33767), .Z(n33769) );
  NOR U46733 ( .A(n33769), .B(n33768), .Z(n37191) );
  NOR U46734 ( .A(n34962), .B(n37191), .Z(n33770) );
  NOR U46735 ( .A(n33770), .B(n34964), .Z(n33771) );
  XOR U46736 ( .A(n34963), .B(n33771), .Z(n34960) );
  XOR U46737 ( .A(n34959), .B(n34960), .Z(n34956) );
  IV U46738 ( .A(n33772), .Z(n33786) );
  NOR U46739 ( .A(n33786), .B(n33773), .Z(n33774) );
  IV U46740 ( .A(n33774), .Z(n34955) );
  NOR U46741 ( .A(n33775), .B(n34955), .Z(n33776) );
  XOR U46742 ( .A(n34956), .B(n33776), .Z(n37199) );
  IV U46743 ( .A(n33777), .Z(n33778) );
  NOR U46744 ( .A(n33778), .B(n33782), .Z(n33779) );
  IV U46745 ( .A(n33779), .Z(n33780) );
  NOR U46746 ( .A(n33786), .B(n33780), .Z(n37197) );
  XOR U46747 ( .A(n37199), .B(n37197), .Z(n37202) );
  IV U46748 ( .A(n33781), .Z(n33783) );
  NOR U46749 ( .A(n33783), .B(n33782), .Z(n33784) );
  IV U46750 ( .A(n33784), .Z(n33785) );
  NOR U46751 ( .A(n33786), .B(n33785), .Z(n37200) );
  XOR U46752 ( .A(n37202), .B(n37200), .Z(n34952) );
  IV U46753 ( .A(n33787), .Z(n33789) );
  NOR U46754 ( .A(n33789), .B(n33788), .Z(n34951) );
  IV U46755 ( .A(n33790), .Z(n33792) );
  NOR U46756 ( .A(n33792), .B(n33791), .Z(n34949) );
  NOR U46757 ( .A(n34951), .B(n34949), .Z(n33793) );
  XOR U46758 ( .A(n34952), .B(n33793), .Z(n34944) );
  XOR U46759 ( .A(n33794), .B(n34944), .Z(n34934) );
  XOR U46760 ( .A(n33795), .B(n34934), .Z(n34928) );
  XOR U46761 ( .A(n34926), .B(n34928), .Z(n34930) );
  XOR U46762 ( .A(n34929), .B(n34930), .Z(n34924) );
  NOR U46763 ( .A(n33797), .B(n33796), .Z(n34923) );
  IV U46764 ( .A(n33798), .Z(n33800) );
  NOR U46765 ( .A(n33800), .B(n33799), .Z(n34921) );
  NOR U46766 ( .A(n34923), .B(n34921), .Z(n33801) );
  XOR U46767 ( .A(n34924), .B(n33801), .Z(n37207) );
  XOR U46768 ( .A(n33802), .B(n37207), .Z(n34920) );
  XOR U46769 ( .A(n34919), .B(n34920), .Z(n33805) );
  NOR U46770 ( .A(n33803), .B(n34912), .Z(n33804) );
  XOR U46771 ( .A(n33805), .B(n33804), .Z(n34905) );
  IV U46772 ( .A(n33806), .Z(n33807) );
  NOR U46773 ( .A(n33807), .B(n34912), .Z(n33808) );
  IV U46774 ( .A(n33808), .Z(n34906) );
  XOR U46775 ( .A(n34905), .B(n34906), .Z(n34909) );
  IV U46776 ( .A(n34909), .Z(n34899) );
  IV U46777 ( .A(n33809), .Z(n33813) );
  IV U46778 ( .A(n33810), .Z(n33811) );
  NOR U46779 ( .A(n33813), .B(n33811), .Z(n34900) );
  NOR U46780 ( .A(n33813), .B(n33812), .Z(n34896) );
  IV U46781 ( .A(n33814), .Z(n33815) );
  NOR U46782 ( .A(n33816), .B(n33815), .Z(n34903) );
  NOR U46783 ( .A(n34908), .B(n34903), .Z(n33817) );
  IV U46784 ( .A(n33817), .Z(n33818) );
  NOR U46785 ( .A(n34896), .B(n33818), .Z(n34898) );
  IV U46786 ( .A(n34898), .Z(n33819) );
  NOR U46787 ( .A(n34900), .B(n33819), .Z(n33820) );
  XOR U46788 ( .A(n34899), .B(n33820), .Z(n34892) );
  XOR U46789 ( .A(n34890), .B(n34892), .Z(n34894) );
  XOR U46790 ( .A(n34893), .B(n34894), .Z(n37225) );
  IV U46791 ( .A(n37225), .Z(n33821) );
  NOR U46792 ( .A(n33822), .B(n33821), .Z(n33832) );
  IV U46793 ( .A(n33823), .Z(n33826) );
  NOR U46794 ( .A(n33824), .B(n34894), .Z(n33825) );
  IV U46795 ( .A(n33825), .Z(n33828) );
  NOR U46796 ( .A(n33826), .B(n33828), .Z(n40508) );
  IV U46797 ( .A(n33827), .Z(n33829) );
  NOR U46798 ( .A(n33829), .B(n33828), .Z(n38430) );
  NOR U46799 ( .A(n40508), .B(n38430), .Z(n33830) );
  IV U46800 ( .A(n33830), .Z(n33831) );
  NOR U46801 ( .A(n33832), .B(n33831), .Z(n33833) );
  IV U46802 ( .A(n33833), .Z(n37231) );
  XOR U46803 ( .A(n33834), .B(n37231), .Z(n37228) );
  IV U46804 ( .A(n33835), .Z(n33836) );
  NOR U46805 ( .A(n33837), .B(n33836), .Z(n40527) );
  IV U46806 ( .A(n33838), .Z(n33839) );
  NOR U46807 ( .A(n33840), .B(n33839), .Z(n40513) );
  NOR U46808 ( .A(n40527), .B(n40513), .Z(n37229) );
  XOR U46809 ( .A(n37228), .B(n37229), .Z(n34885) );
  XOR U46810 ( .A(n34884), .B(n34885), .Z(n34889) );
  IV U46811 ( .A(n33841), .Z(n33842) );
  NOR U46812 ( .A(n33842), .B(n33846), .Z(n34887) );
  XOR U46813 ( .A(n34889), .B(n34887), .Z(n40535) );
  IV U46814 ( .A(n40535), .Z(n33848) );
  NOR U46815 ( .A(n33844), .B(n33843), .Z(n40542) );
  IV U46816 ( .A(n33845), .Z(n33847) );
  NOR U46817 ( .A(n33847), .B(n33846), .Z(n40534) );
  NOR U46818 ( .A(n40542), .B(n40534), .Z(n34883) );
  XOR U46819 ( .A(n33848), .B(n34883), .Z(n34878) );
  XOR U46820 ( .A(n34877), .B(n34878), .Z(n34882) );
  XOR U46821 ( .A(n34880), .B(n34882), .Z(n37242) );
  XOR U46822 ( .A(n37240), .B(n37242), .Z(n34869) );
  XOR U46823 ( .A(n34868), .B(n34869), .Z(n34866) );
  NOR U46824 ( .A(n33855), .B(n34866), .Z(n40560) );
  IV U46825 ( .A(n33849), .Z(n33851) );
  NOR U46826 ( .A(n33851), .B(n33850), .Z(n34865) );
  XOR U46827 ( .A(n34865), .B(n34866), .Z(n37249) );
  IV U46828 ( .A(n33852), .Z(n33854) );
  NOR U46829 ( .A(n33854), .B(n33853), .Z(n33856) );
  IV U46830 ( .A(n33856), .Z(n37248) );
  XOR U46831 ( .A(n37249), .B(n37248), .Z(n33858) );
  NOR U46832 ( .A(n33856), .B(n33855), .Z(n33857) );
  NOR U46833 ( .A(n33858), .B(n33857), .Z(n33859) );
  NOR U46834 ( .A(n40560), .B(n33859), .Z(n37250) );
  XOR U46835 ( .A(n37252), .B(n37250), .Z(n37255) );
  XOR U46836 ( .A(n37254), .B(n37255), .Z(n37262) );
  XOR U46837 ( .A(n33860), .B(n37262), .Z(n33861) );
  IV U46838 ( .A(n33861), .Z(n34862) );
  XOR U46839 ( .A(n34860), .B(n34862), .Z(n37264) );
  IV U46840 ( .A(n33862), .Z(n33864) );
  NOR U46841 ( .A(n33864), .B(n33863), .Z(n34863) );
  IV U46842 ( .A(n33865), .Z(n33867) );
  NOR U46843 ( .A(n33867), .B(n33866), .Z(n37263) );
  NOR U46844 ( .A(n34863), .B(n37263), .Z(n33868) );
  XOR U46845 ( .A(n37264), .B(n33868), .Z(n37266) );
  NOR U46846 ( .A(n33870), .B(n33869), .Z(n37267) );
  NOR U46847 ( .A(n37270), .B(n37267), .Z(n33871) );
  XOR U46848 ( .A(n37266), .B(n33871), .Z(n34851) );
  XOR U46849 ( .A(n34850), .B(n34851), .Z(n37278) );
  XOR U46850 ( .A(n37277), .B(n37278), .Z(n37275) );
  XOR U46851 ( .A(n37274), .B(n37275), .Z(n34846) );
  IV U46852 ( .A(n33872), .Z(n33874) );
  NOR U46853 ( .A(n33874), .B(n33873), .Z(n34848) );
  IV U46854 ( .A(n33875), .Z(n33876) );
  NOR U46855 ( .A(n33879), .B(n33876), .Z(n34845) );
  NOR U46856 ( .A(n34848), .B(n34845), .Z(n33877) );
  XOR U46857 ( .A(n34846), .B(n33877), .Z(n33878) );
  IV U46858 ( .A(n33878), .Z(n34842) );
  NOR U46859 ( .A(n33880), .B(n33879), .Z(n33881) );
  IV U46860 ( .A(n33881), .Z(n34841) );
  NOR U46861 ( .A(n33882), .B(n34841), .Z(n33883) );
  XOR U46862 ( .A(n34842), .B(n33883), .Z(n34838) );
  XOR U46863 ( .A(n34836), .B(n34838), .Z(n34833) );
  NOR U46864 ( .A(n33884), .B(n34833), .Z(n33885) );
  IV U46865 ( .A(n33885), .Z(n41628) );
  NOR U46866 ( .A(n33887), .B(n41628), .Z(n38389) );
  IV U46867 ( .A(n33886), .Z(n33889) );
  NOR U46868 ( .A(n33889), .B(n33887), .Z(n33894) );
  XOR U46869 ( .A(n34832), .B(n34833), .Z(n34831) );
  IV U46870 ( .A(n33888), .Z(n33890) );
  NOR U46871 ( .A(n33890), .B(n33889), .Z(n34829) );
  NOR U46872 ( .A(n33891), .B(n34829), .Z(n33892) );
  XOR U46873 ( .A(n34831), .B(n33892), .Z(n33893) );
  NOR U46874 ( .A(n33894), .B(n33893), .Z(n33895) );
  NOR U46875 ( .A(n38389), .B(n33895), .Z(n33896) );
  IV U46876 ( .A(n33896), .Z(n34820) );
  NOR U46877 ( .A(n33898), .B(n33897), .Z(n33899) );
  NOR U46878 ( .A(n34821), .B(n33899), .Z(n33900) );
  XOR U46879 ( .A(n34820), .B(n33900), .Z(n34818) );
  IV U46880 ( .A(n33901), .Z(n33903) );
  NOR U46881 ( .A(n33903), .B(n33902), .Z(n34816) );
  XOR U46882 ( .A(n34818), .B(n34816), .Z(n37307) );
  XOR U46883 ( .A(n37305), .B(n37307), .Z(n37310) );
  XOR U46884 ( .A(n37308), .B(n37310), .Z(n37313) );
  XOR U46885 ( .A(n37312), .B(n37313), .Z(n37316) );
  XOR U46886 ( .A(n37315), .B(n37316), .Z(n37321) );
  XOR U46887 ( .A(n33904), .B(n37321), .Z(n33905) );
  IV U46888 ( .A(n33905), .Z(n37324) );
  XOR U46889 ( .A(n37323), .B(n37324), .Z(n34812) );
  IV U46890 ( .A(n33906), .Z(n33910) );
  NOR U46891 ( .A(n33908), .B(n33907), .Z(n33909) );
  IV U46892 ( .A(n33909), .Z(n33912) );
  NOR U46893 ( .A(n33910), .B(n33912), .Z(n34810) );
  XOR U46894 ( .A(n34812), .B(n34810), .Z(n37332) );
  IV U46895 ( .A(n33911), .Z(n33913) );
  NOR U46896 ( .A(n33913), .B(n33912), .Z(n37330) );
  XOR U46897 ( .A(n37332), .B(n37330), .Z(n34809) );
  IV U46898 ( .A(n33914), .Z(n33916) );
  NOR U46899 ( .A(n33916), .B(n33915), .Z(n34807) );
  XOR U46900 ( .A(n34809), .B(n34807), .Z(n38363) );
  IV U46901 ( .A(n33917), .Z(n33918) );
  NOR U46902 ( .A(n33923), .B(n33918), .Z(n34803) );
  IV U46903 ( .A(n33919), .Z(n33920) );
  NOR U46904 ( .A(n33921), .B(n33920), .Z(n38361) );
  IV U46905 ( .A(n33922), .Z(n33924) );
  NOR U46906 ( .A(n33924), .B(n33923), .Z(n40624) );
  NOR U46907 ( .A(n38361), .B(n40624), .Z(n34805) );
  IV U46908 ( .A(n34805), .Z(n33925) );
  NOR U46909 ( .A(n34803), .B(n33925), .Z(n33926) );
  XOR U46910 ( .A(n38363), .B(n33926), .Z(n34797) );
  IV U46911 ( .A(n33927), .Z(n33928) );
  NOR U46912 ( .A(n33930), .B(n33928), .Z(n34800) );
  IV U46913 ( .A(n33929), .Z(n33933) );
  NOR U46914 ( .A(n33931), .B(n33930), .Z(n33932) );
  IV U46915 ( .A(n33932), .Z(n33936) );
  NOR U46916 ( .A(n33933), .B(n33936), .Z(n34798) );
  NOR U46917 ( .A(n34800), .B(n34798), .Z(n33934) );
  XOR U46918 ( .A(n34797), .B(n33934), .Z(n37347) );
  IV U46919 ( .A(n33935), .Z(n33937) );
  NOR U46920 ( .A(n33937), .B(n33936), .Z(n37344) );
  IV U46921 ( .A(n33938), .Z(n33939) );
  NOR U46922 ( .A(n33939), .B(n33943), .Z(n37346) );
  NOR U46923 ( .A(n37344), .B(n37346), .Z(n33940) );
  XOR U46924 ( .A(n37347), .B(n33940), .Z(n34789) );
  IV U46925 ( .A(n33941), .Z(n34790) );
  NOR U46926 ( .A(n34792), .B(n34790), .Z(n33945) );
  IV U46927 ( .A(n33942), .Z(n33944) );
  NOR U46928 ( .A(n33944), .B(n33943), .Z(n37340) );
  NOR U46929 ( .A(n33945), .B(n37340), .Z(n33946) );
  XOR U46930 ( .A(n34789), .B(n33946), .Z(n34794) );
  IV U46931 ( .A(n33947), .Z(n33949) );
  NOR U46932 ( .A(n33949), .B(n33948), .Z(n34793) );
  IV U46933 ( .A(n33950), .Z(n33951) );
  NOR U46934 ( .A(n33954), .B(n33951), .Z(n34787) );
  NOR U46935 ( .A(n34793), .B(n34787), .Z(n33952) );
  XOR U46936 ( .A(n34794), .B(n33952), .Z(n34784) );
  IV U46937 ( .A(n33953), .Z(n33955) );
  NOR U46938 ( .A(n33955), .B(n33954), .Z(n34785) );
  NOR U46939 ( .A(n34785), .B(n37355), .Z(n33956) );
  XOR U46940 ( .A(n34784), .B(n33956), .Z(n34782) );
  XOR U46941 ( .A(n33957), .B(n34782), .Z(n33958) );
  IV U46942 ( .A(n33958), .Z(n37360) );
  IV U46943 ( .A(n33959), .Z(n33962) );
  IV U46944 ( .A(n33960), .Z(n33961) );
  NOR U46945 ( .A(n33962), .B(n33961), .Z(n33964) );
  IV U46946 ( .A(n33964), .Z(n44040) );
  NOR U46947 ( .A(n37360), .B(n44040), .Z(n40658) );
  XOR U46948 ( .A(n37358), .B(n37360), .Z(n44043) );
  IV U46949 ( .A(n44043), .Z(n33963) );
  NOR U46950 ( .A(n33964), .B(n33963), .Z(n33965) );
  NOR U46951 ( .A(n40658), .B(n33965), .Z(n34773) );
  IV U46952 ( .A(n33966), .Z(n33969) );
  IV U46953 ( .A(n33967), .Z(n33968) );
  NOR U46954 ( .A(n33969), .B(n33968), .Z(n33970) );
  IV U46955 ( .A(n33970), .Z(n34774) );
  XOR U46956 ( .A(n34773), .B(n34774), .Z(n34777) );
  XOR U46957 ( .A(n34776), .B(n34777), .Z(n37365) );
  IV U46958 ( .A(n33971), .Z(n33973) );
  NOR U46959 ( .A(n33973), .B(n33972), .Z(n37363) );
  XOR U46960 ( .A(n37365), .B(n37363), .Z(n37367) );
  XOR U46961 ( .A(n37366), .B(n37367), .Z(n38320) );
  XOR U46962 ( .A(n33974), .B(n38320), .Z(n34764) );
  NOR U46963 ( .A(n34763), .B(n34769), .Z(n33975) );
  NOR U46964 ( .A(n33975), .B(n34765), .Z(n33976) );
  XOR U46965 ( .A(n34764), .B(n33976), .Z(n34756) );
  NOR U46966 ( .A(n33977), .B(n34756), .Z(n38302) );
  IV U46967 ( .A(n33978), .Z(n41570) );
  NOR U46968 ( .A(n41570), .B(n33979), .Z(n33980) );
  IV U46969 ( .A(n33980), .Z(n34753) );
  IV U46970 ( .A(n33981), .Z(n33982) );
  NOR U46971 ( .A(n34757), .B(n33982), .Z(n33983) );
  XOR U46972 ( .A(n34756), .B(n33983), .Z(n34752) );
  XOR U46973 ( .A(n34753), .B(n34752), .Z(n33984) );
  NOR U46974 ( .A(n33985), .B(n33984), .Z(n33986) );
  NOR U46975 ( .A(n38302), .B(n33986), .Z(n37375) );
  IV U46976 ( .A(n33987), .Z(n33988) );
  NOR U46977 ( .A(n41570), .B(n33988), .Z(n37374) );
  IV U46978 ( .A(n33989), .Z(n37383) );
  NOR U46979 ( .A(n37385), .B(n37383), .Z(n33990) );
  NOR U46980 ( .A(n37374), .B(n33990), .Z(n33991) );
  XOR U46981 ( .A(n37375), .B(n33991), .Z(n37380) );
  IV U46982 ( .A(n33992), .Z(n33994) );
  NOR U46983 ( .A(n33994), .B(n33993), .Z(n33995) );
  IV U46984 ( .A(n33995), .Z(n33997) );
  NOR U46985 ( .A(n33997), .B(n33996), .Z(n37378) );
  XOR U46986 ( .A(n37380), .B(n37378), .Z(n37391) );
  XOR U46987 ( .A(n37389), .B(n37391), .Z(n37396) );
  XOR U46988 ( .A(n33998), .B(n37396), .Z(n34748) );
  XOR U46989 ( .A(n34749), .B(n34748), .Z(n37401) );
  XOR U46990 ( .A(n37400), .B(n37401), .Z(n34746) );
  XOR U46991 ( .A(n34745), .B(n34746), .Z(n34743) );
  XOR U46992 ( .A(n34742), .B(n34743), .Z(n34738) );
  XOR U46993 ( .A(n33999), .B(n34738), .Z(n34732) );
  IV U46994 ( .A(n34000), .Z(n34002) );
  NOR U46995 ( .A(n34002), .B(n34001), .Z(n34728) );
  NOR U46996 ( .A(n34731), .B(n34728), .Z(n34003) );
  XOR U46997 ( .A(n34732), .B(n34003), .Z(n37420) );
  IV U46998 ( .A(n34004), .Z(n34006) );
  NOR U46999 ( .A(n34006), .B(n34005), .Z(n37418) );
  XOR U47000 ( .A(n37420), .B(n37418), .Z(n37422) );
  XOR U47001 ( .A(n37421), .B(n37422), .Z(n34725) );
  XOR U47002 ( .A(n34723), .B(n34725), .Z(n37426) );
  XOR U47003 ( .A(n34007), .B(n37426), .Z(n34720) );
  XOR U47004 ( .A(n34721), .B(n34720), .Z(n37430) );
  XOR U47005 ( .A(n37428), .B(n37430), .Z(n37433) );
  IV U47006 ( .A(n37433), .Z(n34018) );
  IV U47007 ( .A(n34008), .Z(n34013) );
  NOR U47008 ( .A(n34010), .B(n34009), .Z(n34011) );
  IV U47009 ( .A(n34011), .Z(n34012) );
  NOR U47010 ( .A(n34013), .B(n34012), .Z(n34718) );
  IV U47011 ( .A(n34014), .Z(n34016) );
  NOR U47012 ( .A(n34016), .B(n34015), .Z(n37431) );
  NOR U47013 ( .A(n34718), .B(n37431), .Z(n34017) );
  XOR U47014 ( .A(n34018), .B(n34017), .Z(n37440) );
  XOR U47015 ( .A(n37438), .B(n37440), .Z(n37443) );
  XOR U47016 ( .A(n37441), .B(n37443), .Z(n37447) );
  XOR U47017 ( .A(n37445), .B(n37447), .Z(n37449) );
  XOR U47018 ( .A(n37448), .B(n37449), .Z(n37457) );
  XOR U47019 ( .A(n34019), .B(n37457), .Z(n37459) );
  NOR U47020 ( .A(n34020), .B(n37459), .Z(n34022) );
  IV U47021 ( .A(n34020), .Z(n34021) );
  NOR U47022 ( .A(n37457), .B(n34021), .Z(n40749) );
  NOR U47023 ( .A(n34022), .B(n40749), .Z(n34716) );
  XOR U47024 ( .A(n34023), .B(n34716), .Z(n34714) );
  XOR U47025 ( .A(n34024), .B(n34714), .Z(n37474) );
  XOR U47026 ( .A(n34025), .B(n37474), .Z(n37485) );
  NOR U47027 ( .A(n34027), .B(n34026), .Z(n37483) );
  NOR U47028 ( .A(n37480), .B(n37483), .Z(n34028) );
  XOR U47029 ( .A(n37485), .B(n34028), .Z(n34029) );
  IV U47030 ( .A(n34029), .Z(n37487) );
  XOR U47031 ( .A(n37486), .B(n37487), .Z(n34707) );
  XOR U47032 ( .A(n34706), .B(n34707), .Z(n37496) );
  XOR U47033 ( .A(n34030), .B(n37496), .Z(n37503) );
  XOR U47034 ( .A(n34031), .B(n37503), .Z(n34032) );
  IV U47035 ( .A(n34032), .Z(n37507) );
  XOR U47036 ( .A(n37505), .B(n37507), .Z(n37508) );
  XOR U47037 ( .A(n37509), .B(n37508), .Z(n34695) );
  IV U47038 ( .A(n34687), .Z(n34041) );
  IV U47039 ( .A(n34033), .Z(n34686) );
  NOR U47040 ( .A(n34041), .B(n34686), .Z(n34694) );
  IV U47041 ( .A(n34034), .Z(n34036) );
  NOR U47042 ( .A(n34036), .B(n34035), .Z(n34701) );
  NOR U47043 ( .A(n34694), .B(n34701), .Z(n34037) );
  XOR U47044 ( .A(n34695), .B(n34037), .Z(n44182) );
  NOR U47045 ( .A(n34038), .B(n44182), .Z(n40802) );
  IV U47046 ( .A(n34039), .Z(n34040) );
  NOR U47047 ( .A(n34041), .B(n34040), .Z(n34697) );
  XOR U47048 ( .A(n34697), .B(n44182), .Z(n34047) );
  IV U47049 ( .A(n34047), .Z(n34042) );
  NOR U47050 ( .A(n34043), .B(n34042), .Z(n34044) );
  NOR U47051 ( .A(n40802), .B(n34044), .Z(n34688) );
  NOR U47052 ( .A(n34045), .B(n34690), .Z(n34046) );
  NOR U47053 ( .A(n34688), .B(n34046), .Z(n34050) );
  IV U47054 ( .A(n34046), .Z(n34048) );
  NOR U47055 ( .A(n34048), .B(n34047), .Z(n34049) );
  NOR U47056 ( .A(n34050), .B(n34049), .Z(n37514) );
  XOR U47057 ( .A(n34051), .B(n37514), .Z(n34679) );
  XOR U47058 ( .A(n34678), .B(n34679), .Z(n34681) );
  XOR U47059 ( .A(n34052), .B(n34681), .Z(n34053) );
  IV U47060 ( .A(n34053), .Z(n34675) );
  XOR U47061 ( .A(n34673), .B(n34675), .Z(n37522) );
  XOR U47062 ( .A(n37521), .B(n37522), .Z(n37541) );
  IV U47063 ( .A(n37541), .Z(n34058) );
  IV U47064 ( .A(n34054), .Z(n34056) );
  NOR U47065 ( .A(n34056), .B(n34055), .Z(n37532) );
  NOR U47066 ( .A(n37534), .B(n37532), .Z(n34057) );
  XOR U47067 ( .A(n34058), .B(n34057), .Z(n37553) );
  NOR U47068 ( .A(n34059), .B(n37542), .Z(n34063) );
  IV U47069 ( .A(n34060), .Z(n34062) );
  IV U47070 ( .A(n34061), .Z(n34069) );
  NOR U47071 ( .A(n34062), .B(n34069), .Z(n37551) );
  NOR U47072 ( .A(n34063), .B(n37551), .Z(n34064) );
  XOR U47073 ( .A(n37553), .B(n34064), .Z(n34671) );
  IV U47074 ( .A(n34065), .Z(n34066) );
  NOR U47075 ( .A(n34066), .B(n34069), .Z(n37548) );
  IV U47076 ( .A(n34067), .Z(n34068) );
  NOR U47077 ( .A(n34069), .B(n34068), .Z(n34670) );
  NOR U47078 ( .A(n37548), .B(n34670), .Z(n34070) );
  XOR U47079 ( .A(n34671), .B(n34070), .Z(n34664) );
  IV U47080 ( .A(n34071), .Z(n34072) );
  NOR U47081 ( .A(n34073), .B(n34072), .Z(n34662) );
  IV U47082 ( .A(n34074), .Z(n34076) );
  NOR U47083 ( .A(n34076), .B(n34075), .Z(n34660) );
  NOR U47084 ( .A(n34662), .B(n34660), .Z(n34077) );
  XOR U47085 ( .A(n34664), .B(n34077), .Z(n34654) );
  IV U47086 ( .A(n34078), .Z(n34079) );
  NOR U47087 ( .A(n34080), .B(n34079), .Z(n34666) );
  IV U47088 ( .A(n34081), .Z(n34082) );
  NOR U47089 ( .A(n34083), .B(n34082), .Z(n34655) );
  NOR U47090 ( .A(n34666), .B(n34655), .Z(n34084) );
  XOR U47091 ( .A(n34654), .B(n34084), .Z(n34658) );
  XOR U47092 ( .A(n34657), .B(n34658), .Z(n34652) );
  XOR U47093 ( .A(n34085), .B(n34652), .Z(n34086) );
  IV U47094 ( .A(n34086), .Z(n34648) );
  XOR U47095 ( .A(n34646), .B(n34648), .Z(n41476) );
  IV U47096 ( .A(n41476), .Z(n34089) );
  NOR U47097 ( .A(n34087), .B(n41483), .Z(n34638) );
  NOR U47098 ( .A(n34643), .B(n34638), .Z(n34088) );
  XOR U47099 ( .A(n34089), .B(n34088), .Z(n38192) );
  XOR U47100 ( .A(n34090), .B(n38192), .Z(n34633) );
  XOR U47101 ( .A(n34632), .B(n34633), .Z(n34636) );
  XOR U47102 ( .A(n34635), .B(n34636), .Z(n38182) );
  XOR U47103 ( .A(n34627), .B(n38182), .Z(n34628) );
  XOR U47104 ( .A(n34630), .B(n34628), .Z(n34625) );
  XOR U47105 ( .A(n34624), .B(n34625), .Z(n34091) );
  XOR U47106 ( .A(n34092), .B(n34091), .Z(n34614) );
  XOR U47107 ( .A(n34093), .B(n34614), .Z(n34610) );
  XOR U47108 ( .A(n34609), .B(n34610), .Z(n34099) );
  NOR U47109 ( .A(n34094), .B(n34099), .Z(n40856) );
  NOR U47110 ( .A(n34096), .B(n34095), .Z(n34101) );
  IV U47111 ( .A(n34101), .Z(n34097) );
  NOR U47112 ( .A(n34097), .B(n34610), .Z(n38162) );
  NOR U47113 ( .A(n40856), .B(n38162), .Z(n34098) );
  IV U47114 ( .A(n34098), .Z(n34102) );
  NOR U47115 ( .A(n34102), .B(n34099), .Z(n34105) );
  NOR U47116 ( .A(n34101), .B(n34100), .Z(n34103) );
  NOR U47117 ( .A(n34103), .B(n34102), .Z(n34104) );
  NOR U47118 ( .A(n34105), .B(n34104), .Z(n37564) );
  XOR U47119 ( .A(n37562), .B(n37564), .Z(n37566) );
  XOR U47120 ( .A(n37565), .B(n37566), .Z(n34605) );
  XOR U47121 ( .A(n34106), .B(n34605), .Z(n34107) );
  IV U47122 ( .A(n34107), .Z(n34600) );
  XOR U47123 ( .A(n34108), .B(n34600), .Z(n37574) );
  XOR U47124 ( .A(n37572), .B(n37574), .Z(n37577) );
  IV U47125 ( .A(n34109), .Z(n34592) );
  NOR U47126 ( .A(n34110), .B(n34592), .Z(n34114) );
  IV U47127 ( .A(n34111), .Z(n34112) );
  NOR U47128 ( .A(n34113), .B(n34112), .Z(n37575) );
  NOR U47129 ( .A(n34114), .B(n37575), .Z(n34115) );
  XOR U47130 ( .A(n37577), .B(n34115), .Z(n34575) );
  NOR U47131 ( .A(n34116), .B(n34584), .Z(n34576) );
  IV U47132 ( .A(n34117), .Z(n34118) );
  NOR U47133 ( .A(n34118), .B(n34579), .Z(n34119) );
  NOR U47134 ( .A(n34576), .B(n34119), .Z(n34120) );
  XOR U47135 ( .A(n34575), .B(n34120), .Z(n34573) );
  XOR U47136 ( .A(n34571), .B(n34573), .Z(n34128) );
  IV U47137 ( .A(n34121), .Z(n34123) );
  NOR U47138 ( .A(n34123), .B(n34122), .Z(n34577) );
  IV U47139 ( .A(n34124), .Z(n34126) );
  NOR U47140 ( .A(n34126), .B(n34125), .Z(n34572) );
  NOR U47141 ( .A(n34577), .B(n34572), .Z(n34127) );
  XOR U47142 ( .A(n34128), .B(n34127), .Z(n34567) );
  IV U47143 ( .A(n34129), .Z(n34131) );
  NOR U47144 ( .A(n34131), .B(n34130), .Z(n34565) );
  XOR U47145 ( .A(n34567), .B(n34565), .Z(n34569) );
  XOR U47146 ( .A(n34568), .B(n34569), .Z(n37581) );
  XOR U47147 ( .A(n37580), .B(n37581), .Z(n37584) );
  XOR U47148 ( .A(n37583), .B(n37584), .Z(n37588) );
  XOR U47149 ( .A(n34132), .B(n37588), .Z(n34133) );
  IV U47150 ( .A(n34133), .Z(n34559) );
  XOR U47151 ( .A(n34557), .B(n34559), .Z(n34562) );
  IV U47152 ( .A(n34562), .Z(n34138) );
  IV U47153 ( .A(n34134), .Z(n34135) );
  NOR U47154 ( .A(n34136), .B(n34135), .Z(n34560) );
  NOR U47155 ( .A(n34555), .B(n34560), .Z(n34137) );
  XOR U47156 ( .A(n34138), .B(n34137), .Z(n34554) );
  XOR U47157 ( .A(n34552), .B(n34554), .Z(n34548) );
  XOR U47158 ( .A(n34547), .B(n34548), .Z(n34545) );
  XOR U47159 ( .A(n34546), .B(n34545), .Z(n34146) );
  IV U47160 ( .A(n34146), .Z(n34139) );
  NOR U47161 ( .A(n34140), .B(n34139), .Z(n40910) );
  IV U47162 ( .A(n34141), .Z(n34143) );
  NOR U47163 ( .A(n34143), .B(n34142), .Z(n34145) );
  IV U47164 ( .A(n34145), .Z(n34144) );
  NOR U47165 ( .A(n34545), .B(n34144), .Z(n40913) );
  NOR U47166 ( .A(n34146), .B(n34145), .Z(n34147) );
  NOR U47167 ( .A(n40913), .B(n34147), .Z(n34148) );
  NOR U47168 ( .A(n34149), .B(n34148), .Z(n34150) );
  NOR U47169 ( .A(n40910), .B(n34150), .Z(n34151) );
  IV U47170 ( .A(n34151), .Z(n37594) );
  XOR U47171 ( .A(n37594), .B(n37593), .Z(n37601) );
  NOR U47172 ( .A(n34152), .B(n37601), .Z(n38101) );
  IV U47173 ( .A(n34153), .Z(n34157) );
  NOR U47174 ( .A(n34155), .B(n34154), .Z(n34156) );
  IV U47175 ( .A(n34156), .Z(n34159) );
  NOR U47176 ( .A(n34157), .B(n34159), .Z(n37600) );
  IV U47177 ( .A(n34158), .Z(n34160) );
  NOR U47178 ( .A(n34160), .B(n34159), .Z(n37596) );
  NOR U47179 ( .A(n37600), .B(n37596), .Z(n34161) );
  XOR U47180 ( .A(n34161), .B(n37601), .Z(n34541) );
  NOR U47181 ( .A(n34162), .B(n34541), .Z(n34163) );
  NOR U47182 ( .A(n38101), .B(n34163), .Z(n34538) );
  IV U47183 ( .A(n34164), .Z(n34165) );
  NOR U47184 ( .A(n34166), .B(n34165), .Z(n34542) );
  IV U47185 ( .A(n34167), .Z(n34169) );
  NOR U47186 ( .A(n34169), .B(n34168), .Z(n34537) );
  NOR U47187 ( .A(n34542), .B(n34537), .Z(n34170) );
  XOR U47188 ( .A(n34538), .B(n34170), .Z(n34533) );
  IV U47189 ( .A(n34171), .Z(n34173) );
  NOR U47190 ( .A(n34173), .B(n34172), .Z(n34531) );
  XOR U47191 ( .A(n34533), .B(n34531), .Z(n34535) );
  XOR U47192 ( .A(n34534), .B(n34535), .Z(n40938) );
  XOR U47193 ( .A(n34526), .B(n40938), .Z(n34524) );
  IV U47194 ( .A(n34174), .Z(n34176) );
  NOR U47195 ( .A(n34176), .B(n34175), .Z(n34527) );
  NOR U47196 ( .A(n34178), .B(n34177), .Z(n34523) );
  NOR U47197 ( .A(n34527), .B(n34523), .Z(n34179) );
  XOR U47198 ( .A(n34524), .B(n34179), .Z(n34519) );
  XOR U47199 ( .A(n34518), .B(n34519), .Z(n37607) );
  XOR U47200 ( .A(n34521), .B(n37607), .Z(n34184) );
  IV U47201 ( .A(n34180), .Z(n34182) );
  NOR U47202 ( .A(n34182), .B(n34181), .Z(n34190) );
  IV U47203 ( .A(n34190), .Z(n34183) );
  NOR U47204 ( .A(n34184), .B(n34183), .Z(n38088) );
  IV U47205 ( .A(n34185), .Z(n34187) );
  NOR U47206 ( .A(n34187), .B(n34186), .Z(n37606) );
  NOR U47207 ( .A(n34521), .B(n37606), .Z(n34188) );
  XOR U47208 ( .A(n37607), .B(n34188), .Z(n34189) );
  NOR U47209 ( .A(n34190), .B(n34189), .Z(n34191) );
  NOR U47210 ( .A(n38088), .B(n34191), .Z(n37610) );
  XOR U47211 ( .A(n37612), .B(n37610), .Z(n37614) );
  XOR U47212 ( .A(n37613), .B(n37614), .Z(n37618) );
  XOR U47213 ( .A(n37617), .B(n37618), .Z(n37622) );
  XOR U47214 ( .A(n37620), .B(n37622), .Z(n34517) );
  XOR U47215 ( .A(n34192), .B(n34517), .Z(n34193) );
  IV U47216 ( .A(n34193), .Z(n34508) );
  XOR U47217 ( .A(n34500), .B(n34508), .Z(n34498) );
  XOR U47218 ( .A(n34497), .B(n34498), .Z(n37626) );
  XOR U47219 ( .A(n37625), .B(n37626), .Z(n37634) );
  IV U47220 ( .A(n37634), .Z(n34200) );
  IV U47221 ( .A(n34194), .Z(n34198) );
  NOR U47222 ( .A(n34196), .B(n34195), .Z(n34197) );
  IV U47223 ( .A(n34197), .Z(n34202) );
  NOR U47224 ( .A(n34198), .B(n34202), .Z(n37632) );
  NOR U47225 ( .A(n37628), .B(n37632), .Z(n34199) );
  XOR U47226 ( .A(n34200), .B(n34199), .Z(n34495) );
  IV U47227 ( .A(n34201), .Z(n34203) );
  NOR U47228 ( .A(n34203), .B(n34202), .Z(n34493) );
  XOR U47229 ( .A(n34495), .B(n34493), .Z(n37636) );
  XOR U47230 ( .A(n37635), .B(n37636), .Z(n37640) );
  XOR U47231 ( .A(n37638), .B(n37640), .Z(n34492) );
  XOR U47232 ( .A(n34490), .B(n34492), .Z(n37643) );
  XOR U47233 ( .A(n37642), .B(n37643), .Z(n37647) );
  IV U47234 ( .A(n34204), .Z(n34208) );
  NOR U47235 ( .A(n34206), .B(n34205), .Z(n34207) );
  IV U47236 ( .A(n34207), .Z(n34210) );
  NOR U47237 ( .A(n34208), .B(n34210), .Z(n34213) );
  IV U47238 ( .A(n34213), .Z(n41348) );
  NOR U47239 ( .A(n37647), .B(n41348), .Z(n40983) );
  IV U47240 ( .A(n34209), .Z(n34211) );
  NOR U47241 ( .A(n34211), .B(n34210), .Z(n37645) );
  XOR U47242 ( .A(n37647), .B(n37645), .Z(n41345) );
  IV U47243 ( .A(n41345), .Z(n34212) );
  NOR U47244 ( .A(n34213), .B(n34212), .Z(n34214) );
  NOR U47245 ( .A(n40983), .B(n34214), .Z(n37649) );
  IV U47246 ( .A(n34215), .Z(n34217) );
  NOR U47247 ( .A(n34217), .B(n34216), .Z(n34218) );
  IV U47248 ( .A(n34218), .Z(n37650) );
  XOR U47249 ( .A(n37649), .B(n37650), .Z(n37654) );
  XOR U47250 ( .A(n37653), .B(n37654), .Z(n37657) );
  NOR U47251 ( .A(n34219), .B(n34221), .Z(n37656) );
  IV U47252 ( .A(n34220), .Z(n34222) );
  NOR U47253 ( .A(n34222), .B(n34221), .Z(n34487) );
  NOR U47254 ( .A(n37656), .B(n34487), .Z(n34223) );
  XOR U47255 ( .A(n37657), .B(n34223), .Z(n34482) );
  XOR U47256 ( .A(n34224), .B(n34482), .Z(n37663) );
  XOR U47257 ( .A(n37661), .B(n37663), .Z(n37670) );
  IV U47258 ( .A(n34225), .Z(n34227) );
  NOR U47259 ( .A(n34227), .B(n34226), .Z(n37669) );
  NOR U47260 ( .A(n37664), .B(n37669), .Z(n34228) );
  XOR U47261 ( .A(n37670), .B(n34228), .Z(n37667) );
  IV U47262 ( .A(n34229), .Z(n34230) );
  NOR U47263 ( .A(n34230), .B(n34238), .Z(n38059) );
  NOR U47264 ( .A(n34232), .B(n34231), .Z(n41024) );
  NOR U47265 ( .A(n38059), .B(n41024), .Z(n37668) );
  XOR U47266 ( .A(n37667), .B(n37668), .Z(n37675) );
  XOR U47267 ( .A(n37674), .B(n37675), .Z(n37679) );
  IV U47268 ( .A(n37679), .Z(n34240) );
  IV U47269 ( .A(n34233), .Z(n34234) );
  NOR U47270 ( .A(n34235), .B(n34234), .Z(n34479) );
  IV U47271 ( .A(n34236), .Z(n34237) );
  NOR U47272 ( .A(n34238), .B(n34237), .Z(n37677) );
  NOR U47273 ( .A(n34479), .B(n37677), .Z(n34239) );
  XOR U47274 ( .A(n34240), .B(n34239), .Z(n44416) );
  XOR U47275 ( .A(n44415), .B(n44416), .Z(n34478) );
  XOR U47276 ( .A(n34241), .B(n34478), .Z(n34470) );
  XOR U47277 ( .A(n34242), .B(n34470), .Z(n34468) );
  XOR U47278 ( .A(n34243), .B(n34468), .Z(n34244) );
  IV U47279 ( .A(n34244), .Z(n34456) );
  XOR U47280 ( .A(n34454), .B(n34456), .Z(n37685) );
  IV U47281 ( .A(n37685), .Z(n34252) );
  IV U47282 ( .A(n34245), .Z(n34246) );
  NOR U47283 ( .A(n34247), .B(n34246), .Z(n37684) );
  IV U47284 ( .A(n34248), .Z(n34250) );
  NOR U47285 ( .A(n34250), .B(n34249), .Z(n34452) );
  NOR U47286 ( .A(n37684), .B(n34452), .Z(n34251) );
  XOR U47287 ( .A(n34252), .B(n34251), .Z(n34451) );
  IV U47288 ( .A(n34253), .Z(n34254) );
  NOR U47289 ( .A(n34255), .B(n34254), .Z(n34449) );
  XOR U47290 ( .A(n34451), .B(n34449), .Z(n37689) );
  XOR U47291 ( .A(n37687), .B(n37689), .Z(n37693) );
  IV U47292 ( .A(n34256), .Z(n34258) );
  NOR U47293 ( .A(n34258), .B(n34257), .Z(n37692) );
  IV U47294 ( .A(n34259), .Z(n34261) );
  NOR U47295 ( .A(n34261), .B(n34260), .Z(n37690) );
  NOR U47296 ( .A(n37692), .B(n37690), .Z(n34262) );
  XOR U47297 ( .A(n37693), .B(n34262), .Z(n34263) );
  NOR U47298 ( .A(n34264), .B(n34263), .Z(n34267) );
  IV U47299 ( .A(n34264), .Z(n34266) );
  XOR U47300 ( .A(n37692), .B(n37693), .Z(n34265) );
  NOR U47301 ( .A(n34266), .B(n34265), .Z(n44452) );
  NOR U47302 ( .A(n34267), .B(n44452), .Z(n34276) );
  IV U47303 ( .A(n34276), .Z(n37699) );
  IV U47304 ( .A(n34268), .Z(n34271) );
  NOR U47305 ( .A(n34269), .B(n34285), .Z(n34270) );
  IV U47306 ( .A(n34270), .Z(n34273) );
  NOR U47307 ( .A(n34271), .B(n34273), .Z(n34278) );
  IV U47308 ( .A(n34278), .Z(n44460) );
  NOR U47309 ( .A(n37699), .B(n44460), .Z(n38025) );
  IV U47310 ( .A(n34272), .Z(n34274) );
  NOR U47311 ( .A(n34274), .B(n34273), .Z(n34275) );
  IV U47312 ( .A(n34275), .Z(n37698) );
  XOR U47313 ( .A(n34276), .B(n37698), .Z(n44463) );
  IV U47314 ( .A(n44463), .Z(n34277) );
  NOR U47315 ( .A(n34278), .B(n34277), .Z(n34279) );
  NOR U47316 ( .A(n38025), .B(n34279), .Z(n37700) );
  IV U47317 ( .A(n34280), .Z(n34289) );
  IV U47318 ( .A(n34281), .Z(n34282) );
  NOR U47319 ( .A(n34289), .B(n34282), .Z(n37704) );
  IV U47320 ( .A(n34283), .Z(n34284) );
  NOR U47321 ( .A(n34285), .B(n34284), .Z(n37701) );
  NOR U47322 ( .A(n37704), .B(n37701), .Z(n34286) );
  XOR U47323 ( .A(n37700), .B(n34286), .Z(n34448) );
  IV U47324 ( .A(n34287), .Z(n34288) );
  NOR U47325 ( .A(n34289), .B(n34288), .Z(n34290) );
  IV U47326 ( .A(n34290), .Z(n34447) );
  XOR U47327 ( .A(n34448), .B(n34447), .Z(n34295) );
  IV U47328 ( .A(n34295), .Z(n34293) );
  IV U47329 ( .A(n34291), .Z(n34292) );
  NOR U47330 ( .A(n34292), .B(n34304), .Z(n34299) );
  IV U47331 ( .A(n34299), .Z(n41282) );
  NOR U47332 ( .A(n34293), .B(n41282), .Z(n34446) );
  NOR U47333 ( .A(n34304), .B(n34294), .Z(n34296) );
  NOR U47334 ( .A(n34296), .B(n34295), .Z(n34298) );
  IV U47335 ( .A(n34296), .Z(n34297) );
  NOR U47336 ( .A(n34448), .B(n34297), .Z(n41062) );
  NOR U47337 ( .A(n34298), .B(n41062), .Z(n41277) );
  NOR U47338 ( .A(n34299), .B(n41277), .Z(n34300) );
  NOR U47339 ( .A(n34446), .B(n34300), .Z(n34301) );
  IV U47340 ( .A(n34301), .Z(n34445) );
  IV U47341 ( .A(n34302), .Z(n34303) );
  NOR U47342 ( .A(n34304), .B(n34303), .Z(n34443) );
  XOR U47343 ( .A(n34445), .B(n34443), .Z(n38017) );
  XOR U47344 ( .A(n34442), .B(n38017), .Z(n34305) );
  IV U47345 ( .A(n34305), .Z(n34437) );
  XOR U47346 ( .A(n34436), .B(n34437), .Z(n34440) );
  IV U47347 ( .A(n34440), .Z(n34313) );
  IV U47348 ( .A(n34306), .Z(n34308) );
  NOR U47349 ( .A(n34308), .B(n34307), .Z(n34439) );
  IV U47350 ( .A(n34309), .Z(n34310) );
  NOR U47351 ( .A(n34311), .B(n34310), .Z(n34434) );
  NOR U47352 ( .A(n34439), .B(n34434), .Z(n34312) );
  XOR U47353 ( .A(n34313), .B(n34312), .Z(n37712) );
  XOR U47354 ( .A(n37711), .B(n37712), .Z(n37715) );
  XOR U47355 ( .A(n37714), .B(n37715), .Z(n37720) );
  XOR U47356 ( .A(n37718), .B(n37720), .Z(n37722) );
  XOR U47357 ( .A(n34314), .B(n37722), .Z(n37735) );
  NOR U47358 ( .A(n34322), .B(n37735), .Z(n41246) );
  IV U47359 ( .A(n34315), .Z(n34316) );
  NOR U47360 ( .A(n37723), .B(n34316), .Z(n37733) );
  XOR U47361 ( .A(n37735), .B(n37733), .Z(n34430) );
  IV U47362 ( .A(n34317), .Z(n34321) );
  NOR U47363 ( .A(n34319), .B(n34318), .Z(n34320) );
  IV U47364 ( .A(n34320), .Z(n34328) );
  NOR U47365 ( .A(n34321), .B(n34328), .Z(n34323) );
  IV U47366 ( .A(n34323), .Z(n34429) );
  XOR U47367 ( .A(n34430), .B(n34429), .Z(n34325) );
  NOR U47368 ( .A(n34323), .B(n34322), .Z(n34324) );
  NOR U47369 ( .A(n34325), .B(n34324), .Z(n34326) );
  NOR U47370 ( .A(n41246), .B(n34326), .Z(n34431) );
  IV U47371 ( .A(n34327), .Z(n34329) );
  NOR U47372 ( .A(n34329), .B(n34328), .Z(n34330) );
  IV U47373 ( .A(n34330), .Z(n34432) );
  XOR U47374 ( .A(n34431), .B(n34432), .Z(n37739) );
  XOR U47375 ( .A(n34427), .B(n37739), .Z(n37742) );
  IV U47376 ( .A(n37742), .Z(n34339) );
  IV U47377 ( .A(n34331), .Z(n34334) );
  IV U47378 ( .A(n34332), .Z(n34333) );
  NOR U47379 ( .A(n34334), .B(n34333), .Z(n37740) );
  IV U47380 ( .A(n34335), .Z(n34337) );
  NOR U47381 ( .A(n34337), .B(n34336), .Z(n37737) );
  NOR U47382 ( .A(n37740), .B(n37737), .Z(n34338) );
  XOR U47383 ( .A(n34339), .B(n34338), .Z(n34426) );
  IV U47384 ( .A(n34340), .Z(n34341) );
  NOR U47385 ( .A(n34341), .B(n34343), .Z(n34424) );
  IV U47386 ( .A(n34342), .Z(n34346) );
  NOR U47387 ( .A(n34344), .B(n34343), .Z(n34345) );
  IV U47388 ( .A(n34345), .Z(n34349) );
  NOR U47389 ( .A(n34346), .B(n34349), .Z(n34422) );
  NOR U47390 ( .A(n34424), .B(n34422), .Z(n34347) );
  XOR U47391 ( .A(n34426), .B(n34347), .Z(n34351) );
  IV U47392 ( .A(n34348), .Z(n34350) );
  NOR U47393 ( .A(n34350), .B(n34349), .Z(n34352) );
  NOR U47394 ( .A(n34351), .B(n34352), .Z(n34355) );
  XOR U47395 ( .A(n34424), .B(n34426), .Z(n34354) );
  IV U47396 ( .A(n34352), .Z(n34353) );
  NOR U47397 ( .A(n34354), .B(n34353), .Z(n37991) );
  NOR U47398 ( .A(n34355), .B(n37991), .Z(n34418) );
  XOR U47399 ( .A(n34356), .B(n34418), .Z(n34414) );
  XOR U47400 ( .A(n34412), .B(n34414), .Z(n37760) );
  IV U47401 ( .A(n37760), .Z(n34364) );
  IV U47402 ( .A(n34357), .Z(n34358) );
  NOR U47403 ( .A(n34359), .B(n34358), .Z(n34415) );
  IV U47404 ( .A(n34360), .Z(n34362) );
  NOR U47405 ( .A(n34362), .B(n34361), .Z(n37759) );
  NOR U47406 ( .A(n34415), .B(n37759), .Z(n34363) );
  XOR U47407 ( .A(n34364), .B(n34363), .Z(n37756) );
  XOR U47408 ( .A(n37755), .B(n37756), .Z(n34410) );
  XOR U47409 ( .A(n34365), .B(n34410), .Z(n34366) );
  IV U47410 ( .A(n34366), .Z(n37770) );
  IV U47411 ( .A(n34367), .Z(n37773) );
  NOR U47412 ( .A(n37771), .B(n37773), .Z(n34368) );
  XOR U47413 ( .A(n37770), .B(n34368), .Z(n37776) );
  IV U47414 ( .A(n34369), .Z(n34371) );
  NOR U47415 ( .A(n34371), .B(n34370), .Z(n37774) );
  XOR U47416 ( .A(n37776), .B(n37774), .Z(n34401) );
  XOR U47417 ( .A(n34400), .B(n34401), .Z(n34404) );
  XOR U47418 ( .A(n34403), .B(n34404), .Z(n34395) );
  IV U47419 ( .A(n34372), .Z(n34374) );
  NOR U47420 ( .A(n34374), .B(n34373), .Z(n34390) );
  NOR U47421 ( .A(n34375), .B(n34390), .Z(n34377) );
  NOR U47422 ( .A(n34377), .B(n34376), .Z(n34383) );
  XOR U47423 ( .A(n34378), .B(n34377), .Z(n37790) );
  IV U47424 ( .A(n34379), .Z(n34381) );
  NOR U47425 ( .A(n34381), .B(n34380), .Z(n37788) );
  IV U47426 ( .A(n37788), .Z(n34382) );
  NOR U47427 ( .A(n37790), .B(n34382), .Z(n34396) );
  NOR U47428 ( .A(n34383), .B(n34396), .Z(n34384) );
  XOR U47429 ( .A(n34398), .B(n34384), .Z(n37835) );
  IV U47430 ( .A(n37835), .Z(n37816) );
  IV U47431 ( .A(n34385), .Z(n34387) );
  NOR U47432 ( .A(n34387), .B(n34386), .Z(n37787) );
  IV U47433 ( .A(n37787), .Z(n34388) );
  NOR U47434 ( .A(n37790), .B(n34388), .Z(n37834) );
  IV U47435 ( .A(n37834), .Z(n37815) );
  NOR U47436 ( .A(n37816), .B(n37815), .Z(n37783) );
  IV U47437 ( .A(n37783), .Z(n34389) );
  NOR U47438 ( .A(n34395), .B(n34389), .Z(n37952) );
  IV U47439 ( .A(n34390), .Z(n34391) );
  NOR U47440 ( .A(n34392), .B(n34391), .Z(n34394) );
  IV U47441 ( .A(n34394), .Z(n34393) );
  NOR U47442 ( .A(n34395), .B(n34393), .Z(n41128) );
  XOR U47443 ( .A(n34395), .B(n34394), .Z(n37782) );
  IV U47444 ( .A(n34396), .Z(n34397) );
  NOR U47445 ( .A(n34398), .B(n34397), .Z(n37784) );
  IV U47446 ( .A(n37784), .Z(n34399) );
  NOR U47447 ( .A(n37782), .B(n34399), .Z(n37955) );
  NOR U47448 ( .A(n41128), .B(n37955), .Z(n37780) );
  IV U47449 ( .A(n34400), .Z(n34402) );
  NOR U47450 ( .A(n34402), .B(n34401), .Z(n37958) );
  IV U47451 ( .A(n34403), .Z(n34405) );
  NOR U47452 ( .A(n34405), .B(n34404), .Z(n41125) );
  NOR U47453 ( .A(n37958), .B(n41125), .Z(n37779) );
  IV U47454 ( .A(n34406), .Z(n34407) );
  NOR U47455 ( .A(n34407), .B(n34410), .Z(n34408) );
  IV U47456 ( .A(n34408), .Z(n41120) );
  IV U47457 ( .A(n34409), .Z(n34411) );
  NOR U47458 ( .A(n34411), .B(n34410), .Z(n37766) );
  IV U47459 ( .A(n34412), .Z(n34413) );
  NOR U47460 ( .A(n34414), .B(n34413), .Z(n37981) );
  IV U47461 ( .A(n34415), .Z(n34416) );
  NOR U47462 ( .A(n34416), .B(n37760), .Z(n37979) );
  NOR U47463 ( .A(n37981), .B(n37979), .Z(n37753) );
  IV U47464 ( .A(n34417), .Z(n34419) );
  IV U47465 ( .A(n34418), .Z(n37744) );
  NOR U47466 ( .A(n34419), .B(n37744), .Z(n41104) );
  IV U47467 ( .A(n34420), .Z(n34421) );
  NOR U47468 ( .A(n34421), .B(n37744), .Z(n37985) );
  IV U47469 ( .A(n34422), .Z(n34423) );
  NOR U47470 ( .A(n34426), .B(n34423), .Z(n37998) );
  IV U47471 ( .A(n34424), .Z(n34425) );
  NOR U47472 ( .A(n34426), .B(n34425), .Z(n37995) );
  IV U47473 ( .A(n34427), .Z(n34428) );
  NOR U47474 ( .A(n34428), .B(n37739), .Z(n41095) );
  NOR U47475 ( .A(n34430), .B(n34429), .Z(n41090) );
  IV U47476 ( .A(n34431), .Z(n34433) );
  NOR U47477 ( .A(n34433), .B(n34432), .Z(n41098) );
  NOR U47478 ( .A(n41090), .B(n41098), .Z(n37736) );
  IV U47479 ( .A(n34434), .Z(n34435) );
  NOR U47480 ( .A(n34435), .B(n34440), .Z(n38012) );
  IV U47481 ( .A(n34436), .Z(n34438) );
  NOR U47482 ( .A(n34438), .B(n34437), .Z(n41262) );
  IV U47483 ( .A(n34439), .Z(n34441) );
  NOR U47484 ( .A(n34441), .B(n34440), .Z(n44477) );
  NOR U47485 ( .A(n41262), .B(n44477), .Z(n41072) );
  NOR U47486 ( .A(n38017), .B(n34442), .Z(n37709) );
  IV U47487 ( .A(n34443), .Z(n34444) );
  NOR U47488 ( .A(n34445), .B(n34444), .Z(n41273) );
  NOR U47489 ( .A(n34446), .B(n41273), .Z(n41061) );
  NOR U47490 ( .A(n34448), .B(n34447), .Z(n41058) );
  NOR U47491 ( .A(n41058), .B(n41062), .Z(n37708) );
  IV U47492 ( .A(n34449), .Z(n34450) );
  NOR U47493 ( .A(n34451), .B(n34450), .Z(n38032) );
  IV U47494 ( .A(n34452), .Z(n34453) );
  NOR U47495 ( .A(n34456), .B(n34453), .Z(n41041) );
  IV U47496 ( .A(n34454), .Z(n34455) );
  NOR U47497 ( .A(n34456), .B(n34455), .Z(n41038) );
  IV U47498 ( .A(n34457), .Z(n34463) );
  NOR U47499 ( .A(n34458), .B(n34468), .Z(n34459) );
  IV U47500 ( .A(n34459), .Z(n34460) );
  NOR U47501 ( .A(n34461), .B(n34460), .Z(n34462) );
  IV U47502 ( .A(n34462), .Z(n34465) );
  NOR U47503 ( .A(n34463), .B(n34465), .Z(n38040) );
  NOR U47504 ( .A(n41038), .B(n38040), .Z(n37682) );
  IV U47505 ( .A(n34464), .Z(n34466) );
  NOR U47506 ( .A(n34466), .B(n34465), .Z(n38037) );
  IV U47507 ( .A(n34467), .Z(n34469) );
  NOR U47508 ( .A(n34469), .B(n34468), .Z(n38045) );
  IV U47509 ( .A(n34470), .Z(n34475) );
  IV U47510 ( .A(n34471), .Z(n34472) );
  NOR U47511 ( .A(n34475), .B(n34472), .Z(n38042) );
  IV U47512 ( .A(n34473), .Z(n34474) );
  NOR U47513 ( .A(n34475), .B(n34474), .Z(n38051) );
  IV U47514 ( .A(n34476), .Z(n34477) );
  NOR U47515 ( .A(n34478), .B(n34477), .Z(n38048) );
  IV U47516 ( .A(n34479), .Z(n34480) );
  NOR U47517 ( .A(n34480), .B(n37679), .Z(n41027) );
  IV U47518 ( .A(n34481), .Z(n34483) );
  IV U47519 ( .A(n34482), .Z(n34485) );
  NOR U47520 ( .A(n34483), .B(n34485), .Z(n41011) );
  IV U47521 ( .A(n34484), .Z(n34486) );
  NOR U47522 ( .A(n34486), .B(n34485), .Z(n41328) );
  NOR U47523 ( .A(n41011), .B(n41328), .Z(n37660) );
  IV U47524 ( .A(n34487), .Z(n34488) );
  NOR U47525 ( .A(n34488), .B(n37657), .Z(n34489) );
  IV U47526 ( .A(n34489), .Z(n41002) );
  IV U47527 ( .A(n34490), .Z(n34491) );
  NOR U47528 ( .A(n34492), .B(n34491), .Z(n38064) );
  IV U47529 ( .A(n34493), .Z(n34494) );
  NOR U47530 ( .A(n34495), .B(n34494), .Z(n34496) );
  IV U47531 ( .A(n34496), .Z(n40972) );
  IV U47532 ( .A(n34497), .Z(n34499) );
  NOR U47533 ( .A(n34499), .B(n34498), .Z(n40965) );
  IV U47534 ( .A(n34500), .Z(n34501) );
  NOR U47535 ( .A(n34508), .B(n34501), .Z(n34502) );
  IV U47536 ( .A(n34502), .Z(n34503) );
  NOR U47537 ( .A(n34504), .B(n34503), .Z(n40962) );
  IV U47538 ( .A(n34504), .Z(n34506) );
  NOR U47539 ( .A(n34506), .B(n34505), .Z(n34507) );
  IV U47540 ( .A(n34507), .Z(n34512) );
  NOR U47541 ( .A(n34509), .B(n34508), .Z(n34510) );
  IV U47542 ( .A(n34510), .Z(n34511) );
  NOR U47543 ( .A(n34512), .B(n34511), .Z(n38079) );
  IV U47544 ( .A(n34513), .Z(n34514) );
  NOR U47545 ( .A(n34517), .B(n34514), .Z(n40958) );
  NOR U47546 ( .A(n38079), .B(n40958), .Z(n37623) );
  IV U47547 ( .A(n34515), .Z(n34516) );
  NOR U47548 ( .A(n34517), .B(n34516), .Z(n40955) );
  IV U47549 ( .A(n34518), .Z(n34520) );
  NOR U47550 ( .A(n34520), .B(n34519), .Z(n38096) );
  IV U47551 ( .A(n34521), .Z(n34522) );
  NOR U47552 ( .A(n34522), .B(n37607), .Z(n38094) );
  NOR U47553 ( .A(n38096), .B(n38094), .Z(n37605) );
  IV U47554 ( .A(n34523), .Z(n34525) );
  IV U47555 ( .A(n34524), .Z(n34528) );
  NOR U47556 ( .A(n34525), .B(n34528), .Z(n40944) );
  NOR U47557 ( .A(n34526), .B(n40938), .Z(n34530) );
  IV U47558 ( .A(n34527), .Z(n34529) );
  NOR U47559 ( .A(n34529), .B(n34528), .Z(n40947) );
  NOR U47560 ( .A(n34530), .B(n40947), .Z(n37604) );
  IV U47561 ( .A(n34531), .Z(n34532) );
  NOR U47562 ( .A(n34533), .B(n34532), .Z(n40932) );
  IV U47563 ( .A(n34534), .Z(n34536) );
  NOR U47564 ( .A(n34536), .B(n34535), .Z(n38099) );
  NOR U47565 ( .A(n40932), .B(n38099), .Z(n37603) );
  IV U47566 ( .A(n34537), .Z(n34540) );
  IV U47567 ( .A(n34538), .Z(n34539) );
  NOR U47568 ( .A(n34540), .B(n34539), .Z(n40929) );
  IV U47569 ( .A(n34541), .Z(n34544) );
  IV U47570 ( .A(n34542), .Z(n34543) );
  NOR U47571 ( .A(n34544), .B(n34543), .Z(n40917) );
  NOR U47572 ( .A(n34546), .B(n34545), .Z(n38110) );
  IV U47573 ( .A(n34547), .Z(n34549) );
  NOR U47574 ( .A(n34549), .B(n34548), .Z(n38114) );
  NOR U47575 ( .A(n38110), .B(n38114), .Z(n34550) );
  IV U47576 ( .A(n34550), .Z(n34551) );
  NOR U47577 ( .A(n40913), .B(n34551), .Z(n37591) );
  IV U47578 ( .A(n34552), .Z(n34553) );
  NOR U47579 ( .A(n34554), .B(n34553), .Z(n41411) );
  IV U47580 ( .A(n34555), .Z(n34556) );
  NOR U47581 ( .A(n34556), .B(n34562), .Z(n41416) );
  NOR U47582 ( .A(n41411), .B(n41416), .Z(n38113) );
  IV U47583 ( .A(n34557), .Z(n34558) );
  NOR U47584 ( .A(n34559), .B(n34558), .Z(n40894) );
  IV U47585 ( .A(n34560), .Z(n34561) );
  NOR U47586 ( .A(n34562), .B(n34561), .Z(n38117) );
  NOR U47587 ( .A(n40894), .B(n38117), .Z(n37590) );
  IV U47588 ( .A(n34563), .Z(n34564) );
  NOR U47589 ( .A(n37588), .B(n34564), .Z(n40899) );
  IV U47590 ( .A(n34565), .Z(n34566) );
  NOR U47591 ( .A(n34567), .B(n34566), .Z(n41432) );
  IV U47592 ( .A(n34568), .Z(n34570) );
  NOR U47593 ( .A(n34570), .B(n34569), .Z(n41427) );
  NOR U47594 ( .A(n41432), .B(n41427), .Z(n38132) );
  NOR U47595 ( .A(n34571), .B(n34573), .Z(n38129) );
  IV U47596 ( .A(n34572), .Z(n34574) );
  NOR U47597 ( .A(n34574), .B(n34573), .Z(n38137) );
  IV U47598 ( .A(n34575), .Z(n34585) );
  XOR U47599 ( .A(n34576), .B(n34585), .Z(n34580) );
  IV U47600 ( .A(n34577), .Z(n34578) );
  NOR U47601 ( .A(n34580), .B(n34578), .Z(n38134) );
  NOR U47602 ( .A(n34580), .B(n34579), .Z(n34581) );
  IV U47603 ( .A(n34581), .Z(n34582) );
  NOR U47604 ( .A(n34584), .B(n34582), .Z(n38140) );
  IV U47605 ( .A(n34583), .Z(n34587) );
  NOR U47606 ( .A(n34585), .B(n34584), .Z(n34586) );
  IV U47607 ( .A(n34586), .Z(n34589) );
  NOR U47608 ( .A(n34587), .B(n34589), .Z(n38143) );
  IV U47609 ( .A(n34588), .Z(n34590) );
  NOR U47610 ( .A(n34590), .B(n34589), .Z(n38146) );
  IV U47611 ( .A(n34591), .Z(n34594) );
  NOR U47612 ( .A(n37574), .B(n34592), .Z(n34593) );
  IV U47613 ( .A(n34593), .Z(n34596) );
  NOR U47614 ( .A(n34594), .B(n34596), .Z(n38154) );
  IV U47615 ( .A(n34595), .Z(n34597) );
  NOR U47616 ( .A(n34597), .B(n34596), .Z(n38151) );
  IV U47617 ( .A(n34598), .Z(n34602) );
  NOR U47618 ( .A(n34600), .B(n34599), .Z(n34601) );
  IV U47619 ( .A(n34601), .Z(n37569) );
  NOR U47620 ( .A(n34602), .B(n37569), .Z(n40878) );
  IV U47621 ( .A(n34606), .Z(n34603) );
  NOR U47622 ( .A(n34603), .B(n34605), .Z(n44299) );
  IV U47623 ( .A(n34604), .Z(n34608) );
  XOR U47624 ( .A(n34606), .B(n34605), .Z(n34607) );
  NOR U47625 ( .A(n34608), .B(n34607), .Z(n41454) );
  NOR U47626 ( .A(n44299), .B(n41454), .Z(n40869) );
  IV U47627 ( .A(n34609), .Z(n34611) );
  NOR U47628 ( .A(n34611), .B(n34610), .Z(n40860) );
  NOR U47629 ( .A(n40860), .B(n40856), .Z(n34612) );
  IV U47630 ( .A(n34612), .Z(n34613) );
  NOR U47631 ( .A(n38162), .B(n34613), .Z(n37561) );
  IV U47632 ( .A(n34614), .Z(n34619) );
  IV U47633 ( .A(n34615), .Z(n34616) );
  NOR U47634 ( .A(n34619), .B(n34616), .Z(n40842) );
  IV U47635 ( .A(n34617), .Z(n34618) );
  NOR U47636 ( .A(n34619), .B(n34618), .Z(n38165) );
  IV U47637 ( .A(n34620), .Z(n34621) );
  NOR U47638 ( .A(n34625), .B(n34621), .Z(n38172) );
  IV U47639 ( .A(n34622), .Z(n34623) );
  NOR U47640 ( .A(n34623), .B(n34625), .Z(n38169) );
  IV U47641 ( .A(n34624), .Z(n34626) );
  NOR U47642 ( .A(n34626), .B(n34625), .Z(n38175) );
  NOR U47643 ( .A(n34627), .B(n38182), .Z(n34631) );
  IV U47644 ( .A(n34628), .Z(n34629) );
  NOR U47645 ( .A(n34630), .B(n34629), .Z(n38179) );
  NOR U47646 ( .A(n34631), .B(n38179), .Z(n37560) );
  IV U47647 ( .A(n34632), .Z(n34634) );
  NOR U47648 ( .A(n34634), .B(n34633), .Z(n38195) );
  IV U47649 ( .A(n34635), .Z(n34637) );
  NOR U47650 ( .A(n34637), .B(n34636), .Z(n38189) );
  NOR U47651 ( .A(n38195), .B(n38189), .Z(n37559) );
  IV U47652 ( .A(n34638), .Z(n34639) );
  NOR U47653 ( .A(n34639), .B(n41476), .Z(n40832) );
  NOR U47654 ( .A(n34640), .B(n38192), .Z(n34641) );
  NOR U47655 ( .A(n40832), .B(n34641), .Z(n34642) );
  IV U47656 ( .A(n34642), .Z(n34645) );
  IV U47657 ( .A(n34643), .Z(n34644) );
  NOR U47658 ( .A(n34644), .B(n41476), .Z(n38201) );
  NOR U47659 ( .A(n34645), .B(n38201), .Z(n37558) );
  IV U47660 ( .A(n34646), .Z(n34647) );
  NOR U47661 ( .A(n34648), .B(n34647), .Z(n38202) );
  IV U47662 ( .A(n34649), .Z(n34650) );
  NOR U47663 ( .A(n34650), .B(n34652), .Z(n38207) );
  NOR U47664 ( .A(n38202), .B(n38207), .Z(n37557) );
  IV U47665 ( .A(n34651), .Z(n34653) );
  NOR U47666 ( .A(n34653), .B(n34652), .Z(n38204) );
  IV U47667 ( .A(n34654), .Z(n34667) );
  IV U47668 ( .A(n34655), .Z(n34656) );
  NOR U47669 ( .A(n34667), .B(n34656), .Z(n44248) );
  IV U47670 ( .A(n34657), .Z(n34659) );
  NOR U47671 ( .A(n34659), .B(n34658), .Z(n44257) );
  NOR U47672 ( .A(n44248), .B(n44257), .Z(n38211) );
  IV U47673 ( .A(n34660), .Z(n34661) );
  NOR U47674 ( .A(n34664), .B(n34661), .Z(n38214) );
  IV U47675 ( .A(n34662), .Z(n34663) );
  NOR U47676 ( .A(n34664), .B(n34663), .Z(n40824) );
  NOR U47677 ( .A(n38214), .B(n40824), .Z(n34665) );
  IV U47678 ( .A(n34665), .Z(n34669) );
  IV U47679 ( .A(n34666), .Z(n34668) );
  NOR U47680 ( .A(n34668), .B(n34667), .Z(n38212) );
  NOR U47681 ( .A(n34669), .B(n38212), .Z(n37556) );
  IV U47682 ( .A(n34670), .Z(n34672) );
  IV U47683 ( .A(n34671), .Z(n37549) );
  NOR U47684 ( .A(n34672), .B(n37549), .Z(n40821) );
  IV U47685 ( .A(n34673), .Z(n34674) );
  NOR U47686 ( .A(n34675), .B(n34674), .Z(n40812) );
  IV U47687 ( .A(n34676), .Z(n34677) );
  NOR U47688 ( .A(n34677), .B(n34681), .Z(n40809) );
  IV U47689 ( .A(n34678), .Z(n34680) );
  NOR U47690 ( .A(n34680), .B(n34679), .Z(n38241) );
  NOR U47691 ( .A(n34682), .B(n34681), .Z(n34683) );
  IV U47692 ( .A(n34683), .Z(n34684) );
  NOR U47693 ( .A(n34685), .B(n34684), .Z(n38237) );
  NOR U47694 ( .A(n38241), .B(n38237), .Z(n37520) );
  XOR U47695 ( .A(n34687), .B(n34686), .Z(n34693) );
  IV U47696 ( .A(n34688), .Z(n34689) );
  NOR U47697 ( .A(n34690), .B(n34689), .Z(n34691) );
  IV U47698 ( .A(n34691), .Z(n34692) );
  NOR U47699 ( .A(n34693), .B(n34692), .Z(n40799) );
  IV U47700 ( .A(n34694), .Z(n34696) );
  IV U47701 ( .A(n34695), .Z(n34703) );
  NOR U47702 ( .A(n34696), .B(n34703), .Z(n44167) );
  IV U47703 ( .A(n34697), .Z(n34698) );
  NOR U47704 ( .A(n34698), .B(n44182), .Z(n34699) );
  NOR U47705 ( .A(n44167), .B(n34699), .Z(n40798) );
  IV U47706 ( .A(n40798), .Z(n34700) );
  NOR U47707 ( .A(n34700), .B(n40802), .Z(n37512) );
  IV U47708 ( .A(n34701), .Z(n34702) );
  NOR U47709 ( .A(n34703), .B(n34702), .Z(n40788) );
  IV U47710 ( .A(n34704), .Z(n34705) );
  NOR U47711 ( .A(n34705), .B(n37503), .Z(n40784) );
  IV U47712 ( .A(n34706), .Z(n34708) );
  NOR U47713 ( .A(n34708), .B(n34707), .Z(n34709) );
  IV U47714 ( .A(n34709), .Z(n37491) );
  IV U47715 ( .A(n34710), .Z(n34711) );
  NOR U47716 ( .A(n34714), .B(n34711), .Z(n40770) );
  IV U47717 ( .A(n34712), .Z(n34713) );
  NOR U47718 ( .A(n34714), .B(n34713), .Z(n40767) );
  IV U47719 ( .A(n34715), .Z(n34717) );
  IV U47720 ( .A(n34716), .Z(n37471) );
  NOR U47721 ( .A(n34717), .B(n37471), .Z(n40760) );
  IV U47722 ( .A(n34718), .Z(n34719) );
  NOR U47723 ( .A(n37433), .B(n34719), .Z(n37437) );
  IV U47724 ( .A(n37437), .Z(n37435) );
  NOR U47725 ( .A(n34721), .B(n34720), .Z(n34722) );
  NOR U47726 ( .A(n34722), .B(n34721), .Z(n38279) );
  IV U47727 ( .A(n34723), .Z(n34724) );
  NOR U47728 ( .A(n34725), .B(n34724), .Z(n40712) );
  IV U47729 ( .A(n34726), .Z(n34727) );
  NOR U47730 ( .A(n34727), .B(n37426), .Z(n40716) );
  NOR U47731 ( .A(n40712), .B(n40716), .Z(n38283) );
  IV U47732 ( .A(n34728), .Z(n34730) );
  XOR U47733 ( .A(n34737), .B(n34738), .Z(n34729) );
  NOR U47734 ( .A(n34730), .B(n34729), .Z(n40699) );
  IV U47735 ( .A(n34731), .Z(n34734) );
  IV U47736 ( .A(n34732), .Z(n34733) );
  NOR U47737 ( .A(n34734), .B(n34733), .Z(n40702) );
  IV U47738 ( .A(n34735), .Z(n34736) );
  NOR U47739 ( .A(n34736), .B(n34738), .Z(n40697) );
  IV U47740 ( .A(n34737), .Z(n34739) );
  NOR U47741 ( .A(n34739), .B(n34738), .Z(n38286) );
  NOR U47742 ( .A(n40697), .B(n38286), .Z(n34740) );
  IV U47743 ( .A(n34740), .Z(n34741) );
  NOR U47744 ( .A(n40702), .B(n34741), .Z(n37417) );
  IV U47745 ( .A(n34742), .Z(n34744) );
  NOR U47746 ( .A(n34744), .B(n34743), .Z(n37412) );
  IV U47747 ( .A(n34745), .Z(n34747) );
  NOR U47748 ( .A(n34747), .B(n34746), .Z(n37409) );
  IV U47749 ( .A(n37409), .Z(n37399) );
  IV U47750 ( .A(n34748), .Z(n38292) );
  NOR U47751 ( .A(n34749), .B(n38292), .Z(n37398) );
  IV U47752 ( .A(n34750), .Z(n34751) );
  NOR U47753 ( .A(n37396), .B(n34751), .Z(n40691) );
  NOR U47754 ( .A(n34753), .B(n34752), .Z(n34754) );
  IV U47755 ( .A(n34754), .Z(n38301) );
  IV U47756 ( .A(n34755), .Z(n34762) );
  NOR U47757 ( .A(n34757), .B(n34756), .Z(n34758) );
  IV U47758 ( .A(n34758), .Z(n34759) );
  NOR U47759 ( .A(n34760), .B(n34759), .Z(n34761) );
  IV U47760 ( .A(n34761), .Z(n37372) );
  NOR U47761 ( .A(n34762), .B(n37372), .Z(n38305) );
  IV U47762 ( .A(n34763), .Z(n34767) );
  NOR U47763 ( .A(n34765), .B(n34764), .Z(n34766) );
  IV U47764 ( .A(n34766), .Z(n34770) );
  NOR U47765 ( .A(n34767), .B(n34770), .Z(n38311) );
  NOR U47766 ( .A(n34768), .B(n38320), .Z(n34772) );
  IV U47767 ( .A(n34769), .Z(n34771) );
  NOR U47768 ( .A(n34771), .B(n34770), .Z(n38315) );
  NOR U47769 ( .A(n34772), .B(n38315), .Z(n37370) );
  IV U47770 ( .A(n34773), .Z(n34775) );
  NOR U47771 ( .A(n34775), .B(n34774), .Z(n40656) );
  IV U47772 ( .A(n34776), .Z(n34778) );
  NOR U47773 ( .A(n34778), .B(n34777), .Z(n40663) );
  NOR U47774 ( .A(n40656), .B(n40663), .Z(n37362) );
  IV U47775 ( .A(n34779), .Z(n34780) );
  NOR U47776 ( .A(n34780), .B(n34782), .Z(n38334) );
  IV U47777 ( .A(n34781), .Z(n34783) );
  NOR U47778 ( .A(n34783), .B(n34782), .Z(n38331) );
  IV U47779 ( .A(n34784), .Z(n37357) );
  IV U47780 ( .A(n34785), .Z(n34786) );
  NOR U47781 ( .A(n37357), .B(n34786), .Z(n38337) );
  IV U47782 ( .A(n34787), .Z(n34788) );
  NOR U47783 ( .A(n34788), .B(n34794), .Z(n40644) );
  IV U47784 ( .A(n34789), .Z(n37342) );
  NOR U47785 ( .A(n34790), .B(n37342), .Z(n34791) );
  IV U47786 ( .A(n34791), .Z(n38345) );
  NOR U47787 ( .A(n34792), .B(n38345), .Z(n34796) );
  IV U47788 ( .A(n34793), .Z(n34795) );
  NOR U47789 ( .A(n34795), .B(n34794), .Z(n40647) );
  NOR U47790 ( .A(n34796), .B(n40647), .Z(n37354) );
  IV U47791 ( .A(n34797), .Z(n34802) );
  IV U47792 ( .A(n34798), .Z(n34799) );
  NOR U47793 ( .A(n34802), .B(n34799), .Z(n40635) );
  IV U47794 ( .A(n34800), .Z(n34801) );
  NOR U47795 ( .A(n34802), .B(n34801), .Z(n38358) );
  IV U47796 ( .A(n34803), .Z(n34804) );
  NOR U47797 ( .A(n38363), .B(n34804), .Z(n38355) );
  NOR U47798 ( .A(n34805), .B(n38363), .Z(n34806) );
  IV U47799 ( .A(n34806), .Z(n40626) );
  IV U47800 ( .A(n34807), .Z(n34808) );
  NOR U47801 ( .A(n34809), .B(n34808), .Z(n37338) );
  IV U47802 ( .A(n37338), .Z(n37329) );
  IV U47803 ( .A(n34810), .Z(n34811) );
  NOR U47804 ( .A(n34812), .B(n34811), .Z(n34813) );
  IV U47805 ( .A(n34813), .Z(n40618) );
  IV U47806 ( .A(n34814), .Z(n34815) );
  NOR U47807 ( .A(n34815), .B(n37321), .Z(n38367) );
  IV U47808 ( .A(n34816), .Z(n34817) );
  NOR U47809 ( .A(n34818), .B(n34817), .Z(n41609) );
  IV U47810 ( .A(n34819), .Z(n34825) );
  NOR U47811 ( .A(n34821), .B(n34820), .Z(n34822) );
  IV U47812 ( .A(n34822), .Z(n37297) );
  NOR U47813 ( .A(n34823), .B(n37297), .Z(n34824) );
  IV U47814 ( .A(n34824), .Z(n34827) );
  NOR U47815 ( .A(n34825), .B(n34827), .Z(n41614) );
  NOR U47816 ( .A(n41609), .B(n41614), .Z(n40612) );
  IV U47817 ( .A(n34826), .Z(n34828) );
  NOR U47818 ( .A(n34828), .B(n34827), .Z(n38383) );
  IV U47819 ( .A(n34829), .Z(n34830) );
  NOR U47820 ( .A(n34831), .B(n34830), .Z(n37293) );
  IV U47821 ( .A(n34832), .Z(n34834) );
  NOR U47822 ( .A(n34834), .B(n34833), .Z(n40607) );
  NOR U47823 ( .A(n34835), .B(n41628), .Z(n38393) );
  NOR U47824 ( .A(n40607), .B(n38393), .Z(n37291) );
  IV U47825 ( .A(n34836), .Z(n34837) );
  NOR U47826 ( .A(n34838), .B(n34837), .Z(n34839) );
  IV U47827 ( .A(n34839), .Z(n37287) );
  IV U47828 ( .A(n34840), .Z(n34844) );
  NOR U47829 ( .A(n34842), .B(n34841), .Z(n34843) );
  IV U47830 ( .A(n34843), .Z(n37285) );
  NOR U47831 ( .A(n34844), .B(n37285), .Z(n40601) );
  IV U47832 ( .A(n34845), .Z(n34847) );
  NOR U47833 ( .A(n34847), .B(n34846), .Z(n40597) );
  IV U47834 ( .A(n34848), .Z(n34849) );
  NOR U47835 ( .A(n34849), .B(n37275), .Z(n40594) );
  IV U47836 ( .A(n34850), .Z(n34852) );
  NOR U47837 ( .A(n34852), .B(n34851), .Z(n40579) );
  IV U47838 ( .A(n37282), .Z(n34853) );
  NOR U47839 ( .A(n37278), .B(n34853), .Z(n34854) );
  IV U47840 ( .A(n34854), .Z(n34859) );
  NOR U47841 ( .A(n34856), .B(n34855), .Z(n34857) );
  IV U47842 ( .A(n34857), .Z(n34858) );
  NOR U47843 ( .A(n34859), .B(n34858), .Z(n38400) );
  NOR U47844 ( .A(n40579), .B(n38400), .Z(n37273) );
  IV U47845 ( .A(n34860), .Z(n34861) );
  NOR U47846 ( .A(n34862), .B(n34861), .Z(n43962) );
  IV U47847 ( .A(n34863), .Z(n34864) );
  NOR U47848 ( .A(n34864), .B(n37264), .Z(n43967) );
  NOR U47849 ( .A(n43962), .B(n43967), .Z(n38409) );
  IV U47850 ( .A(n34865), .Z(n34867) );
  NOR U47851 ( .A(n34867), .B(n34866), .Z(n38420) );
  NOR U47852 ( .A(n38420), .B(n40560), .Z(n37247) );
  IV U47853 ( .A(n34868), .Z(n34870) );
  NOR U47854 ( .A(n34870), .B(n34869), .Z(n34871) );
  IV U47855 ( .A(n34871), .Z(n38422) );
  IV U47856 ( .A(n34872), .Z(n34873) );
  NOR U47857 ( .A(n34873), .B(n37242), .Z(n34874) );
  IV U47858 ( .A(n34874), .Z(n34875) );
  NOR U47859 ( .A(n34876), .B(n34875), .Z(n40549) );
  IV U47860 ( .A(n34877), .Z(n34879) );
  NOR U47861 ( .A(n34879), .B(n34878), .Z(n40539) );
  IV U47862 ( .A(n34880), .Z(n34881) );
  NOR U47863 ( .A(n34882), .B(n34881), .Z(n40546) );
  NOR U47864 ( .A(n40539), .B(n40546), .Z(n37238) );
  NOR U47865 ( .A(n34883), .B(n40535), .Z(n37237) );
  IV U47866 ( .A(n34884), .Z(n34886) );
  NOR U47867 ( .A(n34886), .B(n34885), .Z(n38423) );
  IV U47868 ( .A(n34887), .Z(n34888) );
  NOR U47869 ( .A(n34889), .B(n34888), .Z(n40531) );
  NOR U47870 ( .A(n38423), .B(n40531), .Z(n37235) );
  IV U47871 ( .A(n34890), .Z(n34891) );
  NOR U47872 ( .A(n34892), .B(n34891), .Z(n41707) );
  IV U47873 ( .A(n34893), .Z(n34895) );
  NOR U47874 ( .A(n34895), .B(n34894), .Z(n41697) );
  NOR U47875 ( .A(n41707), .B(n41697), .Z(n40507) );
  IV U47876 ( .A(n34896), .Z(n34897) );
  NOR U47877 ( .A(n34897), .B(n34909), .Z(n41714) );
  XOR U47878 ( .A(n34899), .B(n34898), .Z(n34902) );
  IV U47879 ( .A(n34900), .Z(n34901) );
  NOR U47880 ( .A(n34902), .B(n34901), .Z(n41710) );
  NOR U47881 ( .A(n41714), .B(n41710), .Z(n38435) );
  IV U47882 ( .A(n38435), .Z(n41698) );
  IV U47883 ( .A(n34903), .Z(n34904) );
  NOR U47884 ( .A(n34904), .B(n34909), .Z(n38432) );
  IV U47885 ( .A(n34905), .Z(n34907) );
  NOR U47886 ( .A(n34907), .B(n34906), .Z(n38439) );
  IV U47887 ( .A(n34908), .Z(n34910) );
  NOR U47888 ( .A(n34910), .B(n34909), .Z(n38436) );
  NOR U47889 ( .A(n38439), .B(n38436), .Z(n37221) );
  IV U47890 ( .A(n34911), .Z(n34914) );
  NOR U47891 ( .A(n34920), .B(n34912), .Z(n34913) );
  IV U47892 ( .A(n34913), .Z(n34917) );
  NOR U47893 ( .A(n34914), .B(n34917), .Z(n34915) );
  IV U47894 ( .A(n34915), .Z(n40501) );
  IV U47895 ( .A(n34916), .Z(n34918) );
  NOR U47896 ( .A(n34918), .B(n34917), .Z(n37217) );
  NOR U47897 ( .A(n34920), .B(n34919), .Z(n37214) );
  IV U47898 ( .A(n37214), .Z(n37209) );
  IV U47899 ( .A(n34921), .Z(n34922) );
  NOR U47900 ( .A(n34922), .B(n34924), .Z(n40489) );
  IV U47901 ( .A(n34923), .Z(n34925) );
  NOR U47902 ( .A(n34925), .B(n34924), .Z(n38445) );
  IV U47903 ( .A(n34926), .Z(n34927) );
  NOR U47904 ( .A(n34928), .B(n34927), .Z(n40481) );
  IV U47905 ( .A(n34929), .Z(n34931) );
  NOR U47906 ( .A(n34931), .B(n34930), .Z(n38448) );
  NOR U47907 ( .A(n40481), .B(n38448), .Z(n37204) );
  IV U47908 ( .A(n34932), .Z(n34939) );
  NOR U47909 ( .A(n34934), .B(n34933), .Z(n34935) );
  IV U47910 ( .A(n34935), .Z(n34936) );
  NOR U47911 ( .A(n34937), .B(n34936), .Z(n34938) );
  IV U47912 ( .A(n34938), .Z(n34941) );
  NOR U47913 ( .A(n34939), .B(n34941), .Z(n40478) );
  IV U47914 ( .A(n34940), .Z(n34942) );
  NOR U47915 ( .A(n34942), .B(n34941), .Z(n38450) );
  IV U47916 ( .A(n34943), .Z(n34946) );
  IV U47917 ( .A(n34944), .Z(n34945) );
  NOR U47918 ( .A(n34946), .B(n34945), .Z(n38456) );
  IV U47919 ( .A(n34947), .Z(n34948) );
  NOR U47920 ( .A(n34948), .B(n34952), .Z(n38453) );
  IV U47921 ( .A(n34949), .Z(n34950) );
  NOR U47922 ( .A(n34950), .B(n34952), .Z(n38462) );
  IV U47923 ( .A(n34951), .Z(n34953) );
  NOR U47924 ( .A(n34953), .B(n34952), .Z(n38459) );
  IV U47925 ( .A(n34954), .Z(n34958) );
  NOR U47926 ( .A(n34956), .B(n34955), .Z(n34957) );
  IV U47927 ( .A(n34957), .Z(n37195) );
  NOR U47928 ( .A(n34958), .B(n37195), .Z(n38465) );
  IV U47929 ( .A(n34959), .Z(n34961) );
  NOR U47930 ( .A(n34961), .B(n34960), .Z(n38470) );
  IV U47931 ( .A(n34962), .Z(n34966) );
  NOR U47932 ( .A(n34964), .B(n34963), .Z(n34965) );
  IV U47933 ( .A(n34965), .Z(n37192) );
  NOR U47934 ( .A(n34966), .B(n37192), .Z(n40466) );
  IV U47935 ( .A(n34967), .Z(n34969) );
  NOR U47936 ( .A(n34969), .B(n34968), .Z(n38476) );
  IV U47937 ( .A(n34970), .Z(n34977) );
  NOR U47938 ( .A(n34977), .B(n34971), .Z(n34972) );
  IV U47939 ( .A(n34972), .Z(n34973) );
  NOR U47940 ( .A(n34974), .B(n34973), .Z(n40462) );
  IV U47941 ( .A(n34975), .Z(n34976) );
  NOR U47942 ( .A(n34977), .B(n34976), .Z(n40459) );
  IV U47943 ( .A(n34978), .Z(n34979) );
  NOR U47944 ( .A(n34979), .B(n34981), .Z(n40455) );
  IV U47945 ( .A(n34980), .Z(n34987) );
  NOR U47946 ( .A(n34982), .B(n34981), .Z(n34983) );
  IV U47947 ( .A(n34983), .Z(n34984) );
  NOR U47948 ( .A(n34985), .B(n34984), .Z(n34986) );
  IV U47949 ( .A(n34986), .Z(n37186) );
  NOR U47950 ( .A(n34987), .B(n37186), .Z(n40447) );
  IV U47951 ( .A(n34988), .Z(n34995) );
  NOR U47952 ( .A(n34990), .B(n34989), .Z(n34991) );
  IV U47953 ( .A(n34991), .Z(n34992) );
  NOR U47954 ( .A(n34993), .B(n34992), .Z(n34994) );
  IV U47955 ( .A(n34994), .Z(n37179) );
  NOR U47956 ( .A(n34995), .B(n37179), .Z(n37172) );
  IV U47957 ( .A(n34996), .Z(n34997) );
  NOR U47958 ( .A(n34997), .B(n35002), .Z(n40439) );
  IV U47959 ( .A(n34998), .Z(n35000) );
  NOR U47960 ( .A(n35000), .B(n34999), .Z(n40431) );
  IV U47961 ( .A(n35001), .Z(n35003) );
  NOR U47962 ( .A(n35003), .B(n35002), .Z(n40436) );
  NOR U47963 ( .A(n40431), .B(n40436), .Z(n37165) );
  IV U47964 ( .A(n35004), .Z(n35005) );
  NOR U47965 ( .A(n35005), .B(n37156), .Z(n43855) );
  IV U47966 ( .A(n35006), .Z(n35008) );
  IV U47967 ( .A(n35007), .Z(n37161) );
  NOR U47968 ( .A(n35008), .B(n37161), .Z(n41774) );
  NOR U47969 ( .A(n43855), .B(n41774), .Z(n40419) );
  IV U47970 ( .A(n35009), .Z(n35010) );
  NOR U47971 ( .A(n35011), .B(n35010), .Z(n38502) );
  IV U47972 ( .A(n35012), .Z(n35014) );
  NOR U47973 ( .A(n35014), .B(n35013), .Z(n38500) );
  NOR U47974 ( .A(n38502), .B(n38500), .Z(n37151) );
  IV U47975 ( .A(n35015), .Z(n35017) );
  NOR U47976 ( .A(n35017), .B(n35016), .Z(n40415) );
  IV U47977 ( .A(n35018), .Z(n35019) );
  NOR U47978 ( .A(n37140), .B(n35019), .Z(n38505) );
  IV U47979 ( .A(n35020), .Z(n35022) );
  IV U47980 ( .A(n35021), .Z(n37133) );
  NOR U47981 ( .A(n35022), .B(n37133), .Z(n38515) );
  IV U47982 ( .A(n35023), .Z(n35024) );
  NOR U47983 ( .A(n35025), .B(n35024), .Z(n38512) );
  IV U47984 ( .A(n35026), .Z(n35035) );
  NOR U47985 ( .A(n35027), .B(n35037), .Z(n35028) );
  IV U47986 ( .A(n35028), .Z(n35029) );
  NOR U47987 ( .A(n35030), .B(n35029), .Z(n35031) );
  IV U47988 ( .A(n35031), .Z(n35032) );
  NOR U47989 ( .A(n35033), .B(n35032), .Z(n35034) );
  IV U47990 ( .A(n35034), .Z(n37124) );
  NOR U47991 ( .A(n35035), .B(n37124), .Z(n40391) );
  IV U47992 ( .A(n35036), .Z(n35040) );
  NOR U47993 ( .A(n35038), .B(n35037), .Z(n35039) );
  IV U47994 ( .A(n35039), .Z(n37121) );
  NOR U47995 ( .A(n35040), .B(n37121), .Z(n38522) );
  IV U47996 ( .A(n35041), .Z(n35042) );
  NOR U47997 ( .A(n35043), .B(n35042), .Z(n38531) );
  IV U47998 ( .A(n35044), .Z(n35045) );
  NOR U47999 ( .A(n35045), .B(n35051), .Z(n38528) );
  IV U48000 ( .A(n35046), .Z(n35047) );
  NOR U48001 ( .A(n35048), .B(n35047), .Z(n40370) );
  IV U48002 ( .A(n35049), .Z(n35050) );
  NOR U48003 ( .A(n35051), .B(n35050), .Z(n40373) );
  NOR U48004 ( .A(n40370), .B(n40373), .Z(n37118) );
  IV U48005 ( .A(n35052), .Z(n35053) );
  NOR U48006 ( .A(n35056), .B(n35053), .Z(n40367) );
  IV U48007 ( .A(n35054), .Z(n35055) );
  NOR U48008 ( .A(n35056), .B(n35055), .Z(n40363) );
  IV U48009 ( .A(n35057), .Z(n35061) );
  NOR U48010 ( .A(n35059), .B(n35058), .Z(n35060) );
  IV U48011 ( .A(n35060), .Z(n35063) );
  NOR U48012 ( .A(n35061), .B(n35063), .Z(n40360) );
  IV U48013 ( .A(n35062), .Z(n35064) );
  NOR U48014 ( .A(n35064), .B(n35063), .Z(n40355) );
  IV U48015 ( .A(n35065), .Z(n35067) );
  IV U48016 ( .A(n35066), .Z(n37104) );
  NOR U48017 ( .A(n35067), .B(n37104), .Z(n37099) );
  IV U48018 ( .A(n35068), .Z(n35069) );
  NOR U48019 ( .A(n35069), .B(n35071), .Z(n38542) );
  IV U48020 ( .A(n35070), .Z(n35072) );
  NOR U48021 ( .A(n35072), .B(n35071), .Z(n40342) );
  NOR U48022 ( .A(n35073), .B(n35078), .Z(n35074) );
  IV U48023 ( .A(n35074), .Z(n35075) );
  NOR U48024 ( .A(n35076), .B(n35075), .Z(n40339) );
  IV U48025 ( .A(n35077), .Z(n35079) );
  NOR U48026 ( .A(n35079), .B(n35078), .Z(n38548) );
  IV U48027 ( .A(n35080), .Z(n35081) );
  NOR U48028 ( .A(n35082), .B(n35081), .Z(n41823) );
  IV U48029 ( .A(n35083), .Z(n35085) );
  NOR U48030 ( .A(n35085), .B(n35084), .Z(n43779) );
  NOR U48031 ( .A(n41823), .B(n43779), .Z(n38547) );
  IV U48032 ( .A(n35086), .Z(n35087) );
  NOR U48033 ( .A(n35088), .B(n35087), .Z(n37064) );
  IV U48034 ( .A(n35089), .Z(n35090) );
  NOR U48035 ( .A(n35092), .B(n35090), .Z(n37060) );
  IV U48036 ( .A(n35091), .Z(n35093) );
  NOR U48037 ( .A(n35093), .B(n35092), .Z(n38561) );
  IV U48038 ( .A(n35094), .Z(n35098) );
  NOR U48039 ( .A(n35098), .B(n35095), .Z(n43764) );
  NOR U48040 ( .A(n41846), .B(n43764), .Z(n38566) );
  IV U48041 ( .A(n38566), .Z(n35099) );
  IV U48042 ( .A(n35096), .Z(n35097) );
  NOR U48043 ( .A(n35098), .B(n35097), .Z(n38564) );
  NOR U48044 ( .A(n35099), .B(n38564), .Z(n37057) );
  IV U48045 ( .A(n35100), .Z(n35101) );
  NOR U48046 ( .A(n35101), .B(n37048), .Z(n40331) );
  IV U48047 ( .A(n35102), .Z(n35104) );
  NOR U48048 ( .A(n35104), .B(n35103), .Z(n43758) );
  IV U48049 ( .A(n35105), .Z(n35109) );
  NOR U48050 ( .A(n35106), .B(n37051), .Z(n35107) );
  IV U48051 ( .A(n35107), .Z(n35108) );
  NOR U48052 ( .A(n35109), .B(n35108), .Z(n41866) );
  NOR U48053 ( .A(n43758), .B(n41866), .Z(n38567) );
  IV U48054 ( .A(n35110), .Z(n35112) );
  NOR U48055 ( .A(n35112), .B(n35111), .Z(n41876) );
  NOR U48056 ( .A(n35114), .B(n35113), .Z(n41871) );
  NOR U48057 ( .A(n41876), .B(n41871), .Z(n40313) );
  IV U48058 ( .A(n35115), .Z(n35116) );
  NOR U48059 ( .A(n35116), .B(n35128), .Z(n40299) );
  NOR U48060 ( .A(n40305), .B(n40299), .Z(n37040) );
  IV U48061 ( .A(n35117), .Z(n35122) );
  IV U48062 ( .A(n35118), .Z(n35119) );
  NOR U48063 ( .A(n35119), .B(n35128), .Z(n35120) );
  IV U48064 ( .A(n35120), .Z(n35121) );
  NOR U48065 ( .A(n35122), .B(n35121), .Z(n40302) );
  IV U48066 ( .A(n35123), .Z(n35130) );
  NOR U48067 ( .A(n35125), .B(n35124), .Z(n35126) );
  IV U48068 ( .A(n35126), .Z(n35127) );
  NOR U48069 ( .A(n35128), .B(n35127), .Z(n35129) );
  IV U48070 ( .A(n35129), .Z(n37038) );
  NOR U48071 ( .A(n35130), .B(n37038), .Z(n40294) );
  IV U48072 ( .A(n35131), .Z(n35133) );
  NOR U48073 ( .A(n35133), .B(n35132), .Z(n40274) );
  IV U48074 ( .A(n35134), .Z(n35138) );
  NOR U48075 ( .A(n35136), .B(n35135), .Z(n35137) );
  IV U48076 ( .A(n35137), .Z(n37027) );
  NOR U48077 ( .A(n35138), .B(n37027), .Z(n40278) );
  NOR U48078 ( .A(n40274), .B(n40278), .Z(n37025) );
  IV U48079 ( .A(n35139), .Z(n35141) );
  NOR U48080 ( .A(n35141), .B(n35140), .Z(n35142) );
  NOR U48081 ( .A(n35142), .B(n43723), .Z(n40273) );
  NOR U48082 ( .A(n35144), .B(n35143), .Z(n40267) );
  IV U48083 ( .A(n35145), .Z(n35147) );
  NOR U48084 ( .A(n35147), .B(n35146), .Z(n45327) );
  IV U48085 ( .A(n35148), .Z(n35149) );
  NOR U48086 ( .A(n35149), .B(n36999), .Z(n45323) );
  NOR U48087 ( .A(n45327), .B(n45323), .Z(n40245) );
  IV U48088 ( .A(n35150), .Z(n35151) );
  NOR U48089 ( .A(n35152), .B(n35151), .Z(n38577) );
  IV U48090 ( .A(n35153), .Z(n35160) );
  IV U48091 ( .A(n35154), .Z(n36987) );
  NOR U48092 ( .A(n35155), .B(n36987), .Z(n35156) );
  IV U48093 ( .A(n35156), .Z(n35157) );
  NOR U48094 ( .A(n35158), .B(n35157), .Z(n35159) );
  IV U48095 ( .A(n35159), .Z(n35164) );
  NOR U48096 ( .A(n35160), .B(n35164), .Z(n38586) );
  IV U48097 ( .A(n35161), .Z(n35162) );
  NOR U48098 ( .A(n35162), .B(n35170), .Z(n38593) );
  IV U48099 ( .A(n35163), .Z(n35165) );
  NOR U48100 ( .A(n35165), .B(n35164), .Z(n38589) );
  NOR U48101 ( .A(n38593), .B(n38589), .Z(n36982) );
  IV U48102 ( .A(n35166), .Z(n35168) );
  NOR U48103 ( .A(n35168), .B(n35167), .Z(n43698) );
  IV U48104 ( .A(n35169), .Z(n35171) );
  NOR U48105 ( .A(n35171), .B(n35170), .Z(n41928) );
  NOR U48106 ( .A(n43698), .B(n41928), .Z(n38592) );
  IV U48107 ( .A(n35172), .Z(n35173) );
  NOR U48108 ( .A(n35174), .B(n35173), .Z(n40228) );
  IV U48109 ( .A(n35175), .Z(n35177) );
  NOR U48110 ( .A(n35177), .B(n35176), .Z(n38597) );
  NOR U48111 ( .A(n40228), .B(n38597), .Z(n36981) );
  IV U48112 ( .A(n35178), .Z(n35179) );
  NOR U48113 ( .A(n35179), .B(n36980), .Z(n40223) );
  IV U48114 ( .A(n35180), .Z(n35181) );
  NOR U48115 ( .A(n35182), .B(n35181), .Z(n36969) );
  IV U48116 ( .A(n36969), .Z(n36958) );
  NOR U48117 ( .A(n35183), .B(n41943), .Z(n36962) );
  IV U48118 ( .A(n35184), .Z(n35186) );
  NOR U48119 ( .A(n35186), .B(n35185), .Z(n38607) );
  NOR U48120 ( .A(n36962), .B(n38607), .Z(n36956) );
  IV U48121 ( .A(n35187), .Z(n35189) );
  NOR U48122 ( .A(n35189), .B(n35188), .Z(n40214) );
  IV U48123 ( .A(n35190), .Z(n35192) );
  NOR U48124 ( .A(n35192), .B(n35191), .Z(n38610) );
  NOR U48125 ( .A(n40214), .B(n38610), .Z(n36955) );
  IV U48126 ( .A(n35193), .Z(n35195) );
  NOR U48127 ( .A(n35195), .B(n35194), .Z(n35196) );
  IV U48128 ( .A(n35196), .Z(n36946) );
  IV U48129 ( .A(n35197), .Z(n35198) );
  NOR U48130 ( .A(n35199), .B(n35198), .Z(n35200) );
  IV U48131 ( .A(n35200), .Z(n40205) );
  NOR U48132 ( .A(n35202), .B(n35201), .Z(n40194) );
  IV U48133 ( .A(n35203), .Z(n35204) );
  NOR U48134 ( .A(n36932), .B(n35204), .Z(n36925) );
  IV U48135 ( .A(n35205), .Z(n35206) );
  NOR U48136 ( .A(n35207), .B(n35206), .Z(n36922) );
  IV U48137 ( .A(n36922), .Z(n36913) );
  IV U48138 ( .A(n35208), .Z(n35209) );
  NOR U48139 ( .A(n35210), .B(n35209), .Z(n38615) );
  IV U48140 ( .A(n35211), .Z(n35212) );
  NOR U48141 ( .A(n35213), .B(n35212), .Z(n38612) );
  IV U48142 ( .A(n35214), .Z(n35215) );
  NOR U48143 ( .A(n35216), .B(n35215), .Z(n38624) );
  NOR U48144 ( .A(n35217), .B(n36902), .Z(n35218) );
  IV U48145 ( .A(n35218), .Z(n35219) );
  NOR U48146 ( .A(n35220), .B(n35219), .Z(n40169) );
  IV U48147 ( .A(n35221), .Z(n35223) );
  IV U48148 ( .A(n35222), .Z(n35227) );
  NOR U48149 ( .A(n35223), .B(n35227), .Z(n40159) );
  IV U48150 ( .A(n35224), .Z(n35225) );
  NOR U48151 ( .A(n35225), .B(n35230), .Z(n40155) );
  IV U48152 ( .A(n35226), .Z(n35228) );
  NOR U48153 ( .A(n35228), .B(n35227), .Z(n40161) );
  NOR U48154 ( .A(n40155), .B(n40161), .Z(n36885) );
  IV U48155 ( .A(n35229), .Z(n35231) );
  NOR U48156 ( .A(n35231), .B(n35230), .Z(n40154) );
  IV U48157 ( .A(n40154), .Z(n40152) );
  IV U48158 ( .A(n35232), .Z(n35233) );
  NOR U48159 ( .A(n35236), .B(n35233), .Z(n38640) );
  IV U48160 ( .A(n35234), .Z(n35235) );
  NOR U48161 ( .A(n35236), .B(n35235), .Z(n36866) );
  IV U48162 ( .A(n35237), .Z(n35239) );
  NOR U48163 ( .A(n35239), .B(n35238), .Z(n36863) );
  IV U48164 ( .A(n36863), .Z(n36858) );
  IV U48165 ( .A(n35240), .Z(n35242) );
  IV U48166 ( .A(n35241), .Z(n36860) );
  NOR U48167 ( .A(n35242), .B(n36860), .Z(n40131) );
  NOR U48168 ( .A(n40127), .B(n40131), .Z(n36857) );
  IV U48169 ( .A(n35243), .Z(n36852) );
  IV U48170 ( .A(n35244), .Z(n35245) );
  NOR U48171 ( .A(n36840), .B(n35245), .Z(n38643) );
  IV U48172 ( .A(n35246), .Z(n35247) );
  NOR U48173 ( .A(n35248), .B(n35247), .Z(n35249) );
  IV U48174 ( .A(n35249), .Z(n36841) );
  IV U48175 ( .A(n35250), .Z(n35251) );
  NOR U48176 ( .A(n35251), .B(n36836), .Z(n38657) );
  IV U48177 ( .A(n35252), .Z(n35253) );
  NOR U48178 ( .A(n35253), .B(n36836), .Z(n35254) );
  IV U48179 ( .A(n35254), .Z(n38656) );
  NOR U48180 ( .A(n35255), .B(n42041), .Z(n35259) );
  IV U48181 ( .A(n35256), .Z(n35257) );
  NOR U48182 ( .A(n35258), .B(n35257), .Z(n42034) );
  NOR U48183 ( .A(n35259), .B(n42034), .Z(n38664) );
  IV U48184 ( .A(n35260), .Z(n35261) );
  NOR U48185 ( .A(n35262), .B(n35261), .Z(n38677) );
  IV U48186 ( .A(n35263), .Z(n35264) );
  NOR U48187 ( .A(n35265), .B(n35264), .Z(n38674) );
  NOR U48188 ( .A(n38677), .B(n38674), .Z(n36818) );
  IV U48189 ( .A(n35266), .Z(n35268) );
  NOR U48190 ( .A(n35268), .B(n35267), .Z(n40116) );
  IV U48191 ( .A(n35269), .Z(n35270) );
  NOR U48192 ( .A(n35271), .B(n35270), .Z(n38679) );
  IV U48193 ( .A(n35272), .Z(n35273) );
  NOR U48194 ( .A(n35274), .B(n35273), .Z(n38683) );
  IV U48195 ( .A(n35275), .Z(n35277) );
  NOR U48196 ( .A(n35277), .B(n35276), .Z(n40099) );
  NOR U48197 ( .A(n38683), .B(n40099), .Z(n36810) );
  IV U48198 ( .A(n35278), .Z(n35282) );
  NOR U48199 ( .A(n35280), .B(n35279), .Z(n35281) );
  IV U48200 ( .A(n35281), .Z(n36798) );
  NOR U48201 ( .A(n35282), .B(n36798), .Z(n38687) );
  IV U48202 ( .A(n35283), .Z(n35290) );
  NOR U48203 ( .A(n35285), .B(n35284), .Z(n35286) );
  IV U48204 ( .A(n35286), .Z(n35287) );
  NOR U48205 ( .A(n35288), .B(n35287), .Z(n35289) );
  IV U48206 ( .A(n35289), .Z(n35292) );
  NOR U48207 ( .A(n35290), .B(n35292), .Z(n38695) );
  NOR U48208 ( .A(n38687), .B(n38695), .Z(n36795) );
  IV U48209 ( .A(n35291), .Z(n35293) );
  NOR U48210 ( .A(n35293), .B(n35292), .Z(n38692) );
  IV U48211 ( .A(n36790), .Z(n43532) );
  IV U48212 ( .A(n35294), .Z(n35301) );
  NOR U48213 ( .A(n35296), .B(n35295), .Z(n35297) );
  IV U48214 ( .A(n35297), .Z(n35298) );
  NOR U48215 ( .A(n35299), .B(n35298), .Z(n35300) );
  IV U48216 ( .A(n35300), .Z(n36776) );
  NOR U48217 ( .A(n35301), .B(n36776), .Z(n35302) );
  IV U48218 ( .A(n35302), .Z(n40082) );
  IV U48219 ( .A(n35303), .Z(n35305) );
  NOR U48220 ( .A(n35305), .B(n35304), .Z(n35306) );
  IV U48221 ( .A(n35306), .Z(n36778) );
  IV U48222 ( .A(n35307), .Z(n35308) );
  NOR U48223 ( .A(n35309), .B(n35308), .Z(n35310) );
  IV U48224 ( .A(n35310), .Z(n36767) );
  IV U48225 ( .A(n35311), .Z(n35312) );
  NOR U48226 ( .A(n35315), .B(n35312), .Z(n40070) );
  IV U48227 ( .A(n35313), .Z(n35314) );
  NOR U48228 ( .A(n35315), .B(n35314), .Z(n35316) );
  IV U48229 ( .A(n35316), .Z(n38715) );
  IV U48230 ( .A(n35317), .Z(n35324) );
  IV U48231 ( .A(n35318), .Z(n35326) );
  NOR U48232 ( .A(n35319), .B(n35326), .Z(n35320) );
  IV U48233 ( .A(n35320), .Z(n35321) );
  NOR U48234 ( .A(n35322), .B(n35321), .Z(n35323) );
  IV U48235 ( .A(n35323), .Z(n36738) );
  NOR U48236 ( .A(n35324), .B(n36738), .Z(n38733) );
  IV U48237 ( .A(n35325), .Z(n35329) );
  NOR U48238 ( .A(n35327), .B(n35326), .Z(n35328) );
  IV U48239 ( .A(n35328), .Z(n35331) );
  NOR U48240 ( .A(n35329), .B(n35331), .Z(n40061) );
  IV U48241 ( .A(n35330), .Z(n35332) );
  NOR U48242 ( .A(n35332), .B(n35331), .Z(n40058) );
  NOR U48243 ( .A(n38739), .B(n40058), .Z(n36735) );
  NOR U48244 ( .A(n35334), .B(n35333), .Z(n38736) );
  IV U48245 ( .A(n35335), .Z(n35342) );
  NOR U48246 ( .A(n35337), .B(n35336), .Z(n35338) );
  IV U48247 ( .A(n35338), .Z(n35339) );
  NOR U48248 ( .A(n35340), .B(n35339), .Z(n35341) );
  IV U48249 ( .A(n35341), .Z(n35344) );
  NOR U48250 ( .A(n35342), .B(n35344), .Z(n38744) );
  IV U48251 ( .A(n35343), .Z(n35345) );
  NOR U48252 ( .A(n35345), .B(n35344), .Z(n38753) );
  IV U48253 ( .A(n35346), .Z(n35348) );
  IV U48254 ( .A(n35347), .Z(n36731) );
  NOR U48255 ( .A(n35348), .B(n36731), .Z(n38750) );
  IV U48256 ( .A(n35349), .Z(n35351) );
  XOR U48257 ( .A(n35356), .B(n35354), .Z(n35350) );
  NOR U48258 ( .A(n35351), .B(n35350), .Z(n40050) );
  IV U48259 ( .A(n35352), .Z(n35353) );
  NOR U48260 ( .A(n35356), .B(n35353), .Z(n40047) );
  IV U48261 ( .A(n35354), .Z(n35355) );
  NOR U48262 ( .A(n35356), .B(n35355), .Z(n38758) );
  NOR U48263 ( .A(n35358), .B(n35357), .Z(n38767) );
  IV U48264 ( .A(n35359), .Z(n35361) );
  NOR U48265 ( .A(n35361), .B(n35360), .Z(n36685) );
  IV U48266 ( .A(n35362), .Z(n35364) );
  NOR U48267 ( .A(n35364), .B(n35363), .Z(n36683) );
  IV U48268 ( .A(n36683), .Z(n36678) );
  IV U48269 ( .A(n35365), .Z(n35366) );
  NOR U48270 ( .A(n36675), .B(n35366), .Z(n36672) );
  IV U48271 ( .A(n36672), .Z(n36652) );
  NOR U48272 ( .A(n35367), .B(n38784), .Z(n36651) );
  IV U48273 ( .A(n35368), .Z(n35369) );
  NOR U48274 ( .A(n35369), .B(n35376), .Z(n39983) );
  IV U48275 ( .A(n35370), .Z(n35374) );
  NOR U48276 ( .A(n35372), .B(n35371), .Z(n35373) );
  IV U48277 ( .A(n35373), .Z(n36640) );
  NOR U48278 ( .A(n35374), .B(n36640), .Z(n39976) );
  IV U48279 ( .A(n35375), .Z(n35377) );
  NOR U48280 ( .A(n35377), .B(n35376), .Z(n39981) );
  NOR U48281 ( .A(n39976), .B(n39981), .Z(n36642) );
  IV U48282 ( .A(n35378), .Z(n35379) );
  NOR U48283 ( .A(n36626), .B(n35379), .Z(n38787) );
  IV U48284 ( .A(n35380), .Z(n35381) );
  NOR U48285 ( .A(n35382), .B(n35381), .Z(n38799) );
  NOR U48286 ( .A(n38801), .B(n38799), .Z(n36624) );
  IV U48287 ( .A(n35383), .Z(n35384) );
  NOR U48288 ( .A(n35386), .B(n35384), .Z(n39968) );
  IV U48289 ( .A(n35385), .Z(n35387) );
  NOR U48290 ( .A(n35387), .B(n35386), .Z(n35388) );
  IV U48291 ( .A(n35388), .Z(n39967) );
  IV U48292 ( .A(n35389), .Z(n35391) );
  NOR U48293 ( .A(n35391), .B(n35390), .Z(n42202) );
  NOR U48294 ( .A(n42207), .B(n42202), .Z(n38809) );
  IV U48295 ( .A(n35392), .Z(n35393) );
  NOR U48296 ( .A(n35393), .B(n35395), .Z(n39946) );
  IV U48297 ( .A(n35394), .Z(n35396) );
  NOR U48298 ( .A(n35396), .B(n35395), .Z(n42224) );
  IV U48299 ( .A(n35397), .Z(n35399) );
  IV U48300 ( .A(n35398), .Z(n42228) );
  NOR U48301 ( .A(n35399), .B(n42228), .Z(n46748) );
  NOR U48302 ( .A(n42224), .B(n46748), .Z(n39944) );
  IV U48303 ( .A(n35400), .Z(n35401) );
  NOR U48304 ( .A(n36606), .B(n35401), .Z(n39938) );
  IV U48305 ( .A(n35402), .Z(n35404) );
  NOR U48306 ( .A(n35404), .B(n35403), .Z(n38829) );
  IV U48307 ( .A(n35405), .Z(n35407) );
  NOR U48308 ( .A(n35407), .B(n35406), .Z(n39935) );
  NOR U48309 ( .A(n38829), .B(n39935), .Z(n36602) );
  IV U48310 ( .A(n35408), .Z(n35409) );
  NOR U48311 ( .A(n35410), .B(n35409), .Z(n35411) );
  IV U48312 ( .A(n35411), .Z(n38835) );
  IV U48313 ( .A(n35412), .Z(n35413) );
  NOR U48314 ( .A(n35413), .B(n35415), .Z(n38842) );
  IV U48315 ( .A(n35414), .Z(n35418) );
  NOR U48316 ( .A(n35416), .B(n35415), .Z(n35417) );
  IV U48317 ( .A(n35417), .Z(n35420) );
  NOR U48318 ( .A(n35418), .B(n35420), .Z(n38847) );
  NOR U48319 ( .A(n38842), .B(n38847), .Z(n36575) );
  IV U48320 ( .A(n35419), .Z(n35421) );
  NOR U48321 ( .A(n35421), .B(n35420), .Z(n38850) );
  NOR U48322 ( .A(n35422), .B(n38850), .Z(n36574) );
  IV U48323 ( .A(n35423), .Z(n38854) );
  NOR U48324 ( .A(n38854), .B(n35424), .Z(n35428) );
  IV U48325 ( .A(n35425), .Z(n35427) );
  NOR U48326 ( .A(n35427), .B(n35426), .Z(n39905) );
  NOR U48327 ( .A(n35428), .B(n39905), .Z(n36573) );
  IV U48328 ( .A(n35429), .Z(n35430) );
  NOR U48329 ( .A(n35431), .B(n35430), .Z(n36569) );
  IV U48330 ( .A(n35432), .Z(n35433) );
  NOR U48331 ( .A(n35436), .B(n35433), .Z(n39884) );
  IV U48332 ( .A(n35434), .Z(n35435) );
  NOR U48333 ( .A(n35436), .B(n35435), .Z(n39896) );
  NOR U48334 ( .A(n39884), .B(n39896), .Z(n36568) );
  IV U48335 ( .A(n35437), .Z(n35440) );
  IV U48336 ( .A(n35438), .Z(n35439) );
  NOR U48337 ( .A(n35440), .B(n35439), .Z(n39880) );
  IV U48338 ( .A(n35441), .Z(n35442) );
  NOR U48339 ( .A(n35442), .B(n50105), .Z(n39887) );
  IV U48340 ( .A(n35443), .Z(n35444) );
  NOR U48341 ( .A(n35444), .B(n35447), .Z(n39867) );
  IV U48342 ( .A(n35445), .Z(n35446) );
  NOR U48343 ( .A(n35447), .B(n35446), .Z(n38860) );
  IV U48344 ( .A(n35448), .Z(n35450) );
  NOR U48345 ( .A(n35450), .B(n35449), .Z(n35451) );
  IV U48346 ( .A(n35451), .Z(n36554) );
  NOR U48347 ( .A(n35452), .B(n35461), .Z(n35453) );
  IV U48348 ( .A(n35453), .Z(n35454) );
  NOR U48349 ( .A(n35455), .B(n35454), .Z(n39852) );
  IV U48350 ( .A(n35456), .Z(n35458) );
  NOR U48351 ( .A(n35458), .B(n35457), .Z(n43281) );
  IV U48352 ( .A(n35459), .Z(n35460) );
  NOR U48353 ( .A(n35461), .B(n35460), .Z(n43301) );
  NOR U48354 ( .A(n43281), .B(n43301), .Z(n38866) );
  IV U48355 ( .A(n35462), .Z(n35464) );
  NOR U48356 ( .A(n35464), .B(n35463), .Z(n39838) );
  IV U48357 ( .A(n35465), .Z(n35467) );
  NOR U48358 ( .A(n35467), .B(n35466), .Z(n39847) );
  NOR U48359 ( .A(n39838), .B(n39847), .Z(n36546) );
  IV U48360 ( .A(n35468), .Z(n35469) );
  NOR U48361 ( .A(n35470), .B(n35469), .Z(n35471) );
  IV U48362 ( .A(n35471), .Z(n39842) );
  IV U48363 ( .A(n35472), .Z(n36541) );
  IV U48364 ( .A(n35473), .Z(n35474) );
  NOR U48365 ( .A(n36535), .B(n35474), .Z(n36530) );
  NOR U48366 ( .A(n35476), .B(n35475), .Z(n39820) );
  IV U48367 ( .A(n35477), .Z(n35479) );
  IV U48368 ( .A(n35478), .Z(n36524) );
  NOR U48369 ( .A(n35479), .B(n36524), .Z(n39823) );
  NOR U48370 ( .A(n39820), .B(n39823), .Z(n36518) );
  IV U48371 ( .A(n35480), .Z(n42302) );
  NOR U48372 ( .A(n35481), .B(n42302), .Z(n38874) );
  IV U48373 ( .A(n35482), .Z(n35483) );
  NOR U48374 ( .A(n35488), .B(n35483), .Z(n38882) );
  IV U48375 ( .A(n35484), .Z(n35485) );
  NOR U48376 ( .A(n35486), .B(n35485), .Z(n42305) );
  IV U48377 ( .A(n35487), .Z(n35489) );
  NOR U48378 ( .A(n35489), .B(n35488), .Z(n43263) );
  NOR U48379 ( .A(n42305), .B(n43263), .Z(n38881) );
  IV U48380 ( .A(n35490), .Z(n35491) );
  NOR U48381 ( .A(n35491), .B(n39797), .Z(n39806) );
  IV U48382 ( .A(n35492), .Z(n35494) );
  NOR U48383 ( .A(n35494), .B(n35493), .Z(n38911) );
  IV U48384 ( .A(n35495), .Z(n35497) );
  NOR U48385 ( .A(n35497), .B(n35496), .Z(n38906) );
  NOR U48386 ( .A(n38911), .B(n38906), .Z(n36497) );
  IV U48387 ( .A(n35498), .Z(n35502) );
  NOR U48388 ( .A(n35506), .B(n35509), .Z(n35499) );
  IV U48389 ( .A(n35499), .Z(n35514) );
  NOR U48390 ( .A(n35500), .B(n35514), .Z(n35501) );
  IV U48391 ( .A(n35501), .Z(n35504) );
  NOR U48392 ( .A(n35502), .B(n35504), .Z(n38908) );
  IV U48393 ( .A(n35503), .Z(n35505) );
  NOR U48394 ( .A(n35505), .B(n35504), .Z(n38917) );
  NOR U48395 ( .A(n35507), .B(n35506), .Z(n35508) );
  IV U48396 ( .A(n35508), .Z(n35510) );
  NOR U48397 ( .A(n35510), .B(n35509), .Z(n35511) );
  IV U48398 ( .A(n35511), .Z(n35512) );
  NOR U48399 ( .A(n35513), .B(n35512), .Z(n38914) );
  IV U48400 ( .A(n35513), .Z(n35518) );
  NOR U48401 ( .A(n35515), .B(n35514), .Z(n35516) );
  IV U48402 ( .A(n35516), .Z(n35517) );
  NOR U48403 ( .A(n35518), .B(n35517), .Z(n35519) );
  IV U48404 ( .A(n35519), .Z(n38923) );
  IV U48405 ( .A(n35520), .Z(n35525) );
  IV U48406 ( .A(n35521), .Z(n35522) );
  NOR U48407 ( .A(n35525), .B(n35522), .Z(n42329) );
  IV U48408 ( .A(n35523), .Z(n35524) );
  NOR U48409 ( .A(n35525), .B(n35524), .Z(n43220) );
  NOR U48410 ( .A(n42329), .B(n43220), .Z(n38920) );
  IV U48411 ( .A(n35526), .Z(n35527) );
  NOR U48412 ( .A(n35532), .B(n35527), .Z(n38927) );
  IV U48413 ( .A(n35528), .Z(n35530) );
  NOR U48414 ( .A(n35530), .B(n35529), .Z(n38933) );
  IV U48415 ( .A(n35531), .Z(n35533) );
  NOR U48416 ( .A(n35533), .B(n35532), .Z(n38925) );
  NOR U48417 ( .A(n38933), .B(n38925), .Z(n36495) );
  IV U48418 ( .A(n35534), .Z(n35535) );
  NOR U48419 ( .A(n35535), .B(n36492), .Z(n43203) );
  IV U48420 ( .A(n35536), .Z(n35539) );
  NOR U48421 ( .A(n35537), .B(n35547), .Z(n35538) );
  IV U48422 ( .A(n35538), .Z(n35541) );
  NOR U48423 ( .A(n35539), .B(n35541), .Z(n43201) );
  NOR U48424 ( .A(n43203), .B(n43201), .Z(n39772) );
  IV U48425 ( .A(n35540), .Z(n35542) );
  NOR U48426 ( .A(n35542), .B(n35541), .Z(n38940) );
  IV U48427 ( .A(n35543), .Z(n35545) );
  NOR U48428 ( .A(n35545), .B(n35544), .Z(n35546) );
  IV U48429 ( .A(n35546), .Z(n35548) );
  NOR U48430 ( .A(n35548), .B(n35547), .Z(n39764) );
  IV U48431 ( .A(n35549), .Z(n35551) );
  IV U48432 ( .A(n35550), .Z(n36485) );
  NOR U48433 ( .A(n35551), .B(n36485), .Z(n39761) );
  IV U48434 ( .A(n36482), .Z(n36474) );
  IV U48435 ( .A(n35552), .Z(n35559) );
  IV U48436 ( .A(n35553), .Z(n36464) );
  NOR U48437 ( .A(n35554), .B(n36464), .Z(n35555) );
  IV U48438 ( .A(n35555), .Z(n35556) );
  NOR U48439 ( .A(n35557), .B(n35556), .Z(n35558) );
  IV U48440 ( .A(n35558), .Z(n36468) );
  NOR U48441 ( .A(n35559), .B(n36468), .Z(n39754) );
  NOR U48442 ( .A(n35561), .B(n35560), .Z(n39751) );
  IV U48443 ( .A(n35562), .Z(n35563) );
  NOR U48444 ( .A(n36462), .B(n35563), .Z(n39747) );
  IV U48445 ( .A(n35564), .Z(n35565) );
  NOR U48446 ( .A(n35565), .B(n35567), .Z(n38960) );
  IV U48447 ( .A(n35566), .Z(n35568) );
  NOR U48448 ( .A(n35568), .B(n35567), .Z(n38955) );
  NOR U48449 ( .A(n38960), .B(n38955), .Z(n36452) );
  IV U48450 ( .A(n35569), .Z(n35573) );
  NOR U48451 ( .A(n35571), .B(n35570), .Z(n35572) );
  IV U48452 ( .A(n35572), .Z(n35578) );
  NOR U48453 ( .A(n35573), .B(n35578), .Z(n38957) );
  IV U48454 ( .A(n35574), .Z(n35576) );
  NOR U48455 ( .A(n35576), .B(n35575), .Z(n46539) );
  IV U48456 ( .A(n35577), .Z(n35579) );
  NOR U48457 ( .A(n35579), .B(n35578), .Z(n45695) );
  NOR U48458 ( .A(n46539), .B(n45695), .Z(n39728) );
  IV U48459 ( .A(n35580), .Z(n35582) );
  IV U48460 ( .A(n35581), .Z(n35587) );
  NOR U48461 ( .A(n35582), .B(n35587), .Z(n35583) );
  IV U48462 ( .A(n35583), .Z(n38967) );
  IV U48463 ( .A(n35584), .Z(n35585) );
  NOR U48464 ( .A(n35585), .B(n35587), .Z(n38964) );
  IV U48465 ( .A(n35586), .Z(n35588) );
  NOR U48466 ( .A(n35588), .B(n35587), .Z(n38972) );
  IV U48467 ( .A(n35589), .Z(n35590) );
  NOR U48468 ( .A(n35590), .B(n35597), .Z(n39696) );
  NOR U48469 ( .A(n35592), .B(n35591), .Z(n35593) );
  IV U48470 ( .A(n35593), .Z(n46503) );
  NOR U48471 ( .A(n35594), .B(n46503), .Z(n42384) );
  IV U48472 ( .A(n35595), .Z(n35596) );
  NOR U48473 ( .A(n35597), .B(n35596), .Z(n42378) );
  NOR U48474 ( .A(n42384), .B(n42378), .Z(n38977) );
  IV U48475 ( .A(n35598), .Z(n49192) );
  NOR U48476 ( .A(n35599), .B(n49192), .Z(n35600) );
  IV U48477 ( .A(n35600), .Z(n36400) );
  IV U48478 ( .A(n35601), .Z(n35602) );
  NOR U48479 ( .A(n35603), .B(n35602), .Z(n35604) );
  IV U48480 ( .A(n35604), .Z(n36388) );
  IV U48481 ( .A(n35605), .Z(n35606) );
  NOR U48482 ( .A(n35607), .B(n35606), .Z(n38989) );
  IV U48483 ( .A(n35608), .Z(n35609) );
  NOR U48484 ( .A(n35609), .B(n36375), .Z(n38991) );
  NOR U48485 ( .A(n38989), .B(n38991), .Z(n36381) );
  IV U48486 ( .A(n35610), .Z(n35611) );
  NOR U48487 ( .A(n35612), .B(n35611), .Z(n39665) );
  IV U48488 ( .A(n35613), .Z(n35620) );
  NOR U48489 ( .A(n35615), .B(n35614), .Z(n35616) );
  IV U48490 ( .A(n35616), .Z(n35617) );
  NOR U48491 ( .A(n35618), .B(n35617), .Z(n35619) );
  IV U48492 ( .A(n35619), .Z(n35625) );
  NOR U48493 ( .A(n35620), .B(n35625), .Z(n35621) );
  IV U48494 ( .A(n35621), .Z(n39664) );
  IV U48495 ( .A(n35622), .Z(n35623) );
  NOR U48496 ( .A(n35623), .B(n35628), .Z(n42409) );
  IV U48497 ( .A(n35624), .Z(n35626) );
  NOR U48498 ( .A(n35626), .B(n35625), .Z(n43085) );
  NOR U48499 ( .A(n42409), .B(n43085), .Z(n39659) );
  IV U48500 ( .A(n35627), .Z(n35629) );
  NOR U48501 ( .A(n35629), .B(n35628), .Z(n39656) );
  IV U48502 ( .A(n35630), .Z(n35632) );
  NOR U48503 ( .A(n35632), .B(n35631), .Z(n38998) );
  IV U48504 ( .A(n35633), .Z(n35635) );
  NOR U48505 ( .A(n35635), .B(n35634), .Z(n39652) );
  NOR U48506 ( .A(n38998), .B(n39652), .Z(n36372) );
  IV U48507 ( .A(n35636), .Z(n35637) );
  NOR U48508 ( .A(n35637), .B(n36362), .Z(n35638) );
  IV U48509 ( .A(n35638), .Z(n38997) );
  IV U48510 ( .A(n35639), .Z(n35644) );
  IV U48511 ( .A(n35640), .Z(n35641) );
  NOR U48512 ( .A(n35644), .B(n35641), .Z(n39638) );
  IV U48513 ( .A(n35642), .Z(n35643) );
  NOR U48514 ( .A(n35644), .B(n35643), .Z(n39641) );
  IV U48515 ( .A(n35645), .Z(n35646) );
  NOR U48516 ( .A(n35646), .B(n35648), .Z(n39020) );
  NOR U48517 ( .A(n39641), .B(n39020), .Z(n36334) );
  IV U48518 ( .A(n35647), .Z(n35652) );
  NOR U48519 ( .A(n35649), .B(n35648), .Z(n35650) );
  IV U48520 ( .A(n35650), .Z(n35651) );
  NOR U48521 ( .A(n35652), .B(n35651), .Z(n39017) );
  IV U48522 ( .A(n35653), .Z(n35659) );
  XOR U48523 ( .A(n35655), .B(n35654), .Z(n35656) );
  NOR U48524 ( .A(n35656), .B(n35661), .Z(n35657) );
  IV U48525 ( .A(n35657), .Z(n35658) );
  NOR U48526 ( .A(n35659), .B(n35658), .Z(n39634) );
  IV U48527 ( .A(n35660), .Z(n35662) );
  NOR U48528 ( .A(n35662), .B(n35661), .Z(n39631) );
  IV U48529 ( .A(n35663), .Z(n35664) );
  NOR U48530 ( .A(n35665), .B(n35664), .Z(n42443) );
  IV U48531 ( .A(n35666), .Z(n35667) );
  NOR U48532 ( .A(n35668), .B(n35667), .Z(n43062) );
  NOR U48533 ( .A(n42443), .B(n43062), .Z(n39625) );
  IV U48534 ( .A(n35669), .Z(n35671) );
  NOR U48535 ( .A(n35671), .B(n35670), .Z(n35672) );
  IV U48536 ( .A(n35672), .Z(n36318) );
  IV U48537 ( .A(n35673), .Z(n35679) );
  IV U48538 ( .A(n35674), .Z(n35675) );
  NOR U48539 ( .A(n35679), .B(n35675), .Z(n35676) );
  IV U48540 ( .A(n35676), .Z(n39612) );
  IV U48541 ( .A(n35677), .Z(n35678) );
  NOR U48542 ( .A(n35679), .B(n35678), .Z(n39608) );
  IV U48543 ( .A(n35680), .Z(n35682) );
  NOR U48544 ( .A(n35682), .B(n35681), .Z(n39605) );
  IV U48545 ( .A(n35683), .Z(n35684) );
  NOR U48546 ( .A(n35684), .B(n36304), .Z(n36300) );
  IV U48547 ( .A(n36300), .Z(n36294) );
  IV U48548 ( .A(n35685), .Z(n36297) );
  IV U48549 ( .A(n35686), .Z(n35687) );
  NOR U48550 ( .A(n36297), .B(n35687), .Z(n39029) );
  IV U48551 ( .A(n35688), .Z(n35690) );
  NOR U48552 ( .A(n35690), .B(n35689), .Z(n39036) );
  IV U48553 ( .A(n35691), .Z(n35692) );
  NOR U48554 ( .A(n35692), .B(n35698), .Z(n39033) );
  IV U48555 ( .A(n35693), .Z(n35694) );
  NOR U48556 ( .A(n35695), .B(n35694), .Z(n42476) );
  IV U48557 ( .A(n35696), .Z(n35697) );
  NOR U48558 ( .A(n35698), .B(n35697), .Z(n42471) );
  NOR U48559 ( .A(n42476), .B(n42471), .Z(n39040) );
  IV U48560 ( .A(n35699), .Z(n35701) );
  IV U48561 ( .A(n35700), .Z(n35703) );
  NOR U48562 ( .A(n35701), .B(n35703), .Z(n39585) );
  IV U48563 ( .A(n35702), .Z(n35704) );
  NOR U48564 ( .A(n35704), .B(n35703), .Z(n39043) );
  NOR U48565 ( .A(n39585), .B(n39043), .Z(n35705) );
  IV U48566 ( .A(n35705), .Z(n35709) );
  IV U48567 ( .A(n35706), .Z(n35707) );
  NOR U48568 ( .A(n35708), .B(n35707), .Z(n39041) );
  NOR U48569 ( .A(n35709), .B(n39041), .Z(n36292) );
  IV U48570 ( .A(n35710), .Z(n35711) );
  NOR U48571 ( .A(n35711), .B(n35713), .Z(n39589) );
  IV U48572 ( .A(n35712), .Z(n35714) );
  NOR U48573 ( .A(n35714), .B(n35713), .Z(n39045) );
  IV U48574 ( .A(n35715), .Z(n35717) );
  IV U48575 ( .A(n35716), .Z(n35719) );
  NOR U48576 ( .A(n35717), .B(n35719), .Z(n39050) );
  IV U48577 ( .A(n35718), .Z(n35720) );
  NOR U48578 ( .A(n35720), .B(n35719), .Z(n39580) );
  NOR U48579 ( .A(n39572), .B(n39580), .Z(n36282) );
  IV U48580 ( .A(n35721), .Z(n35722) );
  NOR U48581 ( .A(n35722), .B(n36272), .Z(n36269) );
  IV U48582 ( .A(n36269), .Z(n36260) );
  IV U48583 ( .A(n35723), .Z(n35725) );
  NOR U48584 ( .A(n35725), .B(n35724), .Z(n35726) );
  IV U48585 ( .A(n35726), .Z(n39060) );
  IV U48586 ( .A(n35727), .Z(n35728) );
  NOR U48587 ( .A(n35728), .B(n35730), .Z(n39062) );
  IV U48588 ( .A(n35729), .Z(n35731) );
  NOR U48589 ( .A(n35731), .B(n35730), .Z(n39554) );
  NOR U48590 ( .A(n39062), .B(n39554), .Z(n36251) );
  IV U48591 ( .A(n35732), .Z(n35736) );
  NOR U48592 ( .A(n35734), .B(n35733), .Z(n35735) );
  IV U48593 ( .A(n35735), .Z(n36247) );
  NOR U48594 ( .A(n35736), .B(n36247), .Z(n39066) );
  IV U48595 ( .A(n35737), .Z(n35738) );
  NOR U48596 ( .A(n35738), .B(n35744), .Z(n39074) );
  IV U48597 ( .A(n35739), .Z(n35740) );
  NOR U48598 ( .A(n35741), .B(n35740), .Z(n39080) );
  IV U48599 ( .A(n35742), .Z(n35743) );
  NOR U48600 ( .A(n35744), .B(n35743), .Z(n39072) );
  NOR U48601 ( .A(n39080), .B(n39072), .Z(n36241) );
  IV U48602 ( .A(n35745), .Z(n35747) );
  IV U48603 ( .A(n35746), .Z(n35749) );
  NOR U48604 ( .A(n35747), .B(n35749), .Z(n39077) );
  IV U48605 ( .A(n35748), .Z(n35750) );
  NOR U48606 ( .A(n35750), .B(n35749), .Z(n39546) );
  IV U48607 ( .A(n35751), .Z(n35756) );
  IV U48608 ( .A(n35752), .Z(n35759) );
  NOR U48609 ( .A(n35753), .B(n35759), .Z(n35754) );
  IV U48610 ( .A(n35754), .Z(n35755) );
  NOR U48611 ( .A(n35756), .B(n35755), .Z(n39543) );
  IV U48612 ( .A(n35757), .Z(n35758) );
  NOR U48613 ( .A(n35766), .B(n35758), .Z(n39084) );
  NOR U48614 ( .A(n35760), .B(n35759), .Z(n35761) );
  IV U48615 ( .A(n35761), .Z(n35762) );
  NOR U48616 ( .A(n35763), .B(n35762), .Z(n39086) );
  NOR U48617 ( .A(n39084), .B(n39086), .Z(n36240) );
  IV U48618 ( .A(n35764), .Z(n35765) );
  NOR U48619 ( .A(n35766), .B(n35765), .Z(n39089) );
  IV U48620 ( .A(n35767), .Z(n35772) );
  IV U48621 ( .A(n35768), .Z(n35769) );
  NOR U48622 ( .A(n35772), .B(n35769), .Z(n39539) );
  NOR U48623 ( .A(n39089), .B(n39539), .Z(n36239) );
  IV U48624 ( .A(n35770), .Z(n35771) );
  NOR U48625 ( .A(n35772), .B(n35771), .Z(n39534) );
  NOR U48626 ( .A(n35774), .B(n35773), .Z(n39094) );
  NOR U48627 ( .A(n39096), .B(n39094), .Z(n36227) );
  IV U48628 ( .A(n35775), .Z(n36214) );
  IV U48629 ( .A(n35776), .Z(n35777) );
  NOR U48630 ( .A(n36214), .B(n35777), .Z(n39513) );
  NOR U48631 ( .A(n35778), .B(n39106), .Z(n35779) );
  NOR U48632 ( .A(n39513), .B(n35779), .Z(n36220) );
  IV U48633 ( .A(n35780), .Z(n35781) );
  NOR U48634 ( .A(n35781), .B(n35786), .Z(n39506) );
  IV U48635 ( .A(n35782), .Z(n35783) );
  NOR U48636 ( .A(n35784), .B(n35783), .Z(n39114) );
  IV U48637 ( .A(n35785), .Z(n35787) );
  NOR U48638 ( .A(n35787), .B(n35786), .Z(n39509) );
  NOR U48639 ( .A(n39114), .B(n39509), .Z(n36210) );
  IV U48640 ( .A(n35788), .Z(n35790) );
  IV U48641 ( .A(n35789), .Z(n36207) );
  NOR U48642 ( .A(n35790), .B(n36207), .Z(n39111) );
  IV U48643 ( .A(n35791), .Z(n35792) );
  NOR U48644 ( .A(n35792), .B(n36207), .Z(n39501) );
  IV U48645 ( .A(n35793), .Z(n35794) );
  NOR U48646 ( .A(n35795), .B(n35794), .Z(n39495) );
  IV U48647 ( .A(n35796), .Z(n35797) );
  NOR U48648 ( .A(n35798), .B(n35797), .Z(n42952) );
  IV U48649 ( .A(n35799), .Z(n35800) );
  NOR U48650 ( .A(n35801), .B(n35800), .Z(n42961) );
  NOR U48651 ( .A(n42952), .B(n42961), .Z(n39494) );
  IV U48652 ( .A(n35802), .Z(n35803) );
  NOR U48653 ( .A(n35804), .B(n35803), .Z(n39490) );
  IV U48654 ( .A(n35805), .Z(n35808) );
  NOR U48655 ( .A(n35806), .B(n36199), .Z(n35807) );
  IV U48656 ( .A(n35807), .Z(n36201) );
  NOR U48657 ( .A(n35808), .B(n36201), .Z(n39487) );
  IV U48658 ( .A(n35809), .Z(n35810) );
  NOR U48659 ( .A(n35811), .B(n35810), .Z(n42944) );
  IV U48660 ( .A(n35812), .Z(n35813) );
  NOR U48661 ( .A(n35813), .B(n35815), .Z(n42586) );
  NOR U48662 ( .A(n42944), .B(n42586), .Z(n39481) );
  IV U48663 ( .A(n35814), .Z(n35816) );
  NOR U48664 ( .A(n35816), .B(n35815), .Z(n35817) );
  IV U48665 ( .A(n35817), .Z(n39478) );
  IV U48666 ( .A(n35818), .Z(n35819) );
  NOR U48667 ( .A(n35820), .B(n35819), .Z(n39468) );
  IV U48668 ( .A(n35821), .Z(n35822) );
  NOR U48669 ( .A(n35823), .B(n35822), .Z(n39474) );
  NOR U48670 ( .A(n39468), .B(n39474), .Z(n36196) );
  IV U48671 ( .A(n35824), .Z(n35825) );
  NOR U48672 ( .A(n35827), .B(n35825), .Z(n39463) );
  IV U48673 ( .A(n35826), .Z(n35828) );
  NOR U48674 ( .A(n35828), .B(n35827), .Z(n39465) );
  NOR U48675 ( .A(n39463), .B(n39465), .Z(n36194) );
  IV U48676 ( .A(n35829), .Z(n35831) );
  NOR U48677 ( .A(n35831), .B(n35830), .Z(n39456) );
  IV U48678 ( .A(n35832), .Z(n35834) );
  NOR U48679 ( .A(n35834), .B(n35833), .Z(n39460) );
  NOR U48680 ( .A(n39456), .B(n39460), .Z(n36193) );
  IV U48681 ( .A(n35835), .Z(n35837) );
  NOR U48682 ( .A(n35837), .B(n35836), .Z(n36191) );
  IV U48683 ( .A(n36191), .Z(n36182) );
  IV U48684 ( .A(n35838), .Z(n35839) );
  NOR U48685 ( .A(n35840), .B(n35839), .Z(n35841) );
  IV U48686 ( .A(n35841), .Z(n39452) );
  IV U48687 ( .A(n35842), .Z(n35844) );
  NOR U48688 ( .A(n35844), .B(n35843), .Z(n39439) );
  IV U48689 ( .A(n35845), .Z(n35849) );
  IV U48690 ( .A(n35846), .Z(n35848) );
  NOR U48691 ( .A(n35848), .B(n35847), .Z(n35854) );
  XOR U48692 ( .A(n35854), .B(n35856), .Z(n35850) );
  NOR U48693 ( .A(n35849), .B(n35850), .Z(n39435) );
  NOR U48694 ( .A(n35851), .B(n35850), .Z(n39432) );
  IV U48695 ( .A(n35852), .Z(n39120) );
  NOR U48696 ( .A(n35853), .B(n39120), .Z(n35857) );
  IV U48697 ( .A(n35854), .Z(n35855) );
  NOR U48698 ( .A(n35856), .B(n35855), .Z(n39429) );
  NOR U48699 ( .A(n35857), .B(n39429), .Z(n36167) );
  IV U48700 ( .A(n35858), .Z(n39134) );
  NOR U48701 ( .A(n39134), .B(n35859), .Z(n39127) );
  IV U48702 ( .A(n35860), .Z(n35861) );
  NOR U48703 ( .A(n35862), .B(n35861), .Z(n39140) );
  IV U48704 ( .A(n35863), .Z(n35864) );
  NOR U48705 ( .A(n35865), .B(n35864), .Z(n42628) );
  IV U48706 ( .A(n35866), .Z(n35867) );
  NOR U48707 ( .A(n35867), .B(n36145), .Z(n42623) );
  NOR U48708 ( .A(n42628), .B(n42623), .Z(n39412) );
  IV U48709 ( .A(n35868), .Z(n36112) );
  NOR U48710 ( .A(n35870), .B(n35869), .Z(n39396) );
  IV U48711 ( .A(n35871), .Z(n35878) );
  NOR U48712 ( .A(n35873), .B(n35872), .Z(n35874) );
  IV U48713 ( .A(n35874), .Z(n35875) );
  NOR U48714 ( .A(n35876), .B(n35875), .Z(n35877) );
  IV U48715 ( .A(n35877), .Z(n35880) );
  NOR U48716 ( .A(n35878), .B(n35880), .Z(n39400) );
  IV U48717 ( .A(n35879), .Z(n35881) );
  NOR U48718 ( .A(n35881), .B(n35880), .Z(n39392) );
  IV U48719 ( .A(n35882), .Z(n35883) );
  NOR U48720 ( .A(n35884), .B(n35883), .Z(n39157) );
  IV U48721 ( .A(n35885), .Z(n35887) );
  NOR U48722 ( .A(n35887), .B(n35886), .Z(n39160) );
  NOR U48723 ( .A(n39157), .B(n39160), .Z(n36098) );
  IV U48724 ( .A(n35888), .Z(n35889) );
  NOR U48725 ( .A(n35889), .B(n35894), .Z(n39373) );
  IV U48726 ( .A(n35890), .Z(n35891) );
  NOR U48727 ( .A(n35892), .B(n35891), .Z(n39164) );
  NOR U48728 ( .A(n39373), .B(n39164), .Z(n36091) );
  IV U48729 ( .A(n35893), .Z(n35895) );
  NOR U48730 ( .A(n35895), .B(n35894), .Z(n39370) );
  IV U48731 ( .A(n35896), .Z(n35897) );
  NOR U48732 ( .A(n35898), .B(n35897), .Z(n39376) );
  IV U48733 ( .A(n35899), .Z(n35901) );
  IV U48734 ( .A(n35900), .Z(n39172) );
  NOR U48735 ( .A(n35901), .B(n39172), .Z(n39169) );
  NOR U48736 ( .A(n39376), .B(n39169), .Z(n36090) );
  NOR U48737 ( .A(n35902), .B(n39172), .Z(n35905) );
  IV U48738 ( .A(n35903), .Z(n35904) );
  NOR U48739 ( .A(n36088), .B(n35904), .Z(n39182) );
  NOR U48740 ( .A(n35905), .B(n39182), .Z(n36089) );
  IV U48741 ( .A(n35906), .Z(n35907) );
  NOR U48742 ( .A(n36088), .B(n35907), .Z(n39179) );
  IV U48743 ( .A(n35908), .Z(n35909) );
  NOR U48744 ( .A(n35909), .B(n36075), .Z(n39190) );
  IV U48745 ( .A(n35910), .Z(n35912) );
  NOR U48746 ( .A(n35912), .B(n35911), .Z(n39197) );
  IV U48747 ( .A(n35913), .Z(n35914) );
  NOR U48748 ( .A(n35914), .B(n36075), .Z(n39195) );
  NOR U48749 ( .A(n39197), .B(n39195), .Z(n36073) );
  NOR U48750 ( .A(n35916), .B(n35915), .Z(n39323) );
  IV U48751 ( .A(n35917), .Z(n36063) );
  IV U48752 ( .A(n36062), .Z(n35918) );
  NOR U48753 ( .A(n36063), .B(n35918), .Z(n39330) );
  NOR U48754 ( .A(n39323), .B(n39330), .Z(n36060) );
  NOR U48755 ( .A(n35920), .B(n35919), .Z(n39202) );
  IV U48756 ( .A(n35921), .Z(n35922) );
  NOR U48757 ( .A(n35922), .B(n36059), .Z(n36052) );
  IV U48758 ( .A(n35923), .Z(n35925) );
  NOR U48759 ( .A(n35925), .B(n35924), .Z(n36049) );
  IV U48760 ( .A(n36049), .Z(n36044) );
  IV U48761 ( .A(n35926), .Z(n35927) );
  NOR U48762 ( .A(n36023), .B(n35927), .Z(n39209) );
  IV U48763 ( .A(n35928), .Z(n35929) );
  NOR U48764 ( .A(n35929), .B(n36023), .Z(n39293) );
  IV U48765 ( .A(n35930), .Z(n35932) );
  NOR U48766 ( .A(n35932), .B(n35931), .Z(n35933) );
  IV U48767 ( .A(n35933), .Z(n36016) );
  IV U48768 ( .A(n35934), .Z(n35935) );
  NOR U48769 ( .A(n35938), .B(n35935), .Z(n39215) );
  IV U48770 ( .A(n35936), .Z(n35937) );
  NOR U48771 ( .A(n35938), .B(n35937), .Z(n42730) );
  IV U48772 ( .A(n35939), .Z(n35941) );
  IV U48773 ( .A(n35940), .Z(n35943) );
  NOR U48774 ( .A(n35941), .B(n35943), .Z(n42683) );
  NOR U48775 ( .A(n42730), .B(n42683), .Z(n39220) );
  IV U48776 ( .A(n39220), .Z(n36007) );
  IV U48777 ( .A(n35942), .Z(n35944) );
  NOR U48778 ( .A(n35944), .B(n35943), .Z(n39217) );
  IV U48779 ( .A(n35945), .Z(n35947) );
  IV U48780 ( .A(n35946), .Z(n35951) );
  NOR U48781 ( .A(n35947), .B(n35951), .Z(n39222) );
  NOR U48782 ( .A(n35949), .B(n35948), .Z(n39262) );
  IV U48783 ( .A(n35950), .Z(n35952) );
  NOR U48784 ( .A(n35952), .B(n35951), .Z(n39225) );
  NOR U48785 ( .A(n39262), .B(n39225), .Z(n36000) );
  IV U48786 ( .A(n39261), .Z(n39254) );
  IV U48787 ( .A(n35953), .Z(n35958) );
  IV U48788 ( .A(n35954), .Z(n35955) );
  NOR U48789 ( .A(n35958), .B(n35955), .Z(n39247) );
  IV U48790 ( .A(n35956), .Z(n35957) );
  NOR U48791 ( .A(n35958), .B(n35957), .Z(n39228) );
  IV U48792 ( .A(n35959), .Z(n35961) );
  NOR U48793 ( .A(n35961), .B(n35960), .Z(n39234) );
  NOR U48794 ( .A(n35963), .B(n35962), .Z(n39243) );
  NOR U48795 ( .A(n39234), .B(n39243), .Z(n35991) );
  IV U48796 ( .A(n35964), .Z(n35965) );
  NOR U48797 ( .A(n35965), .B(n35989), .Z(n35966) );
  IV U48798 ( .A(n35966), .Z(n39233) );
  IV U48799 ( .A(n35967), .Z(n35968) );
  NOR U48800 ( .A(n35969), .B(n35968), .Z(n35983) );
  IV U48801 ( .A(n35983), .Z(n35978) );
  IV U48802 ( .A(n35970), .Z(n35972) );
  NOR U48803 ( .A(n35972), .B(n35971), .Z(n35976) );
  NOR U48804 ( .A(n35974), .B(n35973), .Z(n35975) );
  NOR U48805 ( .A(n35976), .B(n35975), .Z(n35982) );
  IV U48806 ( .A(n35982), .Z(n35977) );
  NOR U48807 ( .A(n35978), .B(n35977), .Z(n39239) );
  IV U48808 ( .A(n35979), .Z(n35980) );
  NOR U48809 ( .A(n35981), .B(n35980), .Z(n35986) );
  NOR U48810 ( .A(n35983), .B(n35982), .Z(n35984) );
  IV U48811 ( .A(n35984), .Z(n35985) );
  NOR U48812 ( .A(n35986), .B(n35985), .Z(n39237) );
  NOR U48813 ( .A(n39239), .B(n39237), .Z(n35990) );
  IV U48814 ( .A(n35987), .Z(n35988) );
  NOR U48815 ( .A(n35989), .B(n35988), .Z(n39235) );
  XOR U48816 ( .A(n35990), .B(n39235), .Z(n39231) );
  XOR U48817 ( .A(n39233), .B(n39231), .Z(n39244) );
  XOR U48818 ( .A(n35991), .B(n39244), .Z(n35992) );
  IV U48819 ( .A(n35992), .Z(n39230) );
  XOR U48820 ( .A(n39228), .B(n39230), .Z(n39248) );
  XOR U48821 ( .A(n39247), .B(n39248), .Z(n39258) );
  IV U48822 ( .A(n35993), .Z(n35994) );
  NOR U48823 ( .A(n35995), .B(n35994), .Z(n39250) );
  IV U48824 ( .A(n35996), .Z(n35998) );
  NOR U48825 ( .A(n35998), .B(n35997), .Z(n39257) );
  NOR U48826 ( .A(n39250), .B(n39257), .Z(n35999) );
  XOR U48827 ( .A(n39258), .B(n35999), .Z(n39260) );
  XOR U48828 ( .A(n39254), .B(n39260), .Z(n39227) );
  XOR U48829 ( .A(n36000), .B(n39227), .Z(n36001) );
  IV U48830 ( .A(n36001), .Z(n39224) );
  XOR U48831 ( .A(n39222), .B(n39224), .Z(n39273) );
  IV U48832 ( .A(n36002), .Z(n36003) );
  NOR U48833 ( .A(n36006), .B(n36003), .Z(n39271) );
  XOR U48834 ( .A(n39273), .B(n39271), .Z(n39276) );
  IV U48835 ( .A(n36004), .Z(n36005) );
  NOR U48836 ( .A(n36006), .B(n36005), .Z(n39274) );
  XOR U48837 ( .A(n39276), .B(n39274), .Z(n39218) );
  XOR U48838 ( .A(n39217), .B(n39218), .Z(n42686) );
  XOR U48839 ( .A(n36007), .B(n42686), .Z(n39280) );
  XOR U48840 ( .A(n39215), .B(n39280), .Z(n36014) );
  NOR U48841 ( .A(n36016), .B(n36014), .Z(n42680) );
  IV U48842 ( .A(n36008), .Z(n36010) );
  NOR U48843 ( .A(n36010), .B(n36009), .Z(n36011) );
  IV U48844 ( .A(n36011), .Z(n39214) );
  IV U48845 ( .A(n36012), .Z(n39281) );
  NOR U48846 ( .A(n36013), .B(n39281), .Z(n36015) );
  XOR U48847 ( .A(n36015), .B(n36014), .Z(n39213) );
  XOR U48848 ( .A(n39214), .B(n39213), .Z(n36019) );
  IV U48849 ( .A(n39213), .Z(n36017) );
  NOR U48850 ( .A(n36017), .B(n36016), .Z(n36018) );
  NOR U48851 ( .A(n36019), .B(n36018), .Z(n36020) );
  NOR U48852 ( .A(n42680), .B(n36020), .Z(n36021) );
  IV U48853 ( .A(n36021), .Z(n39294) );
  XOR U48854 ( .A(n39293), .B(n39294), .Z(n39210) );
  XOR U48855 ( .A(n39209), .B(n39210), .Z(n39291) );
  IV U48856 ( .A(n36022), .Z(n36024) );
  NOR U48857 ( .A(n36024), .B(n36023), .Z(n39289) );
  XOR U48858 ( .A(n39291), .B(n39289), .Z(n39303) );
  IV U48859 ( .A(n36025), .Z(n36026) );
  NOR U48860 ( .A(n36027), .B(n36026), .Z(n39205) );
  IV U48861 ( .A(n36028), .Z(n36031) );
  IV U48862 ( .A(n36029), .Z(n36030) );
  NOR U48863 ( .A(n36031), .B(n36030), .Z(n39301) );
  NOR U48864 ( .A(n39205), .B(n39301), .Z(n36032) );
  XOR U48865 ( .A(n39303), .B(n36032), .Z(n39207) );
  IV U48866 ( .A(n36033), .Z(n36034) );
  NOR U48867 ( .A(n36035), .B(n36034), .Z(n39307) );
  IV U48868 ( .A(n36036), .Z(n36038) );
  NOR U48869 ( .A(n36038), .B(n36037), .Z(n42754) );
  IV U48870 ( .A(n36039), .Z(n36041) );
  NOR U48871 ( .A(n36041), .B(n36040), .Z(n42671) );
  NOR U48872 ( .A(n42754), .B(n42671), .Z(n39208) );
  IV U48873 ( .A(n39208), .Z(n36042) );
  NOR U48874 ( .A(n39307), .B(n36042), .Z(n36043) );
  XOR U48875 ( .A(n39207), .B(n36043), .Z(n39310) );
  NOR U48876 ( .A(n36044), .B(n39310), .Z(n42758) );
  IV U48877 ( .A(n36045), .Z(n36046) );
  NOR U48878 ( .A(n36047), .B(n36046), .Z(n39309) );
  XOR U48879 ( .A(n39309), .B(n39310), .Z(n36053) );
  IV U48880 ( .A(n36053), .Z(n36048) );
  NOR U48881 ( .A(n36049), .B(n36048), .Z(n36050) );
  NOR U48882 ( .A(n42758), .B(n36050), .Z(n36051) );
  NOR U48883 ( .A(n36052), .B(n36051), .Z(n36055) );
  IV U48884 ( .A(n36052), .Z(n36054) );
  NOR U48885 ( .A(n36054), .B(n36053), .Z(n42766) );
  NOR U48886 ( .A(n36055), .B(n42766), .Z(n36056) );
  IV U48887 ( .A(n36056), .Z(n39315) );
  IV U48888 ( .A(n36057), .Z(n36058) );
  NOR U48889 ( .A(n36059), .B(n36058), .Z(n39314) );
  XOR U48890 ( .A(n39315), .B(n39314), .Z(n39203) );
  XOR U48891 ( .A(n39202), .B(n39203), .Z(n39319) );
  XOR U48892 ( .A(n39318), .B(n39319), .Z(n39332) );
  XOR U48893 ( .A(n36060), .B(n39332), .Z(n39327) );
  IV U48894 ( .A(n36061), .Z(n36065) );
  XOR U48895 ( .A(n36063), .B(n36062), .Z(n36064) );
  NOR U48896 ( .A(n36065), .B(n36064), .Z(n36066) );
  IV U48897 ( .A(n36066), .Z(n39328) );
  XOR U48898 ( .A(n39327), .B(n39328), .Z(n39344) );
  IV U48899 ( .A(n36067), .Z(n36068) );
  NOR U48900 ( .A(n36069), .B(n36068), .Z(n39347) );
  IV U48901 ( .A(n36070), .Z(n36072) );
  NOR U48902 ( .A(n36072), .B(n36071), .Z(n39341) );
  NOR U48903 ( .A(n39347), .B(n39341), .Z(n39201) );
  XOR U48904 ( .A(n39344), .B(n39201), .Z(n39194) );
  XOR U48905 ( .A(n36073), .B(n39194), .Z(n39192) );
  XOR U48906 ( .A(n39190), .B(n39192), .Z(n39360) );
  IV U48907 ( .A(n36074), .Z(n36076) );
  NOR U48908 ( .A(n36076), .B(n36075), .Z(n39358) );
  XOR U48909 ( .A(n39360), .B(n39358), .Z(n39354) );
  IV U48910 ( .A(n39354), .Z(n36085) );
  IV U48911 ( .A(n36080), .Z(n36078) );
  IV U48912 ( .A(n36077), .Z(n36081) );
  NOR U48913 ( .A(n36078), .B(n36081), .Z(n39353) );
  IV U48914 ( .A(n36079), .Z(n36083) );
  XOR U48915 ( .A(n36081), .B(n36080), .Z(n36082) );
  NOR U48916 ( .A(n36083), .B(n36082), .Z(n39188) );
  NOR U48917 ( .A(n39353), .B(n39188), .Z(n36084) );
  XOR U48918 ( .A(n36085), .B(n36084), .Z(n39187) );
  IV U48919 ( .A(n36086), .Z(n36087) );
  NOR U48920 ( .A(n36088), .B(n36087), .Z(n39185) );
  XOR U48921 ( .A(n39187), .B(n39185), .Z(n39180) );
  XOR U48922 ( .A(n39179), .B(n39180), .Z(n39184) );
  XOR U48923 ( .A(n36089), .B(n39184), .Z(n39168) );
  XOR U48924 ( .A(n36090), .B(n39168), .Z(n39371) );
  XOR U48925 ( .A(n39370), .B(n39371), .Z(n39374) );
  XOR U48926 ( .A(n36091), .B(n39374), .Z(n42646) );
  IV U48927 ( .A(n36092), .Z(n36093) );
  NOR U48928 ( .A(n36093), .B(n36095), .Z(n39166) );
  IV U48929 ( .A(n36094), .Z(n36096) );
  NOR U48930 ( .A(n36096), .B(n36095), .Z(n39159) );
  NOR U48931 ( .A(n39166), .B(n39159), .Z(n36097) );
  XOR U48932 ( .A(n42646), .B(n36097), .Z(n39162) );
  XOR U48933 ( .A(n36098), .B(n39162), .Z(n39155) );
  IV U48934 ( .A(n36099), .Z(n36100) );
  NOR U48935 ( .A(n36100), .B(n36106), .Z(n39154) );
  IV U48936 ( .A(n36101), .Z(n36103) );
  NOR U48937 ( .A(n36103), .B(n36102), .Z(n39385) );
  NOR U48938 ( .A(n39154), .B(n39385), .Z(n36104) );
  XOR U48939 ( .A(n39155), .B(n36104), .Z(n39391) );
  IV U48940 ( .A(n36105), .Z(n36107) );
  NOR U48941 ( .A(n36107), .B(n36106), .Z(n39389) );
  XOR U48942 ( .A(n39391), .B(n39389), .Z(n39393) );
  XOR U48943 ( .A(n39392), .B(n39393), .Z(n39401) );
  XOR U48944 ( .A(n39400), .B(n39401), .Z(n39151) );
  XOR U48945 ( .A(n39150), .B(n39151), .Z(n39397) );
  XOR U48946 ( .A(n39396), .B(n39397), .Z(n36121) );
  NOR U48947 ( .A(n36117), .B(n36121), .Z(n36108) );
  IV U48948 ( .A(n36108), .Z(n36109) );
  NOR U48949 ( .A(n36110), .B(n36109), .Z(n36111) );
  IV U48950 ( .A(n36111), .Z(n36114) );
  NOR U48951 ( .A(n36112), .B(n36114), .Z(n42856) );
  IV U48952 ( .A(n36113), .Z(n36115) );
  NOR U48953 ( .A(n36115), .B(n36114), .Z(n42848) );
  IV U48954 ( .A(n36116), .Z(n36118) );
  NOR U48955 ( .A(n36118), .B(n36117), .Z(n36124) );
  IV U48956 ( .A(n36119), .Z(n39144) );
  NOR U48957 ( .A(n36120), .B(n39144), .Z(n36122) );
  XOR U48958 ( .A(n36122), .B(n36121), .Z(n36134) );
  IV U48959 ( .A(n36134), .Z(n36123) );
  NOR U48960 ( .A(n36124), .B(n36123), .Z(n36125) );
  NOR U48961 ( .A(n42848), .B(n36125), .Z(n36126) );
  IV U48962 ( .A(n36126), .Z(n36127) );
  NOR U48963 ( .A(n42856), .B(n36127), .Z(n39409) );
  IV U48964 ( .A(n36128), .Z(n36130) );
  NOR U48965 ( .A(n36130), .B(n36129), .Z(n36140) );
  IV U48966 ( .A(n36140), .Z(n39411) );
  NOR U48967 ( .A(n39409), .B(n39411), .Z(n36142) );
  IV U48968 ( .A(n36131), .Z(n36132) );
  NOR U48969 ( .A(n36133), .B(n36132), .Z(n36136) );
  IV U48970 ( .A(n36136), .Z(n36135) );
  NOR U48971 ( .A(n36135), .B(n36134), .Z(n42852) );
  NOR U48972 ( .A(n39409), .B(n36136), .Z(n36137) );
  NOR U48973 ( .A(n42852), .B(n36137), .Z(n36138) );
  IV U48974 ( .A(n36138), .Z(n36139) );
  NOR U48975 ( .A(n36140), .B(n36139), .Z(n36141) );
  NOR U48976 ( .A(n36142), .B(n36141), .Z(n42624) );
  XOR U48977 ( .A(n39412), .B(n42624), .Z(n39137) );
  IV U48978 ( .A(n36143), .Z(n36144) );
  NOR U48979 ( .A(n36145), .B(n36144), .Z(n36146) );
  IV U48980 ( .A(n36146), .Z(n39138) );
  XOR U48981 ( .A(n39137), .B(n39138), .Z(n39141) );
  XOR U48982 ( .A(n39140), .B(n39141), .Z(n36156) );
  IV U48983 ( .A(n36156), .Z(n36154) );
  IV U48984 ( .A(n36147), .Z(n36148) );
  NOR U48985 ( .A(n36149), .B(n36148), .Z(n36158) );
  NOR U48986 ( .A(n36151), .B(n36150), .Z(n36155) );
  NOR U48987 ( .A(n36158), .B(n36155), .Z(n36152) );
  IV U48988 ( .A(n36152), .Z(n36153) );
  NOR U48989 ( .A(n36154), .B(n36153), .Z(n36161) );
  IV U48990 ( .A(n36155), .Z(n36157) );
  NOR U48991 ( .A(n36157), .B(n36156), .Z(n42621) );
  IV U48992 ( .A(n36158), .Z(n36159) );
  NOR U48993 ( .A(n36159), .B(n39141), .Z(n42866) );
  NOR U48994 ( .A(n42621), .B(n42866), .Z(n36160) );
  IV U48995 ( .A(n36160), .Z(n39418) );
  NOR U48996 ( .A(n36161), .B(n39418), .Z(n39133) );
  NOR U48997 ( .A(n36163), .B(n36162), .Z(n36164) );
  NOR U48998 ( .A(n39415), .B(n36164), .Z(n36165) );
  XOR U48999 ( .A(n39133), .B(n36165), .Z(n39129) );
  XOR U49000 ( .A(n39127), .B(n39129), .Z(n39123) );
  XOR U49001 ( .A(n36166), .B(n39123), .Z(n39430) );
  XOR U49002 ( .A(n36167), .B(n39430), .Z(n36168) );
  IV U49003 ( .A(n36168), .Z(n39434) );
  XOR U49004 ( .A(n39432), .B(n39434), .Z(n39436) );
  XOR U49005 ( .A(n39435), .B(n39436), .Z(n39440) );
  XOR U49006 ( .A(n39439), .B(n39440), .Z(n39447) );
  IV U49007 ( .A(n39447), .Z(n36177) );
  IV U49008 ( .A(n36169), .Z(n36170) );
  NOR U49009 ( .A(n36171), .B(n36170), .Z(n39442) );
  NOR U49010 ( .A(n36172), .B(n36179), .Z(n36173) );
  IV U49011 ( .A(n36173), .Z(n36174) );
  NOR U49012 ( .A(n36175), .B(n36174), .Z(n39445) );
  NOR U49013 ( .A(n39442), .B(n39445), .Z(n36176) );
  XOR U49014 ( .A(n36177), .B(n36176), .Z(n39450) );
  IV U49015 ( .A(n36178), .Z(n36180) );
  NOR U49016 ( .A(n36180), .B(n36179), .Z(n39448) );
  XOR U49017 ( .A(n39450), .B(n39448), .Z(n39451) );
  XOR U49018 ( .A(n39452), .B(n39451), .Z(n36187) );
  IV U49019 ( .A(n36187), .Z(n36181) );
  NOR U49020 ( .A(n36182), .B(n36181), .Z(n42604) );
  IV U49021 ( .A(n36183), .Z(n36184) );
  NOR U49022 ( .A(n36185), .B(n36184), .Z(n36188) );
  IV U49023 ( .A(n36188), .Z(n36186) );
  NOR U49024 ( .A(n36186), .B(n39451), .Z(n42607) );
  NOR U49025 ( .A(n36188), .B(n36187), .Z(n36189) );
  NOR U49026 ( .A(n42607), .B(n36189), .Z(n36190) );
  NOR U49027 ( .A(n36191), .B(n36190), .Z(n36192) );
  NOR U49028 ( .A(n42604), .B(n36192), .Z(n39457) );
  XOR U49029 ( .A(n36193), .B(n39457), .Z(n39467) );
  XOR U49030 ( .A(n36194), .B(n39467), .Z(n39117) );
  XOR U49031 ( .A(n36195), .B(n39117), .Z(n39476) );
  XOR U49032 ( .A(n36196), .B(n39476), .Z(n39477) );
  XOR U49033 ( .A(n39478), .B(n39477), .Z(n42588) );
  XOR U49034 ( .A(n39481), .B(n42588), .Z(n39482) );
  IV U49035 ( .A(n36197), .Z(n36198) );
  NOR U49036 ( .A(n36199), .B(n36198), .Z(n42947) );
  IV U49037 ( .A(n36200), .Z(n36202) );
  NOR U49038 ( .A(n36202), .B(n36201), .Z(n42579) );
  NOR U49039 ( .A(n42947), .B(n42579), .Z(n39483) );
  XOR U49040 ( .A(n39482), .B(n39483), .Z(n39489) );
  XOR U49041 ( .A(n39487), .B(n39489), .Z(n39492) );
  XOR U49042 ( .A(n39490), .B(n39492), .Z(n42954) );
  XOR U49043 ( .A(n39494), .B(n42954), .Z(n36203) );
  IV U49044 ( .A(n36203), .Z(n39496) );
  XOR U49045 ( .A(n39495), .B(n39496), .Z(n42570) );
  IV U49046 ( .A(n42570), .Z(n36209) );
  NOR U49047 ( .A(n36205), .B(n36204), .Z(n42574) );
  IV U49048 ( .A(n36206), .Z(n36208) );
  NOR U49049 ( .A(n36208), .B(n36207), .Z(n42569) );
  NOR U49050 ( .A(n42574), .B(n42569), .Z(n39500) );
  XOR U49051 ( .A(n36209), .B(n39500), .Z(n39503) );
  XOR U49052 ( .A(n39501), .B(n39503), .Z(n39112) );
  XOR U49053 ( .A(n39111), .B(n39112), .Z(n39510) );
  XOR U49054 ( .A(n36210), .B(n39510), .Z(n36211) );
  IV U49055 ( .A(n36211), .Z(n39508) );
  XOR U49056 ( .A(n39506), .B(n39508), .Z(n39517) );
  IV U49057 ( .A(n39517), .Z(n36219) );
  IV U49058 ( .A(n36212), .Z(n36213) );
  NOR U49059 ( .A(n36214), .B(n36213), .Z(n39516) );
  IV U49060 ( .A(n36215), .Z(n36217) );
  NOR U49061 ( .A(n36217), .B(n36216), .Z(n39109) );
  NOR U49062 ( .A(n39516), .B(n39109), .Z(n36218) );
  XOR U49063 ( .A(n36219), .B(n36218), .Z(n39515) );
  XOR U49064 ( .A(n36220), .B(n39515), .Z(n39100) );
  IV U49065 ( .A(n36221), .Z(n36223) );
  NOR U49066 ( .A(n36223), .B(n36222), .Z(n39102) );
  NOR U49067 ( .A(n36225), .B(n36224), .Z(n39099) );
  NOR U49068 ( .A(n39102), .B(n39099), .Z(n36226) );
  XOR U49069 ( .A(n39100), .B(n36226), .Z(n39097) );
  XOR U49070 ( .A(n36227), .B(n39097), .Z(n39092) );
  IV U49071 ( .A(n36228), .Z(n36230) );
  IV U49072 ( .A(n36229), .Z(n36231) );
  NOR U49073 ( .A(n36230), .B(n36231), .Z(n39528) );
  NOR U49074 ( .A(n36232), .B(n36231), .Z(n39526) );
  NOR U49075 ( .A(n39091), .B(n39526), .Z(n36233) );
  IV U49076 ( .A(n36233), .Z(n36234) );
  NOR U49077 ( .A(n39528), .B(n36234), .Z(n36235) );
  XOR U49078 ( .A(n39092), .B(n36235), .Z(n39533) );
  IV U49079 ( .A(n36236), .Z(n36238) );
  NOR U49080 ( .A(n36238), .B(n36237), .Z(n39531) );
  XOR U49081 ( .A(n39533), .B(n39531), .Z(n39535) );
  XOR U49082 ( .A(n39534), .B(n39535), .Z(n39541) );
  XOR U49083 ( .A(n36239), .B(n39541), .Z(n39083) );
  XOR U49084 ( .A(n36240), .B(n39083), .Z(n39544) );
  XOR U49085 ( .A(n39543), .B(n39544), .Z(n39547) );
  XOR U49086 ( .A(n39546), .B(n39547), .Z(n39078) );
  XOR U49087 ( .A(n39077), .B(n39078), .Z(n39081) );
  XOR U49088 ( .A(n36241), .B(n39081), .Z(n36242) );
  IV U49089 ( .A(n36242), .Z(n39075) );
  XOR U49090 ( .A(n39074), .B(n39075), .Z(n39070) );
  IV U49091 ( .A(n39070), .Z(n36250) );
  IV U49092 ( .A(n36243), .Z(n36245) );
  NOR U49093 ( .A(n36245), .B(n36244), .Z(n39069) );
  IV U49094 ( .A(n36246), .Z(n36248) );
  NOR U49095 ( .A(n36248), .B(n36247), .Z(n39064) );
  NOR U49096 ( .A(n39069), .B(n39064), .Z(n36249) );
  XOR U49097 ( .A(n36250), .B(n36249), .Z(n39067) );
  XOR U49098 ( .A(n39066), .B(n39067), .Z(n39556) );
  XOR U49099 ( .A(n36251), .B(n39556), .Z(n39558) );
  IV U49100 ( .A(n36252), .Z(n36253) );
  NOR U49101 ( .A(n36254), .B(n36253), .Z(n39562) );
  IV U49102 ( .A(n36255), .Z(n36257) );
  NOR U49103 ( .A(n36257), .B(n36256), .Z(n39557) );
  NOR U49104 ( .A(n39562), .B(n39557), .Z(n36258) );
  XOR U49105 ( .A(n39558), .B(n36258), .Z(n39061) );
  XOR U49106 ( .A(n39060), .B(n39061), .Z(n36265) );
  IV U49107 ( .A(n36265), .Z(n36259) );
  NOR U49108 ( .A(n36260), .B(n36259), .Z(n42501) );
  IV U49109 ( .A(n36261), .Z(n36262) );
  NOR U49110 ( .A(n36263), .B(n36262), .Z(n36266) );
  IV U49111 ( .A(n36266), .Z(n36264) );
  NOR U49112 ( .A(n39061), .B(n36264), .Z(n42507) );
  NOR U49113 ( .A(n36266), .B(n36265), .Z(n36267) );
  NOR U49114 ( .A(n42507), .B(n36267), .Z(n36268) );
  NOR U49115 ( .A(n36269), .B(n36268), .Z(n36270) );
  NOR U49116 ( .A(n42501), .B(n36270), .Z(n39566) );
  IV U49117 ( .A(n36271), .Z(n36273) );
  NOR U49118 ( .A(n36273), .B(n36272), .Z(n36274) );
  IV U49119 ( .A(n36274), .Z(n39567) );
  XOR U49120 ( .A(n39566), .B(n39567), .Z(n42498) );
  IV U49121 ( .A(n42498), .Z(n36281) );
  IV U49122 ( .A(n36275), .Z(n36276) );
  NOR U49123 ( .A(n36277), .B(n36276), .Z(n42496) );
  IV U49124 ( .A(n36278), .Z(n36279) );
  NOR U49125 ( .A(n36280), .B(n36279), .Z(n43023) );
  NOR U49126 ( .A(n42496), .B(n43023), .Z(n39570) );
  XOR U49127 ( .A(n36281), .B(n39570), .Z(n39057) );
  XOR U49128 ( .A(n39056), .B(n39057), .Z(n39582) );
  XOR U49129 ( .A(n36282), .B(n39582), .Z(n36283) );
  IV U49130 ( .A(n36283), .Z(n39052) );
  XOR U49131 ( .A(n39050), .B(n39052), .Z(n39054) );
  IV U49132 ( .A(n39054), .Z(n36291) );
  IV U49133 ( .A(n36284), .Z(n36285) );
  NOR U49134 ( .A(n36286), .B(n36285), .Z(n39053) );
  IV U49135 ( .A(n36287), .Z(n36288) );
  NOR U49136 ( .A(n36289), .B(n36288), .Z(n39048) );
  NOR U49137 ( .A(n39053), .B(n39048), .Z(n36290) );
  XOR U49138 ( .A(n36291), .B(n36290), .Z(n39047) );
  XOR U49139 ( .A(n39045), .B(n39047), .Z(n39590) );
  XOR U49140 ( .A(n39589), .B(n39590), .Z(n39586) );
  XOR U49141 ( .A(n36292), .B(n39586), .Z(n39039) );
  XOR U49142 ( .A(n39040), .B(n39039), .Z(n39035) );
  XOR U49143 ( .A(n39033), .B(n39035), .Z(n39037) );
  XOR U49144 ( .A(n39036), .B(n39037), .Z(n39031) );
  XOR U49145 ( .A(n39029), .B(n39031), .Z(n36293) );
  NOR U49146 ( .A(n36294), .B(n36293), .Z(n45782) );
  IV U49147 ( .A(n36295), .Z(n36296) );
  NOR U49148 ( .A(n36297), .B(n36296), .Z(n39027) );
  NOR U49149 ( .A(n39029), .B(n39027), .Z(n36298) );
  XOR U49150 ( .A(n39031), .B(n36298), .Z(n36299) );
  NOR U49151 ( .A(n36300), .B(n36299), .Z(n36301) );
  NOR U49152 ( .A(n45782), .B(n36301), .Z(n36302) );
  IV U49153 ( .A(n36302), .Z(n39026) );
  IV U49154 ( .A(n36303), .Z(n36305) );
  NOR U49155 ( .A(n36305), .B(n36304), .Z(n39024) );
  XOR U49156 ( .A(n39026), .B(n39024), .Z(n39607) );
  XOR U49157 ( .A(n39605), .B(n39607), .Z(n42451) );
  XOR U49158 ( .A(n39608), .B(n42451), .Z(n39611) );
  XOR U49159 ( .A(n39612), .B(n39611), .Z(n36309) );
  IV U49160 ( .A(n36309), .Z(n36306) );
  NOR U49161 ( .A(n36318), .B(n36306), .Z(n43051) );
  NOR U49162 ( .A(n36307), .B(n42454), .Z(n36310) );
  IV U49163 ( .A(n36310), .Z(n36308) );
  NOR U49164 ( .A(n36308), .B(n42451), .Z(n39613) );
  NOR U49165 ( .A(n36310), .B(n36309), .Z(n36311) );
  NOR U49166 ( .A(n39613), .B(n36311), .Z(n36312) );
  IV U49167 ( .A(n36312), .Z(n39023) );
  IV U49168 ( .A(n36313), .Z(n36317) );
  NOR U49169 ( .A(n36329), .B(n36314), .Z(n36315) );
  IV U49170 ( .A(n36315), .Z(n36316) );
  NOR U49171 ( .A(n36317), .B(n36316), .Z(n36319) );
  IV U49172 ( .A(n36319), .Z(n39022) );
  XOR U49173 ( .A(n39023), .B(n39022), .Z(n36321) );
  NOR U49174 ( .A(n36319), .B(n36318), .Z(n36320) );
  NOR U49175 ( .A(n36321), .B(n36320), .Z(n36322) );
  NOR U49176 ( .A(n43051), .B(n36322), .Z(n36323) );
  IV U49177 ( .A(n36323), .Z(n39619) );
  IV U49178 ( .A(n36324), .Z(n36325) );
  NOR U49179 ( .A(n36326), .B(n36325), .Z(n36327) );
  IV U49180 ( .A(n36327), .Z(n36328) );
  NOR U49181 ( .A(n36329), .B(n36328), .Z(n39617) );
  XOR U49182 ( .A(n39619), .B(n39617), .Z(n39627) );
  IV U49183 ( .A(n36330), .Z(n36332) );
  NOR U49184 ( .A(n36332), .B(n36331), .Z(n39626) );
  NOR U49185 ( .A(n39620), .B(n39626), .Z(n36333) );
  XOR U49186 ( .A(n39627), .B(n36333), .Z(n39624) );
  XOR U49187 ( .A(n39625), .B(n39624), .Z(n39632) );
  XOR U49188 ( .A(n39631), .B(n39632), .Z(n39636) );
  XOR U49189 ( .A(n39634), .B(n39636), .Z(n39019) );
  XOR U49190 ( .A(n39017), .B(n39019), .Z(n39643) );
  XOR U49191 ( .A(n36334), .B(n39643), .Z(n36335) );
  IV U49192 ( .A(n36335), .Z(n39640) );
  XOR U49193 ( .A(n39638), .B(n39640), .Z(n39016) );
  IV U49194 ( .A(n36336), .Z(n36342) );
  NOR U49195 ( .A(n36337), .B(n36347), .Z(n36338) );
  IV U49196 ( .A(n36338), .Z(n36339) );
  NOR U49197 ( .A(n36340), .B(n36339), .Z(n36341) );
  IV U49198 ( .A(n36341), .Z(n36344) );
  NOR U49199 ( .A(n36342), .B(n36344), .Z(n39014) );
  XOR U49200 ( .A(n39016), .B(n39014), .Z(n39011) );
  IV U49201 ( .A(n36343), .Z(n36345) );
  NOR U49202 ( .A(n36345), .B(n36344), .Z(n39009) );
  XOR U49203 ( .A(n39011), .B(n39009), .Z(n39013) );
  IV U49204 ( .A(n36346), .Z(n36348) );
  NOR U49205 ( .A(n36348), .B(n36347), .Z(n36349) );
  IV U49206 ( .A(n36349), .Z(n39012) );
  XOR U49207 ( .A(n39013), .B(n39012), .Z(n39003) );
  IV U49208 ( .A(n36350), .Z(n36352) );
  NOR U49209 ( .A(n36352), .B(n36351), .Z(n39007) );
  IV U49210 ( .A(n36353), .Z(n36354) );
  NOR U49211 ( .A(n36354), .B(n36366), .Z(n39004) );
  NOR U49212 ( .A(n39007), .B(n39004), .Z(n36355) );
  XOR U49213 ( .A(n39003), .B(n36355), .Z(n39648) );
  IV U49214 ( .A(n36356), .Z(n36357) );
  NOR U49215 ( .A(n36358), .B(n36357), .Z(n36359) );
  IV U49216 ( .A(n36359), .Z(n36367) );
  NOR U49217 ( .A(n39648), .B(n36367), .Z(n42424) );
  IV U49218 ( .A(n36360), .Z(n36361) );
  NOR U49219 ( .A(n36362), .B(n36361), .Z(n36363) );
  IV U49220 ( .A(n36363), .Z(n39002) );
  IV U49221 ( .A(n36364), .Z(n36365) );
  NOR U49222 ( .A(n36366), .B(n36365), .Z(n39646) );
  XOR U49223 ( .A(n39646), .B(n39648), .Z(n39001) );
  XOR U49224 ( .A(n39002), .B(n39001), .Z(n36370) );
  IV U49225 ( .A(n39001), .Z(n36368) );
  NOR U49226 ( .A(n36368), .B(n36367), .Z(n36369) );
  NOR U49227 ( .A(n36370), .B(n36369), .Z(n36371) );
  NOR U49228 ( .A(n42424), .B(n36371), .Z(n38996) );
  XOR U49229 ( .A(n38997), .B(n38996), .Z(n39653) );
  XOR U49230 ( .A(n36372), .B(n39653), .Z(n36373) );
  IV U49231 ( .A(n36373), .Z(n39658) );
  XOR U49232 ( .A(n39656), .B(n39658), .Z(n42410) );
  XOR U49233 ( .A(n39659), .B(n42410), .Z(n39662) );
  XOR U49234 ( .A(n39664), .B(n39662), .Z(n39666) );
  XOR U49235 ( .A(n39665), .B(n39666), .Z(n39672) );
  IV U49236 ( .A(n36374), .Z(n36376) );
  NOR U49237 ( .A(n36376), .B(n36375), .Z(n38994) );
  IV U49238 ( .A(n36377), .Z(n36379) );
  NOR U49239 ( .A(n36379), .B(n36378), .Z(n39670) );
  NOR U49240 ( .A(n38994), .B(n39670), .Z(n36380) );
  XOR U49241 ( .A(n39672), .B(n36380), .Z(n38988) );
  XOR U49242 ( .A(n36381), .B(n38988), .Z(n38986) );
  NOR U49243 ( .A(n36388), .B(n38986), .Z(n42394) );
  IV U49244 ( .A(n36382), .Z(n36383) );
  NOR U49245 ( .A(n36383), .B(n49190), .Z(n36384) );
  IV U49246 ( .A(n36384), .Z(n38984) );
  IV U49247 ( .A(n36385), .Z(n36387) );
  NOR U49248 ( .A(n36387), .B(n36386), .Z(n38985) );
  XOR U49249 ( .A(n38985), .B(n38986), .Z(n38983) );
  XOR U49250 ( .A(n38984), .B(n38983), .Z(n36391) );
  IV U49251 ( .A(n38983), .Z(n36389) );
  NOR U49252 ( .A(n36389), .B(n36388), .Z(n36390) );
  NOR U49253 ( .A(n36391), .B(n36390), .Z(n36392) );
  NOR U49254 ( .A(n42394), .B(n36392), .Z(n36393) );
  IV U49255 ( .A(n36393), .Z(n38979) );
  NOR U49256 ( .A(n36400), .B(n38979), .Z(n38982) );
  IV U49257 ( .A(n36394), .Z(n36395) );
  NOR U49258 ( .A(n36395), .B(n36407), .Z(n36396) );
  IV U49259 ( .A(n36396), .Z(n38981) );
  IV U49260 ( .A(n36397), .Z(n36399) );
  NOR U49261 ( .A(n36399), .B(n36398), .Z(n38978) );
  XOR U49262 ( .A(n38978), .B(n38979), .Z(n49193) );
  XOR U49263 ( .A(n38981), .B(n49193), .Z(n36403) );
  IV U49264 ( .A(n49193), .Z(n36401) );
  NOR U49265 ( .A(n36401), .B(n36400), .Z(n36402) );
  NOR U49266 ( .A(n36403), .B(n36402), .Z(n36404) );
  NOR U49267 ( .A(n38982), .B(n36404), .Z(n39685) );
  IV U49268 ( .A(n36405), .Z(n36406) );
  NOR U49269 ( .A(n36407), .B(n36406), .Z(n39684) );
  IV U49270 ( .A(n36408), .Z(n36410) );
  NOR U49271 ( .A(n36410), .B(n36409), .Z(n39688) );
  NOR U49272 ( .A(n39684), .B(n39688), .Z(n36411) );
  XOR U49273 ( .A(n39685), .B(n36411), .Z(n42385) );
  XOR U49274 ( .A(n38977), .B(n42385), .Z(n36412) );
  IV U49275 ( .A(n36412), .Z(n39697) );
  XOR U49276 ( .A(n39696), .B(n39697), .Z(n39710) );
  XOR U49277 ( .A(n36413), .B(n39710), .Z(n39720) );
  IV U49278 ( .A(n36414), .Z(n36415) );
  NOR U49279 ( .A(n36416), .B(n36415), .Z(n39709) );
  IV U49280 ( .A(n36417), .Z(n36418) );
  NOR U49281 ( .A(n36419), .B(n36418), .Z(n39719) );
  NOR U49282 ( .A(n39709), .B(n39719), .Z(n36420) );
  XOR U49283 ( .A(n39720), .B(n36420), .Z(n36421) );
  IV U49284 ( .A(n36421), .Z(n39718) );
  IV U49285 ( .A(n36422), .Z(n36424) );
  NOR U49286 ( .A(n36424), .B(n36423), .Z(n36425) );
  IV U49287 ( .A(n36425), .Z(n36432) );
  NOR U49288 ( .A(n39718), .B(n36432), .Z(n43124) );
  IV U49289 ( .A(n36426), .Z(n36427) );
  NOR U49290 ( .A(n36439), .B(n36427), .Z(n36428) );
  IV U49291 ( .A(n36428), .Z(n38976) );
  IV U49292 ( .A(n36429), .Z(n36430) );
  NOR U49293 ( .A(n36431), .B(n36430), .Z(n39716) );
  XOR U49294 ( .A(n39716), .B(n39718), .Z(n38975) );
  XOR U49295 ( .A(n38976), .B(n38975), .Z(n36435) );
  IV U49296 ( .A(n38975), .Z(n36433) );
  NOR U49297 ( .A(n36433), .B(n36432), .Z(n36434) );
  NOR U49298 ( .A(n36435), .B(n36434), .Z(n36436) );
  NOR U49299 ( .A(n43124), .B(n36436), .Z(n36437) );
  IV U49300 ( .A(n36437), .Z(n38970) );
  IV U49301 ( .A(n36438), .Z(n36440) );
  NOR U49302 ( .A(n36440), .B(n36439), .Z(n38969) );
  XOR U49303 ( .A(n38970), .B(n38969), .Z(n38973) );
  XOR U49304 ( .A(n38972), .B(n38973), .Z(n38965) );
  XOR U49305 ( .A(n38964), .B(n38965), .Z(n38968) );
  XOR U49306 ( .A(n38967), .B(n38968), .Z(n42358) );
  IV U49307 ( .A(n42358), .Z(n42369) );
  IV U49308 ( .A(n36448), .Z(n42365) );
  NOR U49309 ( .A(n42369), .B(n42365), .Z(n39733) );
  IV U49310 ( .A(n36441), .Z(n36442) );
  NOR U49311 ( .A(n36443), .B(n36442), .Z(n42372) );
  IV U49312 ( .A(n36444), .Z(n36445) );
  NOR U49313 ( .A(n36446), .B(n36445), .Z(n42366) );
  NOR U49314 ( .A(n42372), .B(n42366), .Z(n38963) );
  IV U49315 ( .A(n38963), .Z(n42357) );
  XOR U49316 ( .A(n42357), .B(n42358), .Z(n36447) );
  NOR U49317 ( .A(n36448), .B(n36447), .Z(n39732) );
  NOR U49318 ( .A(n36450), .B(n36449), .Z(n39730) );
  XOR U49319 ( .A(n39732), .B(n39730), .Z(n36451) );
  NOR U49320 ( .A(n39733), .B(n36451), .Z(n39726) );
  XOR U49321 ( .A(n39728), .B(n39726), .Z(n38959) );
  XOR U49322 ( .A(n38957), .B(n38959), .Z(n38961) );
  XOR U49323 ( .A(n36452), .B(n38961), .Z(n39739) );
  IV U49324 ( .A(n36453), .Z(n36454) );
  NOR U49325 ( .A(n36455), .B(n36454), .Z(n39741) );
  IV U49326 ( .A(n36456), .Z(n36458) );
  NOR U49327 ( .A(n36458), .B(n36457), .Z(n39738) );
  NOR U49328 ( .A(n39741), .B(n39738), .Z(n36459) );
  XOR U49329 ( .A(n39739), .B(n36459), .Z(n39746) );
  IV U49330 ( .A(n36460), .Z(n36461) );
  NOR U49331 ( .A(n36462), .B(n36461), .Z(n39744) );
  XOR U49332 ( .A(n39746), .B(n39744), .Z(n39749) );
  XOR U49333 ( .A(n39747), .B(n39749), .Z(n39752) );
  XOR U49334 ( .A(n39751), .B(n39752), .Z(n39756) );
  XOR U49335 ( .A(n39754), .B(n39756), .Z(n38954) );
  IV U49336 ( .A(n36463), .Z(n36465) );
  NOR U49337 ( .A(n36465), .B(n36464), .Z(n36470) );
  IV U49338 ( .A(n36470), .Z(n36466) );
  NOR U49339 ( .A(n38954), .B(n36466), .Z(n43177) );
  IV U49340 ( .A(n36467), .Z(n36469) );
  NOR U49341 ( .A(n36469), .B(n36468), .Z(n38952) );
  XOR U49342 ( .A(n38954), .B(n38952), .Z(n36477) );
  IV U49343 ( .A(n36477), .Z(n36471) );
  NOR U49344 ( .A(n36471), .B(n36470), .Z(n36472) );
  NOR U49345 ( .A(n43177), .B(n36472), .Z(n36479) );
  IV U49346 ( .A(n36479), .Z(n36473) );
  NOR U49347 ( .A(n36474), .B(n36473), .Z(n43181) );
  NOR U49348 ( .A(n36476), .B(n36475), .Z(n36480) );
  IV U49349 ( .A(n36480), .Z(n36478) );
  NOR U49350 ( .A(n36478), .B(n36477), .Z(n38951) );
  NOR U49351 ( .A(n36480), .B(n36479), .Z(n36481) );
  NOR U49352 ( .A(n38951), .B(n36481), .Z(n38948) );
  NOR U49353 ( .A(n36482), .B(n38948), .Z(n36483) );
  NOR U49354 ( .A(n43181), .B(n36483), .Z(n38943) );
  IV U49355 ( .A(n36484), .Z(n36486) );
  NOR U49356 ( .A(n36486), .B(n36485), .Z(n38942) );
  NOR U49357 ( .A(n38947), .B(n38942), .Z(n36487) );
  XOR U49358 ( .A(n38943), .B(n36487), .Z(n39763) );
  XOR U49359 ( .A(n39761), .B(n39763), .Z(n39765) );
  XOR U49360 ( .A(n39764), .B(n39765), .Z(n49102) );
  XOR U49361 ( .A(n38940), .B(n49102), .Z(n39770) );
  XOR U49362 ( .A(n39772), .B(n39770), .Z(n38931) );
  IV U49363 ( .A(n36488), .Z(n36490) );
  NOR U49364 ( .A(n36490), .B(n36489), .Z(n38930) );
  IV U49365 ( .A(n36491), .Z(n36493) );
  NOR U49366 ( .A(n36493), .B(n36492), .Z(n38936) );
  NOR U49367 ( .A(n38930), .B(n38936), .Z(n36494) );
  XOR U49368 ( .A(n38931), .B(n36494), .Z(n38934) );
  XOR U49369 ( .A(n36495), .B(n38934), .Z(n36496) );
  IV U49370 ( .A(n36496), .Z(n38928) );
  XOR U49371 ( .A(n38927), .B(n38928), .Z(n42330) );
  XOR U49372 ( .A(n38920), .B(n42330), .Z(n38921) );
  XOR U49373 ( .A(n38923), .B(n38921), .Z(n38915) );
  XOR U49374 ( .A(n38914), .B(n38915), .Z(n38919) );
  XOR U49375 ( .A(n38917), .B(n38919), .Z(n38910) );
  XOR U49376 ( .A(n38908), .B(n38910), .Z(n38912) );
  XOR U49377 ( .A(n36497), .B(n38912), .Z(n36498) );
  IV U49378 ( .A(n36498), .Z(n38899) );
  NOR U49379 ( .A(n36499), .B(n38898), .Z(n36500) );
  XOR U49380 ( .A(n38899), .B(n36500), .Z(n38894) );
  IV U49381 ( .A(n36501), .Z(n36503) );
  NOR U49382 ( .A(n36503), .B(n36502), .Z(n38893) );
  IV U49383 ( .A(n36504), .Z(n36505) );
  NOR U49384 ( .A(n36508), .B(n36505), .Z(n38891) );
  NOR U49385 ( .A(n38893), .B(n38891), .Z(n36506) );
  XOR U49386 ( .A(n38894), .B(n36506), .Z(n39792) );
  IV U49387 ( .A(n36507), .Z(n36509) );
  NOR U49388 ( .A(n36509), .B(n36508), .Z(n39791) );
  IV U49389 ( .A(n36510), .Z(n36511) );
  NOR U49390 ( .A(n36511), .B(n39797), .Z(n36512) );
  NOR U49391 ( .A(n39791), .B(n36512), .Z(n36513) );
  XOR U49392 ( .A(n39792), .B(n36513), .Z(n39808) );
  XOR U49393 ( .A(n39806), .B(n39808), .Z(n39810) );
  NOR U49394 ( .A(n39809), .B(n36514), .Z(n38887) );
  XOR U49395 ( .A(n39810), .B(n38887), .Z(n38880) );
  XOR U49396 ( .A(n38881), .B(n38880), .Z(n38883) );
  XOR U49397 ( .A(n38882), .B(n38883), .Z(n42294) );
  XOR U49398 ( .A(n38874), .B(n42294), .Z(n38876) );
  IV U49399 ( .A(n36515), .Z(n36517) );
  NOR U49400 ( .A(n36517), .B(n36516), .Z(n42298) );
  NOR U49401 ( .A(n42298), .B(n42292), .Z(n38877) );
  XOR U49402 ( .A(n38876), .B(n38877), .Z(n39821) );
  XOR U49403 ( .A(n36518), .B(n39821), .Z(n39818) );
  IV U49404 ( .A(n36519), .Z(n36520) );
  NOR U49405 ( .A(n36521), .B(n36520), .Z(n36527) );
  IV U49406 ( .A(n36527), .Z(n36522) );
  NOR U49407 ( .A(n39818), .B(n36522), .Z(n39831) );
  IV U49408 ( .A(n36523), .Z(n36525) );
  NOR U49409 ( .A(n36525), .B(n36524), .Z(n39816) );
  XOR U49410 ( .A(n39816), .B(n39818), .Z(n36531) );
  IV U49411 ( .A(n36531), .Z(n36526) );
  NOR U49412 ( .A(n36527), .B(n36526), .Z(n36528) );
  NOR U49413 ( .A(n39831), .B(n36528), .Z(n36529) );
  NOR U49414 ( .A(n36530), .B(n36529), .Z(n36533) );
  IV U49415 ( .A(n36530), .Z(n36532) );
  NOR U49416 ( .A(n36532), .B(n36531), .Z(n39833) );
  NOR U49417 ( .A(n36533), .B(n39833), .Z(n38869) );
  IV U49418 ( .A(n36534), .Z(n36536) );
  NOR U49419 ( .A(n36536), .B(n36535), .Z(n36537) );
  IV U49420 ( .A(n36537), .Z(n38870) );
  XOR U49421 ( .A(n38869), .B(n38870), .Z(n49066) );
  NOR U49422 ( .A(n36541), .B(n49066), .Z(n42278) );
  IV U49423 ( .A(n36538), .Z(n38868) );
  NOR U49424 ( .A(n36540), .B(n36539), .Z(n38872) );
  XOR U49425 ( .A(n38872), .B(n49066), .Z(n38867) );
  XOR U49426 ( .A(n38868), .B(n38867), .Z(n36544) );
  IV U49427 ( .A(n38867), .Z(n36542) );
  NOR U49428 ( .A(n36542), .B(n36541), .Z(n36543) );
  NOR U49429 ( .A(n36544), .B(n36543), .Z(n36545) );
  NOR U49430 ( .A(n42278), .B(n36545), .Z(n39839) );
  XOR U49431 ( .A(n39842), .B(n39839), .Z(n39848) );
  XOR U49432 ( .A(n36546), .B(n39848), .Z(n38865) );
  XOR U49433 ( .A(n38866), .B(n38865), .Z(n39854) );
  XOR U49434 ( .A(n39852), .B(n39854), .Z(n39856) );
  NOR U49435 ( .A(n36554), .B(n39856), .Z(n39859) );
  IV U49436 ( .A(n36547), .Z(n36548) );
  NOR U49437 ( .A(n36549), .B(n36548), .Z(n36550) );
  IV U49438 ( .A(n36550), .Z(n38864) );
  IV U49439 ( .A(n36551), .Z(n36552) );
  NOR U49440 ( .A(n36553), .B(n36552), .Z(n39855) );
  XOR U49441 ( .A(n39855), .B(n39856), .Z(n38863) );
  XOR U49442 ( .A(n38864), .B(n38863), .Z(n36557) );
  IV U49443 ( .A(n38863), .Z(n36555) );
  NOR U49444 ( .A(n36555), .B(n36554), .Z(n36556) );
  NOR U49445 ( .A(n36557), .B(n36556), .Z(n36558) );
  NOR U49446 ( .A(n39859), .B(n36558), .Z(n36559) );
  IV U49447 ( .A(n36559), .Z(n38861) );
  XOR U49448 ( .A(n38860), .B(n38861), .Z(n39868) );
  XOR U49449 ( .A(n39867), .B(n39868), .Z(n39871) );
  IV U49450 ( .A(n39871), .Z(n36567) );
  IV U49451 ( .A(n36560), .Z(n36561) );
  NOR U49452 ( .A(n36562), .B(n36561), .Z(n39870) );
  IV U49453 ( .A(n36563), .Z(n36565) );
  NOR U49454 ( .A(n36565), .B(n36564), .Z(n38857) );
  NOR U49455 ( .A(n39870), .B(n38857), .Z(n36566) );
  XOR U49456 ( .A(n36567), .B(n36566), .Z(n42269) );
  XOR U49457 ( .A(n39874), .B(n42269), .Z(n39876) );
  XOR U49458 ( .A(n39875), .B(n39876), .Z(n39889) );
  XOR U49459 ( .A(n39887), .B(n39889), .Z(n39882) );
  XOR U49460 ( .A(n39880), .B(n39882), .Z(n39898) );
  XOR U49461 ( .A(n36568), .B(n39898), .Z(n36570) );
  NOR U49462 ( .A(n36569), .B(n36570), .Z(n38853) );
  IV U49463 ( .A(n36569), .Z(n36572) );
  IV U49464 ( .A(n36570), .Z(n36571) );
  NOR U49465 ( .A(n36572), .B(n36571), .Z(n46701) );
  NOR U49466 ( .A(n38853), .B(n46701), .Z(n39906) );
  XOR U49467 ( .A(n36573), .B(n39906), .Z(n39915) );
  XOR U49468 ( .A(n36574), .B(n39915), .Z(n38841) );
  XOR U49469 ( .A(n36575), .B(n38841), .Z(n38846) );
  IV U49470 ( .A(n36576), .Z(n36577) );
  NOR U49471 ( .A(n36577), .B(n36585), .Z(n36578) );
  IV U49472 ( .A(n36578), .Z(n36579) );
  NOR U49473 ( .A(n36579), .B(n36584), .Z(n38844) );
  XOR U49474 ( .A(n38846), .B(n38844), .Z(n39927) );
  IV U49475 ( .A(n36580), .Z(n36594) );
  IV U49476 ( .A(n36581), .Z(n36582) );
  NOR U49477 ( .A(n36594), .B(n36582), .Z(n39918) );
  IV U49478 ( .A(n36583), .Z(n36588) );
  NOR U49479 ( .A(n36585), .B(n36584), .Z(n36586) );
  IV U49480 ( .A(n36586), .Z(n36587) );
  NOR U49481 ( .A(n36588), .B(n36587), .Z(n39925) );
  NOR U49482 ( .A(n39918), .B(n39925), .Z(n36589) );
  XOR U49483 ( .A(n39927), .B(n36589), .Z(n38837) );
  IV U49484 ( .A(n36590), .Z(n36591) );
  NOR U49485 ( .A(n36591), .B(n36600), .Z(n38838) );
  IV U49486 ( .A(n36592), .Z(n36593) );
  NOR U49487 ( .A(n36594), .B(n36593), .Z(n39921) );
  NOR U49488 ( .A(n38838), .B(n39921), .Z(n36595) );
  XOR U49489 ( .A(n38837), .B(n36595), .Z(n43380) );
  IV U49490 ( .A(n36596), .Z(n36597) );
  NOR U49491 ( .A(n36598), .B(n36597), .Z(n43383) );
  IV U49492 ( .A(n36599), .Z(n36601) );
  NOR U49493 ( .A(n36601), .B(n36600), .Z(n43378) );
  NOR U49494 ( .A(n43383), .B(n43378), .Z(n38832) );
  XOR U49495 ( .A(n43380), .B(n38832), .Z(n38833) );
  XOR U49496 ( .A(n38835), .B(n38833), .Z(n39936) );
  XOR U49497 ( .A(n36602), .B(n39936), .Z(n36603) );
  IV U49498 ( .A(n36603), .Z(n39939) );
  XOR U49499 ( .A(n39938), .B(n39939), .Z(n42231) );
  IV U49500 ( .A(n36604), .Z(n36605) );
  NOR U49501 ( .A(n36606), .B(n36605), .Z(n42238) );
  IV U49502 ( .A(n36607), .Z(n36608) );
  NOR U49503 ( .A(n42228), .B(n36608), .Z(n45568) );
  NOR U49504 ( .A(n42238), .B(n45568), .Z(n39950) );
  XOR U49505 ( .A(n42231), .B(n39950), .Z(n39942) );
  XOR U49506 ( .A(n39944), .B(n39942), .Z(n39947) );
  XOR U49507 ( .A(n39946), .B(n39947), .Z(n39960) );
  IV U49508 ( .A(n36609), .Z(n36610) );
  NOR U49509 ( .A(n36611), .B(n36610), .Z(n39957) );
  IV U49510 ( .A(n36612), .Z(n36613) );
  NOR U49511 ( .A(n36614), .B(n36613), .Z(n39959) );
  NOR U49512 ( .A(n39957), .B(n39959), .Z(n36615) );
  XOR U49513 ( .A(n39960), .B(n36615), .Z(n38814) );
  NOR U49514 ( .A(n36616), .B(n38823), .Z(n36619) );
  NOR U49515 ( .A(n36617), .B(n38816), .Z(n36618) );
  NOR U49516 ( .A(n36619), .B(n36618), .Z(n36620) );
  XOR U49517 ( .A(n38814), .B(n36620), .Z(n38812) );
  XOR U49518 ( .A(n38810), .B(n38812), .Z(n42204) );
  XOR U49519 ( .A(n38809), .B(n42204), .Z(n39965) );
  XOR U49520 ( .A(n39967), .B(n39965), .Z(n39969) );
  XOR U49521 ( .A(n39968), .B(n39969), .Z(n38807) );
  NOR U49522 ( .A(n36622), .B(n36621), .Z(n38806) );
  NOR U49523 ( .A(n38806), .B(n38804), .Z(n36623) );
  XOR U49524 ( .A(n38807), .B(n36623), .Z(n38798) );
  XOR U49525 ( .A(n36624), .B(n38798), .Z(n38796) );
  IV U49526 ( .A(n36625), .Z(n36627) );
  NOR U49527 ( .A(n36627), .B(n36626), .Z(n38795) );
  IV U49528 ( .A(n36628), .Z(n36630) );
  NOR U49529 ( .A(n36630), .B(n36629), .Z(n38793) );
  NOR U49530 ( .A(n38795), .B(n38793), .Z(n36631) );
  XOR U49531 ( .A(n38796), .B(n36631), .Z(n36632) );
  IV U49532 ( .A(n36632), .Z(n38789) );
  XOR U49533 ( .A(n38787), .B(n38789), .Z(n38792) );
  IV U49534 ( .A(n36633), .Z(n36634) );
  NOR U49535 ( .A(n36635), .B(n36634), .Z(n38790) );
  XOR U49536 ( .A(n38792), .B(n38790), .Z(n42180) );
  IV U49537 ( .A(n36636), .Z(n36637) );
  NOR U49538 ( .A(n36638), .B(n36637), .Z(n42178) );
  IV U49539 ( .A(n36639), .Z(n36641) );
  NOR U49540 ( .A(n36641), .B(n36640), .Z(n43430) );
  NOR U49541 ( .A(n42178), .B(n43430), .Z(n39975) );
  IV U49542 ( .A(n39975), .Z(n39973) );
  XOR U49543 ( .A(n42180), .B(n39973), .Z(n43437) );
  XOR U49544 ( .A(n36642), .B(n43437), .Z(n36643) );
  IV U49545 ( .A(n36643), .Z(n39985) );
  XOR U49546 ( .A(n39983), .B(n39985), .Z(n45539) );
  IV U49547 ( .A(n45539), .Z(n36650) );
  IV U49548 ( .A(n36644), .Z(n36646) );
  NOR U49549 ( .A(n36646), .B(n36645), .Z(n46814) );
  IV U49550 ( .A(n36647), .Z(n36648) );
  NOR U49551 ( .A(n36649), .B(n36648), .Z(n45535) );
  NOR U49552 ( .A(n46814), .B(n45535), .Z(n39986) );
  XOR U49553 ( .A(n36650), .B(n39986), .Z(n38783) );
  XOR U49554 ( .A(n36651), .B(n38783), .Z(n36657) );
  NOR U49555 ( .A(n36652), .B(n36657), .Z(n39998) );
  IV U49556 ( .A(n36653), .Z(n36655) );
  IV U49557 ( .A(n36654), .Z(n36662) );
  NOR U49558 ( .A(n36655), .B(n36662), .Z(n36659) );
  IV U49559 ( .A(n36659), .Z(n36656) );
  NOR U49560 ( .A(n38783), .B(n36656), .Z(n42167) );
  IV U49561 ( .A(n36657), .Z(n36658) );
  NOR U49562 ( .A(n36659), .B(n36658), .Z(n36660) );
  NOR U49563 ( .A(n42167), .B(n36660), .Z(n36661) );
  IV U49564 ( .A(n36661), .Z(n39993) );
  NOR U49565 ( .A(n36663), .B(n36662), .Z(n36664) );
  IV U49566 ( .A(n36664), .Z(n36665) );
  NOR U49567 ( .A(n36666), .B(n36665), .Z(n36667) );
  IV U49568 ( .A(n36667), .Z(n36668) );
  NOR U49569 ( .A(n36669), .B(n36668), .Z(n36670) );
  IV U49570 ( .A(n36670), .Z(n39992) );
  XOR U49571 ( .A(n39993), .B(n39992), .Z(n36671) );
  NOR U49572 ( .A(n36672), .B(n36671), .Z(n36673) );
  NOR U49573 ( .A(n39998), .B(n36673), .Z(n38779) );
  IV U49574 ( .A(n36674), .Z(n36676) );
  NOR U49575 ( .A(n36676), .B(n36675), .Z(n36677) );
  IV U49576 ( .A(n36677), .Z(n38780) );
  XOR U49577 ( .A(n38779), .B(n38780), .Z(n38777) );
  NOR U49578 ( .A(n36678), .B(n38777), .Z(n43449) );
  IV U49579 ( .A(n36679), .Z(n36680) );
  NOR U49580 ( .A(n36681), .B(n36680), .Z(n38776) );
  XOR U49581 ( .A(n38776), .B(n38777), .Z(n36686) );
  IV U49582 ( .A(n36686), .Z(n36682) );
  NOR U49583 ( .A(n36683), .B(n36682), .Z(n36684) );
  NOR U49584 ( .A(n43449), .B(n36684), .Z(n38771) );
  NOR U49585 ( .A(n36685), .B(n38771), .Z(n36688) );
  IV U49586 ( .A(n36685), .Z(n36687) );
  NOR U49587 ( .A(n36687), .B(n36686), .Z(n42161) );
  NOR U49588 ( .A(n36688), .B(n42161), .Z(n40011) );
  NOR U49589 ( .A(n36689), .B(n38773), .Z(n36694) );
  XOR U49590 ( .A(n36690), .B(n38773), .Z(n36693) );
  IV U49591 ( .A(n36691), .Z(n36692) );
  NOR U49592 ( .A(n36693), .B(n36692), .Z(n40012) );
  NOR U49593 ( .A(n36694), .B(n40012), .Z(n36695) );
  XOR U49594 ( .A(n40011), .B(n36695), .Z(n40019) );
  IV U49595 ( .A(n40019), .Z(n36708) );
  IV U49596 ( .A(n36696), .Z(n36698) );
  NOR U49597 ( .A(n36698), .B(n36697), .Z(n40009) );
  IV U49598 ( .A(n36699), .Z(n36706) );
  NOR U49599 ( .A(n36701), .B(n36700), .Z(n36702) );
  IV U49600 ( .A(n36702), .Z(n36703) );
  NOR U49601 ( .A(n36704), .B(n36703), .Z(n36705) );
  IV U49602 ( .A(n36705), .Z(n36710) );
  NOR U49603 ( .A(n36706), .B(n36710), .Z(n40017) );
  NOR U49604 ( .A(n40009), .B(n40017), .Z(n36707) );
  XOR U49605 ( .A(n36708), .B(n36707), .Z(n38766) );
  IV U49606 ( .A(n36709), .Z(n36711) );
  NOR U49607 ( .A(n36711), .B(n36710), .Z(n38764) );
  XOR U49608 ( .A(n38766), .B(n38764), .Z(n38768) );
  XOR U49609 ( .A(n38767), .B(n38768), .Z(n43470) );
  NOR U49610 ( .A(n36712), .B(n43468), .Z(n36713) );
  NOR U49611 ( .A(n36714), .B(n36713), .Z(n40021) );
  XOR U49612 ( .A(n43470), .B(n40021), .Z(n40025) );
  IV U49613 ( .A(n36715), .Z(n36718) );
  IV U49614 ( .A(n36716), .Z(n36717) );
  NOR U49615 ( .A(n36718), .B(n36717), .Z(n40023) );
  XOR U49616 ( .A(n40025), .B(n40023), .Z(n40035) );
  IV U49617 ( .A(n36719), .Z(n36720) );
  NOR U49618 ( .A(n36721), .B(n36720), .Z(n40034) );
  IV U49619 ( .A(n36722), .Z(n36724) );
  NOR U49620 ( .A(n36724), .B(n36723), .Z(n40029) );
  NOR U49621 ( .A(n40034), .B(n40029), .Z(n36725) );
  XOR U49622 ( .A(n40035), .B(n36725), .Z(n38755) );
  XOR U49623 ( .A(n38755), .B(n36726), .Z(n38759) );
  XOR U49624 ( .A(n38758), .B(n38759), .Z(n40048) );
  XOR U49625 ( .A(n40047), .B(n40048), .Z(n40051) );
  XOR U49626 ( .A(n40050), .B(n40051), .Z(n38751) );
  XOR U49627 ( .A(n38750), .B(n38751), .Z(n42115) );
  XOR U49628 ( .A(n38753), .B(n42115), .Z(n38745) );
  XOR U49629 ( .A(n38744), .B(n38745), .Z(n38748) );
  IV U49630 ( .A(n38748), .Z(n36734) );
  IV U49631 ( .A(n36727), .Z(n36728) );
  NOR U49632 ( .A(n36729), .B(n36728), .Z(n38741) );
  IV U49633 ( .A(n36730), .Z(n36732) );
  NOR U49634 ( .A(n36732), .B(n36731), .Z(n38746) );
  NOR U49635 ( .A(n38741), .B(n38746), .Z(n36733) );
  XOR U49636 ( .A(n36734), .B(n36733), .Z(n38738) );
  XOR U49637 ( .A(n38736), .B(n38738), .Z(n40060) );
  XOR U49638 ( .A(n36735), .B(n40060), .Z(n36736) );
  IV U49639 ( .A(n36736), .Z(n40063) );
  XOR U49640 ( .A(n40061), .B(n40063), .Z(n40066) );
  IV U49641 ( .A(n36737), .Z(n36739) );
  NOR U49642 ( .A(n36739), .B(n36738), .Z(n40064) );
  XOR U49643 ( .A(n40066), .B(n40064), .Z(n38734) );
  XOR U49644 ( .A(n38733), .B(n38734), .Z(n38730) );
  IV U49645 ( .A(n36740), .Z(n36741) );
  NOR U49646 ( .A(n36742), .B(n36741), .Z(n38731) );
  IV U49647 ( .A(n36743), .Z(n36744) );
  NOR U49648 ( .A(n36744), .B(n36750), .Z(n38728) );
  NOR U49649 ( .A(n38731), .B(n38728), .Z(n36745) );
  XOR U49650 ( .A(n38730), .B(n36745), .Z(n38719) );
  IV U49651 ( .A(n36746), .Z(n36747) );
  NOR U49652 ( .A(n36748), .B(n36747), .Z(n38720) );
  IV U49653 ( .A(n36749), .Z(n36751) );
  NOR U49654 ( .A(n36751), .B(n36750), .Z(n38725) );
  NOR U49655 ( .A(n38720), .B(n38725), .Z(n36752) );
  XOR U49656 ( .A(n38719), .B(n36752), .Z(n38723) );
  IV U49657 ( .A(n36753), .Z(n36754) );
  NOR U49658 ( .A(n36755), .B(n36754), .Z(n38722) );
  IV U49659 ( .A(n36756), .Z(n36758) );
  NOR U49660 ( .A(n36758), .B(n36757), .Z(n38717) );
  NOR U49661 ( .A(n38722), .B(n38717), .Z(n36759) );
  XOR U49662 ( .A(n38723), .B(n36759), .Z(n38714) );
  XOR U49663 ( .A(n38715), .B(n38714), .Z(n40072) );
  XOR U49664 ( .A(n40070), .B(n40072), .Z(n40074) );
  NOR U49665 ( .A(n36767), .B(n40074), .Z(n42072) );
  IV U49666 ( .A(n36760), .Z(n36762) );
  NOR U49667 ( .A(n36762), .B(n36761), .Z(n36763) );
  IV U49668 ( .A(n36763), .Z(n38710) );
  IV U49669 ( .A(n36764), .Z(n36765) );
  NOR U49670 ( .A(n36766), .B(n36765), .Z(n40073) );
  XOR U49671 ( .A(n40073), .B(n40074), .Z(n38709) );
  XOR U49672 ( .A(n38710), .B(n38709), .Z(n36770) );
  IV U49673 ( .A(n38709), .Z(n36768) );
  NOR U49674 ( .A(n36768), .B(n36767), .Z(n36769) );
  NOR U49675 ( .A(n36770), .B(n36769), .Z(n36771) );
  NOR U49676 ( .A(n42072), .B(n36771), .Z(n36772) );
  IV U49677 ( .A(n36772), .Z(n38705) );
  NOR U49678 ( .A(n36778), .B(n38705), .Z(n42066) );
  NOR U49679 ( .A(n36773), .B(n38706), .Z(n36774) );
  XOR U49680 ( .A(n36774), .B(n38705), .Z(n38703) );
  IV U49681 ( .A(n36775), .Z(n36777) );
  NOR U49682 ( .A(n36777), .B(n36776), .Z(n36779) );
  IV U49683 ( .A(n36779), .Z(n38702) );
  XOR U49684 ( .A(n38703), .B(n38702), .Z(n36781) );
  NOR U49685 ( .A(n36779), .B(n36778), .Z(n36780) );
  NOR U49686 ( .A(n36781), .B(n36780), .Z(n36782) );
  NOR U49687 ( .A(n42066), .B(n36782), .Z(n40080) );
  XOR U49688 ( .A(n40082), .B(n40080), .Z(n40088) );
  NOR U49689 ( .A(n43532), .B(n40088), .Z(n38701) );
  IV U49690 ( .A(n36783), .Z(n36785) );
  NOR U49691 ( .A(n36785), .B(n36784), .Z(n40083) );
  IV U49692 ( .A(n36786), .Z(n36788) );
  NOR U49693 ( .A(n36788), .B(n36787), .Z(n40087) );
  NOR U49694 ( .A(n40083), .B(n40087), .Z(n36789) );
  XOR U49695 ( .A(n36789), .B(n40088), .Z(n43527) );
  NOR U49696 ( .A(n36790), .B(n43527), .Z(n36791) );
  NOR U49697 ( .A(n38701), .B(n36791), .Z(n36792) );
  IV U49698 ( .A(n36792), .Z(n38699) );
  NOR U49699 ( .A(n36794), .B(n36793), .Z(n38698) );
  XOR U49700 ( .A(n38699), .B(n38698), .Z(n38693) );
  XOR U49701 ( .A(n38692), .B(n38693), .Z(n38697) );
  XOR U49702 ( .A(n36795), .B(n38697), .Z(n36796) );
  IV U49703 ( .A(n36796), .Z(n38691) );
  IV U49704 ( .A(n36797), .Z(n36799) );
  NOR U49705 ( .A(n36799), .B(n36798), .Z(n38689) );
  XOR U49706 ( .A(n38691), .B(n38689), .Z(n40094) );
  IV U49707 ( .A(n40094), .Z(n36806) );
  IV U49708 ( .A(n36800), .Z(n36801) );
  NOR U49709 ( .A(n36809), .B(n36801), .Z(n38685) );
  IV U49710 ( .A(n36802), .Z(n36804) );
  NOR U49711 ( .A(n36804), .B(n36803), .Z(n40093) );
  NOR U49712 ( .A(n38685), .B(n40093), .Z(n36805) );
  XOR U49713 ( .A(n36806), .B(n36805), .Z(n40098) );
  IV U49714 ( .A(n36807), .Z(n36808) );
  NOR U49715 ( .A(n36809), .B(n36808), .Z(n40096) );
  XOR U49716 ( .A(n40098), .B(n40096), .Z(n40101) );
  XOR U49717 ( .A(n36810), .B(n40101), .Z(n40103) );
  IV U49718 ( .A(n36811), .Z(n36813) );
  NOR U49719 ( .A(n36813), .B(n36812), .Z(n40107) );
  IV U49720 ( .A(n36814), .Z(n36815) );
  NOR U49721 ( .A(n36816), .B(n36815), .Z(n40104) );
  NOR U49722 ( .A(n40107), .B(n40104), .Z(n36817) );
  XOR U49723 ( .A(n40103), .B(n36817), .Z(n38680) );
  XOR U49724 ( .A(n38679), .B(n38680), .Z(n40117) );
  XOR U49725 ( .A(n40116), .B(n40117), .Z(n38675) );
  XOR U49726 ( .A(n36818), .B(n38675), .Z(n36819) );
  IV U49727 ( .A(n36819), .Z(n38670) );
  XOR U49728 ( .A(n38668), .B(n38670), .Z(n38672) );
  IV U49729 ( .A(n36820), .Z(n36822) );
  NOR U49730 ( .A(n36822), .B(n36821), .Z(n38665) );
  NOR U49731 ( .A(n38671), .B(n38665), .Z(n36823) );
  XOR U49732 ( .A(n38672), .B(n36823), .Z(n38663) );
  XOR U49733 ( .A(n38664), .B(n38663), .Z(n42025) );
  IV U49734 ( .A(n36824), .Z(n36830) );
  NOR U49735 ( .A(n36825), .B(n36836), .Z(n36826) );
  IV U49736 ( .A(n36826), .Z(n36827) );
  NOR U49737 ( .A(n36828), .B(n36827), .Z(n36829) );
  IV U49738 ( .A(n36829), .Z(n36832) );
  NOR U49739 ( .A(n36830), .B(n36832), .Z(n42026) );
  IV U49740 ( .A(n36831), .Z(n36833) );
  NOR U49741 ( .A(n36833), .B(n36832), .Z(n38661) );
  NOR U49742 ( .A(n42026), .B(n38661), .Z(n36834) );
  XOR U49743 ( .A(n42025), .B(n36834), .Z(n38654) );
  XOR U49744 ( .A(n38656), .B(n38654), .Z(n38658) );
  XOR U49745 ( .A(n38657), .B(n38658), .Z(n38652) );
  NOR U49746 ( .A(n36841), .B(n38652), .Z(n42017) );
  IV U49747 ( .A(n36835), .Z(n36837) );
  NOR U49748 ( .A(n36837), .B(n36836), .Z(n38651) );
  XOR U49749 ( .A(n38651), .B(n38652), .Z(n38650) );
  IV U49750 ( .A(n36838), .Z(n36839) );
  NOR U49751 ( .A(n36840), .B(n36839), .Z(n36842) );
  IV U49752 ( .A(n36842), .Z(n38649) );
  XOR U49753 ( .A(n38650), .B(n38649), .Z(n36844) );
  NOR U49754 ( .A(n36842), .B(n36841), .Z(n36843) );
  NOR U49755 ( .A(n36844), .B(n36843), .Z(n36845) );
  NOR U49756 ( .A(n42017), .B(n36845), .Z(n36846) );
  IV U49757 ( .A(n36846), .Z(n38644) );
  XOR U49758 ( .A(n38643), .B(n38644), .Z(n38647) );
  NOR U49759 ( .A(n36852), .B(n38647), .Z(n42007) );
  NOR U49760 ( .A(n36848), .B(n36847), .Z(n36849) );
  IV U49761 ( .A(n36849), .Z(n40126) );
  NOR U49762 ( .A(n36851), .B(n36850), .Z(n38646) );
  XOR U49763 ( .A(n38646), .B(n38647), .Z(n40125) );
  XOR U49764 ( .A(n40126), .B(n40125), .Z(n36855) );
  IV U49765 ( .A(n40125), .Z(n36853) );
  NOR U49766 ( .A(n36853), .B(n36852), .Z(n36854) );
  NOR U49767 ( .A(n36855), .B(n36854), .Z(n36856) );
  NOR U49768 ( .A(n42007), .B(n36856), .Z(n40128) );
  XOR U49769 ( .A(n36857), .B(n40128), .Z(n40135) );
  NOR U49770 ( .A(n36858), .B(n40135), .Z(n42005) );
  IV U49771 ( .A(n36859), .Z(n36861) );
  NOR U49772 ( .A(n36861), .B(n36860), .Z(n40134) );
  XOR U49773 ( .A(n40134), .B(n40135), .Z(n36867) );
  IV U49774 ( .A(n36867), .Z(n36862) );
  NOR U49775 ( .A(n36863), .B(n36862), .Z(n36864) );
  NOR U49776 ( .A(n42005), .B(n36864), .Z(n36865) );
  NOR U49777 ( .A(n36866), .B(n36865), .Z(n36869) );
  IV U49778 ( .A(n36866), .Z(n36868) );
  NOR U49779 ( .A(n36868), .B(n36867), .Z(n45420) );
  NOR U49780 ( .A(n36869), .B(n45420), .Z(n36870) );
  IV U49781 ( .A(n36870), .Z(n38641) );
  XOR U49782 ( .A(n38640), .B(n38641), .Z(n40147) );
  IV U49783 ( .A(n36871), .Z(n36872) );
  NOR U49784 ( .A(n36873), .B(n36872), .Z(n40141) );
  IV U49785 ( .A(n36874), .Z(n36878) );
  NOR U49786 ( .A(n36876), .B(n36875), .Z(n36877) );
  IV U49787 ( .A(n36877), .Z(n36882) );
  NOR U49788 ( .A(n36878), .B(n36882), .Z(n40145) );
  NOR U49789 ( .A(n40141), .B(n40145), .Z(n36879) );
  XOR U49790 ( .A(n40147), .B(n36879), .Z(n36880) );
  IV U49791 ( .A(n36880), .Z(n38639) );
  IV U49792 ( .A(n36881), .Z(n36883) );
  NOR U49793 ( .A(n36883), .B(n36882), .Z(n36884) );
  IV U49794 ( .A(n36884), .Z(n38638) );
  XOR U49795 ( .A(n38639), .B(n38638), .Z(n40153) );
  XOR U49796 ( .A(n40152), .B(n40153), .Z(n40162) );
  XOR U49797 ( .A(n36885), .B(n40162), .Z(n36886) );
  IV U49798 ( .A(n36886), .Z(n40168) );
  XOR U49799 ( .A(n40159), .B(n40168), .Z(n38637) );
  IV U49800 ( .A(n36887), .Z(n36889) );
  NOR U49801 ( .A(n36889), .B(n36888), .Z(n40166) );
  IV U49802 ( .A(n36890), .Z(n36891) );
  NOR U49803 ( .A(n36891), .B(n36898), .Z(n38635) );
  NOR U49804 ( .A(n40166), .B(n38635), .Z(n36892) );
  XOR U49805 ( .A(n38637), .B(n36892), .Z(n38629) );
  IV U49806 ( .A(n36893), .Z(n36894) );
  NOR U49807 ( .A(n36895), .B(n36894), .Z(n38630) );
  IV U49808 ( .A(n36896), .Z(n36897) );
  NOR U49809 ( .A(n36898), .B(n36897), .Z(n38632) );
  NOR U49810 ( .A(n38630), .B(n38632), .Z(n36899) );
  XOR U49811 ( .A(n38629), .B(n36899), .Z(n40170) );
  XOR U49812 ( .A(n40169), .B(n40170), .Z(n40174) );
  IV U49813 ( .A(n36900), .Z(n36901) );
  NOR U49814 ( .A(n36902), .B(n36901), .Z(n40172) );
  XOR U49815 ( .A(n40174), .B(n40172), .Z(n38627) );
  XOR U49816 ( .A(n38624), .B(n38627), .Z(n38622) );
  IV U49817 ( .A(n38622), .Z(n36909) );
  IV U49818 ( .A(n36903), .Z(n36904) );
  NOR U49819 ( .A(n36905), .B(n36904), .Z(n38626) );
  IV U49820 ( .A(n36906), .Z(n36907) );
  NOR U49821 ( .A(n36907), .B(n36912), .Z(n38621) );
  NOR U49822 ( .A(n38626), .B(n38621), .Z(n36908) );
  XOR U49823 ( .A(n36909), .B(n36908), .Z(n38620) );
  IV U49824 ( .A(n36910), .Z(n36911) );
  NOR U49825 ( .A(n36912), .B(n36911), .Z(n38618) );
  XOR U49826 ( .A(n38620), .B(n38618), .Z(n38614) );
  XOR U49827 ( .A(n38612), .B(n38614), .Z(n38616) );
  XOR U49828 ( .A(n38615), .B(n38616), .Z(n36918) );
  NOR U49829 ( .A(n36913), .B(n36918), .Z(n40182) );
  IV U49830 ( .A(n36914), .Z(n36916) );
  NOR U49831 ( .A(n36916), .B(n36915), .Z(n36920) );
  IV U49832 ( .A(n36920), .Z(n36917) );
  NOR U49833 ( .A(n36917), .B(n38616), .Z(n40185) );
  IV U49834 ( .A(n36918), .Z(n36919) );
  NOR U49835 ( .A(n36920), .B(n36919), .Z(n36921) );
  NOR U49836 ( .A(n40185), .B(n36921), .Z(n36926) );
  NOR U49837 ( .A(n36922), .B(n36926), .Z(n36923) );
  NOR U49838 ( .A(n40182), .B(n36923), .Z(n36924) );
  NOR U49839 ( .A(n36925), .B(n36924), .Z(n36929) );
  IV U49840 ( .A(n36925), .Z(n36928) );
  IV U49841 ( .A(n36926), .Z(n36927) );
  NOR U49842 ( .A(n36928), .B(n36927), .Z(n41972) );
  NOR U49843 ( .A(n36929), .B(n41972), .Z(n36930) );
  IV U49844 ( .A(n36930), .Z(n40191) );
  IV U49845 ( .A(n36931), .Z(n36933) );
  NOR U49846 ( .A(n36933), .B(n36932), .Z(n40190) );
  XOR U49847 ( .A(n40191), .B(n40190), .Z(n40195) );
  XOR U49848 ( .A(n40194), .B(n40195), .Z(n40198) );
  XOR U49849 ( .A(n40197), .B(n40198), .Z(n40202) );
  XOR U49850 ( .A(n40201), .B(n40202), .Z(n40204) );
  XOR U49851 ( .A(n40205), .B(n40204), .Z(n36943) );
  IV U49852 ( .A(n36943), .Z(n36934) );
  NOR U49853 ( .A(n36946), .B(n36934), .Z(n41956) );
  IV U49854 ( .A(n36935), .Z(n36937) );
  NOR U49855 ( .A(n36937), .B(n36936), .Z(n36938) );
  IV U49856 ( .A(n36938), .Z(n40209) );
  IV U49857 ( .A(n36939), .Z(n36941) );
  NOR U49858 ( .A(n36941), .B(n36940), .Z(n36944) );
  IV U49859 ( .A(n36944), .Z(n36942) );
  NOR U49860 ( .A(n36942), .B(n40204), .Z(n41961) );
  NOR U49861 ( .A(n36944), .B(n36943), .Z(n36945) );
  NOR U49862 ( .A(n41961), .B(n36945), .Z(n36947) );
  IV U49863 ( .A(n36947), .Z(n40208) );
  XOR U49864 ( .A(n40209), .B(n40208), .Z(n36949) );
  NOR U49865 ( .A(n36947), .B(n36946), .Z(n36948) );
  NOR U49866 ( .A(n36949), .B(n36948), .Z(n36950) );
  NOR U49867 ( .A(n41956), .B(n36950), .Z(n36951) );
  IV U49868 ( .A(n36951), .Z(n40211) );
  IV U49869 ( .A(n36952), .Z(n36954) );
  NOR U49870 ( .A(n36954), .B(n36953), .Z(n40210) );
  XOR U49871 ( .A(n40211), .B(n40210), .Z(n40215) );
  XOR U49872 ( .A(n36955), .B(n40215), .Z(n36963) );
  IV U49873 ( .A(n36963), .Z(n41944) );
  XOR U49874 ( .A(n36956), .B(n41944), .Z(n36966) );
  IV U49875 ( .A(n36966), .Z(n36957) );
  NOR U49876 ( .A(n36958), .B(n36957), .Z(n41939) );
  IV U49877 ( .A(n36959), .Z(n36960) );
  NOR U49878 ( .A(n36961), .B(n36960), .Z(n36967) );
  IV U49879 ( .A(n36967), .Z(n36965) );
  IV U49880 ( .A(n36962), .Z(n38609) );
  XOR U49881 ( .A(n38609), .B(n36963), .Z(n36964) );
  NOR U49882 ( .A(n36965), .B(n36964), .Z(n43680) );
  NOR U49883 ( .A(n36967), .B(n36966), .Z(n36968) );
  NOR U49884 ( .A(n43680), .B(n36968), .Z(n38600) );
  NOR U49885 ( .A(n36969), .B(n38600), .Z(n36970) );
  NOR U49886 ( .A(n41939), .B(n36970), .Z(n38604) );
  IV U49887 ( .A(n36971), .Z(n36972) );
  NOR U49888 ( .A(n36973), .B(n36972), .Z(n38603) );
  IV U49889 ( .A(n36974), .Z(n36976) );
  NOR U49890 ( .A(n36976), .B(n36975), .Z(n38599) );
  NOR U49891 ( .A(n38603), .B(n38599), .Z(n36977) );
  XOR U49892 ( .A(n38604), .B(n36977), .Z(n40222) );
  IV U49893 ( .A(n36978), .Z(n36979) );
  NOR U49894 ( .A(n36980), .B(n36979), .Z(n40220) );
  XOR U49895 ( .A(n40222), .B(n40220), .Z(n40224) );
  XOR U49896 ( .A(n40223), .B(n40224), .Z(n40229) );
  XOR U49897 ( .A(n36981), .B(n40229), .Z(n38591) );
  XOR U49898 ( .A(n38592), .B(n38591), .Z(n38594) );
  XOR U49899 ( .A(n36982), .B(n38594), .Z(n36983) );
  IV U49900 ( .A(n36983), .Z(n38588) );
  XOR U49901 ( .A(n38586), .B(n38588), .Z(n38582) );
  IV U49902 ( .A(n36984), .Z(n36985) );
  NOR U49903 ( .A(n36985), .B(n36987), .Z(n38580) );
  XOR U49904 ( .A(n38582), .B(n38580), .Z(n38585) );
  IV U49905 ( .A(n36986), .Z(n36988) );
  NOR U49906 ( .A(n36988), .B(n36987), .Z(n38583) );
  XOR U49907 ( .A(n38585), .B(n38583), .Z(n41911) );
  IV U49908 ( .A(n41911), .Z(n36997) );
  IV U49909 ( .A(n36991), .Z(n36989) );
  NOR U49910 ( .A(n36990), .B(n36989), .Z(n41909) );
  XOR U49911 ( .A(n36991), .B(n36990), .Z(n36992) );
  NOR U49912 ( .A(n36993), .B(n36992), .Z(n36994) );
  IV U49913 ( .A(n36994), .Z(n36995) );
  NOR U49914 ( .A(n36996), .B(n36995), .Z(n43703) );
  NOR U49915 ( .A(n41909), .B(n43703), .Z(n40236) );
  XOR U49916 ( .A(n36997), .B(n40236), .Z(n38578) );
  XOR U49917 ( .A(n38577), .B(n38578), .Z(n40244) );
  XOR U49918 ( .A(n40245), .B(n40244), .Z(n40251) );
  IV U49919 ( .A(n36998), .Z(n37000) );
  NOR U49920 ( .A(n37000), .B(n36999), .Z(n40252) );
  XOR U49921 ( .A(n40251), .B(n40252), .Z(n40256) );
  IV U49922 ( .A(n37001), .Z(n37002) );
  NOR U49923 ( .A(n37003), .B(n37002), .Z(n40255) );
  IV U49924 ( .A(n37004), .Z(n37005) );
  NOR U49925 ( .A(n37006), .B(n37005), .Z(n40261) );
  NOR U49926 ( .A(n40255), .B(n40261), .Z(n37007) );
  XOR U49927 ( .A(n40256), .B(n37007), .Z(n40260) );
  IV U49928 ( .A(n37008), .Z(n37010) );
  NOR U49929 ( .A(n37010), .B(n37009), .Z(n37011) );
  IV U49930 ( .A(n37011), .Z(n37019) );
  NOR U49931 ( .A(n40260), .B(n37019), .Z(n41903) );
  IV U49932 ( .A(n37012), .Z(n37014) );
  NOR U49933 ( .A(n37014), .B(n37013), .Z(n37015) );
  IV U49934 ( .A(n37015), .Z(n38576) );
  IV U49935 ( .A(n37016), .Z(n37018) );
  NOR U49936 ( .A(n37018), .B(n37017), .Z(n40258) );
  XOR U49937 ( .A(n40258), .B(n40260), .Z(n38575) );
  XOR U49938 ( .A(n38576), .B(n38575), .Z(n37022) );
  IV U49939 ( .A(n38575), .Z(n37020) );
  NOR U49940 ( .A(n37020), .B(n37019), .Z(n37021) );
  NOR U49941 ( .A(n37022), .B(n37021), .Z(n37023) );
  NOR U49942 ( .A(n41903), .B(n37023), .Z(n37024) );
  IV U49943 ( .A(n37024), .Z(n40268) );
  XOR U49944 ( .A(n40267), .B(n40268), .Z(n38573) );
  XOR U49945 ( .A(n38572), .B(n38573), .Z(n43726) );
  XOR U49946 ( .A(n40273), .B(n43726), .Z(n40275) );
  XOR U49947 ( .A(n37025), .B(n40275), .Z(n40283) );
  IV U49948 ( .A(n37026), .Z(n37028) );
  NOR U49949 ( .A(n37028), .B(n37027), .Z(n40281) );
  XOR U49950 ( .A(n40283), .B(n40281), .Z(n40289) );
  IV U49951 ( .A(n40289), .Z(n37036) );
  IV U49952 ( .A(n37029), .Z(n37031) );
  NOR U49953 ( .A(n37031), .B(n37030), .Z(n40286) );
  IV U49954 ( .A(n37032), .Z(n37033) );
  NOR U49955 ( .A(n37034), .B(n37033), .Z(n40288) );
  NOR U49956 ( .A(n40286), .B(n40288), .Z(n37035) );
  XOR U49957 ( .A(n37036), .B(n37035), .Z(n40293) );
  IV U49958 ( .A(n37037), .Z(n37039) );
  NOR U49959 ( .A(n37039), .B(n37038), .Z(n40291) );
  XOR U49960 ( .A(n40293), .B(n40291), .Z(n40295) );
  XOR U49961 ( .A(n40294), .B(n40295), .Z(n40303) );
  XOR U49962 ( .A(n40302), .B(n40303), .Z(n40306) );
  XOR U49963 ( .A(n37040), .B(n40306), .Z(n37041) );
  IV U49964 ( .A(n37041), .Z(n43746) );
  XOR U49965 ( .A(n37042), .B(n43746), .Z(n41873) );
  XOR U49966 ( .A(n40313), .B(n41873), .Z(n40315) );
  IV U49967 ( .A(n37043), .Z(n37044) );
  NOR U49968 ( .A(n37045), .B(n37044), .Z(n40320) );
  NOR U49969 ( .A(n40314), .B(n40320), .Z(n37046) );
  XOR U49970 ( .A(n40315), .B(n37046), .Z(n41868) );
  XOR U49971 ( .A(n38567), .B(n41868), .Z(n38569) );
  IV U49972 ( .A(n37047), .Z(n37049) );
  NOR U49973 ( .A(n37049), .B(n37048), .Z(n40325) );
  IV U49974 ( .A(n37050), .Z(n37052) );
  NOR U49975 ( .A(n37052), .B(n37051), .Z(n38568) );
  NOR U49976 ( .A(n40325), .B(n38568), .Z(n37053) );
  XOR U49977 ( .A(n38569), .B(n37053), .Z(n40330) );
  IV U49978 ( .A(n37054), .Z(n37056) );
  NOR U49979 ( .A(n37056), .B(n37055), .Z(n40328) );
  XOR U49980 ( .A(n40330), .B(n40328), .Z(n40333) );
  XOR U49981 ( .A(n40331), .B(n40333), .Z(n41850) );
  XOR U49982 ( .A(n37057), .B(n41850), .Z(n37058) );
  IV U49983 ( .A(n37058), .Z(n38563) );
  XOR U49984 ( .A(n38561), .B(n38563), .Z(n37065) );
  IV U49985 ( .A(n37065), .Z(n37059) );
  NOR U49986 ( .A(n37060), .B(n37059), .Z(n37062) );
  IV U49987 ( .A(n37060), .Z(n37061) );
  NOR U49988 ( .A(n38563), .B(n37061), .Z(n41837) );
  NOR U49989 ( .A(n37062), .B(n41837), .Z(n37063) );
  NOR U49990 ( .A(n37064), .B(n37063), .Z(n37067) );
  IV U49991 ( .A(n37064), .Z(n37066) );
  NOR U49992 ( .A(n37066), .B(n37065), .Z(n41834) );
  NOR U49993 ( .A(n37067), .B(n41834), .Z(n38555) );
  IV U49994 ( .A(n37068), .Z(n37070) );
  NOR U49995 ( .A(n37070), .B(n37069), .Z(n38558) );
  IV U49996 ( .A(n37071), .Z(n37078) );
  NOR U49997 ( .A(n37073), .B(n37072), .Z(n37074) );
  IV U49998 ( .A(n37074), .Z(n37075) );
  NOR U49999 ( .A(n37076), .B(n37075), .Z(n37077) );
  IV U50000 ( .A(n37077), .Z(n37081) );
  NOR U50001 ( .A(n37078), .B(n37081), .Z(n38556) );
  NOR U50002 ( .A(n38558), .B(n38556), .Z(n37079) );
  XOR U50003 ( .A(n38555), .B(n37079), .Z(n38554) );
  IV U50004 ( .A(n37080), .Z(n37082) );
  NOR U50005 ( .A(n37082), .B(n37081), .Z(n38552) );
  XOR U50006 ( .A(n38554), .B(n38552), .Z(n41825) );
  XOR U50007 ( .A(n38547), .B(n41825), .Z(n37083) );
  IV U50008 ( .A(n37083), .Z(n38549) );
  XOR U50009 ( .A(n38548), .B(n38549), .Z(n40340) );
  XOR U50010 ( .A(n40339), .B(n40340), .Z(n40343) );
  XOR U50011 ( .A(n40342), .B(n40343), .Z(n38543) );
  XOR U50012 ( .A(n38542), .B(n38543), .Z(n41820) );
  IV U50013 ( .A(n41820), .Z(n37091) );
  IV U50014 ( .A(n37084), .Z(n37088) );
  IV U50015 ( .A(n37087), .Z(n37085) );
  NOR U50016 ( .A(n37088), .B(n37085), .Z(n43792) );
  IV U50017 ( .A(n37086), .Z(n37090) );
  XOR U50018 ( .A(n37088), .B(n37087), .Z(n37089) );
  NOR U50019 ( .A(n37090), .B(n37089), .Z(n41818) );
  NOR U50020 ( .A(n43792), .B(n41818), .Z(n38545) );
  XOR U50021 ( .A(n37091), .B(n38545), .Z(n38541) );
  IV U50022 ( .A(n37092), .Z(n37093) );
  NOR U50023 ( .A(n37096), .B(n37093), .Z(n38537) );
  IV U50024 ( .A(n37094), .Z(n37095) );
  NOR U50025 ( .A(n37096), .B(n37095), .Z(n38539) );
  NOR U50026 ( .A(n38537), .B(n38539), .Z(n37097) );
  XOR U50027 ( .A(n38541), .B(n37097), .Z(n37098) );
  NOR U50028 ( .A(n37099), .B(n37098), .Z(n37102) );
  IV U50029 ( .A(n37099), .Z(n37101) );
  XOR U50030 ( .A(n38539), .B(n38541), .Z(n37100) );
  NOR U50031 ( .A(n37101), .B(n37100), .Z(n43804) );
  NOR U50032 ( .A(n37102), .B(n43804), .Z(n38534) );
  IV U50033 ( .A(n37103), .Z(n37105) );
  NOR U50034 ( .A(n37105), .B(n37104), .Z(n38535) );
  IV U50035 ( .A(n37106), .Z(n37113) );
  NOR U50036 ( .A(n37108), .B(n37107), .Z(n37109) );
  IV U50037 ( .A(n37109), .Z(n37110) );
  NOR U50038 ( .A(n37111), .B(n37110), .Z(n37112) );
  IV U50039 ( .A(n37112), .Z(n37116) );
  NOR U50040 ( .A(n37113), .B(n37116), .Z(n40349) );
  NOR U50041 ( .A(n38535), .B(n40349), .Z(n37114) );
  XOR U50042 ( .A(n38534), .B(n37114), .Z(n40354) );
  IV U50043 ( .A(n37115), .Z(n37117) );
  NOR U50044 ( .A(n37117), .B(n37116), .Z(n40352) );
  XOR U50045 ( .A(n40354), .B(n40352), .Z(n40357) );
  XOR U50046 ( .A(n40355), .B(n40357), .Z(n40361) );
  XOR U50047 ( .A(n40360), .B(n40361), .Z(n40364) );
  XOR U50048 ( .A(n40363), .B(n40364), .Z(n40368) );
  XOR U50049 ( .A(n40367), .B(n40368), .Z(n40375) );
  XOR U50050 ( .A(n37118), .B(n40375), .Z(n37119) );
  IV U50051 ( .A(n37119), .Z(n38529) );
  XOR U50052 ( .A(n38528), .B(n38529), .Z(n38532) );
  XOR U50053 ( .A(n38531), .B(n38532), .Z(n38523) );
  XOR U50054 ( .A(n38522), .B(n38523), .Z(n38527) );
  IV U50055 ( .A(n37120), .Z(n37122) );
  NOR U50056 ( .A(n37122), .B(n37121), .Z(n38525) );
  XOR U50057 ( .A(n38527), .B(n38525), .Z(n40392) );
  XOR U50058 ( .A(n40391), .B(n40392), .Z(n38520) );
  IV U50059 ( .A(n37123), .Z(n37125) );
  NOR U50060 ( .A(n37125), .B(n37124), .Z(n38518) );
  XOR U50061 ( .A(n38520), .B(n38518), .Z(n40389) );
  IV U50062 ( .A(n37126), .Z(n37127) );
  NOR U50063 ( .A(n37128), .B(n37127), .Z(n40387) );
  XOR U50064 ( .A(n40389), .B(n40387), .Z(n38513) );
  XOR U50065 ( .A(n38512), .B(n38513), .Z(n38516) );
  XOR U50066 ( .A(n38515), .B(n38516), .Z(n40401) );
  IV U50067 ( .A(n37129), .Z(n37130) );
  NOR U50068 ( .A(n37131), .B(n37130), .Z(n40400) );
  IV U50069 ( .A(n37132), .Z(n37134) );
  NOR U50070 ( .A(n37134), .B(n37133), .Z(n38510) );
  NOR U50071 ( .A(n40400), .B(n38510), .Z(n37135) );
  XOR U50072 ( .A(n40401), .B(n37135), .Z(n40404) );
  IV U50073 ( .A(n37136), .Z(n37138) );
  NOR U50074 ( .A(n37138), .B(n37137), .Z(n40403) );
  IV U50075 ( .A(n37139), .Z(n37141) );
  NOR U50076 ( .A(n37141), .B(n37140), .Z(n40408) );
  NOR U50077 ( .A(n40403), .B(n40408), .Z(n37142) );
  XOR U50078 ( .A(n40404), .B(n37142), .Z(n38507) );
  XOR U50079 ( .A(n38505), .B(n38507), .Z(n40413) );
  IV U50080 ( .A(n40413), .Z(n37150) );
  IV U50081 ( .A(n37143), .Z(n37144) );
  NOR U50082 ( .A(n37145), .B(n37144), .Z(n38508) );
  IV U50083 ( .A(n37146), .Z(n37148) );
  NOR U50084 ( .A(n37148), .B(n37147), .Z(n40412) );
  NOR U50085 ( .A(n38508), .B(n40412), .Z(n37149) );
  XOR U50086 ( .A(n37150), .B(n37149), .Z(n40416) );
  XOR U50087 ( .A(n40415), .B(n40416), .Z(n38503) );
  XOR U50088 ( .A(n37151), .B(n38503), .Z(n38495) );
  IV U50089 ( .A(n37152), .Z(n37154) );
  NOR U50090 ( .A(n37154), .B(n37153), .Z(n38497) );
  IV U50091 ( .A(n37155), .Z(n37157) );
  NOR U50092 ( .A(n37157), .B(n37156), .Z(n38494) );
  NOR U50093 ( .A(n38497), .B(n38494), .Z(n37158) );
  XOR U50094 ( .A(n38495), .B(n37158), .Z(n41775) );
  XOR U50095 ( .A(n40419), .B(n41775), .Z(n40432) );
  NOR U50096 ( .A(n37159), .B(n38488), .Z(n37163) );
  IV U50097 ( .A(n37160), .Z(n37162) );
  NOR U50098 ( .A(n37162), .B(n37161), .Z(n38491) );
  NOR U50099 ( .A(n37163), .B(n38491), .Z(n37164) );
  XOR U50100 ( .A(n40432), .B(n37164), .Z(n40437) );
  XOR U50101 ( .A(n37165), .B(n40437), .Z(n37166) );
  IV U50102 ( .A(n37166), .Z(n40441) );
  XOR U50103 ( .A(n40439), .B(n40441), .Z(n40443) );
  IV U50104 ( .A(n37167), .Z(n37169) );
  NOR U50105 ( .A(n37169), .B(n37168), .Z(n37170) );
  IV U50106 ( .A(n37170), .Z(n40442) );
  XOR U50107 ( .A(n40443), .B(n40442), .Z(n37171) );
  NOR U50108 ( .A(n37172), .B(n37171), .Z(n38485) );
  IV U50109 ( .A(n37172), .Z(n37173) );
  NOR U50110 ( .A(n37173), .B(n40443), .Z(n47303) );
  NOR U50111 ( .A(n38485), .B(n47303), .Z(n37174) );
  IV U50112 ( .A(n37174), .Z(n38481) );
  IV U50113 ( .A(n37175), .Z(n37176) );
  NOR U50114 ( .A(n37177), .B(n37176), .Z(n38480) );
  IV U50115 ( .A(n37178), .Z(n37180) );
  NOR U50116 ( .A(n37180), .B(n37179), .Z(n38483) );
  NOR U50117 ( .A(n38480), .B(n38483), .Z(n37181) );
  XOR U50118 ( .A(n38481), .B(n37181), .Z(n40445) );
  IV U50119 ( .A(n37182), .Z(n37184) );
  NOR U50120 ( .A(n37184), .B(n37183), .Z(n43874) );
  IV U50121 ( .A(n37185), .Z(n37187) );
  NOR U50122 ( .A(n37187), .B(n37186), .Z(n41760) );
  NOR U50123 ( .A(n43874), .B(n41760), .Z(n40446) );
  XOR U50124 ( .A(n40445), .B(n40446), .Z(n40448) );
  XOR U50125 ( .A(n40447), .B(n40448), .Z(n40454) );
  IV U50126 ( .A(n37188), .Z(n37190) );
  NOR U50127 ( .A(n37190), .B(n37189), .Z(n40452) );
  XOR U50128 ( .A(n40454), .B(n40452), .Z(n40456) );
  XOR U50129 ( .A(n40455), .B(n40456), .Z(n40460) );
  XOR U50130 ( .A(n40459), .B(n40460), .Z(n40463) );
  XOR U50131 ( .A(n40462), .B(n40463), .Z(n38477) );
  XOR U50132 ( .A(n38476), .B(n38477), .Z(n40467) );
  XOR U50133 ( .A(n40466), .B(n40467), .Z(n40471) );
  IV U50134 ( .A(n37191), .Z(n37193) );
  NOR U50135 ( .A(n37193), .B(n37192), .Z(n40469) );
  XOR U50136 ( .A(n40471), .B(n40469), .Z(n38471) );
  XOR U50137 ( .A(n38470), .B(n38471), .Z(n38475) );
  IV U50138 ( .A(n37194), .Z(n37196) );
  NOR U50139 ( .A(n37196), .B(n37195), .Z(n38473) );
  XOR U50140 ( .A(n38475), .B(n38473), .Z(n38466) );
  XOR U50141 ( .A(n38465), .B(n38466), .Z(n43885) );
  IV U50142 ( .A(n43885), .Z(n37203) );
  IV U50143 ( .A(n37197), .Z(n37198) );
  NOR U50144 ( .A(n37199), .B(n37198), .Z(n43883) );
  IV U50145 ( .A(n37200), .Z(n37201) );
  NOR U50146 ( .A(n37202), .B(n37201), .Z(n43892) );
  NOR U50147 ( .A(n43883), .B(n43892), .Z(n38468) );
  XOR U50148 ( .A(n37203), .B(n38468), .Z(n38460) );
  XOR U50149 ( .A(n38459), .B(n38460), .Z(n38463) );
  XOR U50150 ( .A(n38462), .B(n38463), .Z(n38455) );
  XOR U50151 ( .A(n38453), .B(n38455), .Z(n38458) );
  XOR U50152 ( .A(n38456), .B(n38458), .Z(n38452) );
  XOR U50153 ( .A(n38450), .B(n38452), .Z(n40480) );
  XOR U50154 ( .A(n40478), .B(n40480), .Z(n40482) );
  XOR U50155 ( .A(n37204), .B(n40482), .Z(n37205) );
  IV U50156 ( .A(n37205), .Z(n38447) );
  XOR U50157 ( .A(n38445), .B(n38447), .Z(n40490) );
  XOR U50158 ( .A(n40489), .B(n40490), .Z(n40487) );
  IV U50159 ( .A(n37206), .Z(n37208) );
  IV U50160 ( .A(n37207), .Z(n37211) );
  NOR U50161 ( .A(n37208), .B(n37211), .Z(n40485) );
  XOR U50162 ( .A(n40487), .B(n40485), .Z(n38443) );
  NOR U50163 ( .A(n37209), .B(n38443), .Z(n41722) );
  IV U50164 ( .A(n37210), .Z(n37212) );
  NOR U50165 ( .A(n37212), .B(n37211), .Z(n38442) );
  XOR U50166 ( .A(n38442), .B(n38443), .Z(n37218) );
  IV U50167 ( .A(n37218), .Z(n37213) );
  NOR U50168 ( .A(n37214), .B(n37213), .Z(n37215) );
  NOR U50169 ( .A(n41722), .B(n37215), .Z(n37216) );
  NOR U50170 ( .A(n37217), .B(n37216), .Z(n37220) );
  IV U50171 ( .A(n37217), .Z(n37219) );
  NOR U50172 ( .A(n37219), .B(n37218), .Z(n41720) );
  NOR U50173 ( .A(n37220), .B(n41720), .Z(n38440) );
  XOR U50174 ( .A(n40501), .B(n38440), .Z(n38438) );
  XOR U50175 ( .A(n37221), .B(n38438), .Z(n37222) );
  IV U50176 ( .A(n37222), .Z(n38434) );
  XOR U50177 ( .A(n38432), .B(n38434), .Z(n41711) );
  XOR U50178 ( .A(n41698), .B(n41711), .Z(n40506) );
  XOR U50179 ( .A(n40507), .B(n40506), .Z(n37223) );
  IV U50180 ( .A(n37223), .Z(n40509) );
  XOR U50181 ( .A(n40508), .B(n40509), .Z(n40521) );
  IV U50182 ( .A(n37224), .Z(n37226) );
  NOR U50183 ( .A(n37226), .B(n37225), .Z(n40519) );
  NOR U50184 ( .A(n38430), .B(n40519), .Z(n37227) );
  XOR U50185 ( .A(n40521), .B(n37227), .Z(n38427) );
  IV U50186 ( .A(n37228), .Z(n40515) );
  NOR U50187 ( .A(n40515), .B(n37229), .Z(n37233) );
  IV U50188 ( .A(n37230), .Z(n37232) );
  NOR U50189 ( .A(n37232), .B(n37231), .Z(n38424) );
  NOR U50190 ( .A(n37233), .B(n38424), .Z(n37234) );
  XOR U50191 ( .A(n38427), .B(n37234), .Z(n40533) );
  XOR U50192 ( .A(n37235), .B(n40533), .Z(n37236) );
  IV U50193 ( .A(n37236), .Z(n40540) );
  XOR U50194 ( .A(n37237), .B(n40540), .Z(n40547) );
  XOR U50195 ( .A(n37238), .B(n40547), .Z(n37239) );
  IV U50196 ( .A(n37239), .Z(n40551) );
  XOR U50197 ( .A(n40549), .B(n40551), .Z(n40554) );
  IV U50198 ( .A(n37240), .Z(n37241) );
  NOR U50199 ( .A(n37242), .B(n37241), .Z(n37243) );
  IV U50200 ( .A(n37243), .Z(n37244) );
  NOR U50201 ( .A(n37245), .B(n37244), .Z(n40552) );
  XOR U50202 ( .A(n40554), .B(n40552), .Z(n40561) );
  XOR U50203 ( .A(n38422), .B(n40561), .Z(n37246) );
  XOR U50204 ( .A(n37247), .B(n37246), .Z(n40571) );
  NOR U50205 ( .A(n37249), .B(n37248), .Z(n40557) );
  IV U50206 ( .A(n37250), .Z(n37251) );
  NOR U50207 ( .A(n37252), .B(n37251), .Z(n40569) );
  NOR U50208 ( .A(n40557), .B(n40569), .Z(n37253) );
  XOR U50209 ( .A(n40571), .B(n37253), .Z(n38418) );
  IV U50210 ( .A(n37254), .Z(n37256) );
  NOR U50211 ( .A(n37256), .B(n37255), .Z(n40565) );
  IV U50212 ( .A(n37257), .Z(n37258) );
  NOR U50213 ( .A(n37262), .B(n37258), .Z(n38417) );
  NOR U50214 ( .A(n40565), .B(n38417), .Z(n37259) );
  XOR U50215 ( .A(n38418), .B(n37259), .Z(n38416) );
  IV U50216 ( .A(n37260), .Z(n37261) );
  NOR U50217 ( .A(n37262), .B(n37261), .Z(n38414) );
  XOR U50218 ( .A(n38416), .B(n38414), .Z(n43963) );
  XOR U50219 ( .A(n38409), .B(n43963), .Z(n38410) );
  IV U50220 ( .A(n37263), .Z(n37265) );
  NOR U50221 ( .A(n37265), .B(n37264), .Z(n38411) );
  IV U50222 ( .A(n37266), .Z(n37272) );
  IV U50223 ( .A(n37267), .Z(n37268) );
  NOR U50224 ( .A(n37272), .B(n37268), .Z(n40583) );
  NOR U50225 ( .A(n38411), .B(n40583), .Z(n37269) );
  XOR U50226 ( .A(n38410), .B(n37269), .Z(n38407) );
  IV U50227 ( .A(n37270), .Z(n37271) );
  NOR U50228 ( .A(n37272), .B(n37271), .Z(n38405) );
  XOR U50229 ( .A(n38407), .B(n38405), .Z(n40580) );
  XOR U50230 ( .A(n37273), .B(n40580), .Z(n38398) );
  IV U50231 ( .A(n37274), .Z(n37276) );
  NOR U50232 ( .A(n37276), .B(n37275), .Z(n38397) );
  IV U50233 ( .A(n37277), .Z(n37279) );
  NOR U50234 ( .A(n37279), .B(n37278), .Z(n37280) );
  IV U50235 ( .A(n37280), .Z(n37281) );
  NOR U50236 ( .A(n37282), .B(n37281), .Z(n38402) );
  NOR U50237 ( .A(n38397), .B(n38402), .Z(n37283) );
  XOR U50238 ( .A(n38398), .B(n37283), .Z(n40595) );
  XOR U50239 ( .A(n40594), .B(n40595), .Z(n40599) );
  XOR U50240 ( .A(n40597), .B(n40599), .Z(n40602) );
  XOR U50241 ( .A(n40601), .B(n40602), .Z(n40605) );
  NOR U50242 ( .A(n37287), .B(n40605), .Z(n43982) );
  IV U50243 ( .A(n37284), .Z(n37286) );
  NOR U50244 ( .A(n37286), .B(n37285), .Z(n37288) );
  IV U50245 ( .A(n37288), .Z(n40604) );
  XOR U50246 ( .A(n40605), .B(n40604), .Z(n37290) );
  NOR U50247 ( .A(n37288), .B(n37287), .Z(n37289) );
  NOR U50248 ( .A(n37290), .B(n37289), .Z(n40608) );
  NOR U50249 ( .A(n43982), .B(n40608), .Z(n38392) );
  XOR U50250 ( .A(n37291), .B(n38392), .Z(n37295) );
  IV U50251 ( .A(n37295), .Z(n37292) );
  NOR U50252 ( .A(n37293), .B(n37292), .Z(n38391) );
  IV U50253 ( .A(n37293), .Z(n37294) );
  NOR U50254 ( .A(n37295), .B(n37294), .Z(n43993) );
  NOR U50255 ( .A(n38391), .B(n43993), .Z(n38386) );
  IV U50256 ( .A(n37296), .Z(n37300) );
  NOR U50257 ( .A(n37298), .B(n37297), .Z(n37299) );
  IV U50258 ( .A(n37299), .Z(n37303) );
  NOR U50259 ( .A(n37300), .B(n37303), .Z(n38387) );
  NOR U50260 ( .A(n38389), .B(n38387), .Z(n37301) );
  XOR U50261 ( .A(n38386), .B(n37301), .Z(n38382) );
  IV U50262 ( .A(n37302), .Z(n37304) );
  NOR U50263 ( .A(n37304), .B(n37303), .Z(n38380) );
  XOR U50264 ( .A(n38382), .B(n38380), .Z(n38384) );
  XOR U50265 ( .A(n38383), .B(n38384), .Z(n41610) );
  XOR U50266 ( .A(n40612), .B(n41610), .Z(n38378) );
  IV U50267 ( .A(n37305), .Z(n37306) );
  NOR U50268 ( .A(n37307), .B(n37306), .Z(n40613) );
  IV U50269 ( .A(n37308), .Z(n37309) );
  NOR U50270 ( .A(n37310), .B(n37309), .Z(n38377) );
  NOR U50271 ( .A(n40613), .B(n38377), .Z(n37311) );
  XOR U50272 ( .A(n38378), .B(n37311), .Z(n38376) );
  IV U50273 ( .A(n38376), .Z(n37319) );
  IV U50274 ( .A(n37312), .Z(n37314) );
  NOR U50275 ( .A(n37314), .B(n37313), .Z(n38374) );
  IV U50276 ( .A(n37315), .Z(n37317) );
  NOR U50277 ( .A(n37317), .B(n37316), .Z(n38372) );
  NOR U50278 ( .A(n38374), .B(n38372), .Z(n37318) );
  XOR U50279 ( .A(n37319), .B(n37318), .Z(n40621) );
  XOR U50280 ( .A(n38367), .B(n40621), .Z(n38370) );
  IV U50281 ( .A(n38370), .Z(n37327) );
  IV U50282 ( .A(n37320), .Z(n37322) );
  NOR U50283 ( .A(n37322), .B(n37321), .Z(n38369) );
  IV U50284 ( .A(n37323), .Z(n37325) );
  NOR U50285 ( .A(n37325), .B(n37324), .Z(n40620) );
  NOR U50286 ( .A(n38369), .B(n40620), .Z(n37326) );
  XOR U50287 ( .A(n37327), .B(n37326), .Z(n40619) );
  XOR U50288 ( .A(n40618), .B(n40619), .Z(n37334) );
  IV U50289 ( .A(n37334), .Z(n37328) );
  NOR U50290 ( .A(n37329), .B(n37328), .Z(n52080) );
  IV U50291 ( .A(n37330), .Z(n37331) );
  NOR U50292 ( .A(n37332), .B(n37331), .Z(n37335) );
  IV U50293 ( .A(n37335), .Z(n37333) );
  NOR U50294 ( .A(n40619), .B(n37333), .Z(n44009) );
  NOR U50295 ( .A(n37335), .B(n37334), .Z(n37336) );
  NOR U50296 ( .A(n44009), .B(n37336), .Z(n37337) );
  NOR U50297 ( .A(n37338), .B(n37337), .Z(n37339) );
  NOR U50298 ( .A(n52080), .B(n37339), .Z(n38362) );
  XOR U50299 ( .A(n40626), .B(n38362), .Z(n38356) );
  XOR U50300 ( .A(n38355), .B(n38356), .Z(n38360) );
  XOR U50301 ( .A(n38358), .B(n38360), .Z(n40637) );
  XOR U50302 ( .A(n40635), .B(n40637), .Z(n38353) );
  IV U50303 ( .A(n37340), .Z(n37341) );
  NOR U50304 ( .A(n37342), .B(n37341), .Z(n37343) );
  IV U50305 ( .A(n37343), .Z(n37349) );
  NOR U50306 ( .A(n38353), .B(n37349), .Z(n41592) );
  IV U50307 ( .A(n37344), .Z(n37345) );
  NOR U50308 ( .A(n37345), .B(n37347), .Z(n38351) );
  XOR U50309 ( .A(n38353), .B(n38351), .Z(n40633) );
  IV U50310 ( .A(n37346), .Z(n37348) );
  NOR U50311 ( .A(n37348), .B(n37347), .Z(n37350) );
  IV U50312 ( .A(n37350), .Z(n40632) );
  XOR U50313 ( .A(n40633), .B(n40632), .Z(n37352) );
  NOR U50314 ( .A(n37350), .B(n37349), .Z(n37351) );
  NOR U50315 ( .A(n37352), .B(n37351), .Z(n37353) );
  NOR U50316 ( .A(n41592), .B(n37353), .Z(n38344) );
  XOR U50317 ( .A(n37354), .B(n38344), .Z(n40646) );
  XOR U50318 ( .A(n40644), .B(n40646), .Z(n38338) );
  XOR U50319 ( .A(n38337), .B(n38338), .Z(n38342) );
  IV U50320 ( .A(n37355), .Z(n37356) );
  NOR U50321 ( .A(n37357), .B(n37356), .Z(n38340) );
  XOR U50322 ( .A(n38342), .B(n38340), .Z(n38332) );
  XOR U50323 ( .A(n38331), .B(n38332), .Z(n38335) );
  XOR U50324 ( .A(n38334), .B(n38335), .Z(n44044) );
  IV U50325 ( .A(n37358), .Z(n37359) );
  NOR U50326 ( .A(n37360), .B(n37359), .Z(n40653) );
  NOR U50327 ( .A(n40658), .B(n40653), .Z(n37361) );
  XOR U50328 ( .A(n44044), .B(n37361), .Z(n40655) );
  XOR U50329 ( .A(n37362), .B(n40655), .Z(n38329) );
  IV U50330 ( .A(n37363), .Z(n37364) );
  NOR U50331 ( .A(n37365), .B(n37364), .Z(n38328) );
  IV U50332 ( .A(n37366), .Z(n37368) );
  NOR U50333 ( .A(n37368), .B(n37367), .Z(n38326) );
  NOR U50334 ( .A(n38328), .B(n38326), .Z(n37369) );
  XOR U50335 ( .A(n38329), .B(n37369), .Z(n38314) );
  XOR U50336 ( .A(n37370), .B(n38314), .Z(n38313) );
  XOR U50337 ( .A(n38311), .B(n38313), .Z(n38306) );
  XOR U50338 ( .A(n38305), .B(n38306), .Z(n38310) );
  IV U50339 ( .A(n37371), .Z(n37373) );
  NOR U50340 ( .A(n37373), .B(n37372), .Z(n38308) );
  XOR U50341 ( .A(n38310), .B(n38308), .Z(n38300) );
  XOR U50342 ( .A(n38301), .B(n38300), .Z(n38303) );
  IV U50343 ( .A(n37374), .Z(n37376) );
  IV U50344 ( .A(n37375), .Z(n37382) );
  NOR U50345 ( .A(n37376), .B(n37382), .Z(n40668) );
  NOR U50346 ( .A(n38302), .B(n40668), .Z(n37377) );
  XOR U50347 ( .A(n38303), .B(n37377), .Z(n41567) );
  IV U50348 ( .A(n37378), .Z(n37379) );
  NOR U50349 ( .A(n37380), .B(n37379), .Z(n37387) );
  IV U50350 ( .A(n37387), .Z(n37381) );
  NOR U50351 ( .A(n41567), .B(n37381), .Z(n44080) );
  NOR U50352 ( .A(n37383), .B(n37382), .Z(n37384) );
  IV U50353 ( .A(n37384), .Z(n41569) );
  NOR U50354 ( .A(n37385), .B(n41569), .Z(n38298) );
  XOR U50355 ( .A(n38298), .B(n41567), .Z(n40680) );
  IV U50356 ( .A(n40680), .Z(n37386) );
  NOR U50357 ( .A(n37387), .B(n37386), .Z(n37388) );
  NOR U50358 ( .A(n44080), .B(n37388), .Z(n40684) );
  IV U50359 ( .A(n37389), .Z(n37390) );
  NOR U50360 ( .A(n37391), .B(n37390), .Z(n40679) );
  IV U50361 ( .A(n37392), .Z(n37393) );
  NOR U50362 ( .A(n37396), .B(n37393), .Z(n40685) );
  NOR U50363 ( .A(n40679), .B(n40685), .Z(n37394) );
  XOR U50364 ( .A(n40684), .B(n37394), .Z(n40690) );
  IV U50365 ( .A(n37395), .Z(n37397) );
  NOR U50366 ( .A(n37397), .B(n37396), .Z(n40688) );
  XOR U50367 ( .A(n40690), .B(n40688), .Z(n40692) );
  XOR U50368 ( .A(n40691), .B(n40692), .Z(n37403) );
  XOR U50369 ( .A(n37398), .B(n37403), .Z(n37405) );
  NOR U50370 ( .A(n37399), .B(n37405), .Z(n44092) );
  IV U50371 ( .A(n37400), .Z(n37402) );
  NOR U50372 ( .A(n37402), .B(n37401), .Z(n37407) );
  IV U50373 ( .A(n37407), .Z(n37404) );
  NOR U50374 ( .A(n37404), .B(n37403), .Z(n41552) );
  IV U50375 ( .A(n37405), .Z(n37406) );
  NOR U50376 ( .A(n37407), .B(n37406), .Z(n37408) );
  NOR U50377 ( .A(n41552), .B(n37408), .Z(n37413) );
  NOR U50378 ( .A(n37409), .B(n37413), .Z(n37410) );
  NOR U50379 ( .A(n44092), .B(n37410), .Z(n37411) );
  NOR U50380 ( .A(n37412), .B(n37411), .Z(n37416) );
  IV U50381 ( .A(n37412), .Z(n37415) );
  IV U50382 ( .A(n37413), .Z(n37414) );
  NOR U50383 ( .A(n37415), .B(n37414), .Z(n38289) );
  NOR U50384 ( .A(n37416), .B(n38289), .Z(n38287) );
  XOR U50385 ( .A(n37417), .B(n38287), .Z(n40701) );
  XOR U50386 ( .A(n40699), .B(n40701), .Z(n40707) );
  IV U50387 ( .A(n37418), .Z(n37419) );
  NOR U50388 ( .A(n37420), .B(n37419), .Z(n38284) );
  IV U50389 ( .A(n37421), .Z(n37423) );
  NOR U50390 ( .A(n37423), .B(n37422), .Z(n40706) );
  NOR U50391 ( .A(n38284), .B(n40706), .Z(n37424) );
  XOR U50392 ( .A(n40707), .B(n37424), .Z(n38282) );
  XOR U50393 ( .A(n38283), .B(n38282), .Z(n38278) );
  IV U50394 ( .A(n37425), .Z(n37427) );
  NOR U50395 ( .A(n37427), .B(n37426), .Z(n38276) );
  XOR U50396 ( .A(n38278), .B(n38276), .Z(n38280) );
  XOR U50397 ( .A(n38279), .B(n38280), .Z(n41539) );
  IV U50398 ( .A(n37428), .Z(n37429) );
  NOR U50399 ( .A(n37430), .B(n37429), .Z(n44112) );
  IV U50400 ( .A(n37431), .Z(n37432) );
  NOR U50401 ( .A(n37433), .B(n37432), .Z(n41538) );
  NOR U50402 ( .A(n44112), .B(n41538), .Z(n40725) );
  XOR U50403 ( .A(n41539), .B(n40725), .Z(n37436) );
  IV U50404 ( .A(n37436), .Z(n37434) );
  NOR U50405 ( .A(n37435), .B(n37434), .Z(n41542) );
  NOR U50406 ( .A(n37437), .B(n37436), .Z(n40724) );
  NOR U50407 ( .A(n41542), .B(n40724), .Z(n40732) );
  IV U50408 ( .A(n37438), .Z(n37439) );
  NOR U50409 ( .A(n37440), .B(n37439), .Z(n40722) );
  IV U50410 ( .A(n37441), .Z(n37442) );
  NOR U50411 ( .A(n37443), .B(n37442), .Z(n40731) );
  NOR U50412 ( .A(n40722), .B(n40731), .Z(n37444) );
  XOR U50413 ( .A(n40732), .B(n37444), .Z(n38275) );
  IV U50414 ( .A(n38275), .Z(n37452) );
  IV U50415 ( .A(n37445), .Z(n37446) );
  NOR U50416 ( .A(n37447), .B(n37446), .Z(n38273) );
  IV U50417 ( .A(n37448), .Z(n37450) );
  NOR U50418 ( .A(n37450), .B(n37449), .Z(n38271) );
  NOR U50419 ( .A(n38273), .B(n38271), .Z(n37451) );
  XOR U50420 ( .A(n37452), .B(n37451), .Z(n40738) );
  IV U50421 ( .A(n37453), .Z(n37454) );
  NOR U50422 ( .A(n37454), .B(n37457), .Z(n40736) );
  XOR U50423 ( .A(n40738), .B(n40736), .Z(n38269) );
  IV U50424 ( .A(n37455), .Z(n37456) );
  NOR U50425 ( .A(n37457), .B(n37456), .Z(n38267) );
  XOR U50426 ( .A(n38269), .B(n38267), .Z(n40750) );
  XOR U50427 ( .A(n40749), .B(n40750), .Z(n38266) );
  IV U50428 ( .A(n37458), .Z(n37466) );
  IV U50429 ( .A(n37459), .Z(n37461) );
  NOR U50430 ( .A(n37461), .B(n37460), .Z(n37462) );
  IV U50431 ( .A(n37462), .Z(n37463) );
  NOR U50432 ( .A(n37464), .B(n37463), .Z(n37465) );
  IV U50433 ( .A(n37465), .Z(n37468) );
  NOR U50434 ( .A(n37466), .B(n37468), .Z(n38264) );
  XOR U50435 ( .A(n38266), .B(n38264), .Z(n38263) );
  IV U50436 ( .A(n37467), .Z(n37469) );
  NOR U50437 ( .A(n37469), .B(n37468), .Z(n38261) );
  XOR U50438 ( .A(n38263), .B(n38261), .Z(n40761) );
  XOR U50439 ( .A(n40760), .B(n40761), .Z(n40765) );
  IV U50440 ( .A(n37470), .Z(n37472) );
  NOR U50441 ( .A(n37472), .B(n37471), .Z(n40763) );
  XOR U50442 ( .A(n40765), .B(n40763), .Z(n40768) );
  XOR U50443 ( .A(n40767), .B(n40768), .Z(n40771) );
  XOR U50444 ( .A(n40770), .B(n40771), .Z(n40775) );
  IV U50445 ( .A(n37473), .Z(n37475) );
  IV U50446 ( .A(n37474), .Z(n37478) );
  NOR U50447 ( .A(n37475), .B(n37478), .Z(n37476) );
  IV U50448 ( .A(n37476), .Z(n40774) );
  XOR U50449 ( .A(n40775), .B(n40774), .Z(n38257) );
  IV U50450 ( .A(n37477), .Z(n37479) );
  NOR U50451 ( .A(n37479), .B(n37478), .Z(n40776) );
  IV U50452 ( .A(n37480), .Z(n37481) );
  NOR U50453 ( .A(n37485), .B(n37481), .Z(n38258) );
  NOR U50454 ( .A(n40776), .B(n38258), .Z(n37482) );
  XOR U50455 ( .A(n38257), .B(n37482), .Z(n38253) );
  IV U50456 ( .A(n37483), .Z(n37484) );
  NOR U50457 ( .A(n37485), .B(n37484), .Z(n38251) );
  XOR U50458 ( .A(n38253), .B(n38251), .Z(n38255) );
  NOR U50459 ( .A(n37491), .B(n38255), .Z(n41518) );
  IV U50460 ( .A(n37486), .Z(n37488) );
  NOR U50461 ( .A(n37488), .B(n37487), .Z(n38254) );
  XOR U50462 ( .A(n38254), .B(n38255), .Z(n38250) );
  IV U50463 ( .A(n37489), .Z(n37490) );
  NOR U50464 ( .A(n37490), .B(n37496), .Z(n37492) );
  IV U50465 ( .A(n37492), .Z(n38249) );
  XOR U50466 ( .A(n38250), .B(n38249), .Z(n37494) );
  NOR U50467 ( .A(n37492), .B(n37491), .Z(n37493) );
  NOR U50468 ( .A(n37494), .B(n37493), .Z(n37495) );
  NOR U50469 ( .A(n41518), .B(n37495), .Z(n38246) );
  NOR U50470 ( .A(n37497), .B(n37496), .Z(n37498) );
  IV U50471 ( .A(n37498), .Z(n37499) );
  NOR U50472 ( .A(n37500), .B(n37499), .Z(n37501) );
  IV U50473 ( .A(n37501), .Z(n38247) );
  XOR U50474 ( .A(n38246), .B(n38247), .Z(n40783) );
  IV U50475 ( .A(n37502), .Z(n37504) );
  NOR U50476 ( .A(n37504), .B(n37503), .Z(n40781) );
  XOR U50477 ( .A(n40783), .B(n40781), .Z(n40785) );
  XOR U50478 ( .A(n40784), .B(n40785), .Z(n40793) );
  IV U50479 ( .A(n40793), .Z(n37511) );
  IV U50480 ( .A(n37505), .Z(n37506) );
  NOR U50481 ( .A(n37507), .B(n37506), .Z(n40792) );
  NOR U50482 ( .A(n37509), .B(n37508), .Z(n40790) );
  NOR U50483 ( .A(n40792), .B(n40790), .Z(n37510) );
  XOR U50484 ( .A(n37511), .B(n37510), .Z(n44168) );
  XOR U50485 ( .A(n40788), .B(n44168), .Z(n40803) );
  XOR U50486 ( .A(n37512), .B(n40803), .Z(n37513) );
  IV U50487 ( .A(n37513), .Z(n40801) );
  XOR U50488 ( .A(n40799), .B(n40801), .Z(n44186) );
  IV U50489 ( .A(n37514), .Z(n44184) );
  IV U50490 ( .A(n37515), .Z(n37516) );
  NOR U50491 ( .A(n44184), .B(n37516), .Z(n38239) );
  IV U50492 ( .A(n37517), .Z(n37518) );
  NOR U50493 ( .A(n44184), .B(n37518), .Z(n44187) );
  NOR U50494 ( .A(n38239), .B(n44187), .Z(n37519) );
  XOR U50495 ( .A(n44186), .B(n37519), .Z(n38236) );
  XOR U50496 ( .A(n37520), .B(n38236), .Z(n40810) );
  XOR U50497 ( .A(n40809), .B(n40810), .Z(n40817) );
  XOR U50498 ( .A(n40812), .B(n40817), .Z(n38235) );
  IV U50499 ( .A(n37521), .Z(n37523) );
  NOR U50500 ( .A(n37523), .B(n37522), .Z(n40816) );
  IV U50501 ( .A(n37538), .Z(n37525) );
  NOR U50502 ( .A(n37525), .B(n37524), .Z(n37526) );
  IV U50503 ( .A(n37526), .Z(n37530) );
  NOR U50504 ( .A(n37541), .B(n37527), .Z(n37528) );
  IV U50505 ( .A(n37528), .Z(n37529) );
  NOR U50506 ( .A(n37530), .B(n37529), .Z(n38233) );
  NOR U50507 ( .A(n40816), .B(n38233), .Z(n37531) );
  XOR U50508 ( .A(n38235), .B(n37531), .Z(n38227) );
  IV U50509 ( .A(n37532), .Z(n37533) );
  NOR U50510 ( .A(n37533), .B(n37541), .Z(n38228) );
  IV U50511 ( .A(n37534), .Z(n37535) );
  NOR U50512 ( .A(n37535), .B(n37541), .Z(n37536) );
  IV U50513 ( .A(n37536), .Z(n37537) );
  NOR U50514 ( .A(n37538), .B(n37537), .Z(n38230) );
  NOR U50515 ( .A(n38228), .B(n38230), .Z(n37539) );
  XOR U50516 ( .A(n38227), .B(n37539), .Z(n38226) );
  IV U50517 ( .A(n37540), .Z(n37544) );
  NOR U50518 ( .A(n37542), .B(n37541), .Z(n37543) );
  IV U50519 ( .A(n37543), .Z(n37546) );
  NOR U50520 ( .A(n37544), .B(n37546), .Z(n38224) );
  XOR U50521 ( .A(n38226), .B(n38224), .Z(n38220) );
  IV U50522 ( .A(n37545), .Z(n37547) );
  NOR U50523 ( .A(n37547), .B(n37546), .Z(n38218) );
  XOR U50524 ( .A(n38220), .B(n38218), .Z(n38223) );
  IV U50525 ( .A(n38223), .Z(n37555) );
  IV U50526 ( .A(n37548), .Z(n37550) );
  NOR U50527 ( .A(n37550), .B(n37549), .Z(n38216) );
  IV U50528 ( .A(n37551), .Z(n37552) );
  NOR U50529 ( .A(n37553), .B(n37552), .Z(n38221) );
  NOR U50530 ( .A(n38216), .B(n38221), .Z(n37554) );
  XOR U50531 ( .A(n37555), .B(n37554), .Z(n40823) );
  XOR U50532 ( .A(n40821), .B(n40823), .Z(n40825) );
  XOR U50533 ( .A(n37556), .B(n40825), .Z(n38210) );
  XOR U50534 ( .A(n38211), .B(n38210), .Z(n38206) );
  XOR U50535 ( .A(n38204), .B(n38206), .Z(n38209) );
  XOR U50536 ( .A(n37557), .B(n38209), .Z(n41474) );
  XOR U50537 ( .A(n37558), .B(n41474), .Z(n38196) );
  XOR U50538 ( .A(n37559), .B(n38196), .Z(n38178) );
  XOR U50539 ( .A(n37560), .B(n38178), .Z(n38176) );
  XOR U50540 ( .A(n38175), .B(n38176), .Z(n38171) );
  XOR U50541 ( .A(n38169), .B(n38171), .Z(n38173) );
  XOR U50542 ( .A(n38172), .B(n38173), .Z(n38167) );
  XOR U50543 ( .A(n38165), .B(n38167), .Z(n40843) );
  XOR U50544 ( .A(n40842), .B(n40843), .Z(n40859) );
  XOR U50545 ( .A(n37561), .B(n40859), .Z(n40865) );
  IV U50546 ( .A(n37562), .Z(n37563) );
  NOR U50547 ( .A(n37564), .B(n37563), .Z(n40858) );
  IV U50548 ( .A(n37565), .Z(n37567) );
  NOR U50549 ( .A(n37567), .B(n37566), .Z(n40864) );
  NOR U50550 ( .A(n40858), .B(n40864), .Z(n37568) );
  XOR U50551 ( .A(n40865), .B(n37568), .Z(n41455) );
  XOR U50552 ( .A(n40869), .B(n41455), .Z(n38159) );
  NOR U50553 ( .A(n37570), .B(n37569), .Z(n37571) );
  IV U50554 ( .A(n37571), .Z(n38160) );
  XOR U50555 ( .A(n38159), .B(n38160), .Z(n40879) );
  XOR U50556 ( .A(n40878), .B(n40879), .Z(n40876) );
  IV U50557 ( .A(n40876), .Z(n37579) );
  IV U50558 ( .A(n37572), .Z(n37573) );
  NOR U50559 ( .A(n37574), .B(n37573), .Z(n40875) );
  IV U50560 ( .A(n37575), .Z(n37576) );
  NOR U50561 ( .A(n37577), .B(n37576), .Z(n38157) );
  NOR U50562 ( .A(n40875), .B(n38157), .Z(n37578) );
  XOR U50563 ( .A(n37579), .B(n37578), .Z(n38152) );
  XOR U50564 ( .A(n38151), .B(n38152), .Z(n38155) );
  XOR U50565 ( .A(n38154), .B(n38155), .Z(n38147) );
  XOR U50566 ( .A(n38146), .B(n38147), .Z(n38145) );
  XOR U50567 ( .A(n38143), .B(n38145), .Z(n38142) );
  XOR U50568 ( .A(n38140), .B(n38142), .Z(n38135) );
  XOR U50569 ( .A(n38134), .B(n38135), .Z(n38139) );
  XOR U50570 ( .A(n38137), .B(n38139), .Z(n38130) );
  XOR U50571 ( .A(n38129), .B(n38130), .Z(n41429) );
  XOR U50572 ( .A(n38132), .B(n41429), .Z(n38124) );
  IV U50573 ( .A(n37580), .Z(n37582) );
  NOR U50574 ( .A(n37582), .B(n37581), .Z(n38126) );
  IV U50575 ( .A(n37583), .Z(n37585) );
  NOR U50576 ( .A(n37585), .B(n37584), .Z(n38123) );
  NOR U50577 ( .A(n38126), .B(n38123), .Z(n37586) );
  XOR U50578 ( .A(n38124), .B(n37586), .Z(n38121) );
  IV U50579 ( .A(n37587), .Z(n37589) );
  NOR U50580 ( .A(n37589), .B(n37588), .Z(n38119) );
  XOR U50581 ( .A(n38121), .B(n38119), .Z(n40900) );
  XOR U50582 ( .A(n40899), .B(n40900), .Z(n40895) );
  XOR U50583 ( .A(n37590), .B(n40895), .Z(n38112) );
  XOR U50584 ( .A(n38113), .B(n38112), .Z(n40914) );
  XOR U50585 ( .A(n37591), .B(n40914), .Z(n37592) );
  IV U50586 ( .A(n37592), .Z(n40912) );
  XOR U50587 ( .A(n40910), .B(n40912), .Z(n38107) );
  IV U50588 ( .A(n38107), .Z(n37599) );
  IV U50589 ( .A(n37593), .Z(n37595) );
  NOR U50590 ( .A(n37595), .B(n37594), .Z(n38108) );
  IV U50591 ( .A(n37596), .Z(n37597) );
  NOR U50592 ( .A(n37597), .B(n37601), .Z(n38105) );
  NOR U50593 ( .A(n38108), .B(n38105), .Z(n37598) );
  XOR U50594 ( .A(n37599), .B(n37598), .Z(n40923) );
  IV U50595 ( .A(n37600), .Z(n37602) );
  NOR U50596 ( .A(n37602), .B(n37601), .Z(n40921) );
  XOR U50597 ( .A(n40923), .B(n40921), .Z(n38102) );
  XOR U50598 ( .A(n38101), .B(n38102), .Z(n40918) );
  XOR U50599 ( .A(n40917), .B(n40918), .Z(n40931) );
  XOR U50600 ( .A(n40929), .B(n40931), .Z(n40933) );
  XOR U50601 ( .A(n37603), .B(n40933), .Z(n40937) );
  XOR U50602 ( .A(n37604), .B(n40937), .Z(n40945) );
  XOR U50603 ( .A(n40944), .B(n40945), .Z(n38097) );
  XOR U50604 ( .A(n37605), .B(n38097), .Z(n38089) );
  IV U50605 ( .A(n37606), .Z(n37608) );
  NOR U50606 ( .A(n37608), .B(n37607), .Z(n38091) );
  NOR U50607 ( .A(n38088), .B(n38091), .Z(n37609) );
  XOR U50608 ( .A(n38089), .B(n37609), .Z(n38087) );
  IV U50609 ( .A(n37610), .Z(n37611) );
  NOR U50610 ( .A(n37612), .B(n37611), .Z(n38085) );
  IV U50611 ( .A(n37613), .Z(n37615) );
  NOR U50612 ( .A(n37615), .B(n37614), .Z(n38083) );
  NOR U50613 ( .A(n38085), .B(n38083), .Z(n37616) );
  XOR U50614 ( .A(n38087), .B(n37616), .Z(n38081) );
  IV U50615 ( .A(n37617), .Z(n37619) );
  NOR U50616 ( .A(n37619), .B(n37618), .Z(n41372) );
  IV U50617 ( .A(n37620), .Z(n37621) );
  NOR U50618 ( .A(n37622), .B(n37621), .Z(n41365) );
  NOR U50619 ( .A(n41372), .B(n41365), .Z(n38082) );
  XOR U50620 ( .A(n38081), .B(n38082), .Z(n40956) );
  XOR U50621 ( .A(n40955), .B(n40956), .Z(n40960) );
  XOR U50622 ( .A(n37623), .B(n40960), .Z(n37624) );
  IV U50623 ( .A(n37624), .Z(n40963) );
  XOR U50624 ( .A(n40962), .B(n40963), .Z(n40966) );
  XOR U50625 ( .A(n40965), .B(n40966), .Z(n38076) );
  IV U50626 ( .A(n38076), .Z(n37631) );
  IV U50627 ( .A(n37625), .Z(n37627) );
  NOR U50628 ( .A(n37627), .B(n37626), .Z(n38077) );
  IV U50629 ( .A(n37628), .Z(n37629) );
  NOR U50630 ( .A(n37629), .B(n37634), .Z(n38074) );
  NOR U50631 ( .A(n38077), .B(n38074), .Z(n37630) );
  XOR U50632 ( .A(n37631), .B(n37630), .Z(n40971) );
  IV U50633 ( .A(n37632), .Z(n37633) );
  NOR U50634 ( .A(n37634), .B(n37633), .Z(n40969) );
  XOR U50635 ( .A(n40971), .B(n40969), .Z(n40976) );
  XOR U50636 ( .A(n40972), .B(n40976), .Z(n38071) );
  IV U50637 ( .A(n37635), .Z(n37637) );
  NOR U50638 ( .A(n37637), .B(n37636), .Z(n40975) );
  IV U50639 ( .A(n37638), .Z(n37639) );
  NOR U50640 ( .A(n37640), .B(n37639), .Z(n38070) );
  NOR U50641 ( .A(n40975), .B(n38070), .Z(n37641) );
  XOR U50642 ( .A(n38071), .B(n37641), .Z(n38066) );
  XOR U50643 ( .A(n38064), .B(n38066), .Z(n40980) );
  IV U50644 ( .A(n37642), .Z(n37644) );
  NOR U50645 ( .A(n37644), .B(n37643), .Z(n38067) );
  IV U50646 ( .A(n37645), .Z(n37646) );
  NOR U50647 ( .A(n37647), .B(n37646), .Z(n40979) );
  NOR U50648 ( .A(n38067), .B(n40979), .Z(n37648) );
  XOR U50649 ( .A(n40980), .B(n37648), .Z(n40986) );
  IV U50650 ( .A(n37649), .Z(n37651) );
  NOR U50651 ( .A(n37651), .B(n37650), .Z(n40987) );
  NOR U50652 ( .A(n40983), .B(n40987), .Z(n37652) );
  XOR U50653 ( .A(n40986), .B(n37652), .Z(n40996) );
  IV U50654 ( .A(n37653), .Z(n37655) );
  NOR U50655 ( .A(n37655), .B(n37654), .Z(n40982) );
  IV U50656 ( .A(n37656), .Z(n37658) );
  NOR U50657 ( .A(n37658), .B(n37657), .Z(n40995) );
  NOR U50658 ( .A(n40982), .B(n40995), .Z(n37659) );
  XOR U50659 ( .A(n40996), .B(n37659), .Z(n41001) );
  XOR U50660 ( .A(n41002), .B(n41001), .Z(n41327) );
  XOR U50661 ( .A(n37660), .B(n41327), .Z(n41013) );
  IV U50662 ( .A(n37661), .Z(n37662) );
  NOR U50663 ( .A(n37663), .B(n37662), .Z(n41012) );
  IV U50664 ( .A(n37664), .Z(n37665) );
  NOR U50665 ( .A(n37665), .B(n37670), .Z(n41020) );
  NOR U50666 ( .A(n41012), .B(n41020), .Z(n37666) );
  XOR U50667 ( .A(n41013), .B(n37666), .Z(n41019) );
  IV U50668 ( .A(n37667), .Z(n38060) );
  NOR U50669 ( .A(n38060), .B(n37668), .Z(n37672) );
  IV U50670 ( .A(n37669), .Z(n37671) );
  NOR U50671 ( .A(n37671), .B(n37670), .Z(n41017) );
  NOR U50672 ( .A(n37672), .B(n41017), .Z(n37673) );
  XOR U50673 ( .A(n41019), .B(n37673), .Z(n38057) );
  IV U50674 ( .A(n37674), .Z(n37676) );
  NOR U50675 ( .A(n37676), .B(n37675), .Z(n38056) );
  IV U50676 ( .A(n37677), .Z(n37678) );
  NOR U50677 ( .A(n37679), .B(n37678), .Z(n41030) );
  NOR U50678 ( .A(n38056), .B(n41030), .Z(n37680) );
  XOR U50679 ( .A(n38057), .B(n37680), .Z(n41029) );
  XOR U50680 ( .A(n41027), .B(n41029), .Z(n44419) );
  NOR U50681 ( .A(n44415), .B(n41306), .Z(n37681) );
  NOR U50682 ( .A(n37681), .B(n44416), .Z(n38054) );
  XOR U50683 ( .A(n44419), .B(n38054), .Z(n38050) );
  XOR U50684 ( .A(n38048), .B(n38050), .Z(n38053) );
  XOR U50685 ( .A(n38051), .B(n38053), .Z(n38043) );
  XOR U50686 ( .A(n38042), .B(n38043), .Z(n38047) );
  XOR U50687 ( .A(n38045), .B(n38047), .Z(n38039) );
  XOR U50688 ( .A(n38037), .B(n38039), .Z(n41039) );
  XOR U50689 ( .A(n37682), .B(n41039), .Z(n37683) );
  IV U50690 ( .A(n37683), .Z(n41043) );
  XOR U50691 ( .A(n41041), .B(n41043), .Z(n41046) );
  IV U50692 ( .A(n37684), .Z(n37686) );
  NOR U50693 ( .A(n37686), .B(n37685), .Z(n41044) );
  XOR U50694 ( .A(n41046), .B(n41044), .Z(n38035) );
  XOR U50695 ( .A(n38032), .B(n38035), .Z(n41050) );
  IV U50696 ( .A(n37687), .Z(n37688) );
  NOR U50697 ( .A(n37689), .B(n37688), .Z(n38034) );
  IV U50698 ( .A(n37690), .Z(n37691) );
  NOR U50699 ( .A(n37691), .B(n37693), .Z(n38029) );
  IV U50700 ( .A(n37692), .Z(n37694) );
  NOR U50701 ( .A(n37694), .B(n37693), .Z(n41049) );
  NOR U50702 ( .A(n38029), .B(n41049), .Z(n37695) );
  IV U50703 ( .A(n37695), .Z(n37696) );
  NOR U50704 ( .A(n38034), .B(n37696), .Z(n37697) );
  XOR U50705 ( .A(n41050), .B(n37697), .Z(n38027) );
  NOR U50706 ( .A(n37699), .B(n37698), .Z(n44457) );
  NOR U50707 ( .A(n44452), .B(n44457), .Z(n38028) );
  XOR U50708 ( .A(n38027), .B(n38028), .Z(n44464) );
  IV U50709 ( .A(n37700), .Z(n37706) );
  IV U50710 ( .A(n37701), .Z(n37702) );
  NOR U50711 ( .A(n37706), .B(n37702), .Z(n38023) );
  NOR U50712 ( .A(n38025), .B(n38023), .Z(n37703) );
  XOR U50713 ( .A(n44464), .B(n37703), .Z(n38020) );
  IV U50714 ( .A(n37704), .Z(n37705) );
  NOR U50715 ( .A(n37706), .B(n37705), .Z(n37707) );
  IV U50716 ( .A(n37707), .Z(n38021) );
  XOR U50717 ( .A(n38020), .B(n38021), .Z(n41063) );
  XOR U50718 ( .A(n37708), .B(n41063), .Z(n41060) );
  XOR U50719 ( .A(n41061), .B(n41060), .Z(n41263) );
  XOR U50720 ( .A(n37709), .B(n41263), .Z(n41071) );
  XOR U50721 ( .A(n41072), .B(n41071), .Z(n37710) );
  IV U50722 ( .A(n37710), .Z(n38013) );
  XOR U50723 ( .A(n38012), .B(n38013), .Z(n41074) );
  IV U50724 ( .A(n37711), .Z(n37713) );
  NOR U50725 ( .A(n37713), .B(n37712), .Z(n41073) );
  IV U50726 ( .A(n37714), .Z(n37716) );
  NOR U50727 ( .A(n37716), .B(n37715), .Z(n38010) );
  NOR U50728 ( .A(n41073), .B(n38010), .Z(n37717) );
  XOR U50729 ( .A(n41074), .B(n37717), .Z(n38007) );
  IV U50730 ( .A(n37718), .Z(n37719) );
  NOR U50731 ( .A(n37720), .B(n37719), .Z(n38008) );
  IV U50732 ( .A(n37721), .Z(n37728) );
  NOR U50733 ( .A(n37723), .B(n37722), .Z(n37724) );
  IV U50734 ( .A(n37724), .Z(n37725) );
  NOR U50735 ( .A(n37726), .B(n37725), .Z(n37727) );
  IV U50736 ( .A(n37727), .Z(n37731) );
  NOR U50737 ( .A(n37728), .B(n37731), .Z(n41082) );
  NOR U50738 ( .A(n38008), .B(n41082), .Z(n37729) );
  XOR U50739 ( .A(n38007), .B(n37729), .Z(n41087) );
  IV U50740 ( .A(n37730), .Z(n37732) );
  NOR U50741 ( .A(n37732), .B(n37731), .Z(n41085) );
  XOR U50742 ( .A(n41087), .B(n41085), .Z(n41247) );
  IV U50743 ( .A(n37733), .Z(n37734) );
  NOR U50744 ( .A(n37735), .B(n37734), .Z(n41251) );
  NOR U50745 ( .A(n41251), .B(n41246), .Z(n41089) );
  XOR U50746 ( .A(n41247), .B(n41089), .Z(n41091) );
  XOR U50747 ( .A(n37736), .B(n41091), .Z(n41097) );
  XOR U50748 ( .A(n41095), .B(n41097), .Z(n38003) );
  IV U50749 ( .A(n37737), .Z(n37738) );
  NOR U50750 ( .A(n37739), .B(n37738), .Z(n38001) );
  XOR U50751 ( .A(n38003), .B(n38001), .Z(n38006) );
  IV U50752 ( .A(n37740), .Z(n37741) );
  NOR U50753 ( .A(n37742), .B(n37741), .Z(n38004) );
  XOR U50754 ( .A(n38006), .B(n38004), .Z(n37996) );
  XOR U50755 ( .A(n37995), .B(n37996), .Z(n37999) );
  XOR U50756 ( .A(n37998), .B(n37999), .Z(n37992) );
  IV U50757 ( .A(n37992), .Z(n37749) );
  IV U50758 ( .A(n37743), .Z(n37747) );
  NOR U50759 ( .A(n37745), .B(n37744), .Z(n37746) );
  IV U50760 ( .A(n37746), .Z(n37751) );
  NOR U50761 ( .A(n37747), .B(n37751), .Z(n37989) );
  NOR U50762 ( .A(n37991), .B(n37989), .Z(n37748) );
  XOR U50763 ( .A(n37749), .B(n37748), .Z(n41110) );
  IV U50764 ( .A(n37750), .Z(n37752) );
  NOR U50765 ( .A(n37752), .B(n37751), .Z(n41108) );
  XOR U50766 ( .A(n41110), .B(n41108), .Z(n37987) );
  XOR U50767 ( .A(n37985), .B(n37987), .Z(n41105) );
  XOR U50768 ( .A(n41104), .B(n41105), .Z(n37982) );
  XOR U50769 ( .A(n37753), .B(n37982), .Z(n37754) );
  IV U50770 ( .A(n37754), .Z(n37978) );
  IV U50771 ( .A(n37755), .Z(n37757) );
  NOR U50772 ( .A(n37757), .B(n37756), .Z(n37763) );
  IV U50773 ( .A(n37763), .Z(n37758) );
  NOR U50774 ( .A(n37978), .B(n37758), .Z(n44495) );
  IV U50775 ( .A(n37759), .Z(n37761) );
  NOR U50776 ( .A(n37761), .B(n37760), .Z(n37976) );
  XOR U50777 ( .A(n37976), .B(n37978), .Z(n37767) );
  IV U50778 ( .A(n37767), .Z(n37762) );
  NOR U50779 ( .A(n37763), .B(n37762), .Z(n37764) );
  NOR U50780 ( .A(n44495), .B(n37764), .Z(n37765) );
  NOR U50781 ( .A(n37766), .B(n37765), .Z(n37769) );
  IV U50782 ( .A(n37766), .Z(n37768) );
  NOR U50783 ( .A(n37768), .B(n37767), .Z(n44498) );
  NOR U50784 ( .A(n37769), .B(n44498), .Z(n41118) );
  XOR U50785 ( .A(n41120), .B(n41118), .Z(n37966) );
  NOR U50786 ( .A(n37771), .B(n37770), .Z(n37772) );
  IV U50787 ( .A(n37772), .Z(n37967) );
  NOR U50788 ( .A(n37773), .B(n37967), .Z(n37777) );
  IV U50789 ( .A(n37774), .Z(n37775) );
  NOR U50790 ( .A(n37776), .B(n37775), .Z(n37960) );
  NOR U50791 ( .A(n37777), .B(n37960), .Z(n37778) );
  XOR U50792 ( .A(n37966), .B(n37778), .Z(n37957) );
  XOR U50793 ( .A(n37779), .B(n37957), .Z(n41129) );
  XOR U50794 ( .A(n37780), .B(n41129), .Z(n37781) );
  IV U50795 ( .A(n37781), .Z(n37954) );
  XOR U50796 ( .A(n37952), .B(n37954), .Z(n37951) );
  IV U50797 ( .A(n37782), .Z(n37786) );
  NOR U50798 ( .A(n37784), .B(n37783), .Z(n37785) );
  XOR U50799 ( .A(n37786), .B(n37785), .Z(n37808) );
  NOR U50800 ( .A(n37788), .B(n37787), .Z(n37789) );
  XOR U50801 ( .A(n37790), .B(n37789), .Z(n37813) );
  IV U50802 ( .A(n37813), .Z(n37802) );
  IV U50803 ( .A(n37791), .Z(n37793) );
  NOR U50804 ( .A(n37793), .B(n37792), .Z(n37806) );
  IV U50805 ( .A(n37806), .Z(n37794) );
  NOR U50806 ( .A(n37802), .B(n37794), .Z(n37795) );
  IV U50807 ( .A(n37795), .Z(n37796) );
  NOR U50808 ( .A(n37816), .B(n37796), .Z(n37807) );
  IV U50809 ( .A(n37807), .Z(n37797) );
  NOR U50810 ( .A(n37808), .B(n37797), .Z(n37949) );
  IV U50811 ( .A(n37798), .Z(n37800) );
  NOR U50812 ( .A(n37800), .B(n37799), .Z(n37801) );
  NOR U50813 ( .A(n37806), .B(n37801), .Z(n37814) );
  NOR U50814 ( .A(n37802), .B(n37814), .Z(n37833) );
  IV U50815 ( .A(n37833), .Z(n37803) );
  NOR U50816 ( .A(n37816), .B(n37803), .Z(n37804) );
  IV U50817 ( .A(n37804), .Z(n37805) );
  NOR U50818 ( .A(n37806), .B(n37805), .Z(n37812) );
  IV U50819 ( .A(n37812), .Z(n37809) );
  XOR U50820 ( .A(n37808), .B(n37807), .Z(n37811) );
  NOR U50821 ( .A(n37809), .B(n37811), .Z(n37947) );
  NOR U50822 ( .A(n37949), .B(n37947), .Z(n37810) );
  XOR U50823 ( .A(n37951), .B(n37810), .Z(n41187) );
  XOR U50824 ( .A(n37812), .B(n37811), .Z(n37832) );
  XOR U50825 ( .A(n37814), .B(n37813), .Z(n37850) );
  XOR U50826 ( .A(n37816), .B(n37815), .Z(n37855) );
  IV U50827 ( .A(n37855), .Z(n37817) );
  NOR U50828 ( .A(n37850), .B(n37817), .Z(n37818) );
  IV U50829 ( .A(n37818), .Z(n37828) );
  IV U50830 ( .A(n37819), .Z(n37821) );
  NOR U50831 ( .A(n37821), .B(n37820), .Z(n37837) );
  IV U50832 ( .A(n37837), .Z(n37822) );
  NOR U50833 ( .A(n37828), .B(n37822), .Z(n37823) );
  IV U50834 ( .A(n37823), .Z(n37845) );
  NOR U50835 ( .A(n37832), .B(n37845), .Z(n41132) );
  IV U50836 ( .A(n37824), .Z(n37825) );
  NOR U50837 ( .A(n37826), .B(n37825), .Z(n37838) );
  IV U50838 ( .A(n37838), .Z(n37827) );
  NOR U50839 ( .A(n37828), .B(n37827), .Z(n37831) );
  IV U50840 ( .A(n37831), .Z(n37829) );
  NOR U50841 ( .A(n37832), .B(n37829), .Z(n37945) );
  NOR U50842 ( .A(n41132), .B(n37945), .Z(n37830) );
  XOR U50843 ( .A(n41187), .B(n37830), .Z(n41136) );
  XOR U50844 ( .A(n37832), .B(n37831), .Z(n37844) );
  NOR U50845 ( .A(n37834), .B(n37833), .Z(n37836) );
  XOR U50846 ( .A(n37836), .B(n37835), .Z(n37852) );
  NOR U50847 ( .A(n37838), .B(n37837), .Z(n37851) );
  XOR U50848 ( .A(n37850), .B(n37851), .Z(n37888) );
  IV U50849 ( .A(n37888), .Z(n37862) );
  IV U50850 ( .A(n37839), .Z(n37841) );
  NOR U50851 ( .A(n37841), .B(n37840), .Z(n37886) );
  IV U50852 ( .A(n37886), .Z(n37869) );
  NOR U50853 ( .A(n37862), .B(n37869), .Z(n37866) );
  IV U50854 ( .A(n37866), .Z(n37842) );
  NOR U50855 ( .A(n37852), .B(n37842), .Z(n37846) );
  IV U50856 ( .A(n37846), .Z(n37843) );
  NOR U50857 ( .A(n37844), .B(n37843), .Z(n41134) );
  XOR U50858 ( .A(n41136), .B(n41134), .Z(n41148) );
  XOR U50859 ( .A(n37844), .B(n37843), .Z(n37848) );
  NOR U50860 ( .A(n37846), .B(n37845), .Z(n37847) );
  NOR U50861 ( .A(n37848), .B(n37847), .Z(n37849) );
  NOR U50862 ( .A(n41132), .B(n37849), .Z(n37881) );
  IV U50863 ( .A(n37881), .Z(n37878) );
  NOR U50864 ( .A(n37851), .B(n37850), .Z(n37853) );
  NOR U50865 ( .A(n37853), .B(n37852), .Z(n37857) );
  IV U50866 ( .A(n37853), .Z(n37854) );
  NOR U50867 ( .A(n37855), .B(n37854), .Z(n37856) );
  NOR U50868 ( .A(n37857), .B(n37856), .Z(n37867) );
  IV U50869 ( .A(n37858), .Z(n37860) );
  NOR U50870 ( .A(n37860), .B(n37859), .Z(n37885) );
  IV U50871 ( .A(n37885), .Z(n37861) );
  NOR U50872 ( .A(n37862), .B(n37861), .Z(n37865) );
  IV U50873 ( .A(n37865), .Z(n37863) );
  NOR U50874 ( .A(n37867), .B(n37863), .Z(n37880) );
  IV U50875 ( .A(n37880), .Z(n37864) );
  NOR U50876 ( .A(n37878), .B(n37864), .Z(n41146) );
  XOR U50877 ( .A(n41148), .B(n41146), .Z(n41141) );
  NOR U50878 ( .A(n37866), .B(n37865), .Z(n37868) );
  XOR U50879 ( .A(n37868), .B(n37867), .Z(n37883) );
  IV U50880 ( .A(n37883), .Z(n37876) );
  XOR U50881 ( .A(n37869), .B(n37888), .Z(n37874) );
  IV U50882 ( .A(n37870), .Z(n37872) );
  NOR U50883 ( .A(n37872), .B(n37871), .Z(n37898) );
  IV U50884 ( .A(n37898), .Z(n37873) );
  NOR U50885 ( .A(n37874), .B(n37873), .Z(n37875) );
  IV U50886 ( .A(n37875), .Z(n37884) );
  NOR U50887 ( .A(n37876), .B(n37884), .Z(n37879) );
  IV U50888 ( .A(n37879), .Z(n37877) );
  NOR U50889 ( .A(n37878), .B(n37877), .Z(n41139) );
  XOR U50890 ( .A(n41141), .B(n41139), .Z(n41167) );
  NOR U50891 ( .A(n37880), .B(n37879), .Z(n37882) );
  XOR U50892 ( .A(n37882), .B(n37881), .Z(n37922) );
  XOR U50893 ( .A(n37884), .B(n37883), .Z(n37895) );
  NOR U50894 ( .A(n37886), .B(n37885), .Z(n37887) );
  XOR U50895 ( .A(n37888), .B(n37887), .Z(n37900) );
  IV U50896 ( .A(n37889), .Z(n37891) );
  NOR U50897 ( .A(n37891), .B(n37890), .Z(n37897) );
  IV U50898 ( .A(n37897), .Z(n37892) );
  NOR U50899 ( .A(n37900), .B(n37892), .Z(n37896) );
  IV U50900 ( .A(n37896), .Z(n37893) );
  NOR U50901 ( .A(n37895), .B(n37893), .Z(n37907) );
  IV U50902 ( .A(n37907), .Z(n37894) );
  NOR U50903 ( .A(n37922), .B(n37894), .Z(n41143) );
  XOR U50904 ( .A(n41167), .B(n41143), .Z(n41162) );
  XOR U50905 ( .A(n37896), .B(n37895), .Z(n44547) );
  NOR U50906 ( .A(n37898), .B(n37897), .Z(n37899) );
  XOR U50907 ( .A(n37900), .B(n37899), .Z(n37924) );
  IV U50908 ( .A(n37924), .Z(n37913) );
  IV U50909 ( .A(n37901), .Z(n37903) );
  NOR U50910 ( .A(n37903), .B(n37902), .Z(n37917) );
  IV U50911 ( .A(n37917), .Z(n37904) );
  NOR U50912 ( .A(n37913), .B(n37904), .Z(n37905) );
  IV U50913 ( .A(n37905), .Z(n37906) );
  NOR U50914 ( .A(n44547), .B(n37906), .Z(n37920) );
  NOR U50915 ( .A(n37907), .B(n37920), .Z(n37908) );
  XOR U50916 ( .A(n37908), .B(n37922), .Z(n37934) );
  IV U50917 ( .A(n37934), .Z(n37919) );
  IV U50918 ( .A(n37909), .Z(n37911) );
  NOR U50919 ( .A(n37911), .B(n37910), .Z(n37912) );
  NOR U50920 ( .A(n37917), .B(n37912), .Z(n37925) );
  NOR U50921 ( .A(n37913), .B(n37925), .Z(n44544) );
  IV U50922 ( .A(n44544), .Z(n37914) );
  NOR U50923 ( .A(n44547), .B(n37914), .Z(n37915) );
  IV U50924 ( .A(n37915), .Z(n37916) );
  NOR U50925 ( .A(n37917), .B(n37916), .Z(n37918) );
  IV U50926 ( .A(n37918), .Z(n37935) );
  NOR U50927 ( .A(n37919), .B(n37935), .Z(n41165) );
  IV U50928 ( .A(n37920), .Z(n37921) );
  NOR U50929 ( .A(n37922), .B(n37921), .Z(n41160) );
  NOR U50930 ( .A(n41165), .B(n41160), .Z(n37923) );
  XOR U50931 ( .A(n41162), .B(n37923), .Z(n44586) );
  IV U50932 ( .A(n44586), .Z(n44562) );
  XOR U50933 ( .A(n37925), .B(n37924), .Z(n44553) );
  IV U50934 ( .A(n37926), .Z(n37928) );
  NOR U50935 ( .A(n37928), .B(n37927), .Z(n44551) );
  IV U50936 ( .A(n44551), .Z(n37929) );
  NOR U50937 ( .A(n44553), .B(n37929), .Z(n41154) );
  IV U50938 ( .A(n37930), .Z(n37932) );
  NOR U50939 ( .A(n37932), .B(n37931), .Z(n44550) );
  IV U50940 ( .A(n44550), .Z(n37933) );
  NOR U50941 ( .A(n44553), .B(n37933), .Z(n41174) );
  NOR U50942 ( .A(n41154), .B(n41174), .Z(n44543) );
  NOR U50943 ( .A(n44543), .B(n44547), .Z(n44581) );
  XOR U50944 ( .A(n37935), .B(n37934), .Z(n44583) );
  XOR U50945 ( .A(n44581), .B(n44583), .Z(n44565) );
  XOR U50946 ( .A(n44544), .B(n44547), .Z(n37942) );
  XOR U50947 ( .A(n44551), .B(n44553), .Z(n37940) );
  IV U50948 ( .A(n37936), .Z(n37938) );
  NOR U50949 ( .A(n37938), .B(n37937), .Z(n44569) );
  IV U50950 ( .A(n44569), .Z(n37939) );
  NOR U50951 ( .A(n37940), .B(n37939), .Z(n44571) );
  IV U50952 ( .A(n44571), .Z(n37941) );
  NOR U50953 ( .A(n37942), .B(n37941), .Z(n44566) );
  IV U50954 ( .A(n44566), .Z(n37943) );
  NOR U50955 ( .A(n44565), .B(n37943), .Z(n44579) );
  IV U50956 ( .A(n44579), .Z(n37944) );
  NOR U50957 ( .A(n44562), .B(n37944), .Z(n44540) );
  IV U50958 ( .A(n44540), .Z(n41173) );
  IV U50959 ( .A(n41187), .Z(n41133) );
  IV U50960 ( .A(n37945), .Z(n41186) );
  NOR U50961 ( .A(n41133), .B(n41186), .Z(n37946) );
  IV U50962 ( .A(n37946), .Z(n41197) );
  IV U50963 ( .A(n37947), .Z(n37948) );
  NOR U50964 ( .A(n37951), .B(n37948), .Z(n41193) );
  IV U50965 ( .A(n37949), .Z(n37950) );
  NOR U50966 ( .A(n37951), .B(n37950), .Z(n44513) );
  IV U50967 ( .A(n37952), .Z(n37953) );
  NOR U50968 ( .A(n37954), .B(n37953), .Z(n44516) );
  IV U50969 ( .A(n37955), .Z(n37956) );
  NOR U50970 ( .A(n37956), .B(n41129), .Z(n44509) );
  NOR U50971 ( .A(n44516), .B(n44509), .Z(n41131) );
  IV U50972 ( .A(n37957), .Z(n41127) );
  IV U50973 ( .A(n37958), .Z(n37959) );
  NOR U50974 ( .A(n41127), .B(n37959), .Z(n41198) );
  IV U50975 ( .A(n37960), .Z(n37961) );
  NOR U50976 ( .A(n37961), .B(n37966), .Z(n44503) );
  IV U50977 ( .A(n37962), .Z(n37964) );
  NOR U50978 ( .A(n37964), .B(n37963), .Z(n37965) );
  IV U50979 ( .A(n37965), .Z(n37972) );
  NOR U50980 ( .A(n37967), .B(n37966), .Z(n37968) );
  IV U50981 ( .A(n37968), .Z(n37969) );
  NOR U50982 ( .A(n37970), .B(n37969), .Z(n37971) );
  IV U50983 ( .A(n37971), .Z(n37974) );
  NOR U50984 ( .A(n37972), .B(n37974), .Z(n41203) );
  NOR U50985 ( .A(n44503), .B(n41203), .Z(n41123) );
  IV U50986 ( .A(n37973), .Z(n37975) );
  NOR U50987 ( .A(n37975), .B(n37974), .Z(n41201) );
  IV U50988 ( .A(n37976), .Z(n37977) );
  NOR U50989 ( .A(n37978), .B(n37977), .Z(n41208) );
  IV U50990 ( .A(n37979), .Z(n37980) );
  NOR U50991 ( .A(n37980), .B(n37982), .Z(n41212) );
  NOR U50992 ( .A(n41208), .B(n41212), .Z(n41116) );
  IV U50993 ( .A(n37981), .Z(n37983) );
  NOR U50994 ( .A(n37983), .B(n37982), .Z(n37984) );
  IV U50995 ( .A(n37984), .Z(n41216) );
  IV U50996 ( .A(n37985), .Z(n37986) );
  NOR U50997 ( .A(n37987), .B(n37986), .Z(n37988) );
  IV U50998 ( .A(n37988), .Z(n41111) );
  IV U50999 ( .A(n37989), .Z(n37990) );
  NOR U51000 ( .A(n37992), .B(n37990), .Z(n41224) );
  IV U51001 ( .A(n37991), .Z(n37993) );
  NOR U51002 ( .A(n37993), .B(n37992), .Z(n37994) );
  IV U51003 ( .A(n37994), .Z(n41222) );
  IV U51004 ( .A(n37995), .Z(n37997) );
  NOR U51005 ( .A(n37997), .B(n37996), .Z(n41229) );
  IV U51006 ( .A(n37998), .Z(n38000) );
  NOR U51007 ( .A(n38000), .B(n37999), .Z(n41227) );
  NOR U51008 ( .A(n41229), .B(n41227), .Z(n41103) );
  IV U51009 ( .A(n38001), .Z(n38002) );
  NOR U51010 ( .A(n38003), .B(n38002), .Z(n41235) );
  IV U51011 ( .A(n38004), .Z(n38005) );
  NOR U51012 ( .A(n38006), .B(n38005), .Z(n41232) );
  NOR U51013 ( .A(n41235), .B(n41232), .Z(n41102) );
  IV U51014 ( .A(n38007), .Z(n41084) );
  IV U51015 ( .A(n38008), .Z(n38009) );
  NOR U51016 ( .A(n41084), .B(n38009), .Z(n41259) );
  IV U51017 ( .A(n38010), .Z(n38011) );
  NOR U51018 ( .A(n38011), .B(n41074), .Z(n44486) );
  NOR U51019 ( .A(n41259), .B(n44486), .Z(n41081) );
  IV U51020 ( .A(n38012), .Z(n38014) );
  NOR U51021 ( .A(n38014), .B(n38013), .Z(n38015) );
  IV U51022 ( .A(n38015), .Z(n41076) );
  IV U51023 ( .A(n38016), .Z(n38019) );
  NOR U51024 ( .A(n38017), .B(n41263), .Z(n38018) );
  IV U51025 ( .A(n38018), .Z(n41069) );
  NOR U51026 ( .A(n38019), .B(n41069), .Z(n41270) );
  IV U51027 ( .A(n38020), .Z(n38022) );
  NOR U51028 ( .A(n38022), .B(n38021), .Z(n41283) );
  IV U51029 ( .A(n38023), .Z(n38024) );
  NOR U51030 ( .A(n44464), .B(n38024), .Z(n41285) );
  NOR U51031 ( .A(n41283), .B(n41285), .Z(n41056) );
  IV U51032 ( .A(n38025), .Z(n38026) );
  NOR U51033 ( .A(n38026), .B(n44464), .Z(n41055) );
  IV U51034 ( .A(n38027), .Z(n44454) );
  NOR U51035 ( .A(n44454), .B(n38028), .Z(n38031) );
  IV U51036 ( .A(n38029), .Z(n38030) );
  NOR U51037 ( .A(n38030), .B(n41050), .Z(n44450) );
  NOR U51038 ( .A(n38031), .B(n44450), .Z(n41054) );
  IV U51039 ( .A(n38032), .Z(n38033) );
  NOR U51040 ( .A(n38033), .B(n38035), .Z(n44444) );
  IV U51041 ( .A(n38034), .Z(n38036) );
  NOR U51042 ( .A(n38036), .B(n38035), .Z(n44446) );
  NOR U51043 ( .A(n44444), .B(n44446), .Z(n41053) );
  IV U51044 ( .A(n38037), .Z(n38038) );
  NOR U51045 ( .A(n38039), .B(n38038), .Z(n48200) );
  IV U51046 ( .A(n38040), .Z(n38041) );
  NOR U51047 ( .A(n41039), .B(n38041), .Z(n48192) );
  NOR U51048 ( .A(n48200), .B(n48192), .Z(n41290) );
  IV U51049 ( .A(n38042), .Z(n38044) );
  NOR U51050 ( .A(n38044), .B(n38043), .Z(n41298) );
  IV U51051 ( .A(n38045), .Z(n38046) );
  NOR U51052 ( .A(n38047), .B(n38046), .Z(n41295) );
  NOR U51053 ( .A(n41298), .B(n41295), .Z(n41036) );
  IV U51054 ( .A(n38048), .Z(n38049) );
  NOR U51055 ( .A(n38050), .B(n38049), .Z(n41304) );
  IV U51056 ( .A(n38051), .Z(n38052) );
  NOR U51057 ( .A(n38053), .B(n38052), .Z(n41301) );
  NOR U51058 ( .A(n41304), .B(n41301), .Z(n41035) );
  IV U51059 ( .A(n38054), .Z(n38055) );
  NOR U51060 ( .A(n38055), .B(n44419), .Z(n41307) );
  IV U51061 ( .A(n38056), .Z(n38058) );
  IV U51062 ( .A(n38057), .Z(n41031) );
  NOR U51063 ( .A(n38058), .B(n41031), .Z(n41312) );
  IV U51064 ( .A(n38059), .Z(n38062) );
  NOR U51065 ( .A(n38060), .B(n41019), .Z(n38061) );
  IV U51066 ( .A(n38061), .Z(n41025) );
  NOR U51067 ( .A(n38062), .B(n41025), .Z(n44404) );
  IV U51068 ( .A(n41328), .Z(n38063) );
  NOR U51069 ( .A(n38063), .B(n41327), .Z(n41008) );
  IV U51070 ( .A(n41008), .Z(n41000) );
  IV U51071 ( .A(n38064), .Z(n38065) );
  NOR U51072 ( .A(n38066), .B(n38065), .Z(n41354) );
  IV U51073 ( .A(n38067), .Z(n38068) );
  NOR U51074 ( .A(n38068), .B(n40980), .Z(n41352) );
  NOR U51075 ( .A(n41354), .B(n41352), .Z(n38069) );
  IV U51076 ( .A(n38069), .Z(n40978) );
  IV U51077 ( .A(n38070), .Z(n38073) );
  IV U51078 ( .A(n38071), .Z(n38072) );
  NOR U51079 ( .A(n38073), .B(n38072), .Z(n44393) );
  IV U51080 ( .A(n38074), .Z(n38075) );
  NOR U51081 ( .A(n38076), .B(n38075), .Z(n41357) );
  IV U51082 ( .A(n38077), .Z(n38078) );
  NOR U51083 ( .A(n38078), .B(n40966), .Z(n44378) );
  IV U51084 ( .A(n38079), .Z(n38080) );
  NOR U51085 ( .A(n38080), .B(n40960), .Z(n44365) );
  IV U51086 ( .A(n38081), .Z(n41366) );
  NOR U51087 ( .A(n38082), .B(n41366), .Z(n40954) );
  IV U51088 ( .A(n38083), .Z(n38084) );
  NOR U51089 ( .A(n38087), .B(n38084), .Z(n41369) );
  IV U51090 ( .A(n38085), .Z(n38086) );
  NOR U51091 ( .A(n38087), .B(n38086), .Z(n41375) );
  IV U51092 ( .A(n38088), .Z(n38090) );
  IV U51093 ( .A(n38089), .Z(n38092) );
  NOR U51094 ( .A(n38090), .B(n38092), .Z(n41378) );
  NOR U51095 ( .A(n41375), .B(n41378), .Z(n40952) );
  IV U51096 ( .A(n38091), .Z(n38093) );
  NOR U51097 ( .A(n38093), .B(n38092), .Z(n41380) );
  IV U51098 ( .A(n38094), .Z(n38095) );
  NOR U51099 ( .A(n38095), .B(n38097), .Z(n44354) );
  IV U51100 ( .A(n38096), .Z(n38098) );
  NOR U51101 ( .A(n38098), .B(n38097), .Z(n44351) );
  IV U51102 ( .A(n38099), .Z(n38100) );
  NOR U51103 ( .A(n38100), .B(n40933), .Z(n41391) );
  IV U51104 ( .A(n38101), .Z(n38103) );
  NOR U51105 ( .A(n38103), .B(n38102), .Z(n38104) );
  IV U51106 ( .A(n38104), .Z(n40924) );
  IV U51107 ( .A(n38105), .Z(n38106) );
  NOR U51108 ( .A(n38107), .B(n38106), .Z(n44329) );
  IV U51109 ( .A(n38108), .Z(n38109) );
  NOR U51110 ( .A(n40912), .B(n38109), .Z(n41401) );
  IV U51111 ( .A(n38110), .Z(n38111) );
  NOR U51112 ( .A(n38111), .B(n40914), .Z(n41404) );
  IV U51113 ( .A(n38112), .Z(n41421) );
  NOR U51114 ( .A(n41421), .B(n38113), .Z(n38116) );
  IV U51115 ( .A(n38114), .Z(n38115) );
  NOR U51116 ( .A(n38115), .B(n40914), .Z(n41407) );
  NOR U51117 ( .A(n38116), .B(n41407), .Z(n40909) );
  IV U51118 ( .A(n38117), .Z(n38118) );
  NOR U51119 ( .A(n40895), .B(n38118), .Z(n41422) );
  IV U51120 ( .A(n38119), .Z(n38120) );
  NOR U51121 ( .A(n38121), .B(n38120), .Z(n38122) );
  IV U51122 ( .A(n38122), .Z(n41426) );
  IV U51123 ( .A(n38123), .Z(n38125) );
  IV U51124 ( .A(n38124), .Z(n38127) );
  NOR U51125 ( .A(n38125), .B(n38127), .Z(n44317) );
  IV U51126 ( .A(n38126), .Z(n38128) );
  NOR U51127 ( .A(n38128), .B(n38127), .Z(n44314) );
  IV U51128 ( .A(n38129), .Z(n38131) );
  NOR U51129 ( .A(n38131), .B(n38130), .Z(n41435) );
  NOR U51130 ( .A(n38132), .B(n41429), .Z(n38133) );
  NOR U51131 ( .A(n41435), .B(n38133), .Z(n40893) );
  IV U51132 ( .A(n38134), .Z(n38136) );
  NOR U51133 ( .A(n38136), .B(n38135), .Z(n41440) );
  IV U51134 ( .A(n38137), .Z(n38138) );
  NOR U51135 ( .A(n38139), .B(n38138), .Z(n41438) );
  NOR U51136 ( .A(n41440), .B(n41438), .Z(n40892) );
  IV U51137 ( .A(n38140), .Z(n38141) );
  NOR U51138 ( .A(n38142), .B(n38141), .Z(n41444) );
  IV U51139 ( .A(n38143), .Z(n38144) );
  NOR U51140 ( .A(n38145), .B(n38144), .Z(n41446) );
  IV U51141 ( .A(n38146), .Z(n38148) );
  NOR U51142 ( .A(n38148), .B(n38147), .Z(n41448) );
  NOR U51143 ( .A(n41446), .B(n41448), .Z(n38149) );
  IV U51144 ( .A(n38149), .Z(n38150) );
  NOR U51145 ( .A(n41444), .B(n38150), .Z(n40891) );
  IV U51146 ( .A(n38151), .Z(n38153) );
  NOR U51147 ( .A(n38153), .B(n38152), .Z(n44309) );
  IV U51148 ( .A(n38154), .Z(n38156) );
  NOR U51149 ( .A(n38156), .B(n38155), .Z(n41451) );
  NOR U51150 ( .A(n44309), .B(n41451), .Z(n40890) );
  IV U51151 ( .A(n38157), .Z(n38158) );
  NOR U51152 ( .A(n38158), .B(n40876), .Z(n44306) );
  IV U51153 ( .A(n38159), .Z(n38161) );
  NOR U51154 ( .A(n38161), .B(n38160), .Z(n40873) );
  IV U51155 ( .A(n40873), .Z(n40868) );
  IV U51156 ( .A(n38162), .Z(n38163) );
  NOR U51157 ( .A(n38163), .B(n40859), .Z(n40852) );
  IV U51158 ( .A(n40860), .Z(n38164) );
  NOR U51159 ( .A(n38164), .B(n40859), .Z(n40850) );
  IV U51160 ( .A(n40850), .Z(n40841) );
  IV U51161 ( .A(n38165), .Z(n38166) );
  NOR U51162 ( .A(n38167), .B(n38166), .Z(n38168) );
  IV U51163 ( .A(n38168), .Z(n41459) );
  IV U51164 ( .A(n38169), .Z(n38170) );
  NOR U51165 ( .A(n38171), .B(n38170), .Z(n41463) );
  IV U51166 ( .A(n38172), .Z(n38174) );
  NOR U51167 ( .A(n38174), .B(n38173), .Z(n41461) );
  NOR U51168 ( .A(n41463), .B(n41461), .Z(n40839) );
  IV U51169 ( .A(n38175), .Z(n38177) );
  NOR U51170 ( .A(n38177), .B(n38176), .Z(n44283) );
  IV U51171 ( .A(n38178), .Z(n38183) );
  IV U51172 ( .A(n38179), .Z(n38180) );
  NOR U51173 ( .A(n38183), .B(n38180), .Z(n44277) );
  NOR U51174 ( .A(n44283), .B(n44277), .Z(n40838) );
  IV U51175 ( .A(n38181), .Z(n38185) );
  NOR U51176 ( .A(n38183), .B(n38182), .Z(n38184) );
  IV U51177 ( .A(n38184), .Z(n38187) );
  NOR U51178 ( .A(n38185), .B(n38187), .Z(n44275) );
  IV U51179 ( .A(n38186), .Z(n38188) );
  NOR U51180 ( .A(n38188), .B(n38187), .Z(n44272) );
  IV U51181 ( .A(n38189), .Z(n38190) );
  NOR U51182 ( .A(n38190), .B(n38196), .Z(n44266) );
  NOR U51183 ( .A(n44272), .B(n44266), .Z(n40837) );
  IV U51184 ( .A(n38191), .Z(n38194) );
  IV U51185 ( .A(n41474), .Z(n40834) );
  NOR U51186 ( .A(n40834), .B(n38192), .Z(n38193) );
  IV U51187 ( .A(n38193), .Z(n38199) );
  NOR U51188 ( .A(n38194), .B(n38199), .Z(n41469) );
  IV U51189 ( .A(n38195), .Z(n38197) );
  NOR U51190 ( .A(n38197), .B(n38196), .Z(n44268) );
  NOR U51191 ( .A(n41469), .B(n44268), .Z(n40836) );
  IV U51192 ( .A(n38198), .Z(n38200) );
  NOR U51193 ( .A(n38200), .B(n38199), .Z(n41466) );
  IV U51194 ( .A(n38201), .Z(n41475) );
  NOR U51195 ( .A(n40834), .B(n41475), .Z(n41486) );
  IV U51196 ( .A(n38202), .Z(n38203) );
  NOR U51197 ( .A(n38203), .B(n38209), .Z(n41488) );
  NOR U51198 ( .A(n41486), .B(n41488), .Z(n40831) );
  IV U51199 ( .A(n38204), .Z(n38205) );
  NOR U51200 ( .A(n38206), .B(n38205), .Z(n44254) );
  IV U51201 ( .A(n38207), .Z(n38208) );
  NOR U51202 ( .A(n38209), .B(n38208), .Z(n44262) );
  NOR U51203 ( .A(n44254), .B(n44262), .Z(n40830) );
  IV U51204 ( .A(n38210), .Z(n44250) );
  NOR U51205 ( .A(n44250), .B(n38211), .Z(n40829) );
  IV U51206 ( .A(n38212), .Z(n38213) );
  NOR U51207 ( .A(n38213), .B(n40825), .Z(n41491) );
  IV U51208 ( .A(n38214), .Z(n38215) );
  NOR U51209 ( .A(n38215), .B(n40825), .Z(n44240) );
  IV U51210 ( .A(n38216), .Z(n38217) );
  NOR U51211 ( .A(n38217), .B(n38223), .Z(n44232) );
  IV U51212 ( .A(n38218), .Z(n38219) );
  NOR U51213 ( .A(n38220), .B(n38219), .Z(n44225) );
  IV U51214 ( .A(n38221), .Z(n38222) );
  NOR U51215 ( .A(n38223), .B(n38222), .Z(n44229) );
  NOR U51216 ( .A(n44225), .B(n44229), .Z(n40819) );
  IV U51217 ( .A(n38224), .Z(n38225) );
  NOR U51218 ( .A(n38226), .B(n38225), .Z(n44214) );
  IV U51219 ( .A(n38227), .Z(n38232) );
  IV U51220 ( .A(n38228), .Z(n38229) );
  NOR U51221 ( .A(n38232), .B(n38229), .Z(n44210) );
  IV U51222 ( .A(n38230), .Z(n38231) );
  NOR U51223 ( .A(n38232), .B(n38231), .Z(n44217) );
  IV U51224 ( .A(n38233), .Z(n38234) );
  NOR U51225 ( .A(n38235), .B(n38234), .Z(n44206) );
  IV U51226 ( .A(n38236), .Z(n38242) );
  IV U51227 ( .A(n38237), .Z(n38238) );
  NOR U51228 ( .A(n38242), .B(n38238), .Z(n41500) );
  IV U51229 ( .A(n38239), .Z(n38240) );
  NOR U51230 ( .A(n38240), .B(n44186), .Z(n38244) );
  IV U51231 ( .A(n38241), .Z(n38243) );
  NOR U51232 ( .A(n38243), .B(n38242), .Z(n41506) );
  NOR U51233 ( .A(n38244), .B(n41506), .Z(n40807) );
  IV U51234 ( .A(n44187), .Z(n38245) );
  NOR U51235 ( .A(n38245), .B(n44186), .Z(n41510) );
  IV U51236 ( .A(n38246), .Z(n38248) );
  NOR U51237 ( .A(n38248), .B(n38247), .Z(n44152) );
  NOR U51238 ( .A(n38250), .B(n38249), .Z(n44139) );
  IV U51239 ( .A(n38251), .Z(n38252) );
  NOR U51240 ( .A(n38253), .B(n38252), .Z(n44137) );
  IV U51241 ( .A(n38254), .Z(n38256) );
  NOR U51242 ( .A(n38256), .B(n38255), .Z(n44143) );
  NOR U51243 ( .A(n44137), .B(n44143), .Z(n40779) );
  IV U51244 ( .A(n38257), .Z(n40778) );
  IV U51245 ( .A(n38258), .Z(n38259) );
  NOR U51246 ( .A(n40778), .B(n38259), .Z(n38260) );
  IV U51247 ( .A(n38260), .Z(n44135) );
  IV U51248 ( .A(n38261), .Z(n38262) );
  NOR U51249 ( .A(n38263), .B(n38262), .Z(n44128) );
  IV U51250 ( .A(n38264), .Z(n38265) );
  NOR U51251 ( .A(n38266), .B(n38265), .Z(n40757) );
  IV U51252 ( .A(n40757), .Z(n40748) );
  IV U51253 ( .A(n38267), .Z(n38268) );
  NOR U51254 ( .A(n38269), .B(n38268), .Z(n38270) );
  IV U51255 ( .A(n38270), .Z(n44125) );
  IV U51256 ( .A(n38271), .Z(n38272) );
  NOR U51257 ( .A(n38275), .B(n38272), .Z(n40743) );
  IV U51258 ( .A(n40743), .Z(n40735) );
  IV U51259 ( .A(n38273), .Z(n38274) );
  NOR U51260 ( .A(n38275), .B(n38274), .Z(n44120) );
  IV U51261 ( .A(n38276), .Z(n38277) );
  NOR U51262 ( .A(n38278), .B(n38277), .Z(n47641) );
  IV U51263 ( .A(n38279), .Z(n38281) );
  NOR U51264 ( .A(n38281), .B(n38280), .Z(n45007) );
  NOR U51265 ( .A(n47641), .B(n45007), .Z(n44111) );
  IV U51266 ( .A(n38282), .Z(n40713) );
  NOR U51267 ( .A(n38283), .B(n40713), .Z(n40711) );
  IV U51268 ( .A(n38284), .Z(n38285) );
  NOR U51269 ( .A(n38285), .B(n40707), .Z(n41545) );
  IV U51270 ( .A(n38286), .Z(n38288) );
  IV U51271 ( .A(n38287), .Z(n40704) );
  NOR U51272 ( .A(n38288), .B(n40704), .Z(n44096) );
  IV U51273 ( .A(n38289), .Z(n44094) );
  IV U51274 ( .A(n44092), .Z(n44091) );
  XOR U51275 ( .A(n44094), .B(n44091), .Z(n38290) );
  NOR U51276 ( .A(n44096), .B(n38290), .Z(n40696) );
  IV U51277 ( .A(n38291), .Z(n38294) );
  NOR U51278 ( .A(n38292), .B(n40692), .Z(n38293) );
  IV U51279 ( .A(n38293), .Z(n38296) );
  NOR U51280 ( .A(n38294), .B(n38296), .Z(n41558) );
  IV U51281 ( .A(n38295), .Z(n38297) );
  NOR U51282 ( .A(n38297), .B(n38296), .Z(n41555) );
  IV U51283 ( .A(n38298), .Z(n38299) );
  NOR U51284 ( .A(n41567), .B(n38299), .Z(n40674) );
  NOR U51285 ( .A(n38301), .B(n38300), .Z(n45065) );
  IV U51286 ( .A(n38302), .Z(n38304) );
  IV U51287 ( .A(n38303), .Z(n40670) );
  NOR U51288 ( .A(n38304), .B(n40670), .Z(n45061) );
  NOR U51289 ( .A(n45065), .B(n45061), .Z(n44073) );
  IV U51290 ( .A(n38305), .Z(n38307) );
  NOR U51291 ( .A(n38307), .B(n38306), .Z(n41576) );
  IV U51292 ( .A(n38308), .Z(n38309) );
  NOR U51293 ( .A(n38310), .B(n38309), .Z(n44074) );
  NOR U51294 ( .A(n41576), .B(n44074), .Z(n40667) );
  IV U51295 ( .A(n38311), .Z(n38312) );
  NOR U51296 ( .A(n38313), .B(n38312), .Z(n41578) );
  IV U51297 ( .A(n38314), .Z(n38317) );
  IV U51298 ( .A(n38315), .Z(n38316) );
  NOR U51299 ( .A(n38317), .B(n38316), .Z(n44069) );
  NOR U51300 ( .A(n41578), .B(n44069), .Z(n40666) );
  IV U51301 ( .A(n38318), .Z(n38322) );
  XOR U51302 ( .A(n38328), .B(n38329), .Z(n38319) );
  NOR U51303 ( .A(n38320), .B(n38319), .Z(n38321) );
  IV U51304 ( .A(n38321), .Z(n38324) );
  NOR U51305 ( .A(n38322), .B(n38324), .Z(n44065) );
  IV U51306 ( .A(n38323), .Z(n38325) );
  NOR U51307 ( .A(n38325), .B(n38324), .Z(n44062) );
  IV U51308 ( .A(n38326), .Z(n38327) );
  NOR U51309 ( .A(n38327), .B(n38329), .Z(n44058) );
  IV U51310 ( .A(n38328), .Z(n38330) );
  NOR U51311 ( .A(n38330), .B(n38329), .Z(n44055) );
  IV U51312 ( .A(n38331), .Z(n38333) );
  NOR U51313 ( .A(n38333), .B(n38332), .Z(n41586) );
  IV U51314 ( .A(n38334), .Z(n38336) );
  NOR U51315 ( .A(n38336), .B(n38335), .Z(n41582) );
  NOR U51316 ( .A(n41586), .B(n41582), .Z(n40651) );
  IV U51317 ( .A(n38337), .Z(n38339) );
  NOR U51318 ( .A(n38339), .B(n38338), .Z(n47594) );
  IV U51319 ( .A(n38340), .Z(n38341) );
  NOR U51320 ( .A(n38342), .B(n38341), .Z(n47601) );
  NOR U51321 ( .A(n47594), .B(n47601), .Z(n41585) );
  IV U51322 ( .A(n38343), .Z(n38347) );
  IV U51323 ( .A(n38344), .Z(n40648) );
  NOR U51324 ( .A(n38345), .B(n40648), .Z(n38346) );
  IV U51325 ( .A(n38346), .Z(n38349) );
  NOR U51326 ( .A(n38347), .B(n38349), .Z(n44030) );
  IV U51327 ( .A(n38348), .Z(n38350) );
  NOR U51328 ( .A(n38350), .B(n38349), .Z(n44027) );
  IV U51329 ( .A(n38351), .Z(n38352) );
  NOR U51330 ( .A(n38353), .B(n38352), .Z(n38354) );
  IV U51331 ( .A(n38354), .Z(n40638) );
  IV U51332 ( .A(n38355), .Z(n38357) );
  NOR U51333 ( .A(n38357), .B(n38356), .Z(n47571) );
  IV U51334 ( .A(n38358), .Z(n38359) );
  NOR U51335 ( .A(n38360), .B(n38359), .Z(n45105) );
  NOR U51336 ( .A(n47571), .B(n45105), .Z(n41601) );
  IV U51337 ( .A(n38361), .Z(n38366) );
  IV U51338 ( .A(n38362), .Z(n40625) );
  NOR U51339 ( .A(n38363), .B(n40625), .Z(n38364) );
  IV U51340 ( .A(n38364), .Z(n38365) );
  NOR U51341 ( .A(n38366), .B(n38365), .Z(n52076) );
  NOR U51342 ( .A(n52080), .B(n52076), .Z(n47563) );
  IV U51343 ( .A(n38367), .Z(n38368) );
  NOR U51344 ( .A(n38368), .B(n40621), .Z(n52100) );
  IV U51345 ( .A(n38369), .Z(n38371) );
  NOR U51346 ( .A(n38371), .B(n38370), .Z(n52092) );
  NOR U51347 ( .A(n52100), .B(n52092), .Z(n50901) );
  IV U51348 ( .A(n38372), .Z(n38373) );
  NOR U51349 ( .A(n38376), .B(n38373), .Z(n44001) );
  IV U51350 ( .A(n38374), .Z(n38375) );
  NOR U51351 ( .A(n38376), .B(n38375), .Z(n43998) );
  IV U51352 ( .A(n38377), .Z(n38379) );
  IV U51353 ( .A(n38378), .Z(n40614) );
  NOR U51354 ( .A(n38379), .B(n40614), .Z(n41603) );
  IV U51355 ( .A(n38380), .Z(n38381) );
  NOR U51356 ( .A(n38382), .B(n38381), .Z(n41620) );
  IV U51357 ( .A(n38383), .Z(n38385) );
  NOR U51358 ( .A(n38385), .B(n38384), .Z(n41617) );
  NOR U51359 ( .A(n41620), .B(n41617), .Z(n40611) );
  IV U51360 ( .A(n38386), .Z(n41629) );
  IV U51361 ( .A(n38387), .Z(n38388) );
  NOR U51362 ( .A(n41629), .B(n38388), .Z(n41622) );
  NOR U51363 ( .A(n38389), .B(n43993), .Z(n38390) );
  NOR U51364 ( .A(n38391), .B(n38390), .Z(n40610) );
  IV U51365 ( .A(n38392), .Z(n38395) );
  IV U51366 ( .A(n38393), .Z(n38394) );
  NOR U51367 ( .A(n38395), .B(n38394), .Z(n38396) );
  IV U51368 ( .A(n38396), .Z(n43991) );
  IV U51369 ( .A(n38397), .Z(n38399) );
  IV U51370 ( .A(n38398), .Z(n38404) );
  NOR U51371 ( .A(n38399), .B(n38404), .Z(n41642) );
  IV U51372 ( .A(n38400), .Z(n38401) );
  NOR U51373 ( .A(n40580), .B(n38401), .Z(n41651) );
  IV U51374 ( .A(n38402), .Z(n38403) );
  NOR U51375 ( .A(n38404), .B(n38403), .Z(n41647) );
  NOR U51376 ( .A(n41651), .B(n41647), .Z(n40593) );
  IV U51377 ( .A(n38405), .Z(n38406) );
  NOR U51378 ( .A(n38407), .B(n38406), .Z(n38408) );
  IV U51379 ( .A(n38408), .Z(n40588) );
  NOR U51380 ( .A(n38409), .B(n43963), .Z(n38413) );
  IV U51381 ( .A(n38410), .Z(n40585) );
  IV U51382 ( .A(n38411), .Z(n38412) );
  NOR U51383 ( .A(n40585), .B(n38412), .Z(n41655) );
  NOR U51384 ( .A(n38413), .B(n41655), .Z(n40578) );
  IV U51385 ( .A(n38414), .Z(n38415) );
  NOR U51386 ( .A(n38416), .B(n38415), .Z(n43958) );
  IV U51387 ( .A(n38417), .Z(n38419) );
  IV U51388 ( .A(n38418), .Z(n40566) );
  NOR U51389 ( .A(n38419), .B(n40566), .Z(n41657) );
  NOR U51390 ( .A(n43958), .B(n41657), .Z(n40577) );
  IV U51391 ( .A(n38420), .Z(n38421) );
  NOR U51392 ( .A(n38421), .B(n40561), .Z(n41663) );
  NOR U51393 ( .A(n38422), .B(n40561), .Z(n41668) );
  IV U51394 ( .A(n38423), .Z(n38426) );
  IV U51395 ( .A(n38424), .Z(n38428) );
  XOR U51396 ( .A(n38428), .B(n38427), .Z(n38425) );
  NOR U51397 ( .A(n38426), .B(n38425), .Z(n43950) );
  IV U51398 ( .A(n38427), .Z(n40514) );
  NOR U51399 ( .A(n40514), .B(n38428), .Z(n38429) );
  IV U51400 ( .A(n38429), .Z(n40522) );
  IV U51401 ( .A(n38430), .Z(n38431) );
  NOR U51402 ( .A(n38431), .B(n40521), .Z(n43939) );
  IV U51403 ( .A(n38432), .Z(n38433) );
  NOR U51404 ( .A(n38434), .B(n38433), .Z(n41717) );
  NOR U51405 ( .A(n38435), .B(n41711), .Z(n41701) );
  NOR U51406 ( .A(n41717), .B(n41701), .Z(n40505) );
  IV U51407 ( .A(n38436), .Z(n38437) );
  NOR U51408 ( .A(n38438), .B(n38437), .Z(n43926) );
  IV U51409 ( .A(n38439), .Z(n38441) );
  IV U51410 ( .A(n38440), .Z(n40502) );
  NOR U51411 ( .A(n38441), .B(n40502), .Z(n43920) );
  IV U51412 ( .A(n38442), .Z(n38444) );
  NOR U51413 ( .A(n38444), .B(n38443), .Z(n40496) );
  IV U51414 ( .A(n38445), .Z(n38446) );
  NOR U51415 ( .A(n38447), .B(n38446), .Z(n43909) );
  IV U51416 ( .A(n38448), .Z(n38449) );
  NOR U51417 ( .A(n38449), .B(n40482), .Z(n43906) );
  NOR U51418 ( .A(n43909), .B(n43906), .Z(n40484) );
  IV U51419 ( .A(n38450), .Z(n38451) );
  NOR U51420 ( .A(n38452), .B(n38451), .Z(n41727) );
  IV U51421 ( .A(n38453), .Z(n38454) );
  NOR U51422 ( .A(n38455), .B(n38454), .Z(n43896) );
  IV U51423 ( .A(n38456), .Z(n38457) );
  NOR U51424 ( .A(n38458), .B(n38457), .Z(n41732) );
  NOR U51425 ( .A(n43896), .B(n41732), .Z(n40476) );
  IV U51426 ( .A(n38459), .Z(n38461) );
  NOR U51427 ( .A(n38461), .B(n38460), .Z(n43890) );
  IV U51428 ( .A(n38462), .Z(n38464) );
  NOR U51429 ( .A(n38464), .B(n38463), .Z(n43899) );
  NOR U51430 ( .A(n43890), .B(n43899), .Z(n40475) );
  IV U51431 ( .A(n38465), .Z(n38467) );
  NOR U51432 ( .A(n38467), .B(n38466), .Z(n43881) );
  NOR U51433 ( .A(n38468), .B(n43885), .Z(n38469) );
  NOR U51434 ( .A(n43881), .B(n38469), .Z(n40474) );
  IV U51435 ( .A(n38470), .Z(n38472) );
  NOR U51436 ( .A(n38472), .B(n38471), .Z(n41738) );
  IV U51437 ( .A(n38473), .Z(n38474) );
  NOR U51438 ( .A(n38475), .B(n38474), .Z(n41736) );
  NOR U51439 ( .A(n41738), .B(n41736), .Z(n40473) );
  IV U51440 ( .A(n38476), .Z(n38478) );
  NOR U51441 ( .A(n38478), .B(n38477), .Z(n38479) );
  IV U51442 ( .A(n38479), .Z(n41747) );
  IV U51443 ( .A(n38480), .Z(n38482) );
  NOR U51444 ( .A(n38482), .B(n38481), .Z(n43868) );
  IV U51445 ( .A(n38483), .Z(n38484) );
  NOR U51446 ( .A(n38485), .B(n38484), .Z(n38486) );
  NOR U51447 ( .A(n47303), .B(n38486), .Z(n45201) );
  IV U51448 ( .A(n38487), .Z(n38490) );
  IV U51449 ( .A(n40432), .Z(n38492) );
  NOR U51450 ( .A(n38488), .B(n38492), .Z(n38489) );
  IV U51451 ( .A(n38489), .Z(n40423) );
  NOR U51452 ( .A(n38490), .B(n40423), .Z(n43858) );
  IV U51453 ( .A(n38491), .Z(n40433) );
  NOR U51454 ( .A(n38492), .B(n40433), .Z(n38493) );
  IV U51455 ( .A(n38493), .Z(n40425) );
  IV U51456 ( .A(n38494), .Z(n38496) );
  IV U51457 ( .A(n38495), .Z(n38498) );
  NOR U51458 ( .A(n38496), .B(n38498), .Z(n43852) );
  IV U51459 ( .A(n38497), .Z(n38499) );
  NOR U51460 ( .A(n38499), .B(n38498), .Z(n41781) );
  IV U51461 ( .A(n38500), .Z(n38501) );
  NOR U51462 ( .A(n38501), .B(n38503), .Z(n41778) );
  IV U51463 ( .A(n38502), .Z(n38504) );
  NOR U51464 ( .A(n38504), .B(n38503), .Z(n43845) );
  IV U51465 ( .A(n38505), .Z(n38506) );
  NOR U51466 ( .A(n38507), .B(n38506), .Z(n43841) );
  IV U51467 ( .A(n38508), .Z(n38509) );
  NOR U51468 ( .A(n38509), .B(n40413), .Z(n41787) );
  NOR U51469 ( .A(n43841), .B(n41787), .Z(n40411) );
  IV U51470 ( .A(n38510), .Z(n38511) );
  NOR U51471 ( .A(n40401), .B(n38511), .Z(n41792) );
  IV U51472 ( .A(n38512), .Z(n38514) );
  NOR U51473 ( .A(n38514), .B(n38513), .Z(n43827) );
  IV U51474 ( .A(n38515), .Z(n38517) );
  NOR U51475 ( .A(n38517), .B(n38516), .Z(n41795) );
  NOR U51476 ( .A(n43827), .B(n41795), .Z(n40399) );
  IV U51477 ( .A(n38518), .Z(n38519) );
  NOR U51478 ( .A(n38520), .B(n38519), .Z(n38521) );
  IV U51479 ( .A(n38521), .Z(n40394) );
  IV U51480 ( .A(n38522), .Z(n38524) );
  NOR U51481 ( .A(n38524), .B(n38523), .Z(n41804) );
  IV U51482 ( .A(n38525), .Z(n38526) );
  NOR U51483 ( .A(n38527), .B(n38526), .Z(n41802) );
  NOR U51484 ( .A(n41804), .B(n41802), .Z(n40386) );
  IV U51485 ( .A(n38528), .Z(n38530) );
  NOR U51486 ( .A(n38530), .B(n38529), .Z(n41809) );
  IV U51487 ( .A(n38531), .Z(n38533) );
  NOR U51488 ( .A(n38533), .B(n38532), .Z(n41807) );
  NOR U51489 ( .A(n41809), .B(n41807), .Z(n40385) );
  IV U51490 ( .A(n38534), .Z(n40351) );
  IV U51491 ( .A(n38535), .Z(n38536) );
  NOR U51492 ( .A(n40351), .B(n38536), .Z(n43807) );
  NOR U51493 ( .A(n43804), .B(n43807), .Z(n40347) );
  IV U51494 ( .A(n38537), .Z(n38538) );
  NOR U51495 ( .A(n38538), .B(n38541), .Z(n43801) );
  IV U51496 ( .A(n38539), .Z(n38540) );
  NOR U51497 ( .A(n38541), .B(n38540), .Z(n41815) );
  IV U51498 ( .A(n38542), .Z(n38544) );
  NOR U51499 ( .A(n38544), .B(n38543), .Z(n43785) );
  NOR U51500 ( .A(n38545), .B(n41820), .Z(n38546) );
  NOR U51501 ( .A(n43785), .B(n38546), .Z(n40346) );
  NOR U51502 ( .A(n38547), .B(n41825), .Z(n38551) );
  IV U51503 ( .A(n38548), .Z(n38550) );
  NOR U51504 ( .A(n38550), .B(n38549), .Z(n43776) );
  NOR U51505 ( .A(n38551), .B(n43776), .Z(n40338) );
  IV U51506 ( .A(n38552), .Z(n38553) );
  NOR U51507 ( .A(n38554), .B(n38553), .Z(n43772) );
  IV U51508 ( .A(n38555), .Z(n38559) );
  IV U51509 ( .A(n38556), .Z(n38557) );
  NOR U51510 ( .A(n38559), .B(n38557), .Z(n41832) );
  NOR U51511 ( .A(n43772), .B(n41832), .Z(n40337) );
  IV U51512 ( .A(n38558), .Z(n38560) );
  NOR U51513 ( .A(n38560), .B(n38559), .Z(n41830) );
  NOR U51514 ( .A(n41834), .B(n41830), .Z(n40336) );
  IV U51515 ( .A(n38561), .Z(n38562) );
  NOR U51516 ( .A(n38563), .B(n38562), .Z(n41843) );
  NOR U51517 ( .A(n41843), .B(n41837), .Z(n40335) );
  IV U51518 ( .A(n38564), .Z(n38565) );
  NOR U51519 ( .A(n41850), .B(n38565), .Z(n41840) );
  NOR U51520 ( .A(n38566), .B(n41850), .Z(n43765) );
  NOR U51521 ( .A(n38567), .B(n41868), .Z(n41861) );
  IV U51522 ( .A(n38568), .Z(n41865) );
  IV U51523 ( .A(n38569), .Z(n40326) );
  NOR U51524 ( .A(n41865), .B(n40326), .Z(n38570) );
  NOR U51525 ( .A(n41861), .B(n38570), .Z(n40323) );
  NOR U51526 ( .A(n38571), .B(n43746), .Z(n40312) );
  IV U51527 ( .A(n38572), .Z(n38574) );
  NOR U51528 ( .A(n38574), .B(n38573), .Z(n40271) );
  IV U51529 ( .A(n40271), .Z(n40266) );
  NOR U51530 ( .A(n38576), .B(n38575), .Z(n43713) );
  IV U51531 ( .A(n38577), .Z(n38579) );
  NOR U51532 ( .A(n38579), .B(n38578), .Z(n40241) );
  IV U51533 ( .A(n40241), .Z(n40235) );
  IV U51534 ( .A(n38580), .Z(n38581) );
  NOR U51535 ( .A(n38582), .B(n38581), .Z(n41916) );
  IV U51536 ( .A(n38583), .Z(n38584) );
  NOR U51537 ( .A(n38585), .B(n38584), .Z(n41914) );
  NOR U51538 ( .A(n41916), .B(n41914), .Z(n40233) );
  IV U51539 ( .A(n38586), .Z(n38587) );
  NOR U51540 ( .A(n38588), .B(n38587), .Z(n41920) );
  IV U51541 ( .A(n38589), .Z(n38590) );
  NOR U51542 ( .A(n38594), .B(n38590), .Z(n41922) );
  NOR U51543 ( .A(n41920), .B(n41922), .Z(n40232) );
  IV U51544 ( .A(n38591), .Z(n41929) );
  NOR U51545 ( .A(n41929), .B(n38592), .Z(n38596) );
  IV U51546 ( .A(n38593), .Z(n38595) );
  NOR U51547 ( .A(n38595), .B(n38594), .Z(n41925) );
  NOR U51548 ( .A(n38596), .B(n41925), .Z(n40231) );
  IV U51549 ( .A(n38597), .Z(n38598) );
  NOR U51550 ( .A(n38598), .B(n40229), .Z(n43693) );
  IV U51551 ( .A(n38599), .Z(n38602) );
  IV U51552 ( .A(n38600), .Z(n38601) );
  NOR U51553 ( .A(n38602), .B(n38601), .Z(n41932) );
  IV U51554 ( .A(n38603), .Z(n38606) );
  IV U51555 ( .A(n38604), .Z(n38605) );
  NOR U51556 ( .A(n38606), .B(n38605), .Z(n41937) );
  NOR U51557 ( .A(n41939), .B(n41937), .Z(n40218) );
  IV U51558 ( .A(n38607), .Z(n38608) );
  NOR U51559 ( .A(n41944), .B(n38608), .Z(n43677) );
  NOR U51560 ( .A(n41944), .B(n38609), .Z(n40217) );
  IV U51561 ( .A(n38610), .Z(n38611) );
  NOR U51562 ( .A(n38611), .B(n40215), .Z(n43663) );
  IV U51563 ( .A(n38612), .Z(n38613) );
  NOR U51564 ( .A(n38614), .B(n38613), .Z(n41978) );
  IV U51565 ( .A(n38615), .Z(n38617) );
  NOR U51566 ( .A(n38617), .B(n38616), .Z(n41975) );
  NOR U51567 ( .A(n41978), .B(n41975), .Z(n40178) );
  IV U51568 ( .A(n38618), .Z(n38619) );
  NOR U51569 ( .A(n38620), .B(n38619), .Z(n41981) );
  IV U51570 ( .A(n38621), .Z(n38623) );
  NOR U51571 ( .A(n38623), .B(n38622), .Z(n43637) );
  NOR U51572 ( .A(n41981), .B(n43637), .Z(n40177) );
  IV U51573 ( .A(n38624), .Z(n38625) );
  NOR U51574 ( .A(n38625), .B(n38627), .Z(n43631) );
  IV U51575 ( .A(n38626), .Z(n38628) );
  NOR U51576 ( .A(n38628), .B(n38627), .Z(n43641) );
  NOR U51577 ( .A(n43631), .B(n43641), .Z(n40176) );
  IV U51578 ( .A(n38629), .Z(n38634) );
  IV U51579 ( .A(n38630), .Z(n38631) );
  NOR U51580 ( .A(n38634), .B(n38631), .Z(n43624) );
  IV U51581 ( .A(n38632), .Z(n38633) );
  NOR U51582 ( .A(n38634), .B(n38633), .Z(n41984) );
  IV U51583 ( .A(n38635), .Z(n38636) );
  NOR U51584 ( .A(n38637), .B(n38636), .Z(n41990) );
  NOR U51585 ( .A(n38639), .B(n38638), .Z(n40150) );
  IV U51586 ( .A(n40150), .Z(n40140) );
  IV U51587 ( .A(n38640), .Z(n38642) );
  NOR U51588 ( .A(n38642), .B(n38641), .Z(n45415) );
  NOR U51589 ( .A(n45420), .B(n45415), .Z(n42000) );
  IV U51590 ( .A(n38643), .Z(n38645) );
  NOR U51591 ( .A(n38645), .B(n38644), .Z(n42014) );
  IV U51592 ( .A(n38646), .Z(n38648) );
  NOR U51593 ( .A(n38648), .B(n38647), .Z(n43598) );
  NOR U51594 ( .A(n42014), .B(n43598), .Z(n40123) );
  NOR U51595 ( .A(n38650), .B(n38649), .Z(n42012) );
  IV U51596 ( .A(n38651), .Z(n38653) );
  NOR U51597 ( .A(n38653), .B(n38652), .Z(n42021) );
  IV U51598 ( .A(n38654), .Z(n38655) );
  NOR U51599 ( .A(n38656), .B(n38655), .Z(n43585) );
  IV U51600 ( .A(n38657), .Z(n38659) );
  NOR U51601 ( .A(n38659), .B(n38658), .Z(n43587) );
  NOR U51602 ( .A(n43585), .B(n43587), .Z(n40122) );
  IV U51603 ( .A(n42026), .Z(n38660) );
  NOR U51604 ( .A(n42025), .B(n38660), .Z(n42031) );
  IV U51605 ( .A(n38661), .Z(n42027) );
  NOR U51606 ( .A(n42025), .B(n42027), .Z(n38662) );
  NOR U51607 ( .A(n42031), .B(n38662), .Z(n40121) );
  IV U51608 ( .A(n38663), .Z(n42036) );
  NOR U51609 ( .A(n38664), .B(n42036), .Z(n38667) );
  IV U51610 ( .A(n38665), .Z(n38666) );
  NOR U51611 ( .A(n38666), .B(n38672), .Z(n43577) );
  NOR U51612 ( .A(n38667), .B(n43577), .Z(n40120) );
  IV U51613 ( .A(n38668), .Z(n38669) );
  NOR U51614 ( .A(n38670), .B(n38669), .Z(n43572) );
  IV U51615 ( .A(n38671), .Z(n38673) );
  NOR U51616 ( .A(n38673), .B(n38672), .Z(n43574) );
  NOR U51617 ( .A(n43572), .B(n43574), .Z(n40119) );
  IV U51618 ( .A(n38674), .Z(n38676) );
  NOR U51619 ( .A(n38676), .B(n38675), .Z(n43568) );
  IV U51620 ( .A(n38677), .Z(n38678) );
  NOR U51621 ( .A(n38678), .B(n40117), .Z(n43565) );
  IV U51622 ( .A(n38679), .Z(n38681) );
  NOR U51623 ( .A(n38681), .B(n38680), .Z(n38682) );
  IV U51624 ( .A(n38682), .Z(n40110) );
  IV U51625 ( .A(n38683), .Z(n38684) );
  NOR U51626 ( .A(n38684), .B(n40101), .Z(n42046) );
  IV U51627 ( .A(n38685), .Z(n38686) );
  NOR U51628 ( .A(n38686), .B(n38691), .Z(n42050) );
  IV U51629 ( .A(n38687), .Z(n38688) );
  NOR U51630 ( .A(n38697), .B(n38688), .Z(n48882) );
  IV U51631 ( .A(n38689), .Z(n38690) );
  NOR U51632 ( .A(n38691), .B(n38690), .Z(n48891) );
  NOR U51633 ( .A(n48882), .B(n48891), .Z(n43538) );
  IV U51634 ( .A(n38692), .Z(n38694) );
  NOR U51635 ( .A(n38694), .B(n38693), .Z(n42058) );
  IV U51636 ( .A(n38695), .Z(n38696) );
  NOR U51637 ( .A(n38697), .B(n38696), .Z(n42055) );
  NOR U51638 ( .A(n42058), .B(n42055), .Z(n40091) );
  IV U51639 ( .A(n38698), .Z(n38700) );
  NOR U51640 ( .A(n38700), .B(n38699), .Z(n42061) );
  NOR U51641 ( .A(n38701), .B(n42061), .Z(n40090) );
  NOR U51642 ( .A(n38703), .B(n38702), .Z(n42069) );
  IV U51643 ( .A(n38704), .Z(n38708) );
  NOR U51644 ( .A(n38706), .B(n38705), .Z(n38707) );
  IV U51645 ( .A(n38707), .Z(n38712) );
  NOR U51646 ( .A(n38708), .B(n38712), .Z(n43512) );
  NOR U51647 ( .A(n38710), .B(n38709), .Z(n42075) );
  IV U51648 ( .A(n38711), .Z(n38713) );
  NOR U51649 ( .A(n38713), .B(n38712), .Z(n43515) );
  NOR U51650 ( .A(n42075), .B(n43515), .Z(n40078) );
  IV U51651 ( .A(n38714), .Z(n38716) );
  NOR U51652 ( .A(n38716), .B(n38715), .Z(n42080) );
  IV U51653 ( .A(n38717), .Z(n38718) );
  NOR U51654 ( .A(n38718), .B(n38723), .Z(n43494) );
  IV U51655 ( .A(n38719), .Z(n38727) );
  IV U51656 ( .A(n38720), .Z(n38721) );
  NOR U51657 ( .A(n38727), .B(n38721), .Z(n46900) );
  IV U51658 ( .A(n38722), .Z(n38724) );
  NOR U51659 ( .A(n38724), .B(n38723), .Z(n45469) );
  NOR U51660 ( .A(n46900), .B(n45469), .Z(n42083) );
  IV U51661 ( .A(n38725), .Z(n38726) );
  NOR U51662 ( .A(n38727), .B(n38726), .Z(n42087) );
  IV U51663 ( .A(n38728), .Z(n38729) );
  NOR U51664 ( .A(n38730), .B(n38729), .Z(n42084) );
  IV U51665 ( .A(n38731), .Z(n38732) );
  NOR U51666 ( .A(n38732), .B(n38734), .Z(n42093) );
  IV U51667 ( .A(n38733), .Z(n38735) );
  NOR U51668 ( .A(n38735), .B(n38734), .Z(n42090) );
  IV U51669 ( .A(n38736), .Z(n38737) );
  NOR U51670 ( .A(n38738), .B(n38737), .Z(n42110) );
  IV U51671 ( .A(n38739), .Z(n38740) );
  NOR U51672 ( .A(n38740), .B(n40060), .Z(n42105) );
  NOR U51673 ( .A(n42110), .B(n42105), .Z(n40056) );
  IV U51674 ( .A(n38741), .Z(n38742) );
  NOR U51675 ( .A(n38742), .B(n38748), .Z(n38743) );
  IV U51676 ( .A(n38743), .Z(n42108) );
  IV U51677 ( .A(n38744), .Z(n42119) );
  NOR U51678 ( .A(n42119), .B(n38745), .Z(n38749) );
  IV U51679 ( .A(n38746), .Z(n38747) );
  NOR U51680 ( .A(n38748), .B(n38747), .Z(n42113) );
  NOR U51681 ( .A(n38749), .B(n42113), .Z(n40055) );
  IV U51682 ( .A(n38750), .Z(n38752) );
  NOR U51683 ( .A(n38752), .B(n38751), .Z(n42124) );
  IV U51684 ( .A(n38753), .Z(n38754) );
  NOR U51685 ( .A(n38754), .B(n42115), .Z(n42120) );
  NOR U51686 ( .A(n42124), .B(n42120), .Z(n40054) );
  IV U51687 ( .A(n38755), .Z(n38763) );
  IV U51688 ( .A(n38756), .Z(n38757) );
  NOR U51689 ( .A(n38763), .B(n38757), .Z(n42135) );
  IV U51690 ( .A(n38758), .Z(n38760) );
  NOR U51691 ( .A(n38760), .B(n38759), .Z(n42132) );
  NOR U51692 ( .A(n42135), .B(n42132), .Z(n40046) );
  IV U51693 ( .A(n38761), .Z(n38762) );
  NOR U51694 ( .A(n38763), .B(n38762), .Z(n40044) );
  IV U51695 ( .A(n40044), .Z(n40028) );
  IV U51696 ( .A(n38764), .Z(n38765) );
  NOR U51697 ( .A(n38766), .B(n38765), .Z(n42146) );
  IV U51698 ( .A(n38767), .Z(n38769) );
  NOR U51699 ( .A(n38769), .B(n38768), .Z(n43465) );
  NOR U51700 ( .A(n42146), .B(n43465), .Z(n40020) );
  IV U51701 ( .A(n38770), .Z(n38775) );
  IV U51702 ( .A(n38771), .Z(n38772) );
  NOR U51703 ( .A(n38773), .B(n38772), .Z(n38774) );
  IV U51704 ( .A(n38774), .Z(n40007) );
  NOR U51705 ( .A(n38775), .B(n40007), .Z(n42158) );
  IV U51706 ( .A(n38776), .Z(n38778) );
  NOR U51707 ( .A(n38778), .B(n38777), .Z(n42164) );
  NOR U51708 ( .A(n43449), .B(n42164), .Z(n40005) );
  IV U51709 ( .A(n38779), .Z(n38781) );
  NOR U51710 ( .A(n38781), .B(n38780), .Z(n40001) );
  IV U51711 ( .A(n39998), .Z(n45530) );
  IV U51712 ( .A(n38782), .Z(n38786) );
  NOR U51713 ( .A(n38784), .B(n38783), .Z(n38785) );
  IV U51714 ( .A(n38785), .Z(n39990) );
  NOR U51715 ( .A(n38786), .B(n39990), .Z(n42173) );
  IV U51716 ( .A(n38787), .Z(n38788) );
  NOR U51717 ( .A(n38789), .B(n38788), .Z(n42188) );
  IV U51718 ( .A(n38790), .Z(n38791) );
  NOR U51719 ( .A(n38792), .B(n38791), .Z(n42183) );
  NOR U51720 ( .A(n42188), .B(n42183), .Z(n39972) );
  IV U51721 ( .A(n38793), .Z(n38794) );
  NOR U51722 ( .A(n38794), .B(n38796), .Z(n42185) );
  IV U51723 ( .A(n38795), .Z(n38797) );
  NOR U51724 ( .A(n38797), .B(n38796), .Z(n43425) );
  IV U51725 ( .A(n38798), .Z(n38803) );
  IV U51726 ( .A(n38799), .Z(n38800) );
  NOR U51727 ( .A(n38803), .B(n38800), .Z(n43422) );
  IV U51728 ( .A(n38801), .Z(n38802) );
  NOR U51729 ( .A(n38803), .B(n38802), .Z(n43410) );
  IV U51730 ( .A(n38804), .Z(n38805) );
  NOR U51731 ( .A(n38805), .B(n38807), .Z(n42191) );
  IV U51732 ( .A(n38806), .Z(n38808) );
  NOR U51733 ( .A(n38808), .B(n38807), .Z(n43414) );
  NOR U51734 ( .A(n38809), .B(n42204), .Z(n39964) );
  IV U51735 ( .A(n38810), .Z(n38811) );
  NOR U51736 ( .A(n38812), .B(n38811), .Z(n42210) );
  IV U51737 ( .A(n38813), .Z(n38818) );
  IV U51738 ( .A(n38814), .Z(n38815) );
  NOR U51739 ( .A(n38816), .B(n38815), .Z(n38817) );
  IV U51740 ( .A(n38817), .Z(n38820) );
  NOR U51741 ( .A(n38818), .B(n38820), .Z(n42215) );
  NOR U51742 ( .A(n42210), .B(n42215), .Z(n39963) );
  IV U51743 ( .A(n38819), .Z(n38821) );
  NOR U51744 ( .A(n38821), .B(n38820), .Z(n42212) );
  IV U51745 ( .A(n38822), .Z(n38825) );
  XOR U51746 ( .A(n39957), .B(n39960), .Z(n43407) );
  NOR U51747 ( .A(n38823), .B(n43407), .Z(n38824) );
  IV U51748 ( .A(n38824), .Z(n38827) );
  NOR U51749 ( .A(n38825), .B(n38827), .Z(n42221) );
  IV U51750 ( .A(n38826), .Z(n38828) );
  NOR U51751 ( .A(n38828), .B(n38827), .Z(n42218) );
  IV U51752 ( .A(n38829), .Z(n38830) );
  NOR U51753 ( .A(n38830), .B(n39936), .Z(n38831) );
  IV U51754 ( .A(n38831), .Z(n43386) );
  NOR U51755 ( .A(n38832), .B(n43380), .Z(n38836) );
  IV U51756 ( .A(n38833), .Z(n38834) );
  NOR U51757 ( .A(n38835), .B(n38834), .Z(n43388) );
  NOR U51758 ( .A(n38836), .B(n43388), .Z(n39933) );
  IV U51759 ( .A(n38837), .Z(n39923) );
  IV U51760 ( .A(n38838), .Z(n38839) );
  NOR U51761 ( .A(n39923), .B(n38839), .Z(n38840) );
  IV U51762 ( .A(n38840), .Z(n42244) );
  IV U51763 ( .A(n38841), .Z(n38849) );
  IV U51764 ( .A(n38842), .Z(n38843) );
  NOR U51765 ( .A(n38849), .B(n38843), .Z(n43369) );
  IV U51766 ( .A(n38844), .Z(n38845) );
  NOR U51767 ( .A(n38846), .B(n38845), .Z(n42251) );
  NOR U51768 ( .A(n43369), .B(n42251), .Z(n39917) );
  IV U51769 ( .A(n38847), .Z(n38848) );
  NOR U51770 ( .A(n38849), .B(n38848), .Z(n43364) );
  IV U51771 ( .A(n38850), .Z(n38851) );
  NOR U51772 ( .A(n39915), .B(n38851), .Z(n43357) );
  NOR U51773 ( .A(n43364), .B(n43357), .Z(n39916) );
  IV U51774 ( .A(n38852), .Z(n38856) );
  NOR U51775 ( .A(n38854), .B(n38853), .Z(n38855) );
  IV U51776 ( .A(n38855), .Z(n39901) );
  NOR U51777 ( .A(n38856), .B(n39901), .Z(n45593) );
  NOR U51778 ( .A(n46701), .B(n45593), .Z(n43339) );
  IV U51779 ( .A(n38857), .Z(n38858) );
  NOR U51780 ( .A(n38858), .B(n39871), .Z(n38859) );
  IV U51781 ( .A(n38859), .Z(n42267) );
  IV U51782 ( .A(n38860), .Z(n38862) );
  NOR U51783 ( .A(n38862), .B(n38861), .Z(n43321) );
  NOR U51784 ( .A(n38864), .B(n38863), .Z(n39863) );
  IV U51785 ( .A(n39859), .Z(n39851) );
  IV U51786 ( .A(n38865), .Z(n43282) );
  NOR U51787 ( .A(n43282), .B(n38866), .Z(n39850) );
  NOR U51788 ( .A(n38868), .B(n38867), .Z(n42276) );
  IV U51789 ( .A(n38869), .Z(n38871) );
  NOR U51790 ( .A(n38871), .B(n38870), .Z(n42284) );
  IV U51791 ( .A(n38872), .Z(n38873) );
  NOR U51792 ( .A(n38873), .B(n49066), .Z(n42281) );
  NOR U51793 ( .A(n42284), .B(n42281), .Z(n39837) );
  IV U51794 ( .A(n39831), .Z(n39815) );
  IV U51795 ( .A(n38874), .Z(n38875) );
  NOR U51796 ( .A(n38875), .B(n42294), .Z(n38879) );
  NOR U51797 ( .A(n38877), .B(n38876), .Z(n38878) );
  NOR U51798 ( .A(n38879), .B(n38878), .Z(n39814) );
  IV U51799 ( .A(n38880), .Z(n42306) );
  NOR U51800 ( .A(n38881), .B(n42306), .Z(n38885) );
  IV U51801 ( .A(n38882), .Z(n38884) );
  NOR U51802 ( .A(n38884), .B(n38883), .Z(n43260) );
  NOR U51803 ( .A(n38885), .B(n43260), .Z(n39813) );
  IV U51804 ( .A(n38886), .Z(n38890) );
  NOR U51805 ( .A(n38887), .B(n39810), .Z(n38888) );
  IV U51806 ( .A(n38888), .Z(n38889) );
  NOR U51807 ( .A(n38890), .B(n38889), .Z(n42309) );
  IV U51808 ( .A(n38891), .Z(n38892) );
  NOR U51809 ( .A(n38892), .B(n38894), .Z(n39782) );
  IV U51810 ( .A(n38893), .Z(n38895) );
  NOR U51811 ( .A(n38895), .B(n38894), .Z(n39786) );
  NOR U51812 ( .A(n39782), .B(n39786), .Z(n38896) );
  IV U51813 ( .A(n38896), .Z(n39781) );
  IV U51814 ( .A(n38897), .Z(n38901) );
  NOR U51815 ( .A(n38899), .B(n38898), .Z(n38900) );
  IV U51816 ( .A(n38900), .Z(n38904) );
  NOR U51817 ( .A(n38901), .B(n38904), .Z(n38902) );
  IV U51818 ( .A(n38902), .Z(n42320) );
  IV U51819 ( .A(n38903), .Z(n38905) );
  NOR U51820 ( .A(n38905), .B(n38904), .Z(n42322) );
  IV U51821 ( .A(n38906), .Z(n38907) );
  NOR U51822 ( .A(n38907), .B(n38912), .Z(n43231) );
  NOR U51823 ( .A(n42322), .B(n43231), .Z(n39780) );
  IV U51824 ( .A(n38908), .Z(n38909) );
  NOR U51825 ( .A(n38910), .B(n38909), .Z(n42327) );
  IV U51826 ( .A(n38911), .Z(n38913) );
  NOR U51827 ( .A(n38913), .B(n38912), .Z(n43234) );
  NOR U51828 ( .A(n42327), .B(n43234), .Z(n39779) );
  IV U51829 ( .A(n38914), .Z(n38916) );
  NOR U51830 ( .A(n38916), .B(n38915), .Z(n43223) );
  IV U51831 ( .A(n38917), .Z(n38918) );
  NOR U51832 ( .A(n38919), .B(n38918), .Z(n42325) );
  NOR U51833 ( .A(n43223), .B(n42325), .Z(n39778) );
  NOR U51834 ( .A(n38920), .B(n42330), .Z(n38924) );
  IV U51835 ( .A(n38921), .Z(n38922) );
  NOR U51836 ( .A(n38923), .B(n38922), .Z(n43216) );
  NOR U51837 ( .A(n38924), .B(n43216), .Z(n39777) );
  IV U51838 ( .A(n38925), .Z(n38926) );
  NOR U51839 ( .A(n38926), .B(n38934), .Z(n42336) );
  IV U51840 ( .A(n38927), .Z(n38929) );
  NOR U51841 ( .A(n38929), .B(n38928), .Z(n42334) );
  NOR U51842 ( .A(n42336), .B(n42334), .Z(n39776) );
  IV U51843 ( .A(n38930), .Z(n38932) );
  IV U51844 ( .A(n38931), .Z(n38938) );
  NOR U51845 ( .A(n38932), .B(n38938), .Z(n43208) );
  IV U51846 ( .A(n38933), .Z(n38935) );
  NOR U51847 ( .A(n38935), .B(n38934), .Z(n43213) );
  NOR U51848 ( .A(n43208), .B(n43213), .Z(n39775) );
  IV U51849 ( .A(n38936), .Z(n38937) );
  NOR U51850 ( .A(n38938), .B(n38937), .Z(n38939) );
  IV U51851 ( .A(n38939), .Z(n43207) );
  NOR U51852 ( .A(n39772), .B(n39770), .Z(n39769) );
  IV U51853 ( .A(n38940), .Z(n38941) );
  NOR U51854 ( .A(n38941), .B(n49102), .Z(n42339) );
  IV U51855 ( .A(n38942), .Z(n38945) );
  IV U51856 ( .A(n38943), .Z(n38944) );
  NOR U51857 ( .A(n38945), .B(n38944), .Z(n38946) );
  IV U51858 ( .A(n38946), .Z(n43188) );
  IV U51859 ( .A(n38947), .Z(n38950) );
  IV U51860 ( .A(n38948), .Z(n38949) );
  NOR U51861 ( .A(n38950), .B(n38949), .Z(n43184) );
  NOR U51862 ( .A(n43181), .B(n43184), .Z(n39759) );
  IV U51863 ( .A(n38951), .Z(n43179) );
  IV U51864 ( .A(n38952), .Z(n38953) );
  NOR U51865 ( .A(n38954), .B(n38953), .Z(n49937) );
  NOR U51866 ( .A(n49937), .B(n43177), .Z(n39758) );
  IV U51867 ( .A(n38955), .Z(n38956) );
  NOR U51868 ( .A(n38961), .B(n38956), .Z(n43162) );
  IV U51869 ( .A(n38957), .Z(n38958) );
  NOR U51870 ( .A(n38959), .B(n38958), .Z(n42350) );
  IV U51871 ( .A(n38960), .Z(n38962) );
  NOR U51872 ( .A(n38962), .B(n38961), .Z(n43158) );
  NOR U51873 ( .A(n42350), .B(n43158), .Z(n39737) );
  NOR U51874 ( .A(n38963), .B(n42369), .Z(n42360) );
  IV U51875 ( .A(n38964), .Z(n38966) );
  NOR U51876 ( .A(n38966), .B(n38965), .Z(n42367) );
  NOR U51877 ( .A(n38968), .B(n38967), .Z(n42376) );
  NOR U51878 ( .A(n42367), .B(n42376), .Z(n39725) );
  IV U51879 ( .A(n38969), .Z(n38971) );
  NOR U51880 ( .A(n38971), .B(n38970), .Z(n43135) );
  IV U51881 ( .A(n38972), .Z(n38974) );
  NOR U51882 ( .A(n38974), .B(n38973), .Z(n43152) );
  NOR U51883 ( .A(n43135), .B(n43152), .Z(n39724) );
  NOR U51884 ( .A(n38976), .B(n38975), .Z(n43139) );
  NOR U51885 ( .A(n38977), .B(n42385), .Z(n42379) );
  IV U51886 ( .A(n38978), .Z(n38980) );
  NOR U51887 ( .A(n38980), .B(n38979), .Z(n43100) );
  NOR U51888 ( .A(n38981), .B(n49193), .Z(n43112) );
  NOR U51889 ( .A(n43100), .B(n43112), .Z(n39683) );
  IV U51890 ( .A(n38982), .Z(n42393) );
  NOR U51891 ( .A(n38984), .B(n38983), .Z(n42397) );
  IV U51892 ( .A(n38985), .Z(n38987) );
  NOR U51893 ( .A(n38987), .B(n38986), .Z(n42400) );
  NOR U51894 ( .A(n42400), .B(n42394), .Z(n39681) );
  IV U51895 ( .A(n38988), .Z(n38993) );
  IV U51896 ( .A(n38989), .Z(n38990) );
  NOR U51897 ( .A(n38993), .B(n38990), .Z(n39677) );
  IV U51898 ( .A(n38991), .Z(n38992) );
  NOR U51899 ( .A(n38993), .B(n38992), .Z(n39674) );
  IV U51900 ( .A(n39674), .Z(n39669) );
  IV U51901 ( .A(n38994), .Z(n38995) );
  NOR U51902 ( .A(n38995), .B(n39666), .Z(n43091) );
  IV U51903 ( .A(n38996), .Z(n38999) );
  NOR U51904 ( .A(n38997), .B(n38999), .Z(n42421) );
  IV U51905 ( .A(n38998), .Z(n39000) );
  NOR U51906 ( .A(n39000), .B(n38999), .Z(n42419) );
  NOR U51907 ( .A(n42421), .B(n42419), .Z(n39651) );
  NOR U51908 ( .A(n39002), .B(n39001), .Z(n42426) );
  IV U51909 ( .A(n39003), .Z(n39006) );
  IV U51910 ( .A(n39004), .Z(n39005) );
  NOR U51911 ( .A(n39006), .B(n39005), .Z(n42429) );
  IV U51912 ( .A(n39007), .Z(n39008) );
  NOR U51913 ( .A(n39008), .B(n39013), .Z(n42435) );
  IV U51914 ( .A(n39009), .Z(n39010) );
  NOR U51915 ( .A(n39011), .B(n39010), .Z(n43078) );
  NOR U51916 ( .A(n39013), .B(n39012), .Z(n42438) );
  NOR U51917 ( .A(n43078), .B(n42438), .Z(n39644) );
  IV U51918 ( .A(n39014), .Z(n39015) );
  NOR U51919 ( .A(n39016), .B(n39015), .Z(n43074) );
  IV U51920 ( .A(n39017), .Z(n39018) );
  NOR U51921 ( .A(n39019), .B(n39018), .Z(n53035) );
  IV U51922 ( .A(n39020), .Z(n39021) );
  NOR U51923 ( .A(n39643), .B(n39021), .Z(n53027) );
  NOR U51924 ( .A(n53035), .B(n53027), .Z(n49252) );
  NOR U51925 ( .A(n39023), .B(n39022), .Z(n43048) );
  IV U51926 ( .A(n39024), .Z(n39025) );
  NOR U51927 ( .A(n39026), .B(n39025), .Z(n45775) );
  NOR U51928 ( .A(n45782), .B(n45775), .Z(n43036) );
  IV U51929 ( .A(n39027), .Z(n39028) );
  NOR U51930 ( .A(n39031), .B(n39028), .Z(n42463) );
  IV U51931 ( .A(n39029), .Z(n39030) );
  NOR U51932 ( .A(n39031), .B(n39030), .Z(n39032) );
  IV U51933 ( .A(n39032), .Z(n42462) );
  IV U51934 ( .A(n39033), .Z(n39034) );
  NOR U51935 ( .A(n39035), .B(n39034), .Z(n42469) );
  IV U51936 ( .A(n39036), .Z(n39038) );
  NOR U51937 ( .A(n39038), .B(n39037), .Z(n42466) );
  NOR U51938 ( .A(n42469), .B(n42466), .Z(n39604) );
  IV U51939 ( .A(n39039), .Z(n42473) );
  NOR U51940 ( .A(n42473), .B(n39040), .Z(n39603) );
  IV U51941 ( .A(n39041), .Z(n39042) );
  NOR U51942 ( .A(n39042), .B(n39586), .Z(n43029) );
  IV U51943 ( .A(n39043), .Z(n39044) );
  NOR U51944 ( .A(n39044), .B(n39586), .Z(n42479) );
  NOR U51945 ( .A(n43029), .B(n42479), .Z(n39602) );
  IV U51946 ( .A(n39045), .Z(n39046) );
  NOR U51947 ( .A(n39047), .B(n39046), .Z(n42482) );
  IV U51948 ( .A(n39048), .Z(n39049) );
  NOR U51949 ( .A(n39049), .B(n39054), .Z(n39592) );
  NOR U51950 ( .A(n42482), .B(n39592), .Z(n39584) );
  IV U51951 ( .A(n39050), .Z(n39051) );
  NOR U51952 ( .A(n39052), .B(n39051), .Z(n42491) );
  IV U51953 ( .A(n39053), .Z(n39055) );
  NOR U51954 ( .A(n39055), .B(n39054), .Z(n42486) );
  NOR U51955 ( .A(n42491), .B(n42486), .Z(n39583) );
  IV U51956 ( .A(n39056), .Z(n39058) );
  NOR U51957 ( .A(n39058), .B(n39057), .Z(n39059) );
  IV U51958 ( .A(n39059), .Z(n39574) );
  NOR U51959 ( .A(n39061), .B(n39060), .Z(n42512) );
  NOR U51960 ( .A(n42512), .B(n42507), .Z(n39565) );
  IV U51961 ( .A(n39062), .Z(n39063) );
  NOR U51962 ( .A(n39063), .B(n39556), .Z(n43011) );
  IV U51963 ( .A(n39064), .Z(n39065) );
  NOR U51964 ( .A(n39065), .B(n39070), .Z(n43008) );
  IV U51965 ( .A(n39066), .Z(n39068) );
  NOR U51966 ( .A(n39068), .B(n39067), .Z(n42515) );
  NOR U51967 ( .A(n43008), .B(n42515), .Z(n39552) );
  IV U51968 ( .A(n39069), .Z(n39071) );
  NOR U51969 ( .A(n39071), .B(n39070), .Z(n42517) );
  IV U51970 ( .A(n39072), .Z(n39073) );
  NOR U51971 ( .A(n39073), .B(n39081), .Z(n42524) );
  IV U51972 ( .A(n39074), .Z(n39076) );
  NOR U51973 ( .A(n39076), .B(n39075), .Z(n42521) );
  NOR U51974 ( .A(n42524), .B(n42521), .Z(n39551) );
  IV U51975 ( .A(n39077), .Z(n39079) );
  NOR U51976 ( .A(n39079), .B(n39078), .Z(n42998) );
  IV U51977 ( .A(n39080), .Z(n39082) );
  NOR U51978 ( .A(n39082), .B(n39081), .Z(n43000) );
  NOR U51979 ( .A(n42998), .B(n43000), .Z(n39550) );
  IV U51980 ( .A(n39083), .Z(n39088) );
  IV U51981 ( .A(n39084), .Z(n39085) );
  NOR U51982 ( .A(n39088), .B(n39085), .Z(n42535) );
  IV U51983 ( .A(n39086), .Z(n39087) );
  NOR U51984 ( .A(n39088), .B(n39087), .Z(n42532) );
  NOR U51985 ( .A(n42535), .B(n42532), .Z(n39542) );
  IV U51986 ( .A(n39089), .Z(n39090) );
  NOR U51987 ( .A(n39090), .B(n39535), .Z(n42537) );
  IV U51988 ( .A(n39091), .Z(n39093) );
  IV U51989 ( .A(n39092), .Z(n39529) );
  NOR U51990 ( .A(n39093), .B(n39529), .Z(n42981) );
  IV U51991 ( .A(n39094), .Z(n39095) );
  NOR U51992 ( .A(n39095), .B(n39097), .Z(n42978) );
  IV U51993 ( .A(n39096), .Z(n39098) );
  NOR U51994 ( .A(n39098), .B(n39097), .Z(n42548) );
  IV U51995 ( .A(n39099), .Z(n39101) );
  IV U51996 ( .A(n39100), .Z(n39103) );
  NOR U51997 ( .A(n39101), .B(n39103), .Z(n42545) );
  IV U51998 ( .A(n39102), .Z(n39104) );
  NOR U51999 ( .A(n39104), .B(n39103), .Z(n42974) );
  IV U52000 ( .A(n39105), .Z(n39108) );
  NOR U52001 ( .A(n39515), .B(n39106), .Z(n39107) );
  IV U52002 ( .A(n39107), .Z(n39522) );
  NOR U52003 ( .A(n39108), .B(n39522), .Z(n42970) );
  NOR U52004 ( .A(n42974), .B(n42970), .Z(n39524) );
  IV U52005 ( .A(n39109), .Z(n39110) );
  NOR U52006 ( .A(n39517), .B(n39110), .Z(n42553) );
  IV U52007 ( .A(n39111), .Z(n39113) );
  NOR U52008 ( .A(n39113), .B(n39112), .Z(n46236) );
  IV U52009 ( .A(n39114), .Z(n39115) );
  NOR U52010 ( .A(n39115), .B(n39510), .Z(n46246) );
  NOR U52011 ( .A(n46236), .B(n46246), .Z(n42565) );
  IV U52012 ( .A(n39116), .Z(n39118) );
  IV U52013 ( .A(n39117), .Z(n39471) );
  NOR U52014 ( .A(n39118), .B(n39471), .Z(n42918) );
  IV U52015 ( .A(n39119), .Z(n39122) );
  NOR U52016 ( .A(n39120), .B(n39123), .Z(n39121) );
  IV U52017 ( .A(n39121), .Z(n39427) );
  NOR U52018 ( .A(n39122), .B(n39427), .Z(n42878) );
  NOR U52019 ( .A(n39124), .B(n39123), .Z(n39125) );
  IV U52020 ( .A(n39125), .Z(n39130) );
  NOR U52021 ( .A(n39126), .B(n39130), .Z(n42614) );
  IV U52022 ( .A(n39127), .Z(n39128) );
  NOR U52023 ( .A(n39129), .B(n39128), .Z(n42616) );
  NOR U52024 ( .A(n39131), .B(n39130), .Z(n42881) );
  NOR U52025 ( .A(n42616), .B(n42881), .Z(n39424) );
  IV U52026 ( .A(n39132), .Z(n39136) );
  IV U52027 ( .A(n39133), .Z(n39416) );
  NOR U52028 ( .A(n39134), .B(n39416), .Z(n39135) );
  IV U52029 ( .A(n39135), .Z(n39421) );
  NOR U52030 ( .A(n39136), .B(n39421), .Z(n42618) );
  IV U52031 ( .A(n39137), .Z(n39139) );
  NOR U52032 ( .A(n39139), .B(n39138), .Z(n45901) );
  IV U52033 ( .A(n39140), .Z(n39142) );
  NOR U52034 ( .A(n39142), .B(n39141), .Z(n45896) );
  NOR U52035 ( .A(n45901), .B(n45896), .Z(n42865) );
  IV U52036 ( .A(n39143), .Z(n39146) );
  NOR U52037 ( .A(n39144), .B(n39151), .Z(n39145) );
  IV U52038 ( .A(n39145), .Z(n39148) );
  NOR U52039 ( .A(n39146), .B(n39148), .Z(n42844) );
  IV U52040 ( .A(n39147), .Z(n39149) );
  NOR U52041 ( .A(n39149), .B(n39148), .Z(n42841) );
  IV U52042 ( .A(n39150), .Z(n39152) );
  NOR U52043 ( .A(n39152), .B(n39151), .Z(n39153) );
  IV U52044 ( .A(n39153), .Z(n39403) );
  IV U52045 ( .A(n39154), .Z(n39156) );
  IV U52046 ( .A(n39155), .Z(n39386) );
  NOR U52047 ( .A(n39156), .B(n39386), .Z(n42641) );
  IV U52048 ( .A(n39157), .Z(n39158) );
  NOR U52049 ( .A(n39158), .B(n39162), .Z(n42638) );
  IV U52050 ( .A(n42646), .Z(n39167) );
  IV U52051 ( .A(n39159), .Z(n42649) );
  NOR U52052 ( .A(n39167), .B(n42649), .Z(n39163) );
  IV U52053 ( .A(n39160), .Z(n39161) );
  NOR U52054 ( .A(n39162), .B(n39161), .Z(n42644) );
  NOR U52055 ( .A(n39163), .B(n42644), .Z(n39383) );
  IV U52056 ( .A(n39164), .Z(n39165) );
  NOR U52057 ( .A(n39165), .B(n39374), .Z(n42817) );
  IV U52058 ( .A(n39166), .Z(n42647) );
  NOR U52059 ( .A(n42647), .B(n39167), .Z(n42654) );
  NOR U52060 ( .A(n42817), .B(n42654), .Z(n39382) );
  IV U52061 ( .A(n39168), .Z(n39378) );
  IV U52062 ( .A(n39169), .Z(n39170) );
  NOR U52063 ( .A(n39378), .B(n39170), .Z(n42810) );
  IV U52064 ( .A(n39171), .Z(n39174) );
  NOR U52065 ( .A(n39187), .B(n39172), .Z(n39173) );
  IV U52066 ( .A(n39173), .Z(n39176) );
  NOR U52067 ( .A(n39174), .B(n39176), .Z(n42807) );
  IV U52068 ( .A(n39175), .Z(n39177) );
  NOR U52069 ( .A(n39177), .B(n39176), .Z(n39178) );
  IV U52070 ( .A(n39178), .Z(n42798) );
  IV U52071 ( .A(n39179), .Z(n39181) );
  NOR U52072 ( .A(n39181), .B(n39180), .Z(n42656) );
  IV U52073 ( .A(n39182), .Z(n39183) );
  NOR U52074 ( .A(n39184), .B(n39183), .Z(n42794) );
  NOR U52075 ( .A(n42656), .B(n42794), .Z(n39369) );
  IV U52076 ( .A(n39185), .Z(n39186) );
  NOR U52077 ( .A(n39187), .B(n39186), .Z(n42790) );
  IV U52078 ( .A(n39188), .Z(n39189) );
  NOR U52079 ( .A(n39354), .B(n39189), .Z(n42659) );
  NOR U52080 ( .A(n42790), .B(n42659), .Z(n39368) );
  IV U52081 ( .A(n39190), .Z(n39191) );
  NOR U52082 ( .A(n39192), .B(n39191), .Z(n39193) );
  IV U52083 ( .A(n39193), .Z(n42662) );
  IV U52084 ( .A(n39194), .Z(n39198) );
  IV U52085 ( .A(n39195), .Z(n39196) );
  NOR U52086 ( .A(n39198), .B(n39196), .Z(n42784) );
  IV U52087 ( .A(n39197), .Z(n39199) );
  NOR U52088 ( .A(n39199), .B(n39198), .Z(n39200) );
  IV U52089 ( .A(n39200), .Z(n42783) );
  NOR U52090 ( .A(n39201), .B(n39344), .Z(n39340) );
  IV U52091 ( .A(n39202), .Z(n39204) );
  NOR U52092 ( .A(n39204), .B(n39203), .Z(n42773) );
  IV U52093 ( .A(n39205), .Z(n39206) );
  NOR U52094 ( .A(n39206), .B(n39303), .Z(n42751) );
  IV U52095 ( .A(n39207), .Z(n42673) );
  NOR U52096 ( .A(n42673), .B(n39208), .Z(n39305) );
  IV U52097 ( .A(n39209), .Z(n39211) );
  NOR U52098 ( .A(n39211), .B(n39210), .Z(n39212) );
  IV U52099 ( .A(n39212), .Z(n39296) );
  NOR U52100 ( .A(n39214), .B(n39213), .Z(n42744) );
  IV U52101 ( .A(n39215), .Z(n39216) );
  NOR U52102 ( .A(n39280), .B(n39216), .Z(n42733) );
  IV U52103 ( .A(n39217), .Z(n39219) );
  NOR U52104 ( .A(n39219), .B(n39218), .Z(n42689) );
  NOR U52105 ( .A(n39220), .B(n42686), .Z(n39221) );
  NOR U52106 ( .A(n42689), .B(n39221), .Z(n39278) );
  IV U52107 ( .A(n39222), .Z(n39223) );
  NOR U52108 ( .A(n39224), .B(n39223), .Z(n42699) );
  IV U52109 ( .A(n39225), .Z(n39226) );
  NOR U52110 ( .A(n39227), .B(n39226), .Z(n42704) );
  NOR U52111 ( .A(n42699), .B(n42704), .Z(n39270) );
  IV U52112 ( .A(n39228), .Z(n39229) );
  NOR U52113 ( .A(n39230), .B(n39229), .Z(n42717) );
  IV U52114 ( .A(n39231), .Z(n39232) );
  NOR U52115 ( .A(n39233), .B(n39232), .Z(n39242) );
  NOR U52116 ( .A(n39235), .B(n39234), .Z(n39236) );
  NOR U52117 ( .A(n39237), .B(n39236), .Z(n39238) );
  NOR U52118 ( .A(n39239), .B(n39238), .Z(n39240) );
  IV U52119 ( .A(n39240), .Z(n39241) );
  NOR U52120 ( .A(n39242), .B(n39241), .Z(n42715) );
  IV U52121 ( .A(n42715), .Z(n42712) );
  IV U52122 ( .A(n39243), .Z(n39245) );
  NOR U52123 ( .A(n39245), .B(n39244), .Z(n42713) );
  IV U52124 ( .A(n42713), .Z(n42714) );
  XOR U52125 ( .A(n42712), .B(n42714), .Z(n39246) );
  XOR U52126 ( .A(n42717), .B(n39246), .Z(n42724) );
  IV U52127 ( .A(n39247), .Z(n39249) );
  NOR U52128 ( .A(n39249), .B(n39248), .Z(n42716) );
  IV U52129 ( .A(n39250), .Z(n39251) );
  NOR U52130 ( .A(n39251), .B(n39258), .Z(n42723) );
  NOR U52131 ( .A(n42716), .B(n42723), .Z(n39252) );
  XOR U52132 ( .A(n42724), .B(n39252), .Z(n39253) );
  IV U52133 ( .A(n39253), .Z(n42709) );
  IV U52134 ( .A(n39260), .Z(n39255) );
  NOR U52135 ( .A(n39255), .B(n39254), .Z(n39256) );
  IV U52136 ( .A(n39256), .Z(n39265) );
  NOR U52137 ( .A(n42709), .B(n39265), .Z(n42710) );
  IV U52138 ( .A(n39257), .Z(n39259) );
  NOR U52139 ( .A(n39259), .B(n39258), .Z(n42707) );
  XOR U52140 ( .A(n42707), .B(n42709), .Z(n42703) );
  NOR U52141 ( .A(n39261), .B(n39260), .Z(n39264) );
  IV U52142 ( .A(n39262), .Z(n39263) );
  NOR U52143 ( .A(n39264), .B(n39263), .Z(n39266) );
  IV U52144 ( .A(n39266), .Z(n42702) );
  XOR U52145 ( .A(n42703), .B(n42702), .Z(n39268) );
  NOR U52146 ( .A(n39266), .B(n39265), .Z(n39267) );
  NOR U52147 ( .A(n39268), .B(n39267), .Z(n39269) );
  NOR U52148 ( .A(n42710), .B(n39269), .Z(n42700) );
  XOR U52149 ( .A(n39270), .B(n42700), .Z(n42695) );
  IV U52150 ( .A(n39271), .Z(n39272) );
  NOR U52151 ( .A(n39273), .B(n39272), .Z(n42692) );
  IV U52152 ( .A(n39274), .Z(n39275) );
  NOR U52153 ( .A(n39276), .B(n39275), .Z(n42694) );
  NOR U52154 ( .A(n42692), .B(n42694), .Z(n39277) );
  XOR U52155 ( .A(n42695), .B(n39277), .Z(n42684) );
  XOR U52156 ( .A(n39278), .B(n42684), .Z(n42735) );
  XOR U52157 ( .A(n42733), .B(n42735), .Z(n42738) );
  IV U52158 ( .A(n39279), .Z(n39283) );
  NOR U52159 ( .A(n39281), .B(n39280), .Z(n39282) );
  IV U52160 ( .A(n39282), .Z(n39285) );
  NOR U52161 ( .A(n39283), .B(n39285), .Z(n42736) );
  XOR U52162 ( .A(n42738), .B(n42736), .Z(n42743) );
  IV U52163 ( .A(n39284), .Z(n39286) );
  NOR U52164 ( .A(n39286), .B(n39285), .Z(n42741) );
  NOR U52165 ( .A(n42680), .B(n42741), .Z(n39287) );
  XOR U52166 ( .A(n42743), .B(n39287), .Z(n39288) );
  IV U52167 ( .A(n39288), .Z(n42746) );
  XOR U52168 ( .A(n42744), .B(n42746), .Z(n42748) );
  NOR U52169 ( .A(n39296), .B(n42748), .Z(n45965) );
  IV U52170 ( .A(n39289), .Z(n39290) );
  NOR U52171 ( .A(n39291), .B(n39290), .Z(n39292) );
  IV U52172 ( .A(n39292), .Z(n42679) );
  IV U52173 ( .A(n39293), .Z(n39295) );
  NOR U52174 ( .A(n39295), .B(n39294), .Z(n42747) );
  XOR U52175 ( .A(n42747), .B(n42748), .Z(n42678) );
  XOR U52176 ( .A(n42679), .B(n42678), .Z(n39299) );
  IV U52177 ( .A(n42678), .Z(n39297) );
  NOR U52178 ( .A(n39297), .B(n39296), .Z(n39298) );
  NOR U52179 ( .A(n39299), .B(n39298), .Z(n39300) );
  NOR U52180 ( .A(n45965), .B(n39300), .Z(n42672) );
  IV U52181 ( .A(n39301), .Z(n39302) );
  NOR U52182 ( .A(n39303), .B(n39302), .Z(n39304) );
  IV U52183 ( .A(n39304), .Z(n42676) );
  XOR U52184 ( .A(n42672), .B(n42676), .Z(n42753) );
  XOR U52185 ( .A(n39305), .B(n42753), .Z(n39306) );
  XOR U52186 ( .A(n42751), .B(n39306), .Z(n42759) );
  IV U52187 ( .A(n39307), .Z(n39308) );
  NOR U52188 ( .A(n42673), .B(n39308), .Z(n42669) );
  IV U52189 ( .A(n39309), .Z(n39311) );
  NOR U52190 ( .A(n39311), .B(n39310), .Z(n42666) );
  NOR U52191 ( .A(n42758), .B(n42666), .Z(n39312) );
  XOR U52192 ( .A(n42669), .B(n39312), .Z(n39313) );
  XOR U52193 ( .A(n42759), .B(n39313), .Z(n42765) );
  IV U52194 ( .A(n39314), .Z(n39316) );
  NOR U52195 ( .A(n39316), .B(n39315), .Z(n42769) );
  NOR U52196 ( .A(n42766), .B(n42769), .Z(n39317) );
  XOR U52197 ( .A(n42765), .B(n39317), .Z(n42776) );
  XOR U52198 ( .A(n42773), .B(n42776), .Z(n42664) );
  IV U52199 ( .A(n39318), .Z(n39320) );
  NOR U52200 ( .A(n39320), .B(n39319), .Z(n42775) );
  IV U52201 ( .A(n39323), .Z(n39321) );
  NOR U52202 ( .A(n39321), .B(n39332), .Z(n42663) );
  NOR U52203 ( .A(n42775), .B(n42663), .Z(n39322) );
  XOR U52204 ( .A(n42664), .B(n39322), .Z(n39334) );
  IV U52205 ( .A(n39334), .Z(n39325) );
  XOR U52206 ( .A(n39323), .B(n39332), .Z(n39324) );
  NOR U52207 ( .A(n39325), .B(n39324), .Z(n39326) );
  IV U52208 ( .A(n39326), .Z(n39331) );
  NOR U52209 ( .A(n39328), .B(n39331), .Z(n45950) );
  IV U52210 ( .A(n39327), .Z(n39329) );
  NOR U52211 ( .A(n39329), .B(n39328), .Z(n39337) );
  IV U52212 ( .A(n39330), .Z(n39333) );
  NOR U52213 ( .A(n39333), .B(n39331), .Z(n45955) );
  NOR U52214 ( .A(n39333), .B(n39332), .Z(n39335) );
  NOR U52215 ( .A(n39335), .B(n39334), .Z(n39336) );
  NOR U52216 ( .A(n45955), .B(n39336), .Z(n39342) );
  NOR U52217 ( .A(n39337), .B(n39342), .Z(n39338) );
  NOR U52218 ( .A(n45950), .B(n39338), .Z(n39339) );
  NOR U52219 ( .A(n39340), .B(n39339), .Z(n39352) );
  IV U52220 ( .A(n39341), .Z(n39346) );
  IV U52221 ( .A(n39342), .Z(n39343) );
  NOR U52222 ( .A(n39344), .B(n39343), .Z(n39345) );
  IV U52223 ( .A(n39345), .Z(n39348) );
  NOR U52224 ( .A(n39346), .B(n39348), .Z(n46050) );
  IV U52225 ( .A(n39347), .Z(n39349) );
  NOR U52226 ( .A(n39349), .B(n39348), .Z(n46047) );
  NOR U52227 ( .A(n46050), .B(n46047), .Z(n39350) );
  IV U52228 ( .A(n39350), .Z(n39351) );
  NOR U52229 ( .A(n39352), .B(n39351), .Z(n42781) );
  XOR U52230 ( .A(n42783), .B(n42781), .Z(n42785) );
  XOR U52231 ( .A(n42784), .B(n42785), .Z(n42661) );
  XOR U52232 ( .A(n42662), .B(n42661), .Z(n39362) );
  IV U52233 ( .A(n39362), .Z(n39357) );
  IV U52234 ( .A(n39353), .Z(n39355) );
  NOR U52235 ( .A(n39355), .B(n39354), .Z(n39366) );
  IV U52236 ( .A(n39366), .Z(n39356) );
  NOR U52237 ( .A(n39357), .B(n39356), .Z(n45943) );
  IV U52238 ( .A(n39358), .Z(n39359) );
  NOR U52239 ( .A(n39360), .B(n39359), .Z(n39363) );
  IV U52240 ( .A(n39363), .Z(n39361) );
  NOR U52241 ( .A(n39361), .B(n42661), .Z(n46065) );
  NOR U52242 ( .A(n39363), .B(n39362), .Z(n39364) );
  NOR U52243 ( .A(n46065), .B(n39364), .Z(n39365) );
  NOR U52244 ( .A(n39366), .B(n39365), .Z(n39367) );
  NOR U52245 ( .A(n45943), .B(n39367), .Z(n42658) );
  XOR U52246 ( .A(n39368), .B(n42658), .Z(n42796) );
  XOR U52247 ( .A(n39369), .B(n42796), .Z(n42797) );
  XOR U52248 ( .A(n42798), .B(n42797), .Z(n42809) );
  XOR U52249 ( .A(n42807), .B(n42809), .Z(n42812) );
  XOR U52250 ( .A(n42810), .B(n42812), .Z(n42821) );
  IV U52251 ( .A(n39370), .Z(n39372) );
  NOR U52252 ( .A(n39372), .B(n39371), .Z(n42801) );
  IV U52253 ( .A(n39373), .Z(n39375) );
  NOR U52254 ( .A(n39375), .B(n39374), .Z(n42820) );
  IV U52255 ( .A(n39376), .Z(n39377) );
  NOR U52256 ( .A(n39378), .B(n39377), .Z(n42804) );
  NOR U52257 ( .A(n42820), .B(n42804), .Z(n39379) );
  IV U52258 ( .A(n39379), .Z(n39380) );
  NOR U52259 ( .A(n42801), .B(n39380), .Z(n39381) );
  XOR U52260 ( .A(n42821), .B(n39381), .Z(n42653) );
  XOR U52261 ( .A(n39382), .B(n42653), .Z(n42648) );
  XOR U52262 ( .A(n39383), .B(n42648), .Z(n39384) );
  IV U52263 ( .A(n39384), .Z(n42640) );
  XOR U52264 ( .A(n42638), .B(n42640), .Z(n42642) );
  XOR U52265 ( .A(n42641), .B(n42642), .Z(n42826) );
  IV U52266 ( .A(n39385), .Z(n39387) );
  NOR U52267 ( .A(n39387), .B(n39386), .Z(n39388) );
  IV U52268 ( .A(n39388), .Z(n42825) );
  XOR U52269 ( .A(n42826), .B(n42825), .Z(n42828) );
  IV U52270 ( .A(n39389), .Z(n39390) );
  NOR U52271 ( .A(n39391), .B(n39390), .Z(n42827) );
  IV U52272 ( .A(n39392), .Z(n39394) );
  NOR U52273 ( .A(n39394), .B(n39393), .Z(n42831) );
  NOR U52274 ( .A(n42827), .B(n42831), .Z(n39395) );
  XOR U52275 ( .A(n42828), .B(n39395), .Z(n42835) );
  NOR U52276 ( .A(n39403), .B(n42835), .Z(n45910) );
  IV U52277 ( .A(n39396), .Z(n39398) );
  NOR U52278 ( .A(n39398), .B(n39397), .Z(n39399) );
  IV U52279 ( .A(n39399), .Z(n42636) );
  IV U52280 ( .A(n39400), .Z(n39402) );
  NOR U52281 ( .A(n39402), .B(n39401), .Z(n42834) );
  XOR U52282 ( .A(n42834), .B(n42835), .Z(n42635) );
  XOR U52283 ( .A(n42636), .B(n42635), .Z(n39406) );
  IV U52284 ( .A(n42635), .Z(n39404) );
  NOR U52285 ( .A(n39404), .B(n39403), .Z(n39405) );
  NOR U52286 ( .A(n39406), .B(n39405), .Z(n39407) );
  NOR U52287 ( .A(n45910), .B(n39407), .Z(n39408) );
  IV U52288 ( .A(n39408), .Z(n42842) );
  XOR U52289 ( .A(n42841), .B(n42842), .Z(n42845) );
  XOR U52290 ( .A(n42844), .B(n42845), .Z(n42857) );
  XOR U52291 ( .A(n42856), .B(n42857), .Z(n42849) );
  XOR U52292 ( .A(n42848), .B(n42849), .Z(n42853) );
  XOR U52293 ( .A(n42852), .B(n42853), .Z(n42632) );
  IV U52294 ( .A(n39409), .Z(n39410) );
  NOR U52295 ( .A(n39411), .B(n39410), .Z(n42631) );
  NOR U52296 ( .A(n39412), .B(n42624), .Z(n39413) );
  NOR U52297 ( .A(n42631), .B(n39413), .Z(n39414) );
  XOR U52298 ( .A(n42632), .B(n39414), .Z(n42864) );
  XOR U52299 ( .A(n42865), .B(n42864), .Z(n42874) );
  IV U52300 ( .A(n39415), .Z(n39417) );
  NOR U52301 ( .A(n39417), .B(n39416), .Z(n42872) );
  NOR U52302 ( .A(n42872), .B(n39418), .Z(n39419) );
  XOR U52303 ( .A(n42874), .B(n39419), .Z(n42615) );
  IV U52304 ( .A(n39420), .Z(n39422) );
  NOR U52305 ( .A(n39422), .B(n39421), .Z(n39423) );
  IV U52306 ( .A(n39423), .Z(n42870) );
  XOR U52307 ( .A(n42615), .B(n42870), .Z(n42619) );
  XOR U52308 ( .A(n42618), .B(n42619), .Z(n42883) );
  XOR U52309 ( .A(n39424), .B(n42883), .Z(n39425) );
  IV U52310 ( .A(n39425), .Z(n42885) );
  XOR U52311 ( .A(n42614), .B(n42885), .Z(n42879) );
  XOR U52312 ( .A(n42878), .B(n42879), .Z(n42613) );
  IV U52313 ( .A(n39426), .Z(n39428) );
  NOR U52314 ( .A(n39428), .B(n39427), .Z(n42611) );
  XOR U52315 ( .A(n42613), .B(n42611), .Z(n42895) );
  IV U52316 ( .A(n39429), .Z(n39431) );
  NOR U52317 ( .A(n39431), .B(n39430), .Z(n42893) );
  XOR U52318 ( .A(n42895), .B(n42893), .Z(n42903) );
  IV U52319 ( .A(n39432), .Z(n39433) );
  NOR U52320 ( .A(n39434), .B(n39433), .Z(n42896) );
  IV U52321 ( .A(n39435), .Z(n39437) );
  NOR U52322 ( .A(n39437), .B(n39436), .Z(n42902) );
  NOR U52323 ( .A(n42896), .B(n42902), .Z(n39438) );
  XOR U52324 ( .A(n42903), .B(n39438), .Z(n42899) );
  IV U52325 ( .A(n39439), .Z(n39441) );
  NOR U52326 ( .A(n39441), .B(n39440), .Z(n42900) );
  IV U52327 ( .A(n39442), .Z(n39443) );
  NOR U52328 ( .A(n39443), .B(n39447), .Z(n42909) );
  NOR U52329 ( .A(n42900), .B(n42909), .Z(n39444) );
  XOR U52330 ( .A(n42899), .B(n39444), .Z(n42908) );
  IV U52331 ( .A(n39445), .Z(n39446) );
  NOR U52332 ( .A(n39447), .B(n39446), .Z(n42906) );
  XOR U52333 ( .A(n42908), .B(n42906), .Z(n42914) );
  IV U52334 ( .A(n39448), .Z(n39449) );
  NOR U52335 ( .A(n39450), .B(n39449), .Z(n42913) );
  NOR U52336 ( .A(n39452), .B(n39451), .Z(n42609) );
  NOR U52337 ( .A(n42913), .B(n42609), .Z(n39453) );
  IV U52338 ( .A(n39453), .Z(n39454) );
  NOR U52339 ( .A(n42607), .B(n39454), .Z(n39455) );
  XOR U52340 ( .A(n42914), .B(n39455), .Z(n42601) );
  IV U52341 ( .A(n39456), .Z(n39458) );
  IV U52342 ( .A(n39457), .Z(n39461) );
  NOR U52343 ( .A(n39458), .B(n39461), .Z(n42602) );
  NOR U52344 ( .A(n42604), .B(n42602), .Z(n39459) );
  XOR U52345 ( .A(n42601), .B(n39459), .Z(n42599) );
  IV U52346 ( .A(n39460), .Z(n39462) );
  NOR U52347 ( .A(n39462), .B(n39461), .Z(n42597) );
  XOR U52348 ( .A(n42599), .B(n42597), .Z(n42924) );
  IV U52349 ( .A(n39463), .Z(n39464) );
  NOR U52350 ( .A(n39467), .B(n39464), .Z(n42922) );
  XOR U52351 ( .A(n42924), .B(n42922), .Z(n42595) );
  IV U52352 ( .A(n39465), .Z(n39466) );
  NOR U52353 ( .A(n39467), .B(n39466), .Z(n42593) );
  XOR U52354 ( .A(n42595), .B(n42593), .Z(n42919) );
  XOR U52355 ( .A(n42918), .B(n42919), .Z(n42936) );
  IV U52356 ( .A(n39468), .Z(n39469) );
  NOR U52357 ( .A(n39476), .B(n39469), .Z(n42935) );
  IV U52358 ( .A(n39470), .Z(n39472) );
  NOR U52359 ( .A(n39472), .B(n39471), .Z(n42591) );
  NOR U52360 ( .A(n42935), .B(n42591), .Z(n39473) );
  XOR U52361 ( .A(n42936), .B(n39473), .Z(n42938) );
  IV U52362 ( .A(n39474), .Z(n39475) );
  NOR U52363 ( .A(n39476), .B(n39475), .Z(n42939) );
  IV U52364 ( .A(n39477), .Z(n39479) );
  NOR U52365 ( .A(n39479), .B(n39478), .Z(n42941) );
  NOR U52366 ( .A(n42939), .B(n42941), .Z(n39480) );
  XOR U52367 ( .A(n42938), .B(n39480), .Z(n42587) );
  NOR U52368 ( .A(n39481), .B(n42588), .Z(n39485) );
  IV U52369 ( .A(n39482), .Z(n42580) );
  NOR U52370 ( .A(n39483), .B(n42580), .Z(n39484) );
  NOR U52371 ( .A(n39485), .B(n39484), .Z(n39486) );
  XOR U52372 ( .A(n42587), .B(n39486), .Z(n42583) );
  IV U52373 ( .A(n39487), .Z(n39488) );
  NOR U52374 ( .A(n39489), .B(n39488), .Z(n42584) );
  IV U52375 ( .A(n39490), .Z(n39491) );
  NOR U52376 ( .A(n39492), .B(n39491), .Z(n42957) );
  NOR U52377 ( .A(n42584), .B(n42957), .Z(n39493) );
  XOR U52378 ( .A(n42583), .B(n39493), .Z(n42953) );
  NOR U52379 ( .A(n39494), .B(n42954), .Z(n39498) );
  IV U52380 ( .A(n39495), .Z(n39497) );
  NOR U52381 ( .A(n39497), .B(n39496), .Z(n42577) );
  NOR U52382 ( .A(n39498), .B(n42577), .Z(n39499) );
  XOR U52383 ( .A(n42953), .B(n39499), .Z(n42566) );
  NOR U52384 ( .A(n39500), .B(n42570), .Z(n39504) );
  IV U52385 ( .A(n39501), .Z(n39502) );
  NOR U52386 ( .A(n39503), .B(n39502), .Z(n42567) );
  NOR U52387 ( .A(n39504), .B(n42567), .Z(n39505) );
  XOR U52388 ( .A(n42566), .B(n39505), .Z(n46237) );
  XOR U52389 ( .A(n42565), .B(n46237), .Z(n42560) );
  IV U52390 ( .A(n39506), .Z(n39507) );
  NOR U52391 ( .A(n39508), .B(n39507), .Z(n42559) );
  IV U52392 ( .A(n39509), .Z(n39511) );
  NOR U52393 ( .A(n39511), .B(n39510), .Z(n42563) );
  NOR U52394 ( .A(n42559), .B(n42563), .Z(n39512) );
  XOR U52395 ( .A(n42560), .B(n39512), .Z(n42555) );
  XOR U52396 ( .A(n42553), .B(n42555), .Z(n42558) );
  IV U52397 ( .A(n42558), .Z(n39520) );
  IV U52398 ( .A(n39513), .Z(n39514) );
  NOR U52399 ( .A(n39515), .B(n39514), .Z(n42551) );
  IV U52400 ( .A(n39516), .Z(n39518) );
  NOR U52401 ( .A(n39518), .B(n39517), .Z(n42556) );
  NOR U52402 ( .A(n42551), .B(n42556), .Z(n39519) );
  XOR U52403 ( .A(n39520), .B(n39519), .Z(n42969) );
  IV U52404 ( .A(n39521), .Z(n39523) );
  NOR U52405 ( .A(n39523), .B(n39522), .Z(n42967) );
  XOR U52406 ( .A(n42969), .B(n42967), .Z(n42975) );
  XOR U52407 ( .A(n39524), .B(n42975), .Z(n39525) );
  IV U52408 ( .A(n39525), .Z(n42547) );
  XOR U52409 ( .A(n42545), .B(n42547), .Z(n42549) );
  XOR U52410 ( .A(n42548), .B(n42549), .Z(n42979) );
  XOR U52411 ( .A(n42978), .B(n42979), .Z(n42982) );
  XOR U52412 ( .A(n42981), .B(n42982), .Z(n42542) );
  IV U52413 ( .A(n39526), .Z(n39527) );
  NOR U52414 ( .A(n39527), .B(n39529), .Z(n42540) );
  XOR U52415 ( .A(n42542), .B(n42540), .Z(n42987) );
  IV U52416 ( .A(n39528), .Z(n39530) );
  NOR U52417 ( .A(n39530), .B(n39529), .Z(n42543) );
  XOR U52418 ( .A(n42987), .B(n42543), .Z(n42993) );
  IV U52419 ( .A(n42993), .Z(n39538) );
  IV U52420 ( .A(n39531), .Z(n39532) );
  NOR U52421 ( .A(n39533), .B(n39532), .Z(n42986) );
  IV U52422 ( .A(n39534), .Z(n39536) );
  NOR U52423 ( .A(n39536), .B(n39535), .Z(n42992) );
  NOR U52424 ( .A(n42986), .B(n42992), .Z(n39537) );
  XOR U52425 ( .A(n39538), .B(n39537), .Z(n42991) );
  IV U52426 ( .A(n39539), .Z(n39540) );
  NOR U52427 ( .A(n39541), .B(n39540), .Z(n42989) );
  XOR U52428 ( .A(n42991), .B(n42989), .Z(n42539) );
  XOR U52429 ( .A(n42537), .B(n42539), .Z(n42533) );
  XOR U52430 ( .A(n39542), .B(n42533), .Z(n42526) );
  IV U52431 ( .A(n39543), .Z(n39545) );
  NOR U52432 ( .A(n39545), .B(n39544), .Z(n42530) );
  IV U52433 ( .A(n39546), .Z(n39548) );
  NOR U52434 ( .A(n39548), .B(n39547), .Z(n42527) );
  NOR U52435 ( .A(n42530), .B(n42527), .Z(n39549) );
  XOR U52436 ( .A(n42526), .B(n39549), .Z(n43001) );
  XOR U52437 ( .A(n39550), .B(n43001), .Z(n42520) );
  XOR U52438 ( .A(n39551), .B(n42520), .Z(n42518) );
  XOR U52439 ( .A(n42517), .B(n42518), .Z(n43009) );
  XOR U52440 ( .A(n39552), .B(n43009), .Z(n39553) );
  IV U52441 ( .A(n39553), .Z(n43018) );
  XOR U52442 ( .A(n43011), .B(n43018), .Z(n43015) );
  IV U52443 ( .A(n43015), .Z(n39561) );
  IV U52444 ( .A(n39554), .Z(n39555) );
  NOR U52445 ( .A(n39556), .B(n39555), .Z(n43016) );
  IV U52446 ( .A(n39557), .Z(n39559) );
  IV U52447 ( .A(n39558), .Z(n39563) );
  NOR U52448 ( .A(n39559), .B(n39563), .Z(n43013) );
  NOR U52449 ( .A(n43016), .B(n43013), .Z(n39560) );
  XOR U52450 ( .A(n39561), .B(n39560), .Z(n42511) );
  IV U52451 ( .A(n39562), .Z(n39564) );
  NOR U52452 ( .A(n39564), .B(n39563), .Z(n42509) );
  XOR U52453 ( .A(n42511), .B(n42509), .Z(n42513) );
  XOR U52454 ( .A(n39565), .B(n42513), .Z(n42502) );
  IV U52455 ( .A(n39566), .Z(n39568) );
  NOR U52456 ( .A(n39568), .B(n39567), .Z(n42504) );
  NOR U52457 ( .A(n42501), .B(n42504), .Z(n39569) );
  XOR U52458 ( .A(n42502), .B(n39569), .Z(n42497) );
  NOR U52459 ( .A(n39574), .B(n42497), .Z(n46342) );
  NOR U52460 ( .A(n39570), .B(n42498), .Z(n39571) );
  XOR U52461 ( .A(n39571), .B(n42497), .Z(n42495) );
  IV U52462 ( .A(n39572), .Z(n39573) );
  NOR U52463 ( .A(n39573), .B(n39582), .Z(n39575) );
  IV U52464 ( .A(n39575), .Z(n42494) );
  XOR U52465 ( .A(n42495), .B(n42494), .Z(n39577) );
  NOR U52466 ( .A(n39575), .B(n39574), .Z(n39576) );
  NOR U52467 ( .A(n39577), .B(n39576), .Z(n39578) );
  NOR U52468 ( .A(n46342), .B(n39578), .Z(n39579) );
  IV U52469 ( .A(n39579), .Z(n42490) );
  IV U52470 ( .A(n39580), .Z(n39581) );
  NOR U52471 ( .A(n39582), .B(n39581), .Z(n42488) );
  XOR U52472 ( .A(n42490), .B(n42488), .Z(n42492) );
  XOR U52473 ( .A(n39583), .B(n42492), .Z(n39593) );
  IV U52474 ( .A(n39593), .Z(n42485) );
  XOR U52475 ( .A(n39584), .B(n42485), .Z(n39596) );
  IV U52476 ( .A(n39596), .Z(n42481) );
  IV U52477 ( .A(n39585), .Z(n39587) );
  NOR U52478 ( .A(n39587), .B(n39586), .Z(n39600) );
  IV U52479 ( .A(n39600), .Z(n39588) );
  NOR U52480 ( .A(n42481), .B(n39588), .Z(n46375) );
  IV U52481 ( .A(n39589), .Z(n39591) );
  NOR U52482 ( .A(n39591), .B(n39590), .Z(n39597) );
  IV U52483 ( .A(n39597), .Z(n39595) );
  IV U52484 ( .A(n39592), .Z(n42484) );
  XOR U52485 ( .A(n39593), .B(n42484), .Z(n39594) );
  NOR U52486 ( .A(n39595), .B(n39594), .Z(n46371) );
  NOR U52487 ( .A(n39597), .B(n39596), .Z(n39598) );
  NOR U52488 ( .A(n46371), .B(n39598), .Z(n39599) );
  NOR U52489 ( .A(n39600), .B(n39599), .Z(n39601) );
  NOR U52490 ( .A(n46375), .B(n39601), .Z(n43028) );
  XOR U52491 ( .A(n39602), .B(n43028), .Z(n42472) );
  XOR U52492 ( .A(n39603), .B(n42472), .Z(n42468) );
  XOR U52493 ( .A(n39604), .B(n42468), .Z(n42460) );
  XOR U52494 ( .A(n42462), .B(n42460), .Z(n42464) );
  XOR U52495 ( .A(n42463), .B(n42464), .Z(n45776) );
  XOR U52496 ( .A(n43036), .B(n45776), .Z(n43038) );
  IV U52497 ( .A(n39605), .Z(n39606) );
  NOR U52498 ( .A(n39607), .B(n39606), .Z(n43037) );
  IV U52499 ( .A(n39608), .Z(n39609) );
  NOR U52500 ( .A(n42451), .B(n39609), .Z(n43042) );
  NOR U52501 ( .A(n43037), .B(n43042), .Z(n39610) );
  XOR U52502 ( .A(n43038), .B(n39610), .Z(n43052) );
  IV U52503 ( .A(n43052), .Z(n39616) );
  NOR U52504 ( .A(n39612), .B(n39611), .Z(n43045) );
  NOR U52505 ( .A(n39613), .B(n43051), .Z(n39614) );
  XOR U52506 ( .A(n43045), .B(n39614), .Z(n39615) );
  XOR U52507 ( .A(n39616), .B(n39615), .Z(n43050) );
  XOR U52508 ( .A(n43048), .B(n43050), .Z(n43057) );
  IV U52509 ( .A(n43057), .Z(n39623) );
  IV U52510 ( .A(n39617), .Z(n39618) );
  NOR U52511 ( .A(n39619), .B(n39618), .Z(n43056) );
  IV U52512 ( .A(n39620), .Z(n39621) );
  NOR U52513 ( .A(n39621), .B(n39627), .Z(n42448) );
  NOR U52514 ( .A(n43056), .B(n42448), .Z(n39622) );
  XOR U52515 ( .A(n39623), .B(n39622), .Z(n42444) );
  IV U52516 ( .A(n39624), .Z(n42445) );
  NOR U52517 ( .A(n42445), .B(n39625), .Z(n39629) );
  IV U52518 ( .A(n39626), .Z(n39628) );
  NOR U52519 ( .A(n39628), .B(n39627), .Z(n42441) );
  NOR U52520 ( .A(n39629), .B(n42441), .Z(n39630) );
  XOR U52521 ( .A(n42444), .B(n39630), .Z(n43060) );
  IV U52522 ( .A(n39631), .Z(n39633) );
  NOR U52523 ( .A(n39633), .B(n39632), .Z(n43059) );
  IV U52524 ( .A(n39634), .Z(n39635) );
  NOR U52525 ( .A(n39636), .B(n39635), .Z(n43066) );
  NOR U52526 ( .A(n43059), .B(n43066), .Z(n39637) );
  XOR U52527 ( .A(n43060), .B(n39637), .Z(n49250) );
  XOR U52528 ( .A(n49252), .B(n49250), .Z(n43072) );
  IV U52529 ( .A(n39638), .Z(n39639) );
  NOR U52530 ( .A(n39640), .B(n39639), .Z(n46439) );
  IV U52531 ( .A(n39641), .Z(n39642) );
  NOR U52532 ( .A(n39643), .B(n39642), .Z(n45755) );
  NOR U52533 ( .A(n46439), .B(n45755), .Z(n43073) );
  XOR U52534 ( .A(n43072), .B(n43073), .Z(n43079) );
  XOR U52535 ( .A(n43074), .B(n43079), .Z(n42439) );
  XOR U52536 ( .A(n39644), .B(n42439), .Z(n39645) );
  IV U52537 ( .A(n39645), .Z(n42437) );
  XOR U52538 ( .A(n42435), .B(n42437), .Z(n42430) );
  XOR U52539 ( .A(n42429), .B(n42430), .Z(n42433) );
  IV U52540 ( .A(n42433), .Z(n39650) );
  IV U52541 ( .A(n39646), .Z(n39647) );
  NOR U52542 ( .A(n39648), .B(n39647), .Z(n42432) );
  NOR U52543 ( .A(n42432), .B(n42424), .Z(n39649) );
  XOR U52544 ( .A(n39650), .B(n39649), .Z(n42427) );
  XOR U52545 ( .A(n42426), .B(n42427), .Z(n42422) );
  XOR U52546 ( .A(n39651), .B(n42422), .Z(n42413) );
  IV U52547 ( .A(n39652), .Z(n39654) );
  NOR U52548 ( .A(n39654), .B(n39653), .Z(n39655) );
  IV U52549 ( .A(n39655), .Z(n42414) );
  XOR U52550 ( .A(n42413), .B(n42414), .Z(n42417) );
  IV U52551 ( .A(n39656), .Z(n39657) );
  NOR U52552 ( .A(n39658), .B(n39657), .Z(n42416) );
  NOR U52553 ( .A(n39659), .B(n42410), .Z(n39660) );
  NOR U52554 ( .A(n42416), .B(n39660), .Z(n39661) );
  XOR U52555 ( .A(n42417), .B(n39661), .Z(n42406) );
  IV U52556 ( .A(n39662), .Z(n39663) );
  NOR U52557 ( .A(n39664), .B(n39663), .Z(n42407) );
  IV U52558 ( .A(n39665), .Z(n39667) );
  NOR U52559 ( .A(n39667), .B(n39666), .Z(n43088) );
  NOR U52560 ( .A(n42407), .B(n43088), .Z(n39668) );
  XOR U52561 ( .A(n42406), .B(n39668), .Z(n43092) );
  XOR U52562 ( .A(n43091), .B(n43092), .Z(n42405) );
  NOR U52563 ( .A(n39669), .B(n42405), .Z(n45726) );
  IV U52564 ( .A(n39670), .Z(n39671) );
  NOR U52565 ( .A(n39672), .B(n39671), .Z(n42403) );
  XOR U52566 ( .A(n42405), .B(n42403), .Z(n39678) );
  IV U52567 ( .A(n39678), .Z(n39673) );
  NOR U52568 ( .A(n39674), .B(n39673), .Z(n39675) );
  NOR U52569 ( .A(n45726), .B(n39675), .Z(n39676) );
  NOR U52570 ( .A(n39677), .B(n39676), .Z(n39680) );
  IV U52571 ( .A(n39677), .Z(n39679) );
  NOR U52572 ( .A(n39679), .B(n39678), .Z(n46476) );
  NOR U52573 ( .A(n39680), .B(n46476), .Z(n42395) );
  XOR U52574 ( .A(n39681), .B(n42395), .Z(n42398) );
  XOR U52575 ( .A(n42397), .B(n42398), .Z(n49202) );
  XOR U52576 ( .A(n42393), .B(n49202), .Z(n39682) );
  XOR U52577 ( .A(n39683), .B(n39682), .Z(n42392) );
  IV U52578 ( .A(n39684), .Z(n39686) );
  IV U52579 ( .A(n39685), .Z(n39689) );
  NOR U52580 ( .A(n39686), .B(n39689), .Z(n39687) );
  IV U52581 ( .A(n39687), .Z(n42391) );
  XOR U52582 ( .A(n42392), .B(n42391), .Z(n39694) );
  IV U52583 ( .A(n39694), .Z(n39692) );
  IV U52584 ( .A(n39688), .Z(n39690) );
  NOR U52585 ( .A(n39690), .B(n39689), .Z(n39693) );
  IV U52586 ( .A(n39693), .Z(n39691) );
  NOR U52587 ( .A(n39692), .B(n39691), .Z(n46491) );
  NOR U52588 ( .A(n39694), .B(n39693), .Z(n42389) );
  NOR U52589 ( .A(n46491), .B(n42389), .Z(n39695) );
  IV U52590 ( .A(n39695), .Z(n46504) );
  XOR U52591 ( .A(n42379), .B(n46504), .Z(n43121) );
  IV U52592 ( .A(n39696), .Z(n39698) );
  NOR U52593 ( .A(n39698), .B(n39697), .Z(n43115) );
  IV U52594 ( .A(n39699), .Z(n39702) );
  NOR U52595 ( .A(n39700), .B(n39710), .Z(n39701) );
  IV U52596 ( .A(n39701), .Z(n39706) );
  NOR U52597 ( .A(n39702), .B(n39706), .Z(n43120) );
  NOR U52598 ( .A(n43115), .B(n43120), .Z(n39703) );
  XOR U52599 ( .A(n43121), .B(n39703), .Z(n39704) );
  IV U52600 ( .A(n39704), .Z(n43119) );
  IV U52601 ( .A(n39705), .Z(n39707) );
  NOR U52602 ( .A(n39707), .B(n39706), .Z(n39708) );
  IV U52603 ( .A(n39708), .Z(n43118) );
  XOR U52604 ( .A(n43119), .B(n43118), .Z(n39715) );
  IV U52605 ( .A(n39715), .Z(n39713) );
  IV U52606 ( .A(n39709), .Z(n39711) );
  NOR U52607 ( .A(n39711), .B(n39710), .Z(n39714) );
  IV U52608 ( .A(n39714), .Z(n39712) );
  NOR U52609 ( .A(n39713), .B(n39712), .Z(n46508) );
  NOR U52610 ( .A(n39715), .B(n39714), .Z(n43130) );
  NOR U52611 ( .A(n46508), .B(n43130), .Z(n43125) );
  IV U52612 ( .A(n39716), .Z(n39717) );
  NOR U52613 ( .A(n39718), .B(n39717), .Z(n45710) );
  IV U52614 ( .A(n39719), .Z(n39721) );
  NOR U52615 ( .A(n39721), .B(n39720), .Z(n46515) );
  NOR U52616 ( .A(n45710), .B(n46515), .Z(n39722) );
  IV U52617 ( .A(n39722), .Z(n43128) );
  NOR U52618 ( .A(n43124), .B(n43128), .Z(n39723) );
  XOR U52619 ( .A(n43125), .B(n39723), .Z(n43141) );
  XOR U52620 ( .A(n43139), .B(n43141), .Z(n43153) );
  XOR U52621 ( .A(n39724), .B(n43153), .Z(n42375) );
  XOR U52622 ( .A(n39725), .B(n42375), .Z(n42359) );
  XOR U52623 ( .A(n42360), .B(n42359), .Z(n42356) );
  IV U52624 ( .A(n39726), .Z(n39727) );
  NOR U52625 ( .A(n39728), .B(n39727), .Z(n39735) );
  IV U52626 ( .A(n39735), .Z(n39729) );
  NOR U52627 ( .A(n42356), .B(n39729), .Z(n45696) );
  IV U52628 ( .A(n39730), .Z(n39731) );
  NOR U52629 ( .A(n39732), .B(n39731), .Z(n42354) );
  NOR U52630 ( .A(n42354), .B(n39733), .Z(n39734) );
  XOR U52631 ( .A(n39734), .B(n42356), .Z(n42351) );
  NOR U52632 ( .A(n39735), .B(n42351), .Z(n39736) );
  NOR U52633 ( .A(n45696), .B(n39736), .Z(n43159) );
  XOR U52634 ( .A(n39737), .B(n43159), .Z(n43164) );
  XOR U52635 ( .A(n43162), .B(n43164), .Z(n43167) );
  IV U52636 ( .A(n39738), .Z(n39740) );
  IV U52637 ( .A(n39739), .Z(n39742) );
  NOR U52638 ( .A(n39740), .B(n39742), .Z(n43165) );
  XOR U52639 ( .A(n43167), .B(n43165), .Z(n42346) );
  IV U52640 ( .A(n39741), .Z(n39743) );
  NOR U52641 ( .A(n39743), .B(n39742), .Z(n42344) );
  XOR U52642 ( .A(n42346), .B(n42344), .Z(n42348) );
  IV U52643 ( .A(n39744), .Z(n39745) );
  NOR U52644 ( .A(n39746), .B(n39745), .Z(n42347) );
  IV U52645 ( .A(n39747), .Z(n39748) );
  NOR U52646 ( .A(n39749), .B(n39748), .Z(n42342) );
  NOR U52647 ( .A(n42347), .B(n42342), .Z(n39750) );
  XOR U52648 ( .A(n42348), .B(n39750), .Z(n43170) );
  IV U52649 ( .A(n39751), .Z(n39753) );
  NOR U52650 ( .A(n39753), .B(n39752), .Z(n43169) );
  IV U52651 ( .A(n39754), .Z(n39755) );
  NOR U52652 ( .A(n39756), .B(n39755), .Z(n43173) );
  NOR U52653 ( .A(n43169), .B(n43173), .Z(n39757) );
  XOR U52654 ( .A(n43170), .B(n39757), .Z(n49936) );
  XOR U52655 ( .A(n39758), .B(n49936), .Z(n43178) );
  XOR U52656 ( .A(n43179), .B(n43178), .Z(n43182) );
  XOR U52657 ( .A(n39759), .B(n43182), .Z(n39760) );
  IV U52658 ( .A(n39760), .Z(n43189) );
  XOR U52659 ( .A(n43188), .B(n43189), .Z(n43191) );
  IV U52660 ( .A(n39761), .Z(n39762) );
  NOR U52661 ( .A(n39763), .B(n39762), .Z(n43190) );
  IV U52662 ( .A(n39764), .Z(n39766) );
  NOR U52663 ( .A(n39766), .B(n39765), .Z(n43195) );
  NOR U52664 ( .A(n43190), .B(n43195), .Z(n39767) );
  XOR U52665 ( .A(n43191), .B(n39767), .Z(n42340) );
  XOR U52666 ( .A(n42339), .B(n42340), .Z(n49112) );
  IV U52667 ( .A(n49112), .Z(n39768) );
  NOR U52668 ( .A(n39769), .B(n39768), .Z(n39774) );
  NOR U52669 ( .A(n39770), .B(n42340), .Z(n39771) );
  IV U52670 ( .A(n39771), .Z(n43204) );
  NOR U52671 ( .A(n43204), .B(n39772), .Z(n39773) );
  NOR U52672 ( .A(n39774), .B(n39773), .Z(n43206) );
  XOR U52673 ( .A(n43207), .B(n43206), .Z(n43209) );
  XOR U52674 ( .A(n39775), .B(n43209), .Z(n42333) );
  XOR U52675 ( .A(n39776), .B(n42333), .Z(n43217) );
  XOR U52676 ( .A(n39777), .B(n43217), .Z(n42324) );
  XOR U52677 ( .A(n39778), .B(n42324), .Z(n43235) );
  XOR U52678 ( .A(n39779), .B(n43235), .Z(n42321) );
  XOR U52679 ( .A(n39780), .B(n42321), .Z(n42319) );
  XOR U52680 ( .A(n42320), .B(n42319), .Z(n39783) );
  NOR U52681 ( .A(n39781), .B(n39783), .Z(n39790) );
  IV U52682 ( .A(n39782), .Z(n39785) );
  IV U52683 ( .A(n39783), .Z(n39784) );
  NOR U52684 ( .A(n39785), .B(n39784), .Z(n43239) );
  IV U52685 ( .A(n39786), .Z(n39787) );
  NOR U52686 ( .A(n39787), .B(n42319), .Z(n45652) );
  NOR U52687 ( .A(n43239), .B(n45652), .Z(n39788) );
  IV U52688 ( .A(n39788), .Z(n39789) );
  NOR U52689 ( .A(n39790), .B(n39789), .Z(n42315) );
  IV U52690 ( .A(n39791), .Z(n39793) );
  IV U52691 ( .A(n39792), .Z(n39796) );
  NOR U52692 ( .A(n39793), .B(n39796), .Z(n39794) );
  IV U52693 ( .A(n39794), .Z(n42316) );
  XOR U52694 ( .A(n42315), .B(n42316), .Z(n42314) );
  IV U52695 ( .A(n39795), .Z(n39802) );
  NOR U52696 ( .A(n39797), .B(n39796), .Z(n39798) );
  IV U52697 ( .A(n39798), .Z(n39799) );
  NOR U52698 ( .A(n39800), .B(n39799), .Z(n39801) );
  IV U52699 ( .A(n39801), .Z(n39804) );
  NOR U52700 ( .A(n39802), .B(n39804), .Z(n42312) );
  XOR U52701 ( .A(n42314), .B(n42312), .Z(n43250) );
  IV U52702 ( .A(n39803), .Z(n39805) );
  NOR U52703 ( .A(n39805), .B(n39804), .Z(n43248) );
  XOR U52704 ( .A(n43250), .B(n43248), .Z(n45642) );
  IV U52705 ( .A(n45642), .Z(n39812) );
  IV U52706 ( .A(n39806), .Z(n39807) );
  NOR U52707 ( .A(n39808), .B(n39807), .Z(n45645) );
  IV U52708 ( .A(n39809), .Z(n39811) );
  NOR U52709 ( .A(n39811), .B(n39810), .Z(n45640) );
  NOR U52710 ( .A(n45645), .B(n45640), .Z(n43246) );
  XOR U52711 ( .A(n39812), .B(n43246), .Z(n42310) );
  XOR U52712 ( .A(n42309), .B(n42310), .Z(n43261) );
  XOR U52713 ( .A(n39813), .B(n43261), .Z(n42293) );
  XOR U52714 ( .A(n39814), .B(n42293), .Z(n42289) );
  NOR U52715 ( .A(n39815), .B(n42289), .Z(n46669) );
  IV U52716 ( .A(n39816), .Z(n39817) );
  NOR U52717 ( .A(n39818), .B(n39817), .Z(n39828) );
  IV U52718 ( .A(n39828), .Z(n39819) );
  NOR U52719 ( .A(n39819), .B(n42289), .Z(n46666) );
  IV U52720 ( .A(n39820), .Z(n39822) );
  IV U52721 ( .A(n39821), .Z(n39825) );
  NOR U52722 ( .A(n39822), .B(n39825), .Z(n42287) );
  XOR U52723 ( .A(n42289), .B(n42287), .Z(n42291) );
  IV U52724 ( .A(n39823), .Z(n39824) );
  NOR U52725 ( .A(n39825), .B(n39824), .Z(n39826) );
  IV U52726 ( .A(n39826), .Z(n42290) );
  XOR U52727 ( .A(n42291), .B(n42290), .Z(n39827) );
  NOR U52728 ( .A(n39828), .B(n39827), .Z(n39829) );
  NOR U52729 ( .A(n46666), .B(n39829), .Z(n39830) );
  NOR U52730 ( .A(n39831), .B(n39830), .Z(n39835) );
  NOR U52731 ( .A(n46669), .B(n39835), .Z(n39832) );
  NOR U52732 ( .A(n39833), .B(n39832), .Z(n39836) );
  IV U52733 ( .A(n39833), .Z(n39834) );
  NOR U52734 ( .A(n39835), .B(n39834), .Z(n45626) );
  NOR U52735 ( .A(n39836), .B(n45626), .Z(n42282) );
  XOR U52736 ( .A(n39837), .B(n42282), .Z(n49067) );
  XOR U52737 ( .A(n42276), .B(n49067), .Z(n43280) );
  IV U52738 ( .A(n43280), .Z(n39846) );
  IV U52739 ( .A(n39838), .Z(n39840) );
  IV U52740 ( .A(n39839), .Z(n39841) );
  NOR U52741 ( .A(n39840), .B(n39841), .Z(n43278) );
  NOR U52742 ( .A(n39842), .B(n39841), .Z(n43276) );
  NOR U52743 ( .A(n42278), .B(n43276), .Z(n39843) );
  IV U52744 ( .A(n39843), .Z(n39844) );
  NOR U52745 ( .A(n43278), .B(n39844), .Z(n39845) );
  XOR U52746 ( .A(n39846), .B(n39845), .Z(n43288) );
  IV U52747 ( .A(n39847), .Z(n39849) );
  NOR U52748 ( .A(n39849), .B(n39848), .Z(n43286) );
  XOR U52749 ( .A(n43288), .B(n43286), .Z(n43297) );
  XOR U52750 ( .A(n39850), .B(n43297), .Z(n42273) );
  NOR U52751 ( .A(n39851), .B(n42273), .Z(n43313) );
  IV U52752 ( .A(n39852), .Z(n39853) );
  NOR U52753 ( .A(n39854), .B(n39853), .Z(n43296) );
  IV U52754 ( .A(n39855), .Z(n39857) );
  NOR U52755 ( .A(n39857), .B(n39856), .Z(n42272) );
  NOR U52756 ( .A(n43296), .B(n42272), .Z(n39858) );
  XOR U52757 ( .A(n39858), .B(n42273), .Z(n39862) );
  NOR U52758 ( .A(n39859), .B(n39862), .Z(n39860) );
  NOR U52759 ( .A(n43313), .B(n39860), .Z(n39861) );
  NOR U52760 ( .A(n39863), .B(n39861), .Z(n39866) );
  IV U52761 ( .A(n39862), .Z(n39865) );
  IV U52762 ( .A(n39863), .Z(n39864) );
  NOR U52763 ( .A(n39865), .B(n39864), .Z(n45611) );
  NOR U52764 ( .A(n39866), .B(n45611), .Z(n43319) );
  XOR U52765 ( .A(n43321), .B(n43319), .Z(n43327) );
  IV U52766 ( .A(n39867), .Z(n39869) );
  NOR U52767 ( .A(n39869), .B(n39868), .Z(n43318) );
  IV U52768 ( .A(n39870), .Z(n39872) );
  NOR U52769 ( .A(n39872), .B(n39871), .Z(n43328) );
  NOR U52770 ( .A(n43318), .B(n43328), .Z(n39873) );
  XOR U52771 ( .A(n43327), .B(n39873), .Z(n42268) );
  XOR U52772 ( .A(n42267), .B(n42268), .Z(n42264) );
  IV U52773 ( .A(n39874), .Z(n42271) );
  NOR U52774 ( .A(n42269), .B(n42271), .Z(n39878) );
  IV U52775 ( .A(n39875), .Z(n39877) );
  NOR U52776 ( .A(n39877), .B(n39876), .Z(n42263) );
  NOR U52777 ( .A(n39878), .B(n42263), .Z(n39879) );
  XOR U52778 ( .A(n42264), .B(n39879), .Z(n43335) );
  IV U52779 ( .A(n39880), .Z(n39881) );
  NOR U52780 ( .A(n39882), .B(n39881), .Z(n39883) );
  IV U52781 ( .A(n39883), .Z(n39890) );
  NOR U52782 ( .A(n43335), .B(n39890), .Z(n45597) );
  IV U52783 ( .A(n39884), .Z(n39885) );
  NOR U52784 ( .A(n39885), .B(n39898), .Z(n39886) );
  IV U52785 ( .A(n39886), .Z(n42262) );
  IV U52786 ( .A(n39887), .Z(n39888) );
  NOR U52787 ( .A(n39889), .B(n39888), .Z(n43333) );
  XOR U52788 ( .A(n43333), .B(n43335), .Z(n42261) );
  XOR U52789 ( .A(n42262), .B(n42261), .Z(n39893) );
  IV U52790 ( .A(n42261), .Z(n39891) );
  NOR U52791 ( .A(n39891), .B(n39890), .Z(n39892) );
  NOR U52792 ( .A(n39893), .B(n39892), .Z(n39894) );
  NOR U52793 ( .A(n45597), .B(n39894), .Z(n39895) );
  IV U52794 ( .A(n39895), .Z(n42259) );
  IV U52795 ( .A(n39896), .Z(n39897) );
  NOR U52796 ( .A(n39898), .B(n39897), .Z(n42258) );
  XOR U52797 ( .A(n42259), .B(n42258), .Z(n45594) );
  XOR U52798 ( .A(n43339), .B(n45594), .Z(n39899) );
  IV U52799 ( .A(n39899), .Z(n42256) );
  IV U52800 ( .A(n39900), .Z(n39904) );
  NOR U52801 ( .A(n46701), .B(n39901), .Z(n39902) );
  IV U52802 ( .A(n39902), .Z(n39903) );
  NOR U52803 ( .A(n39904), .B(n39903), .Z(n42254) );
  XOR U52804 ( .A(n42256), .B(n42254), .Z(n43355) );
  IV U52805 ( .A(n43355), .Z(n39912) );
  IV U52806 ( .A(n39905), .Z(n39908) );
  IV U52807 ( .A(n39906), .Z(n39907) );
  NOR U52808 ( .A(n39908), .B(n39907), .Z(n43343) );
  IV U52809 ( .A(n39909), .Z(n39910) );
  NOR U52810 ( .A(n39915), .B(n39910), .Z(n43353) );
  NOR U52811 ( .A(n43343), .B(n43353), .Z(n39911) );
  XOR U52812 ( .A(n39912), .B(n39911), .Z(n43366) );
  IV U52813 ( .A(n39913), .Z(n39914) );
  NOR U52814 ( .A(n39915), .B(n39914), .Z(n43351) );
  XOR U52815 ( .A(n43366), .B(n43351), .Z(n43359) );
  XOR U52816 ( .A(n39916), .B(n43359), .Z(n42250) );
  XOR U52817 ( .A(n39917), .B(n42250), .Z(n42249) );
  IV U52818 ( .A(n39918), .Z(n39919) );
  NOR U52819 ( .A(n39927), .B(n39919), .Z(n39920) );
  IV U52820 ( .A(n39920), .Z(n39928) );
  NOR U52821 ( .A(n42249), .B(n39928), .Z(n46724) );
  IV U52822 ( .A(n39921), .Z(n39922) );
  NOR U52823 ( .A(n39923), .B(n39922), .Z(n39924) );
  IV U52824 ( .A(n39924), .Z(n42246) );
  IV U52825 ( .A(n39925), .Z(n39926) );
  NOR U52826 ( .A(n39927), .B(n39926), .Z(n42247) );
  XOR U52827 ( .A(n42249), .B(n42247), .Z(n42245) );
  XOR U52828 ( .A(n42246), .B(n42245), .Z(n39931) );
  IV U52829 ( .A(n42245), .Z(n39929) );
  NOR U52830 ( .A(n39929), .B(n39928), .Z(n39930) );
  NOR U52831 ( .A(n39931), .B(n39930), .Z(n39932) );
  NOR U52832 ( .A(n46724), .B(n39932), .Z(n42243) );
  XOR U52833 ( .A(n42244), .B(n42243), .Z(n43389) );
  XOR U52834 ( .A(n39933), .B(n43389), .Z(n39934) );
  IV U52835 ( .A(n39934), .Z(n43387) );
  XOR U52836 ( .A(n43386), .B(n43387), .Z(n42236) );
  IV U52837 ( .A(n39935), .Z(n39937) );
  NOR U52838 ( .A(n39937), .B(n39936), .Z(n42240) );
  IV U52839 ( .A(n39938), .Z(n39940) );
  NOR U52840 ( .A(n39940), .B(n39939), .Z(n42235) );
  NOR U52841 ( .A(n42240), .B(n42235), .Z(n39941) );
  XOR U52842 ( .A(n42236), .B(n39941), .Z(n42232) );
  IV U52843 ( .A(n39942), .Z(n39943) );
  NOR U52844 ( .A(n39944), .B(n39943), .Z(n39945) );
  IV U52845 ( .A(n39945), .Z(n39952) );
  NOR U52846 ( .A(n42232), .B(n39952), .Z(n42225) );
  IV U52847 ( .A(n39946), .Z(n39948) );
  NOR U52848 ( .A(n39948), .B(n39947), .Z(n39949) );
  IV U52849 ( .A(n39949), .Z(n43397) );
  NOR U52850 ( .A(n39950), .B(n42231), .Z(n39951) );
  XOR U52851 ( .A(n42232), .B(n39951), .Z(n43396) );
  XOR U52852 ( .A(n43397), .B(n43396), .Z(n39955) );
  IV U52853 ( .A(n43396), .Z(n39953) );
  NOR U52854 ( .A(n39953), .B(n39952), .Z(n39954) );
  NOR U52855 ( .A(n39955), .B(n39954), .Z(n39956) );
  NOR U52856 ( .A(n42225), .B(n39956), .Z(n43399) );
  IV U52857 ( .A(n39957), .Z(n39958) );
  NOR U52858 ( .A(n39958), .B(n39960), .Z(n43398) );
  IV U52859 ( .A(n39959), .Z(n39961) );
  NOR U52860 ( .A(n39961), .B(n39960), .Z(n39962) );
  NOR U52861 ( .A(n43398), .B(n39962), .Z(n43404) );
  XOR U52862 ( .A(n43399), .B(n43404), .Z(n42220) );
  XOR U52863 ( .A(n42218), .B(n42220), .Z(n42223) );
  XOR U52864 ( .A(n42221), .B(n42223), .Z(n42213) );
  XOR U52865 ( .A(n42212), .B(n42213), .Z(n42217) );
  XOR U52866 ( .A(n39963), .B(n42217), .Z(n42200) );
  XOR U52867 ( .A(n39964), .B(n42200), .Z(n42196) );
  IV U52868 ( .A(n39965), .Z(n39966) );
  NOR U52869 ( .A(n39967), .B(n39966), .Z(n42199) );
  IV U52870 ( .A(n39968), .Z(n39970) );
  NOR U52871 ( .A(n39970), .B(n39969), .Z(n42195) );
  NOR U52872 ( .A(n42199), .B(n42195), .Z(n39971) );
  XOR U52873 ( .A(n42196), .B(n39971), .Z(n43416) );
  XOR U52874 ( .A(n43414), .B(n43416), .Z(n42193) );
  XOR U52875 ( .A(n42191), .B(n42193), .Z(n43411) );
  XOR U52876 ( .A(n43410), .B(n43411), .Z(n43424) );
  XOR U52877 ( .A(n43422), .B(n43424), .Z(n43426) );
  XOR U52878 ( .A(n43425), .B(n43426), .Z(n42187) );
  XOR U52879 ( .A(n42185), .B(n42187), .Z(n42189) );
  XOR U52880 ( .A(n39972), .B(n42189), .Z(n42179) );
  IV U52881 ( .A(n42180), .Z(n39974) );
  NOR U52882 ( .A(n39974), .B(n39973), .Z(n39979) );
  NOR U52883 ( .A(n39975), .B(n42180), .Z(n39977) );
  NOR U52884 ( .A(n39977), .B(n39976), .Z(n39978) );
  NOR U52885 ( .A(n39979), .B(n39978), .Z(n39980) );
  IV U52886 ( .A(n39980), .Z(n43433) );
  XOR U52887 ( .A(n42179), .B(n43433), .Z(n43440) );
  IV U52888 ( .A(n39981), .Z(n39982) );
  NOR U52889 ( .A(n43437), .B(n39982), .Z(n43438) );
  XOR U52890 ( .A(n43440), .B(n43438), .Z(n45536) );
  IV U52891 ( .A(n45536), .Z(n39988) );
  IV U52892 ( .A(n39983), .Z(n39984) );
  NOR U52893 ( .A(n39985), .B(n39984), .Z(n43441) );
  NOR U52894 ( .A(n39986), .B(n45539), .Z(n42176) );
  NOR U52895 ( .A(n43441), .B(n42176), .Z(n39987) );
  XOR U52896 ( .A(n39988), .B(n39987), .Z(n42172) );
  IV U52897 ( .A(n39989), .Z(n39991) );
  NOR U52898 ( .A(n39991), .B(n39990), .Z(n42170) );
  XOR U52899 ( .A(n42172), .B(n42170), .Z(n42175) );
  XOR U52900 ( .A(n42173), .B(n42175), .Z(n42168) );
  XOR U52901 ( .A(n42167), .B(n42168), .Z(n45532) );
  NOR U52902 ( .A(n45530), .B(n45532), .Z(n43447) );
  NOR U52903 ( .A(n39993), .B(n39992), .Z(n39996) );
  IV U52904 ( .A(n39996), .Z(n39994) );
  NOR U52905 ( .A(n39994), .B(n42168), .Z(n46846) );
  IV U52906 ( .A(n45532), .Z(n39995) );
  NOR U52907 ( .A(n39996), .B(n39995), .Z(n39997) );
  NOR U52908 ( .A(n46846), .B(n39997), .Z(n40002) );
  NOR U52909 ( .A(n39998), .B(n40002), .Z(n39999) );
  NOR U52910 ( .A(n43447), .B(n39999), .Z(n40000) );
  NOR U52911 ( .A(n40001), .B(n40000), .Z(n40004) );
  IV U52912 ( .A(n40001), .Z(n40003) );
  IV U52913 ( .A(n40002), .Z(n48966) );
  NOR U52914 ( .A(n40003), .B(n48966), .Z(n45525) );
  NOR U52915 ( .A(n40004), .B(n45525), .Z(n42165) );
  XOR U52916 ( .A(n40005), .B(n42165), .Z(n42163) );
  XOR U52917 ( .A(n42161), .B(n42163), .Z(n42157) );
  IV U52918 ( .A(n40006), .Z(n40008) );
  NOR U52919 ( .A(n40008), .B(n40007), .Z(n42155) );
  XOR U52920 ( .A(n42157), .B(n42155), .Z(n42159) );
  XOR U52921 ( .A(n42158), .B(n42159), .Z(n42153) );
  IV U52922 ( .A(n42153), .Z(n40016) );
  IV U52923 ( .A(n40009), .Z(n40010) );
  NOR U52924 ( .A(n40019), .B(n40010), .Z(n42148) );
  IV U52925 ( .A(n40011), .Z(n40014) );
  IV U52926 ( .A(n40012), .Z(n40013) );
  NOR U52927 ( .A(n40014), .B(n40013), .Z(n42151) );
  NOR U52928 ( .A(n42148), .B(n42151), .Z(n40015) );
  XOR U52929 ( .A(n40016), .B(n40015), .Z(n43457) );
  IV U52930 ( .A(n40017), .Z(n40018) );
  NOR U52931 ( .A(n40019), .B(n40018), .Z(n43455) );
  XOR U52932 ( .A(n43457), .B(n43455), .Z(n43466) );
  XOR U52933 ( .A(n40020), .B(n43466), .Z(n40033) );
  IV U52934 ( .A(n40033), .Z(n43469) );
  IV U52935 ( .A(n40021), .Z(n40022) );
  NOR U52936 ( .A(n43470), .B(n40022), .Z(n40032) );
  IV U52937 ( .A(n40023), .Z(n40024) );
  NOR U52938 ( .A(n40025), .B(n40024), .Z(n42141) );
  NOR U52939 ( .A(n40032), .B(n42141), .Z(n40026) );
  XOR U52940 ( .A(n43469), .B(n40026), .Z(n40039) );
  IV U52941 ( .A(n40039), .Z(n40027) );
  NOR U52942 ( .A(n40028), .B(n40027), .Z(n43480) );
  IV U52943 ( .A(n40029), .Z(n40030) );
  NOR U52944 ( .A(n40030), .B(n40035), .Z(n40031) );
  IV U52945 ( .A(n40031), .Z(n42140) );
  IV U52946 ( .A(n40032), .Z(n42143) );
  XOR U52947 ( .A(n42143), .B(n40033), .Z(n40038) );
  IV U52948 ( .A(n40034), .Z(n40036) );
  NOR U52949 ( .A(n40036), .B(n40035), .Z(n40040) );
  IV U52950 ( .A(n40040), .Z(n40037) );
  NOR U52951 ( .A(n40038), .B(n40037), .Z(n46869) );
  NOR U52952 ( .A(n40040), .B(n40039), .Z(n40041) );
  NOR U52953 ( .A(n46869), .B(n40041), .Z(n40042) );
  IV U52954 ( .A(n40042), .Z(n42139) );
  XOR U52955 ( .A(n42140), .B(n42139), .Z(n40043) );
  NOR U52956 ( .A(n40044), .B(n40043), .Z(n40045) );
  NOR U52957 ( .A(n43480), .B(n40045), .Z(n42133) );
  XOR U52958 ( .A(n40046), .B(n42133), .Z(n42130) );
  IV U52959 ( .A(n40047), .Z(n40049) );
  NOR U52960 ( .A(n40049), .B(n40048), .Z(n42129) );
  IV U52961 ( .A(n40050), .Z(n40052) );
  NOR U52962 ( .A(n40052), .B(n40051), .Z(n42127) );
  NOR U52963 ( .A(n42129), .B(n42127), .Z(n40053) );
  XOR U52964 ( .A(n42130), .B(n40053), .Z(n42121) );
  XOR U52965 ( .A(n40054), .B(n42121), .Z(n42116) );
  XOR U52966 ( .A(n40055), .B(n42116), .Z(n42107) );
  XOR U52967 ( .A(n42108), .B(n42107), .Z(n42111) );
  XOR U52968 ( .A(n40056), .B(n42111), .Z(n40057) );
  IV U52969 ( .A(n40057), .Z(n42101) );
  IV U52970 ( .A(n40058), .Z(n40059) );
  NOR U52971 ( .A(n40060), .B(n40059), .Z(n42099) );
  XOR U52972 ( .A(n42101), .B(n42099), .Z(n42103) );
  IV U52973 ( .A(n42103), .Z(n40068) );
  IV U52974 ( .A(n40061), .Z(n40062) );
  NOR U52975 ( .A(n40063), .B(n40062), .Z(n42102) );
  IV U52976 ( .A(n40064), .Z(n40065) );
  NOR U52977 ( .A(n40066), .B(n40065), .Z(n42096) );
  NOR U52978 ( .A(n42102), .B(n42096), .Z(n40067) );
  XOR U52979 ( .A(n40068), .B(n40067), .Z(n42092) );
  XOR U52980 ( .A(n42090), .B(n42092), .Z(n42094) );
  XOR U52981 ( .A(n42093), .B(n42094), .Z(n42085) );
  XOR U52982 ( .A(n42084), .B(n42085), .Z(n42088) );
  XOR U52983 ( .A(n42087), .B(n42088), .Z(n45471) );
  XOR U52984 ( .A(n42083), .B(n45471), .Z(n40069) );
  IV U52985 ( .A(n40069), .Z(n43495) );
  XOR U52986 ( .A(n43494), .B(n43495), .Z(n43492) );
  XOR U52987 ( .A(n42080), .B(n43492), .Z(n42078) );
  IV U52988 ( .A(n42078), .Z(n40077) );
  IV U52989 ( .A(n40070), .Z(n40071) );
  NOR U52990 ( .A(n40072), .B(n40071), .Z(n43491) );
  IV U52991 ( .A(n40073), .Z(n40075) );
  NOR U52992 ( .A(n40075), .B(n40074), .Z(n42077) );
  NOR U52993 ( .A(n43491), .B(n42077), .Z(n40076) );
  XOR U52994 ( .A(n40077), .B(n40076), .Z(n42074) );
  XOR U52995 ( .A(n42072), .B(n42074), .Z(n43517) );
  XOR U52996 ( .A(n40078), .B(n43517), .Z(n40079) );
  IV U52997 ( .A(n40079), .Z(n43514) );
  XOR U52998 ( .A(n43512), .B(n43514), .Z(n42067) );
  XOR U52999 ( .A(n42066), .B(n42067), .Z(n42070) );
  XOR U53000 ( .A(n42069), .B(n42070), .Z(n43524) );
  IV U53001 ( .A(n43524), .Z(n40086) );
  IV U53002 ( .A(n40080), .Z(n40081) );
  NOR U53003 ( .A(n40082), .B(n40081), .Z(n42064) );
  IV U53004 ( .A(n40083), .Z(n40084) );
  NOR U53005 ( .A(n40084), .B(n40088), .Z(n43522) );
  NOR U53006 ( .A(n42064), .B(n43522), .Z(n40085) );
  XOR U53007 ( .A(n40086), .B(n40085), .Z(n43528) );
  IV U53008 ( .A(n40087), .Z(n40089) );
  NOR U53009 ( .A(n40089), .B(n40088), .Z(n43520) );
  XOR U53010 ( .A(n43528), .B(n43520), .Z(n42062) );
  XOR U53011 ( .A(n40090), .B(n42062), .Z(n42054) );
  XOR U53012 ( .A(n40091), .B(n42054), .Z(n48887) );
  XOR U53013 ( .A(n43538), .B(n48887), .Z(n40092) );
  IV U53014 ( .A(n40092), .Z(n42051) );
  XOR U53015 ( .A(n42050), .B(n42051), .Z(n43536) );
  IV U53016 ( .A(n40093), .Z(n40095) );
  NOR U53017 ( .A(n40095), .B(n40094), .Z(n43534) );
  XOR U53018 ( .A(n43536), .B(n43534), .Z(n46943) );
  IV U53019 ( .A(n46943), .Z(n40102) );
  IV U53020 ( .A(n40096), .Z(n40097) );
  NOR U53021 ( .A(n40098), .B(n40097), .Z(n46941) );
  IV U53022 ( .A(n40099), .Z(n40100) );
  NOR U53023 ( .A(n40101), .B(n40100), .Z(n46948) );
  NOR U53024 ( .A(n46941), .B(n46948), .Z(n43553) );
  XOR U53025 ( .A(n40102), .B(n43553), .Z(n42048) );
  XOR U53026 ( .A(n42046), .B(n42048), .Z(n43551) );
  NOR U53027 ( .A(n40110), .B(n43551), .Z(n45437) );
  IV U53028 ( .A(n40103), .Z(n40109) );
  IV U53029 ( .A(n40104), .Z(n40105) );
  NOR U53030 ( .A(n40109), .B(n40105), .Z(n40106) );
  IV U53031 ( .A(n40106), .Z(n42045) );
  IV U53032 ( .A(n40107), .Z(n40108) );
  NOR U53033 ( .A(n40109), .B(n40108), .Z(n43549) );
  XOR U53034 ( .A(n43551), .B(n43549), .Z(n42044) );
  XOR U53035 ( .A(n42045), .B(n42044), .Z(n40113) );
  IV U53036 ( .A(n42044), .Z(n40111) );
  NOR U53037 ( .A(n40111), .B(n40110), .Z(n40112) );
  NOR U53038 ( .A(n40113), .B(n40112), .Z(n40114) );
  NOR U53039 ( .A(n45437), .B(n40114), .Z(n40115) );
  IV U53040 ( .A(n40115), .Z(n43562) );
  IV U53041 ( .A(n40116), .Z(n40118) );
  NOR U53042 ( .A(n40118), .B(n40117), .Z(n43561) );
  XOR U53043 ( .A(n43562), .B(n43561), .Z(n43567) );
  XOR U53044 ( .A(n43565), .B(n43567), .Z(n43569) );
  XOR U53045 ( .A(n43568), .B(n43569), .Z(n43576) );
  XOR U53046 ( .A(n40119), .B(n43576), .Z(n42035) );
  XOR U53047 ( .A(n40120), .B(n42035), .Z(n42032) );
  XOR U53048 ( .A(n40121), .B(n42032), .Z(n43584) );
  XOR U53049 ( .A(n40122), .B(n43584), .Z(n42022) );
  XOR U53050 ( .A(n42021), .B(n42022), .Z(n42018) );
  XOR U53051 ( .A(n42017), .B(n42018), .Z(n42015) );
  XOR U53052 ( .A(n42012), .B(n42015), .Z(n43599) );
  XOR U53053 ( .A(n40123), .B(n43599), .Z(n40124) );
  IV U53054 ( .A(n40124), .Z(n42009) );
  XOR U53055 ( .A(n42007), .B(n42009), .Z(n43604) );
  NOR U53056 ( .A(n40126), .B(n40125), .Z(n42010) );
  IV U53057 ( .A(n40127), .Z(n40129) );
  IV U53058 ( .A(n40128), .Z(n40132) );
  NOR U53059 ( .A(n40129), .B(n40132), .Z(n43603) );
  NOR U53060 ( .A(n42010), .B(n43603), .Z(n40130) );
  XOR U53061 ( .A(n43604), .B(n40130), .Z(n42004) );
  IV U53062 ( .A(n40131), .Z(n40133) );
  NOR U53063 ( .A(n40133), .B(n40132), .Z(n43601) );
  IV U53064 ( .A(n40134), .Z(n40136) );
  NOR U53065 ( .A(n40136), .B(n40135), .Z(n43607) );
  NOR U53066 ( .A(n43601), .B(n43607), .Z(n40137) );
  IV U53067 ( .A(n40137), .Z(n40138) );
  NOR U53068 ( .A(n42005), .B(n40138), .Z(n40139) );
  XOR U53069 ( .A(n42004), .B(n40139), .Z(n45417) );
  XOR U53070 ( .A(n42000), .B(n45417), .Z(n40144) );
  IV U53071 ( .A(n40144), .Z(n42002) );
  NOR U53072 ( .A(n40140), .B(n42002), .Z(n45408) );
  IV U53073 ( .A(n40141), .Z(n40142) );
  NOR U53074 ( .A(n40142), .B(n40147), .Z(n40143) );
  IV U53075 ( .A(n40143), .Z(n42001) );
  XOR U53076 ( .A(n40144), .B(n42001), .Z(n41999) );
  IV U53077 ( .A(n40145), .Z(n40146) );
  NOR U53078 ( .A(n40147), .B(n40146), .Z(n40148) );
  IV U53079 ( .A(n40148), .Z(n41998) );
  XOR U53080 ( .A(n41999), .B(n41998), .Z(n40149) );
  NOR U53081 ( .A(n40150), .B(n40149), .Z(n40151) );
  NOR U53082 ( .A(n45408), .B(n40151), .Z(n43613) );
  IV U53083 ( .A(n40153), .Z(n43618) );
  NOR U53084 ( .A(n40152), .B(n43618), .Z(n43612) );
  NOR U53085 ( .A(n40154), .B(n40153), .Z(n40156) );
  IV U53086 ( .A(n40155), .Z(n43621) );
  NOR U53087 ( .A(n40156), .B(n43621), .Z(n40157) );
  NOR U53088 ( .A(n43612), .B(n40157), .Z(n40158) );
  XOR U53089 ( .A(n43613), .B(n40158), .Z(n41997) );
  IV U53090 ( .A(n41997), .Z(n40165) );
  IV U53091 ( .A(n40159), .Z(n40160) );
  NOR U53092 ( .A(n40168), .B(n40160), .Z(n41993) );
  IV U53093 ( .A(n40161), .Z(n40163) );
  NOR U53094 ( .A(n40163), .B(n40162), .Z(n41995) );
  NOR U53095 ( .A(n41993), .B(n41995), .Z(n40164) );
  XOR U53096 ( .A(n40165), .B(n40164), .Z(n41989) );
  IV U53097 ( .A(n40166), .Z(n40167) );
  NOR U53098 ( .A(n40168), .B(n40167), .Z(n41987) );
  XOR U53099 ( .A(n41989), .B(n41987), .Z(n41991) );
  XOR U53100 ( .A(n41990), .B(n41991), .Z(n41985) );
  XOR U53101 ( .A(n41984), .B(n41985), .Z(n43625) );
  XOR U53102 ( .A(n43624), .B(n43625), .Z(n43632) );
  IV U53103 ( .A(n40169), .Z(n40171) );
  NOR U53104 ( .A(n40171), .B(n40170), .Z(n43633) );
  IV U53105 ( .A(n40172), .Z(n40173) );
  NOR U53106 ( .A(n40174), .B(n40173), .Z(n43629) );
  NOR U53107 ( .A(n43633), .B(n43629), .Z(n40175) );
  XOR U53108 ( .A(n43632), .B(n40175), .Z(n43640) );
  XOR U53109 ( .A(n40176), .B(n43640), .Z(n43639) );
  XOR U53110 ( .A(n40177), .B(n43639), .Z(n40186) );
  XOR U53111 ( .A(n40178), .B(n40186), .Z(n40183) );
  IV U53112 ( .A(n40183), .Z(n40181) );
  NOR U53113 ( .A(n40185), .B(n40182), .Z(n40179) );
  IV U53114 ( .A(n40179), .Z(n40180) );
  NOR U53115 ( .A(n40181), .B(n40180), .Z(n40189) );
  IV U53116 ( .A(n40182), .Z(n40184) );
  NOR U53117 ( .A(n40184), .B(n40183), .Z(n45383) );
  IV U53118 ( .A(n40185), .Z(n40187) );
  IV U53119 ( .A(n40186), .Z(n41979) );
  NOR U53120 ( .A(n40187), .B(n41979), .Z(n45389) );
  NOR U53121 ( .A(n45383), .B(n45389), .Z(n40188) );
  IV U53122 ( .A(n40188), .Z(n41977) );
  NOR U53123 ( .A(n40189), .B(n41977), .Z(n41973) );
  IV U53124 ( .A(n40190), .Z(n40192) );
  NOR U53125 ( .A(n40192), .B(n40191), .Z(n43647) );
  NOR U53126 ( .A(n41972), .B(n43647), .Z(n40193) );
  XOR U53127 ( .A(n41973), .B(n40193), .Z(n43652) );
  IV U53128 ( .A(n40194), .Z(n40196) );
  NOR U53129 ( .A(n40196), .B(n40195), .Z(n43650) );
  IV U53130 ( .A(n40197), .Z(n40199) );
  NOR U53131 ( .A(n40199), .B(n40198), .Z(n41970) );
  NOR U53132 ( .A(n43650), .B(n41970), .Z(n40200) );
  XOR U53133 ( .A(n43652), .B(n40200), .Z(n41965) );
  IV U53134 ( .A(n40201), .Z(n40203) );
  NOR U53135 ( .A(n40203), .B(n40202), .Z(n41967) );
  NOR U53136 ( .A(n40205), .B(n40204), .Z(n41964) );
  NOR U53137 ( .A(n41967), .B(n41964), .Z(n40206) );
  XOR U53138 ( .A(n41965), .B(n40206), .Z(n41963) );
  NOR U53139 ( .A(n41961), .B(n41956), .Z(n40207) );
  XOR U53140 ( .A(n41963), .B(n40207), .Z(n41959) );
  NOR U53141 ( .A(n40209), .B(n40208), .Z(n41958) );
  IV U53142 ( .A(n40210), .Z(n40212) );
  NOR U53143 ( .A(n40212), .B(n40211), .Z(n43657) );
  NOR U53144 ( .A(n41958), .B(n43657), .Z(n40213) );
  XOR U53145 ( .A(n41959), .B(n40213), .Z(n43656) );
  IV U53146 ( .A(n40214), .Z(n40216) );
  NOR U53147 ( .A(n40216), .B(n40215), .Z(n43654) );
  XOR U53148 ( .A(n43656), .B(n43654), .Z(n43664) );
  XOR U53149 ( .A(n43663), .B(n43664), .Z(n41955) );
  XOR U53150 ( .A(n40217), .B(n41955), .Z(n43678) );
  XOR U53151 ( .A(n43677), .B(n43678), .Z(n43681) );
  XOR U53152 ( .A(n43680), .B(n43681), .Z(n41940) );
  XOR U53153 ( .A(n40218), .B(n41940), .Z(n40219) );
  IV U53154 ( .A(n40219), .Z(n41934) );
  XOR U53155 ( .A(n41932), .B(n41934), .Z(n43688) );
  IV U53156 ( .A(n43688), .Z(n40227) );
  IV U53157 ( .A(n40220), .Z(n40221) );
  NOR U53158 ( .A(n40222), .B(n40221), .Z(n41935) );
  IV U53159 ( .A(n40223), .Z(n40225) );
  NOR U53160 ( .A(n40225), .B(n40224), .Z(n43687) );
  NOR U53161 ( .A(n41935), .B(n43687), .Z(n40226) );
  XOR U53162 ( .A(n40227), .B(n40226), .Z(n43692) );
  IV U53163 ( .A(n40228), .Z(n40230) );
  NOR U53164 ( .A(n40230), .B(n40229), .Z(n43690) );
  XOR U53165 ( .A(n43692), .B(n43690), .Z(n43695) );
  XOR U53166 ( .A(n43693), .B(n43695), .Z(n41927) );
  XOR U53167 ( .A(n40231), .B(n41927), .Z(n41919) );
  XOR U53168 ( .A(n40232), .B(n41919), .Z(n41917) );
  XOR U53169 ( .A(n40233), .B(n41917), .Z(n40234) );
  IV U53170 ( .A(n40234), .Z(n41910) );
  NOR U53171 ( .A(n40235), .B(n41910), .Z(n45330) );
  NOR U53172 ( .A(n40236), .B(n41911), .Z(n40237) );
  XOR U53173 ( .A(n40237), .B(n41910), .Z(n40240) );
  NOR U53174 ( .A(n40244), .B(n40240), .Z(n40238) );
  IV U53175 ( .A(n40238), .Z(n45324) );
  NOR U53176 ( .A(n40245), .B(n45324), .Z(n40239) );
  NOR U53177 ( .A(n45330), .B(n40239), .Z(n43706) );
  IV U53178 ( .A(n43706), .Z(n40243) );
  IV U53179 ( .A(n40240), .Z(n40248) );
  NOR U53180 ( .A(n40241), .B(n40248), .Z(n40242) );
  NOR U53181 ( .A(n40243), .B(n40242), .Z(n40250) );
  NOR U53182 ( .A(n40245), .B(n40244), .Z(n40246) );
  IV U53183 ( .A(n40246), .Z(n40247) );
  NOR U53184 ( .A(n40248), .B(n40247), .Z(n40249) );
  NOR U53185 ( .A(n40250), .B(n40249), .Z(n45320) );
  IV U53186 ( .A(n40251), .Z(n40254) );
  IV U53187 ( .A(n40252), .Z(n40253) );
  NOR U53188 ( .A(n40254), .B(n40253), .Z(n45318) );
  IV U53189 ( .A(n40255), .Z(n40257) );
  IV U53190 ( .A(n40256), .Z(n40262) );
  NOR U53191 ( .A(n40257), .B(n40262), .Z(n47104) );
  NOR U53192 ( .A(n45318), .B(n47104), .Z(n43707) );
  XOR U53193 ( .A(n45320), .B(n43707), .Z(n41907) );
  IV U53194 ( .A(n40258), .Z(n40259) );
  NOR U53195 ( .A(n40260), .B(n40259), .Z(n41906) );
  IV U53196 ( .A(n40261), .Z(n40263) );
  NOR U53197 ( .A(n40263), .B(n40262), .Z(n43708) );
  NOR U53198 ( .A(n41906), .B(n43708), .Z(n40264) );
  XOR U53199 ( .A(n41907), .B(n40264), .Z(n41904) );
  XOR U53200 ( .A(n41903), .B(n41904), .Z(n43716) );
  XOR U53201 ( .A(n43713), .B(n43716), .Z(n40265) );
  NOR U53202 ( .A(n40266), .B(n40265), .Z(n43722) );
  IV U53203 ( .A(n40267), .Z(n40269) );
  NOR U53204 ( .A(n40269), .B(n40268), .Z(n43715) );
  NOR U53205 ( .A(n43713), .B(n43715), .Z(n40270) );
  XOR U53206 ( .A(n40270), .B(n43716), .Z(n43724) );
  NOR U53207 ( .A(n40271), .B(n43724), .Z(n40272) );
  NOR U53208 ( .A(n43722), .B(n40272), .Z(n41895) );
  NOR U53209 ( .A(n40273), .B(n43726), .Z(n41897) );
  IV U53210 ( .A(n40274), .Z(n40276) );
  IV U53211 ( .A(n40275), .Z(n40280) );
  NOR U53212 ( .A(n40276), .B(n40280), .Z(n41894) );
  NOR U53213 ( .A(n41897), .B(n41894), .Z(n40277) );
  XOR U53214 ( .A(n41895), .B(n40277), .Z(n41893) );
  IV U53215 ( .A(n41893), .Z(n40285) );
  IV U53216 ( .A(n40278), .Z(n40279) );
  NOR U53217 ( .A(n40280), .B(n40279), .Z(n41891) );
  IV U53218 ( .A(n40281), .Z(n40282) );
  NOR U53219 ( .A(n40283), .B(n40282), .Z(n41889) );
  NOR U53220 ( .A(n41891), .B(n41889), .Z(n40284) );
  XOR U53221 ( .A(n40285), .B(n40284), .Z(n43735) );
  IV U53222 ( .A(n40286), .Z(n40287) );
  NOR U53223 ( .A(n40287), .B(n40289), .Z(n43733) );
  XOR U53224 ( .A(n43735), .B(n43733), .Z(n43738) );
  IV U53225 ( .A(n40288), .Z(n40290) );
  NOR U53226 ( .A(n40290), .B(n40289), .Z(n43736) );
  XOR U53227 ( .A(n43738), .B(n43736), .Z(n41885) );
  IV U53228 ( .A(n41885), .Z(n40298) );
  IV U53229 ( .A(n40291), .Z(n40292) );
  NOR U53230 ( .A(n40293), .B(n40292), .Z(n41887) );
  IV U53231 ( .A(n40294), .Z(n40296) );
  NOR U53232 ( .A(n40296), .B(n40295), .Z(n41884) );
  NOR U53233 ( .A(n41887), .B(n41884), .Z(n40297) );
  XOR U53234 ( .A(n40298), .B(n40297), .Z(n41883) );
  IV U53235 ( .A(n40299), .Z(n40300) );
  NOR U53236 ( .A(n40300), .B(n40306), .Z(n40309) );
  IV U53237 ( .A(n40309), .Z(n40301) );
  NOR U53238 ( .A(n41883), .B(n40301), .Z(n45287) );
  IV U53239 ( .A(n40302), .Z(n40304) );
  NOR U53240 ( .A(n40304), .B(n40303), .Z(n41881) );
  IV U53241 ( .A(n40305), .Z(n40307) );
  NOR U53242 ( .A(n40307), .B(n40306), .Z(n41879) );
  NOR U53243 ( .A(n41881), .B(n41879), .Z(n40308) );
  XOR U53244 ( .A(n41883), .B(n40308), .Z(n43744) );
  NOR U53245 ( .A(n40309), .B(n43744), .Z(n40310) );
  NOR U53246 ( .A(n45287), .B(n40310), .Z(n40311) );
  IV U53247 ( .A(n40311), .Z(n41872) );
  XOR U53248 ( .A(n40312), .B(n41872), .Z(n43753) );
  IV U53249 ( .A(n43753), .Z(n40319) );
  NOR U53250 ( .A(n40313), .B(n41873), .Z(n40317) );
  IV U53251 ( .A(n40314), .Z(n40316) );
  IV U53252 ( .A(n40315), .Z(n40321) );
  NOR U53253 ( .A(n40316), .B(n40321), .Z(n43752) );
  NOR U53254 ( .A(n40317), .B(n43752), .Z(n40318) );
  XOR U53255 ( .A(n40319), .B(n40318), .Z(n43757) );
  IV U53256 ( .A(n40320), .Z(n40322) );
  NOR U53257 ( .A(n40322), .B(n40321), .Z(n43755) );
  XOR U53258 ( .A(n43757), .B(n43755), .Z(n41867) );
  XOR U53259 ( .A(n40323), .B(n41867), .Z(n40324) );
  IV U53260 ( .A(n40324), .Z(n41858) );
  IV U53261 ( .A(n40325), .Z(n40327) );
  NOR U53262 ( .A(n40327), .B(n40326), .Z(n41856) );
  XOR U53263 ( .A(n41858), .B(n41856), .Z(n41859) );
  IV U53264 ( .A(n41859), .Z(n41848) );
  IV U53265 ( .A(n40328), .Z(n40329) );
  NOR U53266 ( .A(n40330), .B(n40329), .Z(n41847) );
  IV U53267 ( .A(n40331), .Z(n40332) );
  NOR U53268 ( .A(n40333), .B(n40332), .Z(n41854) );
  NOR U53269 ( .A(n41847), .B(n41854), .Z(n40334) );
  XOR U53270 ( .A(n41848), .B(n40334), .Z(n43767) );
  XOR U53271 ( .A(n43765), .B(n43767), .Z(n41842) );
  XOR U53272 ( .A(n41840), .B(n41842), .Z(n41844) );
  XOR U53273 ( .A(n40335), .B(n41844), .Z(n41829) );
  XOR U53274 ( .A(n40336), .B(n41829), .Z(n43773) );
  XOR U53275 ( .A(n40337), .B(n43773), .Z(n41824) );
  XOR U53276 ( .A(n40338), .B(n41824), .Z(n43790) );
  IV U53277 ( .A(n40339), .Z(n40341) );
  NOR U53278 ( .A(n40341), .B(n40340), .Z(n43783) );
  IV U53279 ( .A(n40342), .Z(n40344) );
  NOR U53280 ( .A(n40344), .B(n40343), .Z(n43789) );
  NOR U53281 ( .A(n43783), .B(n43789), .Z(n40345) );
  XOR U53282 ( .A(n43790), .B(n40345), .Z(n41819) );
  XOR U53283 ( .A(n40346), .B(n41819), .Z(n41816) );
  XOR U53284 ( .A(n41815), .B(n41816), .Z(n43802) );
  XOR U53285 ( .A(n43801), .B(n43802), .Z(n43809) );
  XOR U53286 ( .A(n40347), .B(n43809), .Z(n40348) );
  IV U53287 ( .A(n40348), .Z(n43812) );
  IV U53288 ( .A(n40349), .Z(n40350) );
  NOR U53289 ( .A(n40351), .B(n40350), .Z(n43810) );
  XOR U53290 ( .A(n43812), .B(n43810), .Z(n43817) );
  IV U53291 ( .A(n43817), .Z(n40359) );
  IV U53292 ( .A(n40352), .Z(n40353) );
  NOR U53293 ( .A(n40354), .B(n40353), .Z(n43814) );
  IV U53294 ( .A(n40355), .Z(n40356) );
  NOR U53295 ( .A(n40357), .B(n40356), .Z(n43816) );
  NOR U53296 ( .A(n43814), .B(n43816), .Z(n40358) );
  XOR U53297 ( .A(n40359), .B(n40358), .Z(n43821) );
  IV U53298 ( .A(n40360), .Z(n40362) );
  NOR U53299 ( .A(n40362), .B(n40361), .Z(n43819) );
  IV U53300 ( .A(n40363), .Z(n40365) );
  NOR U53301 ( .A(n40365), .B(n40364), .Z(n41813) );
  NOR U53302 ( .A(n43819), .B(n41813), .Z(n40366) );
  XOR U53303 ( .A(n43821), .B(n40366), .Z(n40377) );
  IV U53304 ( .A(n40367), .Z(n40369) );
  NOR U53305 ( .A(n40369), .B(n40368), .Z(n47232) );
  IV U53306 ( .A(n40370), .Z(n40371) );
  NOR U53307 ( .A(n40371), .B(n40375), .Z(n47244) );
  NOR U53308 ( .A(n47232), .B(n47244), .Z(n40378) );
  IV U53309 ( .A(n40378), .Z(n40372) );
  NOR U53310 ( .A(n40377), .B(n40372), .Z(n40382) );
  IV U53311 ( .A(n40373), .Z(n40374) );
  NOR U53312 ( .A(n40375), .B(n40374), .Z(n40376) );
  IV U53313 ( .A(n40376), .Z(n40381) );
  NOR U53314 ( .A(n40382), .B(n40381), .Z(n47240) );
  IV U53315 ( .A(n40377), .Z(n47234) );
  NOR U53316 ( .A(n40378), .B(n47234), .Z(n40379) );
  NOR U53317 ( .A(n47240), .B(n40379), .Z(n40380) );
  IV U53318 ( .A(n40380), .Z(n41812) );
  NOR U53319 ( .A(n41812), .B(n40381), .Z(n40384) );
  NOR U53320 ( .A(n40382), .B(n41812), .Z(n40383) );
  NOR U53321 ( .A(n40384), .B(n40383), .Z(n41810) );
  XOR U53322 ( .A(n40385), .B(n41810), .Z(n41801) );
  XOR U53323 ( .A(n40386), .B(n41801), .Z(n41799) );
  NOR U53324 ( .A(n40394), .B(n41799), .Z(n50775) );
  IV U53325 ( .A(n40387), .Z(n40388) );
  NOR U53326 ( .A(n40389), .B(n40388), .Z(n40390) );
  IV U53327 ( .A(n40390), .Z(n43826) );
  IV U53328 ( .A(n40391), .Z(n40393) );
  NOR U53329 ( .A(n40393), .B(n40392), .Z(n41798) );
  XOR U53330 ( .A(n41798), .B(n41799), .Z(n43825) );
  XOR U53331 ( .A(n43826), .B(n43825), .Z(n40397) );
  IV U53332 ( .A(n43825), .Z(n40395) );
  NOR U53333 ( .A(n40395), .B(n40394), .Z(n40396) );
  NOR U53334 ( .A(n40397), .B(n40396), .Z(n40398) );
  NOR U53335 ( .A(n50775), .B(n40398), .Z(n41796) );
  XOR U53336 ( .A(n40399), .B(n41796), .Z(n41793) );
  XOR U53337 ( .A(n41792), .B(n41793), .Z(n43836) );
  IV U53338 ( .A(n43836), .Z(n40407) );
  IV U53339 ( .A(n40400), .Z(n40402) );
  NOR U53340 ( .A(n40402), .B(n40401), .Z(n43835) );
  IV U53341 ( .A(n40403), .Z(n40405) );
  IV U53342 ( .A(n40404), .Z(n40409) );
  NOR U53343 ( .A(n40405), .B(n40409), .Z(n43832) );
  NOR U53344 ( .A(n43835), .B(n43832), .Z(n40406) );
  XOR U53345 ( .A(n40407), .B(n40406), .Z(n43843) );
  IV U53346 ( .A(n40408), .Z(n40410) );
  NOR U53347 ( .A(n40410), .B(n40409), .Z(n41790) );
  XOR U53348 ( .A(n43843), .B(n41790), .Z(n41788) );
  XOR U53349 ( .A(n40411), .B(n41788), .Z(n41784) );
  IV U53350 ( .A(n40412), .Z(n40414) );
  NOR U53351 ( .A(n40414), .B(n40413), .Z(n41785) );
  IV U53352 ( .A(n40415), .Z(n40417) );
  NOR U53353 ( .A(n40417), .B(n40416), .Z(n43848) );
  NOR U53354 ( .A(n41785), .B(n43848), .Z(n40418) );
  XOR U53355 ( .A(n41784), .B(n40418), .Z(n43846) );
  XOR U53356 ( .A(n43845), .B(n43846), .Z(n41779) );
  XOR U53357 ( .A(n41778), .B(n41779), .Z(n41782) );
  XOR U53358 ( .A(n41781), .B(n41782), .Z(n43853) );
  XOR U53359 ( .A(n43852), .B(n43853), .Z(n40420) );
  NOR U53360 ( .A(n40425), .B(n40420), .Z(n48657) );
  NOR U53361 ( .A(n40419), .B(n41775), .Z(n40421) );
  XOR U53362 ( .A(n40421), .B(n40420), .Z(n41773) );
  IV U53363 ( .A(n40422), .Z(n40424) );
  NOR U53364 ( .A(n40424), .B(n40423), .Z(n40426) );
  IV U53365 ( .A(n40426), .Z(n41772) );
  XOR U53366 ( .A(n41773), .B(n41772), .Z(n40428) );
  NOR U53367 ( .A(n40426), .B(n40425), .Z(n40427) );
  NOR U53368 ( .A(n40428), .B(n40427), .Z(n40429) );
  NOR U53369 ( .A(n48657), .B(n40429), .Z(n40430) );
  IV U53370 ( .A(n40430), .Z(n43859) );
  XOR U53371 ( .A(n43858), .B(n43859), .Z(n43863) );
  IV U53372 ( .A(n40431), .Z(n40435) );
  XOR U53373 ( .A(n40433), .B(n40432), .Z(n40434) );
  NOR U53374 ( .A(n40435), .B(n40434), .Z(n43861) );
  XOR U53375 ( .A(n43863), .B(n43861), .Z(n41768) );
  IV U53376 ( .A(n40436), .Z(n40438) );
  NOR U53377 ( .A(n40438), .B(n40437), .Z(n41766) );
  XOR U53378 ( .A(n41768), .B(n41766), .Z(n41770) );
  IV U53379 ( .A(n40439), .Z(n40440) );
  NOR U53380 ( .A(n40441), .B(n40440), .Z(n41769) );
  NOR U53381 ( .A(n40443), .B(n40442), .Z(n41764) );
  NOR U53382 ( .A(n41769), .B(n41764), .Z(n40444) );
  XOR U53383 ( .A(n41770), .B(n40444), .Z(n43867) );
  XOR U53384 ( .A(n45201), .B(n43867), .Z(n43869) );
  XOR U53385 ( .A(n43868), .B(n43869), .Z(n41758) );
  IV U53386 ( .A(n40445), .Z(n41761) );
  NOR U53387 ( .A(n41761), .B(n40446), .Z(n40450) );
  IV U53388 ( .A(n40447), .Z(n40449) );
  NOR U53389 ( .A(n40449), .B(n40448), .Z(n41757) );
  NOR U53390 ( .A(n40450), .B(n41757), .Z(n40451) );
  XOR U53391 ( .A(n41758), .B(n40451), .Z(n41751) );
  IV U53392 ( .A(n40452), .Z(n40453) );
  NOR U53393 ( .A(n40454), .B(n40453), .Z(n41754) );
  IV U53394 ( .A(n40455), .Z(n40457) );
  NOR U53395 ( .A(n40457), .B(n40456), .Z(n41752) );
  NOR U53396 ( .A(n41754), .B(n41752), .Z(n40458) );
  XOR U53397 ( .A(n41751), .B(n40458), .Z(n41749) );
  IV U53398 ( .A(n40459), .Z(n40461) );
  NOR U53399 ( .A(n40461), .B(n40460), .Z(n41748) );
  IV U53400 ( .A(n40462), .Z(n40464) );
  NOR U53401 ( .A(n40464), .B(n40463), .Z(n41744) );
  NOR U53402 ( .A(n41748), .B(n41744), .Z(n40465) );
  XOR U53403 ( .A(n41749), .B(n40465), .Z(n41742) );
  XOR U53404 ( .A(n41747), .B(n41742), .Z(n43879) );
  IV U53405 ( .A(n40466), .Z(n40468) );
  NOR U53406 ( .A(n40468), .B(n40467), .Z(n41741) );
  IV U53407 ( .A(n40469), .Z(n40470) );
  NOR U53408 ( .A(n40471), .B(n40470), .Z(n43878) );
  NOR U53409 ( .A(n41741), .B(n43878), .Z(n40472) );
  XOR U53410 ( .A(n43879), .B(n40472), .Z(n41735) );
  XOR U53411 ( .A(n40473), .B(n41735), .Z(n43884) );
  XOR U53412 ( .A(n40474), .B(n43884), .Z(n43889) );
  XOR U53413 ( .A(n40475), .B(n43889), .Z(n43897) );
  XOR U53414 ( .A(n40476), .B(n43897), .Z(n40477) );
  IV U53415 ( .A(n40477), .Z(n41729) );
  XOR U53416 ( .A(n41727), .B(n41729), .Z(n47377) );
  IV U53417 ( .A(n40478), .Z(n40479) );
  NOR U53418 ( .A(n40480), .B(n40479), .Z(n41730) );
  IV U53419 ( .A(n40481), .Z(n40483) );
  NOR U53420 ( .A(n40483), .B(n40482), .Z(n41725) );
  NOR U53421 ( .A(n41730), .B(n41725), .Z(n47378) );
  XOR U53422 ( .A(n47377), .B(n47378), .Z(n43905) );
  XOR U53423 ( .A(n40484), .B(n43905), .Z(n43914) );
  IV U53424 ( .A(n40485), .Z(n40486) );
  NOR U53425 ( .A(n40487), .B(n40486), .Z(n40493) );
  IV U53426 ( .A(n40493), .Z(n40488) );
  NOR U53427 ( .A(n43914), .B(n40488), .Z(n45181) );
  IV U53428 ( .A(n40489), .Z(n40491) );
  NOR U53429 ( .A(n40491), .B(n40490), .Z(n43912) );
  XOR U53430 ( .A(n43912), .B(n43914), .Z(n40497) );
  IV U53431 ( .A(n40497), .Z(n40492) );
  NOR U53432 ( .A(n40493), .B(n40492), .Z(n40494) );
  NOR U53433 ( .A(n45181), .B(n40494), .Z(n40495) );
  NOR U53434 ( .A(n40496), .B(n40495), .Z(n40499) );
  IV U53435 ( .A(n40496), .Z(n40498) );
  NOR U53436 ( .A(n40498), .B(n40497), .Z(n47387) );
  NOR U53437 ( .A(n40499), .B(n47387), .Z(n40500) );
  IV U53438 ( .A(n40500), .Z(n41723) );
  XOR U53439 ( .A(n41722), .B(n41723), .Z(n43918) );
  IV U53440 ( .A(n43918), .Z(n40504) );
  NOR U53441 ( .A(n40502), .B(n40501), .Z(n43917) );
  NOR U53442 ( .A(n41720), .B(n43917), .Z(n40503) );
  XOR U53443 ( .A(n40504), .B(n40503), .Z(n43921) );
  XOR U53444 ( .A(n43920), .B(n43921), .Z(n43928) );
  XOR U53445 ( .A(n43926), .B(n43928), .Z(n41718) );
  XOR U53446 ( .A(n40505), .B(n41718), .Z(n41692) );
  NOR U53447 ( .A(n40507), .B(n40506), .Z(n40511) );
  IV U53448 ( .A(n40508), .Z(n40510) );
  NOR U53449 ( .A(n40510), .B(n40509), .Z(n41693) );
  NOR U53450 ( .A(n40511), .B(n41693), .Z(n40512) );
  XOR U53451 ( .A(n41692), .B(n40512), .Z(n43940) );
  XOR U53452 ( .A(n43939), .B(n43940), .Z(n43943) );
  NOR U53453 ( .A(n40522), .B(n43943), .Z(n45169) );
  IV U53454 ( .A(n40513), .Z(n40517) );
  NOR U53455 ( .A(n40515), .B(n40514), .Z(n40516) );
  IV U53456 ( .A(n40516), .Z(n40528) );
  NOR U53457 ( .A(n40517), .B(n40528), .Z(n40518) );
  IV U53458 ( .A(n40518), .Z(n41691) );
  IV U53459 ( .A(n40519), .Z(n40520) );
  NOR U53460 ( .A(n40521), .B(n40520), .Z(n43942) );
  XOR U53461 ( .A(n43942), .B(n43943), .Z(n41690) );
  XOR U53462 ( .A(n41691), .B(n41690), .Z(n40525) );
  IV U53463 ( .A(n41690), .Z(n40523) );
  NOR U53464 ( .A(n40523), .B(n40522), .Z(n40524) );
  NOR U53465 ( .A(n40525), .B(n40524), .Z(n40526) );
  NOR U53466 ( .A(n45169), .B(n40526), .Z(n43947) );
  IV U53467 ( .A(n40527), .Z(n40529) );
  NOR U53468 ( .A(n40529), .B(n40528), .Z(n40530) );
  IV U53469 ( .A(n40530), .Z(n43948) );
  XOR U53470 ( .A(n43947), .B(n43948), .Z(n43951) );
  XOR U53471 ( .A(n43950), .B(n43951), .Z(n41689) );
  IV U53472 ( .A(n40531), .Z(n40532) );
  NOR U53473 ( .A(n40533), .B(n40532), .Z(n41687) );
  IV U53474 ( .A(n40534), .Z(n40537) );
  NOR U53475 ( .A(n40535), .B(n40540), .Z(n40536) );
  IV U53476 ( .A(n40536), .Z(n40543) );
  NOR U53477 ( .A(n40537), .B(n40543), .Z(n41685) );
  NOR U53478 ( .A(n41687), .B(n41685), .Z(n40538) );
  XOR U53479 ( .A(n41689), .B(n40538), .Z(n41679) );
  IV U53480 ( .A(n40539), .Z(n40541) );
  NOR U53481 ( .A(n40541), .B(n40540), .Z(n41680) );
  IV U53482 ( .A(n40542), .Z(n40544) );
  NOR U53483 ( .A(n40544), .B(n40543), .Z(n41682) );
  NOR U53484 ( .A(n41680), .B(n41682), .Z(n40545) );
  XOR U53485 ( .A(n41679), .B(n40545), .Z(n41675) );
  IV U53486 ( .A(n40546), .Z(n40548) );
  NOR U53487 ( .A(n40548), .B(n40547), .Z(n41673) );
  XOR U53488 ( .A(n41675), .B(n41673), .Z(n41677) );
  IV U53489 ( .A(n41677), .Z(n40556) );
  IV U53490 ( .A(n40549), .Z(n40550) );
  NOR U53491 ( .A(n40551), .B(n40550), .Z(n41676) );
  IV U53492 ( .A(n40552), .Z(n40553) );
  NOR U53493 ( .A(n40554), .B(n40553), .Z(n41671) );
  NOR U53494 ( .A(n41676), .B(n41671), .Z(n40555) );
  XOR U53495 ( .A(n40556), .B(n40555), .Z(n41670) );
  XOR U53496 ( .A(n41668), .B(n41670), .Z(n41665) );
  XOR U53497 ( .A(n41663), .B(n41665), .Z(n41666) );
  IV U53498 ( .A(n40557), .Z(n40558) );
  NOR U53499 ( .A(n40571), .B(n40558), .Z(n40559) );
  IV U53500 ( .A(n40559), .Z(n41662) );
  IV U53501 ( .A(n40560), .Z(n40562) );
  NOR U53502 ( .A(n40562), .B(n40561), .Z(n40563) );
  IV U53503 ( .A(n40563), .Z(n41667) );
  XOR U53504 ( .A(n41662), .B(n41667), .Z(n40564) );
  XOR U53505 ( .A(n41666), .B(n40564), .Z(n41660) );
  IV U53506 ( .A(n40565), .Z(n40567) );
  NOR U53507 ( .A(n40567), .B(n40566), .Z(n40568) );
  IV U53508 ( .A(n40568), .Z(n40573) );
  NOR U53509 ( .A(n41660), .B(n40573), .Z(n47482) );
  IV U53510 ( .A(n40569), .Z(n40570) );
  NOR U53511 ( .A(n40571), .B(n40570), .Z(n40572) );
  IV U53512 ( .A(n40572), .Z(n41661) );
  XOR U53513 ( .A(n41661), .B(n41660), .Z(n40576) );
  IV U53514 ( .A(n41660), .Z(n40574) );
  NOR U53515 ( .A(n40574), .B(n40573), .Z(n40575) );
  NOR U53516 ( .A(n40576), .B(n40575), .Z(n41659) );
  NOR U53517 ( .A(n47482), .B(n41659), .Z(n43959) );
  XOR U53518 ( .A(n40577), .B(n43959), .Z(n43964) );
  XOR U53519 ( .A(n40578), .B(n43964), .Z(n40587) );
  IV U53520 ( .A(n40587), .Z(n43971) );
  NOR U53521 ( .A(n40588), .B(n43971), .Z(n47495) );
  IV U53522 ( .A(n40579), .Z(n40581) );
  NOR U53523 ( .A(n40581), .B(n40580), .Z(n40582) );
  IV U53524 ( .A(n40582), .Z(n41654) );
  IV U53525 ( .A(n40583), .Z(n40584) );
  NOR U53526 ( .A(n40585), .B(n40584), .Z(n40586) );
  IV U53527 ( .A(n40586), .Z(n43970) );
  XOR U53528 ( .A(n40587), .B(n43970), .Z(n41653) );
  XOR U53529 ( .A(n41654), .B(n41653), .Z(n40591) );
  IV U53530 ( .A(n41653), .Z(n40589) );
  NOR U53531 ( .A(n40589), .B(n40588), .Z(n40590) );
  NOR U53532 ( .A(n40591), .B(n40590), .Z(n40592) );
  NOR U53533 ( .A(n47495), .B(n40592), .Z(n41648) );
  XOR U53534 ( .A(n40593), .B(n41648), .Z(n41644) );
  XOR U53535 ( .A(n41642), .B(n41644), .Z(n43976) );
  IV U53536 ( .A(n40594), .Z(n40596) );
  NOR U53537 ( .A(n40596), .B(n40595), .Z(n41645) );
  IV U53538 ( .A(n40597), .Z(n40598) );
  NOR U53539 ( .A(n40599), .B(n40598), .Z(n43975) );
  NOR U53540 ( .A(n41645), .B(n43975), .Z(n40600) );
  XOR U53541 ( .A(n43976), .B(n40600), .Z(n43978) );
  IV U53542 ( .A(n40601), .Z(n40603) );
  NOR U53543 ( .A(n40603), .B(n40602), .Z(n43979) );
  NOR U53544 ( .A(n40605), .B(n40604), .Z(n43985) );
  NOR U53545 ( .A(n43979), .B(n43985), .Z(n40606) );
  XOR U53546 ( .A(n43978), .B(n40606), .Z(n43983) );
  IV U53547 ( .A(n40607), .Z(n41641) );
  NOR U53548 ( .A(n41641), .B(n40608), .Z(n40609) );
  NOR U53549 ( .A(n43982), .B(n40609), .Z(n41638) );
  XOR U53550 ( .A(n43983), .B(n41638), .Z(n43990) );
  XOR U53551 ( .A(n43991), .B(n43990), .Z(n43994) );
  XOR U53552 ( .A(n40610), .B(n43994), .Z(n41623) );
  XOR U53553 ( .A(n41622), .B(n41623), .Z(n41618) );
  XOR U53554 ( .A(n40611), .B(n41618), .Z(n41606) );
  NOR U53555 ( .A(n40612), .B(n41610), .Z(n40616) );
  IV U53556 ( .A(n40613), .Z(n40615) );
  NOR U53557 ( .A(n40615), .B(n40614), .Z(n41607) );
  NOR U53558 ( .A(n40616), .B(n41607), .Z(n40617) );
  XOR U53559 ( .A(n41606), .B(n40617), .Z(n41605) );
  XOR U53560 ( .A(n41603), .B(n41605), .Z(n43999) );
  XOR U53561 ( .A(n43998), .B(n43999), .Z(n44002) );
  XOR U53562 ( .A(n44001), .B(n44002), .Z(n47546) );
  XOR U53563 ( .A(n50901), .B(n47546), .Z(n44004) );
  NOR U53564 ( .A(n40619), .B(n40618), .Z(n44012) );
  IV U53565 ( .A(n40620), .Z(n40622) );
  NOR U53566 ( .A(n40622), .B(n40621), .Z(n44005) );
  NOR U53567 ( .A(n44012), .B(n44005), .Z(n40623) );
  XOR U53568 ( .A(n44004), .B(n40623), .Z(n44011) );
  XOR U53569 ( .A(n44009), .B(n44011), .Z(n47561) );
  XOR U53570 ( .A(n47563), .B(n47561), .Z(n44018) );
  IV U53571 ( .A(n40624), .Z(n40629) );
  NOR U53572 ( .A(n40626), .B(n40625), .Z(n40627) );
  IV U53573 ( .A(n40627), .Z(n40628) );
  NOR U53574 ( .A(n40629), .B(n40628), .Z(n40630) );
  IV U53575 ( .A(n40630), .Z(n44019) );
  XOR U53576 ( .A(n44018), .B(n44019), .Z(n41600) );
  XOR U53577 ( .A(n41601), .B(n41600), .Z(n40631) );
  IV U53578 ( .A(n40631), .Z(n41598) );
  NOR U53579 ( .A(n40638), .B(n41598), .Z(n47582) );
  NOR U53580 ( .A(n40633), .B(n40632), .Z(n40634) );
  IV U53581 ( .A(n40634), .Z(n41596) );
  IV U53582 ( .A(n40635), .Z(n40636) );
  NOR U53583 ( .A(n40637), .B(n40636), .Z(n41597) );
  XOR U53584 ( .A(n41597), .B(n41598), .Z(n41595) );
  XOR U53585 ( .A(n41596), .B(n41595), .Z(n40641) );
  IV U53586 ( .A(n41595), .Z(n40639) );
  NOR U53587 ( .A(n40639), .B(n40638), .Z(n40640) );
  NOR U53588 ( .A(n40641), .B(n40640), .Z(n40642) );
  NOR U53589 ( .A(n47582), .B(n40642), .Z(n40643) );
  IV U53590 ( .A(n40643), .Z(n41593) );
  XOR U53591 ( .A(n41593), .B(n41592), .Z(n44029) );
  XOR U53592 ( .A(n44027), .B(n44029), .Z(n44031) );
  XOR U53593 ( .A(n44030), .B(n44031), .Z(n44037) );
  IV U53594 ( .A(n40644), .Z(n40645) );
  NOR U53595 ( .A(n40646), .B(n40645), .Z(n41590) );
  IV U53596 ( .A(n40647), .Z(n40649) );
  NOR U53597 ( .A(n40649), .B(n40648), .Z(n44035) );
  NOR U53598 ( .A(n41590), .B(n44035), .Z(n40650) );
  XOR U53599 ( .A(n44037), .B(n40650), .Z(n41584) );
  XOR U53600 ( .A(n41585), .B(n41584), .Z(n41587) );
  XOR U53601 ( .A(n40651), .B(n41587), .Z(n40652) );
  IV U53602 ( .A(n40652), .Z(n44041) );
  IV U53603 ( .A(n40653), .Z(n40654) );
  NOR U53604 ( .A(n40654), .B(n44044), .Z(n41580) );
  XOR U53605 ( .A(n44041), .B(n41580), .Z(n44053) );
  IV U53606 ( .A(n44053), .Z(n40662) );
  IV U53607 ( .A(n40655), .Z(n40665) );
  IV U53608 ( .A(n40656), .Z(n40657) );
  NOR U53609 ( .A(n40665), .B(n40657), .Z(n44051) );
  IV U53610 ( .A(n40658), .Z(n40659) );
  NOR U53611 ( .A(n44044), .B(n40659), .Z(n40660) );
  NOR U53612 ( .A(n44051), .B(n40660), .Z(n40661) );
  XOR U53613 ( .A(n40662), .B(n40661), .Z(n44050) );
  IV U53614 ( .A(n40663), .Z(n40664) );
  NOR U53615 ( .A(n40665), .B(n40664), .Z(n44048) );
  XOR U53616 ( .A(n44050), .B(n44048), .Z(n44056) );
  XOR U53617 ( .A(n44055), .B(n44056), .Z(n44059) );
  XOR U53618 ( .A(n44058), .B(n44059), .Z(n44064) );
  XOR U53619 ( .A(n44062), .B(n44064), .Z(n44066) );
  XOR U53620 ( .A(n44065), .B(n44066), .Z(n44071) );
  XOR U53621 ( .A(n40666), .B(n44071), .Z(n41575) );
  XOR U53622 ( .A(n40667), .B(n41575), .Z(n45062) );
  XOR U53623 ( .A(n44073), .B(n45062), .Z(n40676) );
  IV U53624 ( .A(n40668), .Z(n40669) );
  NOR U53625 ( .A(n40670), .B(n40669), .Z(n40671) );
  NOR U53626 ( .A(n40676), .B(n40671), .Z(n41566) );
  IV U53627 ( .A(n40671), .Z(n40672) );
  NOR U53628 ( .A(n45062), .B(n40672), .Z(n48438) );
  NOR U53629 ( .A(n41566), .B(n48438), .Z(n40673) );
  IV U53630 ( .A(n40673), .Z(n50981) );
  NOR U53631 ( .A(n40674), .B(n50981), .Z(n40678) );
  IV U53632 ( .A(n40674), .Z(n40675) );
  NOR U53633 ( .A(n40676), .B(n40675), .Z(n40677) );
  NOR U53634 ( .A(n40678), .B(n40677), .Z(n44087) );
  IV U53635 ( .A(n40679), .Z(n40681) );
  NOR U53636 ( .A(n40681), .B(n40680), .Z(n44085) );
  NOR U53637 ( .A(n44080), .B(n44085), .Z(n40682) );
  XOR U53638 ( .A(n44087), .B(n40682), .Z(n40683) );
  IV U53639 ( .A(n40683), .Z(n44084) );
  IV U53640 ( .A(n40684), .Z(n40687) );
  IV U53641 ( .A(n40685), .Z(n40686) );
  NOR U53642 ( .A(n40687), .B(n40686), .Z(n44082) );
  XOR U53643 ( .A(n44084), .B(n44082), .Z(n41564) );
  IV U53644 ( .A(n41564), .Z(n40695) );
  IV U53645 ( .A(n40688), .Z(n40689) );
  NOR U53646 ( .A(n40690), .B(n40689), .Z(n41563) );
  IV U53647 ( .A(n40691), .Z(n40693) );
  NOR U53648 ( .A(n40693), .B(n40692), .Z(n41561) );
  NOR U53649 ( .A(n41563), .B(n41561), .Z(n40694) );
  XOR U53650 ( .A(n40695), .B(n40694), .Z(n41557) );
  XOR U53651 ( .A(n41555), .B(n41557), .Z(n41559) );
  XOR U53652 ( .A(n41558), .B(n41559), .Z(n41553) );
  XOR U53653 ( .A(n41552), .B(n41553), .Z(n44097) );
  XOR U53654 ( .A(n40696), .B(n44097), .Z(n44099) );
  IV U53655 ( .A(n40697), .Z(n40698) );
  NOR U53656 ( .A(n40698), .B(n40704), .Z(n44100) );
  XOR U53657 ( .A(n44099), .B(n44100), .Z(n41549) );
  IV U53658 ( .A(n40699), .Z(n40700) );
  NOR U53659 ( .A(n40701), .B(n40700), .Z(n41548) );
  IV U53660 ( .A(n40702), .Z(n40703) );
  NOR U53661 ( .A(n40704), .B(n40703), .Z(n44103) );
  NOR U53662 ( .A(n41548), .B(n44103), .Z(n40705) );
  XOR U53663 ( .A(n41549), .B(n40705), .Z(n41547) );
  XOR U53664 ( .A(n41545), .B(n41547), .Z(n44107) );
  IV U53665 ( .A(n40706), .Z(n40708) );
  NOR U53666 ( .A(n40708), .B(n40707), .Z(n40709) );
  IV U53667 ( .A(n40709), .Z(n44106) );
  XOR U53668 ( .A(n44107), .B(n44106), .Z(n40710) );
  NOR U53669 ( .A(n40711), .B(n40710), .Z(n40721) );
  IV U53670 ( .A(n40712), .Z(n40715) );
  NOR U53671 ( .A(n40713), .B(n41547), .Z(n40714) );
  IV U53672 ( .A(n40714), .Z(n40717) );
  NOR U53673 ( .A(n40715), .B(n40717), .Z(n45011) );
  IV U53674 ( .A(n40716), .Z(n40718) );
  NOR U53675 ( .A(n40718), .B(n40717), .Z(n47638) );
  NOR U53676 ( .A(n45011), .B(n47638), .Z(n40719) );
  IV U53677 ( .A(n40719), .Z(n40720) );
  NOR U53678 ( .A(n40721), .B(n40720), .Z(n44110) );
  XOR U53679 ( .A(n44111), .B(n44110), .Z(n41543) );
  IV U53680 ( .A(n41543), .Z(n40730) );
  IV U53681 ( .A(n40722), .Z(n40723) );
  NOR U53682 ( .A(n40724), .B(n40723), .Z(n41536) );
  NOR U53683 ( .A(n40725), .B(n41539), .Z(n40726) );
  NOR U53684 ( .A(n40726), .B(n41542), .Z(n40727) );
  IV U53685 ( .A(n40727), .Z(n40728) );
  NOR U53686 ( .A(n41536), .B(n40728), .Z(n40729) );
  XOR U53687 ( .A(n40730), .B(n40729), .Z(n44119) );
  IV U53688 ( .A(n40731), .Z(n40734) );
  IV U53689 ( .A(n40732), .Z(n40733) );
  NOR U53690 ( .A(n40734), .B(n40733), .Z(n44117) );
  XOR U53691 ( .A(n44119), .B(n44117), .Z(n44121) );
  XOR U53692 ( .A(n44120), .B(n44121), .Z(n40741) );
  NOR U53693 ( .A(n40735), .B(n40741), .Z(n45002) );
  IV U53694 ( .A(n40736), .Z(n40737) );
  NOR U53695 ( .A(n40738), .B(n40737), .Z(n40742) );
  IV U53696 ( .A(n40742), .Z(n40739) );
  NOR U53697 ( .A(n40739), .B(n44121), .Z(n45000) );
  NOR U53698 ( .A(n45002), .B(n45000), .Z(n40740) );
  IV U53699 ( .A(n40740), .Z(n44126) );
  NOR U53700 ( .A(n44126), .B(n40741), .Z(n40746) );
  NOR U53701 ( .A(n40743), .B(n40742), .Z(n40744) );
  NOR U53702 ( .A(n40744), .B(n44126), .Z(n40745) );
  NOR U53703 ( .A(n40746), .B(n40745), .Z(n44124) );
  XOR U53704 ( .A(n44125), .B(n44124), .Z(n40753) );
  IV U53705 ( .A(n40753), .Z(n40747) );
  NOR U53706 ( .A(n40748), .B(n40747), .Z(n47662) );
  IV U53707 ( .A(n40749), .Z(n40751) );
  NOR U53708 ( .A(n40751), .B(n40750), .Z(n40754) );
  IV U53709 ( .A(n40754), .Z(n40752) );
  NOR U53710 ( .A(n40752), .B(n44124), .Z(n41535) );
  NOR U53711 ( .A(n40754), .B(n40753), .Z(n40755) );
  NOR U53712 ( .A(n41535), .B(n40755), .Z(n40756) );
  NOR U53713 ( .A(n40757), .B(n40756), .Z(n40758) );
  NOR U53714 ( .A(n47662), .B(n40758), .Z(n40759) );
  IV U53715 ( .A(n40759), .Z(n44129) );
  XOR U53716 ( .A(n44128), .B(n44129), .Z(n41531) );
  IV U53717 ( .A(n40760), .Z(n40762) );
  NOR U53718 ( .A(n40762), .B(n40761), .Z(n41533) );
  IV U53719 ( .A(n40763), .Z(n40764) );
  NOR U53720 ( .A(n40765), .B(n40764), .Z(n41530) );
  NOR U53721 ( .A(n41533), .B(n41530), .Z(n40766) );
  XOR U53722 ( .A(n41531), .B(n40766), .Z(n41522) );
  IV U53723 ( .A(n40767), .Z(n40769) );
  NOR U53724 ( .A(n40769), .B(n40768), .Z(n41527) );
  IV U53725 ( .A(n40770), .Z(n40772) );
  NOR U53726 ( .A(n40772), .B(n40771), .Z(n41523) );
  NOR U53727 ( .A(n41527), .B(n41523), .Z(n40773) );
  XOR U53728 ( .A(n41522), .B(n40773), .Z(n44982) );
  NOR U53729 ( .A(n40775), .B(n40774), .Z(n44985) );
  IV U53730 ( .A(n40776), .Z(n40777) );
  NOR U53731 ( .A(n40778), .B(n40777), .Z(n44981) );
  NOR U53732 ( .A(n44985), .B(n44981), .Z(n41526) );
  XOR U53733 ( .A(n44982), .B(n41526), .Z(n44134) );
  XOR U53734 ( .A(n44135), .B(n44134), .Z(n44144) );
  XOR U53735 ( .A(n40779), .B(n44144), .Z(n40780) );
  IV U53736 ( .A(n40780), .Z(n41520) );
  XOR U53737 ( .A(n41518), .B(n41520), .Z(n44140) );
  XOR U53738 ( .A(n44139), .B(n44140), .Z(n44155) );
  XOR U53739 ( .A(n44152), .B(n44155), .Z(n44162) );
  IV U53740 ( .A(n40781), .Z(n40782) );
  NOR U53741 ( .A(n40783), .B(n40782), .Z(n44154) );
  IV U53742 ( .A(n40784), .Z(n40786) );
  NOR U53743 ( .A(n40786), .B(n40785), .Z(n44161) );
  NOR U53744 ( .A(n44154), .B(n44161), .Z(n40787) );
  XOR U53745 ( .A(n44162), .B(n40787), .Z(n44158) );
  IV U53746 ( .A(n40788), .Z(n40789) );
  NOR U53747 ( .A(n40789), .B(n44168), .Z(n44172) );
  IV U53748 ( .A(n40790), .Z(n40791) );
  NOR U53749 ( .A(n40791), .B(n40793), .Z(n44165) );
  IV U53750 ( .A(n40792), .Z(n40794) );
  NOR U53751 ( .A(n40794), .B(n40793), .Z(n44159) );
  NOR U53752 ( .A(n44165), .B(n44159), .Z(n40795) );
  IV U53753 ( .A(n40795), .Z(n40796) );
  NOR U53754 ( .A(n44172), .B(n40796), .Z(n40797) );
  XOR U53755 ( .A(n44158), .B(n40797), .Z(n44179) );
  NOR U53756 ( .A(n40798), .B(n40803), .Z(n44177) );
  XOR U53757 ( .A(n44179), .B(n44177), .Z(n41517) );
  IV U53758 ( .A(n41517), .Z(n40806) );
  IV U53759 ( .A(n40799), .Z(n40800) );
  NOR U53760 ( .A(n40801), .B(n40800), .Z(n41513) );
  IV U53761 ( .A(n40802), .Z(n40804) );
  NOR U53762 ( .A(n40804), .B(n40803), .Z(n41515) );
  NOR U53763 ( .A(n41513), .B(n41515), .Z(n40805) );
  XOR U53764 ( .A(n40806), .B(n40805), .Z(n44183) );
  XOR U53765 ( .A(n41510), .B(n44183), .Z(n41507) );
  XOR U53766 ( .A(n40807), .B(n41507), .Z(n40808) );
  IV U53767 ( .A(n40808), .Z(n41502) );
  XOR U53768 ( .A(n41500), .B(n41502), .Z(n41504) );
  IV U53769 ( .A(n41504), .Z(n40815) );
  IV U53770 ( .A(n40809), .Z(n40811) );
  NOR U53771 ( .A(n40811), .B(n40810), .Z(n41503) );
  IV U53772 ( .A(n40812), .Z(n40813) );
  NOR U53773 ( .A(n40813), .B(n40817), .Z(n41497) );
  NOR U53774 ( .A(n41503), .B(n41497), .Z(n40814) );
  XOR U53775 ( .A(n40815), .B(n40814), .Z(n44205) );
  IV U53776 ( .A(n40816), .Z(n40818) );
  NOR U53777 ( .A(n40818), .B(n40817), .Z(n44203) );
  XOR U53778 ( .A(n44205), .B(n44203), .Z(n44207) );
  XOR U53779 ( .A(n44206), .B(n44207), .Z(n44218) );
  XOR U53780 ( .A(n44217), .B(n44218), .Z(n44211) );
  XOR U53781 ( .A(n44210), .B(n44211), .Z(n44226) );
  XOR U53782 ( .A(n44214), .B(n44226), .Z(n44230) );
  XOR U53783 ( .A(n40819), .B(n44230), .Z(n40820) );
  IV U53784 ( .A(n40820), .Z(n44234) );
  XOR U53785 ( .A(n44232), .B(n44234), .Z(n44236) );
  IV U53786 ( .A(n44236), .Z(n40828) );
  IV U53787 ( .A(n40821), .Z(n40822) );
  NOR U53788 ( .A(n40823), .B(n40822), .Z(n44235) );
  IV U53789 ( .A(n40824), .Z(n40826) );
  NOR U53790 ( .A(n40826), .B(n40825), .Z(n41494) );
  NOR U53791 ( .A(n44235), .B(n41494), .Z(n40827) );
  XOR U53792 ( .A(n40828), .B(n40827), .Z(n44242) );
  XOR U53793 ( .A(n44240), .B(n44242), .Z(n44249) );
  XOR U53794 ( .A(n41491), .B(n44249), .Z(n44255) );
  XOR U53795 ( .A(n40829), .B(n44255), .Z(n44263) );
  XOR U53796 ( .A(n40830), .B(n44263), .Z(n41485) );
  XOR U53797 ( .A(n40831), .B(n41485), .Z(n41472) );
  IV U53798 ( .A(n40832), .Z(n40833) );
  NOR U53799 ( .A(n40834), .B(n40833), .Z(n40835) );
  XOR U53800 ( .A(n41472), .B(n40835), .Z(n41468) );
  XOR U53801 ( .A(n41466), .B(n41468), .Z(n44270) );
  XOR U53802 ( .A(n40836), .B(n44270), .Z(n44265) );
  XOR U53803 ( .A(n40837), .B(n44265), .Z(n44279) );
  XOR U53804 ( .A(n44275), .B(n44279), .Z(n44284) );
  XOR U53805 ( .A(n40838), .B(n44284), .Z(n41460) );
  XOR U53806 ( .A(n40839), .B(n41460), .Z(n41458) );
  XOR U53807 ( .A(n41459), .B(n41458), .Z(n40846) );
  IV U53808 ( .A(n40846), .Z(n40840) );
  NOR U53809 ( .A(n40841), .B(n40840), .Z(n44898) );
  IV U53810 ( .A(n40842), .Z(n40844) );
  NOR U53811 ( .A(n40844), .B(n40843), .Z(n40847) );
  IV U53812 ( .A(n40847), .Z(n40845) );
  NOR U53813 ( .A(n40845), .B(n41458), .Z(n44903) );
  NOR U53814 ( .A(n40847), .B(n40846), .Z(n40848) );
  NOR U53815 ( .A(n44903), .B(n40848), .Z(n40849) );
  NOR U53816 ( .A(n40850), .B(n40849), .Z(n40851) );
  NOR U53817 ( .A(n44898), .B(n40851), .Z(n40853) );
  NOR U53818 ( .A(n40852), .B(n40853), .Z(n44289) );
  IV U53819 ( .A(n40852), .Z(n40855) );
  IV U53820 ( .A(n40853), .Z(n40854) );
  NOR U53821 ( .A(n40855), .B(n40854), .Z(n54685) );
  NOR U53822 ( .A(n44289), .B(n54685), .Z(n44294) );
  IV U53823 ( .A(n40856), .Z(n40857) );
  NOR U53824 ( .A(n40857), .B(n40859), .Z(n44287) );
  IV U53825 ( .A(n40858), .Z(n40862) );
  XOR U53826 ( .A(n40860), .B(n40859), .Z(n40861) );
  NOR U53827 ( .A(n40862), .B(n40861), .Z(n44295) );
  NOR U53828 ( .A(n44287), .B(n44295), .Z(n40863) );
  XOR U53829 ( .A(n44294), .B(n40863), .Z(n44293) );
  IV U53830 ( .A(n40864), .Z(n40867) );
  IV U53831 ( .A(n40865), .Z(n40866) );
  NOR U53832 ( .A(n40867), .B(n40866), .Z(n44291) );
  XOR U53833 ( .A(n44293), .B(n44291), .Z(n40870) );
  NOR U53834 ( .A(n40868), .B(n40870), .Z(n51153) );
  NOR U53835 ( .A(n40869), .B(n41455), .Z(n40871) );
  XOR U53836 ( .A(n40871), .B(n40870), .Z(n40881) );
  IV U53837 ( .A(n40881), .Z(n40872) );
  NOR U53838 ( .A(n40873), .B(n40872), .Z(n40874) );
  NOR U53839 ( .A(n51153), .B(n40874), .Z(n44303) );
  IV U53840 ( .A(n40875), .Z(n40877) );
  NOR U53841 ( .A(n40877), .B(n40876), .Z(n40887) );
  IV U53842 ( .A(n40887), .Z(n44305) );
  NOR U53843 ( .A(n44303), .B(n44305), .Z(n40889) );
  IV U53844 ( .A(n40878), .Z(n40880) );
  NOR U53845 ( .A(n40880), .B(n40879), .Z(n40883) );
  IV U53846 ( .A(n40883), .Z(n40882) );
  NOR U53847 ( .A(n40882), .B(n40881), .Z(n51161) );
  NOR U53848 ( .A(n44303), .B(n40883), .Z(n40884) );
  NOR U53849 ( .A(n51161), .B(n40884), .Z(n40885) );
  IV U53850 ( .A(n40885), .Z(n40886) );
  NOR U53851 ( .A(n40887), .B(n40886), .Z(n40888) );
  NOR U53852 ( .A(n40889), .B(n40888), .Z(n44310) );
  XOR U53853 ( .A(n44306), .B(n44310), .Z(n41452) );
  XOR U53854 ( .A(n40890), .B(n41452), .Z(n41443) );
  XOR U53855 ( .A(n40891), .B(n41443), .Z(n41441) );
  XOR U53856 ( .A(n40892), .B(n41441), .Z(n41428) );
  XOR U53857 ( .A(n40893), .B(n41428), .Z(n44316) );
  XOR U53858 ( .A(n44314), .B(n44316), .Z(n44319) );
  XOR U53859 ( .A(n44317), .B(n44319), .Z(n41425) );
  XOR U53860 ( .A(n41426), .B(n41425), .Z(n40903) );
  IV U53861 ( .A(n40903), .Z(n40898) );
  IV U53862 ( .A(n40894), .Z(n40896) );
  NOR U53863 ( .A(n40896), .B(n40895), .Z(n40907) );
  IV U53864 ( .A(n40907), .Z(n40897) );
  NOR U53865 ( .A(n40898), .B(n40897), .Z(n44886) );
  IV U53866 ( .A(n40899), .Z(n40901) );
  NOR U53867 ( .A(n40901), .B(n40900), .Z(n40904) );
  IV U53868 ( .A(n40904), .Z(n40902) );
  NOR U53869 ( .A(n40902), .B(n41425), .Z(n47838) );
  NOR U53870 ( .A(n40904), .B(n40903), .Z(n40905) );
  NOR U53871 ( .A(n47838), .B(n40905), .Z(n40906) );
  NOR U53872 ( .A(n40907), .B(n40906), .Z(n40908) );
  NOR U53873 ( .A(n44886), .B(n40908), .Z(n41417) );
  XOR U53874 ( .A(n41422), .B(n41417), .Z(n41410) );
  XOR U53875 ( .A(n40909), .B(n41410), .Z(n41406) );
  XOR U53876 ( .A(n41404), .B(n41406), .Z(n44872) );
  IV U53877 ( .A(n44872), .Z(n40916) );
  IV U53878 ( .A(n40910), .Z(n40911) );
  NOR U53879 ( .A(n40912), .B(n40911), .Z(n44871) );
  IV U53880 ( .A(n40913), .Z(n40915) );
  NOR U53881 ( .A(n40915), .B(n40914), .Z(n47844) );
  NOR U53882 ( .A(n44871), .B(n47844), .Z(n41400) );
  XOR U53883 ( .A(n40916), .B(n41400), .Z(n41402) );
  XOR U53884 ( .A(n41401), .B(n41402), .Z(n44330) );
  XOR U53885 ( .A(n44329), .B(n44330), .Z(n41398) );
  NOR U53886 ( .A(n40924), .B(n41398), .Z(n47847) );
  IV U53887 ( .A(n40917), .Z(n40919) );
  NOR U53888 ( .A(n40919), .B(n40918), .Z(n40920) );
  IV U53889 ( .A(n40920), .Z(n44342) );
  IV U53890 ( .A(n40921), .Z(n40922) );
  NOR U53891 ( .A(n40923), .B(n40922), .Z(n41397) );
  XOR U53892 ( .A(n41397), .B(n41398), .Z(n44341) );
  XOR U53893 ( .A(n44342), .B(n44341), .Z(n40927) );
  IV U53894 ( .A(n44341), .Z(n40925) );
  NOR U53895 ( .A(n40925), .B(n40924), .Z(n40926) );
  NOR U53896 ( .A(n40927), .B(n40926), .Z(n40928) );
  NOR U53897 ( .A(n47847), .B(n40928), .Z(n41395) );
  IV U53898 ( .A(n40929), .Z(n40930) );
  NOR U53899 ( .A(n40931), .B(n40930), .Z(n44343) );
  IV U53900 ( .A(n40932), .Z(n40934) );
  NOR U53901 ( .A(n40934), .B(n40933), .Z(n41394) );
  NOR U53902 ( .A(n44343), .B(n41394), .Z(n40935) );
  XOR U53903 ( .A(n41395), .B(n40935), .Z(n41393) );
  XOR U53904 ( .A(n41391), .B(n41393), .Z(n41390) );
  IV U53905 ( .A(n40936), .Z(n40940) );
  IV U53906 ( .A(n40937), .Z(n40949) );
  NOR U53907 ( .A(n40949), .B(n40938), .Z(n40939) );
  IV U53908 ( .A(n40939), .Z(n40942) );
  NOR U53909 ( .A(n40940), .B(n40942), .Z(n41388) );
  XOR U53910 ( .A(n41390), .B(n41388), .Z(n41385) );
  IV U53911 ( .A(n40941), .Z(n40943) );
  NOR U53912 ( .A(n40943), .B(n40942), .Z(n41383) );
  XOR U53913 ( .A(n41385), .B(n41383), .Z(n44349) );
  IV U53914 ( .A(n44349), .Z(n40951) );
  IV U53915 ( .A(n40944), .Z(n40946) );
  NOR U53916 ( .A(n40946), .B(n40945), .Z(n44348) );
  IV U53917 ( .A(n40947), .Z(n40948) );
  NOR U53918 ( .A(n40949), .B(n40948), .Z(n41386) );
  NOR U53919 ( .A(n44348), .B(n41386), .Z(n40950) );
  XOR U53920 ( .A(n40951), .B(n40950), .Z(n44353) );
  XOR U53921 ( .A(n44351), .B(n44353), .Z(n44355) );
  XOR U53922 ( .A(n44354), .B(n44355), .Z(n41382) );
  XOR U53923 ( .A(n41380), .B(n41382), .Z(n41376) );
  XOR U53924 ( .A(n40952), .B(n41376), .Z(n40953) );
  IV U53925 ( .A(n40953), .Z(n41371) );
  XOR U53926 ( .A(n41369), .B(n41371), .Z(n44362) );
  XOR U53927 ( .A(n40954), .B(n44362), .Z(n41362) );
  IV U53928 ( .A(n40955), .Z(n40957) );
  NOR U53929 ( .A(n40957), .B(n40956), .Z(n44361) );
  IV U53930 ( .A(n40958), .Z(n40959) );
  NOR U53931 ( .A(n40960), .B(n40959), .Z(n41361) );
  NOR U53932 ( .A(n44361), .B(n41361), .Z(n40961) );
  XOR U53933 ( .A(n41362), .B(n40961), .Z(n44364) );
  XOR U53934 ( .A(n44365), .B(n44364), .Z(n44372) );
  IV U53935 ( .A(n40962), .Z(n40964) );
  NOR U53936 ( .A(n40964), .B(n40963), .Z(n44367) );
  IV U53937 ( .A(n40965), .Z(n40967) );
  NOR U53938 ( .A(n40967), .B(n40966), .Z(n44371) );
  NOR U53939 ( .A(n44367), .B(n44371), .Z(n40968) );
  XOR U53940 ( .A(n44372), .B(n40968), .Z(n44380) );
  XOR U53941 ( .A(n44378), .B(n44380), .Z(n41358) );
  XOR U53942 ( .A(n41357), .B(n41358), .Z(n44387) );
  IV U53943 ( .A(n44387), .Z(n40974) );
  IV U53944 ( .A(n40969), .Z(n40970) );
  NOR U53945 ( .A(n40971), .B(n40970), .Z(n44375) );
  NOR U53946 ( .A(n40972), .B(n40976), .Z(n44386) );
  NOR U53947 ( .A(n44375), .B(n44386), .Z(n40973) );
  XOR U53948 ( .A(n40974), .B(n40973), .Z(n44392) );
  IV U53949 ( .A(n40975), .Z(n40977) );
  NOR U53950 ( .A(n40977), .B(n40976), .Z(n44390) );
  XOR U53951 ( .A(n44392), .B(n44390), .Z(n44394) );
  XOR U53952 ( .A(n44393), .B(n44394), .Z(n41355) );
  XOR U53953 ( .A(n40978), .B(n41355), .Z(n41351) );
  IV U53954 ( .A(n40979), .Z(n40981) );
  NOR U53955 ( .A(n40981), .B(n40980), .Z(n41349) );
  XOR U53956 ( .A(n41351), .B(n41349), .Z(n41339) );
  IV U53957 ( .A(n40982), .Z(n40985) );
  IV U53958 ( .A(n40983), .Z(n40988) );
  XOR U53959 ( .A(n40988), .B(n40986), .Z(n40984) );
  NOR U53960 ( .A(n40985), .B(n40984), .Z(n41337) );
  IV U53961 ( .A(n40986), .Z(n41341) );
  IV U53962 ( .A(n40987), .Z(n41343) );
  NOR U53963 ( .A(n41341), .B(n41343), .Z(n40990) );
  NOR U53964 ( .A(n41341), .B(n40988), .Z(n40989) );
  NOR U53965 ( .A(n40990), .B(n40989), .Z(n40991) );
  IV U53966 ( .A(n40991), .Z(n40992) );
  NOR U53967 ( .A(n41337), .B(n40992), .Z(n40993) );
  XOR U53968 ( .A(n41339), .B(n40993), .Z(n40994) );
  IV U53969 ( .A(n40994), .Z(n41336) );
  IV U53970 ( .A(n40995), .Z(n40997) );
  NOR U53971 ( .A(n40997), .B(n40996), .Z(n40998) );
  IV U53972 ( .A(n40998), .Z(n41335) );
  XOR U53973 ( .A(n41336), .B(n41335), .Z(n41005) );
  IV U53974 ( .A(n41005), .Z(n40999) );
  NOR U53975 ( .A(n41000), .B(n40999), .Z(n44820) );
  IV U53976 ( .A(n41001), .Z(n41003) );
  NOR U53977 ( .A(n41003), .B(n41002), .Z(n41006) );
  IV U53978 ( .A(n41006), .Z(n41004) );
  NOR U53979 ( .A(n41336), .B(n41004), .Z(n44816) );
  NOR U53980 ( .A(n41006), .B(n41005), .Z(n41007) );
  NOR U53981 ( .A(n44816), .B(n41007), .Z(n41329) );
  NOR U53982 ( .A(n41008), .B(n41329), .Z(n41009) );
  NOR U53983 ( .A(n44820), .B(n41009), .Z(n41010) );
  IV U53984 ( .A(n41010), .Z(n41326) );
  IV U53985 ( .A(n41011), .Z(n41334) );
  NOR U53986 ( .A(n41334), .B(n41327), .Z(n41015) );
  IV U53987 ( .A(n41012), .Z(n41014) );
  IV U53988 ( .A(n41013), .Z(n41022) );
  NOR U53989 ( .A(n41014), .B(n41022), .Z(n41324) );
  NOR U53990 ( .A(n41015), .B(n41324), .Z(n41016) );
  XOR U53991 ( .A(n41326), .B(n41016), .Z(n41318) );
  IV U53992 ( .A(n41017), .Z(n41018) );
  NOR U53993 ( .A(n41019), .B(n41018), .Z(n41319) );
  IV U53994 ( .A(n41020), .Z(n41021) );
  NOR U53995 ( .A(n41022), .B(n41021), .Z(n41321) );
  NOR U53996 ( .A(n41319), .B(n41321), .Z(n41023) );
  XOR U53997 ( .A(n41318), .B(n41023), .Z(n44405) );
  XOR U53998 ( .A(n44404), .B(n44405), .Z(n41317) );
  IV U53999 ( .A(n41024), .Z(n41026) );
  NOR U54000 ( .A(n41026), .B(n41025), .Z(n41315) );
  XOR U54001 ( .A(n41317), .B(n41315), .Z(n41313) );
  XOR U54002 ( .A(n41312), .B(n41313), .Z(n44430) );
  IV U54003 ( .A(n44430), .Z(n41034) );
  IV U54004 ( .A(n41027), .Z(n41028) );
  NOR U54005 ( .A(n41029), .B(n41028), .Z(n44425) );
  IV U54006 ( .A(n41030), .Z(n41032) );
  NOR U54007 ( .A(n41032), .B(n41031), .Z(n44428) );
  NOR U54008 ( .A(n44425), .B(n44428), .Z(n41033) );
  XOR U54009 ( .A(n41034), .B(n41033), .Z(n44420) );
  XOR U54010 ( .A(n41307), .B(n44420), .Z(n41302) );
  XOR U54011 ( .A(n41035), .B(n41302), .Z(n41294) );
  XOR U54012 ( .A(n41036), .B(n41294), .Z(n48204) );
  XOR U54013 ( .A(n41290), .B(n48204), .Z(n41037) );
  IV U54014 ( .A(n41037), .Z(n41293) );
  IV U54015 ( .A(n41038), .Z(n41040) );
  NOR U54016 ( .A(n41040), .B(n41039), .Z(n41291) );
  XOR U54017 ( .A(n41293), .B(n41291), .Z(n44442) );
  IV U54018 ( .A(n44442), .Z(n41048) );
  IV U54019 ( .A(n41041), .Z(n41042) );
  NOR U54020 ( .A(n41043), .B(n41042), .Z(n44438) );
  IV U54021 ( .A(n41044), .Z(n41045) );
  NOR U54022 ( .A(n41046), .B(n41045), .Z(n44441) );
  NOR U54023 ( .A(n44438), .B(n44441), .Z(n41047) );
  XOR U54024 ( .A(n41048), .B(n41047), .Z(n44448) );
  IV U54025 ( .A(n41049), .Z(n41051) );
  NOR U54026 ( .A(n41051), .B(n41050), .Z(n41288) );
  XOR U54027 ( .A(n44448), .B(n41288), .Z(n41052) );
  XOR U54028 ( .A(n41053), .B(n41052), .Z(n44449) );
  XOR U54029 ( .A(n41054), .B(n44449), .Z(n44461) );
  XOR U54030 ( .A(n41055), .B(n44461), .Z(n41287) );
  XOR U54031 ( .A(n41056), .B(n41287), .Z(n41057) );
  IV U54032 ( .A(n41057), .Z(n44470) );
  IV U54033 ( .A(n41058), .Z(n41059) );
  NOR U54034 ( .A(n41059), .B(n41063), .Z(n44468) );
  XOR U54035 ( .A(n44470), .B(n44468), .Z(n44473) );
  IV U54036 ( .A(n44473), .Z(n41067) );
  IV U54037 ( .A(n41060), .Z(n41274) );
  NOR U54038 ( .A(n41274), .B(n41061), .Z(n41065) );
  IV U54039 ( .A(n41062), .Z(n41064) );
  NOR U54040 ( .A(n41064), .B(n41063), .Z(n44471) );
  NOR U54041 ( .A(n41065), .B(n44471), .Z(n41066) );
  XOR U54042 ( .A(n41067), .B(n41066), .Z(n41269) );
  IV U54043 ( .A(n41068), .Z(n41070) );
  NOR U54044 ( .A(n41070), .B(n41069), .Z(n41267) );
  XOR U54045 ( .A(n41269), .B(n41267), .Z(n41271) );
  XOR U54046 ( .A(n41270), .B(n41271), .Z(n44479) );
  NOR U54047 ( .A(n41076), .B(n44479), .Z(n47984) );
  NOR U54048 ( .A(n41072), .B(n41071), .Z(n44478) );
  XOR U54049 ( .A(n44478), .B(n44479), .Z(n44485) );
  IV U54050 ( .A(n41073), .Z(n41075) );
  NOR U54051 ( .A(n41075), .B(n41074), .Z(n41077) );
  IV U54052 ( .A(n41077), .Z(n44484) );
  XOR U54053 ( .A(n44485), .B(n44484), .Z(n41079) );
  NOR U54054 ( .A(n41077), .B(n41076), .Z(n41078) );
  NOR U54055 ( .A(n41079), .B(n41078), .Z(n41080) );
  NOR U54056 ( .A(n47984), .B(n41080), .Z(n41260) );
  XOR U54057 ( .A(n41081), .B(n41260), .Z(n41257) );
  IV U54058 ( .A(n41082), .Z(n41083) );
  NOR U54059 ( .A(n41084), .B(n41083), .Z(n41256) );
  IV U54060 ( .A(n41085), .Z(n41086) );
  NOR U54061 ( .A(n41087), .B(n41086), .Z(n41254) );
  NOR U54062 ( .A(n41256), .B(n41254), .Z(n41088) );
  XOR U54063 ( .A(n41257), .B(n41088), .Z(n41243) );
  NOR U54064 ( .A(n41089), .B(n41247), .Z(n41093) );
  IV U54065 ( .A(n41090), .Z(n41092) );
  IV U54066 ( .A(n41091), .Z(n41099) );
  NOR U54067 ( .A(n41092), .B(n41099), .Z(n41244) );
  NOR U54068 ( .A(n41093), .B(n41244), .Z(n41094) );
  XOR U54069 ( .A(n41243), .B(n41094), .Z(n41242) );
  IV U54070 ( .A(n41095), .Z(n41096) );
  NOR U54071 ( .A(n41097), .B(n41096), .Z(n41238) );
  IV U54072 ( .A(n41098), .Z(n41100) );
  NOR U54073 ( .A(n41100), .B(n41099), .Z(n41240) );
  NOR U54074 ( .A(n41238), .B(n41240), .Z(n41101) );
  XOR U54075 ( .A(n41242), .B(n41101), .Z(n41233) );
  XOR U54076 ( .A(n41102), .B(n41233), .Z(n41231) );
  XOR U54077 ( .A(n41103), .B(n41231), .Z(n41221) );
  XOR U54078 ( .A(n41222), .B(n41221), .Z(n41226) );
  XOR U54079 ( .A(n41224), .B(n41226), .Z(n41219) );
  NOR U54080 ( .A(n41111), .B(n41219), .Z(n44730) );
  IV U54081 ( .A(n41104), .Z(n41106) );
  NOR U54082 ( .A(n41106), .B(n41105), .Z(n41107) );
  IV U54083 ( .A(n41107), .Z(n41215) );
  IV U54084 ( .A(n41108), .Z(n41109) );
  NOR U54085 ( .A(n41110), .B(n41109), .Z(n41218) );
  XOR U54086 ( .A(n41218), .B(n41219), .Z(n41214) );
  XOR U54087 ( .A(n41215), .B(n41214), .Z(n41114) );
  IV U54088 ( .A(n41214), .Z(n41112) );
  NOR U54089 ( .A(n41112), .B(n41111), .Z(n41113) );
  NOR U54090 ( .A(n41114), .B(n41113), .Z(n41115) );
  NOR U54091 ( .A(n44730), .B(n41115), .Z(n41211) );
  XOR U54092 ( .A(n41216), .B(n41211), .Z(n41209) );
  XOR U54093 ( .A(n41116), .B(n41209), .Z(n41117) );
  IV U54094 ( .A(n41117), .Z(n44497) );
  XOR U54095 ( .A(n44495), .B(n44497), .Z(n44499) );
  IV U54096 ( .A(n44499), .Z(n41122) );
  IV U54097 ( .A(n41118), .Z(n41119) );
  NOR U54098 ( .A(n41120), .B(n41119), .Z(n41206) );
  NOR U54099 ( .A(n44498), .B(n41206), .Z(n41121) );
  XOR U54100 ( .A(n41122), .B(n41121), .Z(n41205) );
  XOR U54101 ( .A(n41201), .B(n41205), .Z(n44505) );
  XOR U54102 ( .A(n41123), .B(n44505), .Z(n41124) );
  IV U54103 ( .A(n41124), .Z(n41200) );
  XOR U54104 ( .A(n41198), .B(n41200), .Z(n48026) );
  IV U54105 ( .A(n41125), .Z(n41126) );
  NOR U54106 ( .A(n41127), .B(n41126), .Z(n48024) );
  IV U54107 ( .A(n41128), .Z(n41130) );
  NOR U54108 ( .A(n41130), .B(n41129), .Z(n48030) );
  NOR U54109 ( .A(n48024), .B(n48030), .Z(n44507) );
  XOR U54110 ( .A(n48026), .B(n44507), .Z(n44508) );
  XOR U54111 ( .A(n41131), .B(n44508), .Z(n44515) );
  XOR U54112 ( .A(n44513), .B(n44515), .Z(n41194) );
  XOR U54113 ( .A(n41193), .B(n41194), .Z(n41196) );
  XOR U54114 ( .A(n41197), .B(n41196), .Z(n41183) );
  IV U54115 ( .A(n41132), .Z(n41191) );
  NOR U54116 ( .A(n41133), .B(n41191), .Z(n41137) );
  IV U54117 ( .A(n41134), .Z(n41135) );
  NOR U54118 ( .A(n41136), .B(n41135), .Z(n41182) );
  NOR U54119 ( .A(n41137), .B(n41182), .Z(n41138) );
  XOR U54120 ( .A(n41183), .B(n41138), .Z(n41181) );
  IV U54121 ( .A(n41139), .Z(n41140) );
  NOR U54122 ( .A(n41141), .B(n41140), .Z(n41142) );
  IV U54123 ( .A(n41142), .Z(n41149) );
  NOR U54124 ( .A(n41181), .B(n41149), .Z(n51484) );
  IV U54125 ( .A(n41143), .Z(n41144) );
  NOR U54126 ( .A(n41167), .B(n41144), .Z(n41145) );
  IV U54127 ( .A(n41145), .Z(n44521) );
  IV U54128 ( .A(n41146), .Z(n41147) );
  NOR U54129 ( .A(n41148), .B(n41147), .Z(n41179) );
  XOR U54130 ( .A(n41179), .B(n41181), .Z(n44520) );
  XOR U54131 ( .A(n44521), .B(n44520), .Z(n41152) );
  IV U54132 ( .A(n44520), .Z(n41150) );
  NOR U54133 ( .A(n41150), .B(n41149), .Z(n41151) );
  NOR U54134 ( .A(n41152), .B(n41151), .Z(n41153) );
  NOR U54135 ( .A(n51484), .B(n41153), .Z(n41164) );
  IV U54136 ( .A(n41164), .Z(n44523) );
  IV U54137 ( .A(n41154), .Z(n41158) );
  NOR U54138 ( .A(n44562), .B(n44547), .Z(n41155) );
  IV U54139 ( .A(n41155), .Z(n41156) );
  NOR U54140 ( .A(n44583), .B(n41156), .Z(n41157) );
  IV U54141 ( .A(n41157), .Z(n41175) );
  NOR U54142 ( .A(n41158), .B(n41175), .Z(n41159) );
  IV U54143 ( .A(n41159), .Z(n41168) );
  NOR U54144 ( .A(n44523), .B(n41168), .Z(n44531) );
  IV U54145 ( .A(n41160), .Z(n41161) );
  NOR U54146 ( .A(n41162), .B(n41161), .Z(n41163) );
  IV U54147 ( .A(n41163), .Z(n44522) );
  XOR U54148 ( .A(n41164), .B(n44522), .Z(n44527) );
  IV U54149 ( .A(n41165), .Z(n41166) );
  NOR U54150 ( .A(n41167), .B(n41166), .Z(n41169) );
  IV U54151 ( .A(n41169), .Z(n44526) );
  XOR U54152 ( .A(n44527), .B(n44526), .Z(n41171) );
  NOR U54153 ( .A(n41169), .B(n41168), .Z(n41170) );
  NOR U54154 ( .A(n41171), .B(n41170), .Z(n41172) );
  NOR U54155 ( .A(n44531), .B(n41172), .Z(n44542) );
  IV U54156 ( .A(n44542), .Z(n41177) );
  NOR U54157 ( .A(n41173), .B(n41177), .Z(n44538) );
  IV U54158 ( .A(n44538), .Z(n44535) );
  IV U54159 ( .A(n41174), .Z(n41176) );
  NOR U54160 ( .A(n41176), .B(n41175), .Z(n44539) );
  IV U54161 ( .A(n44539), .Z(n41178) );
  NOR U54162 ( .A(n41178), .B(n41177), .Z(n44530) );
  IV U54163 ( .A(n44530), .Z(n44525) );
  IV U54164 ( .A(n41179), .Z(n41180) );
  NOR U54165 ( .A(n41181), .B(n41180), .Z(n48125) );
  NOR U54166 ( .A(n48125), .B(n51484), .Z(n48035) );
  IV U54167 ( .A(n41182), .Z(n41185) );
  IV U54168 ( .A(n41183), .Z(n41184) );
  NOR U54169 ( .A(n41185), .B(n41184), .Z(n44702) );
  XOR U54170 ( .A(n41187), .B(n41186), .Z(n41188) );
  NOR U54171 ( .A(n41188), .B(n41196), .Z(n41189) );
  IV U54172 ( .A(n41189), .Z(n41190) );
  NOR U54173 ( .A(n41191), .B(n41190), .Z(n41192) );
  IV U54174 ( .A(n41192), .Z(n44707) );
  IV U54175 ( .A(n41193), .Z(n41195) );
  NOR U54176 ( .A(n41195), .B(n41194), .Z(n51459) );
  NOR U54177 ( .A(n41197), .B(n41196), .Z(n48135) );
  NOR U54178 ( .A(n51459), .B(n48135), .Z(n44705) );
  IV U54179 ( .A(n41198), .Z(n41199) );
  NOR U54180 ( .A(n41200), .B(n41199), .Z(n48022) );
  IV U54181 ( .A(n41201), .Z(n41202) );
  NOR U54182 ( .A(n41202), .B(n41205), .Z(n51434) );
  IV U54183 ( .A(n41203), .Z(n41204) );
  NOR U54184 ( .A(n41205), .B(n41204), .Z(n51426) );
  NOR U54185 ( .A(n51434), .B(n51426), .Z(n48017) );
  IV U54186 ( .A(n41206), .Z(n41207) );
  NOR U54187 ( .A(n41207), .B(n44499), .Z(n44722) );
  IV U54188 ( .A(n41208), .Z(n41210) );
  NOR U54189 ( .A(n41210), .B(n41209), .Z(n48007) );
  IV U54190 ( .A(n41211), .Z(n41217) );
  IV U54191 ( .A(n41212), .Z(n41213) );
  NOR U54192 ( .A(n41217), .B(n41213), .Z(n48004) );
  NOR U54193 ( .A(n41215), .B(n41214), .Z(n44732) );
  NOR U54194 ( .A(n41217), .B(n41216), .Z(n44727) );
  NOR U54195 ( .A(n44732), .B(n44727), .Z(n44493) );
  IV U54196 ( .A(n41218), .Z(n41220) );
  NOR U54197 ( .A(n41220), .B(n41219), .Z(n44735) );
  NOR U54198 ( .A(n44735), .B(n44730), .Z(n44492) );
  IV U54199 ( .A(n41221), .Z(n41223) );
  NOR U54200 ( .A(n41223), .B(n41222), .Z(n44743) );
  IV U54201 ( .A(n41224), .Z(n41225) );
  NOR U54202 ( .A(n41226), .B(n41225), .Z(n44738) );
  NOR U54203 ( .A(n44743), .B(n44738), .Z(n44491) );
  IV U54204 ( .A(n41227), .Z(n41228) );
  NOR U54205 ( .A(n41231), .B(n41228), .Z(n44740) );
  IV U54206 ( .A(n41229), .Z(n41230) );
  NOR U54207 ( .A(n41231), .B(n41230), .Z(n47996) );
  IV U54208 ( .A(n41232), .Z(n41234) );
  IV U54209 ( .A(n41233), .Z(n41236) );
  NOR U54210 ( .A(n41234), .B(n41236), .Z(n47993) );
  IV U54211 ( .A(n41235), .Z(n41237) );
  NOR U54212 ( .A(n41237), .B(n41236), .Z(n44749) );
  IV U54213 ( .A(n41238), .Z(n41239) );
  NOR U54214 ( .A(n41239), .B(n41242), .Z(n44746) );
  IV U54215 ( .A(n41240), .Z(n41241) );
  NOR U54216 ( .A(n41242), .B(n41241), .Z(n44755) );
  IV U54217 ( .A(n41243), .Z(n41248) );
  IV U54218 ( .A(n41244), .Z(n41245) );
  NOR U54219 ( .A(n41248), .B(n41245), .Z(n44752) );
  IV U54220 ( .A(n41246), .Z(n41250) );
  NOR U54221 ( .A(n41248), .B(n41247), .Z(n41249) );
  IV U54222 ( .A(n41249), .Z(n41252) );
  NOR U54223 ( .A(n41250), .B(n41252), .Z(n44761) );
  IV U54224 ( .A(n41251), .Z(n41253) );
  NOR U54225 ( .A(n41253), .B(n41252), .Z(n44758) );
  IV U54226 ( .A(n41254), .Z(n41255) );
  NOR U54227 ( .A(n41255), .B(n41257), .Z(n44767) );
  IV U54228 ( .A(n41256), .Z(n41258) );
  NOR U54229 ( .A(n41258), .B(n41257), .Z(n44764) );
  IV U54230 ( .A(n41259), .Z(n41261) );
  IV U54231 ( .A(n41260), .Z(n44488) );
  NOR U54232 ( .A(n41261), .B(n44488), .Z(n44772) );
  IV U54233 ( .A(n41262), .Z(n41266) );
  NOR U54234 ( .A(n41263), .B(n44479), .Z(n41264) );
  IV U54235 ( .A(n41264), .Z(n41265) );
  NOR U54236 ( .A(n41266), .B(n41265), .Z(n44775) );
  IV U54237 ( .A(n41267), .Z(n41268) );
  NOR U54238 ( .A(n41269), .B(n41268), .Z(n48167) );
  IV U54239 ( .A(n41270), .Z(n41272) );
  NOR U54240 ( .A(n41272), .B(n41271), .Z(n48163) );
  NOR U54241 ( .A(n48167), .B(n48163), .Z(n47980) );
  IV U54242 ( .A(n41273), .Z(n41276) );
  NOR U54243 ( .A(n41274), .B(n44470), .Z(n41275) );
  IV U54244 ( .A(n41275), .Z(n41278) );
  NOR U54245 ( .A(n41276), .B(n41278), .Z(n47977) );
  IV U54246 ( .A(n41277), .Z(n41279) );
  NOR U54247 ( .A(n41279), .B(n41278), .Z(n41280) );
  IV U54248 ( .A(n41280), .Z(n41281) );
  NOR U54249 ( .A(n41282), .B(n41281), .Z(n47973) );
  IV U54250 ( .A(n41283), .Z(n41284) );
  NOR U54251 ( .A(n41284), .B(n41287), .Z(n47964) );
  IV U54252 ( .A(n41285), .Z(n41286) );
  NOR U54253 ( .A(n41287), .B(n41286), .Z(n47960) );
  IV U54254 ( .A(n41288), .Z(n41289) );
  NOR U54255 ( .A(n44448), .B(n41289), .Z(n47943) );
  NOR U54256 ( .A(n41290), .B(n48204), .Z(n47933) );
  IV U54257 ( .A(n41291), .Z(n41292) );
  NOR U54258 ( .A(n41293), .B(n41292), .Z(n44784) );
  NOR U54259 ( .A(n47933), .B(n44784), .Z(n44437) );
  IV U54260 ( .A(n41294), .Z(n41300) );
  IV U54261 ( .A(n41295), .Z(n41296) );
  NOR U54262 ( .A(n41300), .B(n41296), .Z(n41297) );
  IV U54263 ( .A(n41297), .Z(n44791) );
  IV U54264 ( .A(n41298), .Z(n41299) );
  NOR U54265 ( .A(n41300), .B(n41299), .Z(n48209) );
  IV U54266 ( .A(n41301), .Z(n41303) );
  NOR U54267 ( .A(n41303), .B(n41302), .Z(n48213) );
  NOR U54268 ( .A(n48209), .B(n48213), .Z(n47926) );
  IV U54269 ( .A(n41304), .Z(n41305) );
  NOR U54270 ( .A(n44420), .B(n41305), .Z(n44793) );
  IV U54271 ( .A(n41306), .Z(n41311) );
  IV U54272 ( .A(n41307), .Z(n41308) );
  NOR U54273 ( .A(n44420), .B(n41308), .Z(n41309) );
  IV U54274 ( .A(n41309), .Z(n41310) );
  NOR U54275 ( .A(n41311), .B(n41310), .Z(n47920) );
  NOR U54276 ( .A(n44793), .B(n47920), .Z(n44436) );
  IV U54277 ( .A(n41312), .Z(n41314) );
  NOR U54278 ( .A(n41314), .B(n41313), .Z(n44411) );
  IV U54279 ( .A(n41315), .Z(n41316) );
  NOR U54280 ( .A(n41317), .B(n41316), .Z(n44408) );
  IV U54281 ( .A(n44408), .Z(n44403) );
  IV U54282 ( .A(n41318), .Z(n41323) );
  IV U54283 ( .A(n41319), .Z(n41320) );
  NOR U54284 ( .A(n41323), .B(n41320), .Z(n44807) );
  IV U54285 ( .A(n41321), .Z(n41322) );
  NOR U54286 ( .A(n41323), .B(n41322), .Z(n44804) );
  IV U54287 ( .A(n41324), .Z(n41325) );
  NOR U54288 ( .A(n41326), .B(n41325), .Z(n44810) );
  XOR U54289 ( .A(n41328), .B(n41327), .Z(n41331) );
  IV U54290 ( .A(n41329), .Z(n41330) );
  NOR U54291 ( .A(n41331), .B(n41330), .Z(n41332) );
  IV U54292 ( .A(n41332), .Z(n41333) );
  NOR U54293 ( .A(n41334), .B(n41333), .Z(n44814) );
  NOR U54294 ( .A(n44820), .B(n44814), .Z(n44402) );
  NOR U54295 ( .A(n41336), .B(n41335), .Z(n44400) );
  IV U54296 ( .A(n44400), .Z(n44398) );
  IV U54297 ( .A(n41337), .Z(n41338) );
  NOR U54298 ( .A(n41339), .B(n41338), .Z(n41340) );
  IV U54299 ( .A(n41340), .Z(n44824) );
  NOR U54300 ( .A(n41341), .B(n41351), .Z(n41342) );
  IV U54301 ( .A(n41342), .Z(n41344) );
  NOR U54302 ( .A(n41343), .B(n41344), .Z(n47906) );
  NOR U54303 ( .A(n41345), .B(n41344), .Z(n41346) );
  IV U54304 ( .A(n41346), .Z(n41347) );
  NOR U54305 ( .A(n41348), .B(n41347), .Z(n44826) );
  IV U54306 ( .A(n41349), .Z(n41350) );
  NOR U54307 ( .A(n41351), .B(n41350), .Z(n47890) );
  IV U54308 ( .A(n41352), .Z(n41353) );
  NOR U54309 ( .A(n41355), .B(n41353), .Z(n47886) );
  IV U54310 ( .A(n41354), .Z(n41356) );
  NOR U54311 ( .A(n41356), .B(n41355), .Z(n47893) );
  IV U54312 ( .A(n41357), .Z(n41359) );
  NOR U54313 ( .A(n41359), .B(n41358), .Z(n41360) );
  IV U54314 ( .A(n41360), .Z(n44381) );
  IV U54315 ( .A(n41361), .Z(n41363) );
  NOR U54316 ( .A(n41363), .B(n41362), .Z(n41364) );
  IV U54317 ( .A(n41364), .Z(n47871) );
  IV U54318 ( .A(n41365), .Z(n41368) );
  NOR U54319 ( .A(n41371), .B(n41366), .Z(n41367) );
  IV U54320 ( .A(n41367), .Z(n41373) );
  NOR U54321 ( .A(n41368), .B(n41373), .Z(n44841) );
  IV U54322 ( .A(n41369), .Z(n41370) );
  NOR U54323 ( .A(n41371), .B(n41370), .Z(n44852) );
  IV U54324 ( .A(n41372), .Z(n41374) );
  NOR U54325 ( .A(n41374), .B(n41373), .Z(n44847) );
  NOR U54326 ( .A(n44852), .B(n44847), .Z(n44359) );
  IV U54327 ( .A(n41375), .Z(n41377) );
  NOR U54328 ( .A(n41377), .B(n41376), .Z(n44849) );
  IV U54329 ( .A(n41378), .Z(n41379) );
  NOR U54330 ( .A(n41379), .B(n41382), .Z(n44858) );
  IV U54331 ( .A(n41380), .Z(n41381) );
  NOR U54332 ( .A(n41382), .B(n41381), .Z(n44855) );
  IV U54333 ( .A(n41383), .Z(n41384) );
  NOR U54334 ( .A(n41385), .B(n41384), .Z(n51233) );
  IV U54335 ( .A(n41386), .Z(n41387) );
  NOR U54336 ( .A(n44349), .B(n41387), .Z(n48266) );
  NOR U54337 ( .A(n51233), .B(n48266), .Z(n47860) );
  IV U54338 ( .A(n41388), .Z(n41389) );
  NOR U54339 ( .A(n41390), .B(n41389), .Z(n44866) );
  IV U54340 ( .A(n41391), .Z(n41392) );
  NOR U54341 ( .A(n41393), .B(n41392), .Z(n51228) );
  IV U54342 ( .A(n41394), .Z(n41396) );
  IV U54343 ( .A(n41395), .Z(n44344) );
  NOR U54344 ( .A(n41396), .B(n44344), .Z(n51220) );
  NOR U54345 ( .A(n51228), .B(n51220), .Z(n47854) );
  IV U54346 ( .A(n41397), .Z(n41399) );
  NOR U54347 ( .A(n41399), .B(n41398), .Z(n44338) );
  IV U54348 ( .A(n44338), .Z(n44327) );
  NOR U54349 ( .A(n41400), .B(n44872), .Z(n44328) );
  IV U54350 ( .A(n41401), .Z(n41403) );
  NOR U54351 ( .A(n41403), .B(n41402), .Z(n44869) );
  NOR U54352 ( .A(n44328), .B(n44869), .Z(n44325) );
  IV U54353 ( .A(n41404), .Z(n41405) );
  NOR U54354 ( .A(n41406), .B(n41405), .Z(n44876) );
  IV U54355 ( .A(n41410), .Z(n41409) );
  IV U54356 ( .A(n41407), .Z(n41408) );
  NOR U54357 ( .A(n41409), .B(n41408), .Z(n44880) );
  NOR U54358 ( .A(n44876), .B(n44880), .Z(n44323) );
  NOR U54359 ( .A(n41416), .B(n41410), .Z(n41415) );
  IV U54360 ( .A(n41411), .Z(n41412) );
  NOR U54361 ( .A(n41421), .B(n41412), .Z(n41413) );
  IV U54362 ( .A(n41413), .Z(n41414) );
  NOR U54363 ( .A(n41415), .B(n41414), .Z(n51190) );
  IV U54364 ( .A(n41416), .Z(n41418) );
  IV U54365 ( .A(n41417), .Z(n41423) );
  NOR U54366 ( .A(n41418), .B(n41423), .Z(n41419) );
  IV U54367 ( .A(n41419), .Z(n41420) );
  NOR U54368 ( .A(n41421), .B(n41420), .Z(n51185) );
  NOR U54369 ( .A(n51190), .B(n51185), .Z(n44879) );
  IV U54370 ( .A(n41422), .Z(n41424) );
  NOR U54371 ( .A(n41424), .B(n41423), .Z(n44884) );
  NOR U54372 ( .A(n44886), .B(n44884), .Z(n44322) );
  NOR U54373 ( .A(n41426), .B(n41425), .Z(n47835) );
  IV U54374 ( .A(n41427), .Z(n41431) );
  IV U54375 ( .A(n41428), .Z(n41437) );
  NOR U54376 ( .A(n41437), .B(n41429), .Z(n41430) );
  IV U54377 ( .A(n41430), .Z(n41433) );
  NOR U54378 ( .A(n41431), .B(n41433), .Z(n47819) );
  IV U54379 ( .A(n41432), .Z(n41434) );
  NOR U54380 ( .A(n41434), .B(n41433), .Z(n47823) );
  IV U54381 ( .A(n41435), .Z(n41436) );
  NOR U54382 ( .A(n41437), .B(n41436), .Z(n47816) );
  NOR U54383 ( .A(n47823), .B(n47816), .Z(n44312) );
  IV U54384 ( .A(n41438), .Z(n41439) );
  NOR U54385 ( .A(n41439), .B(n41441), .Z(n47813) );
  IV U54386 ( .A(n41440), .Z(n41442) );
  NOR U54387 ( .A(n41442), .B(n41441), .Z(n44891) );
  IV U54388 ( .A(n41443), .Z(n41450) );
  IV U54389 ( .A(n41444), .Z(n41445) );
  NOR U54390 ( .A(n41450), .B(n41445), .Z(n47808) );
  IV U54391 ( .A(n41446), .Z(n41447) );
  NOR U54392 ( .A(n41450), .B(n41447), .Z(n47805) );
  IV U54393 ( .A(n41448), .Z(n41449) );
  NOR U54394 ( .A(n41450), .B(n41449), .Z(n47801) );
  IV U54395 ( .A(n41451), .Z(n41453) );
  NOR U54396 ( .A(n41453), .B(n41452), .Z(n47798) );
  NOR U54397 ( .A(n51153), .B(n51161), .Z(n47786) );
  IV U54398 ( .A(n41454), .Z(n41457) );
  NOR U54399 ( .A(n41455), .B(n44293), .Z(n41456) );
  IV U54400 ( .A(n41456), .Z(n44300) );
  NOR U54401 ( .A(n41457), .B(n44300), .Z(n44895) );
  NOR U54402 ( .A(n41459), .B(n41458), .Z(n44900) );
  IV U54403 ( .A(n41460), .Z(n41465) );
  IV U54404 ( .A(n41461), .Z(n41462) );
  NOR U54405 ( .A(n41465), .B(n41462), .Z(n47758) );
  IV U54406 ( .A(n41463), .Z(n41464) );
  NOR U54407 ( .A(n41465), .B(n41464), .Z(n47755) );
  IV U54408 ( .A(n41466), .Z(n41467) );
  NOR U54409 ( .A(n41468), .B(n41467), .Z(n51142) );
  IV U54410 ( .A(n41469), .Z(n41470) );
  NOR U54411 ( .A(n44270), .B(n41470), .Z(n48337) );
  NOR U54412 ( .A(n51142), .B(n48337), .Z(n47732) );
  NOR U54413 ( .A(n41472), .B(n41471), .Z(n41473) );
  IV U54414 ( .A(n41473), .Z(n41480) );
  XOR U54415 ( .A(n41475), .B(n41474), .Z(n41477) );
  NOR U54416 ( .A(n41477), .B(n41476), .Z(n41478) );
  IV U54417 ( .A(n41478), .Z(n41479) );
  NOR U54418 ( .A(n41480), .B(n41479), .Z(n41481) );
  IV U54419 ( .A(n41481), .Z(n41482) );
  NOR U54420 ( .A(n41483), .B(n41482), .Z(n41484) );
  IV U54421 ( .A(n41484), .Z(n44921) );
  IV U54422 ( .A(n41485), .Z(n41490) );
  IV U54423 ( .A(n41486), .Z(n41487) );
  NOR U54424 ( .A(n41490), .B(n41487), .Z(n44918) );
  IV U54425 ( .A(n41488), .Z(n41489) );
  NOR U54426 ( .A(n41490), .B(n41489), .Z(n47727) );
  IV U54427 ( .A(n41491), .Z(n41492) );
  NOR U54428 ( .A(n44249), .B(n41492), .Z(n41493) );
  IV U54429 ( .A(n41493), .Z(n44244) );
  IV U54430 ( .A(n41494), .Z(n41495) );
  NOR U54431 ( .A(n44236), .B(n41495), .Z(n41496) );
  IV U54432 ( .A(n41496), .Z(n44933) );
  IV U54433 ( .A(n41497), .Z(n41498) );
  NOR U54434 ( .A(n41498), .B(n41504), .Z(n41499) );
  IV U54435 ( .A(n41499), .Z(n47706) );
  IV U54436 ( .A(n41500), .Z(n41501) );
  NOR U54437 ( .A(n41502), .B(n41501), .Z(n47691) );
  IV U54438 ( .A(n41503), .Z(n41505) );
  NOR U54439 ( .A(n41505), .B(n41504), .Z(n47702) );
  NOR U54440 ( .A(n47691), .B(n47702), .Z(n44201) );
  IV U54441 ( .A(n41506), .Z(n41508) );
  NOR U54442 ( .A(n41508), .B(n41507), .Z(n41509) );
  IV U54443 ( .A(n41509), .Z(n47697) );
  IV U54444 ( .A(n41510), .Z(n41511) );
  NOR U54445 ( .A(n41511), .B(n44183), .Z(n41512) );
  IV U54446 ( .A(n41512), .Z(n47683) );
  IV U54447 ( .A(n41513), .Z(n41514) );
  NOR U54448 ( .A(n41514), .B(n41517), .Z(n44954) );
  IV U54449 ( .A(n41515), .Z(n41516) );
  NOR U54450 ( .A(n41517), .B(n41516), .Z(n44951) );
  IV U54451 ( .A(n41518), .Z(n41519) );
  NOR U54452 ( .A(n41520), .B(n41519), .Z(n41521) );
  IV U54453 ( .A(n41521), .Z(n44146) );
  IV U54454 ( .A(n41522), .Z(n41529) );
  IV U54455 ( .A(n41523), .Z(n41524) );
  NOR U54456 ( .A(n41529), .B(n41524), .Z(n41525) );
  IV U54457 ( .A(n41525), .Z(n47670) );
  NOR U54458 ( .A(n41526), .B(n44982), .Z(n44132) );
  IV U54459 ( .A(n41527), .Z(n41528) );
  NOR U54460 ( .A(n41529), .B(n41528), .Z(n47667) );
  IV U54461 ( .A(n41530), .Z(n41532) );
  NOR U54462 ( .A(n41532), .B(n41531), .Z(n44991) );
  IV U54463 ( .A(n41533), .Z(n41534) );
  NOR U54464 ( .A(n41534), .B(n44129), .Z(n44988) );
  IV U54465 ( .A(n41535), .Z(n47661) );
  IV U54466 ( .A(n41536), .Z(n41537) );
  NOR U54467 ( .A(n41543), .B(n41537), .Z(n47650) );
  IV U54468 ( .A(n41538), .Z(n41541) );
  NOR U54469 ( .A(n41539), .B(n41543), .Z(n41540) );
  IV U54470 ( .A(n41540), .Z(n44113) );
  NOR U54471 ( .A(n41541), .B(n44113), .Z(n48407) );
  IV U54472 ( .A(n41542), .Z(n41544) );
  NOR U54473 ( .A(n41544), .B(n41543), .Z(n51029) );
  NOR U54474 ( .A(n48407), .B(n51029), .Z(n47649) );
  IV U54475 ( .A(n41545), .Z(n41546) );
  NOR U54476 ( .A(n41547), .B(n41546), .Z(n45015) );
  IV U54477 ( .A(n41548), .Z(n41551) );
  IV U54478 ( .A(n41549), .Z(n41550) );
  NOR U54479 ( .A(n41551), .B(n41550), .Z(n45023) );
  IV U54480 ( .A(n41552), .Z(n41554) );
  NOR U54481 ( .A(n41554), .B(n41553), .Z(n45038) );
  IV U54482 ( .A(n41555), .Z(n41556) );
  NOR U54483 ( .A(n41557), .B(n41556), .Z(n45049) );
  IV U54484 ( .A(n41558), .Z(n41560) );
  NOR U54485 ( .A(n41560), .B(n41559), .Z(n45043) );
  NOR U54486 ( .A(n45049), .B(n45043), .Z(n44089) );
  IV U54487 ( .A(n41561), .Z(n41562) );
  NOR U54488 ( .A(n41562), .B(n41564), .Z(n45046) );
  IV U54489 ( .A(n41563), .Z(n41565) );
  NOR U54490 ( .A(n41565), .B(n41564), .Z(n45052) );
  NOR U54491 ( .A(n41567), .B(n41566), .Z(n41568) );
  IV U54492 ( .A(n41568), .Z(n41573) );
  NOR U54493 ( .A(n41570), .B(n41569), .Z(n41571) );
  IV U54494 ( .A(n41571), .Z(n41572) );
  NOR U54495 ( .A(n41573), .B(n41572), .Z(n41574) );
  NOR U54496 ( .A(n48438), .B(n41574), .Z(n47625) );
  IV U54497 ( .A(n41575), .Z(n44076) );
  IV U54498 ( .A(n41576), .Z(n41577) );
  NOR U54499 ( .A(n44076), .B(n41577), .Z(n45069) );
  IV U54500 ( .A(n41578), .Z(n41579) );
  NOR U54501 ( .A(n41579), .B(n44071), .Z(n47617) );
  IV U54502 ( .A(n41580), .Z(n41581) );
  NOR U54503 ( .A(n44041), .B(n41581), .Z(n47605) );
  IV U54504 ( .A(n41582), .Z(n41583) );
  NOR U54505 ( .A(n41583), .B(n41587), .Z(n45092) );
  IV U54506 ( .A(n41584), .Z(n47596) );
  NOR U54507 ( .A(n41585), .B(n47596), .Z(n41589) );
  IV U54508 ( .A(n41586), .Z(n41588) );
  NOR U54509 ( .A(n41588), .B(n41587), .Z(n45095) );
  NOR U54510 ( .A(n41589), .B(n45095), .Z(n44038) );
  IV U54511 ( .A(n41590), .Z(n41591) );
  NOR U54512 ( .A(n41591), .B(n44037), .Z(n47591) );
  IV U54513 ( .A(n41592), .Z(n41594) );
  NOR U54514 ( .A(n41594), .B(n41593), .Z(n45100) );
  NOR U54515 ( .A(n41596), .B(n41595), .Z(n47585) );
  IV U54516 ( .A(n41597), .Z(n41599) );
  NOR U54517 ( .A(n41599), .B(n41598), .Z(n47579) );
  NOR U54518 ( .A(n47579), .B(n47582), .Z(n44026) );
  NOR U54519 ( .A(n41601), .B(n41600), .Z(n44024) );
  IV U54520 ( .A(n44024), .Z(n44017) );
  NOR U54521 ( .A(n47563), .B(n47561), .Z(n41602) );
  IV U54522 ( .A(n41602), .Z(n47564) );
  IV U54523 ( .A(n41603), .Z(n41604) );
  NOR U54524 ( .A(n41605), .B(n41604), .Z(n50894) );
  IV U54525 ( .A(n41606), .Z(n41611) );
  IV U54526 ( .A(n41607), .Z(n41608) );
  NOR U54527 ( .A(n41611), .B(n41608), .Z(n48482) );
  NOR U54528 ( .A(n50894), .B(n48482), .Z(n47536) );
  IV U54529 ( .A(n41609), .Z(n41613) );
  NOR U54530 ( .A(n41611), .B(n41610), .Z(n41612) );
  IV U54531 ( .A(n41612), .Z(n41615) );
  NOR U54532 ( .A(n41613), .B(n41615), .Z(n45115) );
  IV U54533 ( .A(n41614), .Z(n41616) );
  NOR U54534 ( .A(n41616), .B(n41615), .Z(n45112) );
  IV U54535 ( .A(n41617), .Z(n41619) );
  NOR U54536 ( .A(n41619), .B(n41618), .Z(n45121) );
  IV U54537 ( .A(n41620), .Z(n41621) );
  NOR U54538 ( .A(n41621), .B(n41623), .Z(n45118) );
  IV U54539 ( .A(n41622), .Z(n41624) );
  NOR U54540 ( .A(n41624), .B(n41623), .Z(n45127) );
  IV U54541 ( .A(n41625), .Z(n41634) );
  NOR U54542 ( .A(n43994), .B(n41626), .Z(n41627) );
  IV U54543 ( .A(n41627), .Z(n41632) );
  NOR U54544 ( .A(n41629), .B(n41628), .Z(n41630) );
  IV U54545 ( .A(n41630), .Z(n41631) );
  NOR U54546 ( .A(n41632), .B(n41631), .Z(n41633) );
  IV U54547 ( .A(n41633), .Z(n41636) );
  NOR U54548 ( .A(n41634), .B(n41636), .Z(n45124) );
  IV U54549 ( .A(n41635), .Z(n41637) );
  NOR U54550 ( .A(n41637), .B(n41636), .Z(n45130) );
  NOR U54551 ( .A(n41638), .B(n43983), .Z(n41639) );
  IV U54552 ( .A(n41639), .Z(n41640) );
  NOR U54553 ( .A(n41641), .B(n41640), .Z(n47525) );
  IV U54554 ( .A(n41642), .Z(n41643) );
  NOR U54555 ( .A(n41644), .B(n41643), .Z(n47508) );
  IV U54556 ( .A(n41645), .Z(n41646) );
  NOR U54557 ( .A(n41646), .B(n43976), .Z(n47514) );
  NOR U54558 ( .A(n47508), .B(n47514), .Z(n43974) );
  IV U54559 ( .A(n41647), .Z(n41650) );
  IV U54560 ( .A(n41648), .Z(n41649) );
  NOR U54561 ( .A(n41650), .B(n41649), .Z(n47504) );
  IV U54562 ( .A(n41651), .Z(n41652) );
  NOR U54563 ( .A(n41652), .B(n41653), .Z(n47501) );
  NOR U54564 ( .A(n41654), .B(n41653), .Z(n47498) );
  IV U54565 ( .A(n41655), .Z(n41656) );
  NOR U54566 ( .A(n43964), .B(n41656), .Z(n47489) );
  IV U54567 ( .A(n41657), .Z(n41658) );
  NOR U54568 ( .A(n41659), .B(n41658), .Z(n45149) );
  NOR U54569 ( .A(n41661), .B(n41660), .Z(n47479) );
  NOR U54570 ( .A(n41662), .B(n41666), .Z(n45152) );
  IV U54571 ( .A(n41663), .Z(n41664) );
  NOR U54572 ( .A(n41665), .B(n41664), .Z(n47466) );
  NOR U54573 ( .A(n41667), .B(n41666), .Z(n47470) );
  NOR U54574 ( .A(n47466), .B(n47470), .Z(n45155) );
  IV U54575 ( .A(n41668), .Z(n41669) );
  NOR U54576 ( .A(n41670), .B(n41669), .Z(n45157) );
  IV U54577 ( .A(n41671), .Z(n41672) );
  NOR U54578 ( .A(n41672), .B(n41677), .Z(n45159) );
  NOR U54579 ( .A(n45157), .B(n45159), .Z(n43956) );
  IV U54580 ( .A(n41673), .Z(n41674) );
  NOR U54581 ( .A(n41675), .B(n41674), .Z(n47459) );
  IV U54582 ( .A(n41676), .Z(n41678) );
  NOR U54583 ( .A(n41678), .B(n41677), .Z(n45162) );
  NOR U54584 ( .A(n47459), .B(n45162), .Z(n43955) );
  IV U54585 ( .A(n41679), .Z(n41684) );
  IV U54586 ( .A(n41680), .Z(n41681) );
  NOR U54587 ( .A(n41684), .B(n41681), .Z(n47456) );
  IV U54588 ( .A(n41682), .Z(n41683) );
  NOR U54589 ( .A(n41684), .B(n41683), .Z(n47452) );
  IV U54590 ( .A(n41685), .Z(n41686) );
  NOR U54591 ( .A(n41689), .B(n41686), .Z(n47449) );
  IV U54592 ( .A(n41687), .Z(n41688) );
  NOR U54593 ( .A(n41689), .B(n41688), .Z(n47445) );
  NOR U54594 ( .A(n41691), .B(n41690), .Z(n45164) );
  IV U54595 ( .A(n41692), .Z(n41695) );
  IV U54596 ( .A(n41693), .Z(n41694) );
  NOR U54597 ( .A(n41695), .B(n41694), .Z(n41696) );
  IV U54598 ( .A(n41696), .Z(n47435) );
  IV U54599 ( .A(n41697), .Z(n41706) );
  IV U54600 ( .A(n41711), .Z(n41699) );
  NOR U54601 ( .A(n41699), .B(n41698), .Z(n41704) );
  XOR U54602 ( .A(n41717), .B(n41718), .Z(n41700) );
  NOR U54603 ( .A(n41701), .B(n41700), .Z(n41702) );
  IV U54604 ( .A(n41702), .Z(n41703) );
  NOR U54605 ( .A(n41704), .B(n41703), .Z(n41705) );
  IV U54606 ( .A(n41705), .Z(n41708) );
  NOR U54607 ( .A(n41706), .B(n41708), .Z(n45172) );
  IV U54608 ( .A(n41707), .Z(n41709) );
  NOR U54609 ( .A(n41709), .B(n41708), .Z(n47418) );
  IV U54610 ( .A(n41710), .Z(n41713) );
  NOR U54611 ( .A(n41711), .B(n41718), .Z(n41712) );
  IV U54612 ( .A(n41712), .Z(n41715) );
  NOR U54613 ( .A(n41713), .B(n41715), .Z(n47422) );
  IV U54614 ( .A(n41714), .Z(n41716) );
  NOR U54615 ( .A(n41716), .B(n41715), .Z(n45175) );
  IV U54616 ( .A(n41717), .Z(n41719) );
  NOR U54617 ( .A(n41719), .B(n41718), .Z(n43933) );
  IV U54618 ( .A(n43933), .Z(n43925) );
  IV U54619 ( .A(n41720), .Z(n41721) );
  NOR U54620 ( .A(n41721), .B(n43918), .Z(n47392) );
  IV U54621 ( .A(n41722), .Z(n41724) );
  NOR U54622 ( .A(n41724), .B(n41723), .Z(n47395) );
  NOR U54623 ( .A(n47387), .B(n47395), .Z(n43916) );
  IV U54624 ( .A(n41725), .Z(n41726) );
  NOR U54625 ( .A(n47377), .B(n41726), .Z(n50825) );
  IV U54626 ( .A(n41727), .Z(n41728) );
  NOR U54627 ( .A(n41729), .B(n41728), .Z(n45187) );
  IV U54628 ( .A(n41730), .Z(n41731) );
  NOR U54629 ( .A(n41731), .B(n47377), .Z(n48599) );
  NOR U54630 ( .A(n45187), .B(n48599), .Z(n43903) );
  IV U54631 ( .A(n41732), .Z(n41733) );
  NOR U54632 ( .A(n41733), .B(n43897), .Z(n41734) );
  IV U54633 ( .A(n41734), .Z(n47368) );
  IV U54634 ( .A(n41735), .Z(n41740) );
  IV U54635 ( .A(n41736), .Z(n41737) );
  NOR U54636 ( .A(n41740), .B(n41737), .Z(n45190) );
  IV U54637 ( .A(n41738), .Z(n41739) );
  NOR U54638 ( .A(n41740), .B(n41739), .Z(n47333) );
  IV U54639 ( .A(n41741), .Z(n41743) );
  IV U54640 ( .A(n41742), .Z(n41746) );
  NOR U54641 ( .A(n41743), .B(n41746), .Z(n47337) );
  IV U54642 ( .A(n41744), .Z(n41745) );
  NOR U54643 ( .A(n41745), .B(n41749), .Z(n48622) );
  NOR U54644 ( .A(n41747), .B(n41746), .Z(n50805) );
  NOR U54645 ( .A(n48622), .B(n50805), .Z(n45195) );
  IV U54646 ( .A(n41748), .Z(n41750) );
  NOR U54647 ( .A(n41750), .B(n41749), .Z(n47324) );
  IV U54648 ( .A(n41751), .Z(n41756) );
  IV U54649 ( .A(n41752), .Z(n41753) );
  NOR U54650 ( .A(n41756), .B(n41753), .Z(n47321) );
  IV U54651 ( .A(n41754), .Z(n41755) );
  NOR U54652 ( .A(n41756), .B(n41755), .Z(n47317) );
  IV U54653 ( .A(n41757), .Z(n41759) );
  NOR U54654 ( .A(n41759), .B(n41758), .Z(n47314) );
  IV U54655 ( .A(n41760), .Z(n41763) );
  NOR U54656 ( .A(n41761), .B(n43869), .Z(n41762) );
  IV U54657 ( .A(n41762), .Z(n43875) );
  NOR U54658 ( .A(n41763), .B(n43875), .Z(n47310) );
  IV U54659 ( .A(n41764), .Z(n41765) );
  NOR U54660 ( .A(n41765), .B(n41770), .Z(n47295) );
  IV U54661 ( .A(n41766), .Z(n41767) );
  NOR U54662 ( .A(n41768), .B(n41767), .Z(n45204) );
  IV U54663 ( .A(n41769), .Z(n41771) );
  NOR U54664 ( .A(n41771), .B(n41770), .Z(n47298) );
  NOR U54665 ( .A(n45204), .B(n47298), .Z(n43866) );
  NOR U54666 ( .A(n41773), .B(n41772), .Z(n45207) );
  IV U54667 ( .A(n41774), .Z(n41777) );
  NOR U54668 ( .A(n41775), .B(n41782), .Z(n41776) );
  IV U54669 ( .A(n41776), .Z(n43856) );
  NOR U54670 ( .A(n41777), .B(n43856), .Z(n48664) );
  NOR U54671 ( .A(n48657), .B(n48664), .Z(n45214) );
  IV U54672 ( .A(n41778), .Z(n41780) );
  NOR U54673 ( .A(n41780), .B(n41779), .Z(n48672) );
  IV U54674 ( .A(n41781), .Z(n41783) );
  NOR U54675 ( .A(n41783), .B(n41782), .Z(n50785) );
  NOR U54676 ( .A(n48672), .B(n50785), .Z(n45218) );
  IV U54677 ( .A(n41784), .Z(n43850) );
  IV U54678 ( .A(n41785), .Z(n41786) );
  NOR U54679 ( .A(n43850), .B(n41786), .Z(n47285) );
  IV U54680 ( .A(n41787), .Z(n41789) );
  NOR U54681 ( .A(n41789), .B(n41788), .Z(n45222) );
  IV U54682 ( .A(n41790), .Z(n41791) );
  NOR U54683 ( .A(n43843), .B(n41791), .Z(n43839) );
  IV U54684 ( .A(n43839), .Z(n43831) );
  IV U54685 ( .A(n41792), .Z(n41794) );
  NOR U54686 ( .A(n41794), .B(n41793), .Z(n47264) );
  IV U54687 ( .A(n41795), .Z(n41797) );
  IV U54688 ( .A(n41796), .Z(n43828) );
  NOR U54689 ( .A(n41797), .B(n43828), .Z(n45228) );
  IV U54690 ( .A(n41798), .Z(n41800) );
  NOR U54691 ( .A(n41800), .B(n41799), .Z(n48694) );
  NOR U54692 ( .A(n48694), .B(n50775), .Z(n45237) );
  IV U54693 ( .A(n41801), .Z(n41806) );
  IV U54694 ( .A(n41802), .Z(n41803) );
  NOR U54695 ( .A(n41806), .B(n41803), .Z(n45234) );
  IV U54696 ( .A(n41804), .Z(n41805) );
  NOR U54697 ( .A(n41806), .B(n41805), .Z(n45240) );
  IV U54698 ( .A(n41807), .Z(n41808) );
  NOR U54699 ( .A(n41808), .B(n41810), .Z(n47251) );
  NOR U54700 ( .A(n45240), .B(n47251), .Z(n43824) );
  IV U54701 ( .A(n41809), .Z(n41811) );
  NOR U54702 ( .A(n41811), .B(n41810), .Z(n47237) );
  NOR U54703 ( .A(n41812), .B(n47237), .Z(n43823) );
  IV U54704 ( .A(n41813), .Z(n41814) );
  NOR U54705 ( .A(n43821), .B(n41814), .Z(n47228) );
  IV U54706 ( .A(n41815), .Z(n41817) );
  NOR U54707 ( .A(n41817), .B(n41816), .Z(n47215) );
  IV U54708 ( .A(n41818), .Z(n41822) );
  IV U54709 ( .A(n41819), .Z(n43787) );
  NOR U54710 ( .A(n43787), .B(n41820), .Z(n41821) );
  IV U54711 ( .A(n41821), .Z(n43793) );
  NOR U54712 ( .A(n41822), .B(n43793), .Z(n47207) );
  NOR U54713 ( .A(n47215), .B(n47207), .Z(n43800) );
  IV U54714 ( .A(n41823), .Z(n41827) );
  IV U54715 ( .A(n41824), .Z(n43778) );
  NOR U54716 ( .A(n43778), .B(n41825), .Z(n41826) );
  IV U54717 ( .A(n41826), .Z(n43780) );
  NOR U54718 ( .A(n41827), .B(n43780), .Z(n41828) );
  IV U54719 ( .A(n41828), .Z(n47200) );
  IV U54720 ( .A(n41829), .Z(n41836) );
  IV U54721 ( .A(n41830), .Z(n41831) );
  NOR U54722 ( .A(n41836), .B(n41831), .Z(n45270) );
  IV U54723 ( .A(n41832), .Z(n41833) );
  NOR U54724 ( .A(n43773), .B(n41833), .Z(n45268) );
  NOR U54725 ( .A(n45270), .B(n45268), .Z(n43771) );
  IV U54726 ( .A(n41834), .Z(n41835) );
  NOR U54727 ( .A(n41836), .B(n41835), .Z(n47182) );
  IV U54728 ( .A(n41837), .Z(n41838) );
  NOR U54729 ( .A(n41838), .B(n41844), .Z(n41839) );
  IV U54730 ( .A(n41839), .Z(n47177) );
  IV U54731 ( .A(n41840), .Z(n41841) );
  NOR U54732 ( .A(n41842), .B(n41841), .Z(n54218) );
  IV U54733 ( .A(n41843), .Z(n41845) );
  NOR U54734 ( .A(n41845), .B(n41844), .Z(n54227) );
  NOR U54735 ( .A(n54218), .B(n54227), .Z(n47175) );
  IV U54736 ( .A(n41846), .Z(n41853) );
  IV U54737 ( .A(n41847), .Z(n41860) );
  XOR U54738 ( .A(n41860), .B(n41848), .Z(n41849) );
  NOR U54739 ( .A(n41850), .B(n41849), .Z(n41851) );
  IV U54740 ( .A(n41851), .Z(n41852) );
  NOR U54741 ( .A(n41853), .B(n41852), .Z(n47163) );
  IV U54742 ( .A(n41854), .Z(n41855) );
  NOR U54743 ( .A(n41855), .B(n41859), .Z(n47159) );
  IV U54744 ( .A(n41856), .Z(n41857) );
  NOR U54745 ( .A(n41858), .B(n41857), .Z(n52381) );
  NOR U54746 ( .A(n41860), .B(n41859), .Z(n52372) );
  NOR U54747 ( .A(n52381), .B(n52372), .Z(n47158) );
  XOR U54748 ( .A(n41861), .B(n41867), .Z(n41862) );
  NOR U54749 ( .A(n41868), .B(n41862), .Z(n41863) );
  IV U54750 ( .A(n41863), .Z(n41864) );
  NOR U54751 ( .A(n41865), .B(n41864), .Z(n47153) );
  IV U54752 ( .A(n41866), .Z(n41870) );
  NOR U54753 ( .A(n41868), .B(n41867), .Z(n41869) );
  IV U54754 ( .A(n41869), .Z(n43759) );
  NOR U54755 ( .A(n41870), .B(n43759), .Z(n47150) );
  IV U54756 ( .A(n41871), .Z(n41875) );
  NOR U54757 ( .A(n41873), .B(n41872), .Z(n41874) );
  IV U54758 ( .A(n41874), .Z(n41877) );
  NOR U54759 ( .A(n41875), .B(n41877), .Z(n47145) );
  IV U54760 ( .A(n41876), .Z(n41878) );
  NOR U54761 ( .A(n41878), .B(n41877), .Z(n47142) );
  IV U54762 ( .A(n41879), .Z(n41880) );
  NOR U54763 ( .A(n41883), .B(n41880), .Z(n45289) );
  IV U54764 ( .A(n41881), .Z(n41882) );
  NOR U54765 ( .A(n41883), .B(n41882), .Z(n45295) );
  NOR U54766 ( .A(n45295), .B(n45287), .Z(n43741) );
  IV U54767 ( .A(n41884), .Z(n41886) );
  NOR U54768 ( .A(n41886), .B(n41885), .Z(n45292) );
  IV U54769 ( .A(n41887), .Z(n41888) );
  NOR U54770 ( .A(n41888), .B(n43738), .Z(n45300) );
  IV U54771 ( .A(n41889), .Z(n41890) );
  NOR U54772 ( .A(n41893), .B(n41890), .Z(n45303) );
  IV U54773 ( .A(n41891), .Z(n41892) );
  NOR U54774 ( .A(n41893), .B(n41892), .Z(n47128) );
  IV U54775 ( .A(n41894), .Z(n41896) );
  IV U54776 ( .A(n41895), .Z(n41898) );
  NOR U54777 ( .A(n41896), .B(n41898), .Z(n47120) );
  NOR U54778 ( .A(n47128), .B(n47120), .Z(n43731) );
  IV U54779 ( .A(n41897), .Z(n41899) );
  NOR U54780 ( .A(n41899), .B(n41898), .Z(n41900) );
  IV U54781 ( .A(n41900), .Z(n41901) );
  NOR U54782 ( .A(n43723), .B(n41901), .Z(n41902) );
  IV U54783 ( .A(n41902), .Z(n45311) );
  IV U54784 ( .A(n41903), .Z(n41905) );
  NOR U54785 ( .A(n41905), .B(n41904), .Z(n47112) );
  IV U54786 ( .A(n41906), .Z(n41908) );
  IV U54787 ( .A(n41907), .Z(n43710) );
  NOR U54788 ( .A(n41908), .B(n43710), .Z(n47109) );
  IV U54789 ( .A(n41909), .Z(n41913) );
  NOR U54790 ( .A(n41911), .B(n41910), .Z(n41912) );
  IV U54791 ( .A(n41912), .Z(n43704) );
  NOR U54792 ( .A(n41913), .B(n43704), .Z(n45333) );
  IV U54793 ( .A(n41914), .Z(n41915) );
  NOR U54794 ( .A(n41915), .B(n41917), .Z(n47093) );
  IV U54795 ( .A(n41916), .Z(n41918) );
  NOR U54796 ( .A(n41918), .B(n41917), .Z(n47090) );
  IV U54797 ( .A(n41919), .Z(n41924) );
  IV U54798 ( .A(n41920), .Z(n41921) );
  NOR U54799 ( .A(n41924), .B(n41921), .Z(n45339) );
  IV U54800 ( .A(n41922), .Z(n41923) );
  NOR U54801 ( .A(n41924), .B(n41923), .Z(n45342) );
  IV U54802 ( .A(n41925), .Z(n41926) );
  NOR U54803 ( .A(n41927), .B(n41926), .Z(n47086) );
  NOR U54804 ( .A(n45342), .B(n47086), .Z(n43701) );
  IV U54805 ( .A(n41928), .Z(n41931) );
  NOR U54806 ( .A(n41929), .B(n43692), .Z(n41930) );
  IV U54807 ( .A(n41930), .Z(n43699) );
  NOR U54808 ( .A(n41931), .B(n43699), .Z(n47082) );
  IV U54809 ( .A(n41932), .Z(n41933) );
  NOR U54810 ( .A(n41934), .B(n41933), .Z(n45357) );
  IV U54811 ( .A(n41935), .Z(n41936) );
  NOR U54812 ( .A(n41936), .B(n43688), .Z(n45349) );
  NOR U54813 ( .A(n45357), .B(n45349), .Z(n43685) );
  IV U54814 ( .A(n41937), .Z(n41938) );
  NOR U54815 ( .A(n41940), .B(n41938), .Z(n45354) );
  IV U54816 ( .A(n41939), .Z(n41941) );
  NOR U54817 ( .A(n41941), .B(n41940), .Z(n45360) );
  IV U54818 ( .A(n41942), .Z(n41949) );
  NOR U54819 ( .A(n41944), .B(n41943), .Z(n41945) );
  IV U54820 ( .A(n41945), .Z(n41951) );
  XOR U54821 ( .A(n41950), .B(n41955), .Z(n41946) );
  NOR U54822 ( .A(n41951), .B(n41946), .Z(n41947) );
  IV U54823 ( .A(n41947), .Z(n41948) );
  NOR U54824 ( .A(n41949), .B(n41948), .Z(n47068) );
  IV U54825 ( .A(n41950), .Z(n41952) );
  NOR U54826 ( .A(n41952), .B(n41951), .Z(n41953) );
  IV U54827 ( .A(n41953), .Z(n41954) );
  NOR U54828 ( .A(n41955), .B(n41954), .Z(n43674) );
  IV U54829 ( .A(n43674), .Z(n43662) );
  IV U54830 ( .A(n41956), .Z(n41957) );
  NOR U54831 ( .A(n41963), .B(n41957), .Z(n52486) );
  IV U54832 ( .A(n41958), .Z(n41960) );
  IV U54833 ( .A(n41959), .Z(n43658) );
  NOR U54834 ( .A(n41960), .B(n43658), .Z(n52481) );
  NOR U54835 ( .A(n52486), .B(n52481), .Z(n45370) );
  IV U54836 ( .A(n41961), .Z(n41962) );
  NOR U54837 ( .A(n41963), .B(n41962), .Z(n45374) );
  IV U54838 ( .A(n41964), .Z(n41966) );
  IV U54839 ( .A(n41965), .Z(n41968) );
  NOR U54840 ( .A(n41966), .B(n41968), .Z(n45371) );
  IV U54841 ( .A(n41967), .Z(n41969) );
  NOR U54842 ( .A(n41969), .B(n41968), .Z(n45380) );
  IV U54843 ( .A(n41970), .Z(n41971) );
  NOR U54844 ( .A(n43652), .B(n41971), .Z(n45377) );
  IV U54845 ( .A(n41972), .Z(n41974) );
  IV U54846 ( .A(n41973), .Z(n43648) );
  NOR U54847 ( .A(n41974), .B(n43648), .Z(n47059) );
  IV U54848 ( .A(n41975), .Z(n41976) );
  NOR U54849 ( .A(n41976), .B(n41979), .Z(n45386) );
  NOR U54850 ( .A(n41977), .B(n45386), .Z(n43645) );
  IV U54851 ( .A(n41978), .Z(n41980) );
  NOR U54852 ( .A(n41980), .B(n41979), .Z(n47054) );
  IV U54853 ( .A(n41981), .Z(n41982) );
  NOR U54854 ( .A(n43639), .B(n41982), .Z(n41983) );
  IV U54855 ( .A(n41983), .Z(n47052) );
  IV U54856 ( .A(n41984), .Z(n41986) );
  NOR U54857 ( .A(n41986), .B(n41985), .Z(n47039) );
  IV U54858 ( .A(n41987), .Z(n41988) );
  NOR U54859 ( .A(n41989), .B(n41988), .Z(n45400) );
  IV U54860 ( .A(n41990), .Z(n41992) );
  NOR U54861 ( .A(n41992), .B(n41991), .Z(n47036) );
  NOR U54862 ( .A(n45400), .B(n47036), .Z(n43622) );
  IV U54863 ( .A(n41993), .Z(n41994) );
  NOR U54864 ( .A(n41997), .B(n41994), .Z(n45405) );
  IV U54865 ( .A(n41995), .Z(n41996) );
  NOR U54866 ( .A(n41997), .B(n41996), .Z(n45402) );
  NOR U54867 ( .A(n41999), .B(n41998), .Z(n45410) );
  NOR U54868 ( .A(n42000), .B(n45417), .Z(n42003) );
  NOR U54869 ( .A(n42002), .B(n42001), .Z(n45413) );
  NOR U54870 ( .A(n42003), .B(n45413), .Z(n43610) );
  IV U54871 ( .A(n42004), .Z(n43609) );
  IV U54872 ( .A(n42005), .Z(n42006) );
  NOR U54873 ( .A(n43609), .B(n42006), .Z(n47023) );
  IV U54874 ( .A(n42007), .Z(n42008) );
  NOR U54875 ( .A(n42009), .B(n42008), .Z(n50450) );
  IV U54876 ( .A(n42010), .Z(n42011) );
  NOR U54877 ( .A(n42011), .B(n43604), .Z(n48855) );
  NOR U54878 ( .A(n50450), .B(n48855), .Z(n46998) );
  IV U54879 ( .A(n42012), .Z(n42013) );
  NOR U54880 ( .A(n42013), .B(n42015), .Z(n46990) );
  IV U54881 ( .A(n42014), .Z(n42016) );
  NOR U54882 ( .A(n42016), .B(n42015), .Z(n45423) );
  NOR U54883 ( .A(n46990), .B(n45423), .Z(n43597) );
  IV U54884 ( .A(n42017), .Z(n42019) );
  NOR U54885 ( .A(n42019), .B(n42018), .Z(n42020) );
  IV U54886 ( .A(n42020), .Z(n46989) );
  IV U54887 ( .A(n42021), .Z(n42023) );
  NOR U54888 ( .A(n42023), .B(n42022), .Z(n42024) );
  IV U54889 ( .A(n42024), .Z(n43590) );
  XOR U54890 ( .A(n42026), .B(n42025), .Z(n42030) );
  NOR U54891 ( .A(n42027), .B(n42032), .Z(n42028) );
  IV U54892 ( .A(n42028), .Z(n42029) );
  NOR U54893 ( .A(n42030), .B(n42029), .Z(n46983) );
  IV U54894 ( .A(n42031), .Z(n42033) );
  NOR U54895 ( .A(n42033), .B(n42032), .Z(n45428) );
  IV U54896 ( .A(n42034), .Z(n42038) );
  IV U54897 ( .A(n42035), .Z(n43579) );
  NOR U54898 ( .A(n42036), .B(n43579), .Z(n42037) );
  IV U54899 ( .A(n42037), .Z(n42040) );
  NOR U54900 ( .A(n42038), .B(n42040), .Z(n46973) );
  IV U54901 ( .A(n42039), .Z(n42043) );
  NOR U54902 ( .A(n42041), .B(n42040), .Z(n42042) );
  IV U54903 ( .A(n42042), .Z(n43581) );
  NOR U54904 ( .A(n42043), .B(n43581), .Z(n45431) );
  NOR U54905 ( .A(n42045), .B(n42044), .Z(n45435) );
  IV U54906 ( .A(n42046), .Z(n42047) );
  NOR U54907 ( .A(n42048), .B(n42047), .Z(n42049) );
  IV U54908 ( .A(n42049), .Z(n43555) );
  IV U54909 ( .A(n42050), .Z(n42052) );
  NOR U54910 ( .A(n42052), .B(n42051), .Z(n42053) );
  IV U54911 ( .A(n42053), .Z(n43543) );
  IV U54912 ( .A(n42054), .Z(n42060) );
  IV U54913 ( .A(n42055), .Z(n42056) );
  NOR U54914 ( .A(n42060), .B(n42056), .Z(n42057) );
  IV U54915 ( .A(n42057), .Z(n46936) );
  IV U54916 ( .A(n42058), .Z(n42059) );
  NOR U54917 ( .A(n42060), .B(n42059), .Z(n46932) );
  IV U54918 ( .A(n42061), .Z(n42063) );
  NOR U54919 ( .A(n42063), .B(n42062), .Z(n46929) );
  IV U54920 ( .A(n42064), .Z(n42065) );
  NOR U54921 ( .A(n42065), .B(n43524), .Z(n45446) );
  IV U54922 ( .A(n42066), .Z(n42068) );
  NOR U54923 ( .A(n42068), .B(n42067), .Z(n45455) );
  IV U54924 ( .A(n42069), .Z(n42071) );
  NOR U54925 ( .A(n42071), .B(n42070), .Z(n45451) );
  NOR U54926 ( .A(n45455), .B(n45451), .Z(n43518) );
  IV U54927 ( .A(n42072), .Z(n42073) );
  NOR U54928 ( .A(n42074), .B(n42073), .Z(n46908) );
  IV U54929 ( .A(n42075), .Z(n42076) );
  NOR U54930 ( .A(n42076), .B(n43517), .Z(n45459) );
  NOR U54931 ( .A(n46908), .B(n45459), .Z(n43511) );
  IV U54932 ( .A(n42077), .Z(n42079) );
  NOR U54933 ( .A(n42079), .B(n42078), .Z(n45462) );
  IV U54934 ( .A(n42080), .Z(n42081) );
  NOR U54935 ( .A(n42081), .B(n43492), .Z(n42082) );
  IV U54936 ( .A(n42082), .Z(n43505) );
  NOR U54937 ( .A(n42083), .B(n45471), .Z(n43490) );
  IV U54938 ( .A(n42084), .Z(n42086) );
  NOR U54939 ( .A(n42086), .B(n42085), .Z(n45474) );
  IV U54940 ( .A(n42087), .Z(n42089) );
  NOR U54941 ( .A(n42089), .B(n42088), .Z(n45467) );
  NOR U54942 ( .A(n45474), .B(n45467), .Z(n43489) );
  IV U54943 ( .A(n42090), .Z(n42091) );
  NOR U54944 ( .A(n42092), .B(n42091), .Z(n45480) );
  IV U54945 ( .A(n42093), .Z(n42095) );
  NOR U54946 ( .A(n42095), .B(n42094), .Z(n45477) );
  NOR U54947 ( .A(n45480), .B(n45477), .Z(n43488) );
  IV U54948 ( .A(n42096), .Z(n42097) );
  NOR U54949 ( .A(n42097), .B(n42103), .Z(n42098) );
  IV U54950 ( .A(n42098), .Z(n45484) );
  IV U54951 ( .A(n42099), .Z(n42100) );
  NOR U54952 ( .A(n42101), .B(n42100), .Z(n50313) );
  IV U54953 ( .A(n42102), .Z(n42104) );
  NOR U54954 ( .A(n42104), .B(n42103), .Z(n50318) );
  NOR U54955 ( .A(n50313), .B(n50318), .Z(n45483) );
  IV U54956 ( .A(n42105), .Z(n42106) );
  NOR U54957 ( .A(n42111), .B(n42106), .Z(n46893) );
  IV U54958 ( .A(n42107), .Z(n42109) );
  NOR U54959 ( .A(n42109), .B(n42108), .Z(n46887) );
  IV U54960 ( .A(n42110), .Z(n42112) );
  NOR U54961 ( .A(n42112), .B(n42111), .Z(n46890) );
  NOR U54962 ( .A(n46887), .B(n46890), .Z(n43486) );
  IV U54963 ( .A(n42113), .Z(n42114) );
  NOR U54964 ( .A(n42116), .B(n42114), .Z(n46884) );
  NOR U54965 ( .A(n42116), .B(n42115), .Z(n42117) );
  IV U54966 ( .A(n42117), .Z(n42118) );
  NOR U54967 ( .A(n42119), .B(n42118), .Z(n45490) );
  IV U54968 ( .A(n42120), .Z(n42123) );
  IV U54969 ( .A(n42121), .Z(n42122) );
  NOR U54970 ( .A(n42123), .B(n42122), .Z(n45487) );
  IV U54971 ( .A(n42124), .Z(n42126) );
  XOR U54972 ( .A(n42129), .B(n42130), .Z(n42125) );
  NOR U54973 ( .A(n42126), .B(n42125), .Z(n45496) );
  IV U54974 ( .A(n42127), .Z(n42128) );
  NOR U54975 ( .A(n42128), .B(n42130), .Z(n45493) );
  IV U54976 ( .A(n42129), .Z(n42131) );
  NOR U54977 ( .A(n42131), .B(n42130), .Z(n45502) );
  IV U54978 ( .A(n42132), .Z(n42134) );
  IV U54979 ( .A(n42133), .Z(n42136) );
  NOR U54980 ( .A(n42134), .B(n42136), .Z(n45499) );
  IV U54981 ( .A(n42135), .Z(n42137) );
  NOR U54982 ( .A(n42137), .B(n42136), .Z(n42138) );
  IV U54983 ( .A(n42138), .Z(n43482) );
  NOR U54984 ( .A(n42140), .B(n42139), .Z(n45505) );
  NOR U54985 ( .A(n46869), .B(n45505), .Z(n43475) );
  IV U54986 ( .A(n42141), .Z(n42142) );
  NOR U54987 ( .A(n42142), .B(n43469), .Z(n45507) );
  NOR U54988 ( .A(n42143), .B(n43469), .Z(n42144) );
  IV U54989 ( .A(n42144), .Z(n42145) );
  NOR U54990 ( .A(n43468), .B(n42145), .Z(n46873) );
  IV U54991 ( .A(n42146), .Z(n42147) );
  NOR U54992 ( .A(n42147), .B(n43466), .Z(n43463) );
  IV U54993 ( .A(n43463), .Z(n43454) );
  IV U54994 ( .A(n42148), .Z(n42149) );
  NOR U54995 ( .A(n42153), .B(n42149), .Z(n42150) );
  IV U54996 ( .A(n42150), .Z(n46854) );
  IV U54997 ( .A(n42151), .Z(n42152) );
  NOR U54998 ( .A(n42153), .B(n42152), .Z(n42154) );
  IV U54999 ( .A(n42154), .Z(n45515) );
  IV U55000 ( .A(n42155), .Z(n42156) );
  NOR U55001 ( .A(n42157), .B(n42156), .Z(n48946) );
  IV U55002 ( .A(n42158), .Z(n42160) );
  NOR U55003 ( .A(n42160), .B(n42159), .Z(n48938) );
  NOR U55004 ( .A(n48946), .B(n48938), .Z(n46857) );
  IV U55005 ( .A(n42161), .Z(n42162) );
  NOR U55006 ( .A(n42163), .B(n42162), .Z(n45521) );
  IV U55007 ( .A(n42164), .Z(n42166) );
  IV U55008 ( .A(n42165), .Z(n43450) );
  NOR U55009 ( .A(n42166), .B(n43450), .Z(n45523) );
  NOR U55010 ( .A(n45525), .B(n45523), .Z(n43448) );
  IV U55011 ( .A(n42167), .Z(n42169) );
  NOR U55012 ( .A(n42169), .B(n42168), .Z(n46848) );
  NOR U55013 ( .A(n46848), .B(n46846), .Z(n43446) );
  IV U55014 ( .A(n42170), .Z(n42171) );
  NOR U55015 ( .A(n42172), .B(n42171), .Z(n46835) );
  IV U55016 ( .A(n42173), .Z(n42174) );
  NOR U55017 ( .A(n42175), .B(n42174), .Z(n46829) );
  NOR U55018 ( .A(n46835), .B(n46829), .Z(n43445) );
  IV U55019 ( .A(n42176), .Z(n42177) );
  NOR U55020 ( .A(n42177), .B(n45536), .Z(n43444) );
  IV U55021 ( .A(n42178), .Z(n42182) );
  IV U55022 ( .A(n42179), .Z(n43434) );
  NOR U55023 ( .A(n42180), .B(n43434), .Z(n42181) );
  IV U55024 ( .A(n42181), .Z(n43431) );
  NOR U55025 ( .A(n42182), .B(n43431), .Z(n46793) );
  IV U55026 ( .A(n42183), .Z(n42184) );
  NOR U55027 ( .A(n42184), .B(n42189), .Z(n45543) );
  IV U55028 ( .A(n42185), .Z(n42186) );
  NOR U55029 ( .A(n42187), .B(n42186), .Z(n48968) );
  IV U55030 ( .A(n42188), .Z(n42190) );
  NOR U55031 ( .A(n42190), .B(n42189), .Z(n50223) );
  NOR U55032 ( .A(n48968), .B(n50223), .Z(n46797) );
  IV U55033 ( .A(n42191), .Z(n42192) );
  NOR U55034 ( .A(n42193), .B(n42192), .Z(n42194) );
  IV U55035 ( .A(n42194), .Z(n43417) );
  IV U55036 ( .A(n42195), .Z(n42198) );
  IV U55037 ( .A(n42196), .Z(n42197) );
  NOR U55038 ( .A(n42198), .B(n42197), .Z(n45553) );
  IV U55039 ( .A(n42199), .Z(n42201) );
  IV U55040 ( .A(n42200), .Z(n42203) );
  NOR U55041 ( .A(n42201), .B(n42203), .Z(n45550) );
  IV U55042 ( .A(n42202), .Z(n42206) );
  NOR U55043 ( .A(n42204), .B(n42203), .Z(n42205) );
  IV U55044 ( .A(n42205), .Z(n42208) );
  NOR U55045 ( .A(n42206), .B(n42208), .Z(n45547) );
  IV U55046 ( .A(n42207), .Z(n42209) );
  NOR U55047 ( .A(n42209), .B(n42208), .Z(n45560) );
  IV U55048 ( .A(n42210), .Z(n42211) );
  NOR U55049 ( .A(n42211), .B(n42217), .Z(n45557) );
  IV U55050 ( .A(n42212), .Z(n42214) );
  NOR U55051 ( .A(n42214), .B(n42213), .Z(n46768) );
  IV U55052 ( .A(n42215), .Z(n42216) );
  NOR U55053 ( .A(n42217), .B(n42216), .Z(n45564) );
  NOR U55054 ( .A(n46768), .B(n45564), .Z(n43409) );
  IV U55055 ( .A(n42218), .Z(n42219) );
  NOR U55056 ( .A(n42220), .B(n42219), .Z(n45566) );
  IV U55057 ( .A(n42221), .Z(n42222) );
  NOR U55058 ( .A(n42223), .B(n42222), .Z(n46771) );
  NOR U55059 ( .A(n45566), .B(n46771), .Z(n43408) );
  IV U55060 ( .A(n42224), .Z(n42227) );
  IV U55061 ( .A(n42225), .Z(n42226) );
  NOR U55062 ( .A(n42227), .B(n42226), .Z(n46752) );
  NOR U55063 ( .A(n42229), .B(n42228), .Z(n42230) );
  IV U55064 ( .A(n42230), .Z(n42234) );
  NOR U55065 ( .A(n42232), .B(n42231), .Z(n42233) );
  IV U55066 ( .A(n42233), .Z(n45569) );
  NOR U55067 ( .A(n42234), .B(n45569), .Z(n43395) );
  IV U55068 ( .A(n42235), .Z(n42237) );
  IV U55069 ( .A(n42236), .Z(n42241) );
  NOR U55070 ( .A(n42237), .B(n42241), .Z(n46744) );
  IV U55071 ( .A(n42238), .Z(n42239) );
  NOR U55072 ( .A(n42239), .B(n45569), .Z(n45573) );
  NOR U55073 ( .A(n46744), .B(n45573), .Z(n43393) );
  IV U55074 ( .A(n42240), .Z(n42242) );
  NOR U55075 ( .A(n42242), .B(n42241), .Z(n46741) );
  IV U55076 ( .A(n42243), .Z(n43379) );
  NOR U55077 ( .A(n42244), .B(n43379), .Z(n46731) );
  NOR U55078 ( .A(n42246), .B(n42245), .Z(n46727) );
  IV U55079 ( .A(n42247), .Z(n42248) );
  NOR U55080 ( .A(n42249), .B(n42248), .Z(n43375) );
  IV U55081 ( .A(n43375), .Z(n43373) );
  IV U55082 ( .A(n42250), .Z(n43371) );
  IV U55083 ( .A(n42251), .Z(n42252) );
  NOR U55084 ( .A(n43371), .B(n42252), .Z(n42253) );
  IV U55085 ( .A(n42253), .Z(n46708) );
  IV U55086 ( .A(n42254), .Z(n42255) );
  NOR U55087 ( .A(n42256), .B(n42255), .Z(n42257) );
  IV U55088 ( .A(n42257), .Z(n43345) );
  IV U55089 ( .A(n42258), .Z(n42260) );
  NOR U55090 ( .A(n42260), .B(n42259), .Z(n46696) );
  NOR U55091 ( .A(n42262), .B(n42261), .Z(n46693) );
  IV U55092 ( .A(n42263), .Z(n42266) );
  IV U55093 ( .A(n42264), .Z(n42265) );
  NOR U55094 ( .A(n42266), .B(n42265), .Z(n45599) );
  NOR U55095 ( .A(n42268), .B(n42267), .Z(n45605) );
  NOR U55096 ( .A(n42269), .B(n42268), .Z(n42270) );
  IV U55097 ( .A(n42270), .Z(n50096) );
  NOR U55098 ( .A(n42271), .B(n50096), .Z(n45606) );
  NOR U55099 ( .A(n45605), .B(n45606), .Z(n43331) );
  IV U55100 ( .A(n42272), .Z(n42274) );
  NOR U55101 ( .A(n42274), .B(n42273), .Z(n42275) );
  IV U55102 ( .A(n42275), .Z(n45614) );
  IV U55103 ( .A(n42276), .Z(n42277) );
  NOR U55104 ( .A(n42277), .B(n49067), .Z(n42280) );
  IV U55105 ( .A(n42278), .Z(n42279) );
  NOR U55106 ( .A(n42279), .B(n43280), .Z(n49058) );
  NOR U55107 ( .A(n42280), .B(n49058), .Z(n45621) );
  IV U55108 ( .A(n42281), .Z(n42283) );
  IV U55109 ( .A(n42282), .Z(n42285) );
  NOR U55110 ( .A(n42283), .B(n42285), .Z(n45618) );
  IV U55111 ( .A(n42284), .Z(n42286) );
  NOR U55112 ( .A(n42286), .B(n42285), .Z(n45623) );
  IV U55113 ( .A(n42287), .Z(n42288) );
  NOR U55114 ( .A(n42289), .B(n42288), .Z(n46651) );
  NOR U55115 ( .A(n42291), .B(n42290), .Z(n46647) );
  NOR U55116 ( .A(n46651), .B(n46647), .Z(n43271) );
  IV U55117 ( .A(n42292), .Z(n42297) );
  IV U55118 ( .A(n42293), .Z(n42295) );
  NOR U55119 ( .A(n42295), .B(n42294), .Z(n42296) );
  IV U55120 ( .A(n42296), .Z(n42301) );
  NOR U55121 ( .A(n42297), .B(n42301), .Z(n46655) );
  IV U55122 ( .A(n42298), .Z(n42299) );
  NOR U55123 ( .A(n42299), .B(n42301), .Z(n45628) );
  IV U55124 ( .A(n42300), .Z(n42304) );
  NOR U55125 ( .A(n42302), .B(n42301), .Z(n42303) );
  IV U55126 ( .A(n42303), .Z(n43269) );
  NOR U55127 ( .A(n42304), .B(n43269), .Z(n46642) );
  IV U55128 ( .A(n42305), .Z(n42308) );
  NOR U55129 ( .A(n42306), .B(n42310), .Z(n42307) );
  IV U55130 ( .A(n42307), .Z(n43264) );
  NOR U55131 ( .A(n42308), .B(n43264), .Z(n45632) );
  IV U55132 ( .A(n42309), .Z(n42311) );
  NOR U55133 ( .A(n42311), .B(n42310), .Z(n45637) );
  IV U55134 ( .A(n42312), .Z(n42313) );
  NOR U55135 ( .A(n42314), .B(n42313), .Z(n45648) );
  IV U55136 ( .A(n42315), .Z(n42317) );
  NOR U55137 ( .A(n42317), .B(n42316), .Z(n42318) );
  IV U55138 ( .A(n42318), .Z(n43240) );
  NOR U55139 ( .A(n42320), .B(n42319), .Z(n46620) );
  IV U55140 ( .A(n42321), .Z(n43233) );
  IV U55141 ( .A(n42322), .Z(n42323) );
  NOR U55142 ( .A(n43233), .B(n42323), .Z(n45655) );
  IV U55143 ( .A(n42324), .Z(n43225) );
  IV U55144 ( .A(n42325), .Z(n42326) );
  NOR U55145 ( .A(n43225), .B(n42326), .Z(n49086) );
  IV U55146 ( .A(n42327), .Z(n42328) );
  NOR U55147 ( .A(n42328), .B(n43235), .Z(n49995) );
  NOR U55148 ( .A(n49086), .B(n49995), .Z(n46609) );
  IV U55149 ( .A(n42329), .Z(n42332) );
  NOR U55150 ( .A(n42330), .B(n43217), .Z(n42331) );
  IV U55151 ( .A(n42331), .Z(n43221) );
  NOR U55152 ( .A(n42332), .B(n43221), .Z(n46595) );
  IV U55153 ( .A(n42333), .Z(n42338) );
  IV U55154 ( .A(n42334), .Z(n42335) );
  NOR U55155 ( .A(n42338), .B(n42335), .Z(n45664) );
  IV U55156 ( .A(n42336), .Z(n42337) );
  NOR U55157 ( .A(n42338), .B(n42337), .Z(n46599) );
  IV U55158 ( .A(n42339), .Z(n42341) );
  NOR U55159 ( .A(n42341), .B(n42340), .Z(n43199) );
  IV U55160 ( .A(n43199), .Z(n43194) );
  IV U55161 ( .A(n42342), .Z(n42343) );
  NOR U55162 ( .A(n42343), .B(n42348), .Z(n46560) );
  IV U55163 ( .A(n42344), .Z(n42345) );
  NOR U55164 ( .A(n42346), .B(n42345), .Z(n53721) );
  IV U55165 ( .A(n42347), .Z(n42349) );
  NOR U55166 ( .A(n42349), .B(n42348), .Z(n52923) );
  NOR U55167 ( .A(n53721), .B(n52923), .Z(n49134) );
  IV U55168 ( .A(n42350), .Z(n42353) );
  IV U55169 ( .A(n42351), .Z(n42352) );
  NOR U55170 ( .A(n42353), .B(n42352), .Z(n45691) );
  IV U55171 ( .A(n42354), .Z(n42355) );
  NOR U55172 ( .A(n42356), .B(n42355), .Z(n46536) );
  NOR U55173 ( .A(n42358), .B(n42357), .Z(n42363) );
  NOR U55174 ( .A(n42360), .B(n42359), .Z(n42361) );
  IV U55175 ( .A(n42361), .Z(n42362) );
  NOR U55176 ( .A(n42363), .B(n42362), .Z(n42364) );
  IV U55177 ( .A(n42364), .Z(n46541) );
  NOR U55178 ( .A(n42365), .B(n46541), .Z(n46533) );
  IV U55179 ( .A(n42366), .Z(n42371) );
  IV U55180 ( .A(n42367), .Z(n43150) );
  XOR U55181 ( .A(n43150), .B(n42375), .Z(n42368) );
  NOR U55182 ( .A(n42369), .B(n42368), .Z(n42370) );
  IV U55183 ( .A(n42370), .Z(n42373) );
  NOR U55184 ( .A(n42371), .B(n42373), .Z(n45701) );
  NOR U55185 ( .A(n46533), .B(n45701), .Z(n43156) );
  IV U55186 ( .A(n42372), .Z(n42374) );
  NOR U55187 ( .A(n42374), .B(n42373), .Z(n46520) );
  IV U55188 ( .A(n42375), .Z(n43151) );
  IV U55189 ( .A(n42376), .Z(n42377) );
  NOR U55190 ( .A(n43151), .B(n42377), .Z(n45703) );
  IV U55191 ( .A(n42378), .Z(n42383) );
  IV U55192 ( .A(n42379), .Z(n42380) );
  NOR U55193 ( .A(n42380), .B(n46504), .Z(n42381) );
  IV U55194 ( .A(n42381), .Z(n42382) );
  NOR U55195 ( .A(n42383), .B(n42382), .Z(n46494) );
  IV U55196 ( .A(n42384), .Z(n42386) );
  NOR U55197 ( .A(n42386), .B(n42385), .Z(n42387) );
  IV U55198 ( .A(n42387), .Z(n42388) );
  NOR U55199 ( .A(n42389), .B(n42388), .Z(n42390) );
  NOR U55200 ( .A(n46491), .B(n42390), .Z(n46498) );
  NOR U55201 ( .A(n42392), .B(n42391), .Z(n46488) );
  NOR U55202 ( .A(n42393), .B(n49202), .Z(n43109) );
  IV U55203 ( .A(n43109), .Z(n43099) );
  IV U55204 ( .A(n42394), .Z(n42396) );
  IV U55205 ( .A(n42395), .Z(n42401) );
  NOR U55206 ( .A(n42396), .B(n42401), .Z(n43102) );
  IV U55207 ( .A(n42397), .Z(n42399) );
  NOR U55208 ( .A(n42399), .B(n42398), .Z(n45719) );
  NOR U55209 ( .A(n43102), .B(n45719), .Z(n43097) );
  IV U55210 ( .A(n42400), .Z(n42402) );
  NOR U55211 ( .A(n42402), .B(n42401), .Z(n46479) );
  NOR U55212 ( .A(n46476), .B(n46479), .Z(n43096) );
  IV U55213 ( .A(n42403), .Z(n42404) );
  NOR U55214 ( .A(n42405), .B(n42404), .Z(n45723) );
  IV U55215 ( .A(n42406), .Z(n43090) );
  IV U55216 ( .A(n42407), .Z(n42408) );
  NOR U55217 ( .A(n43090), .B(n42408), .Z(n46468) );
  IV U55218 ( .A(n42409), .Z(n42412) );
  NOR U55219 ( .A(n42410), .B(n42417), .Z(n42411) );
  IV U55220 ( .A(n42411), .Z(n43086) );
  NOR U55221 ( .A(n42412), .B(n43086), .Z(n45731) );
  IV U55222 ( .A(n42413), .Z(n42415) );
  NOR U55223 ( .A(n42415), .B(n42414), .Z(n46465) );
  IV U55224 ( .A(n42416), .Z(n42418) );
  NOR U55225 ( .A(n42418), .B(n42417), .Z(n45737) );
  NOR U55226 ( .A(n46465), .B(n45737), .Z(n43083) );
  IV U55227 ( .A(n42419), .Z(n42420) );
  NOR U55228 ( .A(n42420), .B(n42422), .Z(n46452) );
  IV U55229 ( .A(n42421), .Z(n42423) );
  NOR U55230 ( .A(n42423), .B(n42422), .Z(n45739) );
  IV U55231 ( .A(n42424), .Z(n42425) );
  NOR U55232 ( .A(n42425), .B(n42433), .Z(n46450) );
  IV U55233 ( .A(n42426), .Z(n42428) );
  NOR U55234 ( .A(n42428), .B(n42427), .Z(n46456) );
  NOR U55235 ( .A(n46450), .B(n46456), .Z(n43082) );
  IV U55236 ( .A(n42429), .Z(n42431) );
  NOR U55237 ( .A(n42431), .B(n42430), .Z(n46442) );
  IV U55238 ( .A(n42432), .Z(n42434) );
  NOR U55239 ( .A(n42434), .B(n42433), .Z(n46446) );
  NOR U55240 ( .A(n46442), .B(n46446), .Z(n43081) );
  IV U55241 ( .A(n42435), .Z(n42436) );
  NOR U55242 ( .A(n42437), .B(n42436), .Z(n45746) );
  IV U55243 ( .A(n42438), .Z(n42440) );
  NOR U55244 ( .A(n42440), .B(n42439), .Z(n45743) );
  NOR U55245 ( .A(n49252), .B(n49250), .Z(n43070) );
  IV U55246 ( .A(n43070), .Z(n43065) );
  IV U55247 ( .A(n42441), .Z(n42442) );
  NOR U55248 ( .A(n42444), .B(n42442), .Z(n49261) );
  IV U55249 ( .A(n42443), .Z(n42447) );
  NOR U55250 ( .A(n42445), .B(n42444), .Z(n42446) );
  IV U55251 ( .A(n42446), .Z(n43063) );
  NOR U55252 ( .A(n42447), .B(n43063), .Z(n49256) );
  NOR U55253 ( .A(n49261), .B(n49256), .Z(n45763) );
  IV U55254 ( .A(n42448), .Z(n42449) );
  NOR U55255 ( .A(n43057), .B(n42449), .Z(n46415) );
  IV U55256 ( .A(n42450), .Z(n42456) );
  NOR U55257 ( .A(n42451), .B(n43052), .Z(n42452) );
  IV U55258 ( .A(n42452), .Z(n42453) );
  NOR U55259 ( .A(n42454), .B(n42453), .Z(n42455) );
  IV U55260 ( .A(n42455), .Z(n42458) );
  NOR U55261 ( .A(n42456), .B(n42458), .Z(n45769) );
  IV U55262 ( .A(n42457), .Z(n42459) );
  NOR U55263 ( .A(n42459), .B(n42458), .Z(n45766) );
  IV U55264 ( .A(n42460), .Z(n42461) );
  NOR U55265 ( .A(n42462), .B(n42461), .Z(n46394) );
  IV U55266 ( .A(n42463), .Z(n42465) );
  NOR U55267 ( .A(n42465), .B(n42464), .Z(n45779) );
  NOR U55268 ( .A(n46394), .B(n45779), .Z(n49283) );
  IV U55269 ( .A(n42466), .Z(n42467) );
  NOR U55270 ( .A(n42468), .B(n42467), .Z(n43033) );
  IV U55271 ( .A(n42469), .Z(n42470) );
  NOR U55272 ( .A(n42472), .B(n42470), .Z(n45785) );
  IV U55273 ( .A(n42471), .Z(n42475) );
  NOR U55274 ( .A(n42473), .B(n42472), .Z(n42474) );
  IV U55275 ( .A(n42474), .Z(n42477) );
  NOR U55276 ( .A(n42475), .B(n42477), .Z(n46382) );
  IV U55277 ( .A(n42476), .Z(n42478) );
  NOR U55278 ( .A(n42478), .B(n42477), .Z(n46388) );
  IV U55279 ( .A(n42479), .Z(n42480) );
  NOR U55280 ( .A(n42481), .B(n42480), .Z(n46378) );
  IV U55281 ( .A(n42482), .Z(n42483) );
  NOR U55282 ( .A(n42485), .B(n42483), .Z(n46368) );
  NOR U55283 ( .A(n42485), .B(n42484), .Z(n46364) );
  IV U55284 ( .A(n42486), .Z(n42487) );
  NOR U55285 ( .A(n42492), .B(n42487), .Z(n46361) );
  IV U55286 ( .A(n42488), .Z(n42489) );
  NOR U55287 ( .A(n42490), .B(n42489), .Z(n49306) );
  IV U55288 ( .A(n42491), .Z(n42493) );
  NOR U55289 ( .A(n42493), .B(n42492), .Z(n49798) );
  NOR U55290 ( .A(n49306), .B(n49798), .Z(n46359) );
  NOR U55291 ( .A(n42495), .B(n42494), .Z(n46345) );
  IV U55292 ( .A(n42496), .Z(n42500) );
  NOR U55293 ( .A(n42498), .B(n42497), .Z(n42499) );
  IV U55294 ( .A(n42499), .Z(n43024) );
  NOR U55295 ( .A(n42500), .B(n43024), .Z(n45788) );
  IV U55296 ( .A(n42501), .Z(n42503) );
  IV U55297 ( .A(n42502), .Z(n42505) );
  NOR U55298 ( .A(n42503), .B(n42505), .Z(n45798) );
  IV U55299 ( .A(n42504), .Z(n42506) );
  NOR U55300 ( .A(n42506), .B(n42505), .Z(n45794) );
  NOR U55301 ( .A(n45798), .B(n45794), .Z(n43022) );
  IV U55302 ( .A(n42507), .Z(n42508) );
  NOR U55303 ( .A(n42508), .B(n42513), .Z(n46337) );
  IV U55304 ( .A(n42509), .Z(n42510) );
  NOR U55305 ( .A(n42511), .B(n42510), .Z(n46329) );
  IV U55306 ( .A(n42512), .Z(n42514) );
  NOR U55307 ( .A(n42514), .B(n42513), .Z(n46334) );
  NOR U55308 ( .A(n46329), .B(n46334), .Z(n43021) );
  IV U55309 ( .A(n42515), .Z(n42516) );
  NOR U55310 ( .A(n42516), .B(n42518), .Z(n46323) );
  IV U55311 ( .A(n42517), .Z(n42519) );
  NOR U55312 ( .A(n42519), .B(n42518), .Z(n46308) );
  IV U55313 ( .A(n42520), .Z(n42523) );
  IV U55314 ( .A(n42521), .Z(n42522) );
  NOR U55315 ( .A(n42523), .B(n42522), .Z(n46311) );
  NOR U55316 ( .A(n46308), .B(n46311), .Z(n43007) );
  IV U55317 ( .A(n42524), .Z(n42525) );
  NOR U55318 ( .A(n42525), .B(n43001), .Z(n43005) );
  IV U55319 ( .A(n43005), .Z(n42997) );
  IV U55320 ( .A(n42526), .Z(n42529) );
  IV U55321 ( .A(n42527), .Z(n42528) );
  NOR U55322 ( .A(n42529), .B(n42528), .Z(n45807) );
  IV U55323 ( .A(n42530), .Z(n42531) );
  NOR U55324 ( .A(n42531), .B(n42533), .Z(n46295) );
  IV U55325 ( .A(n42532), .Z(n42534) );
  NOR U55326 ( .A(n42534), .B(n42533), .Z(n46287) );
  IV U55327 ( .A(n42535), .Z(n42536) );
  NOR U55328 ( .A(n42991), .B(n42536), .Z(n46284) );
  IV U55329 ( .A(n42537), .Z(n42538) );
  NOR U55330 ( .A(n42539), .B(n42538), .Z(n45810) );
  IV U55331 ( .A(n42540), .Z(n42541) );
  NOR U55332 ( .A(n42542), .B(n42541), .Z(n46276) );
  IV U55333 ( .A(n42543), .Z(n42544) );
  NOR U55334 ( .A(n42987), .B(n42544), .Z(n45821) );
  NOR U55335 ( .A(n46276), .B(n45821), .Z(n42984) );
  IV U55336 ( .A(n42545), .Z(n42546) );
  NOR U55337 ( .A(n42547), .B(n42546), .Z(n45825) );
  IV U55338 ( .A(n42548), .Z(n42550) );
  NOR U55339 ( .A(n42550), .B(n42549), .Z(n45823) );
  NOR U55340 ( .A(n45825), .B(n45823), .Z(n42977) );
  IV U55341 ( .A(n42551), .Z(n42552) );
  NOR U55342 ( .A(n42558), .B(n42552), .Z(n46257) );
  IV U55343 ( .A(n42553), .Z(n42554) );
  NOR U55344 ( .A(n42555), .B(n42554), .Z(n45835) );
  IV U55345 ( .A(n42556), .Z(n42557) );
  NOR U55346 ( .A(n42558), .B(n42557), .Z(n45830) );
  NOR U55347 ( .A(n45835), .B(n45830), .Z(n42965) );
  IV U55348 ( .A(n42559), .Z(n42562) );
  IV U55349 ( .A(n42560), .Z(n42561) );
  NOR U55350 ( .A(n42562), .B(n42561), .Z(n45833) );
  IV U55351 ( .A(n42563), .Z(n42564) );
  NOR U55352 ( .A(n42564), .B(n46237), .Z(n46242) );
  NOR U55353 ( .A(n42565), .B(n46237), .Z(n46247) );
  IV U55354 ( .A(n42566), .Z(n42571) );
  IV U55355 ( .A(n42567), .Z(n42568) );
  NOR U55356 ( .A(n42571), .B(n42568), .Z(n46233) );
  IV U55357 ( .A(n42569), .Z(n42573) );
  NOR U55358 ( .A(n42571), .B(n42570), .Z(n42572) );
  IV U55359 ( .A(n42572), .Z(n42575) );
  NOR U55360 ( .A(n42573), .B(n42575), .Z(n45838) );
  IV U55361 ( .A(n42574), .Z(n42576) );
  NOR U55362 ( .A(n42576), .B(n42575), .Z(n46222) );
  IV U55363 ( .A(n42577), .Z(n42578) );
  NOR U55364 ( .A(n42578), .B(n42953), .Z(n45841) );
  IV U55365 ( .A(n42579), .Z(n42582) );
  NOR U55366 ( .A(n42580), .B(n42587), .Z(n42581) );
  IV U55367 ( .A(n42581), .Z(n42948) );
  NOR U55368 ( .A(n42582), .B(n42948), .Z(n46198) );
  IV U55369 ( .A(n42583), .Z(n42959) );
  IV U55370 ( .A(n42584), .Z(n42585) );
  NOR U55371 ( .A(n42959), .B(n42585), .Z(n46195) );
  NOR U55372 ( .A(n46198), .B(n46195), .Z(n42951) );
  IV U55373 ( .A(n42586), .Z(n42590) );
  NOR U55374 ( .A(n42588), .B(n42587), .Z(n42589) );
  IV U55375 ( .A(n42589), .Z(n42945) );
  NOR U55376 ( .A(n42590), .B(n42945), .Z(n45846) );
  IV U55377 ( .A(n42591), .Z(n42592) );
  NOR U55378 ( .A(n42924), .B(n42592), .Z(n45860) );
  IV U55379 ( .A(n42593), .Z(n42594) );
  NOR U55380 ( .A(n42595), .B(n42594), .Z(n42596) );
  IV U55381 ( .A(n42596), .Z(n42929) );
  IV U55382 ( .A(n42597), .Z(n42598) );
  NOR U55383 ( .A(n42599), .B(n42598), .Z(n42600) );
  IV U55384 ( .A(n42600), .Z(n46186) );
  IV U55385 ( .A(n42601), .Z(n42606) );
  IV U55386 ( .A(n42602), .Z(n42603) );
  NOR U55387 ( .A(n42606), .B(n42603), .Z(n46182) );
  IV U55388 ( .A(n42604), .Z(n42605) );
  NOR U55389 ( .A(n42606), .B(n42605), .Z(n46178) );
  IV U55390 ( .A(n42607), .Z(n42608) );
  NOR U55391 ( .A(n42608), .B(n42914), .Z(n46175) );
  IV U55392 ( .A(n42609), .Z(n42610) );
  NOR U55393 ( .A(n42610), .B(n42914), .Z(n46171) );
  IV U55394 ( .A(n42611), .Z(n42612) );
  NOR U55395 ( .A(n42613), .B(n42612), .Z(n45878) );
  IV U55396 ( .A(n42614), .Z(n42884) );
  IV U55397 ( .A(n42615), .Z(n42871) );
  IV U55398 ( .A(n42616), .Z(n42617) );
  NOR U55399 ( .A(n42871), .B(n42617), .Z(n46148) );
  IV U55400 ( .A(n42618), .Z(n42620) );
  NOR U55401 ( .A(n42620), .B(n42619), .Z(n45890) );
  IV U55402 ( .A(n42621), .Z(n42622) );
  NOR U55403 ( .A(n42622), .B(n42874), .Z(n46138) );
  IV U55404 ( .A(n42623), .Z(n42626) );
  NOR U55405 ( .A(n42624), .B(n42632), .Z(n42625) );
  IV U55406 ( .A(n42625), .Z(n42629) );
  NOR U55407 ( .A(n42626), .B(n42629), .Z(n42627) );
  IV U55408 ( .A(n42627), .Z(n45904) );
  IV U55409 ( .A(n42628), .Z(n42630) );
  NOR U55410 ( .A(n42630), .B(n42629), .Z(n46130) );
  IV U55411 ( .A(n42631), .Z(n42633) );
  NOR U55412 ( .A(n42633), .B(n42632), .Z(n42634) );
  IV U55413 ( .A(n42634), .Z(n46129) );
  NOR U55414 ( .A(n42636), .B(n42635), .Z(n42637) );
  IV U55415 ( .A(n42637), .Z(n46115) );
  IV U55416 ( .A(n42638), .Z(n42639) );
  NOR U55417 ( .A(n42640), .B(n42639), .Z(n45921) );
  IV U55418 ( .A(n42641), .Z(n42643) );
  NOR U55419 ( .A(n42643), .B(n42642), .Z(n46103) );
  NOR U55420 ( .A(n45921), .B(n46103), .Z(n42824) );
  IV U55421 ( .A(n42644), .Z(n42645) );
  NOR U55422 ( .A(n42645), .B(n42648), .Z(n46086) );
  XOR U55423 ( .A(n42647), .B(n42646), .Z(n42652) );
  NOR U55424 ( .A(n42649), .B(n42648), .Z(n42650) );
  IV U55425 ( .A(n42650), .Z(n42651) );
  NOR U55426 ( .A(n42652), .B(n42651), .Z(n45923) );
  IV U55427 ( .A(n42653), .Z(n42819) );
  IV U55428 ( .A(n42654), .Z(n42655) );
  NOR U55429 ( .A(n42819), .B(n42655), .Z(n46090) );
  IV U55430 ( .A(n42656), .Z(n42657) );
  NOR U55431 ( .A(n42796), .B(n42657), .Z(n46080) );
  IV U55432 ( .A(n42658), .Z(n42791) );
  IV U55433 ( .A(n42659), .Z(n42660) );
  NOR U55434 ( .A(n42791), .B(n42660), .Z(n46061) );
  NOR U55435 ( .A(n45943), .B(n46061), .Z(n42789) );
  NOR U55436 ( .A(n42662), .B(n42661), .Z(n45946) );
  NOR U55437 ( .A(n45950), .B(n46047), .Z(n42779) );
  IV U55438 ( .A(n42663), .Z(n42665) );
  NOR U55439 ( .A(n42665), .B(n42664), .Z(n45952) );
  IV U55440 ( .A(n42666), .Z(n42667) );
  NOR U55441 ( .A(n42667), .B(n42759), .Z(n42668) );
  IV U55442 ( .A(n42668), .Z(n46034) );
  IV U55443 ( .A(n42669), .Z(n42670) );
  NOR U55444 ( .A(n42670), .B(n42759), .Z(n46030) );
  IV U55445 ( .A(n42671), .Z(n42675) );
  IV U55446 ( .A(n42672), .Z(n42677) );
  NOR U55447 ( .A(n42673), .B(n42677), .Z(n42674) );
  IV U55448 ( .A(n42674), .Z(n42755) );
  NOR U55449 ( .A(n42675), .B(n42755), .Z(n46025) );
  NOR U55450 ( .A(n42677), .B(n42676), .Z(n45962) );
  NOR U55451 ( .A(n42679), .B(n42678), .Z(n45959) );
  IV U55452 ( .A(n42680), .Z(n42681) );
  NOR U55453 ( .A(n42681), .B(n42743), .Z(n42682) );
  IV U55454 ( .A(n42682), .Z(n45971) );
  IV U55455 ( .A(n42683), .Z(n42688) );
  IV U55456 ( .A(n42684), .Z(n42685) );
  NOR U55457 ( .A(n42686), .B(n42685), .Z(n42687) );
  IV U55458 ( .A(n42687), .Z(n42731) );
  NOR U55459 ( .A(n42688), .B(n42731), .Z(n45979) );
  IV U55460 ( .A(n42689), .Z(n42691) );
  XOR U55461 ( .A(n42692), .B(n42695), .Z(n42690) );
  NOR U55462 ( .A(n42691), .B(n42690), .Z(n45982) );
  IV U55463 ( .A(n42692), .Z(n42693) );
  NOR U55464 ( .A(n42693), .B(n42695), .Z(n45992) );
  IV U55465 ( .A(n42694), .Z(n42696) );
  NOR U55466 ( .A(n42696), .B(n42695), .Z(n45984) );
  NOR U55467 ( .A(n45992), .B(n45984), .Z(n42697) );
  IV U55468 ( .A(n42697), .Z(n42698) );
  NOR U55469 ( .A(n45982), .B(n42698), .Z(n42728) );
  IV U55470 ( .A(n42699), .Z(n42701) );
  IV U55471 ( .A(n42700), .Z(n42706) );
  NOR U55472 ( .A(n42701), .B(n42706), .Z(n45987) );
  IV U55473 ( .A(n45987), .Z(n45989) );
  NOR U55474 ( .A(n42703), .B(n42702), .Z(n45995) );
  IV U55475 ( .A(n42704), .Z(n42705) );
  NOR U55476 ( .A(n42706), .B(n42705), .Z(n45997) );
  NOR U55477 ( .A(n45995), .B(n45997), .Z(n42727) );
  IV U55478 ( .A(n42707), .Z(n42708) );
  NOR U55479 ( .A(n42709), .B(n42708), .Z(n42711) );
  NOR U55480 ( .A(n42711), .B(n42710), .Z(n46002) );
  NOR U55481 ( .A(n42713), .B(n42712), .Z(n42722) );
  NOR U55482 ( .A(n42715), .B(n42714), .Z(n42720) );
  NOR U55483 ( .A(n42717), .B(n42716), .Z(n42718) );
  IV U55484 ( .A(n42718), .Z(n42719) );
  NOR U55485 ( .A(n42720), .B(n42719), .Z(n42721) );
  NOR U55486 ( .A(n42722), .B(n42721), .Z(n45999) );
  IV U55487 ( .A(n45999), .Z(n46001) );
  IV U55488 ( .A(n42723), .Z(n42725) );
  NOR U55489 ( .A(n42725), .B(n42724), .Z(n45998) );
  IV U55490 ( .A(n45998), .Z(n46000) );
  XOR U55491 ( .A(n46001), .B(n46000), .Z(n42726) );
  XOR U55492 ( .A(n46002), .B(n42726), .Z(n45996) );
  XOR U55493 ( .A(n42727), .B(n45996), .Z(n45988) );
  XOR U55494 ( .A(n45989), .B(n45988), .Z(n45985) );
  XOR U55495 ( .A(n42728), .B(n45985), .Z(n42729) );
  IV U55496 ( .A(n42729), .Z(n45981) );
  XOR U55497 ( .A(n45979), .B(n45981), .Z(n46013) );
  IV U55498 ( .A(n42730), .Z(n42732) );
  NOR U55499 ( .A(n42732), .B(n42731), .Z(n46011) );
  XOR U55500 ( .A(n46013), .B(n46011), .Z(n46020) );
  IV U55501 ( .A(n46020), .Z(n42740) );
  IV U55502 ( .A(n42733), .Z(n42734) );
  NOR U55503 ( .A(n42735), .B(n42734), .Z(n46007) );
  IV U55504 ( .A(n42736), .Z(n42737) );
  NOR U55505 ( .A(n42738), .B(n42737), .Z(n46019) );
  NOR U55506 ( .A(n46007), .B(n46019), .Z(n42739) );
  XOR U55507 ( .A(n42740), .B(n42739), .Z(n45978) );
  IV U55508 ( .A(n42741), .Z(n42742) );
  NOR U55509 ( .A(n42743), .B(n42742), .Z(n45976) );
  XOR U55510 ( .A(n45978), .B(n45976), .Z(n45972) );
  XOR U55511 ( .A(n45971), .B(n45972), .Z(n45969) );
  IV U55512 ( .A(n42744), .Z(n42745) );
  NOR U55513 ( .A(n42746), .B(n42745), .Z(n45973) );
  IV U55514 ( .A(n42747), .Z(n42749) );
  NOR U55515 ( .A(n42749), .B(n42748), .Z(n45968) );
  NOR U55516 ( .A(n45973), .B(n45968), .Z(n42750) );
  XOR U55517 ( .A(n45969), .B(n42750), .Z(n45967) );
  XOR U55518 ( .A(n45965), .B(n45967), .Z(n45960) );
  XOR U55519 ( .A(n45959), .B(n45960), .Z(n45963) );
  XOR U55520 ( .A(n45962), .B(n45963), .Z(n49603) );
  IV U55521 ( .A(n49603), .Z(n42757) );
  IV U55522 ( .A(n42751), .Z(n42752) );
  NOR U55523 ( .A(n42753), .B(n42752), .Z(n53321) );
  IV U55524 ( .A(n42754), .Z(n42756) );
  NOR U55525 ( .A(n42756), .B(n42755), .Z(n53316) );
  NOR U55526 ( .A(n53321), .B(n53316), .Z(n49605) );
  XOR U55527 ( .A(n42757), .B(n49605), .Z(n46027) );
  XOR U55528 ( .A(n46025), .B(n46027), .Z(n46031) );
  XOR U55529 ( .A(n46030), .B(n46031), .Z(n46033) );
  XOR U55530 ( .A(n46034), .B(n46033), .Z(n42764) );
  IV U55531 ( .A(n42764), .Z(n42762) );
  IV U55532 ( .A(n42758), .Z(n42760) );
  NOR U55533 ( .A(n42760), .B(n42759), .Z(n42763) );
  IV U55534 ( .A(n42763), .Z(n42761) );
  NOR U55535 ( .A(n42762), .B(n42761), .Z(n49523) );
  NOR U55536 ( .A(n42764), .B(n42763), .Z(n46041) );
  IV U55537 ( .A(n42765), .Z(n42771) );
  IV U55538 ( .A(n42766), .Z(n42767) );
  NOR U55539 ( .A(n42771), .B(n42767), .Z(n46039) );
  XOR U55540 ( .A(n46041), .B(n46039), .Z(n42768) );
  NOR U55541 ( .A(n49523), .B(n42768), .Z(n46036) );
  IV U55542 ( .A(n42769), .Z(n42770) );
  NOR U55543 ( .A(n42771), .B(n42770), .Z(n42772) );
  IV U55544 ( .A(n42772), .Z(n46037) );
  XOR U55545 ( .A(n46036), .B(n46037), .Z(n53373) );
  IV U55546 ( .A(n53373), .Z(n42778) );
  IV U55547 ( .A(n42773), .Z(n42774) );
  NOR U55548 ( .A(n42774), .B(n42776), .Z(n53379) );
  IV U55549 ( .A(n42775), .Z(n42777) );
  NOR U55550 ( .A(n42777), .B(n42776), .Z(n53368) );
  NOR U55551 ( .A(n53379), .B(n53368), .Z(n45958) );
  XOR U55552 ( .A(n42778), .B(n45958), .Z(n45954) );
  XOR U55553 ( .A(n45952), .B(n45954), .Z(n45956) );
  XOR U55554 ( .A(n45955), .B(n45956), .Z(n46048) );
  XOR U55555 ( .A(n42779), .B(n46048), .Z(n42780) );
  IV U55556 ( .A(n42780), .Z(n46052) );
  XOR U55557 ( .A(n46050), .B(n46052), .Z(n46058) );
  IV U55558 ( .A(n46058), .Z(n42788) );
  IV U55559 ( .A(n42781), .Z(n42782) );
  NOR U55560 ( .A(n42783), .B(n42782), .Z(n46053) );
  IV U55561 ( .A(n42784), .Z(n42786) );
  NOR U55562 ( .A(n42786), .B(n42785), .Z(n46057) );
  NOR U55563 ( .A(n46053), .B(n46057), .Z(n42787) );
  XOR U55564 ( .A(n42788), .B(n42787), .Z(n45948) );
  XOR U55565 ( .A(n45946), .B(n45948), .Z(n46066) );
  XOR U55566 ( .A(n46065), .B(n46066), .Z(n46062) );
  XOR U55567 ( .A(n42789), .B(n46062), .Z(n46077) );
  IV U55568 ( .A(n42790), .Z(n42792) );
  NOR U55569 ( .A(n42792), .B(n42791), .Z(n42793) );
  IV U55570 ( .A(n42793), .Z(n46078) );
  XOR U55571 ( .A(n46077), .B(n46078), .Z(n46081) );
  XOR U55572 ( .A(n46080), .B(n46081), .Z(n45941) );
  IV U55573 ( .A(n42794), .Z(n42795) );
  NOR U55574 ( .A(n42796), .B(n42795), .Z(n45940) );
  IV U55575 ( .A(n42797), .Z(n42799) );
  NOR U55576 ( .A(n42799), .B(n42798), .Z(n45938) );
  NOR U55577 ( .A(n45940), .B(n45938), .Z(n42800) );
  XOR U55578 ( .A(n45941), .B(n42800), .Z(n42813) );
  IV U55579 ( .A(n42813), .Z(n49487) );
  IV U55580 ( .A(n42801), .Z(n42802) );
  NOR U55581 ( .A(n42802), .B(n42821), .Z(n42815) );
  IV U55582 ( .A(n42815), .Z(n42803) );
  NOR U55583 ( .A(n49487), .B(n42803), .Z(n49481) );
  IV U55584 ( .A(n42804), .Z(n42805) );
  NOR U55585 ( .A(n42821), .B(n42805), .Z(n42806) );
  IV U55586 ( .A(n42806), .Z(n45935) );
  IV U55587 ( .A(n42807), .Z(n42808) );
  NOR U55588 ( .A(n42809), .B(n42808), .Z(n49493) );
  IV U55589 ( .A(n42810), .Z(n42811) );
  NOR U55590 ( .A(n42812), .B(n42811), .Z(n49485) );
  NOR U55591 ( .A(n49493), .B(n49485), .Z(n45934) );
  XOR U55592 ( .A(n42813), .B(n45934), .Z(n45936) );
  XOR U55593 ( .A(n45935), .B(n45936), .Z(n42814) );
  NOR U55594 ( .A(n42815), .B(n42814), .Z(n42816) );
  NOR U55595 ( .A(n49481), .B(n42816), .Z(n45928) );
  IV U55596 ( .A(n42817), .Z(n42818) );
  NOR U55597 ( .A(n42819), .B(n42818), .Z(n45927) );
  IV U55598 ( .A(n42820), .Z(n42822) );
  NOR U55599 ( .A(n42822), .B(n42821), .Z(n45931) );
  NOR U55600 ( .A(n45927), .B(n45931), .Z(n42823) );
  XOR U55601 ( .A(n45928), .B(n42823), .Z(n46092) );
  XOR U55602 ( .A(n46090), .B(n46092), .Z(n45924) );
  XOR U55603 ( .A(n45923), .B(n45924), .Z(n46088) );
  XOR U55604 ( .A(n46086), .B(n46088), .Z(n46104) );
  XOR U55605 ( .A(n42824), .B(n46104), .Z(n45919) );
  NOR U55606 ( .A(n42826), .B(n42825), .Z(n46106) );
  IV U55607 ( .A(n42827), .Z(n42829) );
  IV U55608 ( .A(n42828), .Z(n42832) );
  NOR U55609 ( .A(n42829), .B(n42832), .Z(n45918) );
  NOR U55610 ( .A(n46106), .B(n45918), .Z(n42830) );
  XOR U55611 ( .A(n45919), .B(n42830), .Z(n45917) );
  IV U55612 ( .A(n45917), .Z(n42840) );
  IV U55613 ( .A(n42831), .Z(n42833) );
  NOR U55614 ( .A(n42833), .B(n42832), .Z(n45915) );
  IV U55615 ( .A(n42834), .Z(n42836) );
  NOR U55616 ( .A(n42836), .B(n42835), .Z(n45912) );
  NOR U55617 ( .A(n45915), .B(n45912), .Z(n42837) );
  IV U55618 ( .A(n42837), .Z(n42838) );
  NOR U55619 ( .A(n45910), .B(n42838), .Z(n42839) );
  XOR U55620 ( .A(n42840), .B(n42839), .Z(n46118) );
  XOR U55621 ( .A(n46115), .B(n46118), .Z(n45907) );
  IV U55622 ( .A(n42841), .Z(n42843) );
  NOR U55623 ( .A(n42843), .B(n42842), .Z(n46117) );
  IV U55624 ( .A(n42844), .Z(n42846) );
  NOR U55625 ( .A(n42846), .B(n42845), .Z(n45906) );
  NOR U55626 ( .A(n46117), .B(n45906), .Z(n42847) );
  XOR U55627 ( .A(n45907), .B(n42847), .Z(n46123) );
  IV U55628 ( .A(n42848), .Z(n42850) );
  NOR U55629 ( .A(n42850), .B(n42849), .Z(n42851) );
  IV U55630 ( .A(n42851), .Z(n42859) );
  NOR U55631 ( .A(n46123), .B(n42859), .Z(n49461) );
  IV U55632 ( .A(n42852), .Z(n42854) );
  NOR U55633 ( .A(n42854), .B(n42853), .Z(n42855) );
  IV U55634 ( .A(n42855), .Z(n46126) );
  IV U55635 ( .A(n42856), .Z(n42858) );
  NOR U55636 ( .A(n42858), .B(n42857), .Z(n46121) );
  XOR U55637 ( .A(n46121), .B(n46123), .Z(n46125) );
  XOR U55638 ( .A(n46126), .B(n46125), .Z(n42862) );
  IV U55639 ( .A(n46125), .Z(n42860) );
  NOR U55640 ( .A(n42860), .B(n42859), .Z(n42861) );
  NOR U55641 ( .A(n42862), .B(n42861), .Z(n42863) );
  NOR U55642 ( .A(n49461), .B(n42863), .Z(n46127) );
  XOR U55643 ( .A(n46129), .B(n46127), .Z(n46131) );
  XOR U55644 ( .A(n46130), .B(n46131), .Z(n45905) );
  XOR U55645 ( .A(n45904), .B(n45905), .Z(n45897) );
  IV U55646 ( .A(n42864), .Z(n45898) );
  NOR U55647 ( .A(n42865), .B(n45898), .Z(n42868) );
  IV U55648 ( .A(n42866), .Z(n42867) );
  NOR U55649 ( .A(n42867), .B(n42874), .Z(n46135) );
  NOR U55650 ( .A(n42868), .B(n46135), .Z(n42869) );
  XOR U55651 ( .A(n45897), .B(n42869), .Z(n46140) );
  XOR U55652 ( .A(n46138), .B(n46140), .Z(n46143) );
  IV U55653 ( .A(n46143), .Z(n42876) );
  NOR U55654 ( .A(n42871), .B(n42870), .Z(n45894) );
  IV U55655 ( .A(n42872), .Z(n42873) );
  NOR U55656 ( .A(n42874), .B(n42873), .Z(n46141) );
  NOR U55657 ( .A(n45894), .B(n46141), .Z(n42875) );
  XOR U55658 ( .A(n42876), .B(n42875), .Z(n45891) );
  XOR U55659 ( .A(n45890), .B(n45891), .Z(n46150) );
  XOR U55660 ( .A(n46148), .B(n46150), .Z(n45888) );
  NOR U55661 ( .A(n42885), .B(n45888), .Z(n42877) );
  IV U55662 ( .A(n42877), .Z(n49721) );
  NOR U55663 ( .A(n42884), .B(n49721), .Z(n45886) );
  IV U55664 ( .A(n42878), .Z(n49724) );
  NOR U55665 ( .A(n49724), .B(n42879), .Z(n42880) );
  IV U55666 ( .A(n42880), .Z(n45882) );
  IV U55667 ( .A(n42881), .Z(n42882) );
  NOR U55668 ( .A(n42883), .B(n42882), .Z(n45887) );
  XOR U55669 ( .A(n45887), .B(n45888), .Z(n45881) );
  XOR U55670 ( .A(n45882), .B(n45881), .Z(n42890) );
  IV U55671 ( .A(n45881), .Z(n42888) );
  NOR U55672 ( .A(n42885), .B(n42884), .Z(n42886) );
  IV U55673 ( .A(n42886), .Z(n42887) );
  NOR U55674 ( .A(n42888), .B(n42887), .Z(n42889) );
  NOR U55675 ( .A(n42890), .B(n42889), .Z(n42891) );
  NOR U55676 ( .A(n45886), .B(n42891), .Z(n42892) );
  IV U55677 ( .A(n42892), .Z(n45879) );
  XOR U55678 ( .A(n45878), .B(n45879), .Z(n45875) );
  IV U55679 ( .A(n42893), .Z(n42894) );
  NOR U55680 ( .A(n42895), .B(n42894), .Z(n45876) );
  IV U55681 ( .A(n42896), .Z(n42897) );
  NOR U55682 ( .A(n42897), .B(n42903), .Z(n45873) );
  NOR U55683 ( .A(n45876), .B(n45873), .Z(n42898) );
  XOR U55684 ( .A(n45875), .B(n42898), .Z(n45870) );
  IV U55685 ( .A(n42899), .Z(n42911) );
  IV U55686 ( .A(n42900), .Z(n42901) );
  NOR U55687 ( .A(n42911), .B(n42901), .Z(n46160) );
  IV U55688 ( .A(n42902), .Z(n42904) );
  NOR U55689 ( .A(n42904), .B(n42903), .Z(n45871) );
  NOR U55690 ( .A(n46160), .B(n45871), .Z(n42905) );
  XOR U55691 ( .A(n45870), .B(n42905), .Z(n46164) );
  IV U55692 ( .A(n42906), .Z(n42907) );
  NOR U55693 ( .A(n42908), .B(n42907), .Z(n45868) );
  IV U55694 ( .A(n42909), .Z(n42910) );
  NOR U55695 ( .A(n42911), .B(n42910), .Z(n46163) );
  NOR U55696 ( .A(n45868), .B(n46163), .Z(n42912) );
  XOR U55697 ( .A(n46164), .B(n42912), .Z(n46168) );
  IV U55698 ( .A(n42913), .Z(n42915) );
  NOR U55699 ( .A(n42915), .B(n42914), .Z(n42916) );
  IV U55700 ( .A(n42916), .Z(n46169) );
  XOR U55701 ( .A(n46168), .B(n46169), .Z(n46173) );
  XOR U55702 ( .A(n46171), .B(n46173), .Z(n46177) );
  XOR U55703 ( .A(n46175), .B(n46177), .Z(n46180) );
  XOR U55704 ( .A(n46178), .B(n46180), .Z(n46184) );
  XOR U55705 ( .A(n46182), .B(n46184), .Z(n46185) );
  XOR U55706 ( .A(n46186), .B(n46185), .Z(n42926) );
  IV U55707 ( .A(n42926), .Z(n42917) );
  NOR U55708 ( .A(n42929), .B(n42917), .Z(n49748) );
  IV U55709 ( .A(n42918), .Z(n42920) );
  NOR U55710 ( .A(n42920), .B(n42919), .Z(n42921) );
  IV U55711 ( .A(n42921), .Z(n45867) );
  IV U55712 ( .A(n42922), .Z(n42923) );
  NOR U55713 ( .A(n42924), .B(n42923), .Z(n42927) );
  IV U55714 ( .A(n42927), .Z(n42925) );
  NOR U55715 ( .A(n42925), .B(n46185), .Z(n49746) );
  NOR U55716 ( .A(n42927), .B(n42926), .Z(n42928) );
  NOR U55717 ( .A(n49746), .B(n42928), .Z(n42930) );
  IV U55718 ( .A(n42930), .Z(n45866) );
  XOR U55719 ( .A(n45867), .B(n45866), .Z(n42932) );
  NOR U55720 ( .A(n42930), .B(n42929), .Z(n42931) );
  NOR U55721 ( .A(n42932), .B(n42931), .Z(n42933) );
  NOR U55722 ( .A(n49748), .B(n42933), .Z(n42934) );
  IV U55723 ( .A(n42934), .Z(n45861) );
  XOR U55724 ( .A(n45860), .B(n45861), .Z(n45865) );
  IV U55725 ( .A(n42935), .Z(n42937) );
  NOR U55726 ( .A(n42937), .B(n42936), .Z(n45863) );
  XOR U55727 ( .A(n45865), .B(n45863), .Z(n45856) );
  IV U55728 ( .A(n42938), .Z(n42943) );
  IV U55729 ( .A(n42939), .Z(n42940) );
  NOR U55730 ( .A(n42943), .B(n42940), .Z(n45854) );
  XOR U55731 ( .A(n45856), .B(n45854), .Z(n45859) );
  IV U55732 ( .A(n42941), .Z(n42942) );
  NOR U55733 ( .A(n42943), .B(n42942), .Z(n45857) );
  XOR U55734 ( .A(n45859), .B(n45857), .Z(n45847) );
  XOR U55735 ( .A(n45846), .B(n45847), .Z(n45853) );
  IV U55736 ( .A(n42944), .Z(n42946) );
  NOR U55737 ( .A(n42946), .B(n42945), .Z(n45851) );
  IV U55738 ( .A(n42947), .Z(n42949) );
  NOR U55739 ( .A(n42949), .B(n42948), .Z(n45849) );
  NOR U55740 ( .A(n45851), .B(n45849), .Z(n42950) );
  XOR U55741 ( .A(n45853), .B(n42950), .Z(n46194) );
  XOR U55742 ( .A(n42951), .B(n46194), .Z(n46211) );
  IV U55743 ( .A(n42952), .Z(n42956) );
  NOR U55744 ( .A(n42954), .B(n42953), .Z(n42955) );
  IV U55745 ( .A(n42955), .Z(n42962) );
  NOR U55746 ( .A(n42956), .B(n42962), .Z(n46209) );
  IV U55747 ( .A(n42957), .Z(n42958) );
  NOR U55748 ( .A(n42959), .B(n42958), .Z(n45844) );
  NOR U55749 ( .A(n46209), .B(n45844), .Z(n42960) );
  XOR U55750 ( .A(n46211), .B(n42960), .Z(n46214) );
  IV U55751 ( .A(n42961), .Z(n42963) );
  NOR U55752 ( .A(n42963), .B(n42962), .Z(n42964) );
  IV U55753 ( .A(n42964), .Z(n46215) );
  XOR U55754 ( .A(n46214), .B(n46215), .Z(n45842) );
  XOR U55755 ( .A(n45841), .B(n45842), .Z(n46223) );
  XOR U55756 ( .A(n46222), .B(n46223), .Z(n45840) );
  XOR U55757 ( .A(n45838), .B(n45840), .Z(n46235) );
  XOR U55758 ( .A(n46233), .B(n46235), .Z(n46248) );
  XOR U55759 ( .A(n46247), .B(n46248), .Z(n46244) );
  XOR U55760 ( .A(n46242), .B(n46244), .Z(n45836) );
  XOR U55761 ( .A(n45833), .B(n45836), .Z(n45832) );
  XOR U55762 ( .A(n42965), .B(n45832), .Z(n42966) );
  IV U55763 ( .A(n42966), .Z(n46259) );
  XOR U55764 ( .A(n46257), .B(n46259), .Z(n46261) );
  IV U55765 ( .A(n46261), .Z(n42973) );
  IV U55766 ( .A(n42967), .Z(n42968) );
  NOR U55767 ( .A(n42969), .B(n42968), .Z(n46260) );
  IV U55768 ( .A(n42970), .Z(n42971) );
  NOR U55769 ( .A(n42975), .B(n42971), .Z(n45828) );
  NOR U55770 ( .A(n46260), .B(n45828), .Z(n42972) );
  XOR U55771 ( .A(n42973), .B(n42972), .Z(n46268) );
  IV U55772 ( .A(n42974), .Z(n42976) );
  NOR U55773 ( .A(n42976), .B(n42975), .Z(n46266) );
  XOR U55774 ( .A(n46268), .B(n46266), .Z(n45826) );
  XOR U55775 ( .A(n42977), .B(n45826), .Z(n46274) );
  IV U55776 ( .A(n42978), .Z(n42980) );
  NOR U55777 ( .A(n42980), .B(n42979), .Z(n49377) );
  IV U55778 ( .A(n42981), .Z(n42983) );
  NOR U55779 ( .A(n42983), .B(n42982), .Z(n49373) );
  NOR U55780 ( .A(n49377), .B(n49373), .Z(n46275) );
  XOR U55781 ( .A(n46274), .B(n46275), .Z(n46277) );
  XOR U55782 ( .A(n42984), .B(n46277), .Z(n42985) );
  IV U55783 ( .A(n42985), .Z(n45817) );
  IV U55784 ( .A(n42986), .Z(n42988) );
  NOR U55785 ( .A(n42988), .B(n42987), .Z(n45815) );
  XOR U55786 ( .A(n45817), .B(n45815), .Z(n45820) );
  IV U55787 ( .A(n45820), .Z(n42996) );
  IV U55788 ( .A(n42989), .Z(n42990) );
  NOR U55789 ( .A(n42991), .B(n42990), .Z(n45813) );
  IV U55790 ( .A(n42992), .Z(n42994) );
  NOR U55791 ( .A(n42994), .B(n42993), .Z(n45818) );
  NOR U55792 ( .A(n45813), .B(n45818), .Z(n42995) );
  XOR U55793 ( .A(n42996), .B(n42995), .Z(n45811) );
  XOR U55794 ( .A(n45810), .B(n45811), .Z(n46285) );
  XOR U55795 ( .A(n46284), .B(n46285), .Z(n46288) );
  XOR U55796 ( .A(n46287), .B(n46288), .Z(n46297) );
  XOR U55797 ( .A(n46295), .B(n46297), .Z(n45808) );
  XOR U55798 ( .A(n45807), .B(n45808), .Z(n46294) );
  NOR U55799 ( .A(n42997), .B(n46294), .Z(n45804) );
  IV U55800 ( .A(n42998), .Z(n42999) );
  NOR U55801 ( .A(n42999), .B(n43001), .Z(n46292) );
  XOR U55802 ( .A(n46294), .B(n46292), .Z(n45806) );
  IV U55803 ( .A(n43000), .Z(n43002) );
  NOR U55804 ( .A(n43002), .B(n43001), .Z(n43003) );
  IV U55805 ( .A(n43003), .Z(n45805) );
  XOR U55806 ( .A(n45806), .B(n45805), .Z(n43004) );
  NOR U55807 ( .A(n43005), .B(n43004), .Z(n43006) );
  NOR U55808 ( .A(n45804), .B(n43006), .Z(n46309) );
  XOR U55809 ( .A(n43007), .B(n46309), .Z(n45803) );
  IV U55810 ( .A(n43008), .Z(n43010) );
  NOR U55811 ( .A(n43010), .B(n43009), .Z(n45801) );
  XOR U55812 ( .A(n45803), .B(n45801), .Z(n46324) );
  XOR U55813 ( .A(n46323), .B(n46324), .Z(n49331) );
  IV U55814 ( .A(n43011), .Z(n43012) );
  NOR U55815 ( .A(n43018), .B(n43012), .Z(n49332) );
  IV U55816 ( .A(n43013), .Z(n43014) );
  NOR U55817 ( .A(n43015), .B(n43014), .Z(n49330) );
  IV U55818 ( .A(n43016), .Z(n43017) );
  NOR U55819 ( .A(n43018), .B(n43017), .Z(n49337) );
  NOR U55820 ( .A(n49330), .B(n49337), .Z(n46328) );
  IV U55821 ( .A(n46328), .Z(n43019) );
  NOR U55822 ( .A(n49332), .B(n43019), .Z(n43020) );
  XOR U55823 ( .A(n49331), .B(n43020), .Z(n46330) );
  XOR U55824 ( .A(n43021), .B(n46330), .Z(n46338) );
  XOR U55825 ( .A(n46337), .B(n46338), .Z(n45799) );
  XOR U55826 ( .A(n43022), .B(n45799), .Z(n45791) );
  IV U55827 ( .A(n43023), .Z(n43025) );
  NOR U55828 ( .A(n43025), .B(n43024), .Z(n43026) );
  IV U55829 ( .A(n43026), .Z(n45792) );
  XOR U55830 ( .A(n45791), .B(n45792), .Z(n45790) );
  XOR U55831 ( .A(n45788), .B(n45790), .Z(n46343) );
  XOR U55832 ( .A(n46342), .B(n46343), .Z(n46346) );
  XOR U55833 ( .A(n46345), .B(n46346), .Z(n49308) );
  XOR U55834 ( .A(n46359), .B(n49308), .Z(n43027) );
  IV U55835 ( .A(n43027), .Z(n46362) );
  XOR U55836 ( .A(n46361), .B(n46362), .Z(n46365) );
  XOR U55837 ( .A(n46364), .B(n46365), .Z(n46369) );
  XOR U55838 ( .A(n46368), .B(n46369), .Z(n46372) );
  XOR U55839 ( .A(n46371), .B(n46372), .Z(n46376) );
  XOR U55840 ( .A(n46375), .B(n46376), .Z(n46379) );
  XOR U55841 ( .A(n46378), .B(n46379), .Z(n46387) );
  IV U55842 ( .A(n43028), .Z(n43031) );
  IV U55843 ( .A(n43029), .Z(n43030) );
  NOR U55844 ( .A(n43031), .B(n43030), .Z(n46385) );
  XOR U55845 ( .A(n46387), .B(n46385), .Z(n46389) );
  XOR U55846 ( .A(n46388), .B(n46389), .Z(n46383) );
  XOR U55847 ( .A(n46382), .B(n46383), .Z(n45786) );
  XOR U55848 ( .A(n45785), .B(n45786), .Z(n43034) );
  IV U55849 ( .A(n43034), .Z(n43032) );
  NOR U55850 ( .A(n43033), .B(n43032), .Z(n46396) );
  IV U55851 ( .A(n43033), .Z(n43035) );
  NOR U55852 ( .A(n43035), .B(n43034), .Z(n49811) );
  NOR U55853 ( .A(n46396), .B(n49811), .Z(n45780) );
  XOR U55854 ( .A(n49283), .B(n45780), .Z(n46403) );
  NOR U55855 ( .A(n43036), .B(n45776), .Z(n43040) );
  IV U55856 ( .A(n43037), .Z(n43039) );
  IV U55857 ( .A(n43038), .Z(n43043) );
  NOR U55858 ( .A(n43039), .B(n43043), .Z(n46402) );
  NOR U55859 ( .A(n43040), .B(n46402), .Z(n43041) );
  XOR U55860 ( .A(n46403), .B(n43041), .Z(n45772) );
  IV U55861 ( .A(n43042), .Z(n43044) );
  NOR U55862 ( .A(n43044), .B(n43043), .Z(n46399) );
  IV U55863 ( .A(n43045), .Z(n43046) );
  NOR U55864 ( .A(n43046), .B(n43052), .Z(n45773) );
  NOR U55865 ( .A(n46399), .B(n45773), .Z(n43047) );
  XOR U55866 ( .A(n45772), .B(n43047), .Z(n45767) );
  XOR U55867 ( .A(n45766), .B(n45767), .Z(n45770) );
  XOR U55868 ( .A(n45769), .B(n45770), .Z(n46410) );
  IV U55869 ( .A(n46410), .Z(n43055) );
  IV U55870 ( .A(n43048), .Z(n43049) );
  NOR U55871 ( .A(n43050), .B(n43049), .Z(n46409) );
  IV U55872 ( .A(n43051), .Z(n43053) );
  NOR U55873 ( .A(n43053), .B(n43052), .Z(n45764) );
  NOR U55874 ( .A(n46409), .B(n45764), .Z(n43054) );
  XOR U55875 ( .A(n43055), .B(n43054), .Z(n46414) );
  IV U55876 ( .A(n43056), .Z(n43058) );
  NOR U55877 ( .A(n43058), .B(n43057), .Z(n46412) );
  XOR U55878 ( .A(n46414), .B(n46412), .Z(n46417) );
  XOR U55879 ( .A(n46415), .B(n46417), .Z(n49257) );
  XOR U55880 ( .A(n45763), .B(n49257), .Z(n46421) );
  IV U55881 ( .A(n43059), .Z(n43061) );
  IV U55882 ( .A(n43060), .Z(n43067) );
  NOR U55883 ( .A(n43061), .B(n43067), .Z(n46430) );
  IV U55884 ( .A(n43062), .Z(n43064) );
  NOR U55885 ( .A(n43064), .B(n43063), .Z(n46425) );
  NOR U55886 ( .A(n46430), .B(n46425), .Z(n46422) );
  XOR U55887 ( .A(n46421), .B(n46422), .Z(n49247) );
  NOR U55888 ( .A(n43065), .B(n49247), .Z(n45762) );
  IV U55889 ( .A(n43066), .Z(n43068) );
  NOR U55890 ( .A(n43068), .B(n43067), .Z(n45760) );
  XOR U55891 ( .A(n49247), .B(n45760), .Z(n45756) );
  IV U55892 ( .A(n45756), .Z(n43069) );
  NOR U55893 ( .A(n43070), .B(n43069), .Z(n43071) );
  NOR U55894 ( .A(n45762), .B(n43071), .Z(n45752) );
  IV U55895 ( .A(n43072), .Z(n45757) );
  NOR U55896 ( .A(n43073), .B(n45757), .Z(n43076) );
  IV U55897 ( .A(n43074), .Z(n43075) );
  NOR U55898 ( .A(n43075), .B(n43079), .Z(n45751) );
  NOR U55899 ( .A(n43076), .B(n45751), .Z(n43077) );
  XOR U55900 ( .A(n45752), .B(n43077), .Z(n45750) );
  IV U55901 ( .A(n43078), .Z(n43080) );
  NOR U55902 ( .A(n43080), .B(n43079), .Z(n45748) );
  XOR U55903 ( .A(n45750), .B(n45748), .Z(n45744) );
  XOR U55904 ( .A(n45743), .B(n45744), .Z(n46443) );
  XOR U55905 ( .A(n45746), .B(n46443), .Z(n46447) );
  XOR U55906 ( .A(n43081), .B(n46447), .Z(n46449) );
  XOR U55907 ( .A(n43082), .B(n46449), .Z(n45740) );
  XOR U55908 ( .A(n45739), .B(n45740), .Z(n46453) );
  XOR U55909 ( .A(n46452), .B(n46453), .Z(n46466) );
  XOR U55910 ( .A(n43083), .B(n46466), .Z(n43084) );
  IV U55911 ( .A(n43084), .Z(n45733) );
  XOR U55912 ( .A(n45731), .B(n45733), .Z(n45736) );
  IV U55913 ( .A(n43085), .Z(n43087) );
  NOR U55914 ( .A(n43087), .B(n43086), .Z(n45734) );
  XOR U55915 ( .A(n45736), .B(n45734), .Z(n46469) );
  XOR U55916 ( .A(n46468), .B(n46469), .Z(n46472) );
  IV U55917 ( .A(n46472), .Z(n43095) );
  IV U55918 ( .A(n43088), .Z(n43089) );
  NOR U55919 ( .A(n43090), .B(n43089), .Z(n46471) );
  IV U55920 ( .A(n43091), .Z(n43093) );
  NOR U55921 ( .A(n43093), .B(n43092), .Z(n45729) );
  NOR U55922 ( .A(n46471), .B(n45729), .Z(n43094) );
  XOR U55923 ( .A(n43095), .B(n43094), .Z(n45724) );
  XOR U55924 ( .A(n45723), .B(n45724), .Z(n45727) );
  XOR U55925 ( .A(n45726), .B(n45727), .Z(n46480) );
  XOR U55926 ( .A(n43096), .B(n46480), .Z(n43103) );
  IV U55927 ( .A(n43103), .Z(n45722) );
  XOR U55928 ( .A(n43097), .B(n45722), .Z(n43106) );
  IV U55929 ( .A(n43106), .Z(n43098) );
  NOR U55930 ( .A(n43099), .B(n43098), .Z(n46485) );
  IV U55931 ( .A(n43100), .Z(n43101) );
  NOR U55932 ( .A(n43101), .B(n49202), .Z(n43107) );
  IV U55933 ( .A(n43107), .Z(n43105) );
  IV U55934 ( .A(n43102), .Z(n45721) );
  XOR U55935 ( .A(n45721), .B(n43103), .Z(n43104) );
  NOR U55936 ( .A(n43105), .B(n43104), .Z(n49904) );
  NOR U55937 ( .A(n43107), .B(n43106), .Z(n43108) );
  NOR U55938 ( .A(n49904), .B(n43108), .Z(n49189) );
  NOR U55939 ( .A(n43109), .B(n49189), .Z(n43110) );
  NOR U55940 ( .A(n46485), .B(n43110), .Z(n43111) );
  IV U55941 ( .A(n43111), .Z(n46484) );
  IV U55942 ( .A(n43112), .Z(n43113) );
  NOR U55943 ( .A(n43113), .B(n49202), .Z(n46482) );
  XOR U55944 ( .A(n46484), .B(n46482), .Z(n46489) );
  XOR U55945 ( .A(n46488), .B(n46489), .Z(n46497) );
  XOR U55946 ( .A(n46498), .B(n46497), .Z(n43114) );
  IV U55947 ( .A(n43114), .Z(n46495) );
  XOR U55948 ( .A(n46494), .B(n46495), .Z(n45715) );
  IV U55949 ( .A(n43115), .Z(n43116) );
  NOR U55950 ( .A(n43116), .B(n46504), .Z(n43117) );
  IV U55951 ( .A(n43117), .Z(n45714) );
  XOR U55952 ( .A(n45715), .B(n45714), .Z(n45716) );
  NOR U55953 ( .A(n43119), .B(n43118), .Z(n46511) );
  IV U55954 ( .A(n43120), .Z(n43122) );
  NOR U55955 ( .A(n43122), .B(n43121), .Z(n45717) );
  NOR U55956 ( .A(n46511), .B(n45717), .Z(n43123) );
  XOR U55957 ( .A(n45716), .B(n43123), .Z(n46510) );
  IV U55958 ( .A(n43124), .Z(n43126) );
  IV U55959 ( .A(n43125), .Z(n45711) );
  NOR U55960 ( .A(n43126), .B(n45711), .Z(n43133) );
  IV U55961 ( .A(n43133), .Z(n43127) );
  NOR U55962 ( .A(n46510), .B(n43127), .Z(n49167) );
  NOR U55963 ( .A(n46508), .B(n43128), .Z(n43129) );
  NOR U55964 ( .A(n43130), .B(n43129), .Z(n43131) );
  XOR U55965 ( .A(n43131), .B(n46510), .Z(n43143) );
  IV U55966 ( .A(n43143), .Z(n43132) );
  NOR U55967 ( .A(n43133), .B(n43132), .Z(n43134) );
  NOR U55968 ( .A(n49167), .B(n43134), .Z(n43144) );
  IV U55969 ( .A(n43144), .Z(n43138) );
  IV U55970 ( .A(n43135), .Z(n43136) );
  NOR U55971 ( .A(n43136), .B(n43153), .Z(n43148) );
  IV U55972 ( .A(n43148), .Z(n43137) );
  NOR U55973 ( .A(n43138), .B(n43137), .Z(n49155) );
  IV U55974 ( .A(n43139), .Z(n43140) );
  NOR U55975 ( .A(n43141), .B(n43140), .Z(n43145) );
  IV U55976 ( .A(n43145), .Z(n43142) );
  NOR U55977 ( .A(n43143), .B(n43142), .Z(n49165) );
  NOR U55978 ( .A(n43145), .B(n43144), .Z(n43146) );
  NOR U55979 ( .A(n49165), .B(n43146), .Z(n43147) );
  NOR U55980 ( .A(n43148), .B(n43147), .Z(n43149) );
  NOR U55981 ( .A(n49155), .B(n43149), .Z(n45707) );
  NOR U55982 ( .A(n43151), .B(n43150), .Z(n46524) );
  IV U55983 ( .A(n43152), .Z(n43154) );
  NOR U55984 ( .A(n43154), .B(n43153), .Z(n45708) );
  NOR U55985 ( .A(n46524), .B(n45708), .Z(n43155) );
  XOR U55986 ( .A(n45707), .B(n43155), .Z(n45704) );
  XOR U55987 ( .A(n45703), .B(n45704), .Z(n46521) );
  XOR U55988 ( .A(n46520), .B(n46521), .Z(n46535) );
  XOR U55989 ( .A(n43156), .B(n46535), .Z(n43157) );
  IV U55990 ( .A(n43157), .Z(n46538) );
  XOR U55991 ( .A(n46536), .B(n46538), .Z(n46540) );
  XOR U55992 ( .A(n45696), .B(n46540), .Z(n45692) );
  XOR U55993 ( .A(n45691), .B(n45692), .Z(n46550) );
  IV U55994 ( .A(n43158), .Z(n43161) );
  IV U55995 ( .A(n43159), .Z(n43160) );
  NOR U55996 ( .A(n43161), .B(n43160), .Z(n46548) );
  XOR U55997 ( .A(n46550), .B(n46548), .Z(n45689) );
  IV U55998 ( .A(n43162), .Z(n43163) );
  NOR U55999 ( .A(n43164), .B(n43163), .Z(n45688) );
  IV U56000 ( .A(n43165), .Z(n43166) );
  NOR U56001 ( .A(n43167), .B(n43166), .Z(n45686) );
  NOR U56002 ( .A(n45688), .B(n45686), .Z(n43168) );
  XOR U56003 ( .A(n45689), .B(n43168), .Z(n46559) );
  XOR U56004 ( .A(n49134), .B(n46559), .Z(n46561) );
  XOR U56005 ( .A(n46560), .B(n46561), .Z(n46567) );
  IV U56006 ( .A(n43169), .Z(n43171) );
  IV U56007 ( .A(n43170), .Z(n43174) );
  NOR U56008 ( .A(n43171), .B(n43174), .Z(n46565) );
  XOR U56009 ( .A(n46567), .B(n46565), .Z(n46572) );
  IV U56010 ( .A(n49937), .Z(n43172) );
  NOR U56011 ( .A(n49936), .B(n43172), .Z(n46571) );
  IV U56012 ( .A(n43173), .Z(n43175) );
  NOR U56013 ( .A(n43175), .B(n43174), .Z(n46568) );
  NOR U56014 ( .A(n46571), .B(n46568), .Z(n43176) );
  XOR U56015 ( .A(n46572), .B(n43176), .Z(n45683) );
  IV U56016 ( .A(n43177), .Z(n49939) );
  NOR U56017 ( .A(n49936), .B(n49939), .Z(n46574) );
  IV U56018 ( .A(n43178), .Z(n43186) );
  NOR U56019 ( .A(n43179), .B(n43186), .Z(n45684) );
  NOR U56020 ( .A(n46574), .B(n45684), .Z(n43180) );
  XOR U56021 ( .A(n45683), .B(n43180), .Z(n46579) );
  IV U56022 ( .A(n43181), .Z(n43183) );
  NOR U56023 ( .A(n43183), .B(n43182), .Z(n46577) );
  XOR U56024 ( .A(n46579), .B(n46577), .Z(n46581) );
  IV U56025 ( .A(n43184), .Z(n43185) );
  NOR U56026 ( .A(n43186), .B(n43185), .Z(n43187) );
  IV U56027 ( .A(n43187), .Z(n46580) );
  XOR U56028 ( .A(n46581), .B(n46580), .Z(n45678) );
  NOR U56029 ( .A(n43189), .B(n43188), .Z(n45680) );
  IV U56030 ( .A(n43190), .Z(n43192) );
  IV U56031 ( .A(n43191), .Z(n43196) );
  NOR U56032 ( .A(n43192), .B(n43196), .Z(n45677) );
  NOR U56033 ( .A(n45680), .B(n45677), .Z(n43193) );
  XOR U56034 ( .A(n45678), .B(n43193), .Z(n45675) );
  NOR U56035 ( .A(n43194), .B(n45675), .Z(n49096) );
  IV U56036 ( .A(n43195), .Z(n43197) );
  NOR U56037 ( .A(n43197), .B(n43196), .Z(n45674) );
  XOR U56038 ( .A(n45674), .B(n45675), .Z(n49106) );
  IV U56039 ( .A(n49106), .Z(n43198) );
  NOR U56040 ( .A(n43199), .B(n43198), .Z(n43200) );
  NOR U56041 ( .A(n49096), .B(n43200), .Z(n46585) );
  IV U56042 ( .A(n43201), .Z(n49105) );
  NOR U56043 ( .A(n49105), .B(n43204), .Z(n43202) );
  IV U56044 ( .A(n43202), .Z(n46586) );
  XOR U56045 ( .A(n46585), .B(n46586), .Z(n46593) );
  IV U56046 ( .A(n43203), .Z(n43205) );
  NOR U56047 ( .A(n43205), .B(n43204), .Z(n46588) );
  XOR U56048 ( .A(n46593), .B(n46588), .Z(n45673) );
  IV U56049 ( .A(n45673), .Z(n43212) );
  IV U56050 ( .A(n43206), .Z(n43214) );
  NOR U56051 ( .A(n43207), .B(n43214), .Z(n46592) );
  IV U56052 ( .A(n43208), .Z(n43210) );
  NOR U56053 ( .A(n43210), .B(n43209), .Z(n45671) );
  NOR U56054 ( .A(n46592), .B(n45671), .Z(n43211) );
  XOR U56055 ( .A(n43212), .B(n43211), .Z(n45670) );
  IV U56056 ( .A(n43213), .Z(n43215) );
  NOR U56057 ( .A(n43215), .B(n43214), .Z(n45668) );
  XOR U56058 ( .A(n45670), .B(n45668), .Z(n46600) );
  XOR U56059 ( .A(n46599), .B(n46600), .Z(n45665) );
  XOR U56060 ( .A(n45664), .B(n45665), .Z(n46597) );
  XOR U56061 ( .A(n46595), .B(n46597), .Z(n45663) );
  IV U56062 ( .A(n43216), .Z(n43218) );
  NOR U56063 ( .A(n43218), .B(n43217), .Z(n43219) );
  IV U56064 ( .A(n43219), .Z(n43226) );
  NOR U56065 ( .A(n45663), .B(n43226), .Z(n49090) );
  IV U56066 ( .A(n43220), .Z(n43222) );
  NOR U56067 ( .A(n43222), .B(n43221), .Z(n45661) );
  XOR U56068 ( .A(n45663), .B(n45661), .Z(n45660) );
  IV U56069 ( .A(n43223), .Z(n43224) );
  NOR U56070 ( .A(n43225), .B(n43224), .Z(n43227) );
  IV U56071 ( .A(n43227), .Z(n45659) );
  XOR U56072 ( .A(n45660), .B(n45659), .Z(n43229) );
  NOR U56073 ( .A(n43227), .B(n43226), .Z(n43228) );
  NOR U56074 ( .A(n43229), .B(n43228), .Z(n43230) );
  NOR U56075 ( .A(n49090), .B(n43230), .Z(n46608) );
  XOR U56076 ( .A(n46609), .B(n46608), .Z(n46616) );
  IV U56077 ( .A(n46616), .Z(n43238) );
  IV U56078 ( .A(n43231), .Z(n43232) );
  NOR U56079 ( .A(n43233), .B(n43232), .Z(n46615) );
  IV U56080 ( .A(n43234), .Z(n43236) );
  NOR U56081 ( .A(n43236), .B(n43235), .Z(n46610) );
  NOR U56082 ( .A(n46615), .B(n46610), .Z(n43237) );
  XOR U56083 ( .A(n43238), .B(n43237), .Z(n45657) );
  XOR U56084 ( .A(n45655), .B(n45657), .Z(n46621) );
  XOR U56085 ( .A(n46620), .B(n46621), .Z(n45653) );
  NOR U56086 ( .A(n43240), .B(n45653), .Z(n45651) );
  IV U56087 ( .A(n43239), .Z(n46632) );
  XOR U56088 ( .A(n45652), .B(n45653), .Z(n46631) );
  XOR U56089 ( .A(n46632), .B(n46631), .Z(n43243) );
  IV U56090 ( .A(n46631), .Z(n43241) );
  NOR U56091 ( .A(n43241), .B(n43240), .Z(n43242) );
  NOR U56092 ( .A(n43243), .B(n43242), .Z(n43244) );
  NOR U56093 ( .A(n45651), .B(n43244), .Z(n43245) );
  IV U56094 ( .A(n43245), .Z(n45649) );
  XOR U56095 ( .A(n45648), .B(n45649), .Z(n45641) );
  IV U56096 ( .A(n45641), .Z(n43253) );
  NOR U56097 ( .A(n43246), .B(n45642), .Z(n43257) );
  IV U56098 ( .A(n43257), .Z(n43247) );
  NOR U56099 ( .A(n43253), .B(n43247), .Z(n43259) );
  IV U56100 ( .A(n43248), .Z(n43249) );
  NOR U56101 ( .A(n43250), .B(n43249), .Z(n43252) );
  IV U56102 ( .A(n43252), .Z(n43251) );
  NOR U56103 ( .A(n43251), .B(n45649), .Z(n50023) );
  NOR U56104 ( .A(n43253), .B(n43252), .Z(n43254) );
  NOR U56105 ( .A(n50023), .B(n43254), .Z(n43255) );
  IV U56106 ( .A(n43255), .Z(n43256) );
  NOR U56107 ( .A(n43257), .B(n43256), .Z(n43258) );
  NOR U56108 ( .A(n43259), .B(n43258), .Z(n45638) );
  XOR U56109 ( .A(n45637), .B(n45638), .Z(n45633) );
  XOR U56110 ( .A(n45632), .B(n45633), .Z(n46638) );
  IV U56111 ( .A(n46638), .Z(n43267) );
  IV U56112 ( .A(n43260), .Z(n43262) );
  NOR U56113 ( .A(n43262), .B(n43261), .Z(n46636) );
  IV U56114 ( .A(n43263), .Z(n43265) );
  NOR U56115 ( .A(n43265), .B(n43264), .Z(n45635) );
  NOR U56116 ( .A(n46636), .B(n45635), .Z(n43266) );
  XOR U56117 ( .A(n43267), .B(n43266), .Z(n46641) );
  IV U56118 ( .A(n43268), .Z(n43270) );
  NOR U56119 ( .A(n43270), .B(n43269), .Z(n46639) );
  XOR U56120 ( .A(n46641), .B(n46639), .Z(n46643) );
  XOR U56121 ( .A(n46642), .B(n46643), .Z(n45629) );
  XOR U56122 ( .A(n45628), .B(n45629), .Z(n46656) );
  XOR U56123 ( .A(n46655), .B(n46656), .Z(n46652) );
  XOR U56124 ( .A(n43271), .B(n46652), .Z(n43272) );
  IV U56125 ( .A(n43272), .Z(n46668) );
  XOR U56126 ( .A(n46666), .B(n46668), .Z(n46670) );
  IV U56127 ( .A(n46670), .Z(n43274) );
  NOR U56128 ( .A(n46669), .B(n45626), .Z(n43273) );
  XOR U56129 ( .A(n43274), .B(n43273), .Z(n45625) );
  XOR U56130 ( .A(n45623), .B(n45625), .Z(n45619) );
  XOR U56131 ( .A(n45618), .B(n45619), .Z(n49060) );
  XOR U56132 ( .A(n45621), .B(n49060), .Z(n43275) );
  IV U56133 ( .A(n43275), .Z(n49046) );
  IV U56134 ( .A(n43276), .Z(n43277) );
  NOR U56135 ( .A(n43277), .B(n43280), .Z(n49055) );
  IV U56136 ( .A(n43278), .Z(n43279) );
  NOR U56137 ( .A(n43280), .B(n43279), .Z(n49045) );
  NOR U56138 ( .A(n49055), .B(n49045), .Z(n45617) );
  XOR U56139 ( .A(n49046), .B(n45617), .Z(n43290) );
  IV U56140 ( .A(n43290), .Z(n43305) );
  IV U56141 ( .A(n43281), .Z(n43284) );
  NOR U56142 ( .A(n43282), .B(n43297), .Z(n43283) );
  IV U56143 ( .A(n43283), .Z(n43302) );
  NOR U56144 ( .A(n43284), .B(n43302), .Z(n43294) );
  IV U56145 ( .A(n43294), .Z(n43285) );
  NOR U56146 ( .A(n43305), .B(n43285), .Z(n49052) );
  IV U56147 ( .A(n43286), .Z(n43287) );
  NOR U56148 ( .A(n43288), .B(n43287), .Z(n43291) );
  IV U56149 ( .A(n43291), .Z(n43289) );
  NOR U56150 ( .A(n43289), .B(n49046), .Z(n49049) );
  NOR U56151 ( .A(n43291), .B(n43290), .Z(n43292) );
  NOR U56152 ( .A(n49049), .B(n43292), .Z(n43293) );
  NOR U56153 ( .A(n43294), .B(n43293), .Z(n43295) );
  NOR U56154 ( .A(n49052), .B(n43295), .Z(n43307) );
  IV U56155 ( .A(n43307), .Z(n43300) );
  IV U56156 ( .A(n43296), .Z(n43298) );
  NOR U56157 ( .A(n43298), .B(n43297), .Z(n43309) );
  IV U56158 ( .A(n43309), .Z(n43299) );
  NOR U56159 ( .A(n43300), .B(n43299), .Z(n49040) );
  IV U56160 ( .A(n43301), .Z(n43303) );
  NOR U56161 ( .A(n43303), .B(n43302), .Z(n43306) );
  IV U56162 ( .A(n43306), .Z(n43304) );
  NOR U56163 ( .A(n43305), .B(n43304), .Z(n49043) );
  NOR U56164 ( .A(n43307), .B(n43306), .Z(n43308) );
  NOR U56165 ( .A(n49043), .B(n43308), .Z(n43314) );
  NOR U56166 ( .A(n43309), .B(n43314), .Z(n43310) );
  NOR U56167 ( .A(n49040), .B(n43310), .Z(n43311) );
  IV U56168 ( .A(n43311), .Z(n45613) );
  XOR U56169 ( .A(n45614), .B(n45613), .Z(n43312) );
  NOR U56170 ( .A(n43313), .B(n43312), .Z(n43317) );
  IV U56171 ( .A(n43313), .Z(n43316) );
  IV U56172 ( .A(n43314), .Z(n43315) );
  NOR U56173 ( .A(n43316), .B(n43315), .Z(n49036) );
  NOR U56174 ( .A(n43317), .B(n49036), .Z(n45609) );
  IV U56175 ( .A(n43318), .Z(n43320) );
  IV U56176 ( .A(n43319), .Z(n43322) );
  NOR U56177 ( .A(n43320), .B(n43322), .Z(n46686) );
  IV U56178 ( .A(n43321), .Z(n43323) );
  NOR U56179 ( .A(n43323), .B(n43322), .Z(n45608) );
  NOR U56180 ( .A(n45611), .B(n45608), .Z(n43324) );
  IV U56181 ( .A(n43324), .Z(n43325) );
  NOR U56182 ( .A(n46686), .B(n43325), .Z(n43326) );
  XOR U56183 ( .A(n45609), .B(n43326), .Z(n46685) );
  IV U56184 ( .A(n43327), .Z(n43330) );
  IV U56185 ( .A(n43328), .Z(n43329) );
  NOR U56186 ( .A(n43330), .B(n43329), .Z(n46683) );
  XOR U56187 ( .A(n46685), .B(n46683), .Z(n50100) );
  XOR U56188 ( .A(n43331), .B(n50100), .Z(n43332) );
  IV U56189 ( .A(n43332), .Z(n45601) );
  XOR U56190 ( .A(n45599), .B(n45601), .Z(n45603) );
  IV U56191 ( .A(n45603), .Z(n43337) );
  IV U56192 ( .A(n43333), .Z(n43334) );
  NOR U56193 ( .A(n43335), .B(n43334), .Z(n45602) );
  NOR U56194 ( .A(n45602), .B(n45597), .Z(n43336) );
  XOR U56195 ( .A(n43337), .B(n43336), .Z(n46694) );
  XOR U56196 ( .A(n46693), .B(n46694), .Z(n46697) );
  XOR U56197 ( .A(n46696), .B(n46697), .Z(n43338) );
  NOR U56198 ( .A(n43345), .B(n43338), .Z(n49010) );
  NOR U56199 ( .A(n43339), .B(n45594), .Z(n43340) );
  NOR U56200 ( .A(n46696), .B(n43340), .Z(n43341) );
  XOR U56201 ( .A(n43341), .B(n46697), .Z(n43342) );
  IV U56202 ( .A(n43342), .Z(n45589) );
  IV U56203 ( .A(n43343), .Z(n43344) );
  NOR U56204 ( .A(n43355), .B(n43344), .Z(n43346) );
  IV U56205 ( .A(n43346), .Z(n45588) );
  XOR U56206 ( .A(n45589), .B(n45588), .Z(n43348) );
  NOR U56207 ( .A(n43346), .B(n43345), .Z(n43347) );
  NOR U56208 ( .A(n43348), .B(n43347), .Z(n43349) );
  NOR U56209 ( .A(n49010), .B(n43349), .Z(n43350) );
  IV U56210 ( .A(n43350), .Z(n45592) );
  IV U56211 ( .A(n43351), .Z(n43352) );
  NOR U56212 ( .A(n43366), .B(n43352), .Z(n45586) );
  IV U56213 ( .A(n43353), .Z(n43354) );
  NOR U56214 ( .A(n43355), .B(n43354), .Z(n45590) );
  NOR U56215 ( .A(n45586), .B(n45590), .Z(n43356) );
  XOR U56216 ( .A(n45592), .B(n43356), .Z(n43362) );
  IV U56217 ( .A(n43362), .Z(n43361) );
  IV U56218 ( .A(n43357), .Z(n43358) );
  NOR U56219 ( .A(n43359), .B(n43358), .Z(n43363) );
  IV U56220 ( .A(n43363), .Z(n43360) );
  NOR U56221 ( .A(n43361), .B(n43360), .Z(n50141) );
  NOR U56222 ( .A(n43363), .B(n43362), .Z(n45585) );
  IV U56223 ( .A(n43364), .Z(n43365) );
  NOR U56224 ( .A(n43366), .B(n43365), .Z(n45583) );
  XOR U56225 ( .A(n45585), .B(n45583), .Z(n43367) );
  NOR U56226 ( .A(n50141), .B(n43367), .Z(n43368) );
  IV U56227 ( .A(n43368), .Z(n46713) );
  IV U56228 ( .A(n43369), .Z(n43370) );
  NOR U56229 ( .A(n43371), .B(n43370), .Z(n46711) );
  XOR U56230 ( .A(n46713), .B(n46711), .Z(n46707) );
  XOR U56231 ( .A(n46708), .B(n46707), .Z(n43374) );
  IV U56232 ( .A(n43374), .Z(n43372) );
  NOR U56233 ( .A(n43373), .B(n43372), .Z(n46722) );
  NOR U56234 ( .A(n43375), .B(n43374), .Z(n46726) );
  XOR U56235 ( .A(n46726), .B(n46724), .Z(n43376) );
  NOR U56236 ( .A(n46722), .B(n43376), .Z(n43377) );
  IV U56237 ( .A(n43377), .Z(n46728) );
  XOR U56238 ( .A(n46727), .B(n46728), .Z(n46732) );
  XOR U56239 ( .A(n46731), .B(n46732), .Z(n46736) );
  IV U56240 ( .A(n43378), .Z(n43382) );
  NOR U56241 ( .A(n43380), .B(n43379), .Z(n43381) );
  IV U56242 ( .A(n43381), .Z(n43384) );
  NOR U56243 ( .A(n43382), .B(n43384), .Z(n46734) );
  XOR U56244 ( .A(n46736), .B(n46734), .Z(n45579) );
  IV U56245 ( .A(n43383), .Z(n43385) );
  NOR U56246 ( .A(n43385), .B(n43384), .Z(n45577) );
  XOR U56247 ( .A(n45579), .B(n45577), .Z(n45582) );
  IV U56248 ( .A(n45582), .Z(n43392) );
  NOR U56249 ( .A(n43387), .B(n43386), .Z(n45575) );
  IV U56250 ( .A(n43388), .Z(n43390) );
  NOR U56251 ( .A(n43390), .B(n43389), .Z(n45580) );
  NOR U56252 ( .A(n45575), .B(n45580), .Z(n43391) );
  XOR U56253 ( .A(n43392), .B(n43391), .Z(n46743) );
  XOR U56254 ( .A(n46741), .B(n46743), .Z(n46746) );
  XOR U56255 ( .A(n43393), .B(n46746), .Z(n43394) );
  IV U56256 ( .A(n43394), .Z(n45570) );
  XOR U56257 ( .A(n43395), .B(n45570), .Z(n46754) );
  XOR U56258 ( .A(n46752), .B(n46754), .Z(n46760) );
  IV U56259 ( .A(n46760), .Z(n43402) );
  NOR U56260 ( .A(n43397), .B(n43396), .Z(n46755) );
  IV U56261 ( .A(n43398), .Z(n43400) );
  IV U56262 ( .A(n43399), .Z(n43403) );
  NOR U56263 ( .A(n43400), .B(n43403), .Z(n46758) );
  NOR U56264 ( .A(n46755), .B(n46758), .Z(n43401) );
  XOR U56265 ( .A(n43402), .B(n43401), .Z(n46764) );
  NOR U56266 ( .A(n43404), .B(n43403), .Z(n43405) );
  IV U56267 ( .A(n43405), .Z(n43406) );
  NOR U56268 ( .A(n43407), .B(n43406), .Z(n46762) );
  XOR U56269 ( .A(n46764), .B(n46762), .Z(n46772) );
  XOR U56270 ( .A(n43408), .B(n46772), .Z(n45563) );
  XOR U56271 ( .A(n43409), .B(n45563), .Z(n45558) );
  XOR U56272 ( .A(n45557), .B(n45558), .Z(n45562) );
  XOR U56273 ( .A(n45560), .B(n45562), .Z(n45549) );
  XOR U56274 ( .A(n45547), .B(n45549), .Z(n45552) );
  XOR U56275 ( .A(n45550), .B(n45552), .Z(n45555) );
  XOR U56276 ( .A(n45553), .B(n45555), .Z(n46780) );
  NOR U56277 ( .A(n43417), .B(n46780), .Z(n50213) );
  IV U56278 ( .A(n43410), .Z(n43412) );
  NOR U56279 ( .A(n43412), .B(n43411), .Z(n43413) );
  IV U56280 ( .A(n43413), .Z(n46784) );
  IV U56281 ( .A(n43414), .Z(n43415) );
  NOR U56282 ( .A(n43416), .B(n43415), .Z(n46779) );
  XOR U56283 ( .A(n46779), .B(n46780), .Z(n46783) );
  XOR U56284 ( .A(n46784), .B(n46783), .Z(n43420) );
  IV U56285 ( .A(n46783), .Z(n43418) );
  NOR U56286 ( .A(n43418), .B(n43417), .Z(n43419) );
  NOR U56287 ( .A(n43420), .B(n43419), .Z(n43421) );
  NOR U56288 ( .A(n50213), .B(n43421), .Z(n46786) );
  IV U56289 ( .A(n43422), .Z(n43423) );
  NOR U56290 ( .A(n43424), .B(n43423), .Z(n46788) );
  IV U56291 ( .A(n43425), .Z(n43427) );
  NOR U56292 ( .A(n43427), .B(n43426), .Z(n46785) );
  NOR U56293 ( .A(n46788), .B(n46785), .Z(n43428) );
  XOR U56294 ( .A(n46786), .B(n43428), .Z(n48971) );
  XOR U56295 ( .A(n46797), .B(n48971), .Z(n43429) );
  IV U56296 ( .A(n43429), .Z(n45544) );
  XOR U56297 ( .A(n45543), .B(n45544), .Z(n46794) );
  XOR U56298 ( .A(n46793), .B(n46794), .Z(n46805) );
  IV U56299 ( .A(n43430), .Z(n43432) );
  NOR U56300 ( .A(n43432), .B(n43431), .Z(n46803) );
  XOR U56301 ( .A(n46805), .B(n46803), .Z(n46808) );
  NOR U56302 ( .A(n43434), .B(n43433), .Z(n43435) );
  IV U56303 ( .A(n43435), .Z(n43436) );
  NOR U56304 ( .A(n43437), .B(n43436), .Z(n46806) );
  XOR U56305 ( .A(n46808), .B(n46806), .Z(n46812) );
  IV U56306 ( .A(n43438), .Z(n43439) );
  NOR U56307 ( .A(n43440), .B(n43439), .Z(n45542) );
  IV U56308 ( .A(n43441), .Z(n43442) );
  NOR U56309 ( .A(n43442), .B(n45536), .Z(n46818) );
  NOR U56310 ( .A(n45542), .B(n46818), .Z(n46813) );
  XOR U56311 ( .A(n46812), .B(n46813), .Z(n43443) );
  IV U56312 ( .A(n43443), .Z(n46836) );
  XOR U56313 ( .A(n43444), .B(n46836), .Z(n46830) );
  XOR U56314 ( .A(n43445), .B(n46830), .Z(n46845) );
  XOR U56315 ( .A(n43446), .B(n46845), .Z(n45529) );
  XOR U56316 ( .A(n43447), .B(n45529), .Z(n45526) );
  XOR U56317 ( .A(n43448), .B(n45526), .Z(n45518) );
  IV U56318 ( .A(n43449), .Z(n43451) );
  NOR U56319 ( .A(n43451), .B(n43450), .Z(n43452) );
  IV U56320 ( .A(n43452), .Z(n45519) );
  XOR U56321 ( .A(n45518), .B(n45519), .Z(n48948) );
  XOR U56322 ( .A(n45521), .B(n48948), .Z(n46856) );
  XOR U56323 ( .A(n46857), .B(n46856), .Z(n45514) );
  XOR U56324 ( .A(n45515), .B(n45514), .Z(n46853) );
  XOR U56325 ( .A(n46854), .B(n46853), .Z(n43459) );
  IV U56326 ( .A(n43459), .Z(n43453) );
  NOR U56327 ( .A(n43454), .B(n43453), .Z(n50264) );
  IV U56328 ( .A(n43455), .Z(n43456) );
  NOR U56329 ( .A(n43457), .B(n43456), .Z(n43460) );
  IV U56330 ( .A(n43460), .Z(n43458) );
  NOR U56331 ( .A(n43458), .B(n46853), .Z(n50259) );
  NOR U56332 ( .A(n43460), .B(n43459), .Z(n43461) );
  NOR U56333 ( .A(n50259), .B(n43461), .Z(n43462) );
  NOR U56334 ( .A(n43463), .B(n43462), .Z(n43464) );
  NOR U56335 ( .A(n50264), .B(n43464), .Z(n45511) );
  IV U56336 ( .A(n43465), .Z(n43467) );
  NOR U56337 ( .A(n43467), .B(n43466), .Z(n46864) );
  IV U56338 ( .A(n43468), .Z(n43473) );
  NOR U56339 ( .A(n43470), .B(n43469), .Z(n43471) );
  IV U56340 ( .A(n43471), .Z(n43472) );
  NOR U56341 ( .A(n43473), .B(n43472), .Z(n45512) );
  NOR U56342 ( .A(n46864), .B(n45512), .Z(n43474) );
  XOR U56343 ( .A(n45511), .B(n43474), .Z(n46875) );
  XOR U56344 ( .A(n46873), .B(n46875), .Z(n45508) );
  XOR U56345 ( .A(n45507), .B(n45508), .Z(n46870) );
  XOR U56346 ( .A(n43475), .B(n46870), .Z(n43483) );
  IV U56347 ( .A(n43483), .Z(n43476) );
  NOR U56348 ( .A(n43482), .B(n43476), .Z(n50275) );
  IV U56349 ( .A(n43480), .Z(n43478) );
  XOR U56350 ( .A(n46869), .B(n46870), .Z(n43477) );
  NOR U56351 ( .A(n43478), .B(n43477), .Z(n50271) );
  NOR U56352 ( .A(n50275), .B(n50271), .Z(n43479) );
  IV U56353 ( .A(n43479), .Z(n46882) );
  NOR U56354 ( .A(n43480), .B(n43483), .Z(n43481) );
  NOR U56355 ( .A(n46882), .B(n43481), .Z(n43485) );
  NOR U56356 ( .A(n43483), .B(n43482), .Z(n43484) );
  NOR U56357 ( .A(n43485), .B(n43484), .Z(n45501) );
  XOR U56358 ( .A(n45499), .B(n45501), .Z(n45503) );
  XOR U56359 ( .A(n45502), .B(n45503), .Z(n45494) );
  XOR U56360 ( .A(n45493), .B(n45494), .Z(n45498) );
  XOR U56361 ( .A(n45496), .B(n45498), .Z(n45489) );
  XOR U56362 ( .A(n45487), .B(n45489), .Z(n45492) );
  XOR U56363 ( .A(n45490), .B(n45492), .Z(n46885) );
  XOR U56364 ( .A(n46884), .B(n46885), .Z(n46891) );
  XOR U56365 ( .A(n43486), .B(n46891), .Z(n43487) );
  IV U56366 ( .A(n43487), .Z(n46894) );
  XOR U56367 ( .A(n46893), .B(n46894), .Z(n50315) );
  XOR U56368 ( .A(n45483), .B(n50315), .Z(n45481) );
  XOR U56369 ( .A(n45484), .B(n45481), .Z(n45478) );
  XOR U56370 ( .A(n43488), .B(n45478), .Z(n45466) );
  XOR U56371 ( .A(n43489), .B(n45466), .Z(n45470) );
  XOR U56372 ( .A(n43490), .B(n45470), .Z(n43498) );
  NOR U56373 ( .A(n43505), .B(n43498), .Z(n48911) );
  IV U56374 ( .A(n43491), .Z(n43493) );
  NOR U56375 ( .A(n43493), .B(n43492), .Z(n43507) );
  IV U56376 ( .A(n43507), .Z(n43503) );
  IV U56377 ( .A(n43494), .Z(n43496) );
  NOR U56378 ( .A(n43496), .B(n43495), .Z(n43500) );
  IV U56379 ( .A(n43500), .Z(n43497) );
  NOR U56380 ( .A(n43497), .B(n45470), .Z(n48907) );
  IV U56381 ( .A(n43498), .Z(n43499) );
  NOR U56382 ( .A(n43500), .B(n43499), .Z(n43501) );
  NOR U56383 ( .A(n48907), .B(n43501), .Z(n43506) );
  IV U56384 ( .A(n43506), .Z(n43502) );
  NOR U56385 ( .A(n43503), .B(n43502), .Z(n48904) );
  NOR U56386 ( .A(n48911), .B(n48904), .Z(n43504) );
  IV U56387 ( .A(n43504), .Z(n46907) );
  NOR U56388 ( .A(n46907), .B(n43505), .Z(n43510) );
  NOR U56389 ( .A(n43507), .B(n43506), .Z(n43508) );
  NOR U56390 ( .A(n43508), .B(n46907), .Z(n43509) );
  NOR U56391 ( .A(n43510), .B(n43509), .Z(n45464) );
  XOR U56392 ( .A(n45462), .B(n45464), .Z(n46909) );
  XOR U56393 ( .A(n43511), .B(n46909), .Z(n45453) );
  IV U56394 ( .A(n43512), .Z(n43513) );
  NOR U56395 ( .A(n43514), .B(n43513), .Z(n50349) );
  IV U56396 ( .A(n43515), .Z(n43516) );
  NOR U56397 ( .A(n43517), .B(n43516), .Z(n50340) );
  NOR U56398 ( .A(n50349), .B(n50340), .Z(n45454) );
  XOR U56399 ( .A(n45453), .B(n45454), .Z(n45456) );
  XOR U56400 ( .A(n43518), .B(n45456), .Z(n43519) );
  IV U56401 ( .A(n43519), .Z(n45448) );
  XOR U56402 ( .A(n45446), .B(n45448), .Z(n46922) );
  IV U56403 ( .A(n46922), .Z(n43526) );
  IV U56404 ( .A(n43520), .Z(n43521) );
  NOR U56405 ( .A(n43528), .B(n43521), .Z(n46921) );
  IV U56406 ( .A(n43522), .Z(n43523) );
  NOR U56407 ( .A(n43524), .B(n43523), .Z(n45449) );
  NOR U56408 ( .A(n46921), .B(n45449), .Z(n43525) );
  XOR U56409 ( .A(n43526), .B(n43525), .Z(n45444) );
  IV U56410 ( .A(n43527), .Z(n43529) );
  NOR U56411 ( .A(n43529), .B(n43528), .Z(n43530) );
  IV U56412 ( .A(n43530), .Z(n43531) );
  NOR U56413 ( .A(n43532), .B(n43531), .Z(n45442) );
  XOR U56414 ( .A(n45444), .B(n45442), .Z(n46930) );
  XOR U56415 ( .A(n46929), .B(n46930), .Z(n48884) );
  XOR U56416 ( .A(n46932), .B(n48884), .Z(n46935) );
  XOR U56417 ( .A(n46936), .B(n46935), .Z(n43540) );
  IV U56418 ( .A(n43540), .Z(n43533) );
  NOR U56419 ( .A(n43543), .B(n43533), .Z(n50366) );
  IV U56420 ( .A(n43534), .Z(n43535) );
  NOR U56421 ( .A(n43536), .B(n43535), .Z(n43537) );
  IV U56422 ( .A(n43537), .Z(n46940) );
  NOR U56423 ( .A(n43538), .B(n48887), .Z(n43541) );
  IV U56424 ( .A(n43541), .Z(n43539) );
  NOR U56425 ( .A(n43539), .B(n48884), .Z(n46937) );
  NOR U56426 ( .A(n43541), .B(n43540), .Z(n43542) );
  NOR U56427 ( .A(n46937), .B(n43542), .Z(n43544) );
  IV U56428 ( .A(n43544), .Z(n46939) );
  XOR U56429 ( .A(n46940), .B(n46939), .Z(n43546) );
  NOR U56430 ( .A(n43544), .B(n43543), .Z(n43545) );
  NOR U56431 ( .A(n43546), .B(n43545), .Z(n43547) );
  NOR U56432 ( .A(n50366), .B(n43547), .Z(n43548) );
  IV U56433 ( .A(n43548), .Z(n46942) );
  NOR U56434 ( .A(n43555), .B(n46942), .Z(n48878) );
  IV U56435 ( .A(n43549), .Z(n43550) );
  NOR U56436 ( .A(n43551), .B(n43550), .Z(n43552) );
  IV U56437 ( .A(n43552), .Z(n45441) );
  NOR U56438 ( .A(n43553), .B(n46943), .Z(n43554) );
  XOR U56439 ( .A(n43554), .B(n46942), .Z(n45440) );
  XOR U56440 ( .A(n45441), .B(n45440), .Z(n43558) );
  IV U56441 ( .A(n45440), .Z(n43556) );
  NOR U56442 ( .A(n43556), .B(n43555), .Z(n43557) );
  NOR U56443 ( .A(n43558), .B(n43557), .Z(n43559) );
  NOR U56444 ( .A(n48878), .B(n43559), .Z(n43560) );
  IV U56445 ( .A(n43560), .Z(n46955) );
  XOR U56446 ( .A(n45435), .B(n46955), .Z(n45438) );
  IV U56447 ( .A(n43561), .Z(n43563) );
  NOR U56448 ( .A(n43563), .B(n43562), .Z(n46954) );
  NOR U56449 ( .A(n45437), .B(n46954), .Z(n43564) );
  XOR U56450 ( .A(n45438), .B(n43564), .Z(n46951) );
  IV U56451 ( .A(n43565), .Z(n43566) );
  NOR U56452 ( .A(n43567), .B(n43566), .Z(n46952) );
  IV U56453 ( .A(n43568), .Z(n43570) );
  NOR U56454 ( .A(n43570), .B(n43569), .Z(n46961) );
  NOR U56455 ( .A(n46952), .B(n46961), .Z(n43571) );
  XOR U56456 ( .A(n46951), .B(n43571), .Z(n46960) );
  IV U56457 ( .A(n43572), .Z(n43573) );
  NOR U56458 ( .A(n43573), .B(n43576), .Z(n46958) );
  XOR U56459 ( .A(n46960), .B(n46958), .Z(n46967) );
  IV U56460 ( .A(n43574), .Z(n43575) );
  NOR U56461 ( .A(n43576), .B(n43575), .Z(n46965) );
  XOR U56462 ( .A(n46967), .B(n46965), .Z(n48870) );
  IV U56463 ( .A(n48870), .Z(n43583) );
  IV U56464 ( .A(n43577), .Z(n43578) );
  NOR U56465 ( .A(n43579), .B(n43578), .Z(n50418) );
  IV U56466 ( .A(n43580), .Z(n43582) );
  NOR U56467 ( .A(n43582), .B(n43581), .Z(n48868) );
  NOR U56468 ( .A(n50418), .B(n48868), .Z(n46968) );
  XOR U56469 ( .A(n43583), .B(n46968), .Z(n45432) );
  XOR U56470 ( .A(n45431), .B(n45432), .Z(n46974) );
  XOR U56471 ( .A(n46973), .B(n46974), .Z(n45429) );
  XOR U56472 ( .A(n45428), .B(n45429), .Z(n46985) );
  XOR U56473 ( .A(n46983), .B(n46985), .Z(n46988) );
  NOR U56474 ( .A(n43590), .B(n46988), .Z(n50437) );
  IV U56475 ( .A(n43584), .Z(n43589) );
  IV U56476 ( .A(n43585), .Z(n43586) );
  NOR U56477 ( .A(n43589), .B(n43586), .Z(n46986) );
  XOR U56478 ( .A(n46988), .B(n46986), .Z(n45426) );
  IV U56479 ( .A(n43587), .Z(n43588) );
  NOR U56480 ( .A(n43589), .B(n43588), .Z(n43591) );
  IV U56481 ( .A(n43591), .Z(n45425) );
  XOR U56482 ( .A(n45426), .B(n45425), .Z(n43593) );
  NOR U56483 ( .A(n43591), .B(n43590), .Z(n43592) );
  NOR U56484 ( .A(n43593), .B(n43592), .Z(n43594) );
  NOR U56485 ( .A(n50437), .B(n43594), .Z(n43595) );
  IV U56486 ( .A(n43595), .Z(n46991) );
  XOR U56487 ( .A(n46989), .B(n46991), .Z(n43596) );
  XOR U56488 ( .A(n43597), .B(n43596), .Z(n46997) );
  IV U56489 ( .A(n43598), .Z(n43600) );
  NOR U56490 ( .A(n43600), .B(n43599), .Z(n46995) );
  XOR U56491 ( .A(n46997), .B(n46995), .Z(n48856) );
  XOR U56492 ( .A(n46998), .B(n48856), .Z(n47006) );
  IV U56493 ( .A(n43601), .Z(n43602) );
  NOR U56494 ( .A(n43609), .B(n43602), .Z(n47015) );
  IV U56495 ( .A(n43603), .Z(n43605) );
  NOR U56496 ( .A(n43605), .B(n43604), .Z(n47007) );
  NOR U56497 ( .A(n47015), .B(n47007), .Z(n43606) );
  XOR U56498 ( .A(n47006), .B(n43606), .Z(n47003) );
  IV U56499 ( .A(n43607), .Z(n43608) );
  NOR U56500 ( .A(n43609), .B(n43608), .Z(n47001) );
  XOR U56501 ( .A(n47003), .B(n47001), .Z(n47025) );
  XOR U56502 ( .A(n47023), .B(n47025), .Z(n45416) );
  XOR U56503 ( .A(n43610), .B(n45416), .Z(n43611) );
  IV U56504 ( .A(n43611), .Z(n45412) );
  XOR U56505 ( .A(n45410), .B(n45412), .Z(n47033) );
  IV U56506 ( .A(n47033), .Z(n43616) );
  IV U56507 ( .A(n43612), .Z(n43614) );
  IV U56508 ( .A(n43613), .Z(n43617) );
  NOR U56509 ( .A(n43614), .B(n43617), .Z(n47031) );
  NOR U56510 ( .A(n45408), .B(n47031), .Z(n43615) );
  XOR U56511 ( .A(n43616), .B(n43615), .Z(n47030) );
  NOR U56512 ( .A(n43618), .B(n43617), .Z(n43619) );
  IV U56513 ( .A(n43619), .Z(n43620) );
  NOR U56514 ( .A(n43621), .B(n43620), .Z(n47028) );
  XOR U56515 ( .A(n47030), .B(n47028), .Z(n45404) );
  XOR U56516 ( .A(n45402), .B(n45404), .Z(n45407) );
  XOR U56517 ( .A(n45405), .B(n45407), .Z(n47037) );
  XOR U56518 ( .A(n43622), .B(n47037), .Z(n43623) );
  IV U56519 ( .A(n43623), .Z(n47043) );
  XOR U56520 ( .A(n47039), .B(n47043), .Z(n45398) );
  IV U56521 ( .A(n43624), .Z(n43626) );
  NOR U56522 ( .A(n43626), .B(n43625), .Z(n47041) );
  IV U56523 ( .A(n43633), .Z(n43627) );
  NOR U56524 ( .A(n43627), .B(n43632), .Z(n45397) );
  NOR U56525 ( .A(n47041), .B(n45397), .Z(n43628) );
  XOR U56526 ( .A(n45398), .B(n43628), .Z(n45394) );
  IV U56527 ( .A(n43629), .Z(n43630) );
  NOR U56528 ( .A(n43630), .B(n43632), .Z(n45395) );
  IV U56529 ( .A(n43631), .Z(n43635) );
  XOR U56530 ( .A(n43633), .B(n43632), .Z(n43634) );
  NOR U56531 ( .A(n43635), .B(n43634), .Z(n47045) );
  NOR U56532 ( .A(n45395), .B(n47045), .Z(n43636) );
  XOR U56533 ( .A(n45394), .B(n43636), .Z(n47049) );
  IV U56534 ( .A(n43637), .Z(n43638) );
  NOR U56535 ( .A(n43639), .B(n43638), .Z(n45392) );
  IV U56536 ( .A(n43640), .Z(n43643) );
  IV U56537 ( .A(n43641), .Z(n43642) );
  NOR U56538 ( .A(n43643), .B(n43642), .Z(n47048) );
  NOR U56539 ( .A(n45392), .B(n47048), .Z(n43644) );
  XOR U56540 ( .A(n47049), .B(n43644), .Z(n47051) );
  XOR U56541 ( .A(n47052), .B(n47051), .Z(n47055) );
  XOR U56542 ( .A(n47054), .B(n47055), .Z(n45387) );
  XOR U56543 ( .A(n43645), .B(n45387), .Z(n43646) );
  IV U56544 ( .A(n43646), .Z(n47061) );
  XOR U56545 ( .A(n47059), .B(n47061), .Z(n50485) );
  IV U56546 ( .A(n50485), .Z(n43653) );
  IV U56547 ( .A(n43647), .Z(n43649) );
  NOR U56548 ( .A(n43649), .B(n43648), .Z(n50483) );
  IV U56549 ( .A(n43650), .Z(n43651) );
  NOR U56550 ( .A(n43652), .B(n43651), .Z(n50496) );
  NOR U56551 ( .A(n50483), .B(n50496), .Z(n47062) );
  XOR U56552 ( .A(n43653), .B(n47062), .Z(n45378) );
  XOR U56553 ( .A(n45377), .B(n45378), .Z(n45381) );
  XOR U56554 ( .A(n45380), .B(n45381), .Z(n45373) );
  XOR U56555 ( .A(n45371), .B(n45373), .Z(n45376) );
  XOR U56556 ( .A(n45374), .B(n45376), .Z(n52483) );
  XOR U56557 ( .A(n45370), .B(n52483), .Z(n43667) );
  IV U56558 ( .A(n43667), .Z(n45368) );
  IV U56559 ( .A(n43654), .Z(n43655) );
  NOR U56560 ( .A(n43656), .B(n43655), .Z(n45365) );
  IV U56561 ( .A(n43657), .Z(n43659) );
  NOR U56562 ( .A(n43659), .B(n43658), .Z(n43666) );
  NOR U56563 ( .A(n45365), .B(n43666), .Z(n43660) );
  XOR U56564 ( .A(n45368), .B(n43660), .Z(n43670) );
  IV U56565 ( .A(n43670), .Z(n43661) );
  NOR U56566 ( .A(n43662), .B(n43661), .Z(n48788) );
  IV U56567 ( .A(n43663), .Z(n43665) );
  NOR U56568 ( .A(n43665), .B(n43664), .Z(n43671) );
  IV U56569 ( .A(n43671), .Z(n43669) );
  IV U56570 ( .A(n43666), .Z(n45367) );
  XOR U56571 ( .A(n45367), .B(n43667), .Z(n43668) );
  NOR U56572 ( .A(n43669), .B(n43668), .Z(n50519) );
  NOR U56573 ( .A(n43671), .B(n43670), .Z(n43672) );
  NOR U56574 ( .A(n50519), .B(n43672), .Z(n43673) );
  NOR U56575 ( .A(n43674), .B(n43673), .Z(n43675) );
  NOR U56576 ( .A(n48788), .B(n43675), .Z(n43676) );
  IV U56577 ( .A(n43676), .Z(n47069) );
  XOR U56578 ( .A(n47068), .B(n47069), .Z(n47072) );
  IV U56579 ( .A(n47072), .Z(n43684) );
  IV U56580 ( .A(n43677), .Z(n43679) );
  NOR U56581 ( .A(n43679), .B(n43678), .Z(n47071) );
  IV U56582 ( .A(n43680), .Z(n43682) );
  NOR U56583 ( .A(n43682), .B(n43681), .Z(n45363) );
  NOR U56584 ( .A(n47071), .B(n45363), .Z(n43683) );
  XOR U56585 ( .A(n43684), .B(n43683), .Z(n45362) );
  XOR U56586 ( .A(n45360), .B(n45362), .Z(n45355) );
  XOR U56587 ( .A(n45354), .B(n45355), .Z(n45358) );
  XOR U56588 ( .A(n43685), .B(n45358), .Z(n43686) );
  IV U56589 ( .A(n43686), .Z(n45353) );
  IV U56590 ( .A(n43687), .Z(n43689) );
  NOR U56591 ( .A(n43689), .B(n43688), .Z(n45351) );
  XOR U56592 ( .A(n45353), .B(n45351), .Z(n45345) );
  IV U56593 ( .A(n45345), .Z(n43697) );
  IV U56594 ( .A(n43690), .Z(n43691) );
  NOR U56595 ( .A(n43692), .B(n43691), .Z(n45347) );
  IV U56596 ( .A(n43693), .Z(n43694) );
  NOR U56597 ( .A(n43695), .B(n43694), .Z(n45344) );
  NOR U56598 ( .A(n45347), .B(n45344), .Z(n43696) );
  XOR U56599 ( .A(n43697), .B(n43696), .Z(n47081) );
  IV U56600 ( .A(n43698), .Z(n43700) );
  NOR U56601 ( .A(n43700), .B(n43699), .Z(n47079) );
  XOR U56602 ( .A(n47081), .B(n47079), .Z(n47084) );
  XOR U56603 ( .A(n47082), .B(n47084), .Z(n47088) );
  XOR U56604 ( .A(n43701), .B(n47088), .Z(n43702) );
  IV U56605 ( .A(n43702), .Z(n45341) );
  XOR U56606 ( .A(n45339), .B(n45341), .Z(n47091) );
  XOR U56607 ( .A(n47090), .B(n47091), .Z(n47094) );
  XOR U56608 ( .A(n47093), .B(n47094), .Z(n45334) );
  XOR U56609 ( .A(n45333), .B(n45334), .Z(n45338) );
  IV U56610 ( .A(n43703), .Z(n43705) );
  NOR U56611 ( .A(n43705), .B(n43704), .Z(n45336) );
  XOR U56612 ( .A(n45338), .B(n45336), .Z(n45331) );
  XOR U56613 ( .A(n43706), .B(n45331), .Z(n45319) );
  NOR U56614 ( .A(n45320), .B(n43707), .Z(n43711) );
  IV U56615 ( .A(n43708), .Z(n43709) );
  NOR U56616 ( .A(n43710), .B(n43709), .Z(n47100) );
  NOR U56617 ( .A(n43711), .B(n47100), .Z(n43712) );
  XOR U56618 ( .A(n45319), .B(n43712), .Z(n47110) );
  XOR U56619 ( .A(n47109), .B(n47110), .Z(n47113) );
  XOR U56620 ( .A(n47112), .B(n47113), .Z(n45314) );
  IV U56621 ( .A(n43713), .Z(n43714) );
  NOR U56622 ( .A(n43714), .B(n43716), .Z(n45316) );
  IV U56623 ( .A(n43715), .Z(n43717) );
  NOR U56624 ( .A(n43717), .B(n43716), .Z(n45313) );
  NOR U56625 ( .A(n45316), .B(n45313), .Z(n43718) );
  XOR U56626 ( .A(n45314), .B(n43718), .Z(n43721) );
  IV U56627 ( .A(n43721), .Z(n43720) );
  IV U56628 ( .A(n43722), .Z(n43719) );
  NOR U56629 ( .A(n43720), .B(n43719), .Z(n48748) );
  NOR U56630 ( .A(n43722), .B(n43721), .Z(n47117) );
  IV U56631 ( .A(n43723), .Z(n43729) );
  IV U56632 ( .A(n43724), .Z(n43725) );
  NOR U56633 ( .A(n43726), .B(n43725), .Z(n43727) );
  IV U56634 ( .A(n43727), .Z(n43728) );
  NOR U56635 ( .A(n43729), .B(n43728), .Z(n47115) );
  XOR U56636 ( .A(n47117), .B(n47115), .Z(n43730) );
  NOR U56637 ( .A(n48748), .B(n43730), .Z(n45309) );
  XOR U56638 ( .A(n45311), .B(n45309), .Z(n47129) );
  XOR U56639 ( .A(n43731), .B(n47129), .Z(n43732) );
  IV U56640 ( .A(n43732), .Z(n45304) );
  XOR U56641 ( .A(n45303), .B(n45304), .Z(n45307) );
  IV U56642 ( .A(n45307), .Z(n43740) );
  IV U56643 ( .A(n43733), .Z(n43734) );
  NOR U56644 ( .A(n43735), .B(n43734), .Z(n45306) );
  IV U56645 ( .A(n43736), .Z(n43737) );
  NOR U56646 ( .A(n43738), .B(n43737), .Z(n45298) );
  NOR U56647 ( .A(n45306), .B(n45298), .Z(n43739) );
  XOR U56648 ( .A(n43740), .B(n43739), .Z(n45301) );
  XOR U56649 ( .A(n45300), .B(n45301), .Z(n45294) );
  XOR U56650 ( .A(n45292), .B(n45294), .Z(n45296) );
  XOR U56651 ( .A(n43741), .B(n45296), .Z(n43742) );
  IV U56652 ( .A(n43742), .Z(n45290) );
  XOR U56653 ( .A(n45289), .B(n45290), .Z(n47138) );
  IV U56654 ( .A(n43743), .Z(n43748) );
  IV U56655 ( .A(n43744), .Z(n43745) );
  NOR U56656 ( .A(n43746), .B(n43745), .Z(n43747) );
  IV U56657 ( .A(n43747), .Z(n43750) );
  NOR U56658 ( .A(n43748), .B(n43750), .Z(n47136) );
  XOR U56659 ( .A(n47138), .B(n47136), .Z(n45286) );
  IV U56660 ( .A(n43749), .Z(n43751) );
  NOR U56661 ( .A(n43751), .B(n43750), .Z(n45284) );
  XOR U56662 ( .A(n45286), .B(n45284), .Z(n47143) );
  XOR U56663 ( .A(n47142), .B(n47143), .Z(n47146) );
  XOR U56664 ( .A(n47145), .B(n47146), .Z(n45280) );
  IV U56665 ( .A(n43752), .Z(n43754) );
  NOR U56666 ( .A(n43754), .B(n43753), .Z(n45278) );
  XOR U56667 ( .A(n45280), .B(n45278), .Z(n45282) );
  IV U56668 ( .A(n45282), .Z(n43762) );
  IV U56669 ( .A(n43755), .Z(n43756) );
  NOR U56670 ( .A(n43757), .B(n43756), .Z(n45281) );
  IV U56671 ( .A(n43758), .Z(n43760) );
  NOR U56672 ( .A(n43760), .B(n43759), .Z(n45276) );
  NOR U56673 ( .A(n45281), .B(n45276), .Z(n43761) );
  XOR U56674 ( .A(n43762), .B(n43761), .Z(n47151) );
  XOR U56675 ( .A(n47150), .B(n47151), .Z(n47155) );
  XOR U56676 ( .A(n47153), .B(n47155), .Z(n52383) );
  XOR U56677 ( .A(n47158), .B(n52383), .Z(n43763) );
  IV U56678 ( .A(n43763), .Z(n47160) );
  XOR U56679 ( .A(n47159), .B(n47160), .Z(n47164) );
  XOR U56680 ( .A(n47163), .B(n47164), .Z(n45275) );
  IV U56681 ( .A(n43764), .Z(n43770) );
  IV U56682 ( .A(n43765), .Z(n43766) );
  NOR U56683 ( .A(n43767), .B(n43766), .Z(n43768) );
  IV U56684 ( .A(n43768), .Z(n43769) );
  NOR U56685 ( .A(n43770), .B(n43769), .Z(n45273) );
  XOR U56686 ( .A(n45275), .B(n45273), .Z(n54222) );
  XOR U56687 ( .A(n47175), .B(n54222), .Z(n47176) );
  XOR U56688 ( .A(n47177), .B(n47176), .Z(n47183) );
  XOR U56689 ( .A(n47182), .B(n47183), .Z(n45271) );
  XOR U56690 ( .A(n43771), .B(n45271), .Z(n47196) );
  IV U56691 ( .A(n43772), .Z(n43774) );
  NOR U56692 ( .A(n43774), .B(n43773), .Z(n43775) );
  IV U56693 ( .A(n43775), .Z(n47197) );
  XOR U56694 ( .A(n47196), .B(n47197), .Z(n47199) );
  XOR U56695 ( .A(n47200), .B(n47199), .Z(n45261) );
  IV U56696 ( .A(n43776), .Z(n43777) );
  NOR U56697 ( .A(n43778), .B(n43777), .Z(n45262) );
  IV U56698 ( .A(n43779), .Z(n43781) );
  NOR U56699 ( .A(n43781), .B(n43780), .Z(n45265) );
  NOR U56700 ( .A(n45262), .B(n45265), .Z(n43782) );
  XOR U56701 ( .A(n45261), .B(n43782), .Z(n45256) );
  IV U56702 ( .A(n43783), .Z(n43784) );
  NOR U56703 ( .A(n43784), .B(n43790), .Z(n45254) );
  XOR U56704 ( .A(n45256), .B(n45254), .Z(n45258) );
  IV U56705 ( .A(n43785), .Z(n43786) );
  NOR U56706 ( .A(n43787), .B(n43786), .Z(n43788) );
  IV U56707 ( .A(n43788), .Z(n43795) );
  NOR U56708 ( .A(n45258), .B(n43795), .Z(n50712) );
  IV U56709 ( .A(n43789), .Z(n43791) );
  NOR U56710 ( .A(n43791), .B(n43790), .Z(n45257) );
  XOR U56711 ( .A(n45257), .B(n45258), .Z(n47205) );
  IV U56712 ( .A(n43792), .Z(n43794) );
  NOR U56713 ( .A(n43794), .B(n43793), .Z(n43796) );
  IV U56714 ( .A(n43796), .Z(n47204) );
  XOR U56715 ( .A(n47205), .B(n47204), .Z(n43798) );
  NOR U56716 ( .A(n43796), .B(n43795), .Z(n43797) );
  NOR U56717 ( .A(n43798), .B(n43797), .Z(n43799) );
  NOR U56718 ( .A(n50712), .B(n43799), .Z(n47206) );
  XOR U56719 ( .A(n43800), .B(n47206), .Z(n47211) );
  IV U56720 ( .A(n43801), .Z(n43803) );
  NOR U56721 ( .A(n43803), .B(n43802), .Z(n47210) );
  IV U56722 ( .A(n43804), .Z(n43805) );
  NOR U56723 ( .A(n43805), .B(n43809), .Z(n45252) );
  NOR U56724 ( .A(n47210), .B(n45252), .Z(n43806) );
  XOR U56725 ( .A(n47211), .B(n43806), .Z(n45246) );
  IV U56726 ( .A(n43807), .Z(n43808) );
  NOR U56727 ( .A(n43809), .B(n43808), .Z(n45249) );
  IV U56728 ( .A(n43810), .Z(n43811) );
  NOR U56729 ( .A(n43812), .B(n43811), .Z(n45247) );
  NOR U56730 ( .A(n45249), .B(n45247), .Z(n43813) );
  XOR U56731 ( .A(n45246), .B(n43813), .Z(n45244) );
  IV U56732 ( .A(n43814), .Z(n43815) );
  NOR U56733 ( .A(n43815), .B(n43817), .Z(n45242) );
  XOR U56734 ( .A(n45244), .B(n45242), .Z(n48709) );
  IV U56735 ( .A(n48709), .Z(n43822) );
  IV U56736 ( .A(n43816), .Z(n43818) );
  NOR U56737 ( .A(n43818), .B(n43817), .Z(n48713) );
  IV U56738 ( .A(n43819), .Z(n43820) );
  NOR U56739 ( .A(n43821), .B(n43820), .Z(n48708) );
  NOR U56740 ( .A(n48713), .B(n48708), .Z(n47227) );
  XOR U56741 ( .A(n43822), .B(n47227), .Z(n47233) );
  XOR U56742 ( .A(n47228), .B(n47233), .Z(n47241) );
  XOR U56743 ( .A(n43823), .B(n47241), .Z(n45239) );
  XOR U56744 ( .A(n43824), .B(n45239), .Z(n45236) );
  XOR U56745 ( .A(n45234), .B(n45236), .Z(n48695) );
  XOR U56746 ( .A(n45237), .B(n48695), .Z(n45232) );
  NOR U56747 ( .A(n43826), .B(n43825), .Z(n45231) );
  IV U56748 ( .A(n43827), .Z(n43829) );
  NOR U56749 ( .A(n43829), .B(n43828), .Z(n47256) );
  NOR U56750 ( .A(n45231), .B(n47256), .Z(n43830) );
  XOR U56751 ( .A(n45232), .B(n43830), .Z(n45230) );
  XOR U56752 ( .A(n45228), .B(n45230), .Z(n47265) );
  XOR U56753 ( .A(n47264), .B(n47265), .Z(n47269) );
  NOR U56754 ( .A(n43831), .B(n47269), .Z(n47280) );
  IV U56755 ( .A(n43832), .Z(n43833) );
  NOR U56756 ( .A(n43836), .B(n43833), .Z(n43834) );
  IV U56757 ( .A(n43834), .Z(n45226) );
  IV U56758 ( .A(n43835), .Z(n43837) );
  NOR U56759 ( .A(n43837), .B(n43836), .Z(n47267) );
  XOR U56760 ( .A(n47269), .B(n47267), .Z(n45225) );
  XOR U56761 ( .A(n45226), .B(n45225), .Z(n43838) );
  NOR U56762 ( .A(n43839), .B(n43838), .Z(n43840) );
  NOR U56763 ( .A(n47280), .B(n43840), .Z(n47274) );
  IV U56764 ( .A(n43841), .Z(n43842) );
  NOR U56765 ( .A(n43843), .B(n43842), .Z(n43844) );
  IV U56766 ( .A(n43844), .Z(n47275) );
  XOR U56767 ( .A(n47274), .B(n47275), .Z(n45223) );
  XOR U56768 ( .A(n45222), .B(n45223), .Z(n47286) );
  XOR U56769 ( .A(n47285), .B(n47286), .Z(n47290) );
  IV U56770 ( .A(n43845), .Z(n43847) );
  NOR U56771 ( .A(n43847), .B(n43846), .Z(n45219) );
  IV U56772 ( .A(n43848), .Z(n43849) );
  NOR U56773 ( .A(n43850), .B(n43849), .Z(n47288) );
  NOR U56774 ( .A(n45219), .B(n47288), .Z(n43851) );
  XOR U56775 ( .A(n47290), .B(n43851), .Z(n45217) );
  XOR U56776 ( .A(n45218), .B(n45217), .Z(n48668) );
  IV U56777 ( .A(n43852), .Z(n43854) );
  NOR U56778 ( .A(n43854), .B(n43853), .Z(n50788) );
  IV U56779 ( .A(n43855), .Z(n43857) );
  NOR U56780 ( .A(n43857), .B(n43856), .Z(n48667) );
  NOR U56781 ( .A(n50788), .B(n48667), .Z(n45212) );
  XOR U56782 ( .A(n48668), .B(n45212), .Z(n45213) );
  XOR U56783 ( .A(n45214), .B(n45213), .Z(n45208) );
  XOR U56784 ( .A(n45207), .B(n45208), .Z(n45210) );
  IV U56785 ( .A(n43858), .Z(n43860) );
  NOR U56786 ( .A(n43860), .B(n43859), .Z(n43865) );
  IV U56787 ( .A(n43861), .Z(n43862) );
  NOR U56788 ( .A(n43863), .B(n43862), .Z(n43864) );
  NOR U56789 ( .A(n43865), .B(n43864), .Z(n45211) );
  XOR U56790 ( .A(n45210), .B(n45211), .Z(n45205) );
  XOR U56791 ( .A(n43866), .B(n45205), .Z(n47297) );
  XOR U56792 ( .A(n47295), .B(n47297), .Z(n45198) );
  IV U56793 ( .A(n45198), .Z(n43873) );
  IV U56794 ( .A(n43867), .Z(n45199) );
  NOR U56795 ( .A(n45201), .B(n45199), .Z(n43871) );
  IV U56796 ( .A(n43868), .Z(n43870) );
  NOR U56797 ( .A(n43870), .B(n43869), .Z(n45196) );
  NOR U56798 ( .A(n43871), .B(n45196), .Z(n43872) );
  XOR U56799 ( .A(n43873), .B(n43872), .Z(n47309) );
  IV U56800 ( .A(n43874), .Z(n43876) );
  NOR U56801 ( .A(n43876), .B(n43875), .Z(n47307) );
  XOR U56802 ( .A(n47309), .B(n47307), .Z(n47311) );
  XOR U56803 ( .A(n47310), .B(n47311), .Z(n47315) );
  XOR U56804 ( .A(n47314), .B(n47315), .Z(n47319) );
  XOR U56805 ( .A(n47317), .B(n47319), .Z(n47323) );
  XOR U56806 ( .A(n47321), .B(n47323), .Z(n47325) );
  XOR U56807 ( .A(n47324), .B(n47325), .Z(n48623) );
  XOR U56808 ( .A(n45195), .B(n48623), .Z(n43877) );
  IV U56809 ( .A(n43877), .Z(n47338) );
  XOR U56810 ( .A(n47337), .B(n47338), .Z(n47331) );
  IV U56811 ( .A(n43878), .Z(n43880) );
  NOR U56812 ( .A(n43880), .B(n43879), .Z(n47329) );
  XOR U56813 ( .A(n47331), .B(n47329), .Z(n47334) );
  XOR U56814 ( .A(n47333), .B(n47334), .Z(n45194) );
  XOR U56815 ( .A(n45190), .B(n45194), .Z(n47356) );
  IV U56816 ( .A(n43881), .Z(n43882) );
  NOR U56817 ( .A(n43882), .B(n43884), .Z(n45192) );
  IV U56818 ( .A(n43883), .Z(n43887) );
  NOR U56819 ( .A(n43885), .B(n43884), .Z(n43886) );
  IV U56820 ( .A(n43886), .Z(n43893) );
  NOR U56821 ( .A(n43887), .B(n43893), .Z(n47354) );
  NOR U56822 ( .A(n45192), .B(n47354), .Z(n43888) );
  XOR U56823 ( .A(n47356), .B(n43888), .Z(n47351) );
  IV U56824 ( .A(n43889), .Z(n43901) );
  IV U56825 ( .A(n43890), .Z(n43891) );
  NOR U56826 ( .A(n43901), .B(n43891), .Z(n47360) );
  IV U56827 ( .A(n43892), .Z(n43894) );
  NOR U56828 ( .A(n43894), .B(n43893), .Z(n47352) );
  NOR U56829 ( .A(n47360), .B(n47352), .Z(n43895) );
  XOR U56830 ( .A(n47351), .B(n43895), .Z(n47366) );
  IV U56831 ( .A(n43896), .Z(n43898) );
  NOR U56832 ( .A(n43898), .B(n43897), .Z(n47364) );
  IV U56833 ( .A(n43899), .Z(n43900) );
  NOR U56834 ( .A(n43901), .B(n43900), .Z(n47358) );
  NOR U56835 ( .A(n47364), .B(n47358), .Z(n43902) );
  XOR U56836 ( .A(n47366), .B(n43902), .Z(n47367) );
  XOR U56837 ( .A(n47368), .B(n47367), .Z(n48603) );
  XOR U56838 ( .A(n43903), .B(n48603), .Z(n43904) );
  IV U56839 ( .A(n43904), .Z(n50827) );
  XOR U56840 ( .A(n50825), .B(n50827), .Z(n45185) );
  IV U56841 ( .A(n45185), .Z(n47380) );
  IV U56842 ( .A(n43905), .Z(n43910) );
  IV U56843 ( .A(n43906), .Z(n43907) );
  NOR U56844 ( .A(n43910), .B(n43907), .Z(n43908) );
  IV U56845 ( .A(n43908), .Z(n45184) );
  XOR U56846 ( .A(n47380), .B(n45184), .Z(n47373) );
  IV U56847 ( .A(n43909), .Z(n43911) );
  NOR U56848 ( .A(n43911), .B(n43910), .Z(n47371) );
  XOR U56849 ( .A(n47373), .B(n47371), .Z(n48592) );
  IV U56850 ( .A(n43912), .Z(n43913) );
  NOR U56851 ( .A(n43914), .B(n43913), .Z(n45182) );
  NOR U56852 ( .A(n45181), .B(n45182), .Z(n43915) );
  XOR U56853 ( .A(n48592), .B(n43915), .Z(n47386) );
  XOR U56854 ( .A(n43916), .B(n47386), .Z(n47393) );
  XOR U56855 ( .A(n47392), .B(n47393), .Z(n47404) );
  IV U56856 ( .A(n43917), .Z(n43919) );
  NOR U56857 ( .A(n43919), .B(n43918), .Z(n45179) );
  IV U56858 ( .A(n43920), .Z(n43922) );
  NOR U56859 ( .A(n43922), .B(n43921), .Z(n47403) );
  NOR U56860 ( .A(n45179), .B(n47403), .Z(n43923) );
  XOR U56861 ( .A(n47404), .B(n43923), .Z(n43924) );
  IV U56862 ( .A(n43924), .Z(n43932) );
  NOR U56863 ( .A(n43925), .B(n43932), .Z(n47402) );
  IV U56864 ( .A(n43926), .Z(n43927) );
  NOR U56865 ( .A(n43928), .B(n43927), .Z(n43934) );
  IV U56866 ( .A(n43934), .Z(n43930) );
  XOR U56867 ( .A(n45179), .B(n47404), .Z(n43929) );
  NOR U56868 ( .A(n43930), .B(n43929), .Z(n45178) );
  NOR U56869 ( .A(n47402), .B(n45178), .Z(n43931) );
  IV U56870 ( .A(n43931), .Z(n43935) );
  NOR U56871 ( .A(n43935), .B(n43932), .Z(n43938) );
  NOR U56872 ( .A(n43934), .B(n43933), .Z(n43936) );
  NOR U56873 ( .A(n43936), .B(n43935), .Z(n43937) );
  NOR U56874 ( .A(n43938), .B(n43937), .Z(n45176) );
  XOR U56875 ( .A(n45175), .B(n45176), .Z(n47423) );
  XOR U56876 ( .A(n47422), .B(n47423), .Z(n47419) );
  XOR U56877 ( .A(n47418), .B(n47419), .Z(n45173) );
  XOR U56878 ( .A(n45172), .B(n45173), .Z(n47434) );
  XOR U56879 ( .A(n47435), .B(n47434), .Z(n45170) );
  IV U56880 ( .A(n43939), .Z(n43941) );
  NOR U56881 ( .A(n43941), .B(n43940), .Z(n47436) );
  IV U56882 ( .A(n43942), .Z(n43944) );
  NOR U56883 ( .A(n43944), .B(n43943), .Z(n47439) );
  NOR U56884 ( .A(n47439), .B(n45169), .Z(n43945) );
  XOR U56885 ( .A(n47436), .B(n43945), .Z(n43946) );
  XOR U56886 ( .A(n45170), .B(n43946), .Z(n45166) );
  XOR U56887 ( .A(n45164), .B(n45166), .Z(n47443) );
  IV U56888 ( .A(n47443), .Z(n43954) );
  IV U56889 ( .A(n43947), .Z(n43949) );
  NOR U56890 ( .A(n43949), .B(n43948), .Z(n45167) );
  IV U56891 ( .A(n43950), .Z(n43952) );
  NOR U56892 ( .A(n43952), .B(n43951), .Z(n47442) );
  NOR U56893 ( .A(n45167), .B(n47442), .Z(n43953) );
  XOR U56894 ( .A(n43954), .B(n43953), .Z(n47446) );
  XOR U56895 ( .A(n47445), .B(n47446), .Z(n47451) );
  XOR U56896 ( .A(n47449), .B(n47451), .Z(n47454) );
  XOR U56897 ( .A(n47452), .B(n47454), .Z(n47458) );
  XOR U56898 ( .A(n47456), .B(n47458), .Z(n47460) );
  XOR U56899 ( .A(n43955), .B(n47460), .Z(n45156) );
  XOR U56900 ( .A(n43956), .B(n45156), .Z(n47472) );
  XOR U56901 ( .A(n45155), .B(n47472), .Z(n43957) );
  IV U56902 ( .A(n43957), .Z(n45153) );
  XOR U56903 ( .A(n45152), .B(n45153), .Z(n47480) );
  XOR U56904 ( .A(n47479), .B(n47480), .Z(n47483) );
  XOR U56905 ( .A(n47482), .B(n47483), .Z(n45150) );
  XOR U56906 ( .A(n45149), .B(n45150), .Z(n45145) );
  IV U56907 ( .A(n43958), .Z(n43961) );
  IV U56908 ( .A(n43959), .Z(n43960) );
  NOR U56909 ( .A(n43961), .B(n43960), .Z(n45143) );
  XOR U56910 ( .A(n45145), .B(n45143), .Z(n45148) );
  IV U56911 ( .A(n43962), .Z(n43966) );
  NOR U56912 ( .A(n43964), .B(n43963), .Z(n43965) );
  IV U56913 ( .A(n43965), .Z(n43968) );
  NOR U56914 ( .A(n43966), .B(n43968), .Z(n45146) );
  XOR U56915 ( .A(n45148), .B(n45146), .Z(n45142) );
  IV U56916 ( .A(n43967), .Z(n43969) );
  NOR U56917 ( .A(n43969), .B(n43968), .Z(n45140) );
  XOR U56918 ( .A(n45142), .B(n45140), .Z(n47490) );
  XOR U56919 ( .A(n47489), .B(n47490), .Z(n47496) );
  IV U56920 ( .A(n47496), .Z(n43973) );
  NOR U56921 ( .A(n43971), .B(n43970), .Z(n47492) );
  NOR U56922 ( .A(n47492), .B(n47495), .Z(n43972) );
  XOR U56923 ( .A(n43973), .B(n43972), .Z(n47499) );
  XOR U56924 ( .A(n47498), .B(n47499), .Z(n47502) );
  XOR U56925 ( .A(n47501), .B(n47502), .Z(n47505) );
  XOR U56926 ( .A(n47504), .B(n47505), .Z(n47516) );
  XOR U56927 ( .A(n43974), .B(n47516), .Z(n47518) );
  IV U56928 ( .A(n43975), .Z(n43977) );
  NOR U56929 ( .A(n43977), .B(n43976), .Z(n47517) );
  IV U56930 ( .A(n43978), .Z(n43987) );
  IV U56931 ( .A(n43979), .Z(n43980) );
  NOR U56932 ( .A(n43987), .B(n43980), .Z(n47522) );
  NOR U56933 ( .A(n47517), .B(n47522), .Z(n43981) );
  XOR U56934 ( .A(n47518), .B(n43981), .Z(n45139) );
  IV U56935 ( .A(n45139), .Z(n43989) );
  IV U56936 ( .A(n43982), .Z(n43984) );
  NOR U56937 ( .A(n43984), .B(n43983), .Z(n45135) );
  IV U56938 ( .A(n43985), .Z(n43986) );
  NOR U56939 ( .A(n43987), .B(n43986), .Z(n45137) );
  NOR U56940 ( .A(n45135), .B(n45137), .Z(n43988) );
  XOR U56941 ( .A(n43989), .B(n43988), .Z(n47526) );
  XOR U56942 ( .A(n47525), .B(n47526), .Z(n47529) );
  IV U56943 ( .A(n47529), .Z(n43997) );
  IV U56944 ( .A(n43990), .Z(n43992) );
  NOR U56945 ( .A(n43992), .B(n43991), .Z(n47528) );
  IV U56946 ( .A(n43993), .Z(n43995) );
  NOR U56947 ( .A(n43995), .B(n43994), .Z(n45133) );
  NOR U56948 ( .A(n47528), .B(n45133), .Z(n43996) );
  XOR U56949 ( .A(n43997), .B(n43996), .Z(n45132) );
  XOR U56950 ( .A(n45130), .B(n45132), .Z(n45126) );
  XOR U56951 ( .A(n45124), .B(n45126), .Z(n45128) );
  XOR U56952 ( .A(n45127), .B(n45128), .Z(n45120) );
  XOR U56953 ( .A(n45118), .B(n45120), .Z(n45123) );
  XOR U56954 ( .A(n45121), .B(n45123), .Z(n45114) );
  XOR U56955 ( .A(n45112), .B(n45114), .Z(n45117) );
  XOR U56956 ( .A(n45115), .B(n45117), .Z(n48484) );
  XOR U56957 ( .A(n47536), .B(n48484), .Z(n47537) );
  IV U56958 ( .A(n43998), .Z(n44000) );
  NOR U56959 ( .A(n44000), .B(n43999), .Z(n48474) );
  IV U56960 ( .A(n44001), .Z(n44003) );
  NOR U56961 ( .A(n44003), .B(n44002), .Z(n50902) );
  NOR U56962 ( .A(n48474), .B(n50902), .Z(n47538) );
  XOR U56963 ( .A(n47537), .B(n47538), .Z(n47545) );
  IV U56964 ( .A(n44004), .Z(n44013) );
  IV U56965 ( .A(n44005), .Z(n44006) );
  NOR U56966 ( .A(n44013), .B(n44006), .Z(n47542) );
  NOR U56967 ( .A(n47546), .B(n50901), .Z(n44007) );
  NOR U56968 ( .A(n47542), .B(n44007), .Z(n44008) );
  XOR U56969 ( .A(n47545), .B(n44008), .Z(n45110) );
  IV U56970 ( .A(n44009), .Z(n44010) );
  NOR U56971 ( .A(n44011), .B(n44010), .Z(n45109) );
  IV U56972 ( .A(n44012), .Z(n44014) );
  NOR U56973 ( .A(n44014), .B(n44013), .Z(n47549) );
  NOR U56974 ( .A(n45109), .B(n47549), .Z(n44015) );
  XOR U56975 ( .A(n45110), .B(n44015), .Z(n47565) );
  XOR U56976 ( .A(n47564), .B(n47565), .Z(n44021) );
  IV U56977 ( .A(n44021), .Z(n44016) );
  NOR U56978 ( .A(n44017), .B(n44016), .Z(n45106) );
  IV U56979 ( .A(n44018), .Z(n47572) );
  NOR U56980 ( .A(n47572), .B(n44019), .Z(n44022) );
  IV U56981 ( .A(n44022), .Z(n44020) );
  NOR U56982 ( .A(n47565), .B(n44020), .Z(n48462) );
  NOR U56983 ( .A(n44022), .B(n44021), .Z(n47573) );
  NOR U56984 ( .A(n48462), .B(n47573), .Z(n44023) );
  NOR U56985 ( .A(n44024), .B(n44023), .Z(n44025) );
  NOR U56986 ( .A(n45106), .B(n44025), .Z(n47580) );
  XOR U56987 ( .A(n44026), .B(n47580), .Z(n47586) );
  XOR U56988 ( .A(n47585), .B(n47586), .Z(n45103) );
  XOR U56989 ( .A(n45100), .B(n45103), .Z(n47589) );
  IV U56990 ( .A(n47589), .Z(n44034) );
  IV U56991 ( .A(n44027), .Z(n44028) );
  NOR U56992 ( .A(n44029), .B(n44028), .Z(n45102) );
  IV U56993 ( .A(n44030), .Z(n44032) );
  NOR U56994 ( .A(n44032), .B(n44031), .Z(n47588) );
  NOR U56995 ( .A(n45102), .B(n47588), .Z(n44033) );
  XOR U56996 ( .A(n44034), .B(n44033), .Z(n47595) );
  IV U56997 ( .A(n44035), .Z(n44036) );
  NOR U56998 ( .A(n44037), .B(n44036), .Z(n45098) );
  XOR U56999 ( .A(n47595), .B(n45098), .Z(n47593) );
  XOR U57000 ( .A(n47591), .B(n47593), .Z(n45096) );
  XOR U57001 ( .A(n44038), .B(n45096), .Z(n44039) );
  IV U57002 ( .A(n44039), .Z(n45094) );
  XOR U57003 ( .A(n45092), .B(n45094), .Z(n47606) );
  XOR U57004 ( .A(n47605), .B(n47606), .Z(n47610) );
  NOR U57005 ( .A(n44041), .B(n44040), .Z(n44042) );
  IV U57006 ( .A(n44042), .Z(n44047) );
  NOR U57007 ( .A(n44044), .B(n44043), .Z(n44045) );
  IV U57008 ( .A(n44045), .Z(n44046) );
  NOR U57009 ( .A(n44047), .B(n44046), .Z(n47608) );
  XOR U57010 ( .A(n47610), .B(n47608), .Z(n45091) );
  IV U57011 ( .A(n44048), .Z(n44049) );
  NOR U57012 ( .A(n44050), .B(n44049), .Z(n45087) );
  IV U57013 ( .A(n44051), .Z(n44052) );
  NOR U57014 ( .A(n44053), .B(n44052), .Z(n45089) );
  NOR U57015 ( .A(n45087), .B(n45089), .Z(n44054) );
  XOR U57016 ( .A(n45091), .B(n44054), .Z(n45078) );
  IV U57017 ( .A(n44055), .Z(n44057) );
  NOR U57018 ( .A(n44057), .B(n44056), .Z(n45084) );
  IV U57019 ( .A(n44058), .Z(n44060) );
  NOR U57020 ( .A(n44060), .B(n44059), .Z(n45079) );
  NOR U57021 ( .A(n45084), .B(n45079), .Z(n44061) );
  XOR U57022 ( .A(n45078), .B(n44061), .Z(n45082) );
  IV U57023 ( .A(n44062), .Z(n44063) );
  NOR U57024 ( .A(n44064), .B(n44063), .Z(n45081) );
  IV U57025 ( .A(n44065), .Z(n44067) );
  NOR U57026 ( .A(n44067), .B(n44066), .Z(n45076) );
  NOR U57027 ( .A(n45081), .B(n45076), .Z(n44068) );
  XOR U57028 ( .A(n45082), .B(n44068), .Z(n45073) );
  IV U57029 ( .A(n44069), .Z(n44070) );
  NOR U57030 ( .A(n44071), .B(n44070), .Z(n44072) );
  IV U57031 ( .A(n44072), .Z(n45074) );
  XOR U57032 ( .A(n45073), .B(n45074), .Z(n47619) );
  XOR U57033 ( .A(n47617), .B(n47619), .Z(n45071) );
  XOR U57034 ( .A(n45069), .B(n45071), .Z(n47614) );
  NOR U57035 ( .A(n44073), .B(n45062), .Z(n44077) );
  IV U57036 ( .A(n44074), .Z(n44075) );
  NOR U57037 ( .A(n44076), .B(n44075), .Z(n47613) );
  XOR U57038 ( .A(n44077), .B(n47613), .Z(n44078) );
  XOR U57039 ( .A(n47614), .B(n44078), .Z(n48440) );
  XOR U57040 ( .A(n47625), .B(n48440), .Z(n44079) );
  IV U57041 ( .A(n44079), .Z(n45059) );
  IV U57042 ( .A(n44080), .Z(n44081) );
  NOR U57043 ( .A(n44087), .B(n44081), .Z(n45057) );
  XOR U57044 ( .A(n45059), .B(n45057), .Z(n48432) );
  IV U57045 ( .A(n48432), .Z(n44088) );
  IV U57046 ( .A(n44082), .Z(n44083) );
  NOR U57047 ( .A(n44084), .B(n44083), .Z(n45055) );
  IV U57048 ( .A(n44085), .Z(n44086) );
  NOR U57049 ( .A(n44087), .B(n44086), .Z(n47626) );
  NOR U57050 ( .A(n45055), .B(n47626), .Z(n48433) );
  XOR U57051 ( .A(n44088), .B(n48433), .Z(n45053) );
  XOR U57052 ( .A(n45052), .B(n45053), .Z(n45047) );
  XOR U57053 ( .A(n45046), .B(n45047), .Z(n45050) );
  XOR U57054 ( .A(n44089), .B(n45050), .Z(n44090) );
  IV U57055 ( .A(n44090), .Z(n45042) );
  XOR U57056 ( .A(n45038), .B(n45042), .Z(n45034) );
  NOR U57057 ( .A(n44091), .B(n44097), .Z(n45040) );
  XOR U57058 ( .A(n44092), .B(n44097), .Z(n44093) );
  NOR U57059 ( .A(n44094), .B(n44093), .Z(n45033) );
  NOR U57060 ( .A(n45040), .B(n45033), .Z(n44095) );
  XOR U57061 ( .A(n45034), .B(n44095), .Z(n45026) );
  IV U57062 ( .A(n44096), .Z(n44098) );
  NOR U57063 ( .A(n44098), .B(n44097), .Z(n45029) );
  IV U57064 ( .A(n44099), .Z(n44104) );
  IV U57065 ( .A(n44100), .Z(n44101) );
  NOR U57066 ( .A(n44104), .B(n44101), .Z(n45027) );
  NOR U57067 ( .A(n45029), .B(n45027), .Z(n44102) );
  XOR U57068 ( .A(n45026), .B(n44102), .Z(n45022) );
  IV U57069 ( .A(n44103), .Z(n44105) );
  NOR U57070 ( .A(n44105), .B(n44104), .Z(n45020) );
  XOR U57071 ( .A(n45022), .B(n45020), .Z(n45024) );
  XOR U57072 ( .A(n45023), .B(n45024), .Z(n45018) );
  XOR U57073 ( .A(n45015), .B(n45018), .Z(n45012) );
  IV U57074 ( .A(n45012), .Z(n44109) );
  NOR U57075 ( .A(n44107), .B(n44106), .Z(n45017) );
  NOR U57076 ( .A(n45017), .B(n45011), .Z(n44108) );
  XOR U57077 ( .A(n44109), .B(n44108), .Z(n47640) );
  XOR U57078 ( .A(n47638), .B(n47640), .Z(n47647) );
  IV U57079 ( .A(n44110), .Z(n45008) );
  NOR U57080 ( .A(n44111), .B(n45008), .Z(n44115) );
  IV U57081 ( .A(n44112), .Z(n44114) );
  NOR U57082 ( .A(n44114), .B(n44113), .Z(n47645) );
  NOR U57083 ( .A(n44115), .B(n47645), .Z(n44116) );
  XOR U57084 ( .A(n47647), .B(n44116), .Z(n47648) );
  XOR U57085 ( .A(n47649), .B(n47648), .Z(n47651) );
  XOR U57086 ( .A(n47650), .B(n47651), .Z(n47657) );
  IV U57087 ( .A(n44117), .Z(n44118) );
  NOR U57088 ( .A(n44119), .B(n44118), .Z(n47656) );
  IV U57089 ( .A(n44120), .Z(n44122) );
  NOR U57090 ( .A(n44122), .B(n44121), .Z(n45005) );
  NOR U57091 ( .A(n47656), .B(n45005), .Z(n44123) );
  XOR U57092 ( .A(n47657), .B(n44123), .Z(n44997) );
  NOR U57093 ( .A(n44125), .B(n44124), .Z(n44998) );
  NOR U57094 ( .A(n44998), .B(n44126), .Z(n44127) );
  XOR U57095 ( .A(n44997), .B(n44127), .Z(n47660) );
  XOR U57096 ( .A(n47661), .B(n47660), .Z(n44995) );
  IV U57097 ( .A(n44128), .Z(n44130) );
  NOR U57098 ( .A(n44130), .B(n44129), .Z(n44994) );
  NOR U57099 ( .A(n47662), .B(n44994), .Z(n44131) );
  XOR U57100 ( .A(n44995), .B(n44131), .Z(n44990) );
  XOR U57101 ( .A(n44988), .B(n44990), .Z(n44992) );
  XOR U57102 ( .A(n44991), .B(n44992), .Z(n47668) );
  XOR U57103 ( .A(n47667), .B(n47668), .Z(n47671) );
  XOR U57104 ( .A(n44132), .B(n47671), .Z(n44133) );
  XOR U57105 ( .A(n47670), .B(n44133), .Z(n44976) );
  IV U57106 ( .A(n44134), .Z(n44136) );
  NOR U57107 ( .A(n44136), .B(n44135), .Z(n51066) );
  IV U57108 ( .A(n44137), .Z(n44138) );
  NOR U57109 ( .A(n44138), .B(n44144), .Z(n48388) );
  NOR U57110 ( .A(n51066), .B(n48388), .Z(n44977) );
  XOR U57111 ( .A(n44976), .B(n44977), .Z(n44974) );
  NOR U57112 ( .A(n44146), .B(n44974), .Z(n48383) );
  IV U57113 ( .A(n44139), .Z(n44141) );
  NOR U57114 ( .A(n44141), .B(n44140), .Z(n44142) );
  IV U57115 ( .A(n44142), .Z(n44969) );
  IV U57116 ( .A(n44143), .Z(n44145) );
  NOR U57117 ( .A(n44145), .B(n44144), .Z(n44973) );
  XOR U57118 ( .A(n44973), .B(n44974), .Z(n44968) );
  XOR U57119 ( .A(n44969), .B(n44968), .Z(n44149) );
  IV U57120 ( .A(n44968), .Z(n44147) );
  NOR U57121 ( .A(n44147), .B(n44146), .Z(n44148) );
  NOR U57122 ( .A(n44149), .B(n44148), .Z(n44150) );
  NOR U57123 ( .A(n48383), .B(n44150), .Z(n44151) );
  IV U57124 ( .A(n44151), .Z(n44971) );
  IV U57125 ( .A(n44152), .Z(n44153) );
  NOR U57126 ( .A(n44153), .B(n44155), .Z(n44970) );
  IV U57127 ( .A(n44154), .Z(n44156) );
  NOR U57128 ( .A(n44156), .B(n44155), .Z(n44966) );
  NOR U57129 ( .A(n44970), .B(n44966), .Z(n44157) );
  XOR U57130 ( .A(n44971), .B(n44157), .Z(n44957) );
  IV U57131 ( .A(n44158), .Z(n44174) );
  IV U57132 ( .A(n44159), .Z(n44160) );
  NOR U57133 ( .A(n44174), .B(n44160), .Z(n44958) );
  IV U57134 ( .A(n44161), .Z(n44163) );
  NOR U57135 ( .A(n44163), .B(n44162), .Z(n44963) );
  NOR U57136 ( .A(n44958), .B(n44963), .Z(n44164) );
  XOR U57137 ( .A(n44957), .B(n44164), .Z(n44962) );
  IV U57138 ( .A(n44165), .Z(n44166) );
  NOR U57139 ( .A(n44174), .B(n44166), .Z(n44960) );
  XOR U57140 ( .A(n44962), .B(n44960), .Z(n47682) );
  IV U57141 ( .A(n47682), .Z(n44176) );
  IV U57142 ( .A(n44167), .Z(n44171) );
  NOR U57143 ( .A(n44168), .B(n44179), .Z(n44169) );
  IV U57144 ( .A(n44169), .Z(n44170) );
  NOR U57145 ( .A(n44171), .B(n44170), .Z(n47680) );
  IV U57146 ( .A(n44172), .Z(n44173) );
  NOR U57147 ( .A(n44174), .B(n44173), .Z(n47674) );
  NOR U57148 ( .A(n47680), .B(n47674), .Z(n44175) );
  XOR U57149 ( .A(n44176), .B(n44175), .Z(n47679) );
  IV U57150 ( .A(n44177), .Z(n44178) );
  NOR U57151 ( .A(n44179), .B(n44178), .Z(n44180) );
  IV U57152 ( .A(n44180), .Z(n44181) );
  NOR U57153 ( .A(n44182), .B(n44181), .Z(n47677) );
  XOR U57154 ( .A(n47679), .B(n47677), .Z(n44952) );
  XOR U57155 ( .A(n44951), .B(n44952), .Z(n44955) );
  XOR U57156 ( .A(n44954), .B(n44955), .Z(n47685) );
  XOR U57157 ( .A(n47683), .B(n47685), .Z(n44196) );
  NOR U57158 ( .A(n44184), .B(n44183), .Z(n44185) );
  IV U57159 ( .A(n44185), .Z(n44192) );
  XOR U57160 ( .A(n44187), .B(n44186), .Z(n44189) );
  NOR U57161 ( .A(n44189), .B(n44188), .Z(n44190) );
  IV U57162 ( .A(n44190), .Z(n44191) );
  NOR U57163 ( .A(n44192), .B(n44191), .Z(n44193) );
  IV U57164 ( .A(n44193), .Z(n47684) );
  NOR U57165 ( .A(n44194), .B(n47684), .Z(n44195) );
  NOR U57166 ( .A(n44196), .B(n44195), .Z(n44200) );
  NOR U57167 ( .A(n47688), .B(n47685), .Z(n44197) );
  IV U57168 ( .A(n44197), .Z(n44198) );
  NOR U57169 ( .A(n44198), .B(n47684), .Z(n44199) );
  NOR U57170 ( .A(n44200), .B(n44199), .Z(n47695) );
  XOR U57171 ( .A(n47697), .B(n47695), .Z(n47704) );
  XOR U57172 ( .A(n44201), .B(n47704), .Z(n44202) );
  IV U57173 ( .A(n44202), .Z(n47707) );
  XOR U57174 ( .A(n47706), .B(n47707), .Z(n47709) );
  IV U57175 ( .A(n44203), .Z(n44204) );
  NOR U57176 ( .A(n44205), .B(n44204), .Z(n47708) );
  IV U57177 ( .A(n44206), .Z(n44208) );
  NOR U57178 ( .A(n44208), .B(n44207), .Z(n47713) );
  NOR U57179 ( .A(n47708), .B(n47713), .Z(n44209) );
  XOR U57180 ( .A(n47709), .B(n44209), .Z(n44950) );
  IV U57181 ( .A(n44210), .Z(n44212) );
  NOR U57182 ( .A(n44212), .B(n44211), .Z(n44213) );
  IV U57183 ( .A(n44213), .Z(n44220) );
  NOR U57184 ( .A(n44950), .B(n44220), .Z(n48362) );
  IV U57185 ( .A(n44214), .Z(n44215) );
  NOR U57186 ( .A(n44215), .B(n44226), .Z(n44216) );
  IV U57187 ( .A(n44216), .Z(n44944) );
  IV U57188 ( .A(n44217), .Z(n44219) );
  NOR U57189 ( .A(n44219), .B(n44218), .Z(n44948) );
  XOR U57190 ( .A(n44948), .B(n44950), .Z(n44943) );
  XOR U57191 ( .A(n44944), .B(n44943), .Z(n44223) );
  IV U57192 ( .A(n44943), .Z(n44221) );
  NOR U57193 ( .A(n44221), .B(n44220), .Z(n44222) );
  NOR U57194 ( .A(n44223), .B(n44222), .Z(n44224) );
  NOR U57195 ( .A(n48362), .B(n44224), .Z(n44945) );
  IV U57196 ( .A(n44225), .Z(n44227) );
  NOR U57197 ( .A(n44227), .B(n44226), .Z(n44228) );
  IV U57198 ( .A(n44228), .Z(n44946) );
  XOR U57199 ( .A(n44945), .B(n44946), .Z(n44939) );
  IV U57200 ( .A(n44229), .Z(n44231) );
  NOR U57201 ( .A(n44231), .B(n44230), .Z(n44937) );
  XOR U57202 ( .A(n44939), .B(n44937), .Z(n44941) );
  IV U57203 ( .A(n44941), .Z(n44239) );
  IV U57204 ( .A(n44232), .Z(n44233) );
  NOR U57205 ( .A(n44234), .B(n44233), .Z(n44940) );
  IV U57206 ( .A(n44235), .Z(n44237) );
  NOR U57207 ( .A(n44237), .B(n44236), .Z(n44935) );
  NOR U57208 ( .A(n44940), .B(n44935), .Z(n44238) );
  XOR U57209 ( .A(n44239), .B(n44238), .Z(n44934) );
  XOR U57210 ( .A(n44933), .B(n44934), .Z(n44245) );
  IV U57211 ( .A(n44245), .Z(n44931) );
  NOR U57212 ( .A(n44244), .B(n44931), .Z(n44930) );
  IV U57213 ( .A(n44240), .Z(n44241) );
  NOR U57214 ( .A(n44242), .B(n44241), .Z(n44243) );
  IV U57215 ( .A(n44243), .Z(n44932) );
  XOR U57216 ( .A(n44932), .B(n44931), .Z(n44247) );
  NOR U57217 ( .A(n44245), .B(n44244), .Z(n44246) );
  NOR U57218 ( .A(n44247), .B(n44246), .Z(n44925) );
  NOR U57219 ( .A(n44930), .B(n44925), .Z(n44926) );
  IV U57220 ( .A(n44248), .Z(n44252) );
  NOR U57221 ( .A(n44250), .B(n44249), .Z(n44251) );
  IV U57222 ( .A(n44251), .Z(n44258) );
  NOR U57223 ( .A(n44252), .B(n44258), .Z(n44253) );
  IV U57224 ( .A(n44253), .Z(n44927) );
  XOR U57225 ( .A(n44926), .B(n44927), .Z(n47723) );
  IV U57226 ( .A(n47723), .Z(n44261) );
  IV U57227 ( .A(n44254), .Z(n44256) );
  NOR U57228 ( .A(n44256), .B(n44255), .Z(n47721) );
  IV U57229 ( .A(n44257), .Z(n44259) );
  NOR U57230 ( .A(n44259), .B(n44258), .Z(n44923) );
  NOR U57231 ( .A(n47721), .B(n44923), .Z(n44260) );
  XOR U57232 ( .A(n44261), .B(n44260), .Z(n47726) );
  IV U57233 ( .A(n44262), .Z(n44264) );
  NOR U57234 ( .A(n44264), .B(n44263), .Z(n47724) );
  XOR U57235 ( .A(n47726), .B(n47724), .Z(n47729) );
  XOR U57236 ( .A(n47727), .B(n47729), .Z(n44919) );
  XOR U57237 ( .A(n44918), .B(n44919), .Z(n44922) );
  XOR U57238 ( .A(n44921), .B(n44922), .Z(n47734) );
  XOR U57239 ( .A(n47732), .B(n47734), .Z(n44917) );
  IV U57240 ( .A(n44265), .Z(n44274) );
  IV U57241 ( .A(n44266), .Z(n44267) );
  NOR U57242 ( .A(n44274), .B(n44267), .Z(n44915) );
  IV U57243 ( .A(n44268), .Z(n44269) );
  NOR U57244 ( .A(n44270), .B(n44269), .Z(n47735) );
  NOR U57245 ( .A(n44915), .B(n47735), .Z(n44271) );
  XOR U57246 ( .A(n44917), .B(n44271), .Z(n44910) );
  IV U57247 ( .A(n44272), .Z(n44273) );
  NOR U57248 ( .A(n44274), .B(n44273), .Z(n44913) );
  IV U57249 ( .A(n44275), .Z(n44276) );
  NOR U57250 ( .A(n44279), .B(n44276), .Z(n44911) );
  IV U57251 ( .A(n44277), .Z(n44278) );
  NOR U57252 ( .A(n44279), .B(n44278), .Z(n47748) );
  NOR U57253 ( .A(n44911), .B(n47748), .Z(n44280) );
  IV U57254 ( .A(n44280), .Z(n44281) );
  NOR U57255 ( .A(n44913), .B(n44281), .Z(n44282) );
  XOR U57256 ( .A(n44910), .B(n44282), .Z(n44908) );
  IV U57257 ( .A(n44283), .Z(n44285) );
  NOR U57258 ( .A(n44285), .B(n44284), .Z(n44906) );
  XOR U57259 ( .A(n44908), .B(n44906), .Z(n47756) );
  XOR U57260 ( .A(n47755), .B(n47756), .Z(n47759) );
  XOR U57261 ( .A(n47758), .B(n47759), .Z(n44901) );
  XOR U57262 ( .A(n44900), .B(n44901), .Z(n44904) );
  NOR U57263 ( .A(n44898), .B(n44903), .Z(n44286) );
  XOR U57264 ( .A(n44904), .B(n44286), .Z(n47766) );
  IV U57265 ( .A(n44287), .Z(n44288) );
  NOR U57266 ( .A(n44289), .B(n44288), .Z(n44290) );
  NOR U57267 ( .A(n54685), .B(n44290), .Z(n47767) );
  XOR U57268 ( .A(n47766), .B(n47767), .Z(n47772) );
  IV U57269 ( .A(n44291), .Z(n44292) );
  NOR U57270 ( .A(n44293), .B(n44292), .Z(n47771) );
  IV U57271 ( .A(n44294), .Z(n44297) );
  IV U57272 ( .A(n44295), .Z(n44296) );
  NOR U57273 ( .A(n44297), .B(n44296), .Z(n47768) );
  NOR U57274 ( .A(n47771), .B(n47768), .Z(n44298) );
  XOR U57275 ( .A(n47772), .B(n44298), .Z(n47777) );
  IV U57276 ( .A(n44299), .Z(n44301) );
  NOR U57277 ( .A(n44301), .B(n44300), .Z(n44302) );
  IV U57278 ( .A(n44302), .Z(n47778) );
  XOR U57279 ( .A(n47777), .B(n47778), .Z(n44897) );
  XOR U57280 ( .A(n44895), .B(n44897), .Z(n51156) );
  XOR U57281 ( .A(n47786), .B(n51156), .Z(n47788) );
  IV U57282 ( .A(n44303), .Z(n44304) );
  NOR U57283 ( .A(n44305), .B(n44304), .Z(n47787) );
  IV U57284 ( .A(n44306), .Z(n44307) );
  NOR U57285 ( .A(n44307), .B(n44310), .Z(n47795) );
  NOR U57286 ( .A(n47787), .B(n47795), .Z(n44308) );
  XOR U57287 ( .A(n47788), .B(n44308), .Z(n47794) );
  IV U57288 ( .A(n44309), .Z(n44311) );
  NOR U57289 ( .A(n44311), .B(n44310), .Z(n47792) );
  XOR U57290 ( .A(n47794), .B(n47792), .Z(n47799) );
  XOR U57291 ( .A(n47798), .B(n47799), .Z(n47802) );
  XOR U57292 ( .A(n47801), .B(n47802), .Z(n47806) );
  XOR U57293 ( .A(n47805), .B(n47806), .Z(n47809) );
  XOR U57294 ( .A(n47808), .B(n47809), .Z(n44893) );
  XOR U57295 ( .A(n44891), .B(n44893), .Z(n47815) );
  XOR U57296 ( .A(n47813), .B(n47815), .Z(n47824) );
  XOR U57297 ( .A(n44312), .B(n47824), .Z(n44313) );
  IV U57298 ( .A(n44313), .Z(n47820) );
  XOR U57299 ( .A(n47819), .B(n47820), .Z(n47827) );
  IV U57300 ( .A(n47827), .Z(n44321) );
  IV U57301 ( .A(n44314), .Z(n44315) );
  NOR U57302 ( .A(n44316), .B(n44315), .Z(n47826) );
  IV U57303 ( .A(n44317), .Z(n44318) );
  NOR U57304 ( .A(n44319), .B(n44318), .Z(n44889) );
  NOR U57305 ( .A(n47826), .B(n44889), .Z(n44320) );
  XOR U57306 ( .A(n44321), .B(n44320), .Z(n47837) );
  XOR U57307 ( .A(n47835), .B(n47837), .Z(n47839) );
  XOR U57308 ( .A(n47838), .B(n47839), .Z(n44887) );
  XOR U57309 ( .A(n44322), .B(n44887), .Z(n44878) );
  XOR U57310 ( .A(n44879), .B(n44878), .Z(n44882) );
  XOR U57311 ( .A(n44323), .B(n44882), .Z(n44324) );
  IV U57312 ( .A(n44324), .Z(n44873) );
  XOR U57313 ( .A(n44325), .B(n44873), .Z(n44334) );
  IV U57314 ( .A(n44334), .Z(n44326) );
  NOR U57315 ( .A(n44327), .B(n44326), .Z(n48275) );
  XOR U57316 ( .A(n44328), .B(n44873), .Z(n44333) );
  IV U57317 ( .A(n44329), .Z(n44331) );
  NOR U57318 ( .A(n44331), .B(n44330), .Z(n44335) );
  IV U57319 ( .A(n44335), .Z(n44332) );
  NOR U57320 ( .A(n44333), .B(n44332), .Z(n51204) );
  NOR U57321 ( .A(n44335), .B(n44334), .Z(n44336) );
  NOR U57322 ( .A(n51204), .B(n44336), .Z(n44337) );
  NOR U57323 ( .A(n44338), .B(n44337), .Z(n44339) );
  NOR U57324 ( .A(n48275), .B(n44339), .Z(n44340) );
  IV U57325 ( .A(n44340), .Z(n47848) );
  XOR U57326 ( .A(n47848), .B(n47847), .Z(n47857) );
  NOR U57327 ( .A(n44342), .B(n44341), .Z(n47850) );
  IV U57328 ( .A(n44343), .Z(n44345) );
  NOR U57329 ( .A(n44345), .B(n44344), .Z(n47855) );
  NOR U57330 ( .A(n47850), .B(n47855), .Z(n44346) );
  XOR U57331 ( .A(n47857), .B(n44346), .Z(n47853) );
  XOR U57332 ( .A(n47854), .B(n47853), .Z(n44867) );
  XOR U57333 ( .A(n44866), .B(n44867), .Z(n48267) );
  XOR U57334 ( .A(n47860), .B(n48267), .Z(n44347) );
  IV U57335 ( .A(n44347), .Z(n47863) );
  IV U57336 ( .A(n44348), .Z(n44350) );
  NOR U57337 ( .A(n44350), .B(n44349), .Z(n47861) );
  XOR U57338 ( .A(n47863), .B(n47861), .Z(n44864) );
  IV U57339 ( .A(n44864), .Z(n44358) );
  IV U57340 ( .A(n44351), .Z(n44352) );
  NOR U57341 ( .A(n44353), .B(n44352), .Z(n44863) );
  IV U57342 ( .A(n44354), .Z(n44356) );
  NOR U57343 ( .A(n44356), .B(n44355), .Z(n44861) );
  NOR U57344 ( .A(n44863), .B(n44861), .Z(n44357) );
  XOR U57345 ( .A(n44358), .B(n44357), .Z(n44856) );
  XOR U57346 ( .A(n44855), .B(n44856), .Z(n44860) );
  XOR U57347 ( .A(n44858), .B(n44860), .Z(n44851) );
  XOR U57348 ( .A(n44849), .B(n44851), .Z(n44853) );
  XOR U57349 ( .A(n44359), .B(n44853), .Z(n44360) );
  IV U57350 ( .A(n44360), .Z(n44842) );
  XOR U57351 ( .A(n44841), .B(n44842), .Z(n44846) );
  IV U57352 ( .A(n44361), .Z(n44363) );
  NOR U57353 ( .A(n44363), .B(n44362), .Z(n44844) );
  XOR U57354 ( .A(n44846), .B(n44844), .Z(n47870) );
  XOR U57355 ( .A(n47871), .B(n47870), .Z(n44838) );
  IV U57356 ( .A(n44364), .Z(n44369) );
  IV U57357 ( .A(n44365), .Z(n44366) );
  NOR U57358 ( .A(n44369), .B(n44366), .Z(n47872) );
  IV U57359 ( .A(n44367), .Z(n44368) );
  NOR U57360 ( .A(n44369), .B(n44368), .Z(n44839) );
  NOR U57361 ( .A(n47872), .B(n44839), .Z(n44370) );
  XOR U57362 ( .A(n44838), .B(n44370), .Z(n44837) );
  IV U57363 ( .A(n44371), .Z(n44374) );
  IV U57364 ( .A(n44372), .Z(n44373) );
  NOR U57365 ( .A(n44374), .B(n44373), .Z(n44835) );
  XOR U57366 ( .A(n44837), .B(n44835), .Z(n44833) );
  NOR U57367 ( .A(n44381), .B(n44833), .Z(n48244) );
  IV U57368 ( .A(n44375), .Z(n44376) );
  NOR U57369 ( .A(n44376), .B(n44387), .Z(n44377) );
  IV U57370 ( .A(n44377), .Z(n44831) );
  IV U57371 ( .A(n44378), .Z(n44379) );
  NOR U57372 ( .A(n44380), .B(n44379), .Z(n44832) );
  XOR U57373 ( .A(n44832), .B(n44833), .Z(n44830) );
  XOR U57374 ( .A(n44831), .B(n44830), .Z(n44384) );
  IV U57375 ( .A(n44830), .Z(n44382) );
  NOR U57376 ( .A(n44382), .B(n44381), .Z(n44383) );
  NOR U57377 ( .A(n44384), .B(n44383), .Z(n44385) );
  NOR U57378 ( .A(n48244), .B(n44385), .Z(n47879) );
  IV U57379 ( .A(n44386), .Z(n44388) );
  NOR U57380 ( .A(n44388), .B(n44387), .Z(n44389) );
  IV U57381 ( .A(n44389), .Z(n47880) );
  XOR U57382 ( .A(n47879), .B(n47880), .Z(n48241) );
  IV U57383 ( .A(n48241), .Z(n44396) );
  IV U57384 ( .A(n44390), .Z(n44391) );
  NOR U57385 ( .A(n44392), .B(n44391), .Z(n51279) );
  IV U57386 ( .A(n44393), .Z(n44395) );
  NOR U57387 ( .A(n44395), .B(n44394), .Z(n48239) );
  NOR U57388 ( .A(n51279), .B(n48239), .Z(n47882) );
  XOR U57389 ( .A(n44396), .B(n47882), .Z(n47894) );
  XOR U57390 ( .A(n47893), .B(n47894), .Z(n47887) );
  XOR U57391 ( .A(n47886), .B(n47887), .Z(n47891) );
  XOR U57392 ( .A(n47890), .B(n47891), .Z(n44827) );
  XOR U57393 ( .A(n44826), .B(n44827), .Z(n47907) );
  XOR U57394 ( .A(n47906), .B(n47907), .Z(n44825) );
  XOR U57395 ( .A(n44824), .B(n44825), .Z(n44399) );
  IV U57396 ( .A(n44399), .Z(n44397) );
  NOR U57397 ( .A(n44398), .B(n44397), .Z(n48231) );
  NOR U57398 ( .A(n44400), .B(n44399), .Z(n44818) );
  XOR U57399 ( .A(n44818), .B(n44816), .Z(n44401) );
  NOR U57400 ( .A(n48231), .B(n44401), .Z(n44813) );
  XOR U57401 ( .A(n44402), .B(n44813), .Z(n44812) );
  XOR U57402 ( .A(n44810), .B(n44812), .Z(n44805) );
  XOR U57403 ( .A(n44804), .B(n44805), .Z(n44808) );
  XOR U57404 ( .A(n44807), .B(n44808), .Z(n44802) );
  NOR U57405 ( .A(n44403), .B(n44802), .Z(n48224) );
  IV U57406 ( .A(n44404), .Z(n44406) );
  NOR U57407 ( .A(n44406), .B(n44405), .Z(n44801) );
  XOR U57408 ( .A(n44801), .B(n44802), .Z(n44412) );
  IV U57409 ( .A(n44412), .Z(n44407) );
  NOR U57410 ( .A(n44408), .B(n44407), .Z(n44409) );
  NOR U57411 ( .A(n48224), .B(n44409), .Z(n44410) );
  NOR U57412 ( .A(n44411), .B(n44410), .Z(n44414) );
  IV U57413 ( .A(n44411), .Z(n44413) );
  NOR U57414 ( .A(n44413), .B(n44412), .Z(n44800) );
  NOR U57415 ( .A(n44414), .B(n44800), .Z(n44432) );
  IV U57416 ( .A(n44432), .Z(n44798) );
  IV U57417 ( .A(n44415), .Z(n44417) );
  NOR U57418 ( .A(n44417), .B(n44416), .Z(n44418) );
  IV U57419 ( .A(n44418), .Z(n44423) );
  NOR U57420 ( .A(n44420), .B(n44419), .Z(n44421) );
  IV U57421 ( .A(n44421), .Z(n44422) );
  NOR U57422 ( .A(n44423), .B(n44422), .Z(n44434) );
  IV U57423 ( .A(n44434), .Z(n44424) );
  NOR U57424 ( .A(n44798), .B(n44424), .Z(n48217) );
  IV U57425 ( .A(n44425), .Z(n44426) );
  NOR U57426 ( .A(n44426), .B(n44430), .Z(n44427) );
  IV U57427 ( .A(n44427), .Z(n44795) );
  IV U57428 ( .A(n44428), .Z(n44429) );
  NOR U57429 ( .A(n44430), .B(n44429), .Z(n44431) );
  IV U57430 ( .A(n44431), .Z(n44797) );
  XOR U57431 ( .A(n44432), .B(n44797), .Z(n44796) );
  XOR U57432 ( .A(n44795), .B(n44796), .Z(n44433) );
  NOR U57433 ( .A(n44434), .B(n44433), .Z(n44435) );
  NOR U57434 ( .A(n48217), .B(n44435), .Z(n44792) );
  XOR U57435 ( .A(n44436), .B(n44792), .Z(n48210) );
  XOR U57436 ( .A(n47926), .B(n48210), .Z(n44789) );
  XOR U57437 ( .A(n44791), .B(n44789), .Z(n48205) );
  XOR U57438 ( .A(n44437), .B(n48205), .Z(n44786) );
  IV U57439 ( .A(n44438), .Z(n44439) );
  NOR U57440 ( .A(n44439), .B(n44442), .Z(n44440) );
  IV U57441 ( .A(n44440), .Z(n44787) );
  XOR U57442 ( .A(n44786), .B(n44787), .Z(n44783) );
  IV U57443 ( .A(n44441), .Z(n44443) );
  NOR U57444 ( .A(n44443), .B(n44442), .Z(n44781) );
  XOR U57445 ( .A(n44783), .B(n44781), .Z(n47938) );
  IV U57446 ( .A(n44444), .Z(n44445) );
  NOR U57447 ( .A(n44448), .B(n44445), .Z(n47936) );
  XOR U57448 ( .A(n47938), .B(n47936), .Z(n47941) );
  IV U57449 ( .A(n44446), .Z(n44447) );
  NOR U57450 ( .A(n44448), .B(n44447), .Z(n47939) );
  XOR U57451 ( .A(n47941), .B(n47939), .Z(n47944) );
  XOR U57452 ( .A(n47943), .B(n47944), .Z(n47948) );
  IV U57453 ( .A(n44449), .Z(n44453) );
  IV U57454 ( .A(n44450), .Z(n44451) );
  NOR U57455 ( .A(n44453), .B(n44451), .Z(n47946) );
  XOR U57456 ( .A(n47948), .B(n47946), .Z(n47952) );
  IV U57457 ( .A(n44452), .Z(n44456) );
  NOR U57458 ( .A(n44454), .B(n44453), .Z(n44455) );
  IV U57459 ( .A(n44455), .Z(n44458) );
  NOR U57460 ( .A(n44456), .B(n44458), .Z(n47950) );
  XOR U57461 ( .A(n47952), .B(n47950), .Z(n47955) );
  IV U57462 ( .A(n44457), .Z(n44459) );
  NOR U57463 ( .A(n44459), .B(n44458), .Z(n47953) );
  XOR U57464 ( .A(n47955), .B(n47953), .Z(n47959) );
  NOR U57465 ( .A(n44461), .B(n44460), .Z(n44462) );
  IV U57466 ( .A(n44462), .Z(n44467) );
  NOR U57467 ( .A(n44464), .B(n44463), .Z(n44465) );
  IV U57468 ( .A(n44465), .Z(n44466) );
  NOR U57469 ( .A(n44467), .B(n44466), .Z(n47957) );
  XOR U57470 ( .A(n47959), .B(n47957), .Z(n47961) );
  XOR U57471 ( .A(n47960), .B(n47961), .Z(n47965) );
  XOR U57472 ( .A(n47964), .B(n47965), .Z(n47972) );
  IV U57473 ( .A(n47972), .Z(n44475) );
  IV U57474 ( .A(n44468), .Z(n44469) );
  NOR U57475 ( .A(n44470), .B(n44469), .Z(n47967) );
  IV U57476 ( .A(n44471), .Z(n44472) );
  NOR U57477 ( .A(n44473), .B(n44472), .Z(n47970) );
  NOR U57478 ( .A(n47967), .B(n47970), .Z(n44474) );
  XOR U57479 ( .A(n44475), .B(n44474), .Z(n47975) );
  XOR U57480 ( .A(n47973), .B(n47975), .Z(n47979) );
  XOR U57481 ( .A(n47977), .B(n47979), .Z(n48164) );
  XOR U57482 ( .A(n47980), .B(n48164), .Z(n44476) );
  IV U57483 ( .A(n44476), .Z(n44776) );
  XOR U57484 ( .A(n44775), .B(n44776), .Z(n44780) );
  IV U57485 ( .A(n44477), .Z(n44483) );
  IV U57486 ( .A(n44478), .Z(n44480) );
  NOR U57487 ( .A(n44480), .B(n44479), .Z(n44481) );
  IV U57488 ( .A(n44481), .Z(n44482) );
  NOR U57489 ( .A(n44483), .B(n44482), .Z(n44778) );
  XOR U57490 ( .A(n44780), .B(n44778), .Z(n47985) );
  XOR U57491 ( .A(n47984), .B(n47985), .Z(n47988) );
  IV U57492 ( .A(n47988), .Z(n44490) );
  NOR U57493 ( .A(n44485), .B(n44484), .Z(n47987) );
  IV U57494 ( .A(n44486), .Z(n44487) );
  NOR U57495 ( .A(n44488), .B(n44487), .Z(n44770) );
  NOR U57496 ( .A(n47987), .B(n44770), .Z(n44489) );
  XOR U57497 ( .A(n44490), .B(n44489), .Z(n44773) );
  XOR U57498 ( .A(n44772), .B(n44773), .Z(n44766) );
  XOR U57499 ( .A(n44764), .B(n44766), .Z(n44768) );
  XOR U57500 ( .A(n44767), .B(n44768), .Z(n44760) );
  XOR U57501 ( .A(n44758), .B(n44760), .Z(n44763) );
  XOR U57502 ( .A(n44761), .B(n44763), .Z(n44753) );
  XOR U57503 ( .A(n44752), .B(n44753), .Z(n44756) );
  XOR U57504 ( .A(n44755), .B(n44756), .Z(n44747) );
  XOR U57505 ( .A(n44746), .B(n44747), .Z(n44750) );
  XOR U57506 ( .A(n44749), .B(n44750), .Z(n47995) );
  XOR U57507 ( .A(n47993), .B(n47995), .Z(n47997) );
  XOR U57508 ( .A(n47996), .B(n47997), .Z(n44741) );
  XOR U57509 ( .A(n44740), .B(n44741), .Z(n44744) );
  XOR U57510 ( .A(n44491), .B(n44744), .Z(n44729) );
  XOR U57511 ( .A(n44492), .B(n44729), .Z(n44733) );
  XOR U57512 ( .A(n44493), .B(n44733), .Z(n44494) );
  IV U57513 ( .A(n44494), .Z(n48006) );
  XOR U57514 ( .A(n48004), .B(n48006), .Z(n48008) );
  XOR U57515 ( .A(n48007), .B(n48008), .Z(n48013) );
  IV U57516 ( .A(n48013), .Z(n44502) );
  IV U57517 ( .A(n44495), .Z(n44496) );
  NOR U57518 ( .A(n44497), .B(n44496), .Z(n48012) );
  IV U57519 ( .A(n44498), .Z(n44500) );
  NOR U57520 ( .A(n44500), .B(n44499), .Z(n44725) );
  NOR U57521 ( .A(n48012), .B(n44725), .Z(n44501) );
  XOR U57522 ( .A(n44502), .B(n44501), .Z(n44724) );
  XOR U57523 ( .A(n44722), .B(n44724), .Z(n51427) );
  XOR U57524 ( .A(n48017), .B(n51427), .Z(n44719) );
  IV U57525 ( .A(n44503), .Z(n44504) );
  NOR U57526 ( .A(n44505), .B(n44504), .Z(n44506) );
  IV U57527 ( .A(n44506), .Z(n44720) );
  XOR U57528 ( .A(n44719), .B(n44720), .Z(n48025) );
  XOR U57529 ( .A(n48022), .B(n48025), .Z(n44718) );
  NOR U57530 ( .A(n44507), .B(n48026), .Z(n44511) );
  IV U57531 ( .A(n44508), .Z(n44517) );
  IV U57532 ( .A(n44509), .Z(n44510) );
  NOR U57533 ( .A(n44517), .B(n44510), .Z(n44716) );
  NOR U57534 ( .A(n44511), .B(n44716), .Z(n44512) );
  XOR U57535 ( .A(n44718), .B(n44512), .Z(n44710) );
  IV U57536 ( .A(n44513), .Z(n44514) );
  NOR U57537 ( .A(n44515), .B(n44514), .Z(n44711) );
  IV U57538 ( .A(n44516), .Z(n44518) );
  NOR U57539 ( .A(n44518), .B(n44517), .Z(n44713) );
  NOR U57540 ( .A(n44711), .B(n44713), .Z(n44519) );
  XOR U57541 ( .A(n44710), .B(n44519), .Z(n48136) );
  XOR U57542 ( .A(n44705), .B(n48136), .Z(n44706) );
  XOR U57543 ( .A(n44707), .B(n44706), .Z(n44704) );
  XOR U57544 ( .A(n44702), .B(n44704), .Z(n48126) );
  XOR U57545 ( .A(n48035), .B(n48126), .Z(n48037) );
  NOR U57546 ( .A(n44521), .B(n44520), .Z(n48036) );
  NOR U57547 ( .A(n44523), .B(n44522), .Z(n48041) );
  NOR U57548 ( .A(n48036), .B(n48041), .Z(n44524) );
  XOR U57549 ( .A(n48037), .B(n44524), .Z(n48045) );
  NOR U57550 ( .A(n44525), .B(n48045), .Z(n54899) );
  IV U57551 ( .A(n44531), .Z(n44528) );
  NOR U57552 ( .A(n44527), .B(n44526), .Z(n48044) );
  XOR U57553 ( .A(n48044), .B(n48045), .Z(n44529) );
  NOR U57554 ( .A(n44528), .B(n44529), .Z(n51530) );
  NOR U57555 ( .A(n54899), .B(n51530), .Z(n51489) );
  IV U57556 ( .A(n51489), .Z(n48047) );
  NOR U57557 ( .A(n48047), .B(n44529), .Z(n44534) );
  NOR U57558 ( .A(n44531), .B(n44530), .Z(n44532) );
  NOR U57559 ( .A(n44532), .B(n48047), .Z(n44533) );
  NOR U57560 ( .A(n44534), .B(n44533), .Z(n44536) );
  NOR U57561 ( .A(n44535), .B(n44536), .Z(n51494) );
  IV U57562 ( .A(n44536), .Z(n44537) );
  NOR U57563 ( .A(n44538), .B(n44537), .Z(n44696) );
  NOR U57564 ( .A(n44540), .B(n44539), .Z(n44541) );
  XOR U57565 ( .A(n44542), .B(n44541), .Z(n44629) );
  IV U57566 ( .A(n44543), .Z(n44545) );
  NOR U57567 ( .A(n44545), .B(n44544), .Z(n44546) );
  XOR U57568 ( .A(n44547), .B(n44546), .Z(n44548) );
  NOR U57569 ( .A(n44571), .B(n44548), .Z(n44549) );
  NOR U57570 ( .A(n44566), .B(n44549), .Z(n44567) );
  IV U57571 ( .A(n44567), .Z(n44608) );
  NOR U57572 ( .A(n44551), .B(n44550), .Z(n44552) );
  XOR U57573 ( .A(n44553), .B(n44552), .Z(n44568) );
  IV U57574 ( .A(n44568), .Z(n44558) );
  IV U57575 ( .A(n44554), .Z(n44556) );
  NOR U57576 ( .A(n44556), .B(n44555), .Z(n44601) );
  IV U57577 ( .A(n44601), .Z(n44557) );
  NOR U57578 ( .A(n44558), .B(n44557), .Z(n44603) );
  IV U57579 ( .A(n44603), .Z(n44559) );
  NOR U57580 ( .A(n44608), .B(n44559), .Z(n44593) );
  IV U57581 ( .A(n44593), .Z(n44560) );
  NOR U57582 ( .A(n44565), .B(n44560), .Z(n44578) );
  IV U57583 ( .A(n44578), .Z(n44561) );
  NOR U57584 ( .A(n44562), .B(n44561), .Z(n44628) );
  IV U57585 ( .A(n44628), .Z(n44563) );
  NOR U57586 ( .A(n44629), .B(n44563), .Z(n44694) );
  XOR U57587 ( .A(n44696), .B(n44694), .Z(n44564) );
  NOR U57588 ( .A(n51494), .B(n44564), .Z(n44687) );
  XOR U57589 ( .A(n44566), .B(n44565), .Z(n44595) );
  XOR U57590 ( .A(n44567), .B(n44603), .Z(n44657) );
  IV U57591 ( .A(n44657), .Z(n44624) );
  NOR U57592 ( .A(n44569), .B(n44568), .Z(n44570) );
  NOR U57593 ( .A(n44571), .B(n44570), .Z(n44600) );
  IV U57594 ( .A(n44600), .Z(n44576) );
  IV U57595 ( .A(n44572), .Z(n44574) );
  NOR U57596 ( .A(n44574), .B(n44573), .Z(n44619) );
  IV U57597 ( .A(n44619), .Z(n44575) );
  NOR U57598 ( .A(n44576), .B(n44575), .Z(n44639) );
  IV U57599 ( .A(n44639), .Z(n44658) );
  NOR U57600 ( .A(n44624), .B(n44658), .Z(n44592) );
  IV U57601 ( .A(n44592), .Z(n44577) );
  NOR U57602 ( .A(n44595), .B(n44577), .Z(n44591) );
  IV U57603 ( .A(n44591), .Z(n44588) );
  NOR U57604 ( .A(n44579), .B(n44578), .Z(n44580) );
  IV U57605 ( .A(n44580), .Z(n44585) );
  IV U57606 ( .A(n44581), .Z(n44582) );
  NOR U57607 ( .A(n44583), .B(n44582), .Z(n44584) );
  NOR U57608 ( .A(n44585), .B(n44584), .Z(n44587) );
  XOR U57609 ( .A(n44587), .B(n44586), .Z(n44590) );
  NOR U57610 ( .A(n44588), .B(n44590), .Z(n44627) );
  IV U57611 ( .A(n44627), .Z(n44589) );
  NOR U57612 ( .A(n44629), .B(n44589), .Z(n44698) );
  XOR U57613 ( .A(n44591), .B(n44590), .Z(n44611) );
  NOR U57614 ( .A(n44593), .B(n44592), .Z(n44594) );
  XOR U57615 ( .A(n44595), .B(n44594), .Z(n44596) );
  IV U57616 ( .A(n44596), .Z(n44614) );
  IV U57617 ( .A(n44597), .Z(n44599) );
  NOR U57618 ( .A(n44599), .B(n44598), .Z(n44636) );
  IV U57619 ( .A(n44636), .Z(n44605) );
  NOR U57620 ( .A(n44601), .B(n44600), .Z(n44602) );
  NOR U57621 ( .A(n44603), .B(n44602), .Z(n44618) );
  IV U57622 ( .A(n44618), .Z(n44604) );
  NOR U57623 ( .A(n44605), .B(n44604), .Z(n44606) );
  IV U57624 ( .A(n44606), .Z(n44607) );
  NOR U57625 ( .A(n44608), .B(n44607), .Z(n44613) );
  IV U57626 ( .A(n44613), .Z(n44609) );
  NOR U57627 ( .A(n44614), .B(n44609), .Z(n44610) );
  IV U57628 ( .A(n44610), .Z(n44612) );
  NOR U57629 ( .A(n44611), .B(n44612), .Z(n44691) );
  XOR U57630 ( .A(n44612), .B(n44611), .Z(n48085) );
  IV U57631 ( .A(n48085), .Z(n44655) );
  XOR U57632 ( .A(n44614), .B(n44613), .Z(n44654) );
  IV U57633 ( .A(n44615), .Z(n44617) );
  NOR U57634 ( .A(n44617), .B(n44616), .Z(n44635) );
  IV U57635 ( .A(n44635), .Z(n44621) );
  NOR U57636 ( .A(n44619), .B(n44618), .Z(n44620) );
  NOR U57637 ( .A(n44639), .B(n44620), .Z(n44642) );
  IV U57638 ( .A(n44642), .Z(n44637) );
  NOR U57639 ( .A(n44621), .B(n44637), .Z(n44622) );
  IV U57640 ( .A(n44622), .Z(n44623) );
  NOR U57641 ( .A(n44624), .B(n44623), .Z(n44625) );
  IV U57642 ( .A(n44625), .Z(n44652) );
  NOR U57643 ( .A(n44654), .B(n44652), .Z(n44626) );
  IV U57644 ( .A(n44626), .Z(n44649) );
  NOR U57645 ( .A(n44655), .B(n44649), .Z(n44686) );
  NOR U57646 ( .A(n44691), .B(n44686), .Z(n44634) );
  NOR U57647 ( .A(n44628), .B(n44627), .Z(n44630) );
  XOR U57648 ( .A(n44630), .B(n44629), .Z(n44633) );
  IV U57649 ( .A(n44633), .Z(n44688) );
  NOR U57650 ( .A(n44634), .B(n44688), .Z(n44631) );
  NOR U57651 ( .A(n44698), .B(n44631), .Z(n44632) );
  XOR U57652 ( .A(n44687), .B(n44632), .Z(n48054) );
  XOR U57653 ( .A(n44634), .B(n44633), .Z(n48057) );
  NOR U57654 ( .A(n44636), .B(n44635), .Z(n44641) );
  NOR U57655 ( .A(n44641), .B(n44637), .Z(n44638) );
  NOR U57656 ( .A(n44639), .B(n44638), .Z(n44640) );
  XOR U57657 ( .A(n44657), .B(n44640), .Z(n44667) );
  XOR U57658 ( .A(n44642), .B(n44641), .Z(n44672) );
  IV U57659 ( .A(n44643), .Z(n44645) );
  NOR U57660 ( .A(n44645), .B(n44644), .Z(n44674) );
  IV U57661 ( .A(n44674), .Z(n44646) );
  NOR U57662 ( .A(n44672), .B(n44646), .Z(n44647) );
  IV U57663 ( .A(n44647), .Z(n44668) );
  NOR U57664 ( .A(n44667), .B(n44668), .Z(n44648) );
  IV U57665 ( .A(n44648), .Z(n44651) );
  NOR U57666 ( .A(n44654), .B(n44651), .Z(n48061) );
  IV U57667 ( .A(n48061), .Z(n44650) );
  XOR U57668 ( .A(n44649), .B(n48085), .Z(n48060) );
  NOR U57669 ( .A(n44650), .B(n48060), .Z(n48050) );
  XOR U57670 ( .A(n44652), .B(n44651), .Z(n44653) );
  XOR U57671 ( .A(n44654), .B(n44653), .Z(n48082) );
  NOR U57672 ( .A(n44655), .B(n48082), .Z(n44656) );
  IV U57673 ( .A(n44656), .Z(n44683) );
  XOR U57674 ( .A(n44658), .B(n44657), .Z(n44664) );
  IV U57675 ( .A(n44659), .Z(n44661) );
  NOR U57676 ( .A(n44661), .B(n44660), .Z(n44673) );
  IV U57677 ( .A(n44673), .Z(n44662) );
  NOR U57678 ( .A(n44672), .B(n44662), .Z(n44670) );
  IV U57679 ( .A(n44670), .Z(n44663) );
  NOR U57680 ( .A(n44664), .B(n44663), .Z(n48063) );
  IV U57681 ( .A(n48063), .Z(n44665) );
  NOR U57682 ( .A(n44683), .B(n44665), .Z(n48055) );
  NOR U57683 ( .A(n48050), .B(n48055), .Z(n44666) );
  XOR U57684 ( .A(n48057), .B(n44666), .Z(n48104) );
  IV U57685 ( .A(n48104), .Z(n48073) );
  XOR U57686 ( .A(n44668), .B(n44667), .Z(n44669) );
  NOR U57687 ( .A(n44670), .B(n44669), .Z(n44671) );
  NOR U57688 ( .A(n48063), .B(n44671), .Z(n54941) );
  IV U57689 ( .A(n54941), .Z(n48097) );
  IV U57690 ( .A(n44672), .Z(n44676) );
  NOR U57691 ( .A(n44674), .B(n44673), .Z(n44675) );
  XOR U57692 ( .A(n44676), .B(n44675), .Z(n48090) );
  IV U57693 ( .A(n44677), .Z(n44679) );
  NOR U57694 ( .A(n44679), .B(n44678), .Z(n48091) );
  IV U57695 ( .A(n48091), .Z(n44680) );
  NOR U57696 ( .A(n48090), .B(n44680), .Z(n54939) );
  IV U57697 ( .A(n54939), .Z(n44681) );
  NOR U57698 ( .A(n48097), .B(n44681), .Z(n48062) );
  IV U57699 ( .A(n48062), .Z(n44682) );
  NOR U57700 ( .A(n44683), .B(n44682), .Z(n48103) );
  IV U57701 ( .A(n48103), .Z(n44684) );
  NOR U57702 ( .A(n48073), .B(n44684), .Z(n44685) );
  IV U57703 ( .A(n44685), .Z(n48077) );
  NOR U57704 ( .A(n48054), .B(n48077), .Z(n48111) );
  IV U57705 ( .A(n44686), .Z(n44690) );
  IV U57706 ( .A(n44687), .Z(n44700) );
  NOR U57707 ( .A(n44700), .B(n44688), .Z(n44689) );
  IV U57708 ( .A(n44689), .Z(n44692) );
  NOR U57709 ( .A(n44690), .B(n44692), .Z(n51500) );
  IV U57710 ( .A(n44691), .Z(n44693) );
  NOR U57711 ( .A(n44693), .B(n44692), .Z(n48114) );
  IV U57712 ( .A(n44694), .Z(n44695) );
  NOR U57713 ( .A(n44696), .B(n44695), .Z(n48119) );
  NOR U57714 ( .A(n51494), .B(n48119), .Z(n44697) );
  IV U57715 ( .A(n44697), .Z(n44701) );
  IV U57716 ( .A(n44698), .Z(n44699) );
  NOR U57717 ( .A(n44700), .B(n44699), .Z(n48117) );
  NOR U57718 ( .A(n44701), .B(n48117), .Z(n48048) );
  IV U57719 ( .A(n44702), .Z(n44703) );
  NOR U57720 ( .A(n44704), .B(n44703), .Z(n48129) );
  NOR U57721 ( .A(n44705), .B(n48136), .Z(n44709) );
  IV U57722 ( .A(n44706), .Z(n44708) );
  NOR U57723 ( .A(n44708), .B(n44707), .Z(n48132) );
  NOR U57724 ( .A(n44709), .B(n48132), .Z(n48033) );
  IV U57725 ( .A(n44710), .Z(n44715) );
  IV U57726 ( .A(n44711), .Z(n44712) );
  NOR U57727 ( .A(n44715), .B(n44712), .Z(n51464) );
  IV U57728 ( .A(n44713), .Z(n44714) );
  NOR U57729 ( .A(n44715), .B(n44714), .Z(n51468) );
  IV U57730 ( .A(n44716), .Z(n44717) );
  NOR U57731 ( .A(n44718), .B(n44717), .Z(n51455) );
  IV U57732 ( .A(n44719), .Z(n44721) );
  NOR U57733 ( .A(n44721), .B(n44720), .Z(n48020) );
  IV U57734 ( .A(n48020), .Z(n48016) );
  IV U57735 ( .A(n44722), .Z(n44723) );
  NOR U57736 ( .A(n44724), .B(n44723), .Z(n51431) );
  IV U57737 ( .A(n44725), .Z(n44726) );
  NOR U57738 ( .A(n44726), .B(n48013), .Z(n51421) );
  IV U57739 ( .A(n44727), .Z(n44728) );
  NOR U57740 ( .A(n44728), .B(n44733), .Z(n48144) );
  IV U57741 ( .A(n44729), .Z(n44737) );
  IV U57742 ( .A(n44730), .Z(n44731) );
  NOR U57743 ( .A(n44737), .B(n44731), .Z(n48152) );
  IV U57744 ( .A(n44732), .Z(n44734) );
  NOR U57745 ( .A(n44734), .B(n44733), .Z(n48149) );
  NOR U57746 ( .A(n48152), .B(n48149), .Z(n48003) );
  IV U57747 ( .A(n44735), .Z(n44736) );
  NOR U57748 ( .A(n44737), .B(n44736), .Z(n51410) );
  IV U57749 ( .A(n44738), .Z(n44739) );
  NOR U57750 ( .A(n44739), .B(n44744), .Z(n51406) );
  NOR U57751 ( .A(n51410), .B(n51406), .Z(n48002) );
  IV U57752 ( .A(n44740), .Z(n44742) );
  NOR U57753 ( .A(n44742), .B(n44741), .Z(n51399) );
  IV U57754 ( .A(n44743), .Z(n44745) );
  NOR U57755 ( .A(n44745), .B(n44744), .Z(n51403) );
  NOR U57756 ( .A(n51399), .B(n51403), .Z(n48001) );
  IV U57757 ( .A(n44746), .Z(n44748) );
  NOR U57758 ( .A(n44748), .B(n44747), .Z(n51597) );
  IV U57759 ( .A(n44749), .Z(n44751) );
  NOR U57760 ( .A(n44751), .B(n44750), .Z(n51591) );
  NOR U57761 ( .A(n51597), .B(n51591), .Z(n51389) );
  IV U57762 ( .A(n44752), .Z(n44754) );
  NOR U57763 ( .A(n44754), .B(n44753), .Z(n48157) );
  IV U57764 ( .A(n44755), .Z(n44757) );
  NOR U57765 ( .A(n44757), .B(n44756), .Z(n51390) );
  NOR U57766 ( .A(n48157), .B(n51390), .Z(n47992) );
  IV U57767 ( .A(n44758), .Z(n44759) );
  NOR U57768 ( .A(n44760), .B(n44759), .Z(n51385) );
  IV U57769 ( .A(n44761), .Z(n44762) );
  NOR U57770 ( .A(n44763), .B(n44762), .Z(n48159) );
  NOR U57771 ( .A(n51385), .B(n48159), .Z(n47991) );
  IV U57772 ( .A(n44764), .Z(n44765) );
  NOR U57773 ( .A(n44766), .B(n44765), .Z(n51621) );
  IV U57774 ( .A(n44767), .Z(n44769) );
  NOR U57775 ( .A(n44769), .B(n44768), .Z(n51616) );
  NOR U57776 ( .A(n51621), .B(n51616), .Z(n51378) );
  IV U57777 ( .A(n44770), .Z(n44771) );
  NOR U57778 ( .A(n44771), .B(n47988), .Z(n51374) );
  IV U57779 ( .A(n44772), .Z(n44774) );
  NOR U57780 ( .A(n44774), .B(n44773), .Z(n51379) );
  NOR U57781 ( .A(n51374), .B(n51379), .Z(n47990) );
  IV U57782 ( .A(n44775), .Z(n44777) );
  NOR U57783 ( .A(n44777), .B(n44776), .Z(n51356) );
  IV U57784 ( .A(n44778), .Z(n44779) );
  NOR U57785 ( .A(n44780), .B(n44779), .Z(n51358) );
  NOR U57786 ( .A(n51356), .B(n51358), .Z(n47983) );
  IV U57787 ( .A(n44781), .Z(n44782) );
  NOR U57788 ( .A(n44783), .B(n44782), .Z(n51326) );
  IV U57789 ( .A(n44784), .Z(n44785) );
  NOR U57790 ( .A(n44785), .B(n48205), .Z(n51657) );
  IV U57791 ( .A(n44786), .Z(n44788) );
  NOR U57792 ( .A(n44788), .B(n44787), .Z(n51652) );
  NOR U57793 ( .A(n51657), .B(n51652), .Z(n48191) );
  IV U57794 ( .A(n44789), .Z(n44790) );
  NOR U57795 ( .A(n44791), .B(n44790), .Z(n47930) );
  IV U57796 ( .A(n47930), .Z(n47925) );
  IV U57797 ( .A(n44792), .Z(n47922) );
  IV U57798 ( .A(n44793), .Z(n44794) );
  NOR U57799 ( .A(n47922), .B(n44794), .Z(n51319) );
  NOR U57800 ( .A(n44796), .B(n44795), .Z(n51312) );
  NOR U57801 ( .A(n44798), .B(n44797), .Z(n44799) );
  NOR U57802 ( .A(n44800), .B(n44799), .Z(n51311) );
  IV U57803 ( .A(n44801), .Z(n44803) );
  NOR U57804 ( .A(n44803), .B(n44802), .Z(n48219) );
  NOR U57805 ( .A(n48224), .B(n48219), .Z(n47919) );
  IV U57806 ( .A(n44804), .Z(n44806) );
  NOR U57807 ( .A(n44806), .B(n44805), .Z(n51303) );
  IV U57808 ( .A(n44807), .Z(n44809) );
  NOR U57809 ( .A(n44809), .B(n44808), .Z(n48221) );
  NOR U57810 ( .A(n51303), .B(n48221), .Z(n47918) );
  IV U57811 ( .A(n44810), .Z(n44811) );
  NOR U57812 ( .A(n44812), .B(n44811), .Z(n51296) );
  IV U57813 ( .A(n44813), .Z(n44821) );
  IV U57814 ( .A(n44814), .Z(n44815) );
  NOR U57815 ( .A(n44821), .B(n44815), .Z(n51290) );
  NOR U57816 ( .A(n51296), .B(n51290), .Z(n47917) );
  IV U57817 ( .A(n44816), .Z(n44817) );
  NOR U57818 ( .A(n44818), .B(n44817), .Z(n48228) );
  NOR U57819 ( .A(n48231), .B(n48228), .Z(n44819) );
  IV U57820 ( .A(n44819), .Z(n44823) );
  IV U57821 ( .A(n44820), .Z(n44822) );
  NOR U57822 ( .A(n44822), .B(n44821), .Z(n51287) );
  NOR U57823 ( .A(n44823), .B(n51287), .Z(n47916) );
  NOR U57824 ( .A(n44825), .B(n44824), .Z(n47914) );
  IV U57825 ( .A(n47914), .Z(n47905) );
  IV U57826 ( .A(n44826), .Z(n44828) );
  NOR U57827 ( .A(n44828), .B(n44827), .Z(n44829) );
  IV U57828 ( .A(n44829), .Z(n48234) );
  NOR U57829 ( .A(n44831), .B(n44830), .Z(n51272) );
  IV U57830 ( .A(n44832), .Z(n44834) );
  NOR U57831 ( .A(n44834), .B(n44833), .Z(n48248) );
  NOR U57832 ( .A(n48248), .B(n48244), .Z(n47877) );
  IV U57833 ( .A(n44835), .Z(n44836) );
  NOR U57834 ( .A(n44837), .B(n44836), .Z(n48246) );
  IV U57835 ( .A(n44838), .Z(n47873) );
  IV U57836 ( .A(n44839), .Z(n44840) );
  NOR U57837 ( .A(n47873), .B(n44840), .Z(n51267) );
  IV U57838 ( .A(n44841), .Z(n44843) );
  NOR U57839 ( .A(n44843), .B(n44842), .Z(n51254) );
  IV U57840 ( .A(n44844), .Z(n44845) );
  NOR U57841 ( .A(n44846), .B(n44845), .Z(n51257) );
  NOR U57842 ( .A(n51254), .B(n51257), .Z(n47869) );
  IV U57843 ( .A(n44847), .Z(n44848) );
  NOR U57844 ( .A(n44853), .B(n44848), .Z(n51251) );
  IV U57845 ( .A(n44849), .Z(n44850) );
  NOR U57846 ( .A(n44851), .B(n44850), .Z(n51239) );
  IV U57847 ( .A(n44852), .Z(n44854) );
  NOR U57848 ( .A(n44854), .B(n44853), .Z(n48252) );
  NOR U57849 ( .A(n51239), .B(n48252), .Z(n47868) );
  IV U57850 ( .A(n44855), .Z(n44857) );
  NOR U57851 ( .A(n44857), .B(n44856), .Z(n48258) );
  IV U57852 ( .A(n44858), .Z(n44859) );
  NOR U57853 ( .A(n44860), .B(n44859), .Z(n51243) );
  NOR U57854 ( .A(n48258), .B(n51243), .Z(n47867) );
  IV U57855 ( .A(n44861), .Z(n44862) );
  NOR U57856 ( .A(n44862), .B(n44864), .Z(n48255) );
  IV U57857 ( .A(n44863), .Z(n44865) );
  NOR U57858 ( .A(n44865), .B(n44864), .Z(n48260) );
  IV U57859 ( .A(n44866), .Z(n44868) );
  NOR U57860 ( .A(n44868), .B(n44867), .Z(n51225) );
  IV U57861 ( .A(n44869), .Z(n44870) );
  NOR U57862 ( .A(n44873), .B(n44870), .Z(n51200) );
  IV U57863 ( .A(n44871), .Z(n44875) );
  NOR U57864 ( .A(n44873), .B(n44872), .Z(n44874) );
  IV U57865 ( .A(n44874), .Z(n47845) );
  NOR U57866 ( .A(n44875), .B(n47845), .Z(n51208) );
  IV U57867 ( .A(n44876), .Z(n44877) );
  NOR U57868 ( .A(n44877), .B(n44882), .Z(n51193) );
  IV U57869 ( .A(n44878), .Z(n51187) );
  NOR U57870 ( .A(n51187), .B(n44879), .Z(n44883) );
  IV U57871 ( .A(n44880), .Z(n44881) );
  NOR U57872 ( .A(n44882), .B(n44881), .Z(n48278) );
  NOR U57873 ( .A(n44883), .B(n48278), .Z(n47842) );
  IV U57874 ( .A(n44884), .Z(n44885) );
  NOR U57875 ( .A(n44885), .B(n44887), .Z(n51181) );
  IV U57876 ( .A(n44886), .Z(n44888) );
  NOR U57877 ( .A(n44888), .B(n44887), .Z(n51179) );
  IV U57878 ( .A(n44889), .Z(n44890) );
  NOR U57879 ( .A(n44890), .B(n47827), .Z(n54712) );
  IV U57880 ( .A(n44891), .Z(n44892) );
  NOR U57881 ( .A(n44893), .B(n44892), .Z(n44894) );
  IV U57882 ( .A(n44894), .Z(n51170) );
  IV U57883 ( .A(n44895), .Z(n44896) );
  NOR U57884 ( .A(n44897), .B(n44896), .Z(n47784) );
  IV U57885 ( .A(n47784), .Z(n47776) );
  IV U57886 ( .A(n44898), .Z(n44899) );
  NOR U57887 ( .A(n44899), .B(n44901), .Z(n47762) );
  IV U57888 ( .A(n44900), .Z(n44902) );
  NOR U57889 ( .A(n44902), .B(n44901), .Z(n54652) );
  IV U57890 ( .A(n44903), .Z(n44905) );
  NOR U57891 ( .A(n44905), .B(n44904), .Z(n51830) );
  NOR U57892 ( .A(n54652), .B(n51830), .Z(n48314) );
  IV U57893 ( .A(n44906), .Z(n44907) );
  NOR U57894 ( .A(n44908), .B(n44907), .Z(n44909) );
  IV U57895 ( .A(n44909), .Z(n47751) );
  IV U57896 ( .A(n44910), .Z(n47750) );
  IV U57897 ( .A(n44911), .Z(n44912) );
  NOR U57898 ( .A(n47750), .B(n44912), .Z(n48327) );
  IV U57899 ( .A(n44913), .Z(n44914) );
  NOR U57900 ( .A(n47750), .B(n44914), .Z(n48331) );
  IV U57901 ( .A(n44915), .Z(n44916) );
  NOR U57902 ( .A(n44917), .B(n44916), .Z(n48333) );
  NOR U57903 ( .A(n48331), .B(n48333), .Z(n47747) );
  IV U57904 ( .A(n44918), .Z(n44920) );
  NOR U57905 ( .A(n44920), .B(n44919), .Z(n48343) );
  NOR U57906 ( .A(n44922), .B(n44921), .Z(n48340) );
  NOR U57907 ( .A(n48343), .B(n48340), .Z(n47731) );
  IV U57908 ( .A(n44923), .Z(n44924) );
  NOR U57909 ( .A(n44925), .B(n44924), .Z(n48347) );
  IV U57910 ( .A(n44926), .Z(n44928) );
  NOR U57911 ( .A(n44928), .B(n44927), .Z(n44929) );
  NOR U57912 ( .A(n44930), .B(n44929), .Z(n48356) );
  NOR U57913 ( .A(n44932), .B(n44931), .Z(n51130) );
  NOR U57914 ( .A(n44934), .B(n44933), .Z(n51133) );
  IV U57915 ( .A(n44935), .Z(n44936) );
  NOR U57916 ( .A(n44936), .B(n44941), .Z(n51128) );
  NOR U57917 ( .A(n51133), .B(n51128), .Z(n47719) );
  IV U57918 ( .A(n44937), .Z(n44938) );
  NOR U57919 ( .A(n44939), .B(n44938), .Z(n48359) );
  IV U57920 ( .A(n44940), .Z(n44942) );
  NOR U57921 ( .A(n44942), .B(n44941), .Z(n48357) );
  NOR U57922 ( .A(n48359), .B(n48357), .Z(n47718) );
  NOR U57923 ( .A(n44944), .B(n44943), .Z(n51112) );
  IV U57924 ( .A(n44945), .Z(n44947) );
  NOR U57925 ( .A(n44947), .B(n44946), .Z(n51119) );
  NOR U57926 ( .A(n51112), .B(n51119), .Z(n47717) );
  IV U57927 ( .A(n44948), .Z(n44949) );
  NOR U57928 ( .A(n44950), .B(n44949), .Z(n51106) );
  NOR U57929 ( .A(n51106), .B(n48362), .Z(n47716) );
  IV U57930 ( .A(n44951), .Z(n44953) );
  NOR U57931 ( .A(n44953), .B(n44952), .Z(n51883) );
  IV U57932 ( .A(n44954), .Z(n44956) );
  NOR U57933 ( .A(n44956), .B(n44955), .Z(n51878) );
  NOR U57934 ( .A(n51883), .B(n51878), .Z(n51089) );
  IV U57935 ( .A(n44957), .Z(n44965) );
  IV U57936 ( .A(n44958), .Z(n44959) );
  NOR U57937 ( .A(n44965), .B(n44959), .Z(n51084) );
  IV U57938 ( .A(n44960), .Z(n44961) );
  NOR U57939 ( .A(n44962), .B(n44961), .Z(n48377) );
  NOR U57940 ( .A(n51084), .B(n48377), .Z(n47673) );
  IV U57941 ( .A(n44963), .Z(n44964) );
  NOR U57942 ( .A(n44965), .B(n44964), .Z(n51070) );
  IV U57943 ( .A(n44966), .Z(n44967) );
  NOR U57944 ( .A(n44967), .B(n44971), .Z(n48379) );
  NOR U57945 ( .A(n44969), .B(n44968), .Z(n51911) );
  IV U57946 ( .A(n44970), .Z(n44972) );
  NOR U57947 ( .A(n44972), .B(n44971), .Z(n51907) );
  NOR U57948 ( .A(n51911), .B(n51907), .Z(n51075) );
  IV U57949 ( .A(n44973), .Z(n44975) );
  NOR U57950 ( .A(n44975), .B(n44974), .Z(n48385) );
  IV U57951 ( .A(n44976), .Z(n48389) );
  NOR U57952 ( .A(n44977), .B(n48389), .Z(n44978) );
  NOR U57953 ( .A(n48385), .B(n44978), .Z(n44979) );
  IV U57954 ( .A(n44979), .Z(n44980) );
  NOR U57955 ( .A(n48383), .B(n44980), .Z(n47672) );
  IV U57956 ( .A(n44981), .Z(n44984) );
  NOR U57957 ( .A(n44982), .B(n47668), .Z(n44983) );
  IV U57958 ( .A(n44983), .Z(n44986) );
  NOR U57959 ( .A(n44984), .B(n44986), .Z(n51062) );
  IV U57960 ( .A(n44985), .Z(n44987) );
  NOR U57961 ( .A(n44987), .B(n44986), .Z(n51059) );
  IV U57962 ( .A(n44988), .Z(n44989) );
  NOR U57963 ( .A(n44990), .B(n44989), .Z(n51050) );
  IV U57964 ( .A(n44991), .Z(n44993) );
  NOR U57965 ( .A(n44993), .B(n44992), .Z(n51053) );
  NOR U57966 ( .A(n51050), .B(n51053), .Z(n47666) );
  IV U57967 ( .A(n44994), .Z(n44996) );
  IV U57968 ( .A(n44995), .Z(n47663) );
  NOR U57969 ( .A(n44996), .B(n47663), .Z(n51047) );
  IV U57970 ( .A(n44997), .Z(n45004) );
  IV U57971 ( .A(n44998), .Z(n44999) );
  NOR U57972 ( .A(n45004), .B(n44999), .Z(n48395) );
  IV U57973 ( .A(n45000), .Z(n45001) );
  NOR U57974 ( .A(n45004), .B(n45001), .Z(n48400) );
  NOR U57975 ( .A(n48395), .B(n48400), .Z(n47659) );
  IV U57976 ( .A(n45002), .Z(n45003) );
  NOR U57977 ( .A(n45004), .B(n45003), .Z(n48403) );
  IV U57978 ( .A(n45005), .Z(n45006) );
  NOR U57979 ( .A(n45006), .B(n47657), .Z(n51036) );
  IV U57980 ( .A(n45007), .Z(n45010) );
  NOR U57981 ( .A(n47640), .B(n45008), .Z(n45009) );
  IV U57982 ( .A(n45009), .Z(n47642) );
  NOR U57983 ( .A(n45010), .B(n47642), .Z(n51015) );
  IV U57984 ( .A(n45011), .Z(n45013) );
  NOR U57985 ( .A(n45013), .B(n45012), .Z(n45014) );
  IV U57986 ( .A(n45014), .Z(n48417) );
  IV U57987 ( .A(n45015), .Z(n45016) );
  NOR U57988 ( .A(n45016), .B(n45018), .Z(n51967) );
  IV U57989 ( .A(n45017), .Z(n45019) );
  NOR U57990 ( .A(n45019), .B(n45018), .Z(n51963) );
  NOR U57991 ( .A(n51967), .B(n51963), .Z(n48423) );
  IV U57992 ( .A(n45020), .Z(n45021) );
  NOR U57993 ( .A(n45022), .B(n45021), .Z(n51004) );
  IV U57994 ( .A(n45023), .Z(n45025) );
  NOR U57995 ( .A(n45025), .B(n45024), .Z(n51008) );
  NOR U57996 ( .A(n51004), .B(n51008), .Z(n47637) );
  IV U57997 ( .A(n45026), .Z(n45031) );
  IV U57998 ( .A(n45027), .Z(n45028) );
  NOR U57999 ( .A(n45031), .B(n45028), .Z(n51001) );
  IV U58000 ( .A(n45029), .Z(n45030) );
  NOR U58001 ( .A(n45031), .B(n45030), .Z(n45032) );
  IV U58002 ( .A(n45032), .Z(n48424) );
  IV U58003 ( .A(n45033), .Z(n45035) );
  NOR U58004 ( .A(n45035), .B(n45034), .Z(n45036) );
  IV U58005 ( .A(n45036), .Z(n50996) );
  XOR U58006 ( .A(n48424), .B(n50996), .Z(n45037) );
  NOR U58007 ( .A(n51001), .B(n45037), .Z(n47636) );
  IV U58008 ( .A(n45038), .Z(n45039) );
  NOR U58009 ( .A(n45042), .B(n45039), .Z(n50991) );
  IV U58010 ( .A(n45040), .Z(n45041) );
  NOR U58011 ( .A(n45042), .B(n45041), .Z(n50997) );
  NOR U58012 ( .A(n50991), .B(n50997), .Z(n47635) );
  IV U58013 ( .A(n45043), .Z(n45044) );
  NOR U58014 ( .A(n45044), .B(n45050), .Z(n45045) );
  IV U58015 ( .A(n45045), .Z(n50989) );
  IV U58016 ( .A(n45046), .Z(n45048) );
  NOR U58017 ( .A(n45048), .B(n45047), .Z(n48426) );
  IV U58018 ( .A(n45049), .Z(n45051) );
  NOR U58019 ( .A(n45051), .B(n45050), .Z(n50985) );
  NOR U58020 ( .A(n48426), .B(n50985), .Z(n47634) );
  IV U58021 ( .A(n45052), .Z(n45054) );
  NOR U58022 ( .A(n45054), .B(n45053), .Z(n48428) );
  IV U58023 ( .A(n45055), .Z(n45056) );
  NOR U58024 ( .A(n45056), .B(n48432), .Z(n52006) );
  NOR U58025 ( .A(n48428), .B(n52006), .Z(n47633) );
  IV U58026 ( .A(n45057), .Z(n45058) );
  NOR U58027 ( .A(n45059), .B(n45058), .Z(n45060) );
  IV U58028 ( .A(n45060), .Z(n47628) );
  IV U58029 ( .A(n45061), .Z(n45064) );
  NOR U58030 ( .A(n45062), .B(n45071), .Z(n45063) );
  IV U58031 ( .A(n45063), .Z(n45066) );
  NOR U58032 ( .A(n45064), .B(n45066), .Z(n48436) );
  IV U58033 ( .A(n45065), .Z(n45067) );
  NOR U58034 ( .A(n45067), .B(n45066), .Z(n45068) );
  IV U58035 ( .A(n45068), .Z(n48448) );
  IV U58036 ( .A(n45069), .Z(n45070) );
  NOR U58037 ( .A(n45071), .B(n45070), .Z(n45072) );
  IV U58038 ( .A(n45072), .Z(n47620) );
  IV U58039 ( .A(n45073), .Z(n45075) );
  NOR U58040 ( .A(n45075), .B(n45074), .Z(n50964) );
  IV U58041 ( .A(n45076), .Z(n45077) );
  NOR U58042 ( .A(n45077), .B(n45082), .Z(n50961) );
  NOR U58043 ( .A(n50964), .B(n50961), .Z(n47612) );
  IV U58044 ( .A(n45078), .Z(n45086) );
  IV U58045 ( .A(n45079), .Z(n45080) );
  NOR U58046 ( .A(n45086), .B(n45080), .Z(n50954) );
  IV U58047 ( .A(n45081), .Z(n45083) );
  NOR U58048 ( .A(n45083), .B(n45082), .Z(n50957) );
  NOR U58049 ( .A(n50954), .B(n50957), .Z(n47611) );
  IV U58050 ( .A(n45084), .Z(n45085) );
  NOR U58051 ( .A(n45086), .B(n45085), .Z(n50950) );
  IV U58052 ( .A(n45087), .Z(n45088) );
  NOR U58053 ( .A(n45088), .B(n45091), .Z(n50947) );
  IV U58054 ( .A(n45089), .Z(n45090) );
  NOR U58055 ( .A(n45091), .B(n45090), .Z(n50942) );
  IV U58056 ( .A(n45092), .Z(n45093) );
  NOR U58057 ( .A(n45094), .B(n45093), .Z(n48454) );
  IV U58058 ( .A(n45095), .Z(n45097) );
  NOR U58059 ( .A(n45097), .B(n45096), .Z(n48459) );
  NOR U58060 ( .A(n48454), .B(n48459), .Z(n47604) );
  IV U58061 ( .A(n45098), .Z(n45099) );
  NOR U58062 ( .A(n47595), .B(n45099), .Z(n50923) );
  IV U58063 ( .A(n45100), .Z(n45101) );
  NOR U58064 ( .A(n45101), .B(n45103), .Z(n52070) );
  IV U58065 ( .A(n45102), .Z(n45104) );
  NOR U58066 ( .A(n45104), .B(n45103), .Z(n52064) );
  NOR U58067 ( .A(n52070), .B(n52064), .Z(n50921) );
  IV U58068 ( .A(n45105), .Z(n45108) );
  IV U58069 ( .A(n45106), .Z(n45107) );
  NOR U58070 ( .A(n45108), .B(n45107), .Z(n47569) );
  IV U58071 ( .A(n47569), .Z(n47557) );
  IV U58072 ( .A(n45109), .Z(n45111) );
  IV U58073 ( .A(n45110), .Z(n47550) );
  NOR U58074 ( .A(n45111), .B(n47550), .Z(n48469) );
  IV U58075 ( .A(n45112), .Z(n45113) );
  NOR U58076 ( .A(n45114), .B(n45113), .Z(n48487) );
  IV U58077 ( .A(n45115), .Z(n45116) );
  NOR U58078 ( .A(n45117), .B(n45116), .Z(n48480) );
  NOR U58079 ( .A(n48487), .B(n48480), .Z(n47535) );
  IV U58080 ( .A(n45118), .Z(n45119) );
  NOR U58081 ( .A(n45120), .B(n45119), .Z(n48493) );
  IV U58082 ( .A(n45121), .Z(n45122) );
  NOR U58083 ( .A(n45123), .B(n45122), .Z(n48491) );
  NOR U58084 ( .A(n48493), .B(n48491), .Z(n47534) );
  IV U58085 ( .A(n45124), .Z(n45125) );
  NOR U58086 ( .A(n45126), .B(n45125), .Z(n48499) );
  IV U58087 ( .A(n45127), .Z(n45129) );
  NOR U58088 ( .A(n45129), .B(n45128), .Z(n48496) );
  NOR U58089 ( .A(n48499), .B(n48496), .Z(n47533) );
  IV U58090 ( .A(n45130), .Z(n45131) );
  NOR U58091 ( .A(n45132), .B(n45131), .Z(n50883) );
  IV U58092 ( .A(n45133), .Z(n45134) );
  NOR U58093 ( .A(n47529), .B(n45134), .Z(n50880) );
  IV U58094 ( .A(n45135), .Z(n45136) );
  NOR U58095 ( .A(n45139), .B(n45136), .Z(n48506) );
  IV U58096 ( .A(n45137), .Z(n45138) );
  NOR U58097 ( .A(n45139), .B(n45138), .Z(n50876) );
  IV U58098 ( .A(n45140), .Z(n45141) );
  NOR U58099 ( .A(n45142), .B(n45141), .Z(n48511) );
  IV U58100 ( .A(n45143), .Z(n45144) );
  NOR U58101 ( .A(n45145), .B(n45144), .Z(n48518) );
  IV U58102 ( .A(n45146), .Z(n45147) );
  NOR U58103 ( .A(n45148), .B(n45147), .Z(n48513) );
  NOR U58104 ( .A(n48518), .B(n48513), .Z(n47487) );
  IV U58105 ( .A(n45149), .Z(n45151) );
  NOR U58106 ( .A(n45151), .B(n45150), .Z(n48516) );
  IV U58107 ( .A(n45152), .Z(n45154) );
  NOR U58108 ( .A(n45154), .B(n45153), .Z(n48527) );
  NOR U58109 ( .A(n45155), .B(n47472), .Z(n47465) );
  IV U58110 ( .A(n45156), .Z(n45161) );
  IV U58111 ( .A(n45157), .Z(n45158) );
  NOR U58112 ( .A(n45161), .B(n45158), .Z(n48532) );
  IV U58113 ( .A(n45159), .Z(n45160) );
  NOR U58114 ( .A(n45161), .B(n45160), .Z(n48536) );
  IV U58115 ( .A(n45162), .Z(n45163) );
  NOR U58116 ( .A(n47460), .B(n45163), .Z(n48538) );
  NOR U58117 ( .A(n48536), .B(n48538), .Z(n47462) );
  IV U58118 ( .A(n45164), .Z(n45165) );
  NOR U58119 ( .A(n45166), .B(n45165), .Z(n54412) );
  IV U58120 ( .A(n45167), .Z(n45168) );
  NOR U58121 ( .A(n45168), .B(n47443), .Z(n52187) );
  NOR U58122 ( .A(n54412), .B(n52187), .Z(n48556) );
  IV U58123 ( .A(n45169), .Z(n45171) );
  IV U58124 ( .A(n45170), .Z(n47440) );
  NOR U58125 ( .A(n45171), .B(n47440), .Z(n48561) );
  IV U58126 ( .A(n45172), .Z(n45174) );
  NOR U58127 ( .A(n45174), .B(n45173), .Z(n47432) );
  IV U58128 ( .A(n47432), .Z(n47417) );
  IV U58129 ( .A(n45175), .Z(n45177) );
  NOR U58130 ( .A(n45177), .B(n45176), .Z(n48576) );
  IV U58131 ( .A(n45178), .Z(n47411) );
  IV U58132 ( .A(n45179), .Z(n45180) );
  NOR U58133 ( .A(n45180), .B(n47404), .Z(n47399) );
  IV U58134 ( .A(n47399), .Z(n47391) );
  IV U58135 ( .A(n45181), .Z(n48595) );
  NOR U58136 ( .A(n48595), .B(n45185), .Z(n47390) );
  IV U58137 ( .A(n45182), .Z(n45183) );
  NOR U58138 ( .A(n45183), .B(n45185), .Z(n48588) );
  NOR U58139 ( .A(n45185), .B(n45184), .Z(n45186) );
  IV U58140 ( .A(n45186), .Z(n47376) );
  IV U58141 ( .A(n45187), .Z(n45188) );
  NOR U58142 ( .A(n45188), .B(n48603), .Z(n45189) );
  IV U58143 ( .A(n45189), .Z(n48608) );
  IV U58144 ( .A(n45190), .Z(n45191) );
  NOR U58145 ( .A(n45191), .B(n45194), .Z(n50811) );
  IV U58146 ( .A(n45192), .Z(n45193) );
  NOR U58147 ( .A(n45194), .B(n45193), .Z(n50813) );
  NOR U58148 ( .A(n50811), .B(n50813), .Z(n47350) );
  NOR U58149 ( .A(n45195), .B(n48623), .Z(n47328) );
  IV U58150 ( .A(n45196), .Z(n45197) );
  NOR U58151 ( .A(n45197), .B(n45198), .Z(n48643) );
  NOR U58152 ( .A(n45199), .B(n45198), .Z(n45200) );
  IV U58153 ( .A(n45200), .Z(n47304) );
  NOR U58154 ( .A(n45201), .B(n47304), .Z(n45202) );
  IV U58155 ( .A(n45202), .Z(n45203) );
  NOR U58156 ( .A(n47303), .B(n45203), .Z(n50801) );
  NOR U58157 ( .A(n48643), .B(n50801), .Z(n47306) );
  IV U58158 ( .A(n45204), .Z(n45206) );
  IV U58159 ( .A(n45205), .Z(n47299) );
  NOR U58160 ( .A(n45206), .B(n47299), .Z(n48648) );
  IV U58161 ( .A(n45207), .Z(n45209) );
  NOR U58162 ( .A(n45209), .B(n45208), .Z(n48654) );
  NOR U58163 ( .A(n45211), .B(n45210), .Z(n48651) );
  NOR U58164 ( .A(n48654), .B(n48651), .Z(n47293) );
  NOR U58165 ( .A(n45212), .B(n48668), .Z(n45216) );
  IV U58166 ( .A(n45213), .Z(n48659) );
  NOR U58167 ( .A(n45214), .B(n48659), .Z(n45215) );
  NOR U58168 ( .A(n45216), .B(n45215), .Z(n47292) );
  IV U58169 ( .A(n45217), .Z(n48673) );
  NOR U58170 ( .A(n45218), .B(n48673), .Z(n45221) );
  IV U58171 ( .A(n45219), .Z(n45220) );
  NOR U58172 ( .A(n45220), .B(n47290), .Z(n48678) );
  NOR U58173 ( .A(n45221), .B(n48678), .Z(n47291) );
  IV U58174 ( .A(n45222), .Z(n45224) );
  NOR U58175 ( .A(n45224), .B(n45223), .Z(n47284) );
  IV U58176 ( .A(n47284), .Z(n47273) );
  NOR U58177 ( .A(n45226), .B(n45225), .Z(n45227) );
  IV U58178 ( .A(n45227), .Z(n48685) );
  IV U58179 ( .A(n45228), .Z(n45229) );
  NOR U58180 ( .A(n45230), .B(n45229), .Z(n47261) );
  IV U58181 ( .A(n45231), .Z(n45233) );
  IV U58182 ( .A(n45232), .Z(n47257) );
  NOR U58183 ( .A(n45233), .B(n47257), .Z(n48689) );
  IV U58184 ( .A(n45234), .Z(n45235) );
  NOR U58185 ( .A(n45236), .B(n45235), .Z(n50755) );
  NOR U58186 ( .A(n45237), .B(n48695), .Z(n45238) );
  NOR U58187 ( .A(n50755), .B(n45238), .Z(n47254) );
  IV U58188 ( .A(n45239), .Z(n47253) );
  IV U58189 ( .A(n45240), .Z(n45241) );
  NOR U58190 ( .A(n47253), .B(n45241), .Z(n50759) );
  IV U58191 ( .A(n45242), .Z(n45243) );
  NOR U58192 ( .A(n45244), .B(n45243), .Z(n45245) );
  IV U58193 ( .A(n45245), .Z(n50736) );
  IV U58194 ( .A(n45246), .Z(n45251) );
  IV U58195 ( .A(n45247), .Z(n45248) );
  NOR U58196 ( .A(n45251), .B(n45248), .Z(n50723) );
  IV U58197 ( .A(n45249), .Z(n45250) );
  NOR U58198 ( .A(n45251), .B(n45250), .Z(n50727) );
  IV U58199 ( .A(n45252), .Z(n45253) );
  NOR U58200 ( .A(n45253), .B(n47211), .Z(n50720) );
  NOR U58201 ( .A(n50727), .B(n50720), .Z(n47226) );
  IV U58202 ( .A(n45254), .Z(n45255) );
  NOR U58203 ( .A(n45256), .B(n45255), .Z(n50704) );
  IV U58204 ( .A(n45257), .Z(n45259) );
  NOR U58205 ( .A(n45259), .B(n45258), .Z(n50706) );
  NOR U58206 ( .A(n50704), .B(n50706), .Z(n50713) );
  IV U58207 ( .A(n50713), .Z(n45260) );
  NOR U58208 ( .A(n50712), .B(n45260), .Z(n47203) );
  IV U58209 ( .A(n45261), .Z(n45267) );
  IV U58210 ( .A(n45262), .Z(n45263) );
  NOR U58211 ( .A(n45267), .B(n45263), .Z(n45264) );
  IV U58212 ( .A(n45264), .Z(n50703) );
  IV U58213 ( .A(n45265), .Z(n45266) );
  NOR U58214 ( .A(n45267), .B(n45266), .Z(n50698) );
  IV U58215 ( .A(n45268), .Z(n45269) );
  NOR U58216 ( .A(n45271), .B(n45269), .Z(n50690) );
  IV U58217 ( .A(n45270), .Z(n45272) );
  NOR U58218 ( .A(n45272), .B(n45271), .Z(n47193) );
  IV U58219 ( .A(n47193), .Z(n47181) );
  IV U58220 ( .A(n45273), .Z(n45274) );
  NOR U58221 ( .A(n45275), .B(n45274), .Z(n47173) );
  IV U58222 ( .A(n47173), .Z(n47169) );
  IV U58223 ( .A(n45276), .Z(n45277) );
  NOR U58224 ( .A(n45282), .B(n45277), .Z(n50672) );
  IV U58225 ( .A(n45278), .Z(n45279) );
  NOR U58226 ( .A(n45280), .B(n45279), .Z(n52398) );
  IV U58227 ( .A(n45281), .Z(n45283) );
  NOR U58228 ( .A(n45283), .B(n45282), .Z(n54201) );
  NOR U58229 ( .A(n52398), .B(n54201), .Z(n48729) );
  IV U58230 ( .A(n45284), .Z(n45285) );
  NOR U58231 ( .A(n45286), .B(n45285), .Z(n47140) );
  IV U58232 ( .A(n47140), .Z(n47135) );
  IV U58233 ( .A(n45287), .Z(n45288) );
  NOR U58234 ( .A(n45288), .B(n45296), .Z(n48741) );
  IV U58235 ( .A(n45289), .Z(n45291) );
  NOR U58236 ( .A(n45291), .B(n45290), .Z(n50667) );
  NOR U58237 ( .A(n48741), .B(n50667), .Z(n47134) );
  IV U58238 ( .A(n45292), .Z(n45293) );
  NOR U58239 ( .A(n45294), .B(n45293), .Z(n50650) );
  IV U58240 ( .A(n45295), .Z(n45297) );
  NOR U58241 ( .A(n45297), .B(n45296), .Z(n50659) );
  NOR U58242 ( .A(n50650), .B(n50659), .Z(n47133) );
  IV U58243 ( .A(n45298), .Z(n45299) );
  NOR U58244 ( .A(n45299), .B(n45307), .Z(n50639) );
  IV U58245 ( .A(n45300), .Z(n45302) );
  NOR U58246 ( .A(n45302), .B(n45301), .Z(n48744) );
  NOR U58247 ( .A(n50639), .B(n48744), .Z(n47132) );
  IV U58248 ( .A(n45303), .Z(n45305) );
  NOR U58249 ( .A(n45305), .B(n45304), .Z(n50630) );
  IV U58250 ( .A(n45306), .Z(n45308) );
  NOR U58251 ( .A(n45308), .B(n45307), .Z(n50633) );
  NOR U58252 ( .A(n50630), .B(n50633), .Z(n47131) );
  IV U58253 ( .A(n45309), .Z(n45310) );
  NOR U58254 ( .A(n45311), .B(n45310), .Z(n45312) );
  IV U58255 ( .A(n45312), .Z(n47122) );
  IV U58256 ( .A(n45313), .Z(n45315) );
  NOR U58257 ( .A(n45315), .B(n45314), .Z(n48750) );
  IV U58258 ( .A(n45316), .Z(n45317) );
  NOR U58259 ( .A(n45317), .B(n47113), .Z(n50598) );
  IV U58260 ( .A(n45318), .Z(n45322) );
  IV U58261 ( .A(n45319), .Z(n47102) );
  NOR U58262 ( .A(n45320), .B(n47102), .Z(n45321) );
  IV U58263 ( .A(n45321), .Z(n47105) );
  NOR U58264 ( .A(n45322), .B(n47105), .Z(n48760) );
  IV U58265 ( .A(n45323), .Z(n45326) );
  NOR U58266 ( .A(n45324), .B(n45331), .Z(n45325) );
  IV U58267 ( .A(n45325), .Z(n45328) );
  NOR U58268 ( .A(n45326), .B(n45328), .Z(n48762) );
  NOR U58269 ( .A(n48760), .B(n48762), .Z(n47099) );
  IV U58270 ( .A(n45327), .Z(n45329) );
  NOR U58271 ( .A(n45329), .B(n45328), .Z(n48766) );
  IV U58272 ( .A(n45330), .Z(n45332) );
  NOR U58273 ( .A(n45332), .B(n45331), .Z(n48768) );
  NOR U58274 ( .A(n48766), .B(n48768), .Z(n47098) );
  IV U58275 ( .A(n45333), .Z(n45335) );
  NOR U58276 ( .A(n45335), .B(n45334), .Z(n50590) );
  IV U58277 ( .A(n45336), .Z(n45337) );
  NOR U58278 ( .A(n45338), .B(n45337), .Z(n50593) );
  NOR U58279 ( .A(n50590), .B(n50593), .Z(n47097) );
  IV U58280 ( .A(n45339), .Z(n45340) );
  NOR U58281 ( .A(n45341), .B(n45340), .Z(n50578) );
  IV U58282 ( .A(n45342), .Z(n45343) );
  NOR U58283 ( .A(n47088), .B(n45343), .Z(n50573) );
  NOR U58284 ( .A(n50578), .B(n50573), .Z(n47089) );
  IV U58285 ( .A(n45344), .Z(n45346) );
  NOR U58286 ( .A(n45346), .B(n45345), .Z(n50558) );
  IV U58287 ( .A(n45347), .Z(n45348) );
  NOR U58288 ( .A(n45348), .B(n45353), .Z(n48780) );
  NOR U58289 ( .A(n50558), .B(n48780), .Z(n47078) );
  IV U58290 ( .A(n45349), .Z(n45350) );
  NOR U58291 ( .A(n45350), .B(n45358), .Z(n48783) );
  IV U58292 ( .A(n45351), .Z(n45352) );
  NOR U58293 ( .A(n45353), .B(n45352), .Z(n50550) );
  NOR U58294 ( .A(n48783), .B(n50550), .Z(n47077) );
  IV U58295 ( .A(n45354), .Z(n45356) );
  NOR U58296 ( .A(n45356), .B(n45355), .Z(n50535) );
  IV U58297 ( .A(n45357), .Z(n45359) );
  NOR U58298 ( .A(n45359), .B(n45358), .Z(n50546) );
  NOR U58299 ( .A(n50535), .B(n50546), .Z(n47076) );
  IV U58300 ( .A(n45360), .Z(n45361) );
  NOR U58301 ( .A(n45362), .B(n45361), .Z(n50541) );
  IV U58302 ( .A(n45363), .Z(n45364) );
  NOR U58303 ( .A(n45364), .B(n47072), .Z(n50538) );
  IV U58304 ( .A(n45365), .Z(n45366) );
  NOR U58305 ( .A(n45366), .B(n45368), .Z(n52472) );
  NOR U58306 ( .A(n45368), .B(n45367), .Z(n52479) );
  NOR U58307 ( .A(n52472), .B(n52479), .Z(n45369) );
  IV U58308 ( .A(n45369), .Z(n50511) );
  NOR U58309 ( .A(n50511), .B(n50519), .Z(n47066) );
  NOR U58310 ( .A(n45370), .B(n52483), .Z(n50514) );
  IV U58311 ( .A(n45371), .Z(n45372) );
  NOR U58312 ( .A(n45373), .B(n45372), .Z(n52495) );
  IV U58313 ( .A(n45374), .Z(n45375) );
  NOR U58314 ( .A(n45376), .B(n45375), .Z(n52489) );
  NOR U58315 ( .A(n52495), .B(n52489), .Z(n50510) );
  IV U58316 ( .A(n50510), .Z(n50509) );
  IV U58317 ( .A(n45377), .Z(n45379) );
  NOR U58318 ( .A(n45379), .B(n45378), .Z(n50490) );
  IV U58319 ( .A(n45380), .Z(n45382) );
  NOR U58320 ( .A(n45382), .B(n45381), .Z(n48790) );
  NOR U58321 ( .A(n50490), .B(n48790), .Z(n47065) );
  IV U58322 ( .A(n45383), .Z(n45385) );
  XOR U58323 ( .A(n45386), .B(n45387), .Z(n45390) );
  XOR U58324 ( .A(n45389), .B(n45390), .Z(n45384) );
  NOR U58325 ( .A(n45385), .B(n45384), .Z(n48793) );
  IV U58326 ( .A(n45386), .Z(n45388) );
  NOR U58327 ( .A(n45388), .B(n45387), .Z(n48800) );
  IV U58328 ( .A(n45389), .Z(n45391) );
  NOR U58329 ( .A(n45391), .B(n45390), .Z(n48797) );
  NOR U58330 ( .A(n48800), .B(n48797), .Z(n47058) );
  IV U58331 ( .A(n45392), .Z(n45393) );
  NOR U58332 ( .A(n45393), .B(n47049), .Z(n48805) );
  IV U58333 ( .A(n45394), .Z(n47047) );
  IV U58334 ( .A(n45395), .Z(n45396) );
  NOR U58335 ( .A(n47047), .B(n45396), .Z(n54091) );
  IV U58336 ( .A(n45397), .Z(n45399) );
  NOR U58337 ( .A(n45399), .B(n45398), .Z(n54077) );
  NOR U58338 ( .A(n54091), .B(n54077), .Z(n48820) );
  IV U58339 ( .A(n45400), .Z(n45401) );
  NOR U58340 ( .A(n45401), .B(n45407), .Z(n48826) );
  IV U58341 ( .A(n45402), .Z(n45403) );
  NOR U58342 ( .A(n45404), .B(n45403), .Z(n48834) );
  IV U58343 ( .A(n45405), .Z(n45406) );
  NOR U58344 ( .A(n45407), .B(n45406), .Z(n50474) );
  NOR U58345 ( .A(n48834), .B(n50474), .Z(n47035) );
  IV U58346 ( .A(n45408), .Z(n45409) );
  NOR U58347 ( .A(n45409), .B(n47033), .Z(n50463) );
  IV U58348 ( .A(n45410), .Z(n45411) );
  NOR U58349 ( .A(n45412), .B(n45411), .Z(n48839) );
  IV U58350 ( .A(n45413), .Z(n45414) );
  NOR U58351 ( .A(n45414), .B(n45416), .Z(n48847) );
  NOR U58352 ( .A(n48839), .B(n48847), .Z(n47026) );
  IV U58353 ( .A(n45415), .Z(n45419) );
  NOR U58354 ( .A(n45417), .B(n45416), .Z(n45418) );
  IV U58355 ( .A(n45418), .Z(n45421) );
  NOR U58356 ( .A(n45419), .B(n45421), .Z(n48844) );
  IV U58357 ( .A(n45420), .Z(n45422) );
  NOR U58358 ( .A(n45422), .B(n45421), .Z(n48841) );
  IV U58359 ( .A(n45423), .Z(n45424) );
  NOR U58360 ( .A(n46991), .B(n45424), .Z(n50442) );
  NOR U58361 ( .A(n45426), .B(n45425), .Z(n45427) );
  IV U58362 ( .A(n45427), .Z(n48863) );
  IV U58363 ( .A(n45428), .Z(n45430) );
  NOR U58364 ( .A(n45430), .B(n45429), .Z(n46981) );
  IV U58365 ( .A(n46981), .Z(n46972) );
  IV U58366 ( .A(n45431), .Z(n45433) );
  NOR U58367 ( .A(n45433), .B(n45432), .Z(n45434) );
  IV U58368 ( .A(n45434), .Z(n48866) );
  IV U58369 ( .A(n45435), .Z(n45436) );
  NOR U58370 ( .A(n45436), .B(n46955), .Z(n52590) );
  IV U58371 ( .A(n45437), .Z(n45439) );
  NOR U58372 ( .A(n45439), .B(n45438), .Z(n52582) );
  NOR U58373 ( .A(n52590), .B(n52582), .Z(n50388) );
  NOR U58374 ( .A(n45441), .B(n45440), .Z(n50385) );
  IV U58375 ( .A(n45442), .Z(n45443) );
  NOR U58376 ( .A(n45444), .B(n45443), .Z(n45445) );
  IV U58377 ( .A(n45445), .Z(n46924) );
  IV U58378 ( .A(n45446), .Z(n45447) );
  NOR U58379 ( .A(n45448), .B(n45447), .Z(n53998) );
  IV U58380 ( .A(n45449), .Z(n45450) );
  NOR U58381 ( .A(n46922), .B(n45450), .Z(n52608) );
  NOR U58382 ( .A(n53998), .B(n52608), .Z(n50354) );
  IV U58383 ( .A(n45451), .Z(n45452) );
  NOR U58384 ( .A(n45452), .B(n45456), .Z(n46918) );
  IV U58385 ( .A(n45453), .Z(n50342) );
  NOR U58386 ( .A(n45454), .B(n50342), .Z(n45458) );
  IV U58387 ( .A(n45455), .Z(n45457) );
  NOR U58388 ( .A(n45457), .B(n45456), .Z(n50346) );
  NOR U58389 ( .A(n45458), .B(n50346), .Z(n46916) );
  IV U58390 ( .A(n45459), .Z(n45460) );
  NOR U58391 ( .A(n45460), .B(n46909), .Z(n45461) );
  IV U58392 ( .A(n45461), .Z(n50339) );
  IV U58393 ( .A(n45462), .Z(n45463) );
  NOR U58394 ( .A(n45464), .B(n45463), .Z(n45465) );
  IV U58395 ( .A(n45465), .Z(n46911) );
  IV U58396 ( .A(n48907), .Z(n48908) );
  IV U58397 ( .A(n45466), .Z(n45476) );
  IV U58398 ( .A(n45467), .Z(n45468) );
  NOR U58399 ( .A(n45476), .B(n45468), .Z(n50334) );
  IV U58400 ( .A(n45469), .Z(n45473) );
  NOR U58401 ( .A(n45471), .B(n45470), .Z(n45472) );
  IV U58402 ( .A(n45472), .Z(n46901) );
  NOR U58403 ( .A(n45473), .B(n46901), .Z(n48914) );
  NOR U58404 ( .A(n50334), .B(n48914), .Z(n46905) );
  IV U58405 ( .A(n45474), .Z(n45475) );
  NOR U58406 ( .A(n45476), .B(n45475), .Z(n48916) );
  IV U58407 ( .A(n45477), .Z(n45479) );
  NOR U58408 ( .A(n45479), .B(n45478), .Z(n50329) );
  NOR U58409 ( .A(n48916), .B(n50329), .Z(n46898) );
  IV U58410 ( .A(n45480), .Z(n45482) );
  IV U58411 ( .A(n45481), .Z(n45485) );
  NOR U58412 ( .A(n45482), .B(n45485), .Z(n50321) );
  NOR U58413 ( .A(n45483), .B(n50315), .Z(n45486) );
  NOR U58414 ( .A(n45485), .B(n45484), .Z(n50324) );
  NOR U58415 ( .A(n45486), .B(n50324), .Z(n46897) );
  IV U58416 ( .A(n45487), .Z(n45488) );
  NOR U58417 ( .A(n45489), .B(n45488), .Z(n53957) );
  IV U58418 ( .A(n45490), .Z(n45491) );
  NOR U58419 ( .A(n45492), .B(n45491), .Z(n53962) );
  NOR U58420 ( .A(n53957), .B(n53962), .Z(n50294) );
  IV U58421 ( .A(n45493), .Z(n45495) );
  NOR U58422 ( .A(n45495), .B(n45494), .Z(n50283) );
  IV U58423 ( .A(n45496), .Z(n45497) );
  NOR U58424 ( .A(n45498), .B(n45497), .Z(n50287) );
  NOR U58425 ( .A(n50283), .B(n50287), .Z(n48924) );
  IV U58426 ( .A(n45499), .Z(n45500) );
  NOR U58427 ( .A(n45501), .B(n45500), .Z(n48925) );
  IV U58428 ( .A(n45502), .Z(n45504) );
  NOR U58429 ( .A(n45504), .B(n45503), .Z(n50278) );
  NOR U58430 ( .A(n48925), .B(n50278), .Z(n46883) );
  IV U58431 ( .A(n45505), .Z(n45506) );
  NOR U58432 ( .A(n45506), .B(n46870), .Z(n50269) );
  IV U58433 ( .A(n45507), .Z(n45509) );
  NOR U58434 ( .A(n45509), .B(n45508), .Z(n45510) );
  IV U58435 ( .A(n45510), .Z(n46876) );
  IV U58436 ( .A(n45511), .Z(n46865) );
  IV U58437 ( .A(n45512), .Z(n45513) );
  NOR U58438 ( .A(n46865), .B(n45513), .Z(n48930) );
  IV U58439 ( .A(n45514), .Z(n45516) );
  NOR U58440 ( .A(n45516), .B(n45515), .Z(n45517) );
  IV U58441 ( .A(n45517), .Z(n46858) );
  IV U58442 ( .A(n45518), .Z(n45520) );
  NOR U58443 ( .A(n45520), .B(n45519), .Z(n52679) );
  IV U58444 ( .A(n45521), .Z(n45522) );
  NOR U58445 ( .A(n45522), .B(n48948), .Z(n52675) );
  NOR U58446 ( .A(n52679), .B(n52675), .Z(n48945) );
  IV U58447 ( .A(n45523), .Z(n45524) );
  NOR U58448 ( .A(n45524), .B(n45526), .Z(n48953) );
  IV U58449 ( .A(n45525), .Z(n45527) );
  NOR U58450 ( .A(n45527), .B(n45526), .Z(n48956) );
  NOR U58451 ( .A(n48953), .B(n48956), .Z(n45528) );
  IV U58452 ( .A(n45528), .Z(n45534) );
  NOR U58453 ( .A(n45530), .B(n45529), .Z(n45531) );
  IV U58454 ( .A(n45531), .Z(n48963) );
  NOR U58455 ( .A(n45532), .B(n48963), .Z(n45533) );
  NOR U58456 ( .A(n45534), .B(n45533), .Z(n46852) );
  IV U58457 ( .A(n45535), .Z(n45541) );
  NOR U58458 ( .A(n45536), .B(n46812), .Z(n45537) );
  IV U58459 ( .A(n45537), .Z(n45538) );
  NOR U58460 ( .A(n45539), .B(n45538), .Z(n45540) );
  IV U58461 ( .A(n45540), .Z(n46815) );
  NOR U58462 ( .A(n45541), .B(n46815), .Z(n50245) );
  IV U58463 ( .A(n45542), .Z(n46811) );
  IV U58464 ( .A(n45543), .Z(n45545) );
  NOR U58465 ( .A(n45545), .B(n45544), .Z(n45546) );
  IV U58466 ( .A(n45546), .Z(n46798) );
  IV U58467 ( .A(n45547), .Z(n45548) );
  NOR U58468 ( .A(n45549), .B(n45548), .Z(n50204) );
  IV U58469 ( .A(n45550), .Z(n45551) );
  NOR U58470 ( .A(n45552), .B(n45551), .Z(n50192) );
  NOR U58471 ( .A(n50204), .B(n50192), .Z(n46778) );
  IV U58472 ( .A(n45553), .Z(n45554) );
  NOR U58473 ( .A(n45555), .B(n45554), .Z(n45556) );
  IV U58474 ( .A(n45556), .Z(n50212) );
  IV U58475 ( .A(n45557), .Z(n45559) );
  NOR U58476 ( .A(n45559), .B(n45558), .Z(n50189) );
  IV U58477 ( .A(n45560), .Z(n45561) );
  NOR U58478 ( .A(n45562), .B(n45561), .Z(n50196) );
  NOR U58479 ( .A(n50189), .B(n50196), .Z(n46775) );
  IV U58480 ( .A(n45563), .Z(n46770) );
  IV U58481 ( .A(n45564), .Z(n45565) );
  NOR U58482 ( .A(n46770), .B(n45565), .Z(n50186) );
  IV U58483 ( .A(n45566), .Z(n45567) );
  NOR U58484 ( .A(n45567), .B(n46772), .Z(n46766) );
  IV U58485 ( .A(n46766), .Z(n46761) );
  IV U58486 ( .A(n45568), .Z(n45572) );
  NOR U58487 ( .A(n45570), .B(n45569), .Z(n45571) );
  IV U58488 ( .A(n45571), .Z(n46749) );
  NOR U58489 ( .A(n45572), .B(n46749), .Z(n50155) );
  IV U58490 ( .A(n45573), .Z(n45574) );
  NOR U58491 ( .A(n46746), .B(n45574), .Z(n48987) );
  NOR U58492 ( .A(n50155), .B(n48987), .Z(n46747) );
  IV U58493 ( .A(n45575), .Z(n45576) );
  NOR U58494 ( .A(n45576), .B(n45582), .Z(n50148) );
  IV U58495 ( .A(n45577), .Z(n45578) );
  NOR U58496 ( .A(n45579), .B(n45578), .Z(n48991) );
  IV U58497 ( .A(n45580), .Z(n45581) );
  NOR U58498 ( .A(n45582), .B(n45581), .Z(n48989) );
  NOR U58499 ( .A(n48991), .B(n48989), .Z(n46739) );
  IV U58500 ( .A(n45583), .Z(n45584) );
  NOR U58501 ( .A(n45585), .B(n45584), .Z(n49007) );
  NOR U58502 ( .A(n50141), .B(n49007), .Z(n46706) );
  IV U58503 ( .A(n45586), .Z(n45587) );
  NOR U58504 ( .A(n45587), .B(n45592), .Z(n50135) );
  NOR U58505 ( .A(n45589), .B(n45588), .Z(n50132) );
  IV U58506 ( .A(n45590), .Z(n45591) );
  NOR U58507 ( .A(n45592), .B(n45591), .Z(n50137) );
  NOR U58508 ( .A(n50132), .B(n50137), .Z(n46704) );
  IV U58509 ( .A(n45593), .Z(n45596) );
  NOR U58510 ( .A(n45594), .B(n46697), .Z(n45595) );
  IV U58511 ( .A(n45595), .Z(n46702) );
  NOR U58512 ( .A(n45596), .B(n46702), .Z(n50117) );
  IV U58513 ( .A(n45597), .Z(n45598) );
  NOR U58514 ( .A(n45598), .B(n45603), .Z(n49013) );
  IV U58515 ( .A(n45599), .Z(n45600) );
  NOR U58516 ( .A(n45601), .B(n45600), .Z(n49020) );
  IV U58517 ( .A(n45602), .Z(n45604) );
  NOR U58518 ( .A(n45604), .B(n45603), .Z(n49018) );
  NOR U58519 ( .A(n49020), .B(n49018), .Z(n46691) );
  IV U58520 ( .A(n45605), .Z(n50091) );
  XOR U58521 ( .A(n50091), .B(n45606), .Z(n45607) );
  NOR U58522 ( .A(n45607), .B(n50100), .Z(n46690) );
  IV U58523 ( .A(n45608), .Z(n45610) );
  IV U58524 ( .A(n45609), .Z(n46688) );
  NOR U58525 ( .A(n45610), .B(n46688), .Z(n49029) );
  IV U58526 ( .A(n45611), .Z(n45612) );
  NOR U58527 ( .A(n45612), .B(n46688), .Z(n49033) );
  NOR U58528 ( .A(n49036), .B(n49033), .Z(n46682) );
  NOR U58529 ( .A(n45614), .B(n45613), .Z(n46680) );
  IV U58530 ( .A(n46680), .Z(n46678) );
  NOR U58531 ( .A(n49049), .B(n49052), .Z(n45615) );
  IV U58532 ( .A(n45615), .Z(n45616) );
  NOR U58533 ( .A(n49043), .B(n45616), .Z(n46676) );
  NOR U58534 ( .A(n45617), .B(n49046), .Z(n46675) );
  IV U58535 ( .A(n45618), .Z(n45620) );
  NOR U58536 ( .A(n45620), .B(n45619), .Z(n50076) );
  NOR U58537 ( .A(n45621), .B(n49060), .Z(n45622) );
  NOR U58538 ( .A(n50076), .B(n45622), .Z(n46673) );
  IV U58539 ( .A(n45623), .Z(n45624) );
  NOR U58540 ( .A(n45625), .B(n45624), .Z(n50061) );
  IV U58541 ( .A(n45626), .Z(n45627) );
  NOR U58542 ( .A(n45627), .B(n46670), .Z(n50057) );
  IV U58543 ( .A(n45628), .Z(n45630) );
  NOR U58544 ( .A(n45630), .B(n45629), .Z(n45631) );
  IV U58545 ( .A(n45631), .Z(n50044) );
  IV U58546 ( .A(n45632), .Z(n45634) );
  NOR U58547 ( .A(n45634), .B(n45633), .Z(n50032) );
  IV U58548 ( .A(n45635), .Z(n45636) );
  NOR U58549 ( .A(n46638), .B(n45636), .Z(n49075) );
  NOR U58550 ( .A(n50032), .B(n49075), .Z(n46634) );
  IV U58551 ( .A(n45637), .Z(n45639) );
  NOR U58552 ( .A(n45639), .B(n45638), .Z(n52844) );
  IV U58553 ( .A(n45640), .Z(n45644) );
  NOR U58554 ( .A(n45642), .B(n45641), .Z(n45643) );
  IV U58555 ( .A(n45643), .Z(n45646) );
  NOR U58556 ( .A(n45644), .B(n45646), .Z(n52848) );
  NOR U58557 ( .A(n52844), .B(n52848), .Z(n50031) );
  IV U58558 ( .A(n45645), .Z(n45647) );
  NOR U58559 ( .A(n45647), .B(n45646), .Z(n49078) );
  NOR U58560 ( .A(n50023), .B(n49078), .Z(n46633) );
  IV U58561 ( .A(n45648), .Z(n45650) );
  NOR U58562 ( .A(n45650), .B(n45649), .Z(n50025) );
  IV U58563 ( .A(n50025), .Z(n50022) );
  IV U58564 ( .A(n45651), .Z(n49080) );
  IV U58565 ( .A(n45652), .Z(n45654) );
  NOR U58566 ( .A(n45654), .B(n45653), .Z(n46628) );
  IV U58567 ( .A(n46628), .Z(n46619) );
  IV U58568 ( .A(n45655), .Z(n45656) );
  NOR U58569 ( .A(n45657), .B(n45656), .Z(n45658) );
  IV U58570 ( .A(n45658), .Z(n49085) );
  NOR U58571 ( .A(n45660), .B(n45659), .Z(n49999) );
  IV U58572 ( .A(n45661), .Z(n45662) );
  NOR U58573 ( .A(n45663), .B(n45662), .Z(n49988) );
  NOR U58574 ( .A(n49988), .B(n49090), .Z(n46607) );
  IV U58575 ( .A(n45664), .Z(n45666) );
  NOR U58576 ( .A(n45666), .B(n45665), .Z(n45667) );
  IV U58577 ( .A(n45667), .Z(n46602) );
  IV U58578 ( .A(n45668), .Z(n45669) );
  NOR U58579 ( .A(n45670), .B(n45669), .Z(n49977) );
  IV U58580 ( .A(n45671), .Z(n45672) );
  NOR U58581 ( .A(n45673), .B(n45672), .Z(n49969) );
  IV U58582 ( .A(n45674), .Z(n45676) );
  NOR U58583 ( .A(n45676), .B(n45675), .Z(n49098) );
  NOR U58584 ( .A(n49098), .B(n49096), .Z(n46584) );
  IV U58585 ( .A(n45677), .Z(n45679) );
  IV U58586 ( .A(n45678), .Z(n45681) );
  NOR U58587 ( .A(n45679), .B(n45681), .Z(n49959) );
  IV U58588 ( .A(n45680), .Z(n45682) );
  NOR U58589 ( .A(n45682), .B(n45681), .Z(n49956) );
  IV U58590 ( .A(n45683), .Z(n49934) );
  IV U58591 ( .A(n45684), .Z(n45685) );
  NOR U58592 ( .A(n49934), .B(n45685), .Z(n49116) );
  IV U58593 ( .A(n45686), .Z(n45687) );
  NOR U58594 ( .A(n45687), .B(n45689), .Z(n49135) );
  IV U58595 ( .A(n45688), .Z(n45690) );
  NOR U58596 ( .A(n45690), .B(n45689), .Z(n46556) );
  IV U58597 ( .A(n46556), .Z(n46547) );
  IV U58598 ( .A(n45691), .Z(n45693) );
  NOR U58599 ( .A(n45693), .B(n45692), .Z(n45694) );
  IV U58600 ( .A(n45694), .Z(n49919) );
  IV U58601 ( .A(n45695), .Z(n45700) );
  IV U58602 ( .A(n45696), .Z(n45697) );
  NOR U58603 ( .A(n45697), .B(n46540), .Z(n45698) );
  IV U58604 ( .A(n45698), .Z(n45699) );
  NOR U58605 ( .A(n45700), .B(n45699), .Z(n49138) );
  IV U58606 ( .A(n45701), .Z(n45702) );
  NOR U58607 ( .A(n46535), .B(n45702), .Z(n49142) );
  IV U58608 ( .A(n45703), .Z(n45705) );
  NOR U58609 ( .A(n45705), .B(n45704), .Z(n45706) );
  IV U58610 ( .A(n45706), .Z(n46527) );
  IV U58611 ( .A(n45707), .Z(n46525) );
  IV U58612 ( .A(n45708), .Z(n45709) );
  NOR U58613 ( .A(n46525), .B(n45709), .Z(n49153) );
  NOR U58614 ( .A(n49155), .B(n49153), .Z(n46519) );
  NOR U58615 ( .A(n49167), .B(n49165), .Z(n46518) );
  IV U58616 ( .A(n45710), .Z(n45713) );
  NOR U58617 ( .A(n46510), .B(n45711), .Z(n45712) );
  IV U58618 ( .A(n45712), .Z(n46516) );
  NOR U58619 ( .A(n45713), .B(n46516), .Z(n49173) );
  NOR U58620 ( .A(n45715), .B(n45714), .Z(n52976) );
  IV U58621 ( .A(n45716), .Z(n46512) );
  IV U58622 ( .A(n45717), .Z(n45718) );
  NOR U58623 ( .A(n46512), .B(n45718), .Z(n52972) );
  NOR U58624 ( .A(n52976), .B(n52972), .Z(n49907) );
  IV U58625 ( .A(n45719), .Z(n45720) );
  NOR U58626 ( .A(n45722), .B(n45720), .Z(n49203) );
  NOR U58627 ( .A(n45722), .B(n45721), .Z(n49206) );
  IV U58628 ( .A(n45723), .Z(n45725) );
  NOR U58629 ( .A(n45725), .B(n45724), .Z(n49886) );
  IV U58630 ( .A(n45726), .Z(n45728) );
  NOR U58631 ( .A(n45728), .B(n45727), .Z(n49209) );
  NOR U58632 ( .A(n49886), .B(n49209), .Z(n46475) );
  IV U58633 ( .A(n45729), .Z(n45730) );
  NOR U58634 ( .A(n45730), .B(n46472), .Z(n49883) );
  IV U58635 ( .A(n45731), .Z(n45732) );
  NOR U58636 ( .A(n45733), .B(n45732), .Z(n53011) );
  IV U58637 ( .A(n45734), .Z(n45735) );
  NOR U58638 ( .A(n45736), .B(n45735), .Z(n53659) );
  NOR U58639 ( .A(n53011), .B(n53659), .Z(n49217) );
  IV U58640 ( .A(n45737), .Z(n45738) );
  NOR U58641 ( .A(n46466), .B(n45738), .Z(n49225) );
  IV U58642 ( .A(n45739), .Z(n45741) );
  NOR U58643 ( .A(n45741), .B(n45740), .Z(n45742) );
  IV U58644 ( .A(n45742), .Z(n46459) );
  IV U58645 ( .A(n45743), .Z(n45745) );
  NOR U58646 ( .A(n45745), .B(n45744), .Z(n49238) );
  IV U58647 ( .A(n45746), .Z(n45747) );
  NOR U58648 ( .A(n45747), .B(n46443), .Z(n49858) );
  NOR U58649 ( .A(n49238), .B(n49858), .Z(n49853) );
  IV U58650 ( .A(n45748), .Z(n45749) );
  NOR U58651 ( .A(n45750), .B(n45749), .Z(n53643) );
  IV U58652 ( .A(n45751), .Z(n45754) );
  IV U58653 ( .A(n45752), .Z(n45753) );
  NOR U58654 ( .A(n45754), .B(n45753), .Z(n53022) );
  NOR U58655 ( .A(n53643), .B(n53022), .Z(n49854) );
  IV U58656 ( .A(n45755), .Z(n45759) );
  NOR U58657 ( .A(n45757), .B(n45756), .Z(n45758) );
  IV U58658 ( .A(n45758), .Z(n46440) );
  NOR U58659 ( .A(n45759), .B(n46440), .Z(n49239) );
  IV U58660 ( .A(n45760), .Z(n45761) );
  NOR U58661 ( .A(n49247), .B(n45761), .Z(n49245) );
  NOR U58662 ( .A(n45762), .B(n49245), .Z(n46438) );
  NOR U58663 ( .A(n45763), .B(n49257), .Z(n46420) );
  IV U58664 ( .A(n45764), .Z(n45765) );
  NOR U58665 ( .A(n46410), .B(n45765), .Z(n49837) );
  IV U58666 ( .A(n45766), .Z(n45768) );
  NOR U58667 ( .A(n45768), .B(n45767), .Z(n49276) );
  IV U58668 ( .A(n45769), .Z(n45771) );
  NOR U58669 ( .A(n45771), .B(n45770), .Z(n49840) );
  NOR U58670 ( .A(n49276), .B(n49840), .Z(n46407) );
  IV U58671 ( .A(n45772), .Z(n46401) );
  IV U58672 ( .A(n45773), .Z(n45774) );
  NOR U58673 ( .A(n46401), .B(n45774), .Z(n49273) );
  IV U58674 ( .A(n45775), .Z(n45778) );
  NOR U58675 ( .A(n45776), .B(n46403), .Z(n45777) );
  IV U58676 ( .A(n45777), .Z(n45783) );
  NOR U58677 ( .A(n45778), .B(n45783), .Z(n49830) );
  IV U58678 ( .A(n45779), .Z(n45781) );
  IV U58679 ( .A(n45780), .Z(n49282) );
  NOR U58680 ( .A(n45781), .B(n49282), .Z(n53061) );
  IV U58681 ( .A(n45782), .Z(n45784) );
  NOR U58682 ( .A(n45784), .B(n45783), .Z(n49825) );
  NOR U58683 ( .A(n53061), .B(n49825), .Z(n46398) );
  IV U58684 ( .A(n45785), .Z(n45787) );
  NOR U58685 ( .A(n45787), .B(n45786), .Z(n49286) );
  IV U58686 ( .A(n45788), .Z(n45789) );
  NOR U58687 ( .A(n45790), .B(n45789), .Z(n49311) );
  IV U58688 ( .A(n45791), .Z(n45793) );
  NOR U58689 ( .A(n45793), .B(n45792), .Z(n45797) );
  IV U58690 ( .A(n45794), .Z(n45795) );
  NOR U58691 ( .A(n45795), .B(n45799), .Z(n45796) );
  NOR U58692 ( .A(n45797), .B(n45796), .Z(n49316) );
  IV U58693 ( .A(n45798), .Z(n45800) );
  NOR U58694 ( .A(n45800), .B(n45799), .Z(n49320) );
  IV U58695 ( .A(n45801), .Z(n45802) );
  NOR U58696 ( .A(n45803), .B(n45802), .Z(n46321) );
  IV U58697 ( .A(n46321), .Z(n46307) );
  IV U58698 ( .A(n45804), .Z(n49344) );
  NOR U58699 ( .A(n45806), .B(n45805), .Z(n49345) );
  IV U58700 ( .A(n45807), .Z(n45809) );
  NOR U58701 ( .A(n45809), .B(n45808), .Z(n46301) );
  IV U58702 ( .A(n46301), .Z(n46291) );
  IV U58703 ( .A(n45810), .Z(n45812) );
  NOR U58704 ( .A(n45812), .B(n45811), .Z(n56607) );
  IV U58705 ( .A(n45813), .Z(n45814) );
  NOR U58706 ( .A(n45814), .B(n45820), .Z(n49361) );
  IV U58707 ( .A(n45815), .Z(n45816) );
  NOR U58708 ( .A(n45817), .B(n45816), .Z(n49367) );
  IV U58709 ( .A(n45818), .Z(n45819) );
  NOR U58710 ( .A(n45820), .B(n45819), .Z(n49359) );
  NOR U58711 ( .A(n49367), .B(n49359), .Z(n46282) );
  IV U58712 ( .A(n45821), .Z(n45822) );
  NOR U58713 ( .A(n45822), .B(n46277), .Z(n49364) );
  IV U58714 ( .A(n45823), .Z(n45824) );
  NOR U58715 ( .A(n45824), .B(n45826), .Z(n49775) );
  IV U58716 ( .A(n45825), .Z(n45827) );
  NOR U58717 ( .A(n45827), .B(n45826), .Z(n46271) );
  IV U58718 ( .A(n46271), .Z(n46265) );
  IV U58719 ( .A(n45828), .Z(n45829) );
  NOR U58720 ( .A(n46261), .B(n45829), .Z(n49768) );
  IV U58721 ( .A(n45830), .Z(n45831) );
  NOR U58722 ( .A(n45832), .B(n45831), .Z(n49380) );
  IV U58723 ( .A(n45833), .Z(n45834) );
  NOR U58724 ( .A(n45836), .B(n45834), .Z(n49389) );
  IV U58725 ( .A(n45835), .Z(n45837) );
  NOR U58726 ( .A(n45837), .B(n45836), .Z(n49386) );
  NOR U58727 ( .A(n49389), .B(n49386), .Z(n46256) );
  IV U58728 ( .A(n45838), .Z(n45839) );
  NOR U58729 ( .A(n45840), .B(n45839), .Z(n46231) );
  IV U58730 ( .A(n46231), .Z(n46221) );
  IV U58731 ( .A(n45841), .Z(n45843) );
  NOR U58732 ( .A(n45843), .B(n45842), .Z(n46218) );
  IV U58733 ( .A(n46218), .Z(n46213) );
  IV U58734 ( .A(n45844), .Z(n45845) );
  NOR U58735 ( .A(n46211), .B(n45845), .Z(n46205) );
  IV U58736 ( .A(n45846), .Z(n45848) );
  NOR U58737 ( .A(n45848), .B(n45847), .Z(n49411) );
  IV U58738 ( .A(n45849), .Z(n45850) );
  NOR U58739 ( .A(n45853), .B(n45850), .Z(n49756) );
  NOR U58740 ( .A(n49411), .B(n49756), .Z(n46192) );
  IV U58741 ( .A(n45851), .Z(n45852) );
  NOR U58742 ( .A(n45853), .B(n45852), .Z(n49409) );
  IV U58743 ( .A(n45854), .Z(n45855) );
  NOR U58744 ( .A(n45856), .B(n45855), .Z(n49417) );
  IV U58745 ( .A(n45857), .Z(n45858) );
  NOR U58746 ( .A(n45859), .B(n45858), .Z(n49414) );
  NOR U58747 ( .A(n49417), .B(n49414), .Z(n46190) );
  IV U58748 ( .A(n45860), .Z(n45862) );
  NOR U58749 ( .A(n45862), .B(n45861), .Z(n49421) );
  IV U58750 ( .A(n45863), .Z(n45864) );
  NOR U58751 ( .A(n45865), .B(n45864), .Z(n49751) );
  NOR U58752 ( .A(n49421), .B(n49751), .Z(n46189) );
  NOR U58753 ( .A(n45867), .B(n45866), .Z(n49423) );
  NOR U58754 ( .A(n49746), .B(n49748), .Z(n46188) );
  IV U58755 ( .A(n45868), .Z(n45869) );
  NOR U58756 ( .A(n45869), .B(n46164), .Z(n49440) );
  IV U58757 ( .A(n45870), .Z(n46162) );
  IV U58758 ( .A(n45871), .Z(n45872) );
  NOR U58759 ( .A(n46162), .B(n45872), .Z(n49444) );
  IV U58760 ( .A(n45873), .Z(n45874) );
  NOR U58761 ( .A(n45875), .B(n45874), .Z(n49731) );
  IV U58762 ( .A(n45876), .Z(n45877) );
  NOR U58763 ( .A(n45877), .B(n45879), .Z(n49728) );
  IV U58764 ( .A(n45878), .Z(n45880) );
  NOR U58765 ( .A(n45880), .B(n45879), .Z(n49726) );
  NOR U58766 ( .A(n45882), .B(n45881), .Z(n45883) );
  NOR U58767 ( .A(n49726), .B(n45883), .Z(n45884) );
  IV U58768 ( .A(n45884), .Z(n45885) );
  NOR U58769 ( .A(n49728), .B(n45885), .Z(n46158) );
  IV U58770 ( .A(n45886), .Z(n49448) );
  IV U58771 ( .A(n45887), .Z(n45889) );
  NOR U58772 ( .A(n45889), .B(n45888), .Z(n46156) );
  IV U58773 ( .A(n46156), .Z(n46147) );
  IV U58774 ( .A(n45890), .Z(n45892) );
  NOR U58775 ( .A(n45892), .B(n45891), .Z(n45893) );
  IV U58776 ( .A(n45893), .Z(n49450) );
  IV U58777 ( .A(n45894), .Z(n45895) );
  NOR U58778 ( .A(n45895), .B(n46143), .Z(n49711) );
  IV U58779 ( .A(n45896), .Z(n45900) );
  IV U58780 ( .A(n45897), .Z(n46137) );
  NOR U58781 ( .A(n45898), .B(n46137), .Z(n45899) );
  IV U58782 ( .A(n45899), .Z(n45902) );
  NOR U58783 ( .A(n45900), .B(n45902), .Z(n49699) );
  IV U58784 ( .A(n45901), .Z(n45903) );
  NOR U58785 ( .A(n45903), .B(n45902), .Z(n49693) );
  NOR U58786 ( .A(n45905), .B(n45904), .Z(n49690) );
  IV U58787 ( .A(n45906), .Z(n45909) );
  IV U58788 ( .A(n45907), .Z(n45908) );
  NOR U58789 ( .A(n45909), .B(n45908), .Z(n49667) );
  IV U58790 ( .A(n45910), .Z(n45911) );
  NOR U58791 ( .A(n45917), .B(n45911), .Z(n46114) );
  IV U58792 ( .A(n46114), .Z(n46112) );
  IV U58793 ( .A(n45912), .Z(n45913) );
  NOR U58794 ( .A(n45917), .B(n45913), .Z(n45914) );
  IV U58795 ( .A(n45914), .Z(n49467) );
  IV U58796 ( .A(n45915), .Z(n45916) );
  NOR U58797 ( .A(n45917), .B(n45916), .Z(n49471) );
  IV U58798 ( .A(n45918), .Z(n45920) );
  IV U58799 ( .A(n45919), .Z(n46107) );
  NOR U58800 ( .A(n45920), .B(n46107), .Z(n49468) );
  IV U58801 ( .A(n45921), .Z(n45922) );
  NOR U58802 ( .A(n45922), .B(n46104), .Z(n49649) );
  IV U58803 ( .A(n45923), .Z(n45925) );
  NOR U58804 ( .A(n45925), .B(n45924), .Z(n45926) );
  IV U58805 ( .A(n45926), .Z(n46097) );
  IV U58806 ( .A(n45927), .Z(n45929) );
  IV U58807 ( .A(n45928), .Z(n45933) );
  NOR U58808 ( .A(n45929), .B(n45933), .Z(n45930) );
  IV U58809 ( .A(n45930), .Z(n49478) );
  IV U58810 ( .A(n45931), .Z(n45932) );
  NOR U58811 ( .A(n45933), .B(n45932), .Z(n49644) );
  NOR U58812 ( .A(n49481), .B(n49644), .Z(n46084) );
  NOR U58813 ( .A(n49487), .B(n45934), .Z(n45937) );
  NOR U58814 ( .A(n45936), .B(n45935), .Z(n49483) );
  NOR U58815 ( .A(n45937), .B(n49483), .Z(n46083) );
  IV U58816 ( .A(n45938), .Z(n45939) );
  NOR U58817 ( .A(n45939), .B(n46081), .Z(n49490) );
  IV U58818 ( .A(n45940), .Z(n45942) );
  NOR U58819 ( .A(n45942), .B(n45941), .Z(n49498) );
  IV U58820 ( .A(n45943), .Z(n45944) );
  NOR U58821 ( .A(n45944), .B(n46062), .Z(n45945) );
  IV U58822 ( .A(n45945), .Z(n46072) );
  IV U58823 ( .A(n45946), .Z(n45947) );
  NOR U58824 ( .A(n45948), .B(n45947), .Z(n45949) );
  IV U58825 ( .A(n45949), .Z(n49635) );
  IV U58826 ( .A(n45950), .Z(n45951) );
  NOR U58827 ( .A(n45951), .B(n45956), .Z(n49513) );
  IV U58828 ( .A(n45952), .Z(n45953) );
  NOR U58829 ( .A(n45954), .B(n45953), .Z(n49616) );
  IV U58830 ( .A(n45955), .Z(n45957) );
  NOR U58831 ( .A(n45957), .B(n45956), .Z(n49619) );
  NOR U58832 ( .A(n49616), .B(n49619), .Z(n46045) );
  NOR U58833 ( .A(n45958), .B(n53373), .Z(n49516) );
  IV U58834 ( .A(n45959), .Z(n45961) );
  NOR U58835 ( .A(n45961), .B(n45960), .Z(n49577) );
  IV U58836 ( .A(n45962), .Z(n45964) );
  NOR U58837 ( .A(n45964), .B(n45963), .Z(n49531) );
  NOR U58838 ( .A(n49577), .B(n49531), .Z(n46024) );
  IV U58839 ( .A(n45965), .Z(n45966) );
  NOR U58840 ( .A(n45967), .B(n45966), .Z(n49580) );
  IV U58841 ( .A(n45968), .Z(n45970) );
  IV U58842 ( .A(n45969), .Z(n45974) );
  NOR U58843 ( .A(n45970), .B(n45974), .Z(n49534) );
  NOR U58844 ( .A(n49580), .B(n49534), .Z(n46023) );
  NOR U58845 ( .A(n45972), .B(n45971), .Z(n49573) );
  IV U58846 ( .A(n45973), .Z(n45975) );
  NOR U58847 ( .A(n45975), .B(n45974), .Z(n49537) );
  NOR U58848 ( .A(n49573), .B(n49537), .Z(n46022) );
  IV U58849 ( .A(n45976), .Z(n45977) );
  NOR U58850 ( .A(n45978), .B(n45977), .Z(n49569) );
  IV U58851 ( .A(n45979), .Z(n45980) );
  NOR U58852 ( .A(n45981), .B(n45980), .Z(n49558) );
  IV U58853 ( .A(n45982), .Z(n45983) );
  NOR U58854 ( .A(n45985), .B(n45983), .Z(n49555) );
  IV U58855 ( .A(n45984), .Z(n45986) );
  NOR U58856 ( .A(n45986), .B(n45985), .Z(n49552) );
  NOR U58857 ( .A(n45987), .B(n45988), .Z(n45994) );
  IV U58858 ( .A(n45988), .Z(n45990) );
  NOR U58859 ( .A(n45990), .B(n45989), .Z(n45991) );
  NOR U58860 ( .A(n45992), .B(n45991), .Z(n45993) );
  NOR U58861 ( .A(n45994), .B(n45993), .Z(n49547) );
  NOR U58862 ( .A(n45999), .B(n45998), .Z(n46006) );
  NOR U58863 ( .A(n46001), .B(n46000), .Z(n46004) );
  IV U58864 ( .A(n46002), .Z(n46003) );
  NOR U58865 ( .A(n46004), .B(n46003), .Z(n46005) );
  NOR U58866 ( .A(n46006), .B(n46005), .Z(n49544) );
  XOR U58867 ( .A(n49546), .B(n49544), .Z(n49548) );
  XOR U58868 ( .A(n49547), .B(n49548), .Z(n49553) );
  XOR U58869 ( .A(n49552), .B(n49553), .Z(n49557) );
  XOR U58870 ( .A(n49555), .B(n49557), .Z(n49559) );
  XOR U58871 ( .A(n49558), .B(n49559), .Z(n46010) );
  IV U58872 ( .A(n46007), .Z(n46008) );
  NOR U58873 ( .A(n46008), .B(n46020), .Z(n46016) );
  IV U58874 ( .A(n46016), .Z(n46009) );
  NOR U58875 ( .A(n46010), .B(n46009), .Z(n49543) );
  IV U58876 ( .A(n46011), .Z(n46012) );
  NOR U58877 ( .A(n46013), .B(n46012), .Z(n49540) );
  NOR U58878 ( .A(n49558), .B(n49540), .Z(n46014) );
  XOR U58879 ( .A(n49559), .B(n46014), .Z(n46015) );
  NOR U58880 ( .A(n46016), .B(n46015), .Z(n46017) );
  NOR U58881 ( .A(n49543), .B(n46017), .Z(n46018) );
  IV U58882 ( .A(n46018), .Z(n49568) );
  IV U58883 ( .A(n46019), .Z(n46021) );
  NOR U58884 ( .A(n46021), .B(n46020), .Z(n49566) );
  XOR U58885 ( .A(n49568), .B(n49566), .Z(n49574) );
  XOR U58886 ( .A(n49569), .B(n49574), .Z(n49539) );
  XOR U58887 ( .A(n46022), .B(n49539), .Z(n49533) );
  XOR U58888 ( .A(n46023), .B(n49533), .Z(n49578) );
  XOR U58889 ( .A(n46024), .B(n49578), .Z(n49529) );
  NOR U58890 ( .A(n49605), .B(n49603), .Z(n46028) );
  IV U58891 ( .A(n46025), .Z(n46026) );
  NOR U58892 ( .A(n46027), .B(n46026), .Z(n49528) );
  NOR U58893 ( .A(n46028), .B(n49528), .Z(n46029) );
  XOR U58894 ( .A(n49529), .B(n46029), .Z(n49601) );
  IV U58895 ( .A(n46030), .Z(n46032) );
  NOR U58896 ( .A(n46032), .B(n46031), .Z(n49599) );
  NOR U58897 ( .A(n46034), .B(n46033), .Z(n49526) );
  NOR U58898 ( .A(n49599), .B(n49526), .Z(n46035) );
  XOR U58899 ( .A(n49601), .B(n46035), .Z(n49519) );
  IV U58900 ( .A(n46036), .Z(n46038) );
  NOR U58901 ( .A(n46038), .B(n46037), .Z(n49518) );
  IV U58902 ( .A(n46039), .Z(n46040) );
  NOR U58903 ( .A(n46041), .B(n46040), .Z(n49521) );
  NOR U58904 ( .A(n49523), .B(n49521), .Z(n46042) );
  IV U58905 ( .A(n46042), .Z(n46043) );
  NOR U58906 ( .A(n49518), .B(n46043), .Z(n46044) );
  XOR U58907 ( .A(n49519), .B(n46044), .Z(n53370) );
  XOR U58908 ( .A(n49516), .B(n53370), .Z(n49620) );
  XOR U58909 ( .A(n46045), .B(n49620), .Z(n46046) );
  IV U58910 ( .A(n46046), .Z(n49515) );
  XOR U58911 ( .A(n49513), .B(n49515), .Z(n49512) );
  IV U58912 ( .A(n46047), .Z(n46049) );
  NOR U58913 ( .A(n46049), .B(n46048), .Z(n49510) );
  XOR U58914 ( .A(n49512), .B(n49510), .Z(n49506) );
  IV U58915 ( .A(n49506), .Z(n46056) );
  IV U58916 ( .A(n46050), .Z(n46051) );
  NOR U58917 ( .A(n46052), .B(n46051), .Z(n49508) );
  IV U58918 ( .A(n46053), .Z(n46054) );
  NOR U58919 ( .A(n46054), .B(n46058), .Z(n49504) );
  NOR U58920 ( .A(n49508), .B(n49504), .Z(n46055) );
  XOR U58921 ( .A(n46056), .B(n46055), .Z(n49633) );
  IV U58922 ( .A(n46057), .Z(n46059) );
  NOR U58923 ( .A(n46059), .B(n46058), .Z(n49631) );
  XOR U58924 ( .A(n49633), .B(n49631), .Z(n49634) );
  XOR U58925 ( .A(n49635), .B(n49634), .Z(n46069) );
  IV U58926 ( .A(n46069), .Z(n46060) );
  NOR U58927 ( .A(n46072), .B(n46060), .Z(n53292) );
  IV U58928 ( .A(n46061), .Z(n46063) );
  NOR U58929 ( .A(n46063), .B(n46062), .Z(n46064) );
  IV U58930 ( .A(n46064), .Z(n49503) );
  IV U58931 ( .A(n46065), .Z(n46067) );
  NOR U58932 ( .A(n46067), .B(n46066), .Z(n46070) );
  IV U58933 ( .A(n46070), .Z(n46068) );
  NOR U58934 ( .A(n46068), .B(n49634), .Z(n53289) );
  NOR U58935 ( .A(n46070), .B(n46069), .Z(n46071) );
  NOR U58936 ( .A(n53289), .B(n46071), .Z(n46073) );
  IV U58937 ( .A(n46073), .Z(n49502) );
  XOR U58938 ( .A(n49503), .B(n49502), .Z(n46075) );
  NOR U58939 ( .A(n46073), .B(n46072), .Z(n46074) );
  NOR U58940 ( .A(n46075), .B(n46074), .Z(n46076) );
  NOR U58941 ( .A(n53292), .B(n46076), .Z(n49496) );
  IV U58942 ( .A(n46077), .Z(n46079) );
  NOR U58943 ( .A(n46079), .B(n46078), .Z(n53420) );
  IV U58944 ( .A(n46080), .Z(n46082) );
  NOR U58945 ( .A(n46082), .B(n46081), .Z(n53284) );
  NOR U58946 ( .A(n53420), .B(n53284), .Z(n49497) );
  XOR U58947 ( .A(n49496), .B(n49497), .Z(n49500) );
  XOR U58948 ( .A(n49498), .B(n49500), .Z(n49491) );
  XOR U58949 ( .A(n49490), .B(n49491), .Z(n49486) );
  XOR U58950 ( .A(n46083), .B(n49486), .Z(n49480) );
  XOR U58951 ( .A(n46084), .B(n49480), .Z(n49477) );
  XOR U58952 ( .A(n49478), .B(n49477), .Z(n46094) );
  IV U58953 ( .A(n46094), .Z(n46085) );
  NOR U58954 ( .A(n46097), .B(n46085), .Z(n53262) );
  IV U58955 ( .A(n46086), .Z(n46087) );
  NOR U58956 ( .A(n46088), .B(n46087), .Z(n46089) );
  IV U58957 ( .A(n46089), .Z(n49658) );
  IV U58958 ( .A(n46090), .Z(n46091) );
  NOR U58959 ( .A(n46092), .B(n46091), .Z(n46095) );
  IV U58960 ( .A(n46095), .Z(n46093) );
  NOR U58961 ( .A(n46093), .B(n49477), .Z(n53264) );
  NOR U58962 ( .A(n46095), .B(n46094), .Z(n46096) );
  NOR U58963 ( .A(n53264), .B(n46096), .Z(n46098) );
  IV U58964 ( .A(n46098), .Z(n49657) );
  XOR U58965 ( .A(n49658), .B(n49657), .Z(n46100) );
  NOR U58966 ( .A(n46098), .B(n46097), .Z(n46099) );
  NOR U58967 ( .A(n46100), .B(n46099), .Z(n46101) );
  NOR U58968 ( .A(n53262), .B(n46101), .Z(n46102) );
  IV U58969 ( .A(n46102), .Z(n49650) );
  XOR U58970 ( .A(n49649), .B(n49650), .Z(n49654) );
  IV U58971 ( .A(n49654), .Z(n46110) );
  IV U58972 ( .A(n46103), .Z(n46105) );
  NOR U58973 ( .A(n46105), .B(n46104), .Z(n49653) );
  IV U58974 ( .A(n46106), .Z(n46108) );
  NOR U58975 ( .A(n46108), .B(n46107), .Z(n49474) );
  NOR U58976 ( .A(n49653), .B(n49474), .Z(n46109) );
  XOR U58977 ( .A(n46110), .B(n46109), .Z(n49470) );
  XOR U58978 ( .A(n49468), .B(n49470), .Z(n49472) );
  XOR U58979 ( .A(n49471), .B(n49472), .Z(n49466) );
  XOR U58980 ( .A(n49467), .B(n49466), .Z(n46113) );
  IV U58981 ( .A(n46113), .Z(n46111) );
  NOR U58982 ( .A(n46112), .B(n46111), .Z(n53253) );
  NOR U58983 ( .A(n46114), .B(n46113), .Z(n49465) );
  NOR U58984 ( .A(n46115), .B(n46118), .Z(n49463) );
  XOR U58985 ( .A(n49465), .B(n49463), .Z(n46116) );
  NOR U58986 ( .A(n53253), .B(n46116), .Z(n49672) );
  IV U58987 ( .A(n46117), .Z(n46119) );
  NOR U58988 ( .A(n46119), .B(n46118), .Z(n46120) );
  IV U58989 ( .A(n46120), .Z(n49673) );
  XOR U58990 ( .A(n49672), .B(n49673), .Z(n49668) );
  XOR U58991 ( .A(n49667), .B(n49668), .Z(n49684) );
  IV U58992 ( .A(n46121), .Z(n46122) );
  NOR U58993 ( .A(n46123), .B(n46122), .Z(n49683) );
  NOR U58994 ( .A(n49683), .B(n49461), .Z(n46124) );
  XOR U58995 ( .A(n49684), .B(n46124), .Z(n49457) );
  NOR U58996 ( .A(n46126), .B(n46125), .Z(n49456) );
  IV U58997 ( .A(n46127), .Z(n46128) );
  NOR U58998 ( .A(n46129), .B(n46128), .Z(n49459) );
  IV U58999 ( .A(n46130), .Z(n46132) );
  NOR U59000 ( .A(n46132), .B(n46131), .Z(n49686) );
  NOR U59001 ( .A(n49459), .B(n49686), .Z(n46133) );
  XOR U59002 ( .A(n49456), .B(n46133), .Z(n46134) );
  XOR U59003 ( .A(n49457), .B(n46134), .Z(n49692) );
  XOR U59004 ( .A(n49690), .B(n49692), .Z(n49694) );
  XOR U59005 ( .A(n49693), .B(n49694), .Z(n49700) );
  XOR U59006 ( .A(n49699), .B(n49700), .Z(n49455) );
  IV U59007 ( .A(n46135), .Z(n46136) );
  NOR U59008 ( .A(n46137), .B(n46136), .Z(n49453) );
  XOR U59009 ( .A(n49455), .B(n49453), .Z(n49715) );
  IV U59010 ( .A(n49715), .Z(n46145) );
  IV U59011 ( .A(n46138), .Z(n46139) );
  NOR U59012 ( .A(n46140), .B(n46139), .Z(n49451) );
  IV U59013 ( .A(n46141), .Z(n46142) );
  NOR U59014 ( .A(n46143), .B(n46142), .Z(n49714) );
  NOR U59015 ( .A(n49451), .B(n49714), .Z(n46144) );
  XOR U59016 ( .A(n46145), .B(n46144), .Z(n49713) );
  XOR U59017 ( .A(n49711), .B(n49713), .Z(n49449) );
  XOR U59018 ( .A(n49450), .B(n49449), .Z(n46152) );
  IV U59019 ( .A(n46152), .Z(n46146) );
  NOR U59020 ( .A(n46147), .B(n46146), .Z(n53478) );
  IV U59021 ( .A(n46148), .Z(n46149) );
  NOR U59022 ( .A(n46150), .B(n46149), .Z(n46153) );
  IV U59023 ( .A(n46153), .Z(n46151) );
  NOR U59024 ( .A(n46151), .B(n49449), .Z(n53475) );
  NOR U59025 ( .A(n46153), .B(n46152), .Z(n46154) );
  NOR U59026 ( .A(n53475), .B(n46154), .Z(n46155) );
  NOR U59027 ( .A(n46156), .B(n46155), .Z(n46157) );
  NOR U59028 ( .A(n53478), .B(n46157), .Z(n49447) );
  XOR U59029 ( .A(n49448), .B(n49447), .Z(n49720) );
  XOR U59030 ( .A(n46158), .B(n49720), .Z(n46159) );
  IV U59031 ( .A(n46159), .Z(n49733) );
  XOR U59032 ( .A(n49731), .B(n49733), .Z(n49445) );
  XOR U59033 ( .A(n49444), .B(n49445), .Z(n49742) );
  IV U59034 ( .A(n46160), .Z(n46161) );
  NOR U59035 ( .A(n46162), .B(n46161), .Z(n49734) );
  IV U59036 ( .A(n46163), .Z(n46165) );
  NOR U59037 ( .A(n46165), .B(n46164), .Z(n49740) );
  NOR U59038 ( .A(n49734), .B(n49740), .Z(n46166) );
  XOR U59039 ( .A(n49742), .B(n46166), .Z(n46167) );
  IV U59040 ( .A(n46167), .Z(n49443) );
  XOR U59041 ( .A(n49440), .B(n49443), .Z(n49439) );
  IV U59042 ( .A(n46168), .Z(n46170) );
  NOR U59043 ( .A(n46170), .B(n46169), .Z(n49441) );
  IV U59044 ( .A(n46171), .Z(n46172) );
  NOR U59045 ( .A(n46173), .B(n46172), .Z(n49437) );
  NOR U59046 ( .A(n49441), .B(n49437), .Z(n46174) );
  XOR U59047 ( .A(n49439), .B(n46174), .Z(n49429) );
  IV U59048 ( .A(n46175), .Z(n46176) );
  NOR U59049 ( .A(n46177), .B(n46176), .Z(n49434) );
  IV U59050 ( .A(n46178), .Z(n46179) );
  NOR U59051 ( .A(n46180), .B(n46179), .Z(n49428) );
  NOR U59052 ( .A(n49434), .B(n49428), .Z(n46181) );
  XOR U59053 ( .A(n49429), .B(n46181), .Z(n49432) );
  IV U59054 ( .A(n46182), .Z(n46183) );
  NOR U59055 ( .A(n46184), .B(n46183), .Z(n49431) );
  NOR U59056 ( .A(n46186), .B(n46185), .Z(n49426) );
  NOR U59057 ( .A(n49431), .B(n49426), .Z(n46187) );
  XOR U59058 ( .A(n49432), .B(n46187), .Z(n49420) );
  XOR U59059 ( .A(n46188), .B(n49420), .Z(n49424) );
  XOR U59060 ( .A(n49423), .B(n49424), .Z(n49752) );
  XOR U59061 ( .A(n46189), .B(n49752), .Z(n49413) );
  XOR U59062 ( .A(n46190), .B(n49413), .Z(n49757) );
  XOR U59063 ( .A(n49409), .B(n49757), .Z(n46191) );
  XOR U59064 ( .A(n46192), .B(n46191), .Z(n46193) );
  IV U59065 ( .A(n46193), .Z(n49407) );
  IV U59066 ( .A(n46194), .Z(n46200) );
  IV U59067 ( .A(n46195), .Z(n46196) );
  NOR U59068 ( .A(n46200), .B(n46196), .Z(n46202) );
  IV U59069 ( .A(n46202), .Z(n46197) );
  NOR U59070 ( .A(n49407), .B(n46197), .Z(n53174) );
  IV U59071 ( .A(n46198), .Z(n46199) );
  NOR U59072 ( .A(n46200), .B(n46199), .Z(n49405) );
  XOR U59073 ( .A(n49405), .B(n49407), .Z(n46206) );
  IV U59074 ( .A(n46206), .Z(n46201) );
  NOR U59075 ( .A(n46202), .B(n46201), .Z(n46203) );
  NOR U59076 ( .A(n53174), .B(n46203), .Z(n46204) );
  NOR U59077 ( .A(n46205), .B(n46204), .Z(n46208) );
  IV U59078 ( .A(n46205), .Z(n46207) );
  NOR U59079 ( .A(n46207), .B(n46206), .Z(n53179) );
  NOR U59080 ( .A(n46208), .B(n53179), .Z(n49402) );
  IV U59081 ( .A(n46209), .Z(n46210) );
  NOR U59082 ( .A(n46211), .B(n46210), .Z(n46212) );
  IV U59083 ( .A(n46212), .Z(n49403) );
  XOR U59084 ( .A(n49402), .B(n49403), .Z(n49400) );
  NOR U59085 ( .A(n46213), .B(n49400), .Z(n53515) );
  IV U59086 ( .A(n46214), .Z(n46216) );
  NOR U59087 ( .A(n46216), .B(n46215), .Z(n49399) );
  XOR U59088 ( .A(n49399), .B(n49400), .Z(n46225) );
  IV U59089 ( .A(n46225), .Z(n46217) );
  NOR U59090 ( .A(n46218), .B(n46217), .Z(n46219) );
  NOR U59091 ( .A(n53515), .B(n46219), .Z(n46227) );
  IV U59092 ( .A(n46227), .Z(n46220) );
  NOR U59093 ( .A(n46221), .B(n46220), .Z(n53521) );
  IV U59094 ( .A(n46222), .Z(n46224) );
  NOR U59095 ( .A(n46224), .B(n46223), .Z(n46228) );
  IV U59096 ( .A(n46228), .Z(n46226) );
  NOR U59097 ( .A(n46226), .B(n46225), .Z(n53171) );
  NOR U59098 ( .A(n46228), .B(n46227), .Z(n46229) );
  NOR U59099 ( .A(n53171), .B(n46229), .Z(n46230) );
  NOR U59100 ( .A(n46231), .B(n46230), .Z(n46232) );
  NOR U59101 ( .A(n53521), .B(n46232), .Z(n49397) );
  IV U59102 ( .A(n46233), .Z(n46234) );
  NOR U59103 ( .A(n46235), .B(n46234), .Z(n49396) );
  IV U59104 ( .A(n46236), .Z(n46240) );
  NOR U59105 ( .A(n46237), .B(n46248), .Z(n46238) );
  IV U59106 ( .A(n46238), .Z(n46239) );
  NOR U59107 ( .A(n46240), .B(n46239), .Z(n49761) );
  NOR U59108 ( .A(n49396), .B(n49761), .Z(n46241) );
  XOR U59109 ( .A(n49397), .B(n46241), .Z(n49395) );
  IV U59110 ( .A(n46242), .Z(n46243) );
  NOR U59111 ( .A(n46244), .B(n46243), .Z(n46254) );
  IV U59112 ( .A(n46254), .Z(n46245) );
  NOR U59113 ( .A(n49395), .B(n46245), .Z(n53162) );
  IV U59114 ( .A(n46246), .Z(n46252) );
  IV U59115 ( .A(n46247), .Z(n46249) );
  NOR U59116 ( .A(n46249), .B(n46248), .Z(n46250) );
  IV U59117 ( .A(n46250), .Z(n46251) );
  NOR U59118 ( .A(n46252), .B(n46251), .Z(n49393) );
  XOR U59119 ( .A(n49393), .B(n49395), .Z(n49390) );
  IV U59120 ( .A(n49390), .Z(n46253) );
  NOR U59121 ( .A(n46254), .B(n46253), .Z(n46255) );
  NOR U59122 ( .A(n53162), .B(n46255), .Z(n49385) );
  XOR U59123 ( .A(n46256), .B(n49385), .Z(n49382) );
  XOR U59124 ( .A(n49380), .B(n49382), .Z(n53537) );
  IV U59125 ( .A(n53537), .Z(n46263) );
  IV U59126 ( .A(n46257), .Z(n46258) );
  NOR U59127 ( .A(n46259), .B(n46258), .Z(n53542) );
  IV U59128 ( .A(n46260), .Z(n46262) );
  NOR U59129 ( .A(n46262), .B(n46261), .Z(n53543) );
  NOR U59130 ( .A(n53542), .B(n53543), .Z(n49383) );
  XOR U59131 ( .A(n46263), .B(n49383), .Z(n49770) );
  XOR U59132 ( .A(n49768), .B(n49770), .Z(n46264) );
  NOR U59133 ( .A(n46265), .B(n46264), .Z(n53547) );
  IV U59134 ( .A(n46266), .Z(n46267) );
  NOR U59135 ( .A(n46268), .B(n46267), .Z(n49769) );
  NOR U59136 ( .A(n49769), .B(n49768), .Z(n46269) );
  XOR U59137 ( .A(n49770), .B(n46269), .Z(n46270) );
  NOR U59138 ( .A(n46271), .B(n46270), .Z(n46272) );
  NOR U59139 ( .A(n53547), .B(n46272), .Z(n46273) );
  IV U59140 ( .A(n46273), .Z(n49776) );
  XOR U59141 ( .A(n49775), .B(n49776), .Z(n49371) );
  IV U59142 ( .A(n49371), .Z(n46281) );
  IV U59143 ( .A(n46274), .Z(n49374) );
  NOR U59144 ( .A(n46275), .B(n49374), .Z(n46279) );
  IV U59145 ( .A(n46276), .Z(n46278) );
  NOR U59146 ( .A(n46278), .B(n46277), .Z(n49370) );
  NOR U59147 ( .A(n46279), .B(n49370), .Z(n46280) );
  XOR U59148 ( .A(n46281), .B(n46280), .Z(n49366) );
  XOR U59149 ( .A(n49364), .B(n49366), .Z(n49368) );
  XOR U59150 ( .A(n46282), .B(n49368), .Z(n46283) );
  IV U59151 ( .A(n46283), .Z(n49362) );
  XOR U59152 ( .A(n49361), .B(n49362), .Z(n56608) );
  XOR U59153 ( .A(n56607), .B(n56608), .Z(n57030) );
  IV U59154 ( .A(n57030), .Z(n46290) );
  IV U59155 ( .A(n46284), .Z(n46286) );
  NOR U59156 ( .A(n46286), .B(n46285), .Z(n49357) );
  IV U59157 ( .A(n46287), .Z(n46289) );
  NOR U59158 ( .A(n46289), .B(n46288), .Z(n49354) );
  NOR U59159 ( .A(n49357), .B(n49354), .Z(n57031) );
  XOR U59160 ( .A(n46290), .B(n57031), .Z(n49351) );
  NOR U59161 ( .A(n46291), .B(n49351), .Z(n49353) );
  IV U59162 ( .A(n46292), .Z(n46293) );
  NOR U59163 ( .A(n46294), .B(n46293), .Z(n46300) );
  IV U59164 ( .A(n46300), .Z(n46298) );
  IV U59165 ( .A(n46295), .Z(n46296) );
  NOR U59166 ( .A(n46297), .B(n46296), .Z(n49350) );
  XOR U59167 ( .A(n49350), .B(n49351), .Z(n46299) );
  NOR U59168 ( .A(n46298), .B(n46299), .Z(n49348) );
  NOR U59169 ( .A(n49353), .B(n49348), .Z(n53130) );
  IV U59170 ( .A(n53130), .Z(n46302) );
  NOR U59171 ( .A(n46302), .B(n46299), .Z(n46305) );
  NOR U59172 ( .A(n46301), .B(n46300), .Z(n46303) );
  NOR U59173 ( .A(n46303), .B(n46302), .Z(n46304) );
  NOR U59174 ( .A(n46305), .B(n46304), .Z(n49346) );
  XOR U59175 ( .A(n49345), .B(n49346), .Z(n46314) );
  XOR U59176 ( .A(n49344), .B(n46314), .Z(n46316) );
  IV U59177 ( .A(n46316), .Z(n46306) );
  NOR U59178 ( .A(n46307), .B(n46306), .Z(n53118) );
  IV U59179 ( .A(n46308), .Z(n46310) );
  IV U59180 ( .A(n46309), .Z(n46313) );
  NOR U59181 ( .A(n46310), .B(n46313), .Z(n49341) );
  IV U59182 ( .A(n46311), .Z(n46312) );
  NOR U59183 ( .A(n46313), .B(n46312), .Z(n46317) );
  IV U59184 ( .A(n46317), .Z(n46315) );
  NOR U59185 ( .A(n46315), .B(n46314), .Z(n53122) );
  NOR U59186 ( .A(n46317), .B(n46316), .Z(n46318) );
  NOR U59187 ( .A(n53122), .B(n46318), .Z(n46319) );
  IV U59188 ( .A(n46319), .Z(n49342) );
  XOR U59189 ( .A(n49341), .B(n49342), .Z(n49787) );
  IV U59190 ( .A(n49787), .Z(n46320) );
  NOR U59191 ( .A(n46321), .B(n46320), .Z(n46322) );
  NOR U59192 ( .A(n53118), .B(n46322), .Z(n49792) );
  IV U59193 ( .A(n46323), .Z(n46325) );
  NOR U59194 ( .A(n46325), .B(n46324), .Z(n49786) );
  IV U59195 ( .A(n49332), .Z(n46326) );
  NOR U59196 ( .A(n46326), .B(n49331), .Z(n49791) );
  NOR U59197 ( .A(n49786), .B(n49791), .Z(n46327) );
  XOR U59198 ( .A(n49792), .B(n46327), .Z(n49334) );
  NOR U59199 ( .A(n46328), .B(n49331), .Z(n46332) );
  IV U59200 ( .A(n46329), .Z(n46331) );
  IV U59201 ( .A(n46330), .Z(n46335) );
  NOR U59202 ( .A(n46331), .B(n46335), .Z(n49328) );
  NOR U59203 ( .A(n46332), .B(n49328), .Z(n46333) );
  XOR U59204 ( .A(n49334), .B(n46333), .Z(n49318) );
  IV U59205 ( .A(n46334), .Z(n46336) );
  NOR U59206 ( .A(n46336), .B(n46335), .Z(n49325) );
  IV U59207 ( .A(n46337), .Z(n46339) );
  NOR U59208 ( .A(n46339), .B(n46338), .Z(n49317) );
  NOR U59209 ( .A(n49325), .B(n49317), .Z(n46340) );
  XOR U59210 ( .A(n49318), .B(n46340), .Z(n49322) );
  XOR U59211 ( .A(n49320), .B(n49322), .Z(n49315) );
  XOR U59212 ( .A(n49316), .B(n49315), .Z(n46341) );
  IV U59213 ( .A(n46341), .Z(n49312) );
  XOR U59214 ( .A(n49311), .B(n49312), .Z(n46352) );
  IV U59215 ( .A(n46352), .Z(n46350) );
  IV U59216 ( .A(n46342), .Z(n46344) );
  NOR U59217 ( .A(n46344), .B(n46343), .Z(n46354) );
  IV U59218 ( .A(n46345), .Z(n46347) );
  NOR U59219 ( .A(n46347), .B(n46346), .Z(n46351) );
  NOR U59220 ( .A(n46354), .B(n46351), .Z(n46348) );
  IV U59221 ( .A(n46348), .Z(n46349) );
  NOR U59222 ( .A(n46350), .B(n46349), .Z(n46357) );
  IV U59223 ( .A(n46351), .Z(n46353) );
  NOR U59224 ( .A(n46353), .B(n46352), .Z(n53591) );
  IV U59225 ( .A(n46354), .Z(n46355) );
  NOR U59226 ( .A(n46355), .B(n49312), .Z(n53577) );
  NOR U59227 ( .A(n53591), .B(n53577), .Z(n46356) );
  IV U59228 ( .A(n46356), .Z(n49314) );
  NOR U59229 ( .A(n46357), .B(n49314), .Z(n46358) );
  IV U59230 ( .A(n46358), .Z(n49307) );
  NOR U59231 ( .A(n46359), .B(n49308), .Z(n46360) );
  XOR U59232 ( .A(n49307), .B(n46360), .Z(n49805) );
  IV U59233 ( .A(n46361), .Z(n46363) );
  NOR U59234 ( .A(n46363), .B(n46362), .Z(n49304) );
  IV U59235 ( .A(n46364), .Z(n46366) );
  NOR U59236 ( .A(n46366), .B(n46365), .Z(n49804) );
  NOR U59237 ( .A(n49304), .B(n49804), .Z(n46367) );
  XOR U59238 ( .A(n49805), .B(n46367), .Z(n49298) );
  IV U59239 ( .A(n46368), .Z(n46370) );
  NOR U59240 ( .A(n46370), .B(n46369), .Z(n49801) );
  IV U59241 ( .A(n46371), .Z(n46373) );
  NOR U59242 ( .A(n46373), .B(n46372), .Z(n49299) );
  NOR U59243 ( .A(n49801), .B(n49299), .Z(n46374) );
  XOR U59244 ( .A(n49298), .B(n46374), .Z(n49302) );
  IV U59245 ( .A(n46375), .Z(n46377) );
  NOR U59246 ( .A(n46377), .B(n46376), .Z(n49301) );
  IV U59247 ( .A(n46378), .Z(n46380) );
  NOR U59248 ( .A(n46380), .B(n46379), .Z(n49294) );
  NOR U59249 ( .A(n49301), .B(n49294), .Z(n46381) );
  XOR U59250 ( .A(n49302), .B(n46381), .Z(n49290) );
  IV U59251 ( .A(n46382), .Z(n46384) );
  NOR U59252 ( .A(n46384), .B(n46383), .Z(n49814) );
  IV U59253 ( .A(n46385), .Z(n46386) );
  NOR U59254 ( .A(n46387), .B(n46386), .Z(n49296) );
  IV U59255 ( .A(n46388), .Z(n46390) );
  NOR U59256 ( .A(n46390), .B(n46389), .Z(n49291) );
  NOR U59257 ( .A(n49296), .B(n49291), .Z(n46391) );
  IV U59258 ( .A(n46391), .Z(n46392) );
  NOR U59259 ( .A(n49814), .B(n46392), .Z(n46393) );
  XOR U59260 ( .A(n49290), .B(n46393), .Z(n49287) );
  XOR U59261 ( .A(n49286), .B(n49287), .Z(n53067) );
  IV U59262 ( .A(n46394), .Z(n46395) );
  NOR U59263 ( .A(n46396), .B(n46395), .Z(n46397) );
  NOR U59264 ( .A(n49811), .B(n46397), .Z(n53068) );
  XOR U59265 ( .A(n53067), .B(n53068), .Z(n49824) );
  XOR U59266 ( .A(n46398), .B(n49824), .Z(n49832) );
  XOR U59267 ( .A(n49830), .B(n49832), .Z(n49834) );
  IV U59268 ( .A(n49834), .Z(n46406) );
  IV U59269 ( .A(n46399), .Z(n46400) );
  NOR U59270 ( .A(n46401), .B(n46400), .Z(n49280) );
  IV U59271 ( .A(n46402), .Z(n46404) );
  NOR U59272 ( .A(n46404), .B(n46403), .Z(n49833) );
  NOR U59273 ( .A(n49280), .B(n49833), .Z(n46405) );
  XOR U59274 ( .A(n46406), .B(n46405), .Z(n49274) );
  XOR U59275 ( .A(n49273), .B(n49274), .Z(n49841) );
  XOR U59276 ( .A(n46407), .B(n49841), .Z(n46408) );
  IV U59277 ( .A(n46408), .Z(n49839) );
  XOR U59278 ( .A(n49837), .B(n49839), .Z(n49272) );
  IV U59279 ( .A(n46409), .Z(n46411) );
  NOR U59280 ( .A(n46411), .B(n46410), .Z(n49270) );
  XOR U59281 ( .A(n49272), .B(n49270), .Z(n49265) );
  IV U59282 ( .A(n49265), .Z(n46419) );
  IV U59283 ( .A(n46412), .Z(n46413) );
  NOR U59284 ( .A(n46414), .B(n46413), .Z(n49268) );
  IV U59285 ( .A(n46415), .Z(n46416) );
  NOR U59286 ( .A(n46417), .B(n46416), .Z(n49264) );
  NOR U59287 ( .A(n49268), .B(n49264), .Z(n46418) );
  XOR U59288 ( .A(n46419), .B(n46418), .Z(n49258) );
  XOR U59289 ( .A(n46420), .B(n49258), .Z(n46427) );
  IV U59290 ( .A(n46427), .Z(n46424) );
  IV U59291 ( .A(n46421), .Z(n46434) );
  NOR U59292 ( .A(n46422), .B(n46434), .Z(n46423) );
  NOR U59293 ( .A(n46424), .B(n46423), .Z(n46437) );
  IV U59294 ( .A(n46425), .Z(n46426) );
  NOR U59295 ( .A(n46427), .B(n46426), .Z(n46428) );
  IV U59296 ( .A(n46428), .Z(n46429) );
  NOR U59297 ( .A(n46434), .B(n46429), .Z(n53041) );
  IV U59298 ( .A(n46430), .Z(n46431) );
  NOR U59299 ( .A(n49258), .B(n46431), .Z(n46432) );
  IV U59300 ( .A(n46432), .Z(n46433) );
  NOR U59301 ( .A(n46434), .B(n46433), .Z(n53038) );
  NOR U59302 ( .A(n53041), .B(n53038), .Z(n46435) );
  IV U59303 ( .A(n46435), .Z(n46436) );
  NOR U59304 ( .A(n46437), .B(n46436), .Z(n49253) );
  XOR U59305 ( .A(n46438), .B(n49253), .Z(n49241) );
  XOR U59306 ( .A(n49239), .B(n49241), .Z(n49244) );
  IV U59307 ( .A(n46439), .Z(n46441) );
  NOR U59308 ( .A(n46441), .B(n46440), .Z(n49242) );
  XOR U59309 ( .A(n49244), .B(n49242), .Z(n53023) );
  XOR U59310 ( .A(n49854), .B(n53023), .Z(n49849) );
  XOR U59311 ( .A(n49853), .B(n49849), .Z(n49237) );
  IV U59312 ( .A(n46442), .Z(n46444) );
  NOR U59313 ( .A(n46444), .B(n46443), .Z(n46445) );
  IV U59314 ( .A(n46445), .Z(n49236) );
  XOR U59315 ( .A(n49237), .B(n49236), .Z(n49865) );
  IV U59316 ( .A(n46446), .Z(n46448) );
  NOR U59317 ( .A(n46448), .B(n46447), .Z(n49868) );
  IV U59318 ( .A(n46449), .Z(n46458) );
  IV U59319 ( .A(n46450), .Z(n46451) );
  NOR U59320 ( .A(n46458), .B(n46451), .Z(n49235) );
  NOR U59321 ( .A(n49868), .B(n49235), .Z(n49872) );
  XOR U59322 ( .A(n49865), .B(n49872), .Z(n49233) );
  NOR U59323 ( .A(n46459), .B(n49233), .Z(n53016) );
  IV U59324 ( .A(n46452), .Z(n46454) );
  NOR U59325 ( .A(n46454), .B(n46453), .Z(n46455) );
  IV U59326 ( .A(n46455), .Z(n49231) );
  IV U59327 ( .A(n46456), .Z(n46457) );
  NOR U59328 ( .A(n46458), .B(n46457), .Z(n49232) );
  XOR U59329 ( .A(n49232), .B(n49233), .Z(n49230) );
  XOR U59330 ( .A(n49231), .B(n49230), .Z(n46462) );
  IV U59331 ( .A(n49230), .Z(n46460) );
  NOR U59332 ( .A(n46460), .B(n46459), .Z(n46461) );
  NOR U59333 ( .A(n46462), .B(n46461), .Z(n46463) );
  NOR U59334 ( .A(n53016), .B(n46463), .Z(n46464) );
  IV U59335 ( .A(n46464), .Z(n49224) );
  IV U59336 ( .A(n46465), .Z(n46467) );
  NOR U59337 ( .A(n46467), .B(n46466), .Z(n49222) );
  XOR U59338 ( .A(n49224), .B(n49222), .Z(n49227) );
  XOR U59339 ( .A(n49225), .B(n49227), .Z(n53013) );
  XOR U59340 ( .A(n49217), .B(n53013), .Z(n49215) );
  IV U59341 ( .A(n46468), .Z(n46470) );
  NOR U59342 ( .A(n46470), .B(n46469), .Z(n49218) );
  IV U59343 ( .A(n46471), .Z(n46473) );
  NOR U59344 ( .A(n46473), .B(n46472), .Z(n49214) );
  NOR U59345 ( .A(n49218), .B(n49214), .Z(n46474) );
  XOR U59346 ( .A(n49215), .B(n46474), .Z(n49884) );
  XOR U59347 ( .A(n49883), .B(n49884), .Z(n49887) );
  XOR U59348 ( .A(n46475), .B(n49887), .Z(n49211) );
  IV U59349 ( .A(n46476), .Z(n46477) );
  NOR U59350 ( .A(n46477), .B(n46480), .Z(n46478) );
  IV U59351 ( .A(n46478), .Z(n49212) );
  XOR U59352 ( .A(n49211), .B(n49212), .Z(n49894) );
  IV U59353 ( .A(n46479), .Z(n46481) );
  NOR U59354 ( .A(n46481), .B(n46480), .Z(n49892) );
  XOR U59355 ( .A(n49894), .B(n49892), .Z(n49207) );
  XOR U59356 ( .A(n49206), .B(n49207), .Z(n49204) );
  XOR U59357 ( .A(n49203), .B(n49204), .Z(n49905) );
  XOR U59358 ( .A(n49904), .B(n49905), .Z(n49187) );
  IV U59359 ( .A(n49187), .Z(n46487) );
  IV U59360 ( .A(n46482), .Z(n46483) );
  NOR U59361 ( .A(n46484), .B(n46483), .Z(n49186) );
  NOR U59362 ( .A(n46485), .B(n49186), .Z(n46486) );
  XOR U59363 ( .A(n46487), .B(n46486), .Z(n49185) );
  IV U59364 ( .A(n46488), .Z(n46490) );
  NOR U59365 ( .A(n46490), .B(n46489), .Z(n49183) );
  IV U59366 ( .A(n46491), .Z(n46492) );
  NOR U59367 ( .A(n46492), .B(n46497), .Z(n49181) );
  NOR U59368 ( .A(n49183), .B(n49181), .Z(n46493) );
  XOR U59369 ( .A(n49185), .B(n46493), .Z(n49179) );
  IV U59370 ( .A(n46494), .Z(n46496) );
  NOR U59371 ( .A(n46496), .B(n46495), .Z(n52979) );
  NOR U59372 ( .A(n46498), .B(n46497), .Z(n46499) );
  IV U59373 ( .A(n46499), .Z(n46501) );
  NOR U59374 ( .A(n46501), .B(n46500), .Z(n46502) );
  IV U59375 ( .A(n46502), .Z(n46507) );
  NOR U59376 ( .A(n46504), .B(n46503), .Z(n46505) );
  IV U59377 ( .A(n46505), .Z(n46506) );
  NOR U59378 ( .A(n46507), .B(n46506), .Z(n53693) );
  NOR U59379 ( .A(n52979), .B(n53693), .Z(n49180) );
  XOR U59380 ( .A(n49179), .B(n49180), .Z(n52973) );
  XOR U59381 ( .A(n49907), .B(n52973), .Z(n49176) );
  IV U59382 ( .A(n46508), .Z(n46509) );
  NOR U59383 ( .A(n46510), .B(n46509), .Z(n49177) );
  IV U59384 ( .A(n46511), .Z(n46513) );
  NOR U59385 ( .A(n46513), .B(n46512), .Z(n49908) );
  NOR U59386 ( .A(n49177), .B(n49908), .Z(n46514) );
  XOR U59387 ( .A(n49176), .B(n46514), .Z(n49172) );
  IV U59388 ( .A(n46515), .Z(n46517) );
  NOR U59389 ( .A(n46517), .B(n46516), .Z(n49170) );
  XOR U59390 ( .A(n49172), .B(n49170), .Z(n49175) );
  XOR U59391 ( .A(n49173), .B(n49175), .Z(n49168) );
  XOR U59392 ( .A(n46518), .B(n49168), .Z(n49152) );
  XOR U59393 ( .A(n46519), .B(n49152), .Z(n49160) );
  NOR U59394 ( .A(n46527), .B(n49160), .Z(n53703) );
  IV U59395 ( .A(n46520), .Z(n46522) );
  NOR U59396 ( .A(n46522), .B(n46521), .Z(n46523) );
  IV U59397 ( .A(n46523), .Z(n49151) );
  IV U59398 ( .A(n46524), .Z(n46526) );
  NOR U59399 ( .A(n46526), .B(n46525), .Z(n49159) );
  XOR U59400 ( .A(n49159), .B(n49160), .Z(n49150) );
  XOR U59401 ( .A(n49151), .B(n49150), .Z(n46530) );
  IV U59402 ( .A(n49150), .Z(n46528) );
  NOR U59403 ( .A(n46528), .B(n46527), .Z(n46529) );
  NOR U59404 ( .A(n46530), .B(n46529), .Z(n46531) );
  NOR U59405 ( .A(n53703), .B(n46531), .Z(n46532) );
  IV U59406 ( .A(n46532), .Z(n49143) );
  XOR U59407 ( .A(n49142), .B(n49143), .Z(n49147) );
  IV U59408 ( .A(n46533), .Z(n46534) );
  NOR U59409 ( .A(n46535), .B(n46534), .Z(n49145) );
  XOR U59410 ( .A(n49147), .B(n49145), .Z(n52939) );
  IV U59411 ( .A(n52939), .Z(n46545) );
  IV U59412 ( .A(n46536), .Z(n46537) );
  NOR U59413 ( .A(n46538), .B(n46537), .Z(n52942) );
  IV U59414 ( .A(n46539), .Z(n46544) );
  NOR U59415 ( .A(n46541), .B(n46540), .Z(n46542) );
  IV U59416 ( .A(n46542), .Z(n46543) );
  NOR U59417 ( .A(n46544), .B(n46543), .Z(n52937) );
  NOR U59418 ( .A(n52942), .B(n52937), .Z(n49921) );
  XOR U59419 ( .A(n46545), .B(n49921), .Z(n49139) );
  XOR U59420 ( .A(n49138), .B(n49139), .Z(n49918) );
  XOR U59421 ( .A(n49919), .B(n49918), .Z(n46552) );
  IV U59422 ( .A(n46552), .Z(n46546) );
  NOR U59423 ( .A(n46547), .B(n46546), .Z(n52928) );
  IV U59424 ( .A(n46548), .Z(n46549) );
  NOR U59425 ( .A(n46550), .B(n46549), .Z(n46553) );
  IV U59426 ( .A(n46553), .Z(n46551) );
  NOR U59427 ( .A(n46551), .B(n49918), .Z(n52932) );
  NOR U59428 ( .A(n46553), .B(n46552), .Z(n46554) );
  NOR U59429 ( .A(n52932), .B(n46554), .Z(n46555) );
  NOR U59430 ( .A(n46556), .B(n46555), .Z(n46557) );
  NOR U59431 ( .A(n52928), .B(n46557), .Z(n46558) );
  IV U59432 ( .A(n46558), .Z(n49136) );
  XOR U59433 ( .A(n49135), .B(n49136), .Z(n49130) );
  IV U59434 ( .A(n46559), .Z(n49132) );
  NOR U59435 ( .A(n49134), .B(n49132), .Z(n46563) );
  IV U59436 ( .A(n46560), .Z(n46562) );
  NOR U59437 ( .A(n46562), .B(n46561), .Z(n49129) );
  NOR U59438 ( .A(n46563), .B(n49129), .Z(n46564) );
  XOR U59439 ( .A(n49130), .B(n46564), .Z(n49126) );
  IV U59440 ( .A(n46565), .Z(n46566) );
  NOR U59441 ( .A(n46567), .B(n46566), .Z(n49127) );
  IV U59442 ( .A(n46568), .Z(n46569) );
  NOR U59443 ( .A(n46572), .B(n46569), .Z(n49946) );
  NOR U59444 ( .A(n49127), .B(n49946), .Z(n46570) );
  XOR U59445 ( .A(n49126), .B(n46570), .Z(n49124) );
  IV U59446 ( .A(n46571), .Z(n46573) );
  NOR U59447 ( .A(n46573), .B(n46572), .Z(n49122) );
  XOR U59448 ( .A(n49124), .B(n49122), .Z(n49933) );
  IV U59449 ( .A(n46574), .Z(n46575) );
  NOR U59450 ( .A(n49934), .B(n46575), .Z(n46576) );
  XOR U59451 ( .A(n49933), .B(n46576), .Z(n49117) );
  XOR U59452 ( .A(n49116), .B(n49117), .Z(n49120) );
  IV U59453 ( .A(n49120), .Z(n46583) );
  IV U59454 ( .A(n46577), .Z(n46578) );
  NOR U59455 ( .A(n46579), .B(n46578), .Z(n49119) );
  NOR U59456 ( .A(n46581), .B(n46580), .Z(n49114) );
  NOR U59457 ( .A(n49119), .B(n49114), .Z(n46582) );
  XOR U59458 ( .A(n46583), .B(n46582), .Z(n49958) );
  XOR U59459 ( .A(n49956), .B(n49958), .Z(n49960) );
  XOR U59460 ( .A(n49959), .B(n49960), .Z(n49099) );
  XOR U59461 ( .A(n46584), .B(n49099), .Z(n49094) );
  IV U59462 ( .A(n46585), .Z(n46587) );
  NOR U59463 ( .A(n46587), .B(n46586), .Z(n46590) );
  IV U59464 ( .A(n46588), .Z(n46589) );
  NOR U59465 ( .A(n46593), .B(n46589), .Z(n49093) );
  NOR U59466 ( .A(n46590), .B(n49093), .Z(n46591) );
  XOR U59467 ( .A(n49094), .B(n46591), .Z(n49968) );
  IV U59468 ( .A(n46592), .Z(n46594) );
  NOR U59469 ( .A(n46594), .B(n46593), .Z(n49966) );
  XOR U59470 ( .A(n49968), .B(n49966), .Z(n49971) );
  XOR U59471 ( .A(n49969), .B(n49971), .Z(n49978) );
  XOR U59472 ( .A(n49977), .B(n49978), .Z(n49981) );
  NOR U59473 ( .A(n46602), .B(n49981), .Z(n49986) );
  IV U59474 ( .A(n46595), .Z(n46596) );
  NOR U59475 ( .A(n46597), .B(n46596), .Z(n46598) );
  IV U59476 ( .A(n46598), .Z(n49975) );
  IV U59477 ( .A(n46599), .Z(n46601) );
  NOR U59478 ( .A(n46601), .B(n46600), .Z(n49980) );
  XOR U59479 ( .A(n49980), .B(n49981), .Z(n49974) );
  XOR U59480 ( .A(n49975), .B(n49974), .Z(n46605) );
  IV U59481 ( .A(n49974), .Z(n46603) );
  NOR U59482 ( .A(n46603), .B(n46602), .Z(n46604) );
  NOR U59483 ( .A(n46605), .B(n46604), .Z(n46606) );
  NOR U59484 ( .A(n49986), .B(n46606), .Z(n49091) );
  XOR U59485 ( .A(n46607), .B(n49091), .Z(n50001) );
  XOR U59486 ( .A(n49999), .B(n50001), .Z(n49993) );
  IV U59487 ( .A(n49993), .Z(n46614) );
  IV U59488 ( .A(n46608), .Z(n49087) );
  NOR U59489 ( .A(n46609), .B(n49087), .Z(n46612) );
  IV U59490 ( .A(n46610), .Z(n46611) );
  NOR U59491 ( .A(n46616), .B(n46611), .Z(n49991) );
  NOR U59492 ( .A(n46612), .B(n49991), .Z(n46613) );
  XOR U59493 ( .A(n46614), .B(n46613), .Z(n49083) );
  IV U59494 ( .A(n46615), .Z(n46617) );
  NOR U59495 ( .A(n46617), .B(n46616), .Z(n49081) );
  XOR U59496 ( .A(n49083), .B(n49081), .Z(n49084) );
  XOR U59497 ( .A(n49085), .B(n49084), .Z(n46624) );
  IV U59498 ( .A(n46624), .Z(n46618) );
  NOR U59499 ( .A(n46619), .B(n46618), .Z(n52866) );
  IV U59500 ( .A(n46620), .Z(n46622) );
  NOR U59501 ( .A(n46622), .B(n46621), .Z(n46625) );
  IV U59502 ( .A(n46625), .Z(n46623) );
  NOR U59503 ( .A(n46623), .B(n49084), .Z(n52862) );
  NOR U59504 ( .A(n46625), .B(n46624), .Z(n46626) );
  NOR U59505 ( .A(n52862), .B(n46626), .Z(n46627) );
  NOR U59506 ( .A(n46628), .B(n46627), .Z(n46629) );
  NOR U59507 ( .A(n52866), .B(n46629), .Z(n46630) );
  IV U59508 ( .A(n46630), .Z(n50010) );
  NOR U59509 ( .A(n46632), .B(n46631), .Z(n50009) );
  XOR U59510 ( .A(n50010), .B(n50009), .Z(n49079) );
  XOR U59511 ( .A(n49080), .B(n49079), .Z(n50024) );
  XOR U59512 ( .A(n50022), .B(n50024), .Z(n50014) );
  XOR U59513 ( .A(n46633), .B(n50014), .Z(n50030) );
  XOR U59514 ( .A(n50031), .B(n50030), .Z(n50033) );
  XOR U59515 ( .A(n46634), .B(n50033), .Z(n46635) );
  IV U59516 ( .A(n46635), .Z(n50040) );
  IV U59517 ( .A(n46636), .Z(n46637) );
  NOR U59518 ( .A(n46638), .B(n46637), .Z(n50038) );
  XOR U59519 ( .A(n50040), .B(n50038), .Z(n50048) );
  IV U59520 ( .A(n50048), .Z(n46646) );
  IV U59521 ( .A(n46639), .Z(n46640) );
  NOR U59522 ( .A(n46641), .B(n46640), .Z(n50041) );
  IV U59523 ( .A(n46642), .Z(n46644) );
  NOR U59524 ( .A(n46644), .B(n46643), .Z(n50047) );
  NOR U59525 ( .A(n50041), .B(n50047), .Z(n46645) );
  XOR U59526 ( .A(n46646), .B(n46645), .Z(n50045) );
  XOR U59527 ( .A(n50044), .B(n50045), .Z(n46659) );
  IV U59528 ( .A(n46659), .Z(n46650) );
  IV U59529 ( .A(n46647), .Z(n46648) );
  NOR U59530 ( .A(n46648), .B(n46652), .Z(n46664) );
  IV U59531 ( .A(n46664), .Z(n46649) );
  NOR U59532 ( .A(n46650), .B(n46649), .Z(n52827) );
  IV U59533 ( .A(n46651), .Z(n46653) );
  NOR U59534 ( .A(n46653), .B(n46652), .Z(n46654) );
  IV U59535 ( .A(n46654), .Z(n50055) );
  IV U59536 ( .A(n46655), .Z(n46657) );
  NOR U59537 ( .A(n46657), .B(n46656), .Z(n46660) );
  IV U59538 ( .A(n46660), .Z(n46658) );
  NOR U59539 ( .A(n50045), .B(n46658), .Z(n49074) );
  NOR U59540 ( .A(n46660), .B(n46659), .Z(n46661) );
  NOR U59541 ( .A(n49074), .B(n46661), .Z(n46662) );
  IV U59542 ( .A(n46662), .Z(n50054) );
  XOR U59543 ( .A(n50055), .B(n50054), .Z(n46663) );
  NOR U59544 ( .A(n46664), .B(n46663), .Z(n46665) );
  NOR U59545 ( .A(n52827), .B(n46665), .Z(n50064) );
  IV U59546 ( .A(n46666), .Z(n46667) );
  NOR U59547 ( .A(n46668), .B(n46667), .Z(n50067) );
  IV U59548 ( .A(n46669), .Z(n46671) );
  NOR U59549 ( .A(n46671), .B(n46670), .Z(n50065) );
  NOR U59550 ( .A(n50067), .B(n50065), .Z(n46672) );
  XOR U59551 ( .A(n50064), .B(n46672), .Z(n50059) );
  XOR U59552 ( .A(n50057), .B(n50059), .Z(n50077) );
  XOR U59553 ( .A(n50061), .B(n50077), .Z(n49059) );
  XOR U59554 ( .A(n46673), .B(n49059), .Z(n46674) );
  IV U59555 ( .A(n46674), .Z(n49054) );
  XOR U59556 ( .A(n46675), .B(n49054), .Z(n49051) );
  XOR U59557 ( .A(n46676), .B(n49051), .Z(n46677) );
  IV U59558 ( .A(n46677), .Z(n49041) );
  NOR U59559 ( .A(n46678), .B(n49041), .Z(n53815) );
  XOR U59560 ( .A(n49040), .B(n49041), .Z(n49037) );
  IV U59561 ( .A(n49037), .Z(n46679) );
  NOR U59562 ( .A(n46680), .B(n46679), .Z(n46681) );
  NOR U59563 ( .A(n53815), .B(n46681), .Z(n49032) );
  XOR U59564 ( .A(n46682), .B(n49032), .Z(n49031) );
  XOR U59565 ( .A(n49029), .B(n49031), .Z(n49027) );
  IV U59566 ( .A(n46683), .Z(n46684) );
  NOR U59567 ( .A(n46685), .B(n46684), .Z(n49023) );
  IV U59568 ( .A(n46686), .Z(n46687) );
  NOR U59569 ( .A(n46688), .B(n46687), .Z(n49025) );
  NOR U59570 ( .A(n49023), .B(n49025), .Z(n46689) );
  XOR U59571 ( .A(n49027), .B(n46689), .Z(n50092) );
  IV U59572 ( .A(n50092), .Z(n50095) );
  XOR U59573 ( .A(n46690), .B(n50095), .Z(n49021) );
  XOR U59574 ( .A(n46691), .B(n49021), .Z(n46692) );
  IV U59575 ( .A(n46692), .Z(n49015) );
  XOR U59576 ( .A(n49013), .B(n49015), .Z(n50112) );
  IV U59577 ( .A(n50112), .Z(n46700) );
  IV U59578 ( .A(n46693), .Z(n46695) );
  NOR U59579 ( .A(n46695), .B(n46694), .Z(n50111) );
  IV U59580 ( .A(n46696), .Z(n46698) );
  NOR U59581 ( .A(n46698), .B(n46697), .Z(n49016) );
  NOR U59582 ( .A(n50111), .B(n49016), .Z(n46699) );
  XOR U59583 ( .A(n46700), .B(n46699), .Z(n50123) );
  IV U59584 ( .A(n46701), .Z(n46703) );
  NOR U59585 ( .A(n46703), .B(n46702), .Z(n50121) );
  XOR U59586 ( .A(n50123), .B(n50121), .Z(n50118) );
  XOR U59587 ( .A(n50117), .B(n50118), .Z(n49011) );
  XOR U59588 ( .A(n49010), .B(n49011), .Z(n50139) );
  XOR U59589 ( .A(n46704), .B(n50139), .Z(n46705) );
  IV U59590 ( .A(n46705), .Z(n50143) );
  XOR U59591 ( .A(n50135), .B(n50143), .Z(n49008) );
  XOR U59592 ( .A(n46706), .B(n49008), .Z(n46715) );
  IV U59593 ( .A(n46715), .Z(n46710) );
  NOR U59594 ( .A(n46708), .B(n46707), .Z(n46718) );
  IV U59595 ( .A(n46718), .Z(n46709) );
  NOR U59596 ( .A(n46710), .B(n46709), .Z(n52778) );
  IV U59597 ( .A(n46711), .Z(n46712) );
  NOR U59598 ( .A(n46713), .B(n46712), .Z(n46716) );
  IV U59599 ( .A(n46716), .Z(n46714) );
  NOR U59600 ( .A(n46714), .B(n49008), .Z(n52781) );
  NOR U59601 ( .A(n46716), .B(n46715), .Z(n46717) );
  NOR U59602 ( .A(n52781), .B(n46717), .Z(n49004) );
  NOR U59603 ( .A(n46718), .B(n49004), .Z(n46719) );
  NOR U59604 ( .A(n52778), .B(n46719), .Z(n46720) );
  IV U59605 ( .A(n46720), .Z(n46721) );
  NOR U59606 ( .A(n46722), .B(n46721), .Z(n49001) );
  IV U59607 ( .A(n46722), .Z(n49006) );
  NOR U59608 ( .A(n49004), .B(n49006), .Z(n46723) );
  NOR U59609 ( .A(n49001), .B(n46723), .Z(n48999) );
  IV U59610 ( .A(n46724), .Z(n46725) );
  NOR U59611 ( .A(n46726), .B(n46725), .Z(n49000) );
  IV U59612 ( .A(n46727), .Z(n46729) );
  NOR U59613 ( .A(n46729), .B(n46728), .Z(n48997) );
  NOR U59614 ( .A(n49000), .B(n48997), .Z(n46730) );
  XOR U59615 ( .A(n48999), .B(n46730), .Z(n48994) );
  IV U59616 ( .A(n46731), .Z(n46733) );
  NOR U59617 ( .A(n46733), .B(n46732), .Z(n46738) );
  IV U59618 ( .A(n46734), .Z(n46735) );
  NOR U59619 ( .A(n46736), .B(n46735), .Z(n46737) );
  NOR U59620 ( .A(n46738), .B(n46737), .Z(n48996) );
  XOR U59621 ( .A(n48994), .B(n48996), .Z(n48992) );
  XOR U59622 ( .A(n46739), .B(n48992), .Z(n46740) );
  IV U59623 ( .A(n46740), .Z(n50149) );
  XOR U59624 ( .A(n50148), .B(n50149), .Z(n53856) );
  IV U59625 ( .A(n46741), .Z(n46742) );
  NOR U59626 ( .A(n46743), .B(n46742), .Z(n53854) );
  IV U59627 ( .A(n46744), .Z(n46745) );
  NOR U59628 ( .A(n46746), .B(n46745), .Z(n53863) );
  NOR U59629 ( .A(n53854), .B(n53863), .Z(n50151) );
  XOR U59630 ( .A(n53856), .B(n50151), .Z(n48986) );
  XOR U59631 ( .A(n46747), .B(n48986), .Z(n48984) );
  IV U59632 ( .A(n46748), .Z(n46750) );
  NOR U59633 ( .A(n46750), .B(n46749), .Z(n46751) );
  IV U59634 ( .A(n46751), .Z(n48983) );
  XOR U59635 ( .A(n48984), .B(n48983), .Z(n48980) );
  IV U59636 ( .A(n46752), .Z(n46753) );
  NOR U59637 ( .A(n46754), .B(n46753), .Z(n50158) );
  IV U59638 ( .A(n46755), .Z(n46756) );
  NOR U59639 ( .A(n46756), .B(n46760), .Z(n48981) );
  NOR U59640 ( .A(n50158), .B(n48981), .Z(n46757) );
  XOR U59641 ( .A(n48980), .B(n46757), .Z(n50169) );
  IV U59642 ( .A(n46758), .Z(n46759) );
  NOR U59643 ( .A(n46760), .B(n46759), .Z(n50167) );
  XOR U59644 ( .A(n50169), .B(n50167), .Z(n50171) );
  NOR U59645 ( .A(n46761), .B(n50171), .Z(n52745) );
  IV U59646 ( .A(n46762), .Z(n46763) );
  NOR U59647 ( .A(n46764), .B(n46763), .Z(n50170) );
  XOR U59648 ( .A(n50170), .B(n50171), .Z(n48978) );
  IV U59649 ( .A(n48978), .Z(n46765) );
  NOR U59650 ( .A(n46766), .B(n46765), .Z(n46767) );
  NOR U59651 ( .A(n52745), .B(n46767), .Z(n50175) );
  IV U59652 ( .A(n46768), .Z(n46769) );
  NOR U59653 ( .A(n46770), .B(n46769), .Z(n48977) );
  IV U59654 ( .A(n46771), .Z(n46773) );
  NOR U59655 ( .A(n46773), .B(n46772), .Z(n50176) );
  NOR U59656 ( .A(n48977), .B(n50176), .Z(n46774) );
  XOR U59657 ( .A(n50175), .B(n46774), .Z(n50188) );
  XOR U59658 ( .A(n50186), .B(n50188), .Z(n50197) );
  XOR U59659 ( .A(n46775), .B(n50197), .Z(n46776) );
  IV U59660 ( .A(n46776), .Z(n50211) );
  XOR U59661 ( .A(n50212), .B(n50211), .Z(n46777) );
  XOR U59662 ( .A(n46778), .B(n46777), .Z(n50217) );
  IV U59663 ( .A(n46779), .Z(n46781) );
  NOR U59664 ( .A(n46781), .B(n46780), .Z(n50215) );
  NOR U59665 ( .A(n50215), .B(n50213), .Z(n46782) );
  XOR U59666 ( .A(n50217), .B(n46782), .Z(n48975) );
  NOR U59667 ( .A(n46784), .B(n46783), .Z(n48969) );
  IV U59668 ( .A(n46785), .Z(n46787) );
  IV U59669 ( .A(n46786), .Z(n46789) );
  NOR U59670 ( .A(n46787), .B(n46789), .Z(n52723) );
  IV U59671 ( .A(n46788), .Z(n46790) );
  NOR U59672 ( .A(n46790), .B(n46789), .Z(n52728) );
  NOR U59673 ( .A(n52723), .B(n52728), .Z(n48976) );
  IV U59674 ( .A(n48976), .Z(n46791) );
  NOR U59675 ( .A(n48969), .B(n46791), .Z(n46792) );
  XOR U59676 ( .A(n48975), .B(n46792), .Z(n50225) );
  NOR U59677 ( .A(n46798), .B(n50225), .Z(n48967) );
  IV U59678 ( .A(n46793), .Z(n46795) );
  NOR U59679 ( .A(n46795), .B(n46794), .Z(n46796) );
  IV U59680 ( .A(n46796), .Z(n50231) );
  NOR U59681 ( .A(n46797), .B(n48971), .Z(n50224) );
  XOR U59682 ( .A(n50224), .B(n50225), .Z(n50230) );
  XOR U59683 ( .A(n50231), .B(n50230), .Z(n46801) );
  IV U59684 ( .A(n50230), .Z(n46799) );
  NOR U59685 ( .A(n46799), .B(n46798), .Z(n46800) );
  NOR U59686 ( .A(n46801), .B(n46800), .Z(n46802) );
  NOR U59687 ( .A(n48967), .B(n46802), .Z(n50233) );
  IV U59688 ( .A(n46803), .Z(n46804) );
  NOR U59689 ( .A(n46805), .B(n46804), .Z(n50232) );
  IV U59690 ( .A(n46806), .Z(n46807) );
  NOR U59691 ( .A(n46808), .B(n46807), .Z(n50237) );
  NOR U59692 ( .A(n50232), .B(n50237), .Z(n46809) );
  XOR U59693 ( .A(n50233), .B(n46809), .Z(n46825) );
  NOR U59694 ( .A(n46825), .B(n46812), .Z(n46810) );
  IV U59695 ( .A(n46810), .Z(n46819) );
  NOR U59696 ( .A(n46811), .B(n46819), .Z(n50236) );
  NOR U59697 ( .A(n46813), .B(n46812), .Z(n46817) );
  IV U59698 ( .A(n46814), .Z(n46816) );
  NOR U59699 ( .A(n46816), .B(n46815), .Z(n46821) );
  NOR U59700 ( .A(n46817), .B(n46821), .Z(n46824) );
  IV U59701 ( .A(n46818), .Z(n46820) );
  NOR U59702 ( .A(n46820), .B(n46819), .Z(n52707) );
  IV U59703 ( .A(n46821), .Z(n46822) );
  NOR U59704 ( .A(n46825), .B(n46822), .Z(n53914) );
  NOR U59705 ( .A(n52707), .B(n53914), .Z(n46823) );
  IV U59706 ( .A(n46823), .Z(n50248) );
  NOR U59707 ( .A(n46824), .B(n50248), .Z(n46827) );
  NOR U59708 ( .A(n46825), .B(n50248), .Z(n46826) );
  NOR U59709 ( .A(n46827), .B(n46826), .Z(n46828) );
  NOR U59710 ( .A(n50236), .B(n46828), .Z(n46834) );
  XOR U59711 ( .A(n50245), .B(n46834), .Z(n46840) );
  IV U59712 ( .A(n46840), .Z(n46833) );
  IV U59713 ( .A(n46829), .Z(n46831) );
  NOR U59714 ( .A(n46831), .B(n46830), .Z(n46843) );
  IV U59715 ( .A(n46843), .Z(n46832) );
  NOR U59716 ( .A(n46833), .B(n46832), .Z(n52702) );
  IV U59717 ( .A(n46834), .Z(n50246) );
  IV U59718 ( .A(n46835), .Z(n46837) );
  NOR U59719 ( .A(n46837), .B(n46836), .Z(n46839) );
  IV U59720 ( .A(n46839), .Z(n46838) );
  NOR U59721 ( .A(n50246), .B(n46838), .Z(n52701) );
  NOR U59722 ( .A(n46840), .B(n46839), .Z(n46841) );
  NOR U59723 ( .A(n52701), .B(n46841), .Z(n46842) );
  NOR U59724 ( .A(n46843), .B(n46842), .Z(n46844) );
  NOR U59725 ( .A(n52702), .B(n46844), .Z(n48961) );
  IV U59726 ( .A(n46845), .Z(n46850) );
  IV U59727 ( .A(n46846), .Z(n46847) );
  NOR U59728 ( .A(n46850), .B(n46847), .Z(n48960) );
  IV U59729 ( .A(n46848), .Z(n46849) );
  NOR U59730 ( .A(n46850), .B(n46849), .Z(n48957) );
  NOR U59731 ( .A(n48960), .B(n48957), .Z(n46851) );
  XOR U59732 ( .A(n48961), .B(n46851), .Z(n48954) );
  XOR U59733 ( .A(n46852), .B(n48954), .Z(n48944) );
  XOR U59734 ( .A(n48945), .B(n48944), .Z(n48947) );
  NOR U59735 ( .A(n46858), .B(n48947), .Z(n53926) );
  NOR U59736 ( .A(n46854), .B(n46853), .Z(n46855) );
  IV U59737 ( .A(n46855), .Z(n50258) );
  NOR U59738 ( .A(n46857), .B(n46856), .Z(n48939) );
  XOR U59739 ( .A(n48939), .B(n48947), .Z(n50257) );
  XOR U59740 ( .A(n50258), .B(n50257), .Z(n46861) );
  IV U59741 ( .A(n50257), .Z(n46859) );
  NOR U59742 ( .A(n46859), .B(n46858), .Z(n46860) );
  NOR U59743 ( .A(n46861), .B(n46860), .Z(n46862) );
  NOR U59744 ( .A(n53926), .B(n46862), .Z(n46863) );
  IV U59745 ( .A(n46863), .Z(n50260) );
  XOR U59746 ( .A(n50259), .B(n50260), .Z(n50265) );
  IV U59747 ( .A(n46864), .Z(n46866) );
  NOR U59748 ( .A(n46866), .B(n46865), .Z(n48936) );
  NOR U59749 ( .A(n50264), .B(n48936), .Z(n46867) );
  XOR U59750 ( .A(n50265), .B(n46867), .Z(n46868) );
  IV U59751 ( .A(n46868), .Z(n48932) );
  XOR U59752 ( .A(n48930), .B(n48932), .Z(n48934) );
  NOR U59753 ( .A(n46876), .B(n48934), .Z(n53950) );
  IV U59754 ( .A(n46869), .Z(n46871) );
  NOR U59755 ( .A(n46871), .B(n46870), .Z(n46872) );
  IV U59756 ( .A(n46872), .Z(n48928) );
  IV U59757 ( .A(n46873), .Z(n46874) );
  NOR U59758 ( .A(n46875), .B(n46874), .Z(n48933) );
  XOR U59759 ( .A(n48933), .B(n48934), .Z(n48927) );
  XOR U59760 ( .A(n48928), .B(n48927), .Z(n46879) );
  IV U59761 ( .A(n48927), .Z(n46877) );
  NOR U59762 ( .A(n46877), .B(n46876), .Z(n46878) );
  NOR U59763 ( .A(n46879), .B(n46878), .Z(n46880) );
  NOR U59764 ( .A(n53950), .B(n46880), .Z(n46881) );
  IV U59765 ( .A(n46881), .Z(n50276) );
  XOR U59766 ( .A(n50269), .B(n50276), .Z(n50272) );
  XOR U59767 ( .A(n46882), .B(n50272), .Z(n50280) );
  XOR U59768 ( .A(n46883), .B(n50280), .Z(n48923) );
  XOR U59769 ( .A(n48924), .B(n48923), .Z(n53959) );
  XOR U59770 ( .A(n50294), .B(n53959), .Z(n48919) );
  IV U59771 ( .A(n46884), .Z(n46886) );
  NOR U59772 ( .A(n46886), .B(n46885), .Z(n50295) );
  IV U59773 ( .A(n46887), .Z(n46888) );
  NOR U59774 ( .A(n46888), .B(n46891), .Z(n48921) );
  NOR U59775 ( .A(n50295), .B(n48921), .Z(n46889) );
  XOR U59776 ( .A(n48919), .B(n46889), .Z(n50310) );
  IV U59777 ( .A(n46890), .Z(n46892) );
  NOR U59778 ( .A(n46892), .B(n46891), .Z(n48918) );
  IV U59779 ( .A(n46893), .Z(n46895) );
  NOR U59780 ( .A(n46895), .B(n46894), .Z(n50309) );
  NOR U59781 ( .A(n48918), .B(n50309), .Z(n46896) );
  XOR U59782 ( .A(n50310), .B(n46896), .Z(n50314) );
  XOR U59783 ( .A(n46897), .B(n50314), .Z(n50323) );
  XOR U59784 ( .A(n50321), .B(n50323), .Z(n50331) );
  XOR U59785 ( .A(n46898), .B(n50331), .Z(n46899) );
  IV U59786 ( .A(n46899), .Z(n50336) );
  IV U59787 ( .A(n46900), .Z(n46902) );
  NOR U59788 ( .A(n46902), .B(n46901), .Z(n46903) );
  IV U59789 ( .A(n46903), .Z(n50333) );
  XOR U59790 ( .A(n50336), .B(n50333), .Z(n46904) );
  XOR U59791 ( .A(n46905), .B(n46904), .Z(n48909) );
  IV U59792 ( .A(n48909), .Z(n48906) );
  XOR U59793 ( .A(n48908), .B(n48906), .Z(n46906) );
  NOR U59794 ( .A(n46911), .B(n46906), .Z(n52622) );
  XOR U59795 ( .A(n46907), .B(n46906), .Z(n48903) );
  IV U59796 ( .A(n46908), .Z(n46910) );
  NOR U59797 ( .A(n46910), .B(n46909), .Z(n46912) );
  IV U59798 ( .A(n46912), .Z(n48902) );
  XOR U59799 ( .A(n48903), .B(n48902), .Z(n46914) );
  NOR U59800 ( .A(n46912), .B(n46911), .Z(n46913) );
  NOR U59801 ( .A(n46914), .B(n46913), .Z(n46915) );
  NOR U59802 ( .A(n52622), .B(n46915), .Z(n50338) );
  XOR U59803 ( .A(n50339), .B(n50338), .Z(n50348) );
  XOR U59804 ( .A(n46916), .B(n50348), .Z(n46917) );
  NOR U59805 ( .A(n46918), .B(n46917), .Z(n54000) );
  IV U59806 ( .A(n46917), .Z(n46920) );
  IV U59807 ( .A(n46918), .Z(n46919) );
  NOR U59808 ( .A(n46920), .B(n46919), .Z(n53997) );
  NOR U59809 ( .A(n54000), .B(n53997), .Z(n50353) );
  XOR U59810 ( .A(n50354), .B(n50353), .Z(n48901) );
  NOR U59811 ( .A(n46924), .B(n48901), .Z(n48899) );
  IV U59812 ( .A(n46921), .Z(n46923) );
  NOR U59813 ( .A(n46923), .B(n46922), .Z(n46925) );
  IV U59814 ( .A(n46925), .Z(n48900) );
  XOR U59815 ( .A(n48901), .B(n48900), .Z(n46927) );
  NOR U59816 ( .A(n46925), .B(n46924), .Z(n46926) );
  NOR U59817 ( .A(n46927), .B(n46926), .Z(n48896) );
  NOR U59818 ( .A(n48899), .B(n48896), .Z(n46928) );
  IV U59819 ( .A(n46928), .Z(n50359) );
  IV U59820 ( .A(n46929), .Z(n46931) );
  NOR U59821 ( .A(n46931), .B(n46930), .Z(n48895) );
  IV U59822 ( .A(n46932), .Z(n46933) );
  NOR U59823 ( .A(n46933), .B(n48884), .Z(n50358) );
  NOR U59824 ( .A(n48895), .B(n50358), .Z(n46934) );
  XOR U59825 ( .A(n50359), .B(n46934), .Z(n48883) );
  NOR U59826 ( .A(n46936), .B(n46935), .Z(n50362) );
  NOR U59827 ( .A(n46937), .B(n50362), .Z(n46938) );
  XOR U59828 ( .A(n48883), .B(n46938), .Z(n50367) );
  XOR U59829 ( .A(n50366), .B(n50367), .Z(n50375) );
  IV U59830 ( .A(n50375), .Z(n46947) );
  NOR U59831 ( .A(n46940), .B(n46939), .Z(n50369) );
  IV U59832 ( .A(n46941), .Z(n46945) );
  NOR U59833 ( .A(n46943), .B(n46942), .Z(n46944) );
  IV U59834 ( .A(n46944), .Z(n46949) );
  NOR U59835 ( .A(n46945), .B(n46949), .Z(n50373) );
  NOR U59836 ( .A(n50369), .B(n50373), .Z(n46946) );
  XOR U59837 ( .A(n46947), .B(n46946), .Z(n50379) );
  IV U59838 ( .A(n46948), .Z(n46950) );
  NOR U59839 ( .A(n46950), .B(n46949), .Z(n50377) );
  XOR U59840 ( .A(n50379), .B(n50377), .Z(n48879) );
  XOR U59841 ( .A(n48878), .B(n48879), .Z(n50386) );
  XOR U59842 ( .A(n50385), .B(n50386), .Z(n52585) );
  XOR U59843 ( .A(n50388), .B(n52585), .Z(n50391) );
  IV U59844 ( .A(n46951), .Z(n46963) );
  IV U59845 ( .A(n46952), .Z(n46953) );
  NOR U59846 ( .A(n46963), .B(n46953), .Z(n50397) );
  IV U59847 ( .A(n46954), .Z(n46956) );
  NOR U59848 ( .A(n46956), .B(n46955), .Z(n50392) );
  NOR U59849 ( .A(n50397), .B(n50392), .Z(n46957) );
  XOR U59850 ( .A(n50391), .B(n46957), .Z(n50409) );
  IV U59851 ( .A(n46958), .Z(n46959) );
  NOR U59852 ( .A(n46960), .B(n46959), .Z(n50407) );
  IV U59853 ( .A(n46961), .Z(n46962) );
  NOR U59854 ( .A(n46963), .B(n46962), .Z(n48876) );
  NOR U59855 ( .A(n50407), .B(n48876), .Z(n46964) );
  XOR U59856 ( .A(n50409), .B(n46964), .Z(n48869) );
  IV U59857 ( .A(n46965), .Z(n46966) );
  NOR U59858 ( .A(n46967), .B(n46966), .Z(n48873) );
  NOR U59859 ( .A(n46968), .B(n48870), .Z(n46969) );
  NOR U59860 ( .A(n48873), .B(n46969), .Z(n46970) );
  XOR U59861 ( .A(n48869), .B(n46970), .Z(n48867) );
  XOR U59862 ( .A(n48866), .B(n48867), .Z(n46977) );
  IV U59863 ( .A(n46977), .Z(n46971) );
  NOR U59864 ( .A(n46972), .B(n46971), .Z(n52568) );
  IV U59865 ( .A(n46973), .Z(n46975) );
  NOR U59866 ( .A(n46975), .B(n46974), .Z(n46978) );
  IV U59867 ( .A(n46978), .Z(n46976) );
  NOR U59868 ( .A(n48867), .B(n46976), .Z(n52565) );
  NOR U59869 ( .A(n46978), .B(n46977), .Z(n46979) );
  NOR U59870 ( .A(n52565), .B(n46979), .Z(n46980) );
  NOR U59871 ( .A(n46981), .B(n46980), .Z(n46982) );
  NOR U59872 ( .A(n52568), .B(n46982), .Z(n48864) );
  IV U59873 ( .A(n46983), .Z(n46984) );
  NOR U59874 ( .A(n46985), .B(n46984), .Z(n50427) );
  IV U59875 ( .A(n46986), .Z(n46987) );
  NOR U59876 ( .A(n46988), .B(n46987), .Z(n50423) );
  NOR U59877 ( .A(n50427), .B(n50423), .Z(n48865) );
  XOR U59878 ( .A(n48864), .B(n48865), .Z(n48862) );
  XOR U59879 ( .A(n48863), .B(n48862), .Z(n48859) );
  NOR U59880 ( .A(n46989), .B(n46991), .Z(n50439) );
  IV U59881 ( .A(n46990), .Z(n46992) );
  NOR U59882 ( .A(n46992), .B(n46991), .Z(n48860) );
  NOR U59883 ( .A(n50439), .B(n48860), .Z(n46993) );
  XOR U59884 ( .A(n50437), .B(n46993), .Z(n46994) );
  XOR U59885 ( .A(n48859), .B(n46994), .Z(n50444) );
  XOR U59886 ( .A(n50442), .B(n50444), .Z(n50446) );
  IV U59887 ( .A(n46995), .Z(n46996) );
  NOR U59888 ( .A(n46997), .B(n46996), .Z(n50445) );
  NOR U59889 ( .A(n46998), .B(n48856), .Z(n46999) );
  NOR U59890 ( .A(n50445), .B(n46999), .Z(n47000) );
  XOR U59891 ( .A(n50446), .B(n47000), .Z(n47011) );
  IV U59892 ( .A(n47011), .Z(n47005) );
  IV U59893 ( .A(n47001), .Z(n47002) );
  NOR U59894 ( .A(n47003), .B(n47002), .Z(n47020) );
  IV U59895 ( .A(n47020), .Z(n47004) );
  NOR U59896 ( .A(n47005), .B(n47004), .Z(n54053) );
  XOR U59897 ( .A(n50445), .B(n50446), .Z(n47010) );
  IV U59898 ( .A(n47006), .Z(n47017) );
  IV U59899 ( .A(n47007), .Z(n47008) );
  NOR U59900 ( .A(n47017), .B(n47008), .Z(n47012) );
  IV U59901 ( .A(n47012), .Z(n47009) );
  NOR U59902 ( .A(n47010), .B(n47009), .Z(n52542) );
  NOR U59903 ( .A(n47012), .B(n47011), .Z(n47013) );
  NOR U59904 ( .A(n52542), .B(n47013), .Z(n47014) );
  IV U59905 ( .A(n47014), .Z(n48854) );
  IV U59906 ( .A(n47015), .Z(n47016) );
  NOR U59907 ( .A(n47017), .B(n47016), .Z(n47018) );
  IV U59908 ( .A(n47018), .Z(n48853) );
  XOR U59909 ( .A(n48854), .B(n48853), .Z(n47019) );
  NOR U59910 ( .A(n47020), .B(n47019), .Z(n47021) );
  NOR U59911 ( .A(n54053), .B(n47021), .Z(n47022) );
  IV U59912 ( .A(n47022), .Z(n48851) );
  IV U59913 ( .A(n47023), .Z(n47024) );
  NOR U59914 ( .A(n47025), .B(n47024), .Z(n48850) );
  XOR U59915 ( .A(n48851), .B(n48850), .Z(n48843) );
  XOR U59916 ( .A(n48841), .B(n48843), .Z(n48845) );
  XOR U59917 ( .A(n48844), .B(n48845), .Z(n48849) );
  XOR U59918 ( .A(n47026), .B(n48849), .Z(n47027) );
  IV U59919 ( .A(n47027), .Z(n50464) );
  XOR U59920 ( .A(n50463), .B(n50464), .Z(n50462) );
  IV U59921 ( .A(n47028), .Z(n47029) );
  NOR U59922 ( .A(n47030), .B(n47029), .Z(n48837) );
  IV U59923 ( .A(n47031), .Z(n47032) );
  NOR U59924 ( .A(n47033), .B(n47032), .Z(n50460) );
  NOR U59925 ( .A(n48837), .B(n50460), .Z(n47034) );
  XOR U59926 ( .A(n50462), .B(n47034), .Z(n48835) );
  XOR U59927 ( .A(n47035), .B(n48835), .Z(n48828) );
  XOR U59928 ( .A(n48826), .B(n48828), .Z(n48831) );
  IV U59929 ( .A(n47036), .Z(n47038) );
  NOR U59930 ( .A(n47038), .B(n47037), .Z(n48829) );
  XOR U59931 ( .A(n48831), .B(n48829), .Z(n48823) );
  IV U59932 ( .A(n47039), .Z(n47040) );
  NOR U59933 ( .A(n47043), .B(n47040), .Z(n48822) );
  IV U59934 ( .A(n47041), .Z(n47042) );
  NOR U59935 ( .A(n47043), .B(n47042), .Z(n48817) );
  NOR U59936 ( .A(n48822), .B(n48817), .Z(n47044) );
  XOR U59937 ( .A(n48823), .B(n47044), .Z(n48819) );
  XOR U59938 ( .A(n48820), .B(n48819), .Z(n48813) );
  IV U59939 ( .A(n47045), .Z(n47046) );
  NOR U59940 ( .A(n47047), .B(n47046), .Z(n48811) );
  XOR U59941 ( .A(n48813), .B(n48811), .Z(n48816) );
  IV U59942 ( .A(n47048), .Z(n47050) );
  NOR U59943 ( .A(n47050), .B(n47049), .Z(n48814) );
  XOR U59944 ( .A(n48816), .B(n48814), .Z(n48806) );
  XOR U59945 ( .A(n48805), .B(n48806), .Z(n48809) );
  IV U59946 ( .A(n47051), .Z(n47053) );
  NOR U59947 ( .A(n47053), .B(n47052), .Z(n48808) );
  IV U59948 ( .A(n47054), .Z(n47056) );
  NOR U59949 ( .A(n47056), .B(n47055), .Z(n48803) );
  NOR U59950 ( .A(n48808), .B(n48803), .Z(n47057) );
  XOR U59951 ( .A(n48809), .B(n47057), .Z(n48796) );
  XOR U59952 ( .A(n47058), .B(n48796), .Z(n48795) );
  XOR U59953 ( .A(n48793), .B(n48795), .Z(n50484) );
  IV U59954 ( .A(n50484), .Z(n50491) );
  IV U59955 ( .A(n47059), .Z(n47060) );
  NOR U59956 ( .A(n47061), .B(n47060), .Z(n50482) );
  NOR U59957 ( .A(n47062), .B(n50485), .Z(n47063) );
  NOR U59958 ( .A(n50482), .B(n47063), .Z(n47064) );
  XOR U59959 ( .A(n50491), .B(n47064), .Z(n48791) );
  XOR U59960 ( .A(n47065), .B(n48791), .Z(n50508) );
  IV U59961 ( .A(n50508), .Z(n52492) );
  XOR U59962 ( .A(n50509), .B(n52492), .Z(n52474) );
  XOR U59963 ( .A(n50514), .B(n52474), .Z(n50520) );
  XOR U59964 ( .A(n47066), .B(n50520), .Z(n47067) );
  IV U59965 ( .A(n47067), .Z(n50526) );
  XOR U59966 ( .A(n48788), .B(n50526), .Z(n48786) );
  IV U59967 ( .A(n48786), .Z(n47075) );
  IV U59968 ( .A(n47068), .Z(n47070) );
  NOR U59969 ( .A(n47070), .B(n47069), .Z(n50524) );
  IV U59970 ( .A(n47071), .Z(n47073) );
  NOR U59971 ( .A(n47073), .B(n47072), .Z(n48785) );
  NOR U59972 ( .A(n50524), .B(n48785), .Z(n47074) );
  XOR U59973 ( .A(n47075), .B(n47074), .Z(n50540) );
  XOR U59974 ( .A(n50538), .B(n50540), .Z(n50542) );
  XOR U59975 ( .A(n50541), .B(n50542), .Z(n50547) );
  XOR U59976 ( .A(n47076), .B(n50547), .Z(n48782) );
  XOR U59977 ( .A(n47077), .B(n48782), .Z(n50559) );
  XOR U59978 ( .A(n47078), .B(n50559), .Z(n48775) );
  IV U59979 ( .A(n47079), .Z(n47080) );
  NOR U59980 ( .A(n47081), .B(n47080), .Z(n48777) );
  IV U59981 ( .A(n47082), .Z(n47083) );
  NOR U59982 ( .A(n47084), .B(n47083), .Z(n48774) );
  NOR U59983 ( .A(n48777), .B(n48774), .Z(n47085) );
  XOR U59984 ( .A(n48775), .B(n47085), .Z(n50572) );
  IV U59985 ( .A(n47086), .Z(n47087) );
  NOR U59986 ( .A(n47088), .B(n47087), .Z(n50570) );
  XOR U59987 ( .A(n50572), .B(n50570), .Z(n50579) );
  XOR U59988 ( .A(n47089), .B(n50579), .Z(n48772) );
  IV U59989 ( .A(n47090), .Z(n47092) );
  NOR U59990 ( .A(n47092), .B(n47091), .Z(n48771) );
  IV U59991 ( .A(n47093), .Z(n47095) );
  NOR U59992 ( .A(n47095), .B(n47094), .Z(n50587) );
  NOR U59993 ( .A(n48771), .B(n50587), .Z(n47096) );
  XOR U59994 ( .A(n48772), .B(n47096), .Z(n50594) );
  XOR U59995 ( .A(n47097), .B(n50594), .Z(n48765) );
  XOR U59996 ( .A(n47098), .B(n48765), .Z(n48763) );
  XOR U59997 ( .A(n47099), .B(n48763), .Z(n48755) );
  IV U59998 ( .A(n47100), .Z(n47101) );
  NOR U59999 ( .A(n47102), .B(n47101), .Z(n47103) );
  IV U60000 ( .A(n47103), .Z(n48756) );
  IV U60001 ( .A(n47104), .Z(n47106) );
  NOR U60002 ( .A(n47106), .B(n47105), .Z(n47107) );
  IV U60003 ( .A(n47107), .Z(n48757) );
  XOR U60004 ( .A(n48756), .B(n48757), .Z(n47108) );
  XOR U60005 ( .A(n48755), .B(n47108), .Z(n48753) );
  IV U60006 ( .A(n47109), .Z(n47111) );
  NOR U60007 ( .A(n47111), .B(n47110), .Z(n54168) );
  IV U60008 ( .A(n47112), .Z(n47114) );
  NOR U60009 ( .A(n47114), .B(n47113), .Z(n52422) );
  NOR U60010 ( .A(n54168), .B(n52422), .Z(n48754) );
  XOR U60011 ( .A(n48753), .B(n48754), .Z(n50600) );
  XOR U60012 ( .A(n50598), .B(n50600), .Z(n48752) );
  XOR U60013 ( .A(n48750), .B(n48752), .Z(n50616) );
  NOR U60014 ( .A(n47122), .B(n50616), .Z(n50621) );
  IV U60015 ( .A(n47115), .Z(n47116) );
  NOR U60016 ( .A(n47117), .B(n47116), .Z(n50615) );
  NOR U60017 ( .A(n48748), .B(n50615), .Z(n47118) );
  XOR U60018 ( .A(n47118), .B(n50616), .Z(n47119) );
  IV U60019 ( .A(n47119), .Z(n48747) );
  IV U60020 ( .A(n47120), .Z(n47121) );
  NOR U60021 ( .A(n47129), .B(n47121), .Z(n47123) );
  IV U60022 ( .A(n47123), .Z(n48746) );
  XOR U60023 ( .A(n48747), .B(n48746), .Z(n47125) );
  NOR U60024 ( .A(n47123), .B(n47122), .Z(n47124) );
  NOR U60025 ( .A(n47125), .B(n47124), .Z(n47126) );
  NOR U60026 ( .A(n50621), .B(n47126), .Z(n47127) );
  IV U60027 ( .A(n47127), .Z(n50628) );
  IV U60028 ( .A(n47128), .Z(n47130) );
  NOR U60029 ( .A(n47130), .B(n47129), .Z(n50627) );
  XOR U60030 ( .A(n50628), .B(n50627), .Z(n50634) );
  XOR U60031 ( .A(n47131), .B(n50634), .Z(n48743) );
  XOR U60032 ( .A(n47132), .B(n48743), .Z(n50660) );
  XOR U60033 ( .A(n47133), .B(n50660), .Z(n48740) );
  XOR U60034 ( .A(n47134), .B(n48740), .Z(n48738) );
  NOR U60035 ( .A(n47135), .B(n48738), .Z(n54193) );
  IV U60036 ( .A(n47136), .Z(n47137) );
  NOR U60037 ( .A(n47138), .B(n47137), .Z(n48737) );
  XOR U60038 ( .A(n48737), .B(n48738), .Z(n48735) );
  IV U60039 ( .A(n48735), .Z(n47139) );
  NOR U60040 ( .A(n47140), .B(n47139), .Z(n47141) );
  NOR U60041 ( .A(n54193), .B(n47141), .Z(n48731) );
  IV U60042 ( .A(n47142), .Z(n47144) );
  NOR U60043 ( .A(n47144), .B(n47143), .Z(n48734) );
  IV U60044 ( .A(n47145), .Z(n47147) );
  NOR U60045 ( .A(n47147), .B(n47146), .Z(n48730) );
  NOR U60046 ( .A(n48734), .B(n48730), .Z(n47148) );
  XOR U60047 ( .A(n48731), .B(n47148), .Z(n52399) );
  XOR U60048 ( .A(n48729), .B(n52399), .Z(n47149) );
  IV U60049 ( .A(n47149), .Z(n50673) );
  XOR U60050 ( .A(n50672), .B(n50673), .Z(n50679) );
  IV U60051 ( .A(n50679), .Z(n47157) );
  IV U60052 ( .A(n47150), .Z(n47152) );
  NOR U60053 ( .A(n47152), .B(n47151), .Z(n50675) );
  IV U60054 ( .A(n47153), .Z(n47154) );
  NOR U60055 ( .A(n47155), .B(n47154), .Z(n50678) );
  NOR U60056 ( .A(n50675), .B(n50678), .Z(n47156) );
  XOR U60057 ( .A(n47157), .B(n47156), .Z(n52386) );
  NOR U60058 ( .A(n47158), .B(n52383), .Z(n48725) );
  IV U60059 ( .A(n47159), .Z(n47161) );
  NOR U60060 ( .A(n47161), .B(n47160), .Z(n48727) );
  NOR U60061 ( .A(n48725), .B(n48727), .Z(n47162) );
  XOR U60062 ( .A(n52386), .B(n47162), .Z(n47168) );
  IV U60063 ( .A(n47163), .Z(n47165) );
  NOR U60064 ( .A(n47165), .B(n47164), .Z(n47166) );
  IV U60065 ( .A(n47166), .Z(n47171) );
  NOR U60066 ( .A(n48727), .B(n47171), .Z(n47167) );
  NOR U60067 ( .A(n47168), .B(n47167), .Z(n47172) );
  NOR U60068 ( .A(n47169), .B(n47172), .Z(n54215) );
  XOR U60069 ( .A(n48725), .B(n52386), .Z(n47170) );
  NOR U60070 ( .A(n47171), .B(n47170), .Z(n52369) );
  NOR U60071 ( .A(n52369), .B(n47172), .Z(n54221) );
  NOR U60072 ( .A(n47173), .B(n54221), .Z(n47174) );
  NOR U60073 ( .A(n54215), .B(n47174), .Z(n47186) );
  IV U60074 ( .A(n47186), .Z(n50685) );
  NOR U60075 ( .A(n47175), .B(n54222), .Z(n47185) );
  IV U60076 ( .A(n47176), .Z(n47178) );
  NOR U60077 ( .A(n47178), .B(n47177), .Z(n50684) );
  NOR U60078 ( .A(n47185), .B(n50684), .Z(n47179) );
  XOR U60079 ( .A(n50685), .B(n47179), .Z(n47189) );
  IV U60080 ( .A(n47189), .Z(n47180) );
  NOR U60081 ( .A(n47181), .B(n47180), .Z(n50688) );
  IV U60082 ( .A(n47182), .Z(n47184) );
  NOR U60083 ( .A(n47184), .B(n47183), .Z(n47190) );
  IV U60084 ( .A(n47190), .Z(n47188) );
  IV U60085 ( .A(n47185), .Z(n48724) );
  XOR U60086 ( .A(n48724), .B(n47186), .Z(n47187) );
  NOR U60087 ( .A(n47188), .B(n47187), .Z(n54235) );
  NOR U60088 ( .A(n47190), .B(n47189), .Z(n47191) );
  NOR U60089 ( .A(n54235), .B(n47191), .Z(n47192) );
  NOR U60090 ( .A(n47193), .B(n47192), .Z(n47194) );
  NOR U60091 ( .A(n50688), .B(n47194), .Z(n47195) );
  IV U60092 ( .A(n47195), .Z(n50691) );
  XOR U60093 ( .A(n50690), .B(n50691), .Z(n50696) );
  IV U60094 ( .A(n50696), .Z(n47202) );
  IV U60095 ( .A(n47196), .Z(n47198) );
  NOR U60096 ( .A(n47198), .B(n47197), .Z(n48722) );
  NOR U60097 ( .A(n47200), .B(n47199), .Z(n50695) );
  NOR U60098 ( .A(n48722), .B(n50695), .Z(n47201) );
  XOR U60099 ( .A(n47202), .B(n47201), .Z(n50700) );
  XOR U60100 ( .A(n50698), .B(n50700), .Z(n50702) );
  XOR U60101 ( .A(n50703), .B(n50702), .Z(n50714) );
  XOR U60102 ( .A(n47203), .B(n50714), .Z(n48720) );
  NOR U60103 ( .A(n47205), .B(n47204), .Z(n48717) );
  IV U60104 ( .A(n47206), .Z(n47216) );
  IV U60105 ( .A(n47207), .Z(n47208) );
  NOR U60106 ( .A(n47216), .B(n47208), .Z(n48719) );
  NOR U60107 ( .A(n48717), .B(n48719), .Z(n47209) );
  XOR U60108 ( .A(n48720), .B(n47209), .Z(n47220) );
  IV U60109 ( .A(n47220), .Z(n47214) );
  IV U60110 ( .A(n47210), .Z(n47212) );
  NOR U60111 ( .A(n47212), .B(n47211), .Z(n47224) );
  IV U60112 ( .A(n47224), .Z(n47213) );
  NOR U60113 ( .A(n47214), .B(n47213), .Z(n54283) );
  IV U60114 ( .A(n47215), .Z(n47217) );
  NOR U60115 ( .A(n47217), .B(n47216), .Z(n47221) );
  IV U60116 ( .A(n47221), .Z(n47219) );
  XOR U60117 ( .A(n48717), .B(n48720), .Z(n47218) );
  NOR U60118 ( .A(n47219), .B(n47218), .Z(n48716) );
  NOR U60119 ( .A(n47221), .B(n47220), .Z(n47222) );
  NOR U60120 ( .A(n48716), .B(n47222), .Z(n47223) );
  NOR U60121 ( .A(n47224), .B(n47223), .Z(n47225) );
  NOR U60122 ( .A(n54283), .B(n47225), .Z(n50719) );
  XOR U60123 ( .A(n47226), .B(n50719), .Z(n50725) );
  XOR U60124 ( .A(n50723), .B(n50725), .Z(n50735) );
  XOR U60125 ( .A(n50736), .B(n50735), .Z(n48704) );
  NOR U60126 ( .A(n47227), .B(n48709), .Z(n47230) );
  IV U60127 ( .A(n47228), .Z(n47229) );
  NOR U60128 ( .A(n47233), .B(n47229), .Z(n48703) );
  NOR U60129 ( .A(n47230), .B(n48703), .Z(n47231) );
  XOR U60130 ( .A(n48704), .B(n47231), .Z(n50748) );
  IV U60131 ( .A(n47232), .Z(n47236) );
  NOR U60132 ( .A(n47234), .B(n47233), .Z(n47235) );
  IV U60133 ( .A(n47235), .Z(n47245) );
  NOR U60134 ( .A(n47236), .B(n47245), .Z(n50746) );
  XOR U60135 ( .A(n50748), .B(n50746), .Z(n50751) );
  IV U60136 ( .A(n47237), .Z(n47238) );
  NOR U60137 ( .A(n47241), .B(n47238), .Z(n47248) );
  IV U60138 ( .A(n47248), .Z(n47239) );
  NOR U60139 ( .A(n50751), .B(n47239), .Z(n52341) );
  IV U60140 ( .A(n47240), .Z(n47242) );
  NOR U60141 ( .A(n47242), .B(n47241), .Z(n47243) );
  IV U60142 ( .A(n47243), .Z(n48702) );
  IV U60143 ( .A(n47244), .Z(n47246) );
  NOR U60144 ( .A(n47246), .B(n47245), .Z(n50749) );
  XOR U60145 ( .A(n50751), .B(n50749), .Z(n48701) );
  XOR U60146 ( .A(n48702), .B(n48701), .Z(n47247) );
  NOR U60147 ( .A(n47248), .B(n47247), .Z(n47249) );
  NOR U60148 ( .A(n52341), .B(n47249), .Z(n47250) );
  IV U60149 ( .A(n47250), .Z(n48699) );
  IV U60150 ( .A(n47251), .Z(n47252) );
  NOR U60151 ( .A(n47253), .B(n47252), .Z(n48698) );
  XOR U60152 ( .A(n48699), .B(n48698), .Z(n50760) );
  XOR U60153 ( .A(n50759), .B(n50760), .Z(n50756) );
  XOR U60154 ( .A(n47254), .B(n50756), .Z(n47255) );
  IV U60155 ( .A(n47255), .Z(n48691) );
  XOR U60156 ( .A(n48689), .B(n48691), .Z(n48693) );
  IV U60157 ( .A(n47256), .Z(n47258) );
  NOR U60158 ( .A(n47258), .B(n47257), .Z(n47259) );
  IV U60159 ( .A(n47259), .Z(n48692) );
  XOR U60160 ( .A(n48693), .B(n48692), .Z(n47260) );
  NOR U60161 ( .A(n47261), .B(n47260), .Z(n48687) );
  IV U60162 ( .A(n47261), .Z(n47262) );
  NOR U60163 ( .A(n48691), .B(n47262), .Z(n52331) );
  NOR U60164 ( .A(n48687), .B(n52331), .Z(n47263) );
  IV U60165 ( .A(n47263), .Z(n54311) );
  IV U60166 ( .A(n47264), .Z(n47266) );
  NOR U60167 ( .A(n47266), .B(n47265), .Z(n47271) );
  IV U60168 ( .A(n47267), .Z(n47268) );
  NOR U60169 ( .A(n47269), .B(n47268), .Z(n47270) );
  NOR U60170 ( .A(n47271), .B(n47270), .Z(n54312) );
  IV U60171 ( .A(n54312), .Z(n48686) );
  XOR U60172 ( .A(n54311), .B(n48686), .Z(n48684) );
  XOR U60173 ( .A(n48685), .B(n48684), .Z(n47279) );
  IV U60174 ( .A(n47279), .Z(n47272) );
  NOR U60175 ( .A(n47273), .B(n47272), .Z(n54337) );
  IV U60176 ( .A(n47274), .Z(n47276) );
  NOR U60177 ( .A(n47276), .B(n47275), .Z(n47277) );
  IV U60178 ( .A(n47277), .Z(n48683) );
  IV U60179 ( .A(n47280), .Z(n47278) );
  NOR U60180 ( .A(n47278), .B(n48684), .Z(n52330) );
  NOR U60181 ( .A(n47280), .B(n47279), .Z(n47281) );
  NOR U60182 ( .A(n52330), .B(n47281), .Z(n47282) );
  IV U60183 ( .A(n47282), .Z(n48682) );
  XOR U60184 ( .A(n48683), .B(n48682), .Z(n47283) );
  NOR U60185 ( .A(n47284), .B(n47283), .Z(n54341) );
  NOR U60186 ( .A(n54337), .B(n54341), .Z(n48676) );
  IV U60187 ( .A(n47285), .Z(n47287) );
  NOR U60188 ( .A(n47287), .B(n47286), .Z(n54338) );
  IV U60189 ( .A(n47288), .Z(n47289) );
  NOR U60190 ( .A(n47290), .B(n47289), .Z(n52324) );
  NOR U60191 ( .A(n54338), .B(n52324), .Z(n48677) );
  XOR U60192 ( .A(n48676), .B(n48677), .Z(n48680) );
  XOR U60193 ( .A(n47291), .B(n48680), .Z(n48658) );
  XOR U60194 ( .A(n47292), .B(n48658), .Z(n48655) );
  XOR U60195 ( .A(n47293), .B(n48655), .Z(n47294) );
  IV U60196 ( .A(n47294), .Z(n48650) );
  XOR U60197 ( .A(n48648), .B(n48650), .Z(n50792) );
  IV U60198 ( .A(n50792), .Z(n47302) );
  IV U60199 ( .A(n47295), .Z(n47296) );
  NOR U60200 ( .A(n47297), .B(n47296), .Z(n50791) );
  IV U60201 ( .A(n47298), .Z(n47300) );
  NOR U60202 ( .A(n47300), .B(n47299), .Z(n48645) );
  NOR U60203 ( .A(n50791), .B(n48645), .Z(n47301) );
  XOR U60204 ( .A(n47302), .B(n47301), .Z(n50800) );
  IV U60205 ( .A(n47303), .Z(n47305) );
  NOR U60206 ( .A(n47305), .B(n47304), .Z(n50798) );
  XOR U60207 ( .A(n50800), .B(n50798), .Z(n50803) );
  XOR U60208 ( .A(n47306), .B(n50803), .Z(n48638) );
  IV U60209 ( .A(n47307), .Z(n47308) );
  NOR U60210 ( .A(n47309), .B(n47308), .Z(n48640) );
  IV U60211 ( .A(n47310), .Z(n47312) );
  NOR U60212 ( .A(n47312), .B(n47311), .Z(n48637) );
  NOR U60213 ( .A(n48640), .B(n48637), .Z(n47313) );
  XOR U60214 ( .A(n48638), .B(n47313), .Z(n48636) );
  IV U60215 ( .A(n47314), .Z(n47316) );
  NOR U60216 ( .A(n47316), .B(n47315), .Z(n48634) );
  IV U60217 ( .A(n47317), .Z(n47318) );
  NOR U60218 ( .A(n47319), .B(n47318), .Z(n48632) );
  NOR U60219 ( .A(n48634), .B(n48632), .Z(n47320) );
  XOR U60220 ( .A(n48636), .B(n47320), .Z(n48620) );
  IV U60221 ( .A(n47321), .Z(n47322) );
  NOR U60222 ( .A(n47323), .B(n47322), .Z(n48629) );
  IV U60223 ( .A(n47324), .Z(n47326) );
  NOR U60224 ( .A(n47326), .B(n47325), .Z(n48619) );
  NOR U60225 ( .A(n48629), .B(n48619), .Z(n47327) );
  XOR U60226 ( .A(n48620), .B(n47327), .Z(n48624) );
  XOR U60227 ( .A(n47328), .B(n48624), .Z(n47341) );
  IV U60228 ( .A(n47329), .Z(n47330) );
  NOR U60229 ( .A(n47331), .B(n47330), .Z(n47332) );
  IV U60230 ( .A(n47332), .Z(n47345) );
  NOR U60231 ( .A(n47341), .B(n47345), .Z(n52280) );
  IV U60232 ( .A(n47333), .Z(n47335) );
  NOR U60233 ( .A(n47335), .B(n47334), .Z(n47336) );
  IV U60234 ( .A(n47336), .Z(n50810) );
  IV U60235 ( .A(n47337), .Z(n47339) );
  NOR U60236 ( .A(n47339), .B(n47338), .Z(n47343) );
  IV U60237 ( .A(n47343), .Z(n47340) );
  NOR U60238 ( .A(n48624), .B(n47340), .Z(n54384) );
  IV U60239 ( .A(n47341), .Z(n47342) );
  NOR U60240 ( .A(n47343), .B(n47342), .Z(n47344) );
  NOR U60241 ( .A(n54384), .B(n47344), .Z(n47346) );
  IV U60242 ( .A(n47346), .Z(n50809) );
  XOR U60243 ( .A(n50810), .B(n50809), .Z(n47348) );
  NOR U60244 ( .A(n47346), .B(n47345), .Z(n47347) );
  NOR U60245 ( .A(n47348), .B(n47347), .Z(n47349) );
  NOR U60246 ( .A(n52280), .B(n47349), .Z(n52270) );
  XOR U60247 ( .A(n47350), .B(n52270), .Z(n50821) );
  IV U60248 ( .A(n47351), .Z(n47362) );
  IV U60249 ( .A(n47352), .Z(n47353) );
  NOR U60250 ( .A(n47362), .B(n47353), .Z(n50819) );
  IV U60251 ( .A(n47354), .Z(n47355) );
  NOR U60252 ( .A(n47356), .B(n47355), .Z(n50815) );
  NOR U60253 ( .A(n50819), .B(n50815), .Z(n47357) );
  XOR U60254 ( .A(n50821), .B(n47357), .Z(n48613) );
  IV U60255 ( .A(n47358), .Z(n47359) );
  NOR U60256 ( .A(n47366), .B(n47359), .Z(n48614) );
  IV U60257 ( .A(n47360), .Z(n47361) );
  NOR U60258 ( .A(n47362), .B(n47361), .Z(n48616) );
  NOR U60259 ( .A(n48614), .B(n48616), .Z(n47363) );
  XOR U60260 ( .A(n48613), .B(n47363), .Z(n48611) );
  IV U60261 ( .A(n47364), .Z(n47365) );
  NOR U60262 ( .A(n47366), .B(n47365), .Z(n48610) );
  IV U60263 ( .A(n47367), .Z(n47369) );
  NOR U60264 ( .A(n47369), .B(n47368), .Z(n48605) );
  NOR U60265 ( .A(n48610), .B(n48605), .Z(n47370) );
  XOR U60266 ( .A(n48611), .B(n47370), .Z(n48607) );
  XOR U60267 ( .A(n48608), .B(n48607), .Z(n50829) );
  NOR U60268 ( .A(n47376), .B(n50829), .Z(n55806) );
  IV U60269 ( .A(n47371), .Z(n47372) );
  NOR U60270 ( .A(n47373), .B(n47372), .Z(n48596) );
  NOR U60271 ( .A(n55806), .B(n48596), .Z(n47374) );
  IV U60272 ( .A(n47374), .Z(n47375) );
  NOR U60273 ( .A(n47376), .B(n47375), .Z(n47385) );
  NOR U60274 ( .A(n47378), .B(n47377), .Z(n47379) );
  IV U60275 ( .A(n47379), .Z(n47381) );
  NOR U60276 ( .A(n47381), .B(n47380), .Z(n47382) );
  XOR U60277 ( .A(n47382), .B(n50829), .Z(n48597) );
  XOR U60278 ( .A(n48596), .B(n48597), .Z(n47383) );
  NOR U60279 ( .A(n55806), .B(n47383), .Z(n47384) );
  NOR U60280 ( .A(n47385), .B(n47384), .Z(n48589) );
  XOR U60281 ( .A(n48588), .B(n48589), .Z(n48591) );
  IV U60282 ( .A(n47386), .Z(n47397) );
  IV U60283 ( .A(n47387), .Z(n47388) );
  NOR U60284 ( .A(n47397), .B(n47388), .Z(n48585) );
  XOR U60285 ( .A(n48591), .B(n48585), .Z(n47389) );
  XOR U60286 ( .A(n47390), .B(n47389), .Z(n48581) );
  NOR U60287 ( .A(n47391), .B(n48581), .Z(n52220) );
  IV U60288 ( .A(n47392), .Z(n47394) );
  NOR U60289 ( .A(n47394), .B(n47393), .Z(n48582) );
  IV U60290 ( .A(n47395), .Z(n47396) );
  NOR U60291 ( .A(n47397), .B(n47396), .Z(n48579) );
  XOR U60292 ( .A(n48581), .B(n48579), .Z(n48583) );
  XOR U60293 ( .A(n48582), .B(n48583), .Z(n47406) );
  IV U60294 ( .A(n47406), .Z(n47398) );
  NOR U60295 ( .A(n47399), .B(n47398), .Z(n47400) );
  NOR U60296 ( .A(n52220), .B(n47400), .Z(n47408) );
  IV U60297 ( .A(n47408), .Z(n47401) );
  NOR U60298 ( .A(n47411), .B(n47401), .Z(n52212) );
  IV U60299 ( .A(n47402), .Z(n48575) );
  IV U60300 ( .A(n47403), .Z(n47405) );
  NOR U60301 ( .A(n47405), .B(n47404), .Z(n47409) );
  IV U60302 ( .A(n47409), .Z(n47407) );
  NOR U60303 ( .A(n47407), .B(n47406), .Z(n52223) );
  NOR U60304 ( .A(n47409), .B(n47408), .Z(n47410) );
  NOR U60305 ( .A(n52223), .B(n47410), .Z(n47412) );
  IV U60306 ( .A(n47412), .Z(n48574) );
  XOR U60307 ( .A(n48575), .B(n48574), .Z(n47414) );
  NOR U60308 ( .A(n47412), .B(n47411), .Z(n47413) );
  NOR U60309 ( .A(n47414), .B(n47413), .Z(n47415) );
  NOR U60310 ( .A(n52212), .B(n47415), .Z(n47425) );
  XOR U60311 ( .A(n48576), .B(n47425), .Z(n47427) );
  IV U60312 ( .A(n47427), .Z(n47416) );
  NOR U60313 ( .A(n47417), .B(n47416), .Z(n52204) );
  IV U60314 ( .A(n47418), .Z(n47420) );
  NOR U60315 ( .A(n47420), .B(n47419), .Z(n47421) );
  IV U60316 ( .A(n47421), .Z(n50841) );
  IV U60317 ( .A(n47422), .Z(n47424) );
  NOR U60318 ( .A(n47424), .B(n47423), .Z(n47428) );
  IV U60319 ( .A(n47428), .Z(n47426) );
  IV U60320 ( .A(n47425), .Z(n48577) );
  NOR U60321 ( .A(n47426), .B(n48577), .Z(n50843) );
  NOR U60322 ( .A(n47428), .B(n47427), .Z(n47429) );
  NOR U60323 ( .A(n50843), .B(n47429), .Z(n47430) );
  IV U60324 ( .A(n47430), .Z(n50840) );
  XOR U60325 ( .A(n50841), .B(n50840), .Z(n47431) );
  NOR U60326 ( .A(n47432), .B(n47431), .Z(n47433) );
  NOR U60327 ( .A(n52204), .B(n47433), .Z(n48569) );
  NOR U60328 ( .A(n47435), .B(n47434), .Z(n48571) );
  IV U60329 ( .A(n47436), .Z(n47437) );
  NOR U60330 ( .A(n47437), .B(n47440), .Z(n48568) );
  NOR U60331 ( .A(n48571), .B(n48568), .Z(n47438) );
  XOR U60332 ( .A(n48569), .B(n47438), .Z(n48567) );
  IV U60333 ( .A(n47439), .Z(n47441) );
  NOR U60334 ( .A(n47441), .B(n47440), .Z(n48565) );
  XOR U60335 ( .A(n48567), .B(n48565), .Z(n48562) );
  XOR U60336 ( .A(n48561), .B(n48562), .Z(n52189) );
  XOR U60337 ( .A(n48556), .B(n52189), .Z(n48554) );
  IV U60338 ( .A(n47442), .Z(n47444) );
  NOR U60339 ( .A(n47444), .B(n47443), .Z(n48557) );
  IV U60340 ( .A(n47445), .Z(n47447) );
  NOR U60341 ( .A(n47447), .B(n47446), .Z(n48553) );
  NOR U60342 ( .A(n48557), .B(n48553), .Z(n47448) );
  XOR U60343 ( .A(n48554), .B(n47448), .Z(n48552) );
  IV U60344 ( .A(n47449), .Z(n47450) );
  NOR U60345 ( .A(n47451), .B(n47450), .Z(n48550) );
  IV U60346 ( .A(n47452), .Z(n47453) );
  NOR U60347 ( .A(n47454), .B(n47453), .Z(n48545) );
  NOR U60348 ( .A(n48550), .B(n48545), .Z(n47455) );
  XOR U60349 ( .A(n48552), .B(n47455), .Z(n48541) );
  IV U60350 ( .A(n47456), .Z(n47457) );
  NOR U60351 ( .A(n47458), .B(n47457), .Z(n48547) );
  IV U60352 ( .A(n47459), .Z(n47461) );
  NOR U60353 ( .A(n47461), .B(n47460), .Z(n48542) );
  NOR U60354 ( .A(n48547), .B(n48542), .Z(n52170) );
  XOR U60355 ( .A(n48541), .B(n52170), .Z(n48540) );
  XOR U60356 ( .A(n47462), .B(n48540), .Z(n47463) );
  IV U60357 ( .A(n47463), .Z(n48533) );
  XOR U60358 ( .A(n48532), .B(n48533), .Z(n47471) );
  IV U60359 ( .A(n47471), .Z(n47464) );
  NOR U60360 ( .A(n47465), .B(n47464), .Z(n47477) );
  IV U60361 ( .A(n47466), .Z(n47469) );
  NOR U60362 ( .A(n47472), .B(n48533), .Z(n47467) );
  IV U60363 ( .A(n47467), .Z(n47468) );
  NOR U60364 ( .A(n47469), .B(n47468), .Z(n52164) );
  IV U60365 ( .A(n47470), .Z(n47475) );
  NOR U60366 ( .A(n47472), .B(n47471), .Z(n47473) );
  IV U60367 ( .A(n47473), .Z(n47474) );
  NOR U60368 ( .A(n47475), .B(n47474), .Z(n52162) );
  NOR U60369 ( .A(n52164), .B(n52162), .Z(n47476) );
  IV U60370 ( .A(n47476), .Z(n48535) );
  NOR U60371 ( .A(n47477), .B(n48535), .Z(n47478) );
  IV U60372 ( .A(n47478), .Z(n48528) );
  XOR U60373 ( .A(n48527), .B(n48528), .Z(n48522) );
  IV U60374 ( .A(n48522), .Z(n47486) );
  IV U60375 ( .A(n47479), .Z(n47481) );
  NOR U60376 ( .A(n47481), .B(n47480), .Z(n48524) );
  IV U60377 ( .A(n47482), .Z(n47484) );
  NOR U60378 ( .A(n47484), .B(n47483), .Z(n48521) );
  NOR U60379 ( .A(n48524), .B(n48521), .Z(n47485) );
  XOR U60380 ( .A(n47486), .B(n47485), .Z(n48520) );
  XOR U60381 ( .A(n48516), .B(n48520), .Z(n48514) );
  XOR U60382 ( .A(n47487), .B(n48514), .Z(n47488) );
  IV U60383 ( .A(n47488), .Z(n50858) );
  XOR U60384 ( .A(n48511), .B(n50858), .Z(n50860) );
  IV U60385 ( .A(n47489), .Z(n47491) );
  NOR U60386 ( .A(n47491), .B(n47490), .Z(n50856) );
  IV U60387 ( .A(n47492), .Z(n47493) );
  NOR U60388 ( .A(n47493), .B(n47496), .Z(n50859) );
  NOR U60389 ( .A(n50856), .B(n50859), .Z(n47494) );
  XOR U60390 ( .A(n50860), .B(n47494), .Z(n50862) );
  IV U60391 ( .A(n47495), .Z(n47497) );
  NOR U60392 ( .A(n47497), .B(n47496), .Z(n52146) );
  IV U60393 ( .A(n47498), .Z(n47500) );
  NOR U60394 ( .A(n47500), .B(n47499), .Z(n52139) );
  NOR U60395 ( .A(n52146), .B(n52139), .Z(n50863) );
  XOR U60396 ( .A(n50862), .B(n50863), .Z(n50865) );
  IV U60397 ( .A(n47501), .Z(n47503) );
  NOR U60398 ( .A(n47503), .B(n47502), .Z(n50864) );
  IV U60399 ( .A(n47504), .Z(n47506) );
  NOR U60400 ( .A(n47506), .B(n47505), .Z(n48509) );
  NOR U60401 ( .A(n50864), .B(n48509), .Z(n47507) );
  XOR U60402 ( .A(n50865), .B(n47507), .Z(n47512) );
  IV U60403 ( .A(n47512), .Z(n47511) );
  IV U60404 ( .A(n47508), .Z(n47509) );
  NOR U60405 ( .A(n47509), .B(n47516), .Z(n47513) );
  IV U60406 ( .A(n47513), .Z(n47510) );
  NOR U60407 ( .A(n47511), .B(n47510), .Z(n52133) );
  NOR U60408 ( .A(n47513), .B(n47512), .Z(n50870) );
  NOR U60409 ( .A(n52133), .B(n50870), .Z(n52126) );
  IV U60410 ( .A(n47514), .Z(n47515) );
  NOR U60411 ( .A(n47516), .B(n47515), .Z(n47521) );
  IV U60412 ( .A(n47517), .Z(n47519) );
  IV U60413 ( .A(n47518), .Z(n47523) );
  NOR U60414 ( .A(n47519), .B(n47523), .Z(n47520) );
  NOR U60415 ( .A(n47521), .B(n47520), .Z(n52128) );
  XOR U60416 ( .A(n52126), .B(n52128), .Z(n50875) );
  IV U60417 ( .A(n47522), .Z(n47524) );
  NOR U60418 ( .A(n47524), .B(n47523), .Z(n50873) );
  XOR U60419 ( .A(n50875), .B(n50873), .Z(n50877) );
  XOR U60420 ( .A(n50876), .B(n50877), .Z(n48507) );
  XOR U60421 ( .A(n48506), .B(n48507), .Z(n48502) );
  IV U60422 ( .A(n48502), .Z(n47532) );
  IV U60423 ( .A(n47525), .Z(n47527) );
  NOR U60424 ( .A(n47527), .B(n47526), .Z(n48504) );
  IV U60425 ( .A(n47528), .Z(n47530) );
  NOR U60426 ( .A(n47530), .B(n47529), .Z(n48501) );
  NOR U60427 ( .A(n48504), .B(n48501), .Z(n47531) );
  XOR U60428 ( .A(n47532), .B(n47531), .Z(n50882) );
  XOR U60429 ( .A(n50880), .B(n50882), .Z(n50884) );
  XOR U60430 ( .A(n50883), .B(n50884), .Z(n48497) );
  XOR U60431 ( .A(n47533), .B(n48497), .Z(n48490) );
  XOR U60432 ( .A(n47534), .B(n48490), .Z(n48488) );
  XOR U60433 ( .A(n47535), .B(n48488), .Z(n48475) );
  NOR U60434 ( .A(n47536), .B(n48484), .Z(n47540) );
  IV U60435 ( .A(n47537), .Z(n48476) );
  NOR U60436 ( .A(n47538), .B(n48476), .Z(n47539) );
  NOR U60437 ( .A(n47540), .B(n47539), .Z(n47541) );
  XOR U60438 ( .A(n48475), .B(n47541), .Z(n50899) );
  IV U60439 ( .A(n47542), .Z(n47543) );
  NOR U60440 ( .A(n47545), .B(n47543), .Z(n47544) );
  IV U60441 ( .A(n47544), .Z(n47552) );
  NOR U60442 ( .A(n50899), .B(n47552), .Z(n52086) );
  NOR U60443 ( .A(n47546), .B(n47545), .Z(n47547) );
  IV U60444 ( .A(n47547), .Z(n50898) );
  NOR U60445 ( .A(n50901), .B(n50898), .Z(n47548) );
  XOR U60446 ( .A(n50899), .B(n47548), .Z(n48473) );
  IV U60447 ( .A(n47549), .Z(n47551) );
  NOR U60448 ( .A(n47551), .B(n47550), .Z(n47553) );
  IV U60449 ( .A(n47553), .Z(n48472) );
  XOR U60450 ( .A(n48473), .B(n48472), .Z(n47555) );
  NOR U60451 ( .A(n47553), .B(n47552), .Z(n47554) );
  NOR U60452 ( .A(n47555), .B(n47554), .Z(n47556) );
  NOR U60453 ( .A(n52086), .B(n47556), .Z(n47558) );
  XOR U60454 ( .A(n48469), .B(n47558), .Z(n47566) );
  IV U60455 ( .A(n47566), .Z(n48463) );
  NOR U60456 ( .A(n47557), .B(n48463), .Z(n54490) );
  IV U60457 ( .A(n47558), .Z(n48471) );
  NOR U60458 ( .A(n47565), .B(n48471), .Z(n47559) );
  IV U60459 ( .A(n47559), .Z(n47560) );
  NOR U60460 ( .A(n47561), .B(n47560), .Z(n47562) );
  IV U60461 ( .A(n47562), .Z(n52077) );
  NOR U60462 ( .A(n47563), .B(n52077), .Z(n50907) );
  NOR U60463 ( .A(n47565), .B(n47564), .Z(n47567) );
  NOR U60464 ( .A(n47567), .B(n47566), .Z(n47568) );
  NOR U60465 ( .A(n50907), .B(n47568), .Z(n48465) );
  NOR U60466 ( .A(n47569), .B(n48465), .Z(n47570) );
  NOR U60467 ( .A(n54490), .B(n47570), .Z(n47578) );
  IV U60468 ( .A(n47571), .Z(n47576) );
  NOR U60469 ( .A(n47573), .B(n47572), .Z(n47574) );
  IV U60470 ( .A(n47574), .Z(n47575) );
  NOR U60471 ( .A(n47576), .B(n47575), .Z(n48466) );
  NOR U60472 ( .A(n48462), .B(n48466), .Z(n47577) );
  XOR U60473 ( .A(n47578), .B(n47577), .Z(n50911) );
  IV U60474 ( .A(n47579), .Z(n47581) );
  IV U60475 ( .A(n47580), .Z(n47583) );
  NOR U60476 ( .A(n47581), .B(n47583), .Z(n50909) );
  XOR U60477 ( .A(n50911), .B(n50909), .Z(n54499) );
  IV U60478 ( .A(n47582), .Z(n47584) );
  NOR U60479 ( .A(n47584), .B(n47583), .Z(n54497) );
  IV U60480 ( .A(n47585), .Z(n47587) );
  NOR U60481 ( .A(n47587), .B(n47586), .Z(n54502) );
  NOR U60482 ( .A(n54497), .B(n54502), .Z(n50912) );
  XOR U60483 ( .A(n54499), .B(n50912), .Z(n50920) );
  XOR U60484 ( .A(n50921), .B(n50920), .Z(n50918) );
  IV U60485 ( .A(n47588), .Z(n47590) );
  NOR U60486 ( .A(n47590), .B(n47589), .Z(n50916) );
  XOR U60487 ( .A(n50918), .B(n50916), .Z(n50931) );
  XOR U60488 ( .A(n50923), .B(n50931), .Z(n50935) );
  IV U60489 ( .A(n50935), .Z(n47600) );
  IV U60490 ( .A(n47591), .Z(n47592) );
  NOR U60491 ( .A(n47593), .B(n47592), .Z(n50930) );
  IV U60492 ( .A(n47594), .Z(n47598) );
  NOR U60493 ( .A(n47596), .B(n47595), .Z(n47597) );
  IV U60494 ( .A(n47597), .Z(n47602) );
  NOR U60495 ( .A(n47598), .B(n47602), .Z(n50933) );
  NOR U60496 ( .A(n50930), .B(n50933), .Z(n47599) );
  XOR U60497 ( .A(n47600), .B(n47599), .Z(n48458) );
  IV U60498 ( .A(n47601), .Z(n47603) );
  NOR U60499 ( .A(n47603), .B(n47602), .Z(n48456) );
  XOR U60500 ( .A(n48458), .B(n48456), .Z(n48461) );
  XOR U60501 ( .A(n47604), .B(n48461), .Z(n50940) );
  IV U60502 ( .A(n47605), .Z(n47607) );
  NOR U60503 ( .A(n47607), .B(n47606), .Z(n52049) );
  IV U60504 ( .A(n47608), .Z(n47609) );
  NOR U60505 ( .A(n47610), .B(n47609), .Z(n52056) );
  NOR U60506 ( .A(n52049), .B(n52056), .Z(n50941) );
  XOR U60507 ( .A(n50940), .B(n50941), .Z(n50944) );
  XOR U60508 ( .A(n50942), .B(n50944), .Z(n50949) );
  XOR U60509 ( .A(n50947), .B(n50949), .Z(n50956) );
  XOR U60510 ( .A(n50950), .B(n50956), .Z(n50959) );
  XOR U60511 ( .A(n47611), .B(n50959), .Z(n50960) );
  XOR U60512 ( .A(n47612), .B(n50960), .Z(n48452) );
  NOR U60513 ( .A(n47620), .B(n48452), .Z(n50971) );
  IV U60514 ( .A(n47613), .Z(n47615) );
  NOR U60515 ( .A(n47615), .B(n47614), .Z(n47616) );
  IV U60516 ( .A(n47616), .Z(n48445) );
  IV U60517 ( .A(n47617), .Z(n47618) );
  NOR U60518 ( .A(n47619), .B(n47618), .Z(n48451) );
  XOR U60519 ( .A(n48451), .B(n48452), .Z(n48444) );
  XOR U60520 ( .A(n48445), .B(n48444), .Z(n47623) );
  IV U60521 ( .A(n48444), .Z(n47621) );
  NOR U60522 ( .A(n47621), .B(n47620), .Z(n47622) );
  NOR U60523 ( .A(n47623), .B(n47622), .Z(n47624) );
  NOR U60524 ( .A(n50971), .B(n47624), .Z(n48446) );
  XOR U60525 ( .A(n48448), .B(n48446), .Z(n48439) );
  XOR U60526 ( .A(n48436), .B(n48439), .Z(n50977) );
  NOR U60527 ( .A(n47628), .B(n50977), .Z(n54524) );
  NOR U60528 ( .A(n47625), .B(n48440), .Z(n50976) );
  XOR U60529 ( .A(n50976), .B(n50977), .Z(n52013) );
  IV U60530 ( .A(n47626), .Z(n47627) );
  NOR U60531 ( .A(n48432), .B(n47627), .Z(n47629) );
  IV U60532 ( .A(n47629), .Z(n52012) );
  XOR U60533 ( .A(n52013), .B(n52012), .Z(n47631) );
  NOR U60534 ( .A(n47629), .B(n47628), .Z(n47630) );
  NOR U60535 ( .A(n47631), .B(n47630), .Z(n47632) );
  NOR U60536 ( .A(n54524), .B(n47632), .Z(n48429) );
  XOR U60537 ( .A(n47633), .B(n48429), .Z(n50987) );
  XOR U60538 ( .A(n47634), .B(n50987), .Z(n50988) );
  XOR U60539 ( .A(n50989), .B(n50988), .Z(n50999) );
  XOR U60540 ( .A(n47635), .B(n50999), .Z(n50995) );
  XOR U60541 ( .A(n47636), .B(n50995), .Z(n51009) );
  XOR U60542 ( .A(n47637), .B(n51009), .Z(n48422) );
  XOR U60543 ( .A(n48423), .B(n48422), .Z(n48418) );
  XOR U60544 ( .A(n48417), .B(n48418), .Z(n48414) );
  IV U60545 ( .A(n47638), .Z(n47639) );
  NOR U60546 ( .A(n47640), .B(n47639), .Z(n48419) );
  IV U60547 ( .A(n47641), .Z(n47643) );
  NOR U60548 ( .A(n47643), .B(n47642), .Z(n48415) );
  NOR U60549 ( .A(n48419), .B(n48415), .Z(n47644) );
  XOR U60550 ( .A(n48414), .B(n47644), .Z(n51017) );
  XOR U60551 ( .A(n51015), .B(n51017), .Z(n48413) );
  IV U60552 ( .A(n47645), .Z(n47646) );
  NOR U60553 ( .A(n47647), .B(n47646), .Z(n48411) );
  XOR U60554 ( .A(n48413), .B(n48411), .Z(n51027) );
  IV U60555 ( .A(n51027), .Z(n47655) );
  IV U60556 ( .A(n47648), .Z(n48408) );
  NOR U60557 ( .A(n48408), .B(n47649), .Z(n47653) );
  IV U60558 ( .A(n47650), .Z(n47652) );
  NOR U60559 ( .A(n47652), .B(n47651), .Z(n51026) );
  NOR U60560 ( .A(n47653), .B(n51026), .Z(n47654) );
  XOR U60561 ( .A(n47655), .B(n47654), .Z(n51035) );
  IV U60562 ( .A(n47656), .Z(n47658) );
  NOR U60563 ( .A(n47658), .B(n47657), .Z(n51033) );
  XOR U60564 ( .A(n51035), .B(n51033), .Z(n51037) );
  XOR U60565 ( .A(n51036), .B(n51037), .Z(n48404) );
  XOR U60566 ( .A(n48403), .B(n48404), .Z(n48402) );
  XOR U60567 ( .A(n47659), .B(n48402), .Z(n48393) );
  NOR U60568 ( .A(n47661), .B(n47660), .Z(n48397) );
  IV U60569 ( .A(n47662), .Z(n47664) );
  NOR U60570 ( .A(n47664), .B(n47663), .Z(n48392) );
  NOR U60571 ( .A(n48397), .B(n48392), .Z(n47665) );
  XOR U60572 ( .A(n48393), .B(n47665), .Z(n51048) );
  XOR U60573 ( .A(n51047), .B(n51048), .Z(n51054) );
  XOR U60574 ( .A(n47666), .B(n51054), .Z(n51056) );
  IV U60575 ( .A(n47667), .Z(n47669) );
  NOR U60576 ( .A(n47669), .B(n47668), .Z(n51937) );
  NOR U60577 ( .A(n47671), .B(n47670), .Z(n54564) );
  NOR U60578 ( .A(n51937), .B(n54564), .Z(n51057) );
  XOR U60579 ( .A(n51056), .B(n51057), .Z(n51061) );
  XOR U60580 ( .A(n51059), .B(n51061), .Z(n51063) );
  XOR U60581 ( .A(n51062), .B(n51063), .Z(n48386) );
  XOR U60582 ( .A(n47672), .B(n48386), .Z(n51074) );
  XOR U60583 ( .A(n51075), .B(n51074), .Z(n48381) );
  XOR U60584 ( .A(n48379), .B(n48381), .Z(n51071) );
  XOR U60585 ( .A(n51070), .B(n51071), .Z(n51085) );
  XOR U60586 ( .A(n47673), .B(n51085), .Z(n48372) );
  IV U60587 ( .A(n47674), .Z(n47675) );
  NOR U60588 ( .A(n47682), .B(n47675), .Z(n47676) );
  IV U60589 ( .A(n47676), .Z(n48373) );
  XOR U60590 ( .A(n48372), .B(n48373), .Z(n51887) );
  IV U60591 ( .A(n47677), .Z(n47678) );
  NOR U60592 ( .A(n47679), .B(n47678), .Z(n51886) );
  IV U60593 ( .A(n47680), .Z(n47681) );
  NOR U60594 ( .A(n47682), .B(n47681), .Z(n51890) );
  NOR U60595 ( .A(n51886), .B(n51890), .Z(n48375) );
  XOR U60596 ( .A(n51887), .B(n48375), .Z(n51088) );
  XOR U60597 ( .A(n51089), .B(n51088), .Z(n51873) );
  NOR U60598 ( .A(n47683), .B(n47685), .Z(n47690) );
  NOR U60599 ( .A(n47685), .B(n47684), .Z(n47686) );
  IV U60600 ( .A(n47686), .Z(n47687) );
  NOR U60601 ( .A(n47688), .B(n47687), .Z(n47689) );
  NOR U60602 ( .A(n47690), .B(n47689), .Z(n51874) );
  IV U60603 ( .A(n51874), .Z(n51090) );
  XOR U60604 ( .A(n51873), .B(n51090), .Z(n47694) );
  IV U60605 ( .A(n47691), .Z(n47692) );
  NOR U60606 ( .A(n47692), .B(n47704), .Z(n47700) );
  IV U60607 ( .A(n47700), .Z(n47693) );
  NOR U60608 ( .A(n47694), .B(n47693), .Z(n54595) );
  IV U60609 ( .A(n47695), .Z(n47696) );
  NOR U60610 ( .A(n47697), .B(n47696), .Z(n48370) );
  NOR U60611 ( .A(n48370), .B(n51090), .Z(n47698) );
  XOR U60612 ( .A(n51873), .B(n47698), .Z(n47699) );
  NOR U60613 ( .A(n47700), .B(n47699), .Z(n47701) );
  NOR U60614 ( .A(n54595), .B(n47701), .Z(n48365) );
  IV U60615 ( .A(n47702), .Z(n47703) );
  NOR U60616 ( .A(n47704), .B(n47703), .Z(n47705) );
  IV U60617 ( .A(n47705), .Z(n48366) );
  XOR U60618 ( .A(n48365), .B(n48366), .Z(n51104) );
  IV U60619 ( .A(n51104), .Z(n47712) );
  NOR U60620 ( .A(n47707), .B(n47706), .Z(n48368) );
  IV U60621 ( .A(n47708), .Z(n47710) );
  IV U60622 ( .A(n47709), .Z(n47714) );
  NOR U60623 ( .A(n47710), .B(n47714), .Z(n51102) );
  NOR U60624 ( .A(n48368), .B(n51102), .Z(n47711) );
  XOR U60625 ( .A(n47712), .B(n47711), .Z(n51101) );
  IV U60626 ( .A(n47713), .Z(n47715) );
  NOR U60627 ( .A(n47715), .B(n47714), .Z(n51099) );
  XOR U60628 ( .A(n51101), .B(n51099), .Z(n51107) );
  XOR U60629 ( .A(n47716), .B(n51107), .Z(n51111) );
  XOR U60630 ( .A(n47717), .B(n51111), .Z(n48360) );
  XOR U60631 ( .A(n47718), .B(n48360), .Z(n51127) );
  XOR U60632 ( .A(n47719), .B(n51127), .Z(n51131) );
  XOR U60633 ( .A(n51130), .B(n51131), .Z(n48355) );
  XOR U60634 ( .A(n48356), .B(n48355), .Z(n47720) );
  IV U60635 ( .A(n47720), .Z(n48348) );
  XOR U60636 ( .A(n48347), .B(n48348), .Z(n48352) );
  IV U60637 ( .A(n47721), .Z(n47722) );
  NOR U60638 ( .A(n47723), .B(n47722), .Z(n48350) );
  XOR U60639 ( .A(n48352), .B(n48350), .Z(n51858) );
  IV U60640 ( .A(n51858), .Z(n47730) );
  IV U60641 ( .A(n47724), .Z(n47725) );
  NOR U60642 ( .A(n47726), .B(n47725), .Z(n51861) );
  IV U60643 ( .A(n47727), .Z(n47728) );
  NOR U60644 ( .A(n47729), .B(n47728), .Z(n51857) );
  NOR U60645 ( .A(n51861), .B(n51857), .Z(n48339) );
  XOR U60646 ( .A(n47730), .B(n48339), .Z(n48344) );
  XOR U60647 ( .A(n47731), .B(n48344), .Z(n47740) );
  IV U60648 ( .A(n47734), .Z(n47742) );
  NOR U60649 ( .A(n47732), .B(n47742), .Z(n47738) );
  IV U60650 ( .A(n47732), .Z(n47733) );
  NOR U60651 ( .A(n47734), .B(n47733), .Z(n47736) );
  IV U60652 ( .A(n47735), .Z(n48336) );
  NOR U60653 ( .A(n47736), .B(n48336), .Z(n47737) );
  NOR U60654 ( .A(n47738), .B(n47737), .Z(n47744) );
  IV U60655 ( .A(n47744), .Z(n47739) );
  NOR U60656 ( .A(n47740), .B(n47739), .Z(n47746) );
  IV U60657 ( .A(n47740), .Z(n47741) );
  NOR U60658 ( .A(n47742), .B(n47741), .Z(n47743) );
  IV U60659 ( .A(n47743), .Z(n51143) );
  NOR U60660 ( .A(n47744), .B(n51143), .Z(n47745) );
  NOR U60661 ( .A(n47746), .B(n47745), .Z(n48330) );
  XOR U60662 ( .A(n47747), .B(n48330), .Z(n48329) );
  XOR U60663 ( .A(n48327), .B(n48329), .Z(n48326) );
  NOR U60664 ( .A(n47751), .B(n48326), .Z(n48324) );
  IV U60665 ( .A(n47748), .Z(n47749) );
  NOR U60666 ( .A(n47750), .B(n47749), .Z(n47752) );
  IV U60667 ( .A(n47752), .Z(n48325) );
  XOR U60668 ( .A(n48326), .B(n48325), .Z(n47754) );
  NOR U60669 ( .A(n47752), .B(n47751), .Z(n47753) );
  NOR U60670 ( .A(n47754), .B(n47753), .Z(n48321) );
  NOR U60671 ( .A(n48324), .B(n48321), .Z(n48317) );
  IV U60672 ( .A(n47755), .Z(n47757) );
  NOR U60673 ( .A(n47757), .B(n47756), .Z(n48320) );
  IV U60674 ( .A(n47758), .Z(n47760) );
  NOR U60675 ( .A(n47760), .B(n47759), .Z(n48316) );
  NOR U60676 ( .A(n48320), .B(n48316), .Z(n47761) );
  XOR U60677 ( .A(n48317), .B(n47761), .Z(n54653) );
  XOR U60678 ( .A(n48314), .B(n54653), .Z(n47763) );
  NOR U60679 ( .A(n47762), .B(n47763), .Z(n48312) );
  IV U60680 ( .A(n47762), .Z(n47765) );
  IV U60681 ( .A(n47763), .Z(n47764) );
  NOR U60682 ( .A(n47765), .B(n47764), .Z(n51827) );
  NOR U60683 ( .A(n48312), .B(n51827), .Z(n48309) );
  IV U60684 ( .A(n47766), .Z(n54666) );
  NOR U60685 ( .A(n54666), .B(n47767), .Z(n54680) );
  IV U60686 ( .A(n47768), .Z(n47769) );
  NOR U60687 ( .A(n47772), .B(n47769), .Z(n48310) );
  NOR U60688 ( .A(n54680), .B(n48310), .Z(n47770) );
  XOR U60689 ( .A(n48309), .B(n47770), .Z(n48308) );
  IV U60690 ( .A(n47771), .Z(n47773) );
  NOR U60691 ( .A(n47773), .B(n47772), .Z(n47774) );
  IV U60692 ( .A(n47774), .Z(n48307) );
  XOR U60693 ( .A(n48308), .B(n48307), .Z(n47781) );
  IV U60694 ( .A(n47781), .Z(n47775) );
  NOR U60695 ( .A(n47776), .B(n47775), .Z(n51819) );
  IV U60696 ( .A(n47777), .Z(n47779) );
  NOR U60697 ( .A(n47779), .B(n47778), .Z(n47782) );
  IV U60698 ( .A(n47782), .Z(n47780) );
  NOR U60699 ( .A(n48308), .B(n47780), .Z(n51815) );
  NOR U60700 ( .A(n47782), .B(n47781), .Z(n47783) );
  NOR U60701 ( .A(n51815), .B(n47783), .Z(n51154) );
  NOR U60702 ( .A(n47784), .B(n51154), .Z(n47785) );
  NOR U60703 ( .A(n51819), .B(n47785), .Z(n48303) );
  NOR U60704 ( .A(n47786), .B(n51156), .Z(n47790) );
  IV U60705 ( .A(n47787), .Z(n47789) );
  IV U60706 ( .A(n47788), .Z(n47796) );
  NOR U60707 ( .A(n47789), .B(n47796), .Z(n48304) );
  NOR U60708 ( .A(n47790), .B(n48304), .Z(n47791) );
  XOR U60709 ( .A(n48303), .B(n47791), .Z(n51799) );
  IV U60710 ( .A(n47792), .Z(n47793) );
  NOR U60711 ( .A(n47794), .B(n47793), .Z(n51798) );
  IV U60712 ( .A(n47795), .Z(n47797) );
  NOR U60713 ( .A(n47797), .B(n47796), .Z(n51802) );
  NOR U60714 ( .A(n51798), .B(n51802), .Z(n48298) );
  XOR U60715 ( .A(n51799), .B(n48298), .Z(n48296) );
  IV U60716 ( .A(n47798), .Z(n47800) );
  NOR U60717 ( .A(n47800), .B(n47799), .Z(n48299) );
  IV U60718 ( .A(n47801), .Z(n47803) );
  NOR U60719 ( .A(n47803), .B(n47802), .Z(n48295) );
  NOR U60720 ( .A(n48299), .B(n48295), .Z(n47804) );
  XOR U60721 ( .A(n48296), .B(n47804), .Z(n51168) );
  IV U60722 ( .A(n47805), .Z(n47807) );
  NOR U60723 ( .A(n47807), .B(n47806), .Z(n48293) );
  IV U60724 ( .A(n47808), .Z(n47810) );
  NOR U60725 ( .A(n47810), .B(n47809), .Z(n51166) );
  NOR U60726 ( .A(n48293), .B(n51166), .Z(n47811) );
  XOR U60727 ( .A(n51168), .B(n47811), .Z(n47812) );
  IV U60728 ( .A(n47812), .Z(n51169) );
  XOR U60729 ( .A(n51170), .B(n51169), .Z(n48288) );
  IV U60730 ( .A(n47813), .Z(n47814) );
  NOR U60731 ( .A(n47815), .B(n47814), .Z(n48291) );
  IV U60732 ( .A(n47816), .Z(n47817) );
  NOR U60733 ( .A(n47824), .B(n47817), .Z(n48287) );
  NOR U60734 ( .A(n48291), .B(n48287), .Z(n47818) );
  XOR U60735 ( .A(n48288), .B(n47818), .Z(n48286) );
  IV U60736 ( .A(n47819), .Z(n47821) );
  NOR U60737 ( .A(n47821), .B(n47820), .Z(n47822) );
  IV U60738 ( .A(n47822), .Z(n47829) );
  NOR U60739 ( .A(n48286), .B(n47829), .Z(n54708) );
  IV U60740 ( .A(n47823), .Z(n47825) );
  NOR U60741 ( .A(n47825), .B(n47824), .Z(n48284) );
  XOR U60742 ( .A(n48284), .B(n48286), .Z(n48283) );
  IV U60743 ( .A(n47826), .Z(n47828) );
  NOR U60744 ( .A(n47828), .B(n47827), .Z(n47830) );
  IV U60745 ( .A(n47830), .Z(n48282) );
  XOR U60746 ( .A(n48283), .B(n48282), .Z(n47832) );
  NOR U60747 ( .A(n47830), .B(n47829), .Z(n47831) );
  NOR U60748 ( .A(n47832), .B(n47831), .Z(n47833) );
  NOR U60749 ( .A(n54708), .B(n47833), .Z(n47834) );
  IV U60750 ( .A(n47834), .Z(n54714) );
  XOR U60751 ( .A(n54712), .B(n54714), .Z(n51175) );
  IV U60752 ( .A(n51175), .Z(n47841) );
  IV U60753 ( .A(n47835), .Z(n47836) );
  NOR U60754 ( .A(n47837), .B(n47836), .Z(n54713) );
  IV U60755 ( .A(n47838), .Z(n47840) );
  NOR U60756 ( .A(n47840), .B(n47839), .Z(n54723) );
  NOR U60757 ( .A(n54713), .B(n54723), .Z(n51176) );
  XOR U60758 ( .A(n47841), .B(n51176), .Z(n51186) );
  XOR U60759 ( .A(n51179), .B(n51186), .Z(n51182) );
  XOR U60760 ( .A(n51181), .B(n51182), .Z(n48280) );
  XOR U60761 ( .A(n47842), .B(n48280), .Z(n47843) );
  IV U60762 ( .A(n47843), .Z(n51195) );
  XOR U60763 ( .A(n51193), .B(n51195), .Z(n51198) );
  IV U60764 ( .A(n47844), .Z(n47846) );
  NOR U60765 ( .A(n47846), .B(n47845), .Z(n51196) );
  XOR U60766 ( .A(n51198), .B(n51196), .Z(n51209) );
  XOR U60767 ( .A(n51208), .B(n51209), .Z(n51201) );
  XOR U60768 ( .A(n51200), .B(n51201), .Z(n51205) );
  XOR U60769 ( .A(n51204), .B(n51205), .Z(n48276) );
  XOR U60770 ( .A(n48275), .B(n48276), .Z(n48272) );
  IV U60771 ( .A(n47847), .Z(n47849) );
  NOR U60772 ( .A(n47849), .B(n47848), .Z(n48273) );
  IV U60773 ( .A(n47850), .Z(n47851) );
  NOR U60774 ( .A(n47851), .B(n47857), .Z(n48270) );
  NOR U60775 ( .A(n48273), .B(n48270), .Z(n47852) );
  XOR U60776 ( .A(n48272), .B(n47852), .Z(n51217) );
  IV U60777 ( .A(n47853), .Z(n51222) );
  NOR U60778 ( .A(n51222), .B(n47854), .Z(n47858) );
  IV U60779 ( .A(n47855), .Z(n47856) );
  NOR U60780 ( .A(n47857), .B(n47856), .Z(n51218) );
  NOR U60781 ( .A(n47858), .B(n51218), .Z(n47859) );
  XOR U60782 ( .A(n51217), .B(n47859), .Z(n51226) );
  XOR U60783 ( .A(n51225), .B(n51226), .Z(n48264) );
  IV U60784 ( .A(n48264), .Z(n47866) );
  NOR U60785 ( .A(n47860), .B(n48267), .Z(n47864) );
  IV U60786 ( .A(n47861), .Z(n47862) );
  NOR U60787 ( .A(n47863), .B(n47862), .Z(n48263) );
  NOR U60788 ( .A(n47864), .B(n48263), .Z(n47865) );
  XOR U60789 ( .A(n47866), .B(n47865), .Z(n48262) );
  XOR U60790 ( .A(n48260), .B(n48262), .Z(n48256) );
  XOR U60791 ( .A(n48255), .B(n48256), .Z(n51244) );
  XOR U60792 ( .A(n47867), .B(n51244), .Z(n48251) );
  XOR U60793 ( .A(n47868), .B(n48251), .Z(n51252) );
  XOR U60794 ( .A(n51251), .B(n51252), .Z(n51258) );
  XOR U60795 ( .A(n47869), .B(n51258), .Z(n51261) );
  NOR U60796 ( .A(n47871), .B(n47870), .Z(n51260) );
  IV U60797 ( .A(n47872), .Z(n47874) );
  NOR U60798 ( .A(n47874), .B(n47873), .Z(n51264) );
  NOR U60799 ( .A(n51260), .B(n51264), .Z(n47875) );
  XOR U60800 ( .A(n51261), .B(n47875), .Z(n51268) );
  XOR U60801 ( .A(n51267), .B(n51268), .Z(n48249) );
  XOR U60802 ( .A(n48246), .B(n48249), .Z(n47876) );
  XOR U60803 ( .A(n47877), .B(n47876), .Z(n47878) );
  IV U60804 ( .A(n47878), .Z(n51276) );
  XOR U60805 ( .A(n51272), .B(n51276), .Z(n48240) );
  IV U60806 ( .A(n48240), .Z(n47885) );
  IV U60807 ( .A(n47879), .Z(n47881) );
  NOR U60808 ( .A(n47881), .B(n47880), .Z(n51274) );
  NOR U60809 ( .A(n47882), .B(n48241), .Z(n47883) );
  NOR U60810 ( .A(n51274), .B(n47883), .Z(n47884) );
  XOR U60811 ( .A(n47885), .B(n47884), .Z(n48238) );
  IV U60812 ( .A(n47886), .Z(n47888) );
  NOR U60813 ( .A(n47888), .B(n47887), .Z(n47900) );
  IV U60814 ( .A(n47900), .Z(n47889) );
  NOR U60815 ( .A(n48238), .B(n47889), .Z(n51700) );
  IV U60816 ( .A(n47890), .Z(n47892) );
  NOR U60817 ( .A(n47892), .B(n47891), .Z(n47899) );
  IV U60818 ( .A(n47899), .Z(n47896) );
  IV U60819 ( .A(n47893), .Z(n47895) );
  NOR U60820 ( .A(n47895), .B(n47894), .Z(n48236) );
  XOR U60821 ( .A(n48236), .B(n48238), .Z(n47898) );
  NOR U60822 ( .A(n47896), .B(n47898), .Z(n51698) );
  NOR U60823 ( .A(n51700), .B(n51698), .Z(n47897) );
  IV U60824 ( .A(n47897), .Z(n48235) );
  NOR U60825 ( .A(n48235), .B(n47898), .Z(n47903) );
  NOR U60826 ( .A(n47900), .B(n47899), .Z(n47901) );
  NOR U60827 ( .A(n47901), .B(n48235), .Z(n47902) );
  NOR U60828 ( .A(n47903), .B(n47902), .Z(n48233) );
  XOR U60829 ( .A(n48234), .B(n48233), .Z(n47910) );
  IV U60830 ( .A(n47910), .Z(n47904) );
  NOR U60831 ( .A(n47905), .B(n47904), .Z(n54776) );
  IV U60832 ( .A(n47906), .Z(n47908) );
  NOR U60833 ( .A(n47908), .B(n47907), .Z(n47911) );
  IV U60834 ( .A(n47911), .Z(n47909) );
  NOR U60835 ( .A(n47909), .B(n48233), .Z(n54775) );
  NOR U60836 ( .A(n47911), .B(n47910), .Z(n47912) );
  NOR U60837 ( .A(n54775), .B(n47912), .Z(n47913) );
  NOR U60838 ( .A(n47914), .B(n47913), .Z(n47915) );
  NOR U60839 ( .A(n54776), .B(n47915), .Z(n48229) );
  XOR U60840 ( .A(n47916), .B(n48229), .Z(n51298) );
  XOR U60841 ( .A(n47917), .B(n51298), .Z(n48222) );
  XOR U60842 ( .A(n47918), .B(n48222), .Z(n48226) );
  XOR U60843 ( .A(n47919), .B(n48226), .Z(n51309) );
  XOR U60844 ( .A(n51311), .B(n51309), .Z(n51313) );
  XOR U60845 ( .A(n51312), .B(n51313), .Z(n51317) );
  IV U60846 ( .A(n47920), .Z(n47921) );
  NOR U60847 ( .A(n47922), .B(n47921), .Z(n51316) );
  NOR U60848 ( .A(n48217), .B(n51316), .Z(n47923) );
  XOR U60849 ( .A(n51317), .B(n47923), .Z(n47924) );
  IV U60850 ( .A(n47924), .Z(n51320) );
  XOR U60851 ( .A(n51319), .B(n51320), .Z(n47927) );
  NOR U60852 ( .A(n47925), .B(n47927), .Z(n54797) );
  NOR U60853 ( .A(n47926), .B(n48210), .Z(n47928) );
  XOR U60854 ( .A(n47928), .B(n47927), .Z(n48202) );
  IV U60855 ( .A(n48202), .Z(n47929) );
  NOR U60856 ( .A(n47930), .B(n47929), .Z(n47931) );
  NOR U60857 ( .A(n54797), .B(n47931), .Z(n47932) );
  IV U60858 ( .A(n47932), .Z(n48194) );
  IV U60859 ( .A(n47933), .Z(n47934) );
  NOR U60860 ( .A(n47934), .B(n48205), .Z(n48193) );
  XOR U60861 ( .A(n48194), .B(n48193), .Z(n51654) );
  XOR U60862 ( .A(n48191), .B(n51654), .Z(n47935) );
  IV U60863 ( .A(n47935), .Z(n51329) );
  XOR U60864 ( .A(n51326), .B(n51329), .Z(n48189) );
  IV U60865 ( .A(n47936), .Z(n47937) );
  NOR U60866 ( .A(n47938), .B(n47937), .Z(n51328) );
  IV U60867 ( .A(n47939), .Z(n47940) );
  NOR U60868 ( .A(n47941), .B(n47940), .Z(n48188) );
  NOR U60869 ( .A(n51328), .B(n48188), .Z(n47942) );
  XOR U60870 ( .A(n48189), .B(n47942), .Z(n51335) );
  IV U60871 ( .A(n47943), .Z(n47945) );
  NOR U60872 ( .A(n47945), .B(n47944), .Z(n51339) );
  IV U60873 ( .A(n47946), .Z(n47947) );
  NOR U60874 ( .A(n47948), .B(n47947), .Z(n51336) );
  NOR U60875 ( .A(n51339), .B(n51336), .Z(n47949) );
  XOR U60876 ( .A(n51335), .B(n47949), .Z(n51345) );
  IV U60877 ( .A(n47950), .Z(n47951) );
  NOR U60878 ( .A(n47952), .B(n47951), .Z(n48186) );
  IV U60879 ( .A(n47953), .Z(n47954) );
  NOR U60880 ( .A(n47955), .B(n47954), .Z(n51344) );
  NOR U60881 ( .A(n48186), .B(n51344), .Z(n47956) );
  XOR U60882 ( .A(n51345), .B(n47956), .Z(n51347) );
  IV U60883 ( .A(n47957), .Z(n47958) );
  NOR U60884 ( .A(n47959), .B(n47958), .Z(n48183) );
  IV U60885 ( .A(n47960), .Z(n47962) );
  NOR U60886 ( .A(n47962), .B(n47961), .Z(n51348) );
  NOR U60887 ( .A(n48183), .B(n51348), .Z(n47963) );
  XOR U60888 ( .A(n51347), .B(n47963), .Z(n48180) );
  IV U60889 ( .A(n47964), .Z(n47966) );
  NOR U60890 ( .A(n47966), .B(n47965), .Z(n48182) );
  IV U60891 ( .A(n47967), .Z(n47968) );
  NOR U60892 ( .A(n47968), .B(n47972), .Z(n48179) );
  NOR U60893 ( .A(n48182), .B(n48179), .Z(n47969) );
  XOR U60894 ( .A(n48180), .B(n47969), .Z(n48173) );
  IV U60895 ( .A(n47970), .Z(n47971) );
  NOR U60896 ( .A(n47972), .B(n47971), .Z(n48176) );
  IV U60897 ( .A(n47973), .Z(n47974) );
  NOR U60898 ( .A(n47975), .B(n47974), .Z(n48174) );
  NOR U60899 ( .A(n48176), .B(n48174), .Z(n47976) );
  XOR U60900 ( .A(n48173), .B(n47976), .Z(n48171) );
  IV U60901 ( .A(n47977), .Z(n47978) );
  NOR U60902 ( .A(n47979), .B(n47978), .Z(n48170) );
  NOR U60903 ( .A(n47980), .B(n48164), .Z(n47981) );
  NOR U60904 ( .A(n48170), .B(n47981), .Z(n47982) );
  XOR U60905 ( .A(n48171), .B(n47982), .Z(n51355) );
  XOR U60906 ( .A(n47983), .B(n51355), .Z(n51365) );
  IV U60907 ( .A(n47984), .Z(n47986) );
  NOR U60908 ( .A(n47986), .B(n47985), .Z(n51368) );
  IV U60909 ( .A(n47987), .Z(n47989) );
  NOR U60910 ( .A(n47989), .B(n47988), .Z(n51364) );
  NOR U60911 ( .A(n51368), .B(n51364), .Z(n48162) );
  XOR U60912 ( .A(n51365), .B(n48162), .Z(n51375) );
  XOR U60913 ( .A(n47990), .B(n51375), .Z(n51618) );
  XOR U60914 ( .A(n51378), .B(n51618), .Z(n48160) );
  XOR U60915 ( .A(n47991), .B(n48160), .Z(n51392) );
  XOR U60916 ( .A(n47992), .B(n51392), .Z(n51388) );
  XOR U60917 ( .A(n51389), .B(n51388), .Z(n48155) );
  IV U60918 ( .A(n47993), .Z(n47994) );
  NOR U60919 ( .A(n47995), .B(n47994), .Z(n48000) );
  IV U60920 ( .A(n47996), .Z(n47998) );
  NOR U60921 ( .A(n47998), .B(n47997), .Z(n47999) );
  NOR U60922 ( .A(n48000), .B(n47999), .Z(n48156) );
  XOR U60923 ( .A(n48155), .B(n48156), .Z(n51400) );
  XOR U60924 ( .A(n48001), .B(n51400), .Z(n51412) );
  XOR U60925 ( .A(n48002), .B(n51412), .Z(n48150) );
  XOR U60926 ( .A(n48003), .B(n48150), .Z(n48146) );
  XOR U60927 ( .A(n48144), .B(n48146), .Z(n51416) );
  IV U60928 ( .A(n51416), .Z(n48011) );
  IV U60929 ( .A(n48004), .Z(n48005) );
  NOR U60930 ( .A(n48006), .B(n48005), .Z(n48147) );
  IV U60931 ( .A(n48007), .Z(n48009) );
  NOR U60932 ( .A(n48009), .B(n48008), .Z(n51415) );
  NOR U60933 ( .A(n48147), .B(n51415), .Z(n48010) );
  XOR U60934 ( .A(n48011), .B(n48010), .Z(n51420) );
  IV U60935 ( .A(n48012), .Z(n48014) );
  NOR U60936 ( .A(n48014), .B(n48013), .Z(n51418) );
  XOR U60937 ( .A(n51420), .B(n51418), .Z(n51423) );
  XOR U60938 ( .A(n51421), .B(n51423), .Z(n51432) );
  XOR U60939 ( .A(n51431), .B(n51432), .Z(n48015) );
  NOR U60940 ( .A(n48016), .B(n48015), .Z(n51442) );
  NOR U60941 ( .A(n48017), .B(n51427), .Z(n48018) );
  NOR U60942 ( .A(n51431), .B(n48018), .Z(n48019) );
  XOR U60943 ( .A(n48019), .B(n51432), .Z(n51443) );
  NOR U60944 ( .A(n48020), .B(n51443), .Z(n48021) );
  NOR U60945 ( .A(n51442), .B(n48021), .Z(n48140) );
  IV U60946 ( .A(n48022), .Z(n48023) );
  NOR U60947 ( .A(n48023), .B(n48025), .Z(n51444) );
  IV U60948 ( .A(n48024), .Z(n48028) );
  NOR U60949 ( .A(n48026), .B(n48025), .Z(n48027) );
  IV U60950 ( .A(n48027), .Z(n48031) );
  NOR U60951 ( .A(n48028), .B(n48031), .Z(n48141) );
  NOR U60952 ( .A(n51444), .B(n48141), .Z(n48029) );
  XOR U60953 ( .A(n48140), .B(n48029), .Z(n51454) );
  IV U60954 ( .A(n48030), .Z(n48032) );
  NOR U60955 ( .A(n48032), .B(n48031), .Z(n51452) );
  XOR U60956 ( .A(n51454), .B(n51452), .Z(n51456) );
  XOR U60957 ( .A(n51455), .B(n51456), .Z(n51470) );
  XOR U60958 ( .A(n51468), .B(n51470), .Z(n51466) );
  XOR U60959 ( .A(n51464), .B(n51466), .Z(n48133) );
  XOR U60960 ( .A(n48033), .B(n48133), .Z(n48034) );
  IV U60961 ( .A(n48034), .Z(n48131) );
  XOR U60962 ( .A(n48129), .B(n48131), .Z(n48123) );
  NOR U60963 ( .A(n48035), .B(n48126), .Z(n48039) );
  IV U60964 ( .A(n48036), .Z(n48038) );
  IV U60965 ( .A(n48037), .Z(n48042) );
  NOR U60966 ( .A(n48038), .B(n48042), .Z(n48122) );
  NOR U60967 ( .A(n48039), .B(n48122), .Z(n48040) );
  XOR U60968 ( .A(n48123), .B(n48040), .Z(n51487) );
  IV U60969 ( .A(n48041), .Z(n48043) );
  NOR U60970 ( .A(n48043), .B(n48042), .Z(n54891) );
  IV U60971 ( .A(n48044), .Z(n48046) );
  NOR U60972 ( .A(n48046), .B(n48045), .Z(n54896) );
  NOR U60973 ( .A(n54891), .B(n54896), .Z(n51488) );
  XOR U60974 ( .A(n51487), .B(n51488), .Z(n51532) );
  XOR U60975 ( .A(n48047), .B(n51532), .Z(n48120) );
  XOR U60976 ( .A(n48048), .B(n48120), .Z(n48049) );
  IV U60977 ( .A(n48049), .Z(n48116) );
  XOR U60978 ( .A(n48114), .B(n48116), .Z(n51501) );
  XOR U60979 ( .A(n51500), .B(n51501), .Z(n51506) );
  IV U60980 ( .A(n51506), .Z(n48059) );
  IV U60981 ( .A(n48050), .Z(n48051) );
  NOR U60982 ( .A(n48057), .B(n48051), .Z(n48053) );
  IV U60983 ( .A(n48053), .Z(n48052) );
  NOR U60984 ( .A(n48054), .B(n48052), .Z(n51504) );
  XOR U60985 ( .A(n48054), .B(n48053), .Z(n48076) );
  IV U60986 ( .A(n48055), .Z(n48056) );
  NOR U60987 ( .A(n48057), .B(n48056), .Z(n48078) );
  IV U60988 ( .A(n48078), .Z(n48075) );
  NOR U60989 ( .A(n48076), .B(n48075), .Z(n51496) );
  NOR U60990 ( .A(n51504), .B(n51496), .Z(n48058) );
  XOR U60991 ( .A(n48059), .B(n48058), .Z(n48113) );
  XOR U60992 ( .A(n48111), .B(n48113), .Z(n54916) );
  XOR U60993 ( .A(n48061), .B(n48060), .Z(n48086) );
  NOR U60994 ( .A(n48063), .B(n48062), .Z(n48083) );
  XOR U60995 ( .A(n48082), .B(n48083), .Z(n48098) );
  IV U60996 ( .A(n48098), .Z(n48070) );
  IV U60997 ( .A(n48064), .Z(n48066) );
  NOR U60998 ( .A(n48066), .B(n48065), .Z(n54929) );
  IV U60999 ( .A(n54929), .Z(n48067) );
  NOR U61000 ( .A(n48090), .B(n48067), .Z(n54938) );
  IV U61001 ( .A(n54938), .Z(n48068) );
  NOR U61002 ( .A(n48097), .B(n48068), .Z(n48069) );
  IV U61003 ( .A(n48069), .Z(n48099) );
  NOR U61004 ( .A(n48070), .B(n48099), .Z(n54923) );
  IV U61005 ( .A(n54923), .Z(n48071) );
  NOR U61006 ( .A(n48086), .B(n48071), .Z(n48102) );
  IV U61007 ( .A(n48102), .Z(n48072) );
  NOR U61008 ( .A(n48073), .B(n48072), .Z(n48074) );
  IV U61009 ( .A(n48074), .Z(n48110) );
  XOR U61010 ( .A(n48076), .B(n48075), .Z(n48080) );
  NOR U61011 ( .A(n48078), .B(n48077), .Z(n48079) );
  NOR U61012 ( .A(n48080), .B(n48079), .Z(n48081) );
  NOR U61013 ( .A(n48111), .B(n48081), .Z(n48108) );
  XOR U61014 ( .A(n48110), .B(n48108), .Z(n54972) );
  NOR U61015 ( .A(n48083), .B(n48082), .Z(n48087) );
  IV U61016 ( .A(n48087), .Z(n48084) );
  NOR U61017 ( .A(n48085), .B(n48084), .Z(n48089) );
  NOR U61018 ( .A(n48087), .B(n48086), .Z(n48088) );
  NOR U61019 ( .A(n48089), .B(n48088), .Z(n54921) );
  XOR U61020 ( .A(n48091), .B(n48090), .Z(n54928) );
  IV U61021 ( .A(n48092), .Z(n48094) );
  NOR U61022 ( .A(n48094), .B(n48093), .Z(n54944) );
  IV U61023 ( .A(n54944), .Z(n48095) );
  NOR U61024 ( .A(n54928), .B(n48095), .Z(n54937) );
  IV U61025 ( .A(n54937), .Z(n48096) );
  NOR U61026 ( .A(n48097), .B(n48096), .Z(n54927) );
  IV U61027 ( .A(n54927), .Z(n48100) );
  XOR U61028 ( .A(n48099), .B(n48098), .Z(n54926) );
  NOR U61029 ( .A(n48100), .B(n54926), .Z(n54922) );
  IV U61030 ( .A(n54922), .Z(n48101) );
  NOR U61031 ( .A(n54921), .B(n48101), .Z(n54919) );
  IV U61032 ( .A(n54919), .Z(n48106) );
  NOR U61033 ( .A(n48103), .B(n48102), .Z(n48105) );
  XOR U61034 ( .A(n48105), .B(n48104), .Z(n54918) );
  NOR U61035 ( .A(n48106), .B(n54918), .Z(n54970) );
  IV U61036 ( .A(n54970), .Z(n48107) );
  NOR U61037 ( .A(n54972), .B(n48107), .Z(n54913) );
  IV U61038 ( .A(n48108), .Z(n48109) );
  NOR U61039 ( .A(n48110), .B(n48109), .Z(n54914) );
  IV U61040 ( .A(n48111), .Z(n48112) );
  NOR U61041 ( .A(n48113), .B(n48112), .Z(n51514) );
  IV U61042 ( .A(n48114), .Z(n48115) );
  NOR U61043 ( .A(n48116), .B(n48115), .Z(n51524) );
  IV U61044 ( .A(n48117), .Z(n48118) );
  NOR U61045 ( .A(n48118), .B(n48120), .Z(n54905) );
  IV U61046 ( .A(n48119), .Z(n48121) );
  NOR U61047 ( .A(n48121), .B(n48120), .Z(n54902) );
  IV U61048 ( .A(n48122), .Z(n48124) );
  NOR U61049 ( .A(n48124), .B(n48123), .Z(n51538) );
  IV U61050 ( .A(n48125), .Z(n48128) );
  NOR U61051 ( .A(n48131), .B(n48126), .Z(n48127) );
  IV U61052 ( .A(n48127), .Z(n51485) );
  NOR U61053 ( .A(n48128), .B(n51485), .Z(n54876) );
  IV U61054 ( .A(n48129), .Z(n48130) );
  NOR U61055 ( .A(n48131), .B(n48130), .Z(n54880) );
  IV U61056 ( .A(n48132), .Z(n48134) );
  NOR U61057 ( .A(n48134), .B(n48133), .Z(n54883) );
  NOR U61058 ( .A(n54880), .B(n54883), .Z(n51482) );
  IV U61059 ( .A(n48135), .Z(n48138) );
  NOR U61060 ( .A(n48136), .B(n51470), .Z(n48137) );
  IV U61061 ( .A(n48137), .Z(n51460) );
  NOR U61062 ( .A(n48138), .B(n51460), .Z(n48139) );
  IV U61063 ( .A(n48139), .Z(n54874) );
  IV U61064 ( .A(n48140), .Z(n48143) );
  IV U61065 ( .A(n48141), .Z(n48142) );
  NOR U61066 ( .A(n48143), .B(n48142), .Z(n51450) );
  IV U61067 ( .A(n51450), .Z(n51441) );
  IV U61068 ( .A(n48144), .Z(n48145) );
  NOR U61069 ( .A(n48146), .B(n48145), .Z(n51567) );
  IV U61070 ( .A(n48147), .Z(n48148) );
  NOR U61071 ( .A(n48148), .B(n51416), .Z(n51565) );
  NOR U61072 ( .A(n51567), .B(n51565), .Z(n51413) );
  IV U61073 ( .A(n48149), .Z(n48151) );
  IV U61074 ( .A(n48150), .Z(n48153) );
  NOR U61075 ( .A(n48151), .B(n48153), .Z(n51573) );
  IV U61076 ( .A(n48152), .Z(n48154) );
  NOR U61077 ( .A(n48154), .B(n48153), .Z(n51570) );
  NOR U61078 ( .A(n48156), .B(n48155), .Z(n51395) );
  IV U61079 ( .A(n48157), .Z(n48158) );
  NOR U61080 ( .A(n51392), .B(n48158), .Z(n51608) );
  IV U61081 ( .A(n48159), .Z(n48161) );
  IV U61082 ( .A(n48160), .Z(n51386) );
  NOR U61083 ( .A(n48161), .B(n51386), .Z(n51605) );
  NOR U61084 ( .A(n48162), .B(n51365), .Z(n51363) );
  IV U61085 ( .A(n48163), .Z(n48166) );
  NOR U61086 ( .A(n48164), .B(n48171), .Z(n48165) );
  IV U61087 ( .A(n48165), .Z(n48168) );
  NOR U61088 ( .A(n48166), .B(n48168), .Z(n51629) );
  IV U61089 ( .A(n48167), .Z(n48169) );
  NOR U61090 ( .A(n48169), .B(n48168), .Z(n51636) );
  IV U61091 ( .A(n48170), .Z(n48172) );
  NOR U61092 ( .A(n48172), .B(n48171), .Z(n51633) );
  IV U61093 ( .A(n48173), .Z(n48178) );
  IV U61094 ( .A(n48174), .Z(n48175) );
  NOR U61095 ( .A(n48178), .B(n48175), .Z(n54826) );
  IV U61096 ( .A(n48176), .Z(n48177) );
  NOR U61097 ( .A(n48178), .B(n48177), .Z(n54823) );
  IV U61098 ( .A(n48179), .Z(n48181) );
  NOR U61099 ( .A(n48181), .B(n48180), .Z(n54818) );
  IV U61100 ( .A(n48182), .Z(n48185) );
  IV U61101 ( .A(n48183), .Z(n51350) );
  XOR U61102 ( .A(n51350), .B(n51347), .Z(n48184) );
  NOR U61103 ( .A(n48185), .B(n48184), .Z(n54815) );
  IV U61104 ( .A(n48186), .Z(n48187) );
  NOR U61105 ( .A(n48187), .B(n51345), .Z(n54802) );
  IV U61106 ( .A(n48188), .Z(n48190) );
  NOR U61107 ( .A(n48190), .B(n48189), .Z(n51332) );
  IV U61108 ( .A(n51332), .Z(n51325) );
  NOR U61109 ( .A(n48191), .B(n51654), .Z(n48199) );
  IV U61110 ( .A(n48192), .Z(n48198) );
  IV U61111 ( .A(n48193), .Z(n48195) );
  NOR U61112 ( .A(n48195), .B(n48194), .Z(n48196) );
  IV U61113 ( .A(n48196), .Z(n48197) );
  NOR U61114 ( .A(n48198), .B(n48197), .Z(n51649) );
  NOR U61115 ( .A(n48199), .B(n51649), .Z(n51324) );
  IV U61116 ( .A(n48200), .Z(n48201) );
  NOR U61117 ( .A(n48202), .B(n48201), .Z(n48203) );
  IV U61118 ( .A(n48203), .Z(n48208) );
  NOR U61119 ( .A(n48205), .B(n48204), .Z(n48206) );
  IV U61120 ( .A(n48206), .Z(n48207) );
  NOR U61121 ( .A(n48208), .B(n48207), .Z(n51662) );
  NOR U61122 ( .A(n54797), .B(n51662), .Z(n51323) );
  IV U61123 ( .A(n48209), .Z(n48212) );
  NOR U61124 ( .A(n48210), .B(n51320), .Z(n48211) );
  IV U61125 ( .A(n48211), .Z(n48214) );
  NOR U61126 ( .A(n48212), .B(n48214), .Z(n54795) );
  IV U61127 ( .A(n54795), .Z(n54793) );
  IV U61128 ( .A(n48213), .Z(n48215) );
  NOR U61129 ( .A(n48215), .B(n48214), .Z(n48216) );
  IV U61130 ( .A(n48216), .Z(n51665) );
  IV U61131 ( .A(n48217), .Z(n48218) );
  NOR U61132 ( .A(n48218), .B(n51317), .Z(n51673) );
  IV U61133 ( .A(n48219), .Z(n48220) );
  NOR U61134 ( .A(n48226), .B(n48220), .Z(n51684) );
  IV U61135 ( .A(n48221), .Z(n48223) );
  IV U61136 ( .A(n48222), .Z(n51304) );
  NOR U61137 ( .A(n48223), .B(n51304), .Z(n51687) );
  NOR U61138 ( .A(n51684), .B(n51687), .Z(n51308) );
  IV U61139 ( .A(n48224), .Z(n48225) );
  NOR U61140 ( .A(n48226), .B(n48225), .Z(n48227) );
  IV U61141 ( .A(n48227), .Z(n51683) );
  IV U61142 ( .A(n48228), .Z(n48230) );
  IV U61143 ( .A(n48229), .Z(n51289) );
  NOR U61144 ( .A(n48230), .B(n51289), .Z(n54785) );
  IV U61145 ( .A(n48231), .Z(n48232) );
  NOR U61146 ( .A(n48232), .B(n51289), .Z(n51694) );
  NOR U61147 ( .A(n54776), .B(n51694), .Z(n51285) );
  IV U61148 ( .A(n54775), .Z(n54773) );
  NOR U61149 ( .A(n48234), .B(n48233), .Z(n51697) );
  NOR U61150 ( .A(n48235), .B(n51697), .Z(n51284) );
  IV U61151 ( .A(n48236), .Z(n48237) );
  NOR U61152 ( .A(n48238), .B(n48237), .Z(n51703) );
  IV U61153 ( .A(n48239), .Z(n48243) );
  NOR U61154 ( .A(n48241), .B(n48240), .Z(n48242) );
  IV U61155 ( .A(n48242), .Z(n51280) );
  NOR U61156 ( .A(n48243), .B(n51280), .Z(n51706) );
  NOR U61157 ( .A(n51703), .B(n51706), .Z(n51282) );
  IV U61158 ( .A(n48244), .Z(n48245) );
  NOR U61159 ( .A(n48245), .B(n48249), .Z(n54765) );
  IV U61160 ( .A(n48246), .Z(n48247) );
  NOR U61161 ( .A(n48247), .B(n48249), .Z(n51717) );
  IV U61162 ( .A(n48248), .Z(n48250) );
  NOR U61163 ( .A(n48250), .B(n48249), .Z(n51714) );
  NOR U61164 ( .A(n51717), .B(n51714), .Z(n51271) );
  IV U61165 ( .A(n48251), .Z(n51241) );
  IV U61166 ( .A(n48252), .Z(n48253) );
  NOR U61167 ( .A(n51241), .B(n48253), .Z(n48254) );
  IV U61168 ( .A(n48254), .Z(n51246) );
  IV U61169 ( .A(n48255), .Z(n48257) );
  NOR U61170 ( .A(n48257), .B(n48256), .Z(n54746) );
  IV U61171 ( .A(n48258), .Z(n48259) );
  NOR U61172 ( .A(n48259), .B(n51244), .Z(n51738) );
  NOR U61173 ( .A(n54746), .B(n51738), .Z(n51238) );
  IV U61174 ( .A(n48260), .Z(n48261) );
  NOR U61175 ( .A(n48262), .B(n48261), .Z(n51740) );
  IV U61176 ( .A(n48263), .Z(n48265) );
  NOR U61177 ( .A(n48265), .B(n48264), .Z(n51747) );
  NOR U61178 ( .A(n51740), .B(n51747), .Z(n51237) );
  IV U61179 ( .A(n48266), .Z(n48269) );
  NOR U61180 ( .A(n48267), .B(n51226), .Z(n48268) );
  IV U61181 ( .A(n48268), .Z(n51234) );
  NOR U61182 ( .A(n48269), .B(n51234), .Z(n51743) );
  IV U61183 ( .A(n51743), .Z(n51746) );
  IV U61184 ( .A(n48270), .Z(n48271) );
  NOR U61185 ( .A(n48272), .B(n48271), .Z(n51764) );
  IV U61186 ( .A(n48273), .Z(n48274) );
  NOR U61187 ( .A(n48274), .B(n48276), .Z(n54739) );
  IV U61188 ( .A(n48275), .Z(n48277) );
  NOR U61189 ( .A(n48277), .B(n48276), .Z(n54736) );
  IV U61190 ( .A(n48278), .Z(n48279) );
  NOR U61191 ( .A(n48280), .B(n48279), .Z(n48281) );
  IV U61192 ( .A(n48281), .Z(n51786) );
  NOR U61193 ( .A(n48283), .B(n48282), .Z(n54706) );
  IV U61194 ( .A(n48284), .Z(n48285) );
  NOR U61195 ( .A(n48286), .B(n48285), .Z(n51790) );
  NOR U61196 ( .A(n51790), .B(n54708), .Z(n51173) );
  IV U61197 ( .A(n48287), .Z(n48290) );
  IV U61198 ( .A(n48288), .Z(n48289) );
  NOR U61199 ( .A(n48290), .B(n48289), .Z(n54702) );
  IV U61200 ( .A(n48291), .Z(n48292) );
  NOR U61201 ( .A(n48292), .B(n51169), .Z(n54699) );
  IV U61202 ( .A(n48293), .Z(n48294) );
  NOR U61203 ( .A(n51168), .B(n48294), .Z(n54691) );
  IV U61204 ( .A(n48295), .Z(n48297) );
  IV U61205 ( .A(n48296), .Z(n48300) );
  NOR U61206 ( .A(n48297), .B(n48300), .Z(n51795) );
  NOR U61207 ( .A(n51799), .B(n48298), .Z(n48302) );
  IV U61208 ( .A(n48299), .Z(n48301) );
  NOR U61209 ( .A(n48301), .B(n48300), .Z(n54688) );
  NOR U61210 ( .A(n48302), .B(n54688), .Z(n51164) );
  IV U61211 ( .A(n48303), .Z(n48306) );
  IV U61212 ( .A(n48304), .Z(n48305) );
  NOR U61213 ( .A(n48306), .B(n48305), .Z(n51808) );
  NOR U61214 ( .A(n48308), .B(n48307), .Z(n51822) );
  IV U61215 ( .A(n48309), .Z(n54664) );
  IV U61216 ( .A(n48310), .Z(n48311) );
  NOR U61217 ( .A(n54664), .B(n48311), .Z(n51824) );
  NOR U61218 ( .A(n51822), .B(n51824), .Z(n51152) );
  NOR U61219 ( .A(n54680), .B(n51827), .Z(n48313) );
  NOR U61220 ( .A(n48313), .B(n48312), .Z(n51151) );
  NOR U61221 ( .A(n48314), .B(n54653), .Z(n48315) );
  IV U61222 ( .A(n48315), .Z(n51832) );
  IV U61223 ( .A(n48316), .Z(n48319) );
  IV U61224 ( .A(n48317), .Z(n48318) );
  NOR U61225 ( .A(n48319), .B(n48318), .Z(n51147) );
  IV U61226 ( .A(n48320), .Z(n48322) );
  NOR U61227 ( .A(n48322), .B(n48321), .Z(n48323) );
  NOR U61228 ( .A(n48324), .B(n48323), .Z(n54651) );
  NOR U61229 ( .A(n48326), .B(n48325), .Z(n54646) );
  IV U61230 ( .A(n48327), .Z(n48328) );
  NOR U61231 ( .A(n48329), .B(n48328), .Z(n51836) );
  IV U61232 ( .A(n48330), .Z(n48335) );
  IV U61233 ( .A(n48331), .Z(n48332) );
  NOR U61234 ( .A(n48335), .B(n48332), .Z(n51838) );
  NOR U61235 ( .A(n51836), .B(n51838), .Z(n51146) );
  IV U61236 ( .A(n48333), .Z(n48334) );
  NOR U61237 ( .A(n48335), .B(n48334), .Z(n51842) );
  NOR U61238 ( .A(n48336), .B(n51143), .Z(n51844) );
  NOR U61239 ( .A(n51842), .B(n51844), .Z(n51145) );
  IV U61240 ( .A(n48337), .Z(n48338) );
  NOR U61241 ( .A(n48338), .B(n51143), .Z(n51851) );
  NOR U61242 ( .A(n48339), .B(n51858), .Z(n48342) );
  IV U61243 ( .A(n48340), .Z(n48341) );
  NOR U61244 ( .A(n48341), .B(n48344), .Z(n54639) );
  NOR U61245 ( .A(n48342), .B(n54639), .Z(n51141) );
  IV U61246 ( .A(n48343), .Z(n48345) );
  NOR U61247 ( .A(n48345), .B(n48344), .Z(n48346) );
  IV U61248 ( .A(n48346), .Z(n51856) );
  IV U61249 ( .A(n48347), .Z(n48349) );
  NOR U61250 ( .A(n48349), .B(n48348), .Z(n48354) );
  IV U61251 ( .A(n48350), .Z(n48351) );
  NOR U61252 ( .A(n48352), .B(n48351), .Z(n48353) );
  NOR U61253 ( .A(n48354), .B(n48353), .Z(n54626) );
  NOR U61254 ( .A(n48356), .B(n48355), .Z(n54627) );
  IV U61255 ( .A(n48357), .Z(n48358) );
  NOR U61256 ( .A(n48358), .B(n48360), .Z(n54615) );
  IV U61257 ( .A(n48359), .Z(n48361) );
  NOR U61258 ( .A(n48361), .B(n48360), .Z(n51124) );
  IV U61259 ( .A(n51124), .Z(n51110) );
  IV U61260 ( .A(n48362), .Z(n48363) );
  NOR U61261 ( .A(n48363), .B(n51107), .Z(n48364) );
  IV U61262 ( .A(n48364), .Z(n54606) );
  IV U61263 ( .A(n48365), .Z(n48367) );
  NOR U61264 ( .A(n48367), .B(n48366), .Z(n51868) );
  IV U61265 ( .A(n48368), .Z(n48369) );
  NOR U61266 ( .A(n48369), .B(n51104), .Z(n51866) );
  NOR U61267 ( .A(n51868), .B(n51866), .Z(n51098) );
  IV U61268 ( .A(n48370), .Z(n48371) );
  NOR U61269 ( .A(n48371), .B(n51873), .Z(n51871) );
  NOR U61270 ( .A(n54595), .B(n51871), .Z(n51097) );
  IV U61271 ( .A(n48372), .Z(n48374) );
  NOR U61272 ( .A(n48374), .B(n48373), .Z(n51893) );
  NOR U61273 ( .A(n48375), .B(n51887), .Z(n48376) );
  NOR U61274 ( .A(n51893), .B(n48376), .Z(n51096) );
  IV U61275 ( .A(n48377), .Z(n48378) );
  NOR U61276 ( .A(n48378), .B(n51085), .Z(n51900) );
  IV U61277 ( .A(n48379), .Z(n48380) );
  NOR U61278 ( .A(n48381), .B(n48380), .Z(n48382) );
  IV U61279 ( .A(n48382), .Z(n51078) );
  IV U61280 ( .A(n48383), .Z(n48384) );
  NOR U61281 ( .A(n48384), .B(n48386), .Z(n51923) );
  IV U61282 ( .A(n48385), .Z(n48387) );
  NOR U61283 ( .A(n48387), .B(n48386), .Z(n51917) );
  IV U61284 ( .A(n48388), .Z(n48391) );
  NOR U61285 ( .A(n48389), .B(n51061), .Z(n48390) );
  IV U61286 ( .A(n48390), .Z(n51067) );
  NOR U61287 ( .A(n48391), .B(n51067), .Z(n51914) );
  IV U61288 ( .A(n48392), .Z(n48394) );
  IV U61289 ( .A(n48393), .Z(n48398) );
  NOR U61290 ( .A(n48394), .B(n48398), .Z(n54548) );
  IV U61291 ( .A(n48395), .Z(n48396) );
  NOR U61292 ( .A(n48396), .B(n48402), .Z(n51943) );
  IV U61293 ( .A(n48397), .Z(n48399) );
  NOR U61294 ( .A(n48399), .B(n48398), .Z(n54551) );
  NOR U61295 ( .A(n51943), .B(n54551), .Z(n51046) );
  IV U61296 ( .A(n48400), .Z(n48401) );
  NOR U61297 ( .A(n48402), .B(n48401), .Z(n51041) );
  IV U61298 ( .A(n48403), .Z(n48405) );
  NOR U61299 ( .A(n48405), .B(n48404), .Z(n48406) );
  IV U61300 ( .A(n48406), .Z(n51949) );
  IV U61301 ( .A(n48407), .Z(n48410) );
  NOR U61302 ( .A(n48408), .B(n48413), .Z(n48409) );
  IV U61303 ( .A(n48409), .Z(n51030) );
  NOR U61304 ( .A(n48410), .B(n51030), .Z(n51022) );
  IV U61305 ( .A(n48411), .Z(n48412) );
  NOR U61306 ( .A(n48413), .B(n48412), .Z(n51019) );
  IV U61307 ( .A(n51019), .Z(n51014) );
  IV U61308 ( .A(n48414), .Z(n48420) );
  IV U61309 ( .A(n48415), .Z(n48416) );
  NOR U61310 ( .A(n48420), .B(n48416), .Z(n54535) );
  NOR U61311 ( .A(n48418), .B(n48417), .Z(n54528) );
  IV U61312 ( .A(n48419), .Z(n48421) );
  NOR U61313 ( .A(n48421), .B(n48420), .Z(n51960) );
  NOR U61314 ( .A(n54528), .B(n51960), .Z(n51012) );
  IV U61315 ( .A(n48422), .Z(n51964) );
  NOR U61316 ( .A(n48423), .B(n51964), .Z(n51011) );
  XOR U61317 ( .A(n50995), .B(n50996), .Z(n48425) );
  NOR U61318 ( .A(n48425), .B(n48424), .Z(n51980) );
  IV U61319 ( .A(n48426), .Z(n48427) );
  NOR U61320 ( .A(n50987), .B(n48427), .Z(n51996) );
  IV U61321 ( .A(n48428), .Z(n48431) );
  IV U61322 ( .A(n48429), .Z(n48430) );
  NOR U61323 ( .A(n48431), .B(n48430), .Z(n52003) );
  NOR U61324 ( .A(n51996), .B(n52003), .Z(n50983) );
  NOR U61325 ( .A(n48433), .B(n48432), .Z(n48434) );
  IV U61326 ( .A(n48434), .Z(n48435) );
  NOR U61327 ( .A(n48435), .B(n52013), .Z(n52007) );
  IV U61328 ( .A(n48436), .Z(n48437) );
  NOR U61329 ( .A(n48439), .B(n48437), .Z(n52020) );
  IV U61330 ( .A(n48438), .Z(n48443) );
  NOR U61331 ( .A(n48440), .B(n48439), .Z(n48441) );
  IV U61332 ( .A(n48441), .Z(n48442) );
  NOR U61333 ( .A(n48443), .B(n48442), .Z(n54521) );
  NOR U61334 ( .A(n52020), .B(n54521), .Z(n50975) );
  NOR U61335 ( .A(n48445), .B(n48444), .Z(n48450) );
  IV U61336 ( .A(n48446), .Z(n48447) );
  NOR U61337 ( .A(n48448), .B(n48447), .Z(n48449) );
  NOR U61338 ( .A(n48450), .B(n48449), .Z(n52024) );
  IV U61339 ( .A(n48451), .Z(n48453) );
  NOR U61340 ( .A(n48453), .B(n48452), .Z(n50968) );
  IV U61341 ( .A(n50968), .Z(n50963) );
  IV U61342 ( .A(n48454), .Z(n48455) );
  NOR U61343 ( .A(n48455), .B(n48461), .Z(n52047) );
  IV U61344 ( .A(n48456), .Z(n48457) );
  NOR U61345 ( .A(n48458), .B(n48457), .Z(n52059) );
  IV U61346 ( .A(n48459), .Z(n48460) );
  NOR U61347 ( .A(n48461), .B(n48460), .Z(n52060) );
  NOR U61348 ( .A(n52059), .B(n52060), .Z(n58217) );
  IV U61349 ( .A(n48462), .Z(n48464) );
  NOR U61350 ( .A(n48464), .B(n48463), .Z(n54486) );
  IV U61351 ( .A(n48465), .Z(n48468) );
  IV U61352 ( .A(n48466), .Z(n48467) );
  NOR U61353 ( .A(n48468), .B(n48467), .Z(n52073) );
  NOR U61354 ( .A(n54486), .B(n52073), .Z(n50908) );
  IV U61355 ( .A(n48469), .Z(n48470) );
  NOR U61356 ( .A(n48471), .B(n48470), .Z(n52083) );
  NOR U61357 ( .A(n48473), .B(n48472), .Z(n52089) );
  IV U61358 ( .A(n48474), .Z(n48478) );
  IV U61359 ( .A(n48475), .Z(n48483) );
  NOR U61360 ( .A(n48476), .B(n48483), .Z(n48477) );
  IV U61361 ( .A(n48477), .Z(n50903) );
  NOR U61362 ( .A(n48478), .B(n50903), .Z(n48479) );
  IV U61363 ( .A(n48479), .Z(n52111) );
  IV U61364 ( .A(n48480), .Z(n48481) );
  NOR U61365 ( .A(n48481), .B(n48488), .Z(n54478) );
  IV U61366 ( .A(n48482), .Z(n48486) );
  NOR U61367 ( .A(n48484), .B(n48483), .Z(n48485) );
  IV U61368 ( .A(n48485), .Z(n50895) );
  NOR U61369 ( .A(n48486), .B(n50895), .Z(n52112) );
  NOR U61370 ( .A(n54478), .B(n52112), .Z(n50893) );
  IV U61371 ( .A(n48487), .Z(n48489) );
  NOR U61372 ( .A(n48489), .B(n48488), .Z(n54479) );
  IV U61373 ( .A(n48490), .Z(n48495) );
  IV U61374 ( .A(n48491), .Z(n48492) );
  NOR U61375 ( .A(n48495), .B(n48492), .Z(n54469) );
  IV U61376 ( .A(n48493), .Z(n48494) );
  NOR U61377 ( .A(n48495), .B(n48494), .Z(n54473) );
  IV U61378 ( .A(n48496), .Z(n48498) );
  NOR U61379 ( .A(n48498), .B(n48497), .Z(n52115) );
  NOR U61380 ( .A(n54473), .B(n52115), .Z(n50891) );
  IV U61381 ( .A(n48499), .Z(n48500) );
  NOR U61382 ( .A(n48500), .B(n50884), .Z(n50889) );
  IV U61383 ( .A(n48501), .Z(n48503) );
  NOR U61384 ( .A(n48503), .B(n48502), .Z(n54464) );
  IV U61385 ( .A(n48504), .Z(n48505) );
  NOR U61386 ( .A(n48505), .B(n48507), .Z(n54461) );
  IV U61387 ( .A(n48506), .Z(n48508) );
  NOR U61388 ( .A(n48508), .B(n48507), .Z(n52123) );
  IV U61389 ( .A(n48509), .Z(n48510) );
  NOR U61390 ( .A(n48510), .B(n50865), .Z(n52132) );
  IV U61391 ( .A(n48511), .Z(n48512) );
  NOR U61392 ( .A(n50858), .B(n48512), .Z(n52152) );
  IV U61393 ( .A(n48513), .Z(n48515) );
  NOR U61394 ( .A(n48515), .B(n48514), .Z(n52149) );
  IV U61395 ( .A(n48516), .Z(n48517) );
  NOR U61396 ( .A(n48520), .B(n48517), .Z(n52160) );
  IV U61397 ( .A(n48518), .Z(n48519) );
  NOR U61398 ( .A(n48520), .B(n48519), .Z(n54443) );
  NOR U61399 ( .A(n52160), .B(n54443), .Z(n50854) );
  IV U61400 ( .A(n48521), .Z(n48523) );
  NOR U61401 ( .A(n48523), .B(n48522), .Z(n54430) );
  IV U61402 ( .A(n48524), .Z(n48525) );
  NOR U61403 ( .A(n48525), .B(n48528), .Z(n48526) );
  IV U61404 ( .A(n48526), .Z(n54436) );
  IV U61405 ( .A(n48527), .Z(n48529) );
  NOR U61406 ( .A(n48529), .B(n48528), .Z(n48530) );
  IV U61407 ( .A(n48530), .Z(n54435) );
  XOR U61408 ( .A(n54436), .B(n54435), .Z(n48531) );
  NOR U61409 ( .A(n54430), .B(n48531), .Z(n50853) );
  IV U61410 ( .A(n48532), .Z(n48534) );
  NOR U61411 ( .A(n48534), .B(n48533), .Z(n52166) );
  NOR U61412 ( .A(n48535), .B(n52166), .Z(n50852) );
  IV U61413 ( .A(n48536), .Z(n48537) );
  NOR U61414 ( .A(n48537), .B(n48540), .Z(n54418) );
  IV U61415 ( .A(n48538), .Z(n48539) );
  NOR U61416 ( .A(n48540), .B(n48539), .Z(n54422) );
  IV U61417 ( .A(n48541), .Z(n52169) );
  IV U61418 ( .A(n48542), .Z(n48543) );
  NOR U61419 ( .A(n52169), .B(n48543), .Z(n48544) );
  NOR U61420 ( .A(n54422), .B(n48544), .Z(n50851) );
  IV U61421 ( .A(n48545), .Z(n48546) );
  NOR U61422 ( .A(n48552), .B(n48546), .Z(n52180) );
  IV U61423 ( .A(n48547), .Z(n48548) );
  NOR U61424 ( .A(n48548), .B(n52169), .Z(n48549) );
  NOR U61425 ( .A(n52180), .B(n48549), .Z(n50850) );
  IV U61426 ( .A(n48550), .Z(n48551) );
  NOR U61427 ( .A(n48552), .B(n48551), .Z(n52174) );
  IV U61428 ( .A(n48553), .Z(n48555) );
  IV U61429 ( .A(n48554), .Z(n48558) );
  NOR U61430 ( .A(n48555), .B(n48558), .Z(n52176) );
  NOR U61431 ( .A(n52174), .B(n52176), .Z(n50849) );
  NOR U61432 ( .A(n48556), .B(n52189), .Z(n48560) );
  IV U61433 ( .A(n48557), .Z(n48559) );
  NOR U61434 ( .A(n48559), .B(n48558), .Z(n52184) );
  NOR U61435 ( .A(n48560), .B(n52184), .Z(n50848) );
  IV U61436 ( .A(n48561), .Z(n48563) );
  NOR U61437 ( .A(n48563), .B(n48562), .Z(n48564) );
  IV U61438 ( .A(n48564), .Z(n54409) );
  IV U61439 ( .A(n48565), .Z(n48566) );
  NOR U61440 ( .A(n48567), .B(n48566), .Z(n52193) );
  IV U61441 ( .A(n48568), .Z(n48570) );
  IV U61442 ( .A(n48569), .Z(n48572) );
  NOR U61443 ( .A(n48570), .B(n48572), .Z(n52195) );
  NOR U61444 ( .A(n52193), .B(n52195), .Z(n50847) );
  IV U61445 ( .A(n48571), .Z(n48573) );
  NOR U61446 ( .A(n48573), .B(n48572), .Z(n52200) );
  NOR U61447 ( .A(n52204), .B(n52200), .Z(n50846) );
  NOR U61448 ( .A(n48575), .B(n48574), .Z(n52216) );
  IV U61449 ( .A(n48576), .Z(n48578) );
  NOR U61450 ( .A(n48578), .B(n48577), .Z(n52209) );
  NOR U61451 ( .A(n52216), .B(n52209), .Z(n50839) );
  IV U61452 ( .A(n52212), .Z(n52214) );
  IV U61453 ( .A(n48579), .Z(n48580) );
  NOR U61454 ( .A(n48581), .B(n48580), .Z(n55828) );
  IV U61455 ( .A(n48582), .Z(n48584) );
  NOR U61456 ( .A(n48584), .B(n48583), .Z(n55842) );
  NOR U61457 ( .A(n55828), .B(n55842), .Z(n52228) );
  IV U61458 ( .A(n48585), .Z(n48586) );
  NOR U61459 ( .A(n48591), .B(n48586), .Z(n48587) );
  IV U61460 ( .A(n48587), .Z(n52231) );
  IV U61461 ( .A(n48588), .Z(n48590) );
  NOR U61462 ( .A(n48590), .B(n48589), .Z(n52237) );
  NOR U61463 ( .A(n48592), .B(n48591), .Z(n48593) );
  IV U61464 ( .A(n48593), .Z(n48594) );
  NOR U61465 ( .A(n48595), .B(n48594), .Z(n52232) );
  NOR U61466 ( .A(n52237), .B(n52232), .Z(n50836) );
  IV U61467 ( .A(n48596), .Z(n48598) );
  NOR U61468 ( .A(n48598), .B(n48597), .Z(n52238) );
  NOR U61469 ( .A(n55806), .B(n52238), .Z(n50835) );
  IV U61470 ( .A(n48599), .Z(n48600) );
  NOR U61471 ( .A(n48600), .B(n50829), .Z(n48601) );
  IV U61472 ( .A(n48601), .Z(n48602) );
  NOR U61473 ( .A(n48603), .B(n48602), .Z(n48604) );
  IV U61474 ( .A(n48604), .Z(n52244) );
  IV U61475 ( .A(n48605), .Z(n48606) );
  NOR U61476 ( .A(n48606), .B(n48611), .Z(n52249) );
  IV U61477 ( .A(n48607), .Z(n48609) );
  NOR U61478 ( .A(n48609), .B(n48608), .Z(n52247) );
  NOR U61479 ( .A(n52249), .B(n52247), .Z(n50824) );
  IV U61480 ( .A(n48610), .Z(n48612) );
  NOR U61481 ( .A(n48612), .B(n48611), .Z(n52252) );
  IV U61482 ( .A(n48613), .Z(n48618) );
  IV U61483 ( .A(n48614), .Z(n48615) );
  NOR U61484 ( .A(n48618), .B(n48615), .Z(n52254) );
  NOR U61485 ( .A(n52252), .B(n52254), .Z(n50823) );
  IV U61486 ( .A(n48616), .Z(n48617) );
  NOR U61487 ( .A(n48618), .B(n48617), .Z(n52260) );
  IV U61488 ( .A(n48619), .Z(n48621) );
  IV U61489 ( .A(n48620), .Z(n48630) );
  NOR U61490 ( .A(n48621), .B(n48630), .Z(n48628) );
  IV U61491 ( .A(n48622), .Z(n48626) );
  NOR U61492 ( .A(n48624), .B(n48623), .Z(n48625) );
  IV U61493 ( .A(n48625), .Z(n50806) );
  NOR U61494 ( .A(n48626), .B(n50806), .Z(n48627) );
  NOR U61495 ( .A(n48628), .B(n48627), .Z(n52283) );
  IV U61496 ( .A(n48629), .Z(n48631) );
  NOR U61497 ( .A(n48631), .B(n48630), .Z(n54370) );
  IV U61498 ( .A(n48632), .Z(n48633) );
  NOR U61499 ( .A(n48636), .B(n48633), .Z(n54373) );
  IV U61500 ( .A(n48634), .Z(n48635) );
  NOR U61501 ( .A(n48636), .B(n48635), .Z(n52284) );
  IV U61502 ( .A(n48637), .Z(n48639) );
  IV U61503 ( .A(n48638), .Z(n48641) );
  NOR U61504 ( .A(n48639), .B(n48641), .Z(n52290) );
  IV U61505 ( .A(n48640), .Z(n48642) );
  NOR U61506 ( .A(n48642), .B(n48641), .Z(n52287) );
  IV U61507 ( .A(n48643), .Z(n48644) );
  NOR U61508 ( .A(n48644), .B(n50803), .Z(n54360) );
  IV U61509 ( .A(n48645), .Z(n48646) );
  NOR U61510 ( .A(n48650), .B(n48646), .Z(n48647) );
  IV U61511 ( .A(n48647), .Z(n54352) );
  IV U61512 ( .A(n48648), .Z(n48649) );
  NOR U61513 ( .A(n48650), .B(n48649), .Z(n54349) );
  IV U61514 ( .A(n48651), .Z(n48652) );
  NOR U61515 ( .A(n48652), .B(n48655), .Z(n48653) );
  IV U61516 ( .A(n48653), .Z(n52297) );
  IV U61517 ( .A(n48654), .Z(n48656) );
  NOR U61518 ( .A(n48656), .B(n48655), .Z(n48663) );
  IV U61519 ( .A(n48657), .Z(n48661) );
  IV U61520 ( .A(n48658), .Z(n48669) );
  NOR U61521 ( .A(n48669), .B(n48659), .Z(n48660) );
  IV U61522 ( .A(n48660), .Z(n48665) );
  NOR U61523 ( .A(n48661), .B(n48665), .Z(n48662) );
  NOR U61524 ( .A(n48663), .B(n48662), .Z(n52302) );
  IV U61525 ( .A(n48664), .Z(n48666) );
  NOR U61526 ( .A(n48666), .B(n48665), .Z(n52298) );
  IV U61527 ( .A(n48667), .Z(n48671) );
  NOR U61528 ( .A(n48669), .B(n48668), .Z(n48670) );
  IV U61529 ( .A(n48670), .Z(n50789) );
  NOR U61530 ( .A(n48671), .B(n50789), .Z(n52308) );
  IV U61531 ( .A(n48672), .Z(n48675) );
  NOR U61532 ( .A(n48673), .B(n48680), .Z(n48674) );
  IV U61533 ( .A(n48674), .Z(n50786) );
  NOR U61534 ( .A(n48675), .B(n50786), .Z(n52313) );
  IV U61535 ( .A(n48676), .Z(n52329) );
  NOR U61536 ( .A(n48677), .B(n52329), .Z(n48681) );
  IV U61537 ( .A(n48678), .Z(n48679) );
  NOR U61538 ( .A(n48680), .B(n48679), .Z(n52321) );
  NOR U61539 ( .A(n48681), .B(n52321), .Z(n50783) );
  NOR U61540 ( .A(n48683), .B(n48682), .Z(n54340) );
  IV U61541 ( .A(n54340), .Z(n54336) );
  NOR U61542 ( .A(n48685), .B(n48684), .Z(n58026) );
  NOR U61543 ( .A(n58026), .B(n52330), .Z(n54332) );
  NOR U61544 ( .A(n52331), .B(n48686), .Z(n48688) );
  NOR U61545 ( .A(n48688), .B(n48687), .Z(n50782) );
  IV U61546 ( .A(n48689), .Z(n48690) );
  NOR U61547 ( .A(n48691), .B(n48690), .Z(n54306) );
  NOR U61548 ( .A(n48693), .B(n48692), .Z(n52333) );
  NOR U61549 ( .A(n54306), .B(n52333), .Z(n50780) );
  IV U61550 ( .A(n48694), .Z(n48697) );
  NOR U61551 ( .A(n48695), .B(n50756), .Z(n48696) );
  IV U61552 ( .A(n48696), .Z(n50776) );
  NOR U61553 ( .A(n48697), .B(n50776), .Z(n50770) );
  IV U61554 ( .A(n48698), .Z(n48700) );
  NOR U61555 ( .A(n48700), .B(n48699), .Z(n52337) );
  NOR U61556 ( .A(n52341), .B(n52337), .Z(n50754) );
  NOR U61557 ( .A(n48702), .B(n48701), .Z(n54296) );
  IV U61558 ( .A(n48703), .Z(n48706) );
  IV U61559 ( .A(n48704), .Z(n48705) );
  NOR U61560 ( .A(n48706), .B(n48705), .Z(n48707) );
  IV U61561 ( .A(n48707), .Z(n52346) );
  IV U61562 ( .A(n48708), .Z(n48711) );
  NOR U61563 ( .A(n48709), .B(n50735), .Z(n48710) );
  IV U61564 ( .A(n48710), .Z(n48714) );
  NOR U61565 ( .A(n48711), .B(n48714), .Z(n48712) );
  IV U61566 ( .A(n48712), .Z(n52350) );
  IV U61567 ( .A(n48713), .Z(n48715) );
  NOR U61568 ( .A(n48715), .B(n48714), .Z(n50742) );
  IV U61569 ( .A(n50742), .Z(n50734) );
  IV U61570 ( .A(n48716), .Z(n52354) );
  IV U61571 ( .A(n48717), .Z(n48718) );
  NOR U61572 ( .A(n48718), .B(n48720), .Z(n52358) );
  IV U61573 ( .A(n48719), .Z(n48721) );
  NOR U61574 ( .A(n48721), .B(n48720), .Z(n52356) );
  NOR U61575 ( .A(n52358), .B(n52356), .Z(n50717) );
  IV U61576 ( .A(n48722), .Z(n48723) );
  NOR U61577 ( .A(n48723), .B(n50696), .Z(n54257) );
  IV U61578 ( .A(n50688), .Z(n50683) );
  NOR U61579 ( .A(n48724), .B(n50685), .Z(n54228) );
  NOR U61580 ( .A(n52369), .B(n54215), .Z(n50682) );
  IV U61581 ( .A(n48725), .Z(n48726) );
  NOR U61582 ( .A(n52386), .B(n48726), .Z(n52373) );
  IV U61583 ( .A(n48727), .Z(n48728) );
  NOR U61584 ( .A(n52386), .B(n48728), .Z(n54211) );
  NOR U61585 ( .A(n52373), .B(n54211), .Z(n50681) );
  NOR U61586 ( .A(n48729), .B(n52399), .Z(n54202) );
  IV U61587 ( .A(n48730), .Z(n48733) );
  IV U61588 ( .A(n48731), .Z(n48732) );
  NOR U61589 ( .A(n48733), .B(n48732), .Z(n52397) );
  IV U61590 ( .A(n48734), .Z(n48736) );
  NOR U61591 ( .A(n48736), .B(n48735), .Z(n54196) );
  IV U61592 ( .A(n48737), .Z(n48739) );
  NOR U61593 ( .A(n48739), .B(n48738), .Z(n52406) );
  NOR U61594 ( .A(n54193), .B(n52406), .Z(n50670) );
  IV U61595 ( .A(n48740), .Z(n50669) );
  IV U61596 ( .A(n48741), .Z(n48742) );
  NOR U61597 ( .A(n50669), .B(n48742), .Z(n50664) );
  IV U61598 ( .A(n50664), .Z(n50649) );
  IV U61599 ( .A(n48743), .Z(n50641) );
  IV U61600 ( .A(n48744), .Z(n48745) );
  NOR U61601 ( .A(n50641), .B(n48745), .Z(n50646) );
  IV U61602 ( .A(n50646), .Z(n50638) );
  NOR U61603 ( .A(n48747), .B(n48746), .Z(n50624) );
  IV U61604 ( .A(n50621), .Z(n50614) );
  IV U61605 ( .A(n48748), .Z(n48749) );
  NOR U61606 ( .A(n48749), .B(n50616), .Z(n50609) );
  IV U61607 ( .A(n48750), .Z(n48751) );
  NOR U61608 ( .A(n48752), .B(n48751), .Z(n50606) );
  IV U61609 ( .A(n50606), .Z(n50597) );
  IV U61610 ( .A(n48753), .Z(n54170) );
  NOR U61611 ( .A(n48754), .B(n54170), .Z(n50596) );
  IV U61612 ( .A(n48755), .Z(n48758) );
  NOR U61613 ( .A(n48758), .B(n48756), .Z(n54166) );
  NOR U61614 ( .A(n48758), .B(n48757), .Z(n48759) );
  IV U61615 ( .A(n48759), .Z(n54162) );
  IV U61616 ( .A(n48760), .Z(n48761) );
  NOR U61617 ( .A(n48761), .B(n48763), .Z(n54158) );
  IV U61618 ( .A(n48762), .Z(n48764) );
  NOR U61619 ( .A(n48764), .B(n48763), .Z(n52430) );
  IV U61620 ( .A(n48765), .Z(n48770) );
  IV U61621 ( .A(n48766), .Z(n48767) );
  NOR U61622 ( .A(n48770), .B(n48767), .Z(n52427) );
  IV U61623 ( .A(n48768), .Z(n48769) );
  NOR U61624 ( .A(n48770), .B(n48769), .Z(n52438) );
  IV U61625 ( .A(n48771), .Z(n48773) );
  IV U61626 ( .A(n48772), .Z(n50588) );
  NOR U61627 ( .A(n48773), .B(n50588), .Z(n50585) );
  IV U61628 ( .A(n50585), .Z(n50577) );
  IV U61629 ( .A(n48774), .Z(n48776) );
  IV U61630 ( .A(n48775), .Z(n48778) );
  NOR U61631 ( .A(n48776), .B(n48778), .Z(n52452) );
  IV U61632 ( .A(n48777), .Z(n48779) );
  NOR U61633 ( .A(n48779), .B(n48778), .Z(n50567) );
  IV U61634 ( .A(n50567), .Z(n50557) );
  IV U61635 ( .A(n48780), .Z(n48781) );
  NOR U61636 ( .A(n50559), .B(n48781), .Z(n50554) );
  IV U61637 ( .A(n50554), .Z(n50549) );
  IV U61638 ( .A(n48782), .Z(n50552) );
  IV U61639 ( .A(n48783), .Z(n48784) );
  NOR U61640 ( .A(n50552), .B(n48784), .Z(n54147) );
  IV U61641 ( .A(n48785), .Z(n48787) );
  NOR U61642 ( .A(n48787), .B(n48786), .Z(n52464) );
  IV U61643 ( .A(n48788), .Z(n48789) );
  NOR U61644 ( .A(n50526), .B(n48789), .Z(n50527) );
  IV U61645 ( .A(n48790), .Z(n48792) );
  NOR U61646 ( .A(n48792), .B(n48791), .Z(n50503) );
  IV U61647 ( .A(n48793), .Z(n48794) );
  NOR U61648 ( .A(n48795), .B(n48794), .Z(n54119) );
  IV U61649 ( .A(n48796), .Z(n48799) );
  IV U61650 ( .A(n48797), .Z(n48798) );
  NOR U61651 ( .A(n48799), .B(n48798), .Z(n52504) );
  IV U61652 ( .A(n48800), .Z(n48802) );
  XOR U61653 ( .A(n48808), .B(n48809), .Z(n48801) );
  NOR U61654 ( .A(n48802), .B(n48801), .Z(n52501) );
  IV U61655 ( .A(n48803), .Z(n48804) );
  NOR U61656 ( .A(n48804), .B(n48809), .Z(n54110) );
  IV U61657 ( .A(n48805), .Z(n48807) );
  NOR U61658 ( .A(n48807), .B(n48806), .Z(n54096) );
  IV U61659 ( .A(n48808), .Z(n48810) );
  NOR U61660 ( .A(n48810), .B(n48809), .Z(n54113) );
  NOR U61661 ( .A(n54096), .B(n54113), .Z(n50480) );
  IV U61662 ( .A(n48811), .Z(n48812) );
  NOR U61663 ( .A(n48813), .B(n48812), .Z(n54090) );
  IV U61664 ( .A(n48814), .Z(n48815) );
  NOR U61665 ( .A(n48816), .B(n48815), .Z(n54102) );
  NOR U61666 ( .A(n54090), .B(n54102), .Z(n50479) );
  IV U61667 ( .A(n48817), .Z(n48818) );
  NOR U61668 ( .A(n48818), .B(n48823), .Z(n52507) );
  IV U61669 ( .A(n48819), .Z(n54079) );
  NOR U61670 ( .A(n48820), .B(n54079), .Z(n48821) );
  NOR U61671 ( .A(n52507), .B(n48821), .Z(n50478) );
  IV U61672 ( .A(n48822), .Z(n48824) );
  NOR U61673 ( .A(n48824), .B(n48823), .Z(n48825) );
  IV U61674 ( .A(n48825), .Z(n52511) );
  IV U61675 ( .A(n48826), .Z(n48827) );
  NOR U61676 ( .A(n48828), .B(n48827), .Z(n48833) );
  IV U61677 ( .A(n48829), .Z(n48830) );
  NOR U61678 ( .A(n48831), .B(n48830), .Z(n48832) );
  NOR U61679 ( .A(n48833), .B(n48832), .Z(n54072) );
  IV U61680 ( .A(n48834), .Z(n48836) );
  IV U61681 ( .A(n48835), .Z(n50475) );
  NOR U61682 ( .A(n48836), .B(n50475), .Z(n50470) );
  IV U61683 ( .A(n48837), .Z(n48838) );
  NOR U61684 ( .A(n48838), .B(n50462), .Z(n50467) );
  IV U61685 ( .A(n50467), .Z(n50459) );
  IV U61686 ( .A(n48839), .Z(n48840) );
  NOR U61687 ( .A(n48840), .B(n48849), .Z(n52520) );
  IV U61688 ( .A(n48841), .Z(n48842) );
  NOR U61689 ( .A(n48843), .B(n48842), .Z(n52529) );
  IV U61690 ( .A(n48844), .Z(n48846) );
  NOR U61691 ( .A(n48846), .B(n48845), .Z(n52525) );
  NOR U61692 ( .A(n52529), .B(n52525), .Z(n50457) );
  IV U61693 ( .A(n48847), .Z(n48848) );
  NOR U61694 ( .A(n48849), .B(n48848), .Z(n52523) );
  IV U61695 ( .A(n48850), .Z(n48852) );
  NOR U61696 ( .A(n48852), .B(n48851), .Z(n52531) );
  NOR U61697 ( .A(n54053), .B(n52531), .Z(n50455) );
  NOR U61698 ( .A(n48854), .B(n48853), .Z(n52534) );
  NOR U61699 ( .A(n52542), .B(n52534), .Z(n50454) );
  IV U61700 ( .A(n48855), .Z(n48858) );
  NOR U61701 ( .A(n48856), .B(n50446), .Z(n48857) );
  IV U61702 ( .A(n48857), .Z(n50451) );
  NOR U61703 ( .A(n48858), .B(n50451), .Z(n52537) );
  IV U61704 ( .A(n52537), .Z(n52539) );
  IV U61705 ( .A(n48859), .Z(n57725) );
  IV U61706 ( .A(n48860), .Z(n48861) );
  NOR U61707 ( .A(n57725), .B(n48861), .Z(n52553) );
  NOR U61708 ( .A(n48863), .B(n48862), .Z(n50434) );
  IV U61709 ( .A(n48864), .Z(n50424) );
  NOR U61710 ( .A(n48865), .B(n50424), .Z(n50422) );
  NOR U61711 ( .A(n48867), .B(n48866), .Z(n52574) );
  IV U61712 ( .A(n48868), .Z(n48872) );
  IV U61713 ( .A(n48869), .Z(n48874) );
  NOR U61714 ( .A(n48870), .B(n48874), .Z(n48871) );
  IV U61715 ( .A(n48871), .Z(n50419) );
  NOR U61716 ( .A(n48872), .B(n50419), .Z(n52577) );
  IV U61717 ( .A(n48873), .Z(n48875) );
  NOR U61718 ( .A(n48875), .B(n48874), .Z(n50412) );
  IV U61719 ( .A(n48876), .Z(n48877) );
  NOR U61720 ( .A(n50409), .B(n48877), .Z(n50404) );
  IV U61721 ( .A(n50404), .Z(n50396) );
  IV U61722 ( .A(n48878), .Z(n48880) );
  NOR U61723 ( .A(n48880), .B(n48879), .Z(n48881) );
  IV U61724 ( .A(n48881), .Z(n50381) );
  IV U61725 ( .A(n48882), .Z(n48889) );
  IV U61726 ( .A(n48883), .Z(n50364) );
  NOR U61727 ( .A(n50364), .B(n48884), .Z(n48885) );
  IV U61728 ( .A(n48885), .Z(n48886) );
  NOR U61729 ( .A(n48887), .B(n48886), .Z(n48888) );
  IV U61730 ( .A(n48888), .Z(n48892) );
  NOR U61731 ( .A(n48889), .B(n48892), .Z(n48890) );
  IV U61732 ( .A(n48890), .Z(n54010) );
  IV U61733 ( .A(n48891), .Z(n48893) );
  NOR U61734 ( .A(n48893), .B(n48892), .Z(n48894) );
  IV U61735 ( .A(n48894), .Z(n52604) );
  IV U61736 ( .A(n48895), .Z(n48897) );
  NOR U61737 ( .A(n48897), .B(n48896), .Z(n48898) );
  NOR U61738 ( .A(n48899), .B(n48898), .Z(n54008) );
  NOR U61739 ( .A(n48901), .B(n48900), .Z(n54004) );
  NOR U61740 ( .A(n48903), .B(n48902), .Z(n53991) );
  IV U61741 ( .A(n48904), .Z(n48905) );
  NOR U61742 ( .A(n48909), .B(n48905), .Z(n52619) );
  NOR U61743 ( .A(n48907), .B(n48906), .Z(n48913) );
  NOR U61744 ( .A(n48909), .B(n48908), .Z(n48910) );
  NOR U61745 ( .A(n48911), .B(n48910), .Z(n48912) );
  NOR U61746 ( .A(n48913), .B(n48912), .Z(n53986) );
  IV U61747 ( .A(n48914), .Z(n48915) );
  NOR U61748 ( .A(n50336), .B(n48915), .Z(n53983) );
  IV U61749 ( .A(n48916), .Z(n48917) );
  NOR U61750 ( .A(n48917), .B(n50331), .Z(n52630) );
  IV U61751 ( .A(n48918), .Z(n48920) );
  IV U61752 ( .A(n48919), .Z(n50296) );
  NOR U61753 ( .A(n48920), .B(n50296), .Z(n50305) );
  IV U61754 ( .A(n48921), .Z(n48922) );
  NOR U61755 ( .A(n48922), .B(n50296), .Z(n50302) );
  IV U61756 ( .A(n50302), .Z(n50293) );
  IV U61757 ( .A(n48923), .Z(n50284) );
  NOR U61758 ( .A(n48924), .B(n50284), .Z(n50282) );
  IV U61759 ( .A(n48925), .Z(n48926) );
  NOR U61760 ( .A(n50280), .B(n48926), .Z(n52651) );
  NOR U61761 ( .A(n48928), .B(n48927), .Z(n48929) );
  IV U61762 ( .A(n48929), .Z(n53954) );
  IV U61763 ( .A(n48930), .Z(n48931) );
  NOR U61764 ( .A(n48932), .B(n48931), .Z(n52668) );
  IV U61765 ( .A(n48933), .Z(n48935) );
  NOR U61766 ( .A(n48935), .B(n48934), .Z(n53939) );
  NOR U61767 ( .A(n52668), .B(n53939), .Z(n50267) );
  IV U61768 ( .A(n48936), .Z(n48937) );
  NOR U61769 ( .A(n48937), .B(n50265), .Z(n53934) );
  IV U61770 ( .A(n48938), .Z(n48943) );
  IV U61771 ( .A(n48939), .Z(n48940) );
  NOR U61772 ( .A(n48940), .B(n48947), .Z(n48941) );
  IV U61773 ( .A(n48941), .Z(n48942) );
  NOR U61774 ( .A(n48943), .B(n48942), .Z(n53923) );
  IV U61775 ( .A(n48944), .Z(n52676) );
  NOR U61776 ( .A(n52676), .B(n48945), .Z(n48952) );
  IV U61777 ( .A(n48946), .Z(n48951) );
  NOR U61778 ( .A(n48948), .B(n48947), .Z(n48949) );
  IV U61779 ( .A(n48949), .Z(n48950) );
  NOR U61780 ( .A(n48951), .B(n48950), .Z(n53920) );
  NOR U61781 ( .A(n48952), .B(n53920), .Z(n50255) );
  IV U61782 ( .A(n48953), .Z(n48955) );
  NOR U61783 ( .A(n48955), .B(n48954), .Z(n52685) );
  IV U61784 ( .A(n48956), .Z(n48959) );
  IV U61785 ( .A(n48957), .Z(n50251) );
  XOR U61786 ( .A(n50251), .B(n48961), .Z(n48958) );
  NOR U61787 ( .A(n48959), .B(n48958), .Z(n52682) );
  IV U61788 ( .A(n48960), .Z(n48962) );
  IV U61789 ( .A(n48961), .Z(n50250) );
  NOR U61790 ( .A(n48962), .B(n50250), .Z(n52691) );
  NOR U61791 ( .A(n48963), .B(n50250), .Z(n48964) );
  IV U61792 ( .A(n48964), .Z(n48965) );
  NOR U61793 ( .A(n48966), .B(n48965), .Z(n52689) );
  NOR U61794 ( .A(n52691), .B(n52689), .Z(n50254) );
  IV U61795 ( .A(n52701), .Z(n52698) );
  IV U61796 ( .A(n48967), .Z(n53900) );
  IV U61797 ( .A(n48968), .Z(n48974) );
  IV U61798 ( .A(n48969), .Z(n50218) );
  XOR U61799 ( .A(n50218), .B(n48975), .Z(n48970) );
  NOR U61800 ( .A(n48971), .B(n48970), .Z(n48972) );
  IV U61801 ( .A(n48972), .Z(n48973) );
  NOR U61802 ( .A(n48974), .B(n48973), .Z(n52720) );
  IV U61803 ( .A(n48975), .Z(n52724) );
  NOR U61804 ( .A(n48976), .B(n52724), .Z(n50222) );
  IV U61805 ( .A(n48977), .Z(n48979) );
  NOR U61806 ( .A(n48979), .B(n48978), .Z(n50181) );
  IV U61807 ( .A(n48980), .Z(n50159) );
  IV U61808 ( .A(n48981), .Z(n48982) );
  NOR U61809 ( .A(n50159), .B(n48982), .Z(n52751) );
  NOR U61810 ( .A(n48984), .B(n48983), .Z(n48985) );
  IV U61811 ( .A(n48985), .Z(n50161) );
  IV U61812 ( .A(n48986), .Z(n50157) );
  IV U61813 ( .A(n48987), .Z(n48988) );
  NOR U61814 ( .A(n50157), .B(n48988), .Z(n53860) );
  IV U61815 ( .A(n48989), .Z(n48990) );
  NOR U61816 ( .A(n48990), .B(n48992), .Z(n52762) );
  IV U61817 ( .A(n48991), .Z(n48993) );
  NOR U61818 ( .A(n48993), .B(n48992), .Z(n52759) );
  IV U61819 ( .A(n48994), .Z(n48995) );
  NOR U61820 ( .A(n48996), .B(n48995), .Z(n52767) );
  IV U61821 ( .A(n48997), .Z(n48998) );
  NOR U61822 ( .A(n48999), .B(n48998), .Z(n52772) );
  NOR U61823 ( .A(n52767), .B(n52772), .Z(n50146) );
  IV U61824 ( .A(n49000), .Z(n49003) );
  IV U61825 ( .A(n49001), .Z(n49002) );
  NOR U61826 ( .A(n49003), .B(n49002), .Z(n52769) );
  IV U61827 ( .A(n49004), .Z(n49005) );
  NOR U61828 ( .A(n49006), .B(n49005), .Z(n52776) );
  NOR U61829 ( .A(n52778), .B(n52776), .Z(n50145) );
  IV U61830 ( .A(n49007), .Z(n49009) );
  NOR U61831 ( .A(n49009), .B(n49008), .Z(n52790) );
  NOR U61832 ( .A(n52781), .B(n52790), .Z(n50144) );
  IV U61833 ( .A(n49010), .Z(n49012) );
  NOR U61834 ( .A(n49012), .B(n49011), .Z(n50128) );
  IV U61835 ( .A(n49013), .Z(n49014) );
  NOR U61836 ( .A(n49015), .B(n49014), .Z(n53834) );
  IV U61837 ( .A(n49016), .Z(n49017) );
  NOR U61838 ( .A(n49017), .B(n50112), .Z(n53838) );
  NOR U61839 ( .A(n53834), .B(n53838), .Z(n50115) );
  IV U61840 ( .A(n49018), .Z(n49019) );
  NOR U61841 ( .A(n49019), .B(n49021), .Z(n53831) );
  IV U61842 ( .A(n49020), .Z(n49022) );
  NOR U61843 ( .A(n49022), .B(n49021), .Z(n52803) );
  IV U61844 ( .A(n49023), .Z(n49024) );
  NOR U61845 ( .A(n49024), .B(n49027), .Z(n50086) );
  IV U61846 ( .A(n49025), .Z(n49026) );
  NOR U61847 ( .A(n49027), .B(n49026), .Z(n49028) );
  IV U61848 ( .A(n49028), .Z(n52809) );
  IV U61849 ( .A(n49029), .Z(n49030) );
  NOR U61850 ( .A(n49031), .B(n49030), .Z(n52806) );
  IV U61851 ( .A(n49032), .Z(n49035) );
  IV U61852 ( .A(n49033), .Z(n49034) );
  NOR U61853 ( .A(n49035), .B(n49034), .Z(n53821) );
  NOR U61854 ( .A(n52806), .B(n53821), .Z(n50083) );
  IV U61855 ( .A(n49036), .Z(n49038) );
  NOR U61856 ( .A(n49038), .B(n49037), .Z(n49039) );
  IV U61857 ( .A(n49039), .Z(n53819) );
  IV U61858 ( .A(n49040), .Z(n49042) );
  NOR U61859 ( .A(n49042), .B(n49041), .Z(n53812) );
  NOR U61860 ( .A(n53815), .B(n53812), .Z(n50082) );
  IV U61861 ( .A(n49043), .Z(n49044) );
  NOR U61862 ( .A(n49051), .B(n49044), .Z(n53811) );
  IV U61863 ( .A(n49045), .Z(n49048) );
  NOR U61864 ( .A(n49054), .B(n49046), .Z(n49047) );
  IV U61865 ( .A(n49047), .Z(n49056) );
  NOR U61866 ( .A(n49048), .B(n49056), .Z(n52816) );
  IV U61867 ( .A(n49049), .Z(n49050) );
  NOR U61868 ( .A(n49051), .B(n49050), .Z(n52814) );
  NOR U61869 ( .A(n52816), .B(n52814), .Z(n50080) );
  IV U61870 ( .A(n49052), .Z(n49053) );
  NOR U61871 ( .A(n49054), .B(n49053), .Z(n52812) );
  IV U61872 ( .A(n49055), .Z(n49057) );
  NOR U61873 ( .A(n49057), .B(n49056), .Z(n53799) );
  IV U61874 ( .A(n49058), .Z(n49062) );
  NOR U61875 ( .A(n49060), .B(n49059), .Z(n49061) );
  IV U61876 ( .A(n49061), .Z(n49064) );
  NOR U61877 ( .A(n49062), .B(n49064), .Z(n53796) );
  NOR U61878 ( .A(n49064), .B(n49063), .Z(n49065) );
  IV U61879 ( .A(n49065), .Z(n49070) );
  NOR U61880 ( .A(n49067), .B(n49066), .Z(n49068) );
  IV U61881 ( .A(n49068), .Z(n49069) );
  NOR U61882 ( .A(n49070), .B(n49069), .Z(n49071) );
  IV U61883 ( .A(n49071), .Z(n49072) );
  NOR U61884 ( .A(n49073), .B(n49072), .Z(n53785) );
  IV U61885 ( .A(n49074), .Z(n52833) );
  IV U61886 ( .A(n49075), .Z(n49076) );
  NOR U61887 ( .A(n49076), .B(n50033), .Z(n49077) );
  IV U61888 ( .A(n49077), .Z(n53762) );
  IV U61889 ( .A(n49078), .Z(n50017) );
  NOR U61890 ( .A(n49080), .B(n49079), .Z(n52855) );
  IV U61891 ( .A(n49081), .Z(n49082) );
  NOR U61892 ( .A(n49083), .B(n49082), .Z(n53753) );
  NOR U61893 ( .A(n49085), .B(n49084), .Z(n53758) );
  NOR U61894 ( .A(n53753), .B(n53758), .Z(n50008) );
  IV U61895 ( .A(n49086), .Z(n49089) );
  NOR U61896 ( .A(n50001), .B(n49087), .Z(n49088) );
  IV U61897 ( .A(n49088), .Z(n49996) );
  NOR U61898 ( .A(n49089), .B(n49996), .Z(n52871) );
  IV U61899 ( .A(n49090), .Z(n49092) );
  IV U61900 ( .A(n49091), .Z(n49989) );
  NOR U61901 ( .A(n49092), .B(n49989), .Z(n52876) );
  IV U61902 ( .A(n52876), .Z(n52874) );
  IV U61903 ( .A(n49093), .Z(n49095) );
  IV U61904 ( .A(n49094), .Z(n49103) );
  NOR U61905 ( .A(n49095), .B(n49103), .Z(n52900) );
  IV U61906 ( .A(n49096), .Z(n49097) );
  NOR U61907 ( .A(n49097), .B(n49099), .Z(n52909) );
  IV U61908 ( .A(n49098), .Z(n49100) );
  NOR U61909 ( .A(n49100), .B(n49099), .Z(n52914) );
  NOR U61910 ( .A(n52909), .B(n52914), .Z(n49101) );
  IV U61911 ( .A(n49101), .Z(n49113) );
  NOR U61912 ( .A(n49103), .B(n49102), .Z(n49104) );
  IV U61913 ( .A(n49104), .Z(n49109) );
  NOR U61914 ( .A(n49106), .B(n49105), .Z(n49107) );
  IV U61915 ( .A(n49107), .Z(n49108) );
  NOR U61916 ( .A(n49109), .B(n49108), .Z(n49110) );
  IV U61917 ( .A(n49110), .Z(n49111) );
  NOR U61918 ( .A(n49112), .B(n49111), .Z(n52907) );
  NOR U61919 ( .A(n49113), .B(n52907), .Z(n49965) );
  IV U61920 ( .A(n49114), .Z(n49115) );
  NOR U61921 ( .A(n49115), .B(n49120), .Z(n52917) );
  IV U61922 ( .A(n49116), .Z(n49118) );
  NOR U61923 ( .A(n49118), .B(n49117), .Z(n53744) );
  IV U61924 ( .A(n49119), .Z(n49121) );
  NOR U61925 ( .A(n49121), .B(n49120), .Z(n53739) );
  NOR U61926 ( .A(n53744), .B(n53739), .Z(n49954) );
  IV U61927 ( .A(n49122), .Z(n49123) );
  NOR U61928 ( .A(n49124), .B(n49123), .Z(n49125) );
  IV U61929 ( .A(n49125), .Z(n49945) );
  IV U61930 ( .A(n49126), .Z(n49948) );
  IV U61931 ( .A(n49127), .Z(n49128) );
  NOR U61932 ( .A(n49948), .B(n49128), .Z(n53732) );
  IV U61933 ( .A(n49129), .Z(n49131) );
  NOR U61934 ( .A(n49131), .B(n49130), .Z(n52920) );
  NOR U61935 ( .A(n53732), .B(n52920), .Z(n49932) );
  NOR U61936 ( .A(n49132), .B(n49136), .Z(n49133) );
  IV U61937 ( .A(n49133), .Z(n52924) );
  NOR U61938 ( .A(n52924), .B(n49134), .Z(n49931) );
  IV U61939 ( .A(n49135), .Z(n49137) );
  NOR U61940 ( .A(n49137), .B(n49136), .Z(n53718) );
  NOR U61941 ( .A(n52928), .B(n53718), .Z(n49929) );
  IV U61942 ( .A(n49138), .Z(n49140) );
  NOR U61943 ( .A(n49140), .B(n49139), .Z(n49141) );
  IV U61944 ( .A(n49141), .Z(n49923) );
  IV U61945 ( .A(n49142), .Z(n49144) );
  NOR U61946 ( .A(n49144), .B(n49143), .Z(n49149) );
  IV U61947 ( .A(n49145), .Z(n49146) );
  NOR U61948 ( .A(n49147), .B(n49146), .Z(n49148) );
  NOR U61949 ( .A(n49149), .B(n49148), .Z(n52949) );
  NOR U61950 ( .A(n49151), .B(n49150), .Z(n52945) );
  IV U61951 ( .A(n49152), .Z(n49157) );
  IV U61952 ( .A(n49153), .Z(n49154) );
  NOR U61953 ( .A(n49157), .B(n49154), .Z(n52953) );
  IV U61954 ( .A(n49155), .Z(n49156) );
  NOR U61955 ( .A(n49157), .B(n49156), .Z(n52958) );
  NOR U61956 ( .A(n52953), .B(n52958), .Z(n49158) );
  IV U61957 ( .A(n49158), .Z(n49164) );
  IV U61958 ( .A(n49159), .Z(n49161) );
  NOR U61959 ( .A(n49161), .B(n49160), .Z(n52952) );
  NOR U61960 ( .A(n52952), .B(n53703), .Z(n49162) );
  IV U61961 ( .A(n49162), .Z(n49163) );
  NOR U61962 ( .A(n49164), .B(n49163), .Z(n49915) );
  IV U61963 ( .A(n49165), .Z(n49166) );
  NOR U61964 ( .A(n49166), .B(n49175), .Z(n52955) );
  IV U61965 ( .A(n49167), .Z(n49169) );
  NOR U61966 ( .A(n49169), .B(n49168), .Z(n52963) );
  IV U61967 ( .A(n49170), .Z(n49171) );
  NOR U61968 ( .A(n49172), .B(n49171), .Z(n52967) );
  IV U61969 ( .A(n49173), .Z(n49174) );
  NOR U61970 ( .A(n49175), .B(n49174), .Z(n52961) );
  NOR U61971 ( .A(n52967), .B(n52961), .Z(n49914) );
  IV U61972 ( .A(n49176), .Z(n49910) );
  IV U61973 ( .A(n49177), .Z(n49178) );
  NOR U61974 ( .A(n49910), .B(n49178), .Z(n52970) );
  IV U61975 ( .A(n49179), .Z(n53698) );
  NOR U61976 ( .A(n49180), .B(n53698), .Z(n52980) );
  IV U61977 ( .A(n49181), .Z(n49182) );
  NOR U61978 ( .A(n49185), .B(n49182), .Z(n52986) );
  IV U61979 ( .A(n49183), .Z(n49184) );
  NOR U61980 ( .A(n49185), .B(n49184), .Z(n52992) );
  IV U61981 ( .A(n49186), .Z(n49188) );
  NOR U61982 ( .A(n49188), .B(n49187), .Z(n52989) );
  IV U61983 ( .A(n49189), .Z(n49199) );
  NOR U61984 ( .A(n49905), .B(n49190), .Z(n49191) );
  IV U61985 ( .A(n49191), .Z(n49196) );
  NOR U61986 ( .A(n49193), .B(n49192), .Z(n49194) );
  IV U61987 ( .A(n49194), .Z(n49195) );
  NOR U61988 ( .A(n49196), .B(n49195), .Z(n49197) );
  IV U61989 ( .A(n49197), .Z(n49198) );
  NOR U61990 ( .A(n49199), .B(n49198), .Z(n49200) );
  IV U61991 ( .A(n49200), .Z(n49201) );
  NOR U61992 ( .A(n49202), .B(n49201), .Z(n53689) );
  IV U61993 ( .A(n49203), .Z(n49205) );
  NOR U61994 ( .A(n49205), .B(n49204), .Z(n49899) );
  IV U61995 ( .A(n49206), .Z(n49208) );
  NOR U61996 ( .A(n49208), .B(n49207), .Z(n49896) );
  IV U61997 ( .A(n49896), .Z(n49891) );
  IV U61998 ( .A(n49209), .Z(n49210) );
  NOR U61999 ( .A(n49210), .B(n49887), .Z(n53682) );
  IV U62000 ( .A(n49211), .Z(n49213) );
  NOR U62001 ( .A(n49213), .B(n49212), .Z(n53004) );
  NOR U62002 ( .A(n53682), .B(n53004), .Z(n49890) );
  IV U62003 ( .A(n49214), .Z(n49216) );
  IV U62004 ( .A(n49215), .Z(n49219) );
  NOR U62005 ( .A(n49216), .B(n49219), .Z(n53665) );
  NOR U62006 ( .A(n49217), .B(n53013), .Z(n49221) );
  IV U62007 ( .A(n49218), .Z(n49220) );
  NOR U62008 ( .A(n49220), .B(n49219), .Z(n53662) );
  NOR U62009 ( .A(n49221), .B(n53662), .Z(n49882) );
  IV U62010 ( .A(n49222), .Z(n49223) );
  NOR U62011 ( .A(n49224), .B(n49223), .Z(n49229) );
  IV U62012 ( .A(n49225), .Z(n49226) );
  NOR U62013 ( .A(n49227), .B(n49226), .Z(n49228) );
  NOR U62014 ( .A(n49229), .B(n49228), .Z(n53657) );
  NOR U62015 ( .A(n49231), .B(n49230), .Z(n53653) );
  IV U62016 ( .A(n49232), .Z(n49234) );
  NOR U62017 ( .A(n49234), .B(n49233), .Z(n53648) );
  NOR U62018 ( .A(n53648), .B(n53016), .Z(n49881) );
  IV U62019 ( .A(n49235), .Z(n49867) );
  NOR U62020 ( .A(n49237), .B(n49236), .Z(n49873) );
  IV U62021 ( .A(n49238), .Z(n49851) );
  IV U62022 ( .A(n49239), .Z(n49240) );
  NOR U62023 ( .A(n49241), .B(n49240), .Z(n53638) );
  IV U62024 ( .A(n49242), .Z(n49243) );
  NOR U62025 ( .A(n49244), .B(n49243), .Z(n53640) );
  NOR U62026 ( .A(n53638), .B(n53640), .Z(n49847) );
  IV U62027 ( .A(n49245), .Z(n49255) );
  XOR U62028 ( .A(n49255), .B(n49253), .Z(n49246) );
  NOR U62029 ( .A(n49247), .B(n49246), .Z(n49248) );
  IV U62030 ( .A(n49248), .Z(n49249) );
  NOR U62031 ( .A(n49250), .B(n49249), .Z(n49251) );
  IV U62032 ( .A(n49251), .Z(n53029) );
  NOR U62033 ( .A(n53029), .B(n49252), .Z(n49846) );
  IV U62034 ( .A(n49253), .Z(n49254) );
  NOR U62035 ( .A(n49255), .B(n49254), .Z(n53033) );
  NOR U62036 ( .A(n53038), .B(n53033), .Z(n49845) );
  IV U62037 ( .A(n49256), .Z(n49260) );
  NOR U62038 ( .A(n49258), .B(n49257), .Z(n49259) );
  IV U62039 ( .A(n49259), .Z(n49262) );
  NOR U62040 ( .A(n49260), .B(n49262), .Z(n53631) );
  NOR U62041 ( .A(n53041), .B(n53631), .Z(n49844) );
  IV U62042 ( .A(n49261), .Z(n49263) );
  NOR U62043 ( .A(n49263), .B(n49262), .Z(n53630) );
  IV U62044 ( .A(n53630), .Z(n53628) );
  IV U62045 ( .A(n49264), .Z(n49266) );
  NOR U62046 ( .A(n49266), .B(n49265), .Z(n49267) );
  IV U62047 ( .A(n49267), .Z(n53624) );
  IV U62048 ( .A(n49268), .Z(n49269) );
  NOR U62049 ( .A(n49269), .B(n49272), .Z(n53621) );
  IV U62050 ( .A(n49270), .Z(n49271) );
  NOR U62051 ( .A(n49272), .B(n49271), .Z(n53044) );
  IV U62052 ( .A(n49273), .Z(n49275) );
  NOR U62053 ( .A(n49275), .B(n49274), .Z(n49279) );
  IV U62054 ( .A(n49276), .Z(n49277) );
  NOR U62055 ( .A(n49277), .B(n49841), .Z(n49278) );
  NOR U62056 ( .A(n49279), .B(n49278), .Z(n53615) );
  IV U62057 ( .A(n49280), .Z(n49281) );
  NOR U62058 ( .A(n49281), .B(n49834), .Z(n53050) );
  NOR U62059 ( .A(n49283), .B(n49282), .Z(n49284) );
  IV U62060 ( .A(n49284), .Z(n49285) );
  NOR U62061 ( .A(n53067), .B(n49285), .Z(n49829) );
  IV U62062 ( .A(n49286), .Z(n49288) );
  NOR U62063 ( .A(n49288), .B(n49287), .Z(n49289) );
  IV U62064 ( .A(n49289), .Z(n49810) );
  IV U62065 ( .A(n49290), .Z(n49816) );
  IV U62066 ( .A(n49291), .Z(n49292) );
  NOR U62067 ( .A(n49816), .B(n49292), .Z(n49293) );
  IV U62068 ( .A(n49293), .Z(n53073) );
  IV U62069 ( .A(n49294), .Z(n49295) );
  NOR U62070 ( .A(n49295), .B(n49302), .Z(n53081) );
  IV U62071 ( .A(n49296), .Z(n49297) );
  NOR U62072 ( .A(n49816), .B(n49297), .Z(n53078) );
  NOR U62073 ( .A(n53081), .B(n53078), .Z(n49809) );
  IV U62074 ( .A(n49298), .Z(n49803) );
  IV U62075 ( .A(n49299), .Z(n49300) );
  NOR U62076 ( .A(n49803), .B(n49300), .Z(n53087) );
  IV U62077 ( .A(n49301), .Z(n49303) );
  NOR U62078 ( .A(n49303), .B(n49302), .Z(n53085) );
  NOR U62079 ( .A(n53087), .B(n53085), .Z(n49808) );
  IV U62080 ( .A(n49304), .Z(n49305) );
  NOR U62081 ( .A(n49305), .B(n49307), .Z(n53599) );
  IV U62082 ( .A(n49306), .Z(n49310) );
  NOR U62083 ( .A(n49308), .B(n49307), .Z(n49309) );
  IV U62084 ( .A(n49309), .Z(n49799) );
  NOR U62085 ( .A(n49310), .B(n49799), .Z(n53588) );
  IV U62086 ( .A(n49311), .Z(n49313) );
  NOR U62087 ( .A(n49313), .B(n49312), .Z(n53095) );
  NOR U62088 ( .A(n49314), .B(n53095), .Z(n49796) );
  NOR U62089 ( .A(n49316), .B(n49315), .Z(n53573) );
  IV U62090 ( .A(n49317), .Z(n49319) );
  IV U62091 ( .A(n49318), .Z(n49326) );
  NOR U62092 ( .A(n49319), .B(n49326), .Z(n49324) );
  IV U62093 ( .A(n49320), .Z(n49321) );
  NOR U62094 ( .A(n49322), .B(n49321), .Z(n49323) );
  NOR U62095 ( .A(n49324), .B(n49323), .Z(n53572) );
  IV U62096 ( .A(n49325), .Z(n49327) );
  NOR U62097 ( .A(n49327), .B(n49326), .Z(n53097) );
  IV U62098 ( .A(n49328), .Z(n49329) );
  NOR U62099 ( .A(n49334), .B(n49329), .Z(n53104) );
  NOR U62100 ( .A(n53097), .B(n53104), .Z(n49795) );
  IV U62101 ( .A(n49330), .Z(n49336) );
  XOR U62102 ( .A(n49332), .B(n49331), .Z(n49333) );
  NOR U62103 ( .A(n49334), .B(n49333), .Z(n49335) );
  IV U62104 ( .A(n49335), .Z(n49338) );
  NOR U62105 ( .A(n49336), .B(n49338), .Z(n53103) );
  IV U62106 ( .A(n53103), .Z(n53101) );
  IV U62107 ( .A(n49337), .Z(n49339) );
  NOR U62108 ( .A(n49339), .B(n49338), .Z(n49340) );
  IV U62109 ( .A(n49340), .Z(n53113) );
  IV U62110 ( .A(n49341), .Z(n49343) );
  NOR U62111 ( .A(n49343), .B(n49342), .Z(n49784) );
  IV U62112 ( .A(n49784), .Z(n49782) );
  NOR U62113 ( .A(n49344), .B(n49346), .Z(n53127) );
  IV U62114 ( .A(n49345), .Z(n49347) );
  NOR U62115 ( .A(n49347), .B(n49346), .Z(n53567) );
  NOR U62116 ( .A(n49348), .B(n53567), .Z(n49349) );
  IV U62117 ( .A(n49349), .Z(n49781) );
  IV U62118 ( .A(n49350), .Z(n49352) );
  NOR U62119 ( .A(n49352), .B(n49351), .Z(n53133) );
  NOR U62120 ( .A(n53133), .B(n49353), .Z(n49780) );
  IV U62121 ( .A(n49354), .Z(n49355) );
  NOR U62122 ( .A(n49355), .B(n57030), .Z(n49356) );
  IV U62123 ( .A(n49356), .Z(n53131) );
  NOR U62124 ( .A(n56607), .B(n49357), .Z(n49358) );
  NOR U62125 ( .A(n49358), .B(n56608), .Z(n53562) );
  IV U62126 ( .A(n49359), .Z(n49360) );
  NOR U62127 ( .A(n49360), .B(n49368), .Z(n53142) );
  IV U62128 ( .A(n49361), .Z(n49363) );
  NOR U62129 ( .A(n49363), .B(n49362), .Z(n53138) );
  NOR U62130 ( .A(n53142), .B(n53138), .Z(n49779) );
  IV U62131 ( .A(n49364), .Z(n49365) );
  NOR U62132 ( .A(n49366), .B(n49365), .Z(n53145) );
  IV U62133 ( .A(n49367), .Z(n49369) );
  NOR U62134 ( .A(n49369), .B(n49368), .Z(n53141) );
  NOR U62135 ( .A(n53145), .B(n53141), .Z(n49778) );
  IV U62136 ( .A(n49370), .Z(n49372) );
  NOR U62137 ( .A(n49372), .B(n49371), .Z(n53154) );
  IV U62138 ( .A(n49373), .Z(n49376) );
  NOR U62139 ( .A(n49374), .B(n49776), .Z(n49375) );
  IV U62140 ( .A(n49375), .Z(n49378) );
  NOR U62141 ( .A(n49376), .B(n49378), .Z(n53151) );
  IV U62142 ( .A(n49377), .Z(n49379) );
  NOR U62143 ( .A(n49379), .B(n49378), .Z(n53148) );
  IV U62144 ( .A(n49380), .Z(n49381) );
  NOR U62145 ( .A(n49382), .B(n49381), .Z(n53541) );
  NOR U62146 ( .A(n49383), .B(n53537), .Z(n49384) );
  NOR U62147 ( .A(n53541), .B(n49384), .Z(n49767) );
  IV U62148 ( .A(n49385), .Z(n49388) );
  IV U62149 ( .A(n49386), .Z(n49387) );
  NOR U62150 ( .A(n49388), .B(n49387), .Z(n53540) );
  IV U62151 ( .A(n53540), .Z(n53538) );
  IV U62152 ( .A(n49389), .Z(n49391) );
  NOR U62153 ( .A(n49391), .B(n49390), .Z(n49392) );
  IV U62154 ( .A(n49392), .Z(n53157) );
  IV U62155 ( .A(n49393), .Z(n49394) );
  NOR U62156 ( .A(n49395), .B(n49394), .Z(n53159) );
  IV U62157 ( .A(n49396), .Z(n49398) );
  IV U62158 ( .A(n49397), .Z(n49763) );
  NOR U62159 ( .A(n49398), .B(n49763), .Z(n53168) );
  NOR U62160 ( .A(n53521), .B(n53168), .Z(n49766) );
  IV U62161 ( .A(n49399), .Z(n49401) );
  NOR U62162 ( .A(n49401), .B(n49400), .Z(n53512) );
  IV U62163 ( .A(n49402), .Z(n49404) );
  NOR U62164 ( .A(n49404), .B(n49403), .Z(n53509) );
  NOR U62165 ( .A(n53179), .B(n53509), .Z(n49759) );
  IV U62166 ( .A(n53174), .Z(n53177) );
  IV U62167 ( .A(n49405), .Z(n49406) );
  NOR U62168 ( .A(n49407), .B(n49406), .Z(n49408) );
  IV U62169 ( .A(n49408), .Z(n53186) );
  IV U62170 ( .A(n49409), .Z(n49410) );
  NOR U62171 ( .A(n49410), .B(n49757), .Z(n53189) );
  IV U62172 ( .A(n49411), .Z(n49412) );
  NOR U62173 ( .A(n49412), .B(n49757), .Z(n53506) );
  NOR U62174 ( .A(n53189), .B(n53506), .Z(n49755) );
  IV U62175 ( .A(n49413), .Z(n49419) );
  IV U62176 ( .A(n49414), .Z(n49415) );
  NOR U62177 ( .A(n49419), .B(n49415), .Z(n49416) );
  IV U62178 ( .A(n49416), .Z(n53192) );
  IV U62179 ( .A(n49417), .Z(n49418) );
  NOR U62180 ( .A(n49419), .B(n49418), .Z(n53502) );
  IV U62181 ( .A(n49420), .Z(n49750) );
  IV U62182 ( .A(n49421), .Z(n49422) );
  NOR U62183 ( .A(n49750), .B(n49422), .Z(n53495) );
  IV U62184 ( .A(n49423), .Z(n49425) );
  NOR U62185 ( .A(n49425), .B(n49424), .Z(n53492) );
  IV U62186 ( .A(n49426), .Z(n49427) );
  NOR U62187 ( .A(n49427), .B(n49432), .Z(n53196) );
  IV U62188 ( .A(n49428), .Z(n49430) );
  IV U62189 ( .A(n49429), .Z(n49435) );
  NOR U62190 ( .A(n49430), .B(n49435), .Z(n53201) );
  IV U62191 ( .A(n49431), .Z(n49433) );
  NOR U62192 ( .A(n49433), .B(n49432), .Z(n53199) );
  NOR U62193 ( .A(n53201), .B(n53199), .Z(n49744) );
  IV U62194 ( .A(n49434), .Z(n49436) );
  NOR U62195 ( .A(n49436), .B(n49435), .Z(n53206) );
  IV U62196 ( .A(n49437), .Z(n49438) );
  NOR U62197 ( .A(n49439), .B(n49438), .Z(n53203) );
  NOR U62198 ( .A(n49441), .B(n49440), .Z(n49442) );
  NOR U62199 ( .A(n49443), .B(n49442), .Z(n53214) );
  IV U62200 ( .A(n49444), .Z(n49446) );
  NOR U62201 ( .A(n49446), .B(n49445), .Z(n53220) );
  IV U62202 ( .A(n49447), .Z(n49730) );
  NOR U62203 ( .A(n49448), .B(n49730), .Z(n53230) );
  NOR U62204 ( .A(n53478), .B(n53230), .Z(n49719) );
  NOR U62205 ( .A(n49450), .B(n49449), .Z(n53237) );
  IV U62206 ( .A(n49451), .Z(n49452) );
  NOR U62207 ( .A(n49452), .B(n49715), .Z(n53470) );
  IV U62208 ( .A(n49453), .Z(n49454) );
  NOR U62209 ( .A(n49455), .B(n49454), .Z(n49708) );
  IV U62210 ( .A(n49708), .Z(n49698) );
  IV U62211 ( .A(n49456), .Z(n49458) );
  IV U62212 ( .A(n49457), .Z(n49687) );
  NOR U62213 ( .A(n49458), .B(n49687), .Z(n53459) );
  IV U62214 ( .A(n49459), .Z(n49460) );
  NOR U62215 ( .A(n49460), .B(n49687), .Z(n53465) );
  NOR U62216 ( .A(n53459), .B(n53465), .Z(n56873) );
  IV U62217 ( .A(n49461), .Z(n49462) );
  NOR U62218 ( .A(n49462), .B(n49684), .Z(n56869) );
  IV U62219 ( .A(n49463), .Z(n49464) );
  NOR U62220 ( .A(n49465), .B(n49464), .Z(n53250) );
  NOR U62221 ( .A(n53253), .B(n53250), .Z(n49666) );
  NOR U62222 ( .A(n49467), .B(n49466), .Z(n53255) );
  IV U62223 ( .A(n49468), .Z(n49469) );
  NOR U62224 ( .A(n49470), .B(n49469), .Z(n53447) );
  IV U62225 ( .A(n49471), .Z(n49473) );
  NOR U62226 ( .A(n49473), .B(n49472), .Z(n53450) );
  NOR U62227 ( .A(n53447), .B(n53450), .Z(n49664) );
  IV U62228 ( .A(n49474), .Z(n49475) );
  NOR U62229 ( .A(n49654), .B(n49475), .Z(n49476) );
  IV U62230 ( .A(n49476), .Z(n53259) );
  NOR U62231 ( .A(n53264), .B(n53262), .Z(n49648) );
  NOR U62232 ( .A(n49478), .B(n49477), .Z(n49479) );
  IV U62233 ( .A(n49479), .Z(n53434) );
  IV U62234 ( .A(n49480), .Z(n49646) );
  IV U62235 ( .A(n49481), .Z(n49482) );
  NOR U62236 ( .A(n49646), .B(n49482), .Z(n53267) );
  IV U62237 ( .A(n49483), .Z(n49484) );
  NOR U62238 ( .A(n49484), .B(n49486), .Z(n53426) );
  IV U62239 ( .A(n49485), .Z(n49489) );
  NOR U62240 ( .A(n49487), .B(n49486), .Z(n49488) );
  IV U62241 ( .A(n49488), .Z(n49494) );
  NOR U62242 ( .A(n49489), .B(n49494), .Z(n53272) );
  NOR U62243 ( .A(n53426), .B(n53272), .Z(n49643) );
  IV U62244 ( .A(n49490), .Z(n49492) );
  NOR U62245 ( .A(n49492), .B(n49491), .Z(n53277) );
  IV U62246 ( .A(n49493), .Z(n49495) );
  NOR U62247 ( .A(n49495), .B(n49494), .Z(n53270) );
  NOR U62248 ( .A(n53277), .B(n53270), .Z(n49642) );
  IV U62249 ( .A(n49496), .Z(n53286) );
  NOR U62250 ( .A(n49497), .B(n53286), .Z(n49501) );
  IV U62251 ( .A(n49498), .Z(n49499) );
  NOR U62252 ( .A(n49500), .B(n49499), .Z(n53280) );
  NOR U62253 ( .A(n49501), .B(n53280), .Z(n49641) );
  NOR U62254 ( .A(n49503), .B(n49502), .Z(n49639) );
  IV U62255 ( .A(n49639), .Z(n49637) );
  IV U62256 ( .A(n49504), .Z(n49505) );
  NOR U62257 ( .A(n49506), .B(n49505), .Z(n49507) );
  IV U62258 ( .A(n49507), .Z(n53409) );
  IV U62259 ( .A(n49508), .Z(n49509) );
  NOR U62260 ( .A(n49509), .B(n49512), .Z(n53393) );
  IV U62261 ( .A(n49510), .Z(n49511) );
  NOR U62262 ( .A(n49512), .B(n49511), .Z(n53301) );
  IV U62263 ( .A(n49513), .Z(n49514) );
  NOR U62264 ( .A(n49515), .B(n49514), .Z(n53304) );
  IV U62265 ( .A(n49516), .Z(n49517) );
  NOR U62266 ( .A(n53370), .B(n49517), .Z(n49615) );
  IV U62267 ( .A(n49518), .Z(n49520) );
  IV U62268 ( .A(n49519), .Z(n49524) );
  NOR U62269 ( .A(n49520), .B(n49524), .Z(n53362) );
  IV U62270 ( .A(n49521), .Z(n49522) );
  NOR U62271 ( .A(n49522), .B(n49524), .Z(n53359) );
  IV U62272 ( .A(n49523), .Z(n49525) );
  NOR U62273 ( .A(n49525), .B(n49524), .Z(n53311) );
  IV U62274 ( .A(n49526), .Z(n49527) );
  NOR U62275 ( .A(n49601), .B(n49527), .Z(n53308) );
  IV U62276 ( .A(n49528), .Z(n49530) );
  IV U62277 ( .A(n49529), .Z(n49602) );
  NOR U62278 ( .A(n49530), .B(n49602), .Z(n49609) );
  IV U62279 ( .A(n49609), .Z(n49598) );
  IV U62280 ( .A(n49531), .Z(n49532) );
  NOR U62281 ( .A(n49532), .B(n49578), .Z(n49595) );
  IV U62282 ( .A(n49595), .Z(n49576) );
  IV U62283 ( .A(n49533), .Z(n49582) );
  IV U62284 ( .A(n49534), .Z(n49535) );
  NOR U62285 ( .A(n49582), .B(n49535), .Z(n49536) );
  IV U62286 ( .A(n49536), .Z(n53355) );
  IV U62287 ( .A(n49537), .Z(n49538) );
  NOR U62288 ( .A(n49539), .B(n49538), .Z(n53324) );
  IV U62289 ( .A(n49540), .Z(n49541) );
  NOR U62290 ( .A(n49541), .B(n49559), .Z(n49542) );
  NOR U62291 ( .A(n49543), .B(n49542), .Z(n53332) );
  IV U62292 ( .A(n49544), .Z(n49545) );
  NOR U62293 ( .A(n49546), .B(n49545), .Z(n49551) );
  IV U62294 ( .A(n49547), .Z(n49549) );
  NOR U62295 ( .A(n49549), .B(n49548), .Z(n49550) );
  NOR U62296 ( .A(n49551), .B(n49550), .Z(n53333) );
  IV U62297 ( .A(n49552), .Z(n49554) );
  NOR U62298 ( .A(n49554), .B(n49553), .Z(n49564) );
  IV U62299 ( .A(n49555), .Z(n49556) );
  NOR U62300 ( .A(n49557), .B(n49556), .Z(n49562) );
  IV U62301 ( .A(n49558), .Z(n49560) );
  NOR U62302 ( .A(n49560), .B(n49559), .Z(n49561) );
  NOR U62303 ( .A(n49562), .B(n49561), .Z(n53334) );
  IV U62304 ( .A(n53334), .Z(n49563) );
  NOR U62305 ( .A(n49564), .B(n49563), .Z(n49565) );
  XOR U62306 ( .A(n53333), .B(n49565), .Z(n53330) );
  XOR U62307 ( .A(n53332), .B(n53330), .Z(n53338) );
  IV U62308 ( .A(n49566), .Z(n49567) );
  NOR U62309 ( .A(n49568), .B(n49567), .Z(n53337) );
  IV U62310 ( .A(n49569), .Z(n49570) );
  NOR U62311 ( .A(n49570), .B(n49574), .Z(n53328) );
  NOR U62312 ( .A(n53337), .B(n53328), .Z(n49571) );
  XOR U62313 ( .A(n53338), .B(n49571), .Z(n49572) );
  IV U62314 ( .A(n49572), .Z(n53342) );
  IV U62315 ( .A(n49573), .Z(n49575) );
  NOR U62316 ( .A(n49575), .B(n49574), .Z(n53340) );
  XOR U62317 ( .A(n53342), .B(n53340), .Z(n53326) );
  XOR U62318 ( .A(n53324), .B(n53326), .Z(n53354) );
  XOR U62319 ( .A(n53355), .B(n53354), .Z(n49583) );
  IV U62320 ( .A(n49583), .Z(n49586) );
  NOR U62321 ( .A(n49576), .B(n49586), .Z(n56742) );
  IV U62322 ( .A(n49577), .Z(n49579) );
  NOR U62323 ( .A(n49579), .B(n49578), .Z(n49592) );
  IV U62324 ( .A(n49592), .Z(n49584) );
  IV U62325 ( .A(n49580), .Z(n49581) );
  NOR U62326 ( .A(n49582), .B(n49581), .Z(n49585) );
  NOR U62327 ( .A(n49585), .B(n49583), .Z(n49590) );
  NOR U62328 ( .A(n49584), .B(n49590), .Z(n49589) );
  IV U62329 ( .A(n49585), .Z(n49587) );
  NOR U62330 ( .A(n49587), .B(n49586), .Z(n49588) );
  NOR U62331 ( .A(n49589), .B(n49588), .Z(n56741) );
  IV U62332 ( .A(n56741), .Z(n56744) );
  IV U62333 ( .A(n49590), .Z(n49591) );
  NOR U62334 ( .A(n49592), .B(n49591), .Z(n49593) );
  NOR U62335 ( .A(n56744), .B(n49593), .Z(n49594) );
  NOR U62336 ( .A(n49595), .B(n49594), .Z(n49596) );
  NOR U62337 ( .A(n56742), .B(n49596), .Z(n49597) );
  IV U62338 ( .A(n49597), .Z(n53318) );
  NOR U62339 ( .A(n49598), .B(n53318), .Z(n56756) );
  IV U62340 ( .A(n49599), .Z(n49600) );
  NOR U62341 ( .A(n49601), .B(n49600), .Z(n49610) );
  IV U62342 ( .A(n49610), .Z(n49607) );
  NOR U62343 ( .A(n49603), .B(n49602), .Z(n49604) );
  IV U62344 ( .A(n49604), .Z(n53317) );
  NOR U62345 ( .A(n53317), .B(n49605), .Z(n49606) );
  XOR U62346 ( .A(n49606), .B(n53318), .Z(n49608) );
  NOR U62347 ( .A(n49607), .B(n49608), .Z(n56757) );
  NOR U62348 ( .A(n56756), .B(n56757), .Z(n53358) );
  IV U62349 ( .A(n53358), .Z(n49611) );
  NOR U62350 ( .A(n49611), .B(n49608), .Z(n49614) );
  NOR U62351 ( .A(n49610), .B(n49609), .Z(n49612) );
  NOR U62352 ( .A(n49612), .B(n49611), .Z(n49613) );
  NOR U62353 ( .A(n49614), .B(n49613), .Z(n53310) );
  XOR U62354 ( .A(n53308), .B(n53310), .Z(n53312) );
  XOR U62355 ( .A(n53311), .B(n53312), .Z(n53361) );
  XOR U62356 ( .A(n53359), .B(n53361), .Z(n53364) );
  XOR U62357 ( .A(n53362), .B(n53364), .Z(n53369) );
  XOR U62358 ( .A(n49615), .B(n53369), .Z(n49623) );
  IV U62359 ( .A(n49616), .Z(n49617) );
  NOR U62360 ( .A(n53370), .B(n49617), .Z(n49627) );
  IV U62361 ( .A(n49627), .Z(n49618) );
  NOR U62362 ( .A(n49623), .B(n49618), .Z(n53389) );
  IV U62363 ( .A(n49619), .Z(n49621) );
  NOR U62364 ( .A(n49621), .B(n49620), .Z(n49625) );
  IV U62365 ( .A(n49625), .Z(n49622) );
  NOR U62366 ( .A(n49622), .B(n53369), .Z(n56708) );
  IV U62367 ( .A(n49623), .Z(n49624) );
  NOR U62368 ( .A(n49625), .B(n49624), .Z(n49626) );
  NOR U62369 ( .A(n56708), .B(n49626), .Z(n49628) );
  NOR U62370 ( .A(n49628), .B(n49627), .Z(n49629) );
  NOR U62371 ( .A(n53389), .B(n49629), .Z(n49630) );
  IV U62372 ( .A(n49630), .Z(n53305) );
  XOR U62373 ( .A(n53304), .B(n53305), .Z(n53302) );
  XOR U62374 ( .A(n53301), .B(n53302), .Z(n53394) );
  XOR U62375 ( .A(n53393), .B(n53394), .Z(n53408) );
  XOR U62376 ( .A(n53409), .B(n53408), .Z(n53298) );
  IV U62377 ( .A(n49631), .Z(n49632) );
  NOR U62378 ( .A(n49633), .B(n49632), .Z(n53297) );
  NOR U62379 ( .A(n49635), .B(n49634), .Z(n53404) );
  NOR U62380 ( .A(n53297), .B(n53404), .Z(n49636) );
  XOR U62381 ( .A(n53298), .B(n49636), .Z(n53290) );
  NOR U62382 ( .A(n49637), .B(n53290), .Z(n53424) );
  XOR U62383 ( .A(n53289), .B(n53290), .Z(n53293) );
  XOR U62384 ( .A(n53292), .B(n53293), .Z(n53285) );
  IV U62385 ( .A(n53285), .Z(n49638) );
  NOR U62386 ( .A(n49639), .B(n49638), .Z(n49640) );
  NOR U62387 ( .A(n53424), .B(n49640), .Z(n53281) );
  XOR U62388 ( .A(n49641), .B(n53281), .Z(n53279) );
  XOR U62389 ( .A(n49642), .B(n53279), .Z(n53273) );
  XOR U62390 ( .A(n49643), .B(n53273), .Z(n53269) );
  XOR U62391 ( .A(n53267), .B(n53269), .Z(n53432) );
  IV U62392 ( .A(n49644), .Z(n49645) );
  NOR U62393 ( .A(n49646), .B(n49645), .Z(n53430) );
  XOR U62394 ( .A(n53432), .B(n53430), .Z(n53433) );
  XOR U62395 ( .A(n53434), .B(n53433), .Z(n49647) );
  XOR U62396 ( .A(n49648), .B(n49647), .Z(n53444) );
  IV U62397 ( .A(n49649), .Z(n49651) );
  NOR U62398 ( .A(n49651), .B(n49650), .Z(n49652) );
  IV U62399 ( .A(n49652), .Z(n49659) );
  NOR U62400 ( .A(n53444), .B(n49659), .Z(n56688) );
  IV U62401 ( .A(n49653), .Z(n49655) );
  NOR U62402 ( .A(n49655), .B(n49654), .Z(n49656) );
  IV U62403 ( .A(n49656), .Z(n53261) );
  NOR U62404 ( .A(n49658), .B(n49657), .Z(n53442) );
  XOR U62405 ( .A(n53442), .B(n53444), .Z(n53260) );
  XOR U62406 ( .A(n53261), .B(n53260), .Z(n49662) );
  IV U62407 ( .A(n53260), .Z(n49660) );
  NOR U62408 ( .A(n49660), .B(n49659), .Z(n49661) );
  NOR U62409 ( .A(n49662), .B(n49661), .Z(n49663) );
  NOR U62410 ( .A(n56688), .B(n49663), .Z(n53258) );
  XOR U62411 ( .A(n53259), .B(n53258), .Z(n53451) );
  XOR U62412 ( .A(n49664), .B(n53451), .Z(n49665) );
  IV U62413 ( .A(n49665), .Z(n53257) );
  XOR U62414 ( .A(n53255), .B(n53257), .Z(n53251) );
  XOR U62415 ( .A(n49666), .B(n53251), .Z(n49676) );
  IV U62416 ( .A(n49676), .Z(n49671) );
  IV U62417 ( .A(n49667), .Z(n49669) );
  NOR U62418 ( .A(n49669), .B(n49668), .Z(n49680) );
  IV U62419 ( .A(n49680), .Z(n49670) );
  NOR U62420 ( .A(n49671), .B(n49670), .Z(n53457) );
  IV U62421 ( .A(n49672), .Z(n49674) );
  NOR U62422 ( .A(n49674), .B(n49673), .Z(n49677) );
  IV U62423 ( .A(n49677), .Z(n49675) );
  NOR U62424 ( .A(n49675), .B(n53251), .Z(n56856) );
  NOR U62425 ( .A(n49677), .B(n49676), .Z(n49678) );
  NOR U62426 ( .A(n56856), .B(n49678), .Z(n49679) );
  NOR U62427 ( .A(n49680), .B(n49679), .Z(n49681) );
  NOR U62428 ( .A(n53457), .B(n49681), .Z(n49682) );
  IV U62429 ( .A(n49682), .Z(n53454) );
  IV U62430 ( .A(n49683), .Z(n49685) );
  NOR U62431 ( .A(n49685), .B(n49684), .Z(n53453) );
  XOR U62432 ( .A(n53454), .B(n53453), .Z(n56870) );
  XOR U62433 ( .A(n56869), .B(n56870), .Z(n56872) );
  XOR U62434 ( .A(n56873), .B(n56872), .Z(n53462) );
  IV U62435 ( .A(n49686), .Z(n49688) );
  NOR U62436 ( .A(n49688), .B(n49687), .Z(n49689) );
  IV U62437 ( .A(n49689), .Z(n53463) );
  XOR U62438 ( .A(n53462), .B(n53463), .Z(n53248) );
  IV U62439 ( .A(n49690), .Z(n49691) );
  NOR U62440 ( .A(n49692), .B(n49691), .Z(n53247) );
  IV U62441 ( .A(n49693), .Z(n49695) );
  NOR U62442 ( .A(n49695), .B(n49694), .Z(n53245) );
  NOR U62443 ( .A(n53247), .B(n53245), .Z(n49696) );
  XOR U62444 ( .A(n53248), .B(n49696), .Z(n49704) );
  IV U62445 ( .A(n49704), .Z(n49697) );
  NOR U62446 ( .A(n49698), .B(n49697), .Z(n56893) );
  IV U62447 ( .A(n49699), .Z(n49701) );
  NOR U62448 ( .A(n49701), .B(n49700), .Z(n49705) );
  IV U62449 ( .A(n49705), .Z(n49703) );
  XOR U62450 ( .A(n53247), .B(n53248), .Z(n49702) );
  NOR U62451 ( .A(n49703), .B(n49702), .Z(n56672) );
  NOR U62452 ( .A(n49705), .B(n49704), .Z(n49706) );
  NOR U62453 ( .A(n56672), .B(n49706), .Z(n49707) );
  NOR U62454 ( .A(n49708), .B(n49707), .Z(n49709) );
  NOR U62455 ( .A(n56893), .B(n49709), .Z(n49710) );
  IV U62456 ( .A(n49710), .Z(n53471) );
  XOR U62457 ( .A(n53470), .B(n53471), .Z(n53244) );
  IV U62458 ( .A(n53244), .Z(n49718) );
  IV U62459 ( .A(n49711), .Z(n49712) );
  NOR U62460 ( .A(n49713), .B(n49712), .Z(n53240) );
  IV U62461 ( .A(n49714), .Z(n49716) );
  NOR U62462 ( .A(n49716), .B(n49715), .Z(n53242) );
  NOR U62463 ( .A(n53240), .B(n53242), .Z(n49717) );
  XOR U62464 ( .A(n49718), .B(n49717), .Z(n53238) );
  XOR U62465 ( .A(n53237), .B(n53238), .Z(n53476) );
  XOR U62466 ( .A(n53475), .B(n53476), .Z(n53479) );
  XOR U62467 ( .A(n49719), .B(n53479), .Z(n53232) );
  NOR U62468 ( .A(n49721), .B(n49720), .Z(n49722) );
  IV U62469 ( .A(n49722), .Z(n49723) );
  NOR U62470 ( .A(n49724), .B(n49723), .Z(n49725) );
  IV U62471 ( .A(n49725), .Z(n53233) );
  XOR U62472 ( .A(n53232), .B(n53233), .Z(n53229) );
  IV U62473 ( .A(n49726), .Z(n49727) );
  NOR U62474 ( .A(n49727), .B(n49730), .Z(n53227) );
  XOR U62475 ( .A(n53229), .B(n53227), .Z(n53223) );
  XOR U62476 ( .A(n53220), .B(n53223), .Z(n53219) );
  IV U62477 ( .A(n53219), .Z(n49739) );
  IV U62478 ( .A(n49728), .Z(n49729) );
  NOR U62479 ( .A(n49730), .B(n49729), .Z(n53225) );
  IV U62480 ( .A(n49731), .Z(n49732) );
  NOR U62481 ( .A(n49733), .B(n49732), .Z(n53222) );
  IV U62482 ( .A(n49734), .Z(n49735) );
  NOR U62483 ( .A(n49735), .B(n49742), .Z(n53217) );
  NOR U62484 ( .A(n53222), .B(n53217), .Z(n49736) );
  IV U62485 ( .A(n49736), .Z(n49737) );
  NOR U62486 ( .A(n53225), .B(n49737), .Z(n49738) );
  XOR U62487 ( .A(n49739), .B(n49738), .Z(n53213) );
  IV U62488 ( .A(n49740), .Z(n49741) );
  NOR U62489 ( .A(n49742), .B(n49741), .Z(n53211) );
  XOR U62490 ( .A(n53213), .B(n53211), .Z(n53215) );
  XOR U62491 ( .A(n53214), .B(n53215), .Z(n53205) );
  XOR U62492 ( .A(n53203), .B(n53205), .Z(n53207) );
  XOR U62493 ( .A(n53206), .B(n53207), .Z(n49743) );
  XOR U62494 ( .A(n49744), .B(n49743), .Z(n49745) );
  IV U62495 ( .A(n49745), .Z(n53198) );
  XOR U62496 ( .A(n53196), .B(n53198), .Z(n53487) );
  IV U62497 ( .A(n49746), .Z(n49747) );
  NOR U62498 ( .A(n49750), .B(n49747), .Z(n53485) );
  XOR U62499 ( .A(n53487), .B(n53485), .Z(n53195) );
  IV U62500 ( .A(n49748), .Z(n49749) );
  NOR U62501 ( .A(n49750), .B(n49749), .Z(n53193) );
  XOR U62502 ( .A(n53195), .B(n53193), .Z(n53493) );
  XOR U62503 ( .A(n53492), .B(n53493), .Z(n53496) );
  XOR U62504 ( .A(n53495), .B(n53496), .Z(n53501) );
  IV U62505 ( .A(n49751), .Z(n49753) );
  NOR U62506 ( .A(n49753), .B(n49752), .Z(n53499) );
  XOR U62507 ( .A(n53501), .B(n53499), .Z(n53508) );
  XOR U62508 ( .A(n53502), .B(n53508), .Z(n53191) );
  XOR U62509 ( .A(n53192), .B(n53191), .Z(n49754) );
  XOR U62510 ( .A(n49755), .B(n49754), .Z(n53184) );
  IV U62511 ( .A(n49756), .Z(n49758) );
  NOR U62512 ( .A(n49758), .B(n49757), .Z(n53182) );
  XOR U62513 ( .A(n53184), .B(n53182), .Z(n53185) );
  XOR U62514 ( .A(n53186), .B(n53185), .Z(n53175) );
  XOR U62515 ( .A(n53177), .B(n53175), .Z(n53510) );
  XOR U62516 ( .A(n49759), .B(n53510), .Z(n49760) );
  IV U62517 ( .A(n49760), .Z(n53514) );
  XOR U62518 ( .A(n53512), .B(n53514), .Z(n53522) );
  XOR U62519 ( .A(n53515), .B(n53522), .Z(n53172) );
  XOR U62520 ( .A(n53171), .B(n53172), .Z(n53169) );
  IV U62521 ( .A(n49761), .Z(n49762) );
  NOR U62522 ( .A(n49763), .B(n49762), .Z(n49764) );
  IV U62523 ( .A(n49764), .Z(n53167) );
  XOR U62524 ( .A(n53169), .B(n53167), .Z(n49765) );
  XOR U62525 ( .A(n49766), .B(n49765), .Z(n53161) );
  XOR U62526 ( .A(n53159), .B(n53161), .Z(n53163) );
  XOR U62527 ( .A(n53162), .B(n53163), .Z(n53158) );
  XOR U62528 ( .A(n53157), .B(n53158), .Z(n53539) );
  XOR U62529 ( .A(n53538), .B(n53539), .Z(n53536) );
  XOR U62530 ( .A(n49767), .B(n53536), .Z(n49772) );
  IV U62531 ( .A(n49773), .Z(n49771) );
  NOR U62532 ( .A(n49772), .B(n49771), .Z(n53551) );
  IV U62533 ( .A(n49772), .Z(n49774) );
  NOR U62534 ( .A(n49774), .B(n49773), .Z(n56629) );
  NOR U62535 ( .A(n53551), .B(n56629), .Z(n56625) );
  IV U62536 ( .A(n49775), .Z(n49777) );
  NOR U62537 ( .A(n49777), .B(n49776), .Z(n53548) );
  NOR U62538 ( .A(n53547), .B(n53548), .Z(n56627) );
  XOR U62539 ( .A(n56625), .B(n56627), .Z(n53149) );
  XOR U62540 ( .A(n53148), .B(n53149), .Z(n53153) );
  XOR U62541 ( .A(n53151), .B(n53153), .Z(n53156) );
  XOR U62542 ( .A(n53154), .B(n53156), .Z(n53146) );
  XOR U62543 ( .A(n49778), .B(n53146), .Z(n53137) );
  XOR U62544 ( .A(n49779), .B(n53137), .Z(n56596) );
  XOR U62545 ( .A(n53562), .B(n56596), .Z(n53132) );
  XOR U62546 ( .A(n53131), .B(n53132), .Z(n57034) );
  XOR U62547 ( .A(n49780), .B(n57034), .Z(n53569) );
  XOR U62548 ( .A(n49781), .B(n53569), .Z(n53129) );
  XOR U62549 ( .A(n53127), .B(n53129), .Z(n53123) );
  NOR U62550 ( .A(n49782), .B(n53123), .Z(n53126) );
  XOR U62551 ( .A(n53122), .B(n53123), .Z(n53119) );
  IV U62552 ( .A(n53119), .Z(n49783) );
  NOR U62553 ( .A(n49784), .B(n49783), .Z(n49785) );
  NOR U62554 ( .A(n53126), .B(n49785), .Z(n49790) );
  IV U62555 ( .A(n49786), .Z(n49788) );
  NOR U62556 ( .A(n49788), .B(n49787), .Z(n53116) );
  NOR U62557 ( .A(n53118), .B(n53116), .Z(n49789) );
  XOR U62558 ( .A(n49790), .B(n49789), .Z(n53111) );
  IV U62559 ( .A(n49791), .Z(n49794) );
  IV U62560 ( .A(n49792), .Z(n49793) );
  NOR U62561 ( .A(n49794), .B(n49793), .Z(n53109) );
  XOR U62562 ( .A(n53111), .B(n53109), .Z(n53112) );
  XOR U62563 ( .A(n53113), .B(n53112), .Z(n53102) );
  XOR U62564 ( .A(n53101), .B(n53102), .Z(n53098) );
  XOR U62565 ( .A(n49795), .B(n53098), .Z(n53570) );
  XOR U62566 ( .A(n53572), .B(n53570), .Z(n53578) );
  XOR U62567 ( .A(n53573), .B(n53578), .Z(n53593) );
  XOR U62568 ( .A(n49796), .B(n53593), .Z(n49797) );
  IV U62569 ( .A(n49797), .Z(n53590) );
  XOR U62570 ( .A(n53588), .B(n53590), .Z(n53598) );
  IV U62571 ( .A(n49798), .Z(n49800) );
  NOR U62572 ( .A(n49800), .B(n49799), .Z(n53596) );
  XOR U62573 ( .A(n53598), .B(n53596), .Z(n53600) );
  XOR U62574 ( .A(n53599), .B(n53600), .Z(n53094) );
  IV U62575 ( .A(n49801), .Z(n49802) );
  NOR U62576 ( .A(n49803), .B(n49802), .Z(n53090) );
  IV U62577 ( .A(n49804), .Z(n49806) );
  NOR U62578 ( .A(n49806), .B(n49805), .Z(n53092) );
  NOR U62579 ( .A(n53090), .B(n53092), .Z(n49807) );
  XOR U62580 ( .A(n53094), .B(n49807), .Z(n53082) );
  XOR U62581 ( .A(n49808), .B(n53082), .Z(n53080) );
  XOR U62582 ( .A(n49809), .B(n53080), .Z(n53072) );
  XOR U62583 ( .A(n53073), .B(n53072), .Z(n53077) );
  NOR U62584 ( .A(n49810), .B(n53077), .Z(n57125) );
  NOR U62585 ( .A(n57125), .B(n49810), .Z(n49813) );
  IV U62586 ( .A(n49811), .Z(n49812) );
  NOR U62587 ( .A(n49812), .B(n53067), .Z(n49819) );
  NOR U62588 ( .A(n49813), .B(n49819), .Z(n49818) );
  IV U62589 ( .A(n49814), .Z(n49815) );
  NOR U62590 ( .A(n49816), .B(n49815), .Z(n53075) );
  XOR U62591 ( .A(n53077), .B(n53075), .Z(n53070) );
  IV U62592 ( .A(n53070), .Z(n49817) );
  NOR U62593 ( .A(n49818), .B(n49817), .Z(n49823) );
  NOR U62594 ( .A(n57125), .B(n49819), .Z(n49820) );
  IV U62595 ( .A(n49820), .Z(n49821) );
  NOR U62596 ( .A(n53070), .B(n49821), .Z(n49822) );
  NOR U62597 ( .A(n49823), .B(n49822), .Z(n53062) );
  IV U62598 ( .A(n49824), .Z(n53066) );
  IV U62599 ( .A(n49825), .Z(n49826) );
  NOR U62600 ( .A(n53066), .B(n49826), .Z(n49827) );
  IV U62601 ( .A(n49827), .Z(n53060) );
  XOR U62602 ( .A(n53062), .B(n53060), .Z(n49828) );
  XOR U62603 ( .A(n49829), .B(n49828), .Z(n53054) );
  IV U62604 ( .A(n49830), .Z(n49831) );
  NOR U62605 ( .A(n49832), .B(n49831), .Z(n53056) );
  IV U62606 ( .A(n49833), .Z(n49835) );
  NOR U62607 ( .A(n49835), .B(n49834), .Z(n53053) );
  NOR U62608 ( .A(n53056), .B(n53053), .Z(n49836) );
  XOR U62609 ( .A(n53054), .B(n49836), .Z(n53052) );
  XOR U62610 ( .A(n53050), .B(n53052), .Z(n53614) );
  XOR U62611 ( .A(n53615), .B(n53614), .Z(n53048) );
  IV U62612 ( .A(n49837), .Z(n49838) );
  NOR U62613 ( .A(n49839), .B(n49838), .Z(n53047) );
  IV U62614 ( .A(n49840), .Z(n49842) );
  NOR U62615 ( .A(n49842), .B(n49841), .Z(n53616) );
  NOR U62616 ( .A(n53047), .B(n53616), .Z(n49843) );
  XOR U62617 ( .A(n53048), .B(n49843), .Z(n53045) );
  XOR U62618 ( .A(n53044), .B(n53045), .Z(n53623) );
  XOR U62619 ( .A(n53621), .B(n53623), .Z(n53625) );
  XOR U62620 ( .A(n53624), .B(n53625), .Z(n53629) );
  XOR U62621 ( .A(n53628), .B(n53629), .Z(n53042) );
  XOR U62622 ( .A(n49844), .B(n53042), .Z(n53032) );
  XOR U62623 ( .A(n49845), .B(n53032), .Z(n53028) );
  XOR U62624 ( .A(n49846), .B(n53028), .Z(n53641) );
  XOR U62625 ( .A(n49847), .B(n53641), .Z(n49848) );
  IV U62626 ( .A(n49848), .Z(n53024) );
  IV U62627 ( .A(n49849), .Z(n49852) );
  NOR U62628 ( .A(n53024), .B(n49852), .Z(n49850) );
  IV U62629 ( .A(n49850), .Z(n49859) );
  NOR U62630 ( .A(n49851), .B(n49859), .Z(n53646) );
  NOR U62631 ( .A(n49853), .B(n49852), .Z(n49857) );
  NOR U62632 ( .A(n49854), .B(n53023), .Z(n49855) );
  XOR U62633 ( .A(n53024), .B(n49855), .Z(n49874) );
  IV U62634 ( .A(n49874), .Z(n49856) );
  NOR U62635 ( .A(n49857), .B(n49856), .Z(n49861) );
  IV U62636 ( .A(n49858), .Z(n49860) );
  NOR U62637 ( .A(n49860), .B(n49859), .Z(n53021) );
  NOR U62638 ( .A(n49861), .B(n53021), .Z(n49862) );
  IV U62639 ( .A(n49862), .Z(n49863) );
  NOR U62640 ( .A(n53646), .B(n49863), .Z(n49864) );
  NOR U62641 ( .A(n49873), .B(n49864), .Z(n49876) );
  IV U62642 ( .A(n49865), .Z(n49871) );
  NOR U62643 ( .A(n49876), .B(n49871), .Z(n49866) );
  IV U62644 ( .A(n49866), .Z(n49869) );
  NOR U62645 ( .A(n49867), .B(n49869), .Z(n53652) );
  IV U62646 ( .A(n49868), .Z(n49870) );
  NOR U62647 ( .A(n49870), .B(n49869), .Z(n57188) );
  NOR U62648 ( .A(n49872), .B(n49871), .Z(n49878) );
  IV U62649 ( .A(n49873), .Z(n49875) );
  NOR U62650 ( .A(n49875), .B(n49874), .Z(n53020) );
  NOR U62651 ( .A(n49876), .B(n53020), .Z(n49877) );
  NOR U62652 ( .A(n49878), .B(n49877), .Z(n49879) );
  NOR U62653 ( .A(n57188), .B(n49879), .Z(n49880) );
  IV U62654 ( .A(n49880), .Z(n53649) );
  NOR U62655 ( .A(n53652), .B(n53649), .Z(n53017) );
  XOR U62656 ( .A(n49881), .B(n53017), .Z(n53655) );
  XOR U62657 ( .A(n53653), .B(n53655), .Z(n53656) );
  XOR U62658 ( .A(n53657), .B(n53656), .Z(n53012) );
  XOR U62659 ( .A(n49882), .B(n53012), .Z(n53667) );
  XOR U62660 ( .A(n53665), .B(n53667), .Z(n53680) );
  IV U62661 ( .A(n49883), .Z(n49885) );
  NOR U62662 ( .A(n49885), .B(n49884), .Z(n53008) );
  IV U62663 ( .A(n49886), .Z(n49888) );
  NOR U62664 ( .A(n49888), .B(n49887), .Z(n53679) );
  NOR U62665 ( .A(n53008), .B(n53679), .Z(n49889) );
  XOR U62666 ( .A(n53680), .B(n49889), .Z(n53005) );
  XOR U62667 ( .A(n49890), .B(n53005), .Z(n53002) );
  NOR U62668 ( .A(n49891), .B(n53002), .Z(n57255) );
  IV U62669 ( .A(n49892), .Z(n49893) );
  NOR U62670 ( .A(n49894), .B(n49893), .Z(n53001) );
  XOR U62671 ( .A(n53001), .B(n53002), .Z(n49900) );
  IV U62672 ( .A(n49900), .Z(n49895) );
  NOR U62673 ( .A(n49896), .B(n49895), .Z(n49897) );
  NOR U62674 ( .A(n57255), .B(n49897), .Z(n49898) );
  NOR U62675 ( .A(n49899), .B(n49898), .Z(n49902) );
  IV U62676 ( .A(n49899), .Z(n49901) );
  NOR U62677 ( .A(n49901), .B(n49900), .Z(n52999) );
  NOR U62678 ( .A(n49902), .B(n52999), .Z(n49903) );
  IV U62679 ( .A(n49903), .Z(n52997) );
  IV U62680 ( .A(n49904), .Z(n49906) );
  NOR U62681 ( .A(n49906), .B(n49905), .Z(n52996) );
  XOR U62682 ( .A(n52997), .B(n52996), .Z(n53690) );
  XOR U62683 ( .A(n53689), .B(n53690), .Z(n52990) );
  XOR U62684 ( .A(n52989), .B(n52990), .Z(n53694) );
  XOR U62685 ( .A(n52992), .B(n53694), .Z(n52988) );
  XOR U62686 ( .A(n52986), .B(n52988), .Z(n52981) );
  XOR U62687 ( .A(n52980), .B(n52981), .Z(n53700) );
  XOR U62688 ( .A(n52970), .B(n53700), .Z(n49913) );
  NOR U62689 ( .A(n49907), .B(n52973), .Z(n49911) );
  IV U62690 ( .A(n49908), .Z(n49909) );
  NOR U62691 ( .A(n49910), .B(n49909), .Z(n53699) );
  NOR U62692 ( .A(n49911), .B(n53699), .Z(n49912) );
  XOR U62693 ( .A(n49913), .B(n49912), .Z(n52960) );
  XOR U62694 ( .A(n49914), .B(n52960), .Z(n52964) );
  XOR U62695 ( .A(n52963), .B(n52964), .Z(n52957) );
  XOR U62696 ( .A(n52955), .B(n52957), .Z(n53704) );
  XOR U62697 ( .A(n49915), .B(n53704), .Z(n49916) );
  IV U62698 ( .A(n49916), .Z(n52947) );
  XOR U62699 ( .A(n52945), .B(n52947), .Z(n52948) );
  XOR U62700 ( .A(n52949), .B(n52948), .Z(n49917) );
  IV U62701 ( .A(n49917), .Z(n52938) );
  NOR U62702 ( .A(n49923), .B(n52938), .Z(n56486) );
  NOR U62703 ( .A(n49919), .B(n49918), .Z(n49920) );
  IV U62704 ( .A(n49920), .Z(n52931) );
  NOR U62705 ( .A(n49921), .B(n52939), .Z(n49922) );
  XOR U62706 ( .A(n49922), .B(n52938), .Z(n52930) );
  XOR U62707 ( .A(n52931), .B(n52930), .Z(n49926) );
  IV U62708 ( .A(n52930), .Z(n49924) );
  NOR U62709 ( .A(n49924), .B(n49923), .Z(n49925) );
  NOR U62710 ( .A(n49926), .B(n49925), .Z(n49927) );
  NOR U62711 ( .A(n56486), .B(n49927), .Z(n49928) );
  IV U62712 ( .A(n49928), .Z(n52933) );
  XOR U62713 ( .A(n52933), .B(n52932), .Z(n53719) );
  XOR U62714 ( .A(n49929), .B(n53719), .Z(n49930) );
  IV U62715 ( .A(n49930), .Z(n52925) );
  XOR U62716 ( .A(n49931), .B(n52925), .Z(n53734) );
  XOR U62717 ( .A(n49932), .B(n53734), .Z(n49950) );
  IV U62718 ( .A(n49950), .Z(n53736) );
  NOR U62719 ( .A(n49945), .B(n53736), .Z(n57342) );
  NOR U62720 ( .A(n49934), .B(n49933), .Z(n49935) );
  IV U62721 ( .A(n49935), .Z(n49942) );
  XOR U62722 ( .A(n49937), .B(n49936), .Z(n49938) );
  NOR U62723 ( .A(n49939), .B(n49938), .Z(n49940) );
  IV U62724 ( .A(n49940), .Z(n49941) );
  NOR U62725 ( .A(n49942), .B(n49941), .Z(n53741) );
  NOR U62726 ( .A(n57342), .B(n53741), .Z(n49943) );
  IV U62727 ( .A(n49943), .Z(n49944) );
  NOR U62728 ( .A(n49945), .B(n49944), .Z(n49953) );
  IV U62729 ( .A(n49946), .Z(n49947) );
  NOR U62730 ( .A(n49948), .B(n49947), .Z(n49949) );
  IV U62731 ( .A(n49949), .Z(n53735) );
  XOR U62732 ( .A(n53735), .B(n49950), .Z(n53742) );
  XOR U62733 ( .A(n53741), .B(n53742), .Z(n49951) );
  NOR U62734 ( .A(n57342), .B(n49951), .Z(n49952) );
  NOR U62735 ( .A(n49953), .B(n49952), .Z(n53745) );
  XOR U62736 ( .A(n49954), .B(n53745), .Z(n49955) );
  IV U62737 ( .A(n49955), .Z(n52918) );
  XOR U62738 ( .A(n52917), .B(n52918), .Z(n52912) );
  IV U62739 ( .A(n52912), .Z(n49964) );
  IV U62740 ( .A(n49956), .Z(n49957) );
  NOR U62741 ( .A(n49958), .B(n49957), .Z(n49963) );
  IV U62742 ( .A(n49959), .Z(n49961) );
  NOR U62743 ( .A(n49961), .B(n49960), .Z(n49962) );
  NOR U62744 ( .A(n49963), .B(n49962), .Z(n52913) );
  XOR U62745 ( .A(n49964), .B(n52913), .Z(n52915) );
  XOR U62746 ( .A(n49965), .B(n52915), .Z(n52899) );
  IV U62747 ( .A(n52899), .Z(n52902) );
  XOR U62748 ( .A(n52900), .B(n52902), .Z(n52897) );
  IV U62749 ( .A(n49966), .Z(n49967) );
  NOR U62750 ( .A(n49968), .B(n49967), .Z(n52904) );
  IV U62751 ( .A(n49969), .Z(n49970) );
  NOR U62752 ( .A(n49971), .B(n49970), .Z(n52896) );
  NOR U62753 ( .A(n52904), .B(n52896), .Z(n49972) );
  XOR U62754 ( .A(n52897), .B(n49972), .Z(n49984) );
  IV U62755 ( .A(n49984), .Z(n52895) );
  IV U62756 ( .A(n49986), .Z(n49973) );
  NOR U62757 ( .A(n52895), .B(n49973), .Z(n57385) );
  NOR U62758 ( .A(n49975), .B(n49974), .Z(n49976) );
  IV U62759 ( .A(n49976), .Z(n52888) );
  IV U62760 ( .A(n49977), .Z(n49979) );
  NOR U62761 ( .A(n49979), .B(n49978), .Z(n52893) );
  IV U62762 ( .A(n49980), .Z(n49982) );
  NOR U62763 ( .A(n49982), .B(n49981), .Z(n52891) );
  NOR U62764 ( .A(n52893), .B(n52891), .Z(n49983) );
  XOR U62765 ( .A(n49984), .B(n49983), .Z(n52887) );
  XOR U62766 ( .A(n52888), .B(n52887), .Z(n49985) );
  NOR U62767 ( .A(n49986), .B(n49985), .Z(n49987) );
  NOR U62768 ( .A(n57385), .B(n49987), .Z(n52883) );
  IV U62769 ( .A(n49988), .Z(n49990) );
  NOR U62770 ( .A(n49990), .B(n49989), .Z(n52884) );
  XOR U62771 ( .A(n52883), .B(n52884), .Z(n52877) );
  XOR U62772 ( .A(n52874), .B(n52877), .Z(n52873) );
  XOR U62773 ( .A(n52871), .B(n52873), .Z(n50002) );
  IV U62774 ( .A(n49991), .Z(n49992) );
  NOR U62775 ( .A(n49993), .B(n49992), .Z(n49994) );
  IV U62776 ( .A(n49994), .Z(n50003) );
  NOR U62777 ( .A(n50002), .B(n50003), .Z(n57430) );
  IV U62778 ( .A(n49995), .Z(n49997) );
  NOR U62779 ( .A(n49997), .B(n49996), .Z(n49998) );
  IV U62780 ( .A(n49998), .Z(n52870) );
  IV U62781 ( .A(n49999), .Z(n50000) );
  NOR U62782 ( .A(n50001), .B(n50000), .Z(n52878) );
  XOR U62783 ( .A(n52878), .B(n50002), .Z(n52869) );
  XOR U62784 ( .A(n52870), .B(n52869), .Z(n50006) );
  IV U62785 ( .A(n52869), .Z(n50004) );
  NOR U62786 ( .A(n50004), .B(n50003), .Z(n50005) );
  NOR U62787 ( .A(n50006), .B(n50005), .Z(n50007) );
  NOR U62788 ( .A(n57430), .B(n50007), .Z(n53754) );
  XOR U62789 ( .A(n50008), .B(n53754), .Z(n52864) );
  XOR U62790 ( .A(n52862), .B(n52864), .Z(n52859) );
  IV U62791 ( .A(n52859), .Z(n50013) );
  IV U62792 ( .A(n50009), .Z(n50011) );
  NOR U62793 ( .A(n50011), .B(n50010), .Z(n52858) );
  NOR U62794 ( .A(n52866), .B(n52858), .Z(n50012) );
  XOR U62795 ( .A(n50013), .B(n50012), .Z(n52857) );
  XOR U62796 ( .A(n52855), .B(n52857), .Z(n50016) );
  NOR U62797 ( .A(n50016), .B(n50014), .Z(n50015) );
  IV U62798 ( .A(n50015), .Z(n52852) );
  NOR U62799 ( .A(n50017), .B(n52852), .Z(n57417) );
  IV U62800 ( .A(n50016), .Z(n50019) );
  IV U62801 ( .A(n50024), .Z(n50021) );
  NOR U62802 ( .A(n50017), .B(n50021), .Z(n50018) );
  NOR U62803 ( .A(n50019), .B(n50018), .Z(n50020) );
  NOR U62804 ( .A(n57417), .B(n50020), .Z(n50029) );
  NOR U62805 ( .A(n50022), .B(n50021), .Z(n52854) );
  IV U62806 ( .A(n50023), .Z(n52853) );
  NOR U62807 ( .A(n50025), .B(n50024), .Z(n50026) );
  NOR U62808 ( .A(n52853), .B(n50026), .Z(n50027) );
  NOR U62809 ( .A(n52854), .B(n50027), .Z(n50028) );
  XOR U62810 ( .A(n50029), .B(n50028), .Z(n53765) );
  IV U62811 ( .A(n50030), .Z(n52845) );
  NOR U62812 ( .A(n52845), .B(n50031), .Z(n50035) );
  IV U62813 ( .A(n50032), .Z(n50034) );
  NOR U62814 ( .A(n50034), .B(n50033), .Z(n53763) );
  NOR U62815 ( .A(n50035), .B(n53763), .Z(n50036) );
  XOR U62816 ( .A(n53765), .B(n50036), .Z(n50037) );
  IV U62817 ( .A(n50037), .Z(n53761) );
  XOR U62818 ( .A(n53762), .B(n53761), .Z(n52838) );
  IV U62819 ( .A(n50038), .Z(n50039) );
  NOR U62820 ( .A(n50040), .B(n50039), .Z(n52841) );
  IV U62821 ( .A(n50041), .Z(n50042) );
  NOR U62822 ( .A(n50042), .B(n50048), .Z(n52839) );
  NOR U62823 ( .A(n52841), .B(n52839), .Z(n50043) );
  XOR U62824 ( .A(n52838), .B(n50043), .Z(n52837) );
  NOR U62825 ( .A(n50045), .B(n50044), .Z(n50051) );
  IV U62826 ( .A(n50051), .Z(n50046) );
  NOR U62827 ( .A(n52837), .B(n50046), .Z(n52834) );
  IV U62828 ( .A(n50047), .Z(n50049) );
  NOR U62829 ( .A(n50049), .B(n50048), .Z(n52835) );
  XOR U62830 ( .A(n52835), .B(n52837), .Z(n53769) );
  IV U62831 ( .A(n53769), .Z(n50050) );
  NOR U62832 ( .A(n50051), .B(n50050), .Z(n50052) );
  NOR U62833 ( .A(n52834), .B(n50052), .Z(n50053) );
  IV U62834 ( .A(n50053), .Z(n52832) );
  XOR U62835 ( .A(n52833), .B(n52832), .Z(n52826) );
  NOR U62836 ( .A(n50055), .B(n50054), .Z(n53768) );
  NOR U62837 ( .A(n52827), .B(n53768), .Z(n50056) );
  XOR U62838 ( .A(n52826), .B(n50056), .Z(n52825) );
  IV U62839 ( .A(n50057), .Z(n50058) );
  NOR U62840 ( .A(n50059), .B(n50058), .Z(n50060) );
  IV U62841 ( .A(n50060), .Z(n50070) );
  NOR U62842 ( .A(n52825), .B(n50070), .Z(n53783) );
  IV U62843 ( .A(n50061), .Z(n50062) );
  NOR U62844 ( .A(n50062), .B(n50077), .Z(n50063) );
  IV U62845 ( .A(n50063), .Z(n53790) );
  IV U62846 ( .A(n50064), .Z(n50068) );
  IV U62847 ( .A(n50065), .Z(n50066) );
  NOR U62848 ( .A(n50068), .B(n50066), .Z(n53780) );
  IV U62849 ( .A(n50067), .Z(n50069) );
  NOR U62850 ( .A(n50069), .B(n50068), .Z(n52823) );
  XOR U62851 ( .A(n52823), .B(n52825), .Z(n53781) );
  XOR U62852 ( .A(n53780), .B(n53781), .Z(n53789) );
  XOR U62853 ( .A(n53790), .B(n53789), .Z(n50073) );
  IV U62854 ( .A(n53789), .Z(n50071) );
  NOR U62855 ( .A(n50071), .B(n50070), .Z(n50072) );
  NOR U62856 ( .A(n50073), .B(n50072), .Z(n50074) );
  NOR U62857 ( .A(n53783), .B(n50074), .Z(n50075) );
  IV U62858 ( .A(n50075), .Z(n52821) );
  IV U62859 ( .A(n50076), .Z(n50078) );
  NOR U62860 ( .A(n50078), .B(n50077), .Z(n52819) );
  XOR U62861 ( .A(n52821), .B(n52819), .Z(n53787) );
  XOR U62862 ( .A(n53785), .B(n53787), .Z(n53798) );
  XOR U62863 ( .A(n53796), .B(n53798), .Z(n53801) );
  XOR U62864 ( .A(n53799), .B(n53801), .Z(n52817) );
  XOR U62865 ( .A(n52812), .B(n52817), .Z(n50079) );
  XOR U62866 ( .A(n50080), .B(n50079), .Z(n50081) );
  IV U62867 ( .A(n50081), .Z(n53814) );
  XOR U62868 ( .A(n53811), .B(n53814), .Z(n53817) );
  XOR U62869 ( .A(n50082), .B(n53817), .Z(n53818) );
  XOR U62870 ( .A(n53819), .B(n53818), .Z(n53823) );
  XOR U62871 ( .A(n50083), .B(n53823), .Z(n50084) );
  IV U62872 ( .A(n50084), .Z(n52808) );
  XOR U62873 ( .A(n52809), .B(n52808), .Z(n50085) );
  NOR U62874 ( .A(n50086), .B(n50085), .Z(n50089) );
  IV U62875 ( .A(n50086), .Z(n50088) );
  XOR U62876 ( .A(n53821), .B(n53823), .Z(n50087) );
  NOR U62877 ( .A(n50088), .B(n50087), .Z(n56430) );
  NOR U62878 ( .A(n50089), .B(n56430), .Z(n50090) );
  IV U62879 ( .A(n50090), .Z(n53828) );
  NOR U62880 ( .A(n50091), .B(n50100), .Z(n50093) );
  NOR U62881 ( .A(n50092), .B(n50093), .Z(n50110) );
  IV U62882 ( .A(n50093), .Z(n50094) );
  NOR U62883 ( .A(n50095), .B(n50094), .Z(n50108) );
  NOR U62884 ( .A(n50097), .B(n50096), .Z(n50098) );
  IV U62885 ( .A(n50098), .Z(n50103) );
  NOR U62886 ( .A(n50100), .B(n50099), .Z(n50101) );
  IV U62887 ( .A(n50101), .Z(n50102) );
  NOR U62888 ( .A(n50103), .B(n50102), .Z(n50104) );
  IV U62889 ( .A(n50104), .Z(n50106) );
  NOR U62890 ( .A(n50106), .B(n50105), .Z(n50107) );
  NOR U62891 ( .A(n50108), .B(n50107), .Z(n50109) );
  NOR U62892 ( .A(n50110), .B(n50109), .Z(n53826) );
  XOR U62893 ( .A(n53828), .B(n53826), .Z(n52805) );
  XOR U62894 ( .A(n52803), .B(n52805), .Z(n53833) );
  XOR U62895 ( .A(n53831), .B(n53833), .Z(n53839) );
  IV U62896 ( .A(n50111), .Z(n50113) );
  NOR U62897 ( .A(n50113), .B(n50112), .Z(n52801) );
  XOR U62898 ( .A(n53839), .B(n52801), .Z(n50114) );
  XOR U62899 ( .A(n50115), .B(n50114), .Z(n50116) );
  IV U62900 ( .A(n50116), .Z(n52800) );
  IV U62901 ( .A(n50117), .Z(n50119) );
  NOR U62902 ( .A(n50119), .B(n50118), .Z(n50125) );
  IV U62903 ( .A(n50125), .Z(n50120) );
  NOR U62904 ( .A(n52800), .B(n50120), .Z(n56372) );
  IV U62905 ( .A(n50121), .Z(n50122) );
  NOR U62906 ( .A(n50123), .B(n50122), .Z(n52798) );
  XOR U62907 ( .A(n52798), .B(n52800), .Z(n50129) );
  IV U62908 ( .A(n50129), .Z(n50124) );
  NOR U62909 ( .A(n50125), .B(n50124), .Z(n50126) );
  NOR U62910 ( .A(n56372), .B(n50126), .Z(n50127) );
  NOR U62911 ( .A(n50128), .B(n50127), .Z(n50131) );
  IV U62912 ( .A(n50128), .Z(n50130) );
  NOR U62913 ( .A(n50130), .B(n50129), .Z(n56375) );
  NOR U62914 ( .A(n50131), .B(n56375), .Z(n53841) );
  IV U62915 ( .A(n50132), .Z(n50133) );
  NOR U62916 ( .A(n50133), .B(n50139), .Z(n50134) );
  IV U62917 ( .A(n50134), .Z(n53842) );
  XOR U62918 ( .A(n53841), .B(n53842), .Z(n52796) );
  IV U62919 ( .A(n50135), .Z(n50136) );
  NOR U62920 ( .A(n50143), .B(n50136), .Z(n52795) );
  IV U62921 ( .A(n50137), .Z(n50138) );
  NOR U62922 ( .A(n50139), .B(n50138), .Z(n53845) );
  NOR U62923 ( .A(n52795), .B(n53845), .Z(n50140) );
  XOR U62924 ( .A(n52796), .B(n50140), .Z(n52788) );
  IV U62925 ( .A(n50141), .Z(n50142) );
  NOR U62926 ( .A(n50143), .B(n50142), .Z(n52789) );
  IV U62927 ( .A(n52789), .Z(n52786) );
  XOR U62928 ( .A(n52788), .B(n52786), .Z(n52782) );
  XOR U62929 ( .A(n50144), .B(n52782), .Z(n52775) );
  XOR U62930 ( .A(n50145), .B(n52775), .Z(n52771) );
  XOR U62931 ( .A(n52769), .B(n52771), .Z(n52774) );
  XOR U62932 ( .A(n50146), .B(n52774), .Z(n50147) );
  IV U62933 ( .A(n50147), .Z(n52761) );
  XOR U62934 ( .A(n52759), .B(n52761), .Z(n52763) );
  XOR U62935 ( .A(n52762), .B(n52763), .Z(n53855) );
  IV U62936 ( .A(n50148), .Z(n50150) );
  NOR U62937 ( .A(n50150), .B(n50149), .Z(n52757) );
  NOR U62938 ( .A(n50151), .B(n53856), .Z(n50152) );
  NOR U62939 ( .A(n52757), .B(n50152), .Z(n50153) );
  XOR U62940 ( .A(n53855), .B(n50153), .Z(n50154) );
  IV U62941 ( .A(n50154), .Z(n53862) );
  XOR U62942 ( .A(n53860), .B(n53862), .Z(n53871) );
  NOR U62943 ( .A(n50161), .B(n53871), .Z(n53869) );
  IV U62944 ( .A(n50155), .Z(n50156) );
  NOR U62945 ( .A(n50157), .B(n50156), .Z(n53870) );
  XOR U62946 ( .A(n53870), .B(n53871), .Z(n52756) );
  IV U62947 ( .A(n50158), .Z(n50160) );
  NOR U62948 ( .A(n50160), .B(n50159), .Z(n50162) );
  IV U62949 ( .A(n50162), .Z(n52755) );
  XOR U62950 ( .A(n52756), .B(n52755), .Z(n50164) );
  NOR U62951 ( .A(n50162), .B(n50161), .Z(n50163) );
  NOR U62952 ( .A(n50164), .B(n50163), .Z(n50165) );
  NOR U62953 ( .A(n53869), .B(n50165), .Z(n50166) );
  IV U62954 ( .A(n50166), .Z(n52753) );
  XOR U62955 ( .A(n52751), .B(n52753), .Z(n52749) );
  IV U62956 ( .A(n52749), .Z(n50174) );
  IV U62957 ( .A(n50167), .Z(n50168) );
  NOR U62958 ( .A(n50169), .B(n50168), .Z(n52752) );
  IV U62959 ( .A(n50170), .Z(n50172) );
  NOR U62960 ( .A(n50172), .B(n50171), .Z(n52748) );
  NOR U62961 ( .A(n52752), .B(n52748), .Z(n50173) );
  XOR U62962 ( .A(n50174), .B(n50173), .Z(n52747) );
  IV U62963 ( .A(n50175), .Z(n50178) );
  IV U62964 ( .A(n50176), .Z(n50177) );
  NOR U62965 ( .A(n50178), .B(n50177), .Z(n52742) );
  NOR U62966 ( .A(n52745), .B(n52742), .Z(n50179) );
  XOR U62967 ( .A(n52747), .B(n50179), .Z(n50180) );
  NOR U62968 ( .A(n50181), .B(n50180), .Z(n50184) );
  IV U62969 ( .A(n50181), .Z(n50183) );
  XOR U62970 ( .A(n52745), .B(n52747), .Z(n50182) );
  NOR U62971 ( .A(n50183), .B(n50182), .Z(n52741) );
  NOR U62972 ( .A(n50184), .B(n52741), .Z(n50185) );
  IV U62973 ( .A(n50185), .Z(n53888) );
  IV U62974 ( .A(n50186), .Z(n50187) );
  NOR U62975 ( .A(n50188), .B(n50187), .Z(n52739) );
  IV U62976 ( .A(n50189), .Z(n50190) );
  NOR U62977 ( .A(n50190), .B(n50197), .Z(n53887) );
  NOR U62978 ( .A(n52739), .B(n53887), .Z(n50191) );
  XOR U62979 ( .A(n53888), .B(n50191), .Z(n50200) );
  IV U62980 ( .A(n50200), .Z(n50195) );
  IV U62981 ( .A(n50192), .Z(n50193) );
  NOR U62982 ( .A(n50193), .B(n50211), .Z(n50208) );
  IV U62983 ( .A(n50208), .Z(n50194) );
  NOR U62984 ( .A(n50195), .B(n50194), .Z(n57530) );
  IV U62985 ( .A(n50196), .Z(n50198) );
  NOR U62986 ( .A(n50198), .B(n50197), .Z(n50201) );
  IV U62987 ( .A(n50201), .Z(n50199) );
  NOR U62988 ( .A(n50199), .B(n53888), .Z(n52738) );
  NOR U62989 ( .A(n50201), .B(n50200), .Z(n50202) );
  NOR U62990 ( .A(n52738), .B(n50202), .Z(n50203) );
  IV U62991 ( .A(n50203), .Z(n52736) );
  IV U62992 ( .A(n50204), .Z(n50205) );
  NOR U62993 ( .A(n50205), .B(n50211), .Z(n50206) );
  IV U62994 ( .A(n50206), .Z(n52735) );
  XOR U62995 ( .A(n52736), .B(n52735), .Z(n50207) );
  NOR U62996 ( .A(n50208), .B(n50207), .Z(n50209) );
  NOR U62997 ( .A(n57530), .B(n50209), .Z(n50210) );
  IV U62998 ( .A(n50210), .Z(n53892) );
  NOR U62999 ( .A(n50212), .B(n50211), .Z(n53891) );
  XOR U63000 ( .A(n53892), .B(n53891), .Z(n53895) );
  IV U63001 ( .A(n50213), .Z(n50214) );
  NOR U63002 ( .A(n50217), .B(n50214), .Z(n52733) );
  IV U63003 ( .A(n50215), .Z(n50216) );
  NOR U63004 ( .A(n50217), .B(n50216), .Z(n53894) );
  NOR U63005 ( .A(n50218), .B(n52724), .Z(n52731) );
  NOR U63006 ( .A(n53894), .B(n52731), .Z(n50219) );
  XOR U63007 ( .A(n52733), .B(n50219), .Z(n50220) );
  XOR U63008 ( .A(n53895), .B(n50220), .Z(n50221) );
  IV U63009 ( .A(n50221), .Z(n52725) );
  XOR U63010 ( .A(n50222), .B(n52725), .Z(n52722) );
  XOR U63011 ( .A(n52720), .B(n52722), .Z(n53903) );
  IV U63012 ( .A(n50223), .Z(n50229) );
  IV U63013 ( .A(n50224), .Z(n50226) );
  NOR U63014 ( .A(n50226), .B(n50225), .Z(n50227) );
  IV U63015 ( .A(n50227), .Z(n50228) );
  NOR U63016 ( .A(n50229), .B(n50228), .Z(n53901) );
  XOR U63017 ( .A(n53903), .B(n53901), .Z(n53899) );
  XOR U63018 ( .A(n53900), .B(n53899), .Z(n52717) );
  NOR U63019 ( .A(n50231), .B(n50230), .Z(n52716) );
  IV U63020 ( .A(n50232), .Z(n50234) );
  IV U63021 ( .A(n50233), .Z(n50238) );
  NOR U63022 ( .A(n50234), .B(n50238), .Z(n52714) );
  NOR U63023 ( .A(n52716), .B(n52714), .Z(n50235) );
  XOR U63024 ( .A(n52717), .B(n50235), .Z(n52713) );
  IV U63025 ( .A(n50236), .Z(n50240) );
  NOR U63026 ( .A(n52713), .B(n50240), .Z(n52711) );
  IV U63027 ( .A(n50237), .Z(n50239) );
  NOR U63028 ( .A(n50239), .B(n50238), .Z(n50241) );
  IV U63029 ( .A(n50241), .Z(n52712) );
  XOR U63030 ( .A(n52713), .B(n52712), .Z(n50243) );
  NOR U63031 ( .A(n50241), .B(n50240), .Z(n50242) );
  NOR U63032 ( .A(n50243), .B(n50242), .Z(n52708) );
  NOR U63033 ( .A(n52711), .B(n52708), .Z(n50244) );
  IV U63034 ( .A(n50244), .Z(n53915) );
  IV U63035 ( .A(n50245), .Z(n50247) );
  NOR U63036 ( .A(n50247), .B(n50246), .Z(n53913) );
  NOR U63037 ( .A(n53913), .B(n50248), .Z(n50249) );
  XOR U63038 ( .A(n53915), .B(n50249), .Z(n52700) );
  XOR U63039 ( .A(n52698), .B(n52700), .Z(n50253) );
  NOR U63040 ( .A(n50251), .B(n50250), .Z(n52695) );
  NOR U63041 ( .A(n52702), .B(n52695), .Z(n50252) );
  XOR U63042 ( .A(n50253), .B(n50252), .Z(n52688) );
  XOR U63043 ( .A(n50254), .B(n52688), .Z(n52684) );
  XOR U63044 ( .A(n52682), .B(n52684), .Z(n52687) );
  XOR U63045 ( .A(n52685), .B(n52687), .Z(n53922) );
  XOR U63046 ( .A(n50255), .B(n53922), .Z(n50256) );
  IV U63047 ( .A(n50256), .Z(n53925) );
  XOR U63048 ( .A(n53923), .B(n53925), .Z(n53927) );
  XOR U63049 ( .A(n53926), .B(n53927), .Z(n52673) );
  IV U63050 ( .A(n52673), .Z(n50263) );
  NOR U63051 ( .A(n50258), .B(n50257), .Z(n52672) );
  IV U63052 ( .A(n50259), .Z(n50261) );
  NOR U63053 ( .A(n50261), .B(n50260), .Z(n52670) );
  NOR U63054 ( .A(n52672), .B(n52670), .Z(n50262) );
  XOR U63055 ( .A(n50263), .B(n50262), .Z(n53933) );
  IV U63056 ( .A(n50264), .Z(n50266) );
  NOR U63057 ( .A(n50266), .B(n50265), .Z(n53931) );
  XOR U63058 ( .A(n53933), .B(n53931), .Z(n53936) );
  XOR U63059 ( .A(n53934), .B(n53936), .Z(n53940) );
  XOR U63060 ( .A(n50267), .B(n53940), .Z(n50268) );
  IV U63061 ( .A(n50268), .Z(n53952) );
  XOR U63062 ( .A(n53950), .B(n53952), .Z(n53953) );
  XOR U63063 ( .A(n53954), .B(n53953), .Z(n52662) );
  IV U63064 ( .A(n50269), .Z(n50270) );
  NOR U63065 ( .A(n50270), .B(n50276), .Z(n52666) );
  IV U63066 ( .A(n50271), .Z(n50273) );
  NOR U63067 ( .A(n50273), .B(n50272), .Z(n52663) );
  NOR U63068 ( .A(n52666), .B(n52663), .Z(n50274) );
  XOR U63069 ( .A(n52662), .B(n50274), .Z(n52661) );
  IV U63070 ( .A(n50275), .Z(n50277) );
  NOR U63071 ( .A(n50277), .B(n50276), .Z(n52659) );
  XOR U63072 ( .A(n52661), .B(n52659), .Z(n52652) );
  XOR U63073 ( .A(n52651), .B(n52652), .Z(n52656) );
  IV U63074 ( .A(n50278), .Z(n50279) );
  NOR U63075 ( .A(n50280), .B(n50279), .Z(n52654) );
  XOR U63076 ( .A(n52656), .B(n52654), .Z(n53958) );
  IV U63077 ( .A(n53958), .Z(n50281) );
  NOR U63078 ( .A(n50282), .B(n50281), .Z(n50292) );
  IV U63079 ( .A(n50283), .Z(n50286) );
  NOR U63080 ( .A(n50284), .B(n52652), .Z(n50285) );
  IV U63081 ( .A(n50285), .Z(n50288) );
  NOR U63082 ( .A(n50286), .B(n50288), .Z(n57581) );
  IV U63083 ( .A(n50287), .Z(n50289) );
  NOR U63084 ( .A(n50289), .B(n50288), .Z(n56199) );
  NOR U63085 ( .A(n57581), .B(n56199), .Z(n50290) );
  IV U63086 ( .A(n50290), .Z(n50291) );
  NOR U63087 ( .A(n50292), .B(n50291), .Z(n50299) );
  IV U63088 ( .A(n50299), .Z(n53966) );
  NOR U63089 ( .A(n50293), .B(n53966), .Z(n57600) );
  NOR U63090 ( .A(n50294), .B(n53959), .Z(n50298) );
  IV U63091 ( .A(n50295), .Z(n50297) );
  NOR U63092 ( .A(n50297), .B(n50296), .Z(n53965) );
  NOR U63093 ( .A(n50298), .B(n53965), .Z(n50300) );
  XOR U63094 ( .A(n50300), .B(n50299), .Z(n50307) );
  IV U63095 ( .A(n50307), .Z(n50301) );
  NOR U63096 ( .A(n50302), .B(n50301), .Z(n50303) );
  NOR U63097 ( .A(n57600), .B(n50303), .Z(n50304) );
  NOR U63098 ( .A(n50305), .B(n50304), .Z(n50308) );
  IV U63099 ( .A(n50305), .Z(n50306) );
  NOR U63100 ( .A(n50307), .B(n50306), .Z(n57603) );
  NOR U63101 ( .A(n50308), .B(n57603), .Z(n52643) );
  IV U63102 ( .A(n50309), .Z(n50311) );
  NOR U63103 ( .A(n50311), .B(n50310), .Z(n50312) );
  IV U63104 ( .A(n50312), .Z(n52644) );
  XOR U63105 ( .A(n52643), .B(n52644), .Z(n52648) );
  IV U63106 ( .A(n50313), .Z(n50317) );
  IV U63107 ( .A(n50314), .Z(n50326) );
  NOR U63108 ( .A(n50326), .B(n50315), .Z(n50316) );
  IV U63109 ( .A(n50316), .Z(n50319) );
  NOR U63110 ( .A(n50317), .B(n50319), .Z(n52646) );
  XOR U63111 ( .A(n52648), .B(n52646), .Z(n53973) );
  IV U63112 ( .A(n53973), .Z(n53971) );
  IV U63113 ( .A(n50318), .Z(n50320) );
  NOR U63114 ( .A(n50320), .B(n50319), .Z(n53970) );
  IV U63115 ( .A(n53970), .Z(n53972) );
  XOR U63116 ( .A(n53971), .B(n53972), .Z(n52640) );
  IV U63117 ( .A(n50321), .Z(n50322) );
  NOR U63118 ( .A(n50323), .B(n50322), .Z(n52638) );
  IV U63119 ( .A(n50324), .Z(n50325) );
  NOR U63120 ( .A(n50326), .B(n50325), .Z(n53974) );
  NOR U63121 ( .A(n52638), .B(n53974), .Z(n50327) );
  XOR U63122 ( .A(n52640), .B(n50327), .Z(n50328) );
  IV U63123 ( .A(n50328), .Z(n52637) );
  IV U63124 ( .A(n50329), .Z(n50330) );
  NOR U63125 ( .A(n50331), .B(n50330), .Z(n50332) );
  IV U63126 ( .A(n50332), .Z(n52636) );
  XOR U63127 ( .A(n52637), .B(n52636), .Z(n52629) );
  XOR U63128 ( .A(n52630), .B(n52629), .Z(n53980) );
  NOR U63129 ( .A(n50336), .B(n50333), .Z(n53979) );
  IV U63130 ( .A(n50334), .Z(n50335) );
  NOR U63131 ( .A(n50336), .B(n50335), .Z(n52631) );
  NOR U63132 ( .A(n53979), .B(n52631), .Z(n50337) );
  XOR U63133 ( .A(n53980), .B(n50337), .Z(n53985) );
  XOR U63134 ( .A(n53983), .B(n53985), .Z(n53987) );
  XOR U63135 ( .A(n53986), .B(n53987), .Z(n52620) );
  XOR U63136 ( .A(n52619), .B(n52620), .Z(n52623) );
  XOR U63137 ( .A(n52622), .B(n52623), .Z(n53992) );
  XOR U63138 ( .A(n53991), .B(n53992), .Z(n52617) );
  IV U63139 ( .A(n50338), .Z(n50341) );
  NOR U63140 ( .A(n50339), .B(n50341), .Z(n53990) );
  IV U63141 ( .A(n50340), .Z(n50344) );
  NOR U63142 ( .A(n50342), .B(n50341), .Z(n50343) );
  IV U63143 ( .A(n50343), .Z(n50350) );
  NOR U63144 ( .A(n50344), .B(n50350), .Z(n52616) );
  NOR U63145 ( .A(n53990), .B(n52616), .Z(n50345) );
  XOR U63146 ( .A(n52617), .B(n50345), .Z(n52613) );
  IV U63147 ( .A(n50346), .Z(n50347) );
  NOR U63148 ( .A(n50348), .B(n50347), .Z(n52614) );
  IV U63149 ( .A(n50349), .Z(n50351) );
  NOR U63150 ( .A(n50351), .B(n50350), .Z(n53994) );
  NOR U63151 ( .A(n52614), .B(n53994), .Z(n50352) );
  XOR U63152 ( .A(n52613), .B(n50352), .Z(n53999) );
  IV U63153 ( .A(n50353), .Z(n52609) );
  NOR U63154 ( .A(n50354), .B(n52609), .Z(n50355) );
  NOR U63155 ( .A(n53997), .B(n50355), .Z(n50356) );
  XOR U63156 ( .A(n53999), .B(n50356), .Z(n50357) );
  IV U63157 ( .A(n50357), .Z(n54006) );
  XOR U63158 ( .A(n54004), .B(n54006), .Z(n54007) );
  XOR U63159 ( .A(n54008), .B(n54007), .Z(n52605) );
  IV U63160 ( .A(n50358), .Z(n50360) );
  NOR U63161 ( .A(n50360), .B(n50359), .Z(n50361) );
  IV U63162 ( .A(n50361), .Z(n52606) );
  XOR U63163 ( .A(n52605), .B(n52606), .Z(n54014) );
  IV U63164 ( .A(n50362), .Z(n50363) );
  NOR U63165 ( .A(n50364), .B(n50363), .Z(n54012) );
  XOR U63166 ( .A(n54014), .B(n54012), .Z(n54011) );
  XOR U63167 ( .A(n52604), .B(n54011), .Z(n50365) );
  XOR U63168 ( .A(n54010), .B(n50365), .Z(n52601) );
  IV U63169 ( .A(n50366), .Z(n50368) );
  NOR U63170 ( .A(n50368), .B(n50367), .Z(n52600) );
  IV U63171 ( .A(n50369), .Z(n50370) );
  NOR U63172 ( .A(n50370), .B(n50375), .Z(n52598) );
  NOR U63173 ( .A(n52600), .B(n52598), .Z(n50371) );
  XOR U63174 ( .A(n52601), .B(n50371), .Z(n50372) );
  IV U63175 ( .A(n50372), .Z(n54025) );
  IV U63176 ( .A(n50373), .Z(n50374) );
  NOR U63177 ( .A(n50375), .B(n50374), .Z(n50376) );
  IV U63178 ( .A(n50376), .Z(n54024) );
  XOR U63179 ( .A(n54025), .B(n54024), .Z(n50382) );
  IV U63180 ( .A(n50382), .Z(n54026) );
  NOR U63181 ( .A(n50381), .B(n54026), .Z(n52597) );
  IV U63182 ( .A(n50377), .Z(n50378) );
  NOR U63183 ( .A(n50379), .B(n50378), .Z(n50380) );
  IV U63184 ( .A(n50380), .Z(n54027) );
  XOR U63185 ( .A(n54027), .B(n54026), .Z(n50384) );
  NOR U63186 ( .A(n50382), .B(n50381), .Z(n50383) );
  NOR U63187 ( .A(n50384), .B(n50383), .Z(n52594) );
  NOR U63188 ( .A(n52597), .B(n52594), .Z(n52583) );
  IV U63189 ( .A(n50385), .Z(n50387) );
  NOR U63190 ( .A(n50387), .B(n50386), .Z(n52593) );
  NOR U63191 ( .A(n50388), .B(n52585), .Z(n50389) );
  NOR U63192 ( .A(n52593), .B(n50389), .Z(n50390) );
  XOR U63193 ( .A(n52583), .B(n50390), .Z(n52581) );
  IV U63194 ( .A(n50391), .Z(n50399) );
  IV U63195 ( .A(n50392), .Z(n50393) );
  NOR U63196 ( .A(n50399), .B(n50393), .Z(n50394) );
  IV U63197 ( .A(n50394), .Z(n52580) );
  XOR U63198 ( .A(n52581), .B(n52580), .Z(n50401) );
  IV U63199 ( .A(n50401), .Z(n50395) );
  NOR U63200 ( .A(n50396), .B(n50395), .Z(n54033) );
  IV U63201 ( .A(n50397), .Z(n50398) );
  NOR U63202 ( .A(n50399), .B(n50398), .Z(n50402) );
  IV U63203 ( .A(n50402), .Z(n50400) );
  NOR U63204 ( .A(n52581), .B(n50400), .Z(n56147) );
  NOR U63205 ( .A(n50402), .B(n50401), .Z(n50403) );
  NOR U63206 ( .A(n56147), .B(n50403), .Z(n50413) );
  NOR U63207 ( .A(n50404), .B(n50413), .Z(n50405) );
  NOR U63208 ( .A(n54033), .B(n50405), .Z(n50406) );
  IV U63209 ( .A(n50406), .Z(n54031) );
  IV U63210 ( .A(n50407), .Z(n50408) );
  NOR U63211 ( .A(n50409), .B(n50408), .Z(n50410) );
  IV U63212 ( .A(n50410), .Z(n54030) );
  XOR U63213 ( .A(n54031), .B(n54030), .Z(n50411) );
  NOR U63214 ( .A(n50412), .B(n50411), .Z(n50416) );
  IV U63215 ( .A(n50412), .Z(n50415) );
  IV U63216 ( .A(n50413), .Z(n50414) );
  NOR U63217 ( .A(n50415), .B(n50414), .Z(n57705) );
  NOR U63218 ( .A(n50416), .B(n57705), .Z(n50417) );
  IV U63219 ( .A(n50417), .Z(n54039) );
  IV U63220 ( .A(n50418), .Z(n50420) );
  NOR U63221 ( .A(n50420), .B(n50419), .Z(n54037) );
  XOR U63222 ( .A(n54039), .B(n54037), .Z(n52578) );
  XOR U63223 ( .A(n52577), .B(n52578), .Z(n52575) );
  XOR U63224 ( .A(n52574), .B(n52575), .Z(n52566) );
  XOR U63225 ( .A(n52565), .B(n52566), .Z(n52569) );
  XOR U63226 ( .A(n52568), .B(n52569), .Z(n50435) );
  IV U63227 ( .A(n50435), .Z(n50421) );
  NOR U63228 ( .A(n50422), .B(n50421), .Z(n50432) );
  IV U63229 ( .A(n50423), .Z(n50426) );
  NOR U63230 ( .A(n50424), .B(n52569), .Z(n50425) );
  IV U63231 ( .A(n50425), .Z(n50428) );
  NOR U63232 ( .A(n50426), .B(n50428), .Z(n56133) );
  IV U63233 ( .A(n50427), .Z(n50429) );
  NOR U63234 ( .A(n50429), .B(n50428), .Z(n57719) );
  NOR U63235 ( .A(n56133), .B(n57719), .Z(n50430) );
  IV U63236 ( .A(n50430), .Z(n50431) );
  NOR U63237 ( .A(n50432), .B(n50431), .Z(n50433) );
  NOR U63238 ( .A(n50434), .B(n50433), .Z(n52563) );
  IV U63239 ( .A(n50434), .Z(n50436) );
  NOR U63240 ( .A(n50436), .B(n50435), .Z(n56137) );
  NOR U63241 ( .A(n52563), .B(n56137), .Z(n52556) );
  IV U63242 ( .A(n50437), .Z(n50438) );
  NOR U63243 ( .A(n50438), .B(n57725), .Z(n52561) );
  IV U63244 ( .A(n50439), .Z(n50440) );
  NOR U63245 ( .A(n50440), .B(n57725), .Z(n52557) );
  NOR U63246 ( .A(n52561), .B(n52557), .Z(n50441) );
  XOR U63247 ( .A(n52556), .B(n50441), .Z(n52555) );
  XOR U63248 ( .A(n52553), .B(n52555), .Z(n52549) );
  IV U63249 ( .A(n50442), .Z(n50443) );
  NOR U63250 ( .A(n50444), .B(n50443), .Z(n52551) );
  IV U63251 ( .A(n50445), .Z(n50447) );
  NOR U63252 ( .A(n50447), .B(n50446), .Z(n52548) );
  NOR U63253 ( .A(n52551), .B(n52548), .Z(n50448) );
  XOR U63254 ( .A(n52549), .B(n50448), .Z(n50449) );
  IV U63255 ( .A(n50449), .Z(n52547) );
  IV U63256 ( .A(n50450), .Z(n50452) );
  NOR U63257 ( .A(n50452), .B(n50451), .Z(n50453) );
  IV U63258 ( .A(n50453), .Z(n52546) );
  XOR U63259 ( .A(n52547), .B(n52546), .Z(n52538) );
  XOR U63260 ( .A(n52539), .B(n52538), .Z(n52535) );
  XOR U63261 ( .A(n50454), .B(n52535), .Z(n52528) );
  XOR U63262 ( .A(n50455), .B(n52528), .Z(n52526) );
  XOR U63263 ( .A(n52523), .B(n52526), .Z(n50456) );
  XOR U63264 ( .A(n50457), .B(n50456), .Z(n50458) );
  IV U63265 ( .A(n50458), .Z(n52522) );
  XOR U63266 ( .A(n52520), .B(n52522), .Z(n54060) );
  NOR U63267 ( .A(n50459), .B(n54060), .Z(n54066) );
  IV U63268 ( .A(n50460), .Z(n50461) );
  NOR U63269 ( .A(n50462), .B(n50461), .Z(n52517) );
  IV U63270 ( .A(n50463), .Z(n50465) );
  NOR U63271 ( .A(n50465), .B(n50464), .Z(n54059) );
  XOR U63272 ( .A(n54059), .B(n54060), .Z(n52518) );
  XOR U63273 ( .A(n52517), .B(n52518), .Z(n50471) );
  IV U63274 ( .A(n50471), .Z(n50466) );
  NOR U63275 ( .A(n50467), .B(n50466), .Z(n50468) );
  NOR U63276 ( .A(n54066), .B(n50468), .Z(n50469) );
  NOR U63277 ( .A(n50470), .B(n50469), .Z(n50473) );
  IV U63278 ( .A(n50470), .Z(n50472) );
  NOR U63279 ( .A(n50472), .B(n50471), .Z(n52516) );
  NOR U63280 ( .A(n50473), .B(n52516), .Z(n52512) );
  IV U63281 ( .A(n50474), .Z(n50476) );
  NOR U63282 ( .A(n50476), .B(n50475), .Z(n50477) );
  IV U63283 ( .A(n50477), .Z(n52513) );
  XOR U63284 ( .A(n52512), .B(n52513), .Z(n54071) );
  XOR U63285 ( .A(n54072), .B(n54071), .Z(n52510) );
  XOR U63286 ( .A(n52511), .B(n52510), .Z(n52508) );
  XOR U63287 ( .A(n50478), .B(n52508), .Z(n54097) );
  XOR U63288 ( .A(n50479), .B(n54097), .Z(n54114) );
  XOR U63289 ( .A(n50480), .B(n54114), .Z(n50481) );
  IV U63290 ( .A(n50481), .Z(n54112) );
  XOR U63291 ( .A(n54110), .B(n54112), .Z(n52502) );
  XOR U63292 ( .A(n52501), .B(n52502), .Z(n52505) );
  XOR U63293 ( .A(n52504), .B(n52505), .Z(n54120) );
  XOR U63294 ( .A(n54119), .B(n54120), .Z(n52499) );
  IV U63295 ( .A(n50482), .Z(n50492) );
  NOR U63296 ( .A(n50492), .B(n50484), .Z(n54118) );
  IV U63297 ( .A(n50483), .Z(n50487) );
  NOR U63298 ( .A(n50485), .B(n50484), .Z(n50486) );
  IV U63299 ( .A(n50486), .Z(n50497) );
  NOR U63300 ( .A(n50487), .B(n50497), .Z(n52498) );
  NOR U63301 ( .A(n54118), .B(n52498), .Z(n50488) );
  XOR U63302 ( .A(n52499), .B(n50488), .Z(n50489) );
  IV U63303 ( .A(n50489), .Z(n54125) );
  IV U63304 ( .A(n50490), .Z(n50494) );
  XOR U63305 ( .A(n50492), .B(n50491), .Z(n50493) );
  NOR U63306 ( .A(n50494), .B(n50493), .Z(n50495) );
  IV U63307 ( .A(n50495), .Z(n50499) );
  NOR U63308 ( .A(n54125), .B(n50499), .Z(n54138) );
  IV U63309 ( .A(n50496), .Z(n50498) );
  NOR U63310 ( .A(n50498), .B(n50497), .Z(n50500) );
  IV U63311 ( .A(n50500), .Z(n54124) );
  XOR U63312 ( .A(n54125), .B(n54124), .Z(n50502) );
  NOR U63313 ( .A(n50500), .B(n50499), .Z(n50501) );
  NOR U63314 ( .A(n50502), .B(n50501), .Z(n50504) );
  NOR U63315 ( .A(n54138), .B(n50504), .Z(n52490) );
  NOR U63316 ( .A(n50503), .B(n52490), .Z(n50506) );
  IV U63317 ( .A(n50503), .Z(n50505) );
  NOR U63318 ( .A(n50505), .B(n50504), .Z(n54137) );
  NOR U63319 ( .A(n50506), .B(n54137), .Z(n50507) );
  IV U63320 ( .A(n50507), .Z(n52473) );
  NOR U63321 ( .A(n50509), .B(n50508), .Z(n50517) );
  NOR U63322 ( .A(n50510), .B(n52492), .Z(n50512) );
  NOR U63323 ( .A(n50512), .B(n50511), .Z(n50513) );
  IV U63324 ( .A(n50513), .Z(n50515) );
  NOR U63325 ( .A(n50515), .B(n50514), .Z(n50516) );
  NOR U63326 ( .A(n50517), .B(n50516), .Z(n50518) );
  XOR U63327 ( .A(n52473), .B(n50518), .Z(n52471) );
  IV U63328 ( .A(n50519), .Z(n50521) );
  NOR U63329 ( .A(n50521), .B(n50520), .Z(n50522) );
  IV U63330 ( .A(n50522), .Z(n52470) );
  XOR U63331 ( .A(n52471), .B(n52470), .Z(n50523) );
  NOR U63332 ( .A(n50527), .B(n50523), .Z(n50531) );
  IV U63333 ( .A(n50524), .Z(n50525) );
  NOR U63334 ( .A(n50526), .B(n50525), .Z(n50533) );
  IV U63335 ( .A(n50527), .Z(n50528) );
  NOR U63336 ( .A(n52471), .B(n50528), .Z(n50529) );
  NOR U63337 ( .A(n50533), .B(n50529), .Z(n50530) );
  NOR U63338 ( .A(n50531), .B(n50530), .Z(n56040) );
  IV U63339 ( .A(n50531), .Z(n50532) );
  NOR U63340 ( .A(n50533), .B(n50532), .Z(n50534) );
  NOR U63341 ( .A(n56040), .B(n50534), .Z(n52463) );
  IV U63342 ( .A(n52463), .Z(n52461) );
  XOR U63343 ( .A(n52464), .B(n52461), .Z(n54141) );
  IV U63344 ( .A(n50535), .Z(n50536) );
  NOR U63345 ( .A(n50536), .B(n50542), .Z(n50537) );
  IV U63346 ( .A(n50537), .Z(n52460) );
  XOR U63347 ( .A(n54141), .B(n52460), .Z(n50545) );
  IV U63348 ( .A(n50538), .Z(n50539) );
  NOR U63349 ( .A(n50540), .B(n50539), .Z(n52465) );
  IV U63350 ( .A(n50541), .Z(n50543) );
  NOR U63351 ( .A(n50543), .B(n50542), .Z(n54140) );
  NOR U63352 ( .A(n52465), .B(n54140), .Z(n50544) );
  XOR U63353 ( .A(n50545), .B(n50544), .Z(n54146) );
  IV U63354 ( .A(n50546), .Z(n50548) );
  NOR U63355 ( .A(n50548), .B(n50547), .Z(n54144) );
  XOR U63356 ( .A(n54146), .B(n54144), .Z(n54149) );
  XOR U63357 ( .A(n54147), .B(n54149), .Z(n52458) );
  NOR U63358 ( .A(n50549), .B(n52458), .Z(n56075) );
  IV U63359 ( .A(n50550), .Z(n50551) );
  NOR U63360 ( .A(n50552), .B(n50551), .Z(n52457) );
  XOR U63361 ( .A(n52457), .B(n52458), .Z(n50561) );
  IV U63362 ( .A(n50561), .Z(n50553) );
  NOR U63363 ( .A(n50554), .B(n50553), .Z(n50555) );
  NOR U63364 ( .A(n56075), .B(n50555), .Z(n50563) );
  IV U63365 ( .A(n50563), .Z(n50556) );
  NOR U63366 ( .A(n50557), .B(n50556), .Z(n52456) );
  IV U63367 ( .A(n50558), .Z(n50560) );
  NOR U63368 ( .A(n50560), .B(n50559), .Z(n50564) );
  IV U63369 ( .A(n50564), .Z(n50562) );
  NOR U63370 ( .A(n50562), .B(n50561), .Z(n56028) );
  NOR U63371 ( .A(n50564), .B(n50563), .Z(n50565) );
  NOR U63372 ( .A(n56028), .B(n50565), .Z(n50566) );
  NOR U63373 ( .A(n50567), .B(n50566), .Z(n50568) );
  NOR U63374 ( .A(n52456), .B(n50568), .Z(n50569) );
  IV U63375 ( .A(n50569), .Z(n52453) );
  XOR U63376 ( .A(n52452), .B(n52453), .Z(n52450) );
  IV U63377 ( .A(n50570), .Z(n50571) );
  NOR U63378 ( .A(n50572), .B(n50571), .Z(n52449) );
  IV U63379 ( .A(n50573), .Z(n50574) );
  NOR U63380 ( .A(n50579), .B(n50574), .Z(n52447) );
  NOR U63381 ( .A(n52449), .B(n52447), .Z(n50575) );
  XOR U63382 ( .A(n52450), .B(n50575), .Z(n50582) );
  IV U63383 ( .A(n50582), .Z(n50576) );
  NOR U63384 ( .A(n50577), .B(n50576), .Z(n56007) );
  IV U63385 ( .A(n50578), .Z(n50580) );
  NOR U63386 ( .A(n50580), .B(n50579), .Z(n50583) );
  IV U63387 ( .A(n50583), .Z(n50581) );
  NOR U63388 ( .A(n50581), .B(n52450), .Z(n56023) );
  NOR U63389 ( .A(n50583), .B(n50582), .Z(n50584) );
  NOR U63390 ( .A(n56023), .B(n50584), .Z(n52444) );
  NOR U63391 ( .A(n50585), .B(n52444), .Z(n50586) );
  NOR U63392 ( .A(n56007), .B(n50586), .Z(n54154) );
  IV U63393 ( .A(n50587), .Z(n50589) );
  NOR U63394 ( .A(n50589), .B(n50588), .Z(n52443) );
  IV U63395 ( .A(n50590), .Z(n50591) );
  NOR U63396 ( .A(n50591), .B(n50594), .Z(n54155) );
  NOR U63397 ( .A(n52443), .B(n54155), .Z(n50592) );
  XOR U63398 ( .A(n54154), .B(n50592), .Z(n52437) );
  IV U63399 ( .A(n50593), .Z(n50595) );
  NOR U63400 ( .A(n50595), .B(n50594), .Z(n52435) );
  XOR U63401 ( .A(n52437), .B(n52435), .Z(n52439) );
  XOR U63402 ( .A(n52438), .B(n52439), .Z(n52428) );
  XOR U63403 ( .A(n52427), .B(n52428), .Z(n52432) );
  XOR U63404 ( .A(n52430), .B(n52432), .Z(n54160) );
  XOR U63405 ( .A(n54158), .B(n54160), .Z(n54161) );
  XOR U63406 ( .A(n54162), .B(n54161), .Z(n54167) );
  IV U63407 ( .A(n54167), .Z(n54165) );
  XOR U63408 ( .A(n54166), .B(n54165), .Z(n52423) );
  XOR U63409 ( .A(n50596), .B(n52423), .Z(n50602) );
  NOR U63410 ( .A(n50597), .B(n50602), .Z(n55975) );
  IV U63411 ( .A(n50598), .Z(n50599) );
  NOR U63412 ( .A(n50600), .B(n50599), .Z(n50604) );
  IV U63413 ( .A(n50604), .Z(n50601) );
  NOR U63414 ( .A(n50601), .B(n52423), .Z(n57868) );
  IV U63415 ( .A(n50602), .Z(n50603) );
  NOR U63416 ( .A(n50604), .B(n50603), .Z(n50605) );
  NOR U63417 ( .A(n57868), .B(n50605), .Z(n50610) );
  NOR U63418 ( .A(n50606), .B(n50610), .Z(n50607) );
  NOR U63419 ( .A(n55975), .B(n50607), .Z(n50608) );
  NOR U63420 ( .A(n50609), .B(n50608), .Z(n50613) );
  IV U63421 ( .A(n50609), .Z(n50612) );
  IV U63422 ( .A(n50610), .Z(n50611) );
  NOR U63423 ( .A(n50612), .B(n50611), .Z(n55976) );
  NOR U63424 ( .A(n50613), .B(n55976), .Z(n50619) );
  IV U63425 ( .A(n50619), .Z(n54177) );
  NOR U63426 ( .A(n50614), .B(n54177), .Z(n55983) );
  IV U63427 ( .A(n50615), .Z(n50617) );
  NOR U63428 ( .A(n50617), .B(n50616), .Z(n50618) );
  IV U63429 ( .A(n50618), .Z(n54176) );
  XOR U63430 ( .A(n50619), .B(n54176), .Z(n50625) );
  IV U63431 ( .A(n50625), .Z(n50620) );
  NOR U63432 ( .A(n50621), .B(n50620), .Z(n50622) );
  NOR U63433 ( .A(n55983), .B(n50622), .Z(n50623) );
  NOR U63434 ( .A(n50624), .B(n50623), .Z(n52421) );
  IV U63435 ( .A(n50624), .Z(n50626) );
  NOR U63436 ( .A(n50626), .B(n50625), .Z(n52418) );
  NOR U63437 ( .A(n52421), .B(n52418), .Z(n52414) );
  IV U63438 ( .A(n50627), .Z(n50629) );
  NOR U63439 ( .A(n50629), .B(n50628), .Z(n52419) );
  IV U63440 ( .A(n50630), .Z(n50631) );
  NOR U63441 ( .A(n50631), .B(n50634), .Z(n52415) );
  NOR U63442 ( .A(n52419), .B(n52415), .Z(n50632) );
  XOR U63443 ( .A(n52414), .B(n50632), .Z(n52413) );
  IV U63444 ( .A(n50633), .Z(n50635) );
  NOR U63445 ( .A(n50635), .B(n50634), .Z(n50636) );
  IV U63446 ( .A(n50636), .Z(n52412) );
  XOR U63447 ( .A(n52413), .B(n52412), .Z(n50643) );
  IV U63448 ( .A(n50643), .Z(n50637) );
  NOR U63449 ( .A(n50638), .B(n50637), .Z(n52411) );
  IV U63450 ( .A(n50639), .Z(n50640) );
  NOR U63451 ( .A(n50641), .B(n50640), .Z(n50644) );
  IV U63452 ( .A(n50644), .Z(n50642) );
  NOR U63453 ( .A(n52413), .B(n50642), .Z(n55967) );
  NOR U63454 ( .A(n50644), .B(n50643), .Z(n50645) );
  NOR U63455 ( .A(n55967), .B(n50645), .Z(n50652) );
  NOR U63456 ( .A(n50646), .B(n50652), .Z(n50647) );
  NOR U63457 ( .A(n52411), .B(n50647), .Z(n50655) );
  IV U63458 ( .A(n50655), .Z(n50648) );
  NOR U63459 ( .A(n50649), .B(n50648), .Z(n57879) );
  IV U63460 ( .A(n50650), .Z(n50651) );
  NOR U63461 ( .A(n50651), .B(n50660), .Z(n50656) );
  IV U63462 ( .A(n50656), .Z(n50654) );
  IV U63463 ( .A(n50652), .Z(n50653) );
  NOR U63464 ( .A(n50654), .B(n50653), .Z(n54185) );
  NOR U63465 ( .A(n50656), .B(n50655), .Z(n50657) );
  NOR U63466 ( .A(n54185), .B(n50657), .Z(n50658) );
  IV U63467 ( .A(n50658), .Z(n54183) );
  IV U63468 ( .A(n50659), .Z(n50661) );
  NOR U63469 ( .A(n50661), .B(n50660), .Z(n50662) );
  IV U63470 ( .A(n50662), .Z(n54182) );
  XOR U63471 ( .A(n54183), .B(n54182), .Z(n50663) );
  NOR U63472 ( .A(n50664), .B(n50663), .Z(n50665) );
  NOR U63473 ( .A(n57879), .B(n50665), .Z(n50666) );
  IV U63474 ( .A(n50666), .Z(n52409) );
  IV U63475 ( .A(n50667), .Z(n50668) );
  NOR U63476 ( .A(n50669), .B(n50668), .Z(n52408) );
  XOR U63477 ( .A(n52409), .B(n52408), .Z(n54194) );
  XOR U63478 ( .A(n50670), .B(n54194), .Z(n50671) );
  IV U63479 ( .A(n50671), .Z(n54197) );
  XOR U63480 ( .A(n54196), .B(n54197), .Z(n52395) );
  XOR U63481 ( .A(n52397), .B(n52395), .Z(n54209) );
  XOR U63482 ( .A(n54202), .B(n54209), .Z(n52392) );
  IV U63483 ( .A(n50672), .Z(n50674) );
  NOR U63484 ( .A(n50674), .B(n50673), .Z(n54208) );
  IV U63485 ( .A(n50675), .Z(n50676) );
  NOR U63486 ( .A(n50676), .B(n50679), .Z(n52391) );
  NOR U63487 ( .A(n54208), .B(n52391), .Z(n50677) );
  XOR U63488 ( .A(n52392), .B(n50677), .Z(n52378) );
  IV U63489 ( .A(n50678), .Z(n50680) );
  NOR U63490 ( .A(n50680), .B(n50679), .Z(n52379) );
  IV U63491 ( .A(n52379), .Z(n52380) );
  XOR U63492 ( .A(n52378), .B(n52380), .Z(n52370) );
  XOR U63493 ( .A(n50681), .B(n52370), .Z(n54214) );
  XOR U63494 ( .A(n50682), .B(n54214), .Z(n54236) );
  XOR U63495 ( .A(n54228), .B(n54236), .Z(n52367) );
  NOR U63496 ( .A(n50683), .B(n52367), .Z(n55946) );
  IV U63497 ( .A(n50684), .Z(n50686) );
  NOR U63498 ( .A(n50686), .B(n50685), .Z(n52366) );
  XOR U63499 ( .A(n52366), .B(n52367), .Z(n54254) );
  IV U63500 ( .A(n54254), .Z(n50687) );
  NOR U63501 ( .A(n50688), .B(n50687), .Z(n50689) );
  NOR U63502 ( .A(n55946), .B(n50689), .Z(n50694) );
  IV U63503 ( .A(n50690), .Z(n50692) );
  NOR U63504 ( .A(n50692), .B(n50691), .Z(n54253) );
  NOR U63505 ( .A(n54235), .B(n54253), .Z(n50693) );
  XOR U63506 ( .A(n50694), .B(n50693), .Z(n54258) );
  XOR U63507 ( .A(n54257), .B(n54258), .Z(n54263) );
  IV U63508 ( .A(n50695), .Z(n50697) );
  NOR U63509 ( .A(n50697), .B(n50696), .Z(n54256) );
  IV U63510 ( .A(n50698), .Z(n50699) );
  NOR U63511 ( .A(n50700), .B(n50699), .Z(n54261) );
  NOR U63512 ( .A(n54256), .B(n54261), .Z(n50701) );
  XOR U63513 ( .A(n54263), .B(n50701), .Z(n52362) );
  NOR U63514 ( .A(n50703), .B(n50702), .Z(n52364) );
  IV U63515 ( .A(n50704), .Z(n50705) );
  IV U63516 ( .A(n50714), .Z(n50707) );
  NOR U63517 ( .A(n50705), .B(n50707), .Z(n52361) );
  IV U63518 ( .A(n50706), .Z(n50708) );
  NOR U63519 ( .A(n50708), .B(n50707), .Z(n54277) );
  NOR U63520 ( .A(n52361), .B(n54277), .Z(n50709) );
  IV U63521 ( .A(n50709), .Z(n50710) );
  NOR U63522 ( .A(n52364), .B(n50710), .Z(n50711) );
  XOR U63523 ( .A(n52362), .B(n50711), .Z(n54276) );
  IV U63524 ( .A(n50712), .Z(n50716) );
  XOR U63525 ( .A(n50714), .B(n50713), .Z(n50715) );
  NOR U63526 ( .A(n50716), .B(n50715), .Z(n54274) );
  XOR U63527 ( .A(n54276), .B(n54274), .Z(n52359) );
  XOR U63528 ( .A(n50717), .B(n52359), .Z(n50718) );
  IV U63529 ( .A(n50718), .Z(n54285) );
  XOR U63530 ( .A(n52354), .B(n54285), .Z(n54290) );
  IV U63531 ( .A(n50719), .Z(n50729) );
  IV U63532 ( .A(n50720), .Z(n50721) );
  NOR U63533 ( .A(n50729), .B(n50721), .Z(n54291) );
  NOR U63534 ( .A(n54283), .B(n54291), .Z(n50722) );
  XOR U63535 ( .A(n54290), .B(n50722), .Z(n52353) );
  IV U63536 ( .A(n50723), .Z(n50724) );
  NOR U63537 ( .A(n50725), .B(n50724), .Z(n50731) );
  IV U63538 ( .A(n50731), .Z(n50726) );
  NOR U63539 ( .A(n52353), .B(n50726), .Z(n57933) );
  IV U63540 ( .A(n50727), .Z(n50728) );
  NOR U63541 ( .A(n50729), .B(n50728), .Z(n52351) );
  XOR U63542 ( .A(n52351), .B(n52353), .Z(n50739) );
  IV U63543 ( .A(n50739), .Z(n50730) );
  NOR U63544 ( .A(n50731), .B(n50730), .Z(n50732) );
  NOR U63545 ( .A(n57933), .B(n50732), .Z(n50737) );
  IV U63546 ( .A(n50737), .Z(n50733) );
  NOR U63547 ( .A(n50734), .B(n50733), .Z(n57946) );
  NOR U63548 ( .A(n50736), .B(n50735), .Z(n50738) );
  NOR U63549 ( .A(n50738), .B(n50737), .Z(n50741) );
  IV U63550 ( .A(n50738), .Z(n50740) );
  NOR U63551 ( .A(n50740), .B(n50739), .Z(n57930) );
  NOR U63552 ( .A(n50741), .B(n57930), .Z(n52348) );
  NOR U63553 ( .A(n50742), .B(n52348), .Z(n50743) );
  NOR U63554 ( .A(n57946), .B(n50743), .Z(n50744) );
  IV U63555 ( .A(n50744), .Z(n52347) );
  XOR U63556 ( .A(n52350), .B(n52347), .Z(n50745) );
  XOR U63557 ( .A(n52346), .B(n50745), .Z(n54301) );
  IV U63558 ( .A(n54301), .Z(n50753) );
  IV U63559 ( .A(n50746), .Z(n50747) );
  NOR U63560 ( .A(n50748), .B(n50747), .Z(n52344) );
  IV U63561 ( .A(n50749), .Z(n50750) );
  NOR U63562 ( .A(n50751), .B(n50750), .Z(n54299) );
  NOR U63563 ( .A(n52344), .B(n54299), .Z(n50752) );
  XOR U63564 ( .A(n50753), .B(n50752), .Z(n54298) );
  XOR U63565 ( .A(n54296), .B(n54298), .Z(n52342) );
  XOR U63566 ( .A(n50754), .B(n52342), .Z(n50764) );
  IV U63567 ( .A(n50764), .Z(n52335) );
  IV U63568 ( .A(n50755), .Z(n50757) );
  NOR U63569 ( .A(n50757), .B(n50756), .Z(n50767) );
  IV U63570 ( .A(n50767), .Z(n50758) );
  NOR U63571 ( .A(n52335), .B(n50758), .Z(n55882) );
  IV U63572 ( .A(n50759), .Z(n50761) );
  NOR U63573 ( .A(n50761), .B(n50760), .Z(n50765) );
  IV U63574 ( .A(n50765), .Z(n50763) );
  XOR U63575 ( .A(n52341), .B(n52342), .Z(n50762) );
  NOR U63576 ( .A(n50763), .B(n50762), .Z(n52339) );
  NOR U63577 ( .A(n50765), .B(n50764), .Z(n50766) );
  NOR U63578 ( .A(n52339), .B(n50766), .Z(n50771) );
  NOR U63579 ( .A(n50767), .B(n50771), .Z(n50768) );
  NOR U63580 ( .A(n55882), .B(n50768), .Z(n50769) );
  NOR U63581 ( .A(n50770), .B(n50769), .Z(n50774) );
  IV U63582 ( .A(n50770), .Z(n50773) );
  IV U63583 ( .A(n50771), .Z(n50772) );
  NOR U63584 ( .A(n50773), .B(n50772), .Z(n55885) );
  NOR U63585 ( .A(n50774), .B(n55885), .Z(n50779) );
  IV U63586 ( .A(n50775), .Z(n50777) );
  NOR U63587 ( .A(n50777), .B(n50776), .Z(n50778) );
  IV U63588 ( .A(n50778), .Z(n52336) );
  XOR U63589 ( .A(n50779), .B(n52336), .Z(n54307) );
  XOR U63590 ( .A(n50780), .B(n54307), .Z(n50781) );
  IV U63591 ( .A(n50781), .Z(n54315) );
  XOR U63592 ( .A(n50782), .B(n54315), .Z(n58025) );
  XOR U63593 ( .A(n54332), .B(n58025), .Z(n54339) );
  XOR U63594 ( .A(n54336), .B(n54339), .Z(n52325) );
  XOR U63595 ( .A(n54337), .B(n52325), .Z(n52322) );
  XOR U63596 ( .A(n50783), .B(n52322), .Z(n50784) );
  IV U63597 ( .A(n50784), .Z(n52315) );
  XOR U63598 ( .A(n52313), .B(n52315), .Z(n52318) );
  IV U63599 ( .A(n50785), .Z(n50787) );
  NOR U63600 ( .A(n50787), .B(n50786), .Z(n52316) );
  XOR U63601 ( .A(n52318), .B(n52316), .Z(n52307) );
  IV U63602 ( .A(n50788), .Z(n50790) );
  NOR U63603 ( .A(n50790), .B(n50789), .Z(n52305) );
  XOR U63604 ( .A(n52307), .B(n52305), .Z(n52309) );
  XOR U63605 ( .A(n52308), .B(n52309), .Z(n52299) );
  XOR U63606 ( .A(n52298), .B(n52299), .Z(n52301) );
  XOR U63607 ( .A(n52302), .B(n52301), .Z(n52295) );
  XOR U63608 ( .A(n52297), .B(n52295), .Z(n54350) );
  XOR U63609 ( .A(n54349), .B(n54350), .Z(n54353) );
  XOR U63610 ( .A(n54352), .B(n54353), .Z(n50797) );
  IV U63611 ( .A(n50797), .Z(n50795) );
  IV U63612 ( .A(n50791), .Z(n50793) );
  NOR U63613 ( .A(n50793), .B(n50792), .Z(n50796) );
  IV U63614 ( .A(n50796), .Z(n50794) );
  NOR U63615 ( .A(n50795), .B(n50794), .Z(n57992) );
  NOR U63616 ( .A(n50797), .B(n50796), .Z(n54358) );
  NOR U63617 ( .A(n57992), .B(n54358), .Z(n54363) );
  IV U63618 ( .A(n50798), .Z(n50799) );
  NOR U63619 ( .A(n50800), .B(n50799), .Z(n54356) );
  IV U63620 ( .A(n50801), .Z(n50802) );
  NOR U63621 ( .A(n50803), .B(n50802), .Z(n54364) );
  NOR U63622 ( .A(n54356), .B(n54364), .Z(n55871) );
  XOR U63623 ( .A(n54363), .B(n55871), .Z(n54361) );
  XOR U63624 ( .A(n54360), .B(n54361), .Z(n52288) );
  XOR U63625 ( .A(n52287), .B(n52288), .Z(n52291) );
  XOR U63626 ( .A(n52290), .B(n52291), .Z(n52285) );
  XOR U63627 ( .A(n52284), .B(n52285), .Z(n54374) );
  XOR U63628 ( .A(n54373), .B(n54374), .Z(n54371) );
  XOR U63629 ( .A(n54370), .B(n54371), .Z(n52282) );
  XOR U63630 ( .A(n52283), .B(n52282), .Z(n50804) );
  IV U63631 ( .A(n50804), .Z(n54383) );
  IV U63632 ( .A(n50805), .Z(n50807) );
  NOR U63633 ( .A(n50807), .B(n50806), .Z(n54381) );
  XOR U63634 ( .A(n54383), .B(n54381), .Z(n54385) );
  NOR U63635 ( .A(n54384), .B(n52280), .Z(n50808) );
  XOR U63636 ( .A(n54385), .B(n50808), .Z(n52267) );
  NOR U63637 ( .A(n50810), .B(n50809), .Z(n52277) );
  IV U63638 ( .A(n50811), .Z(n52271) );
  IV U63639 ( .A(n52270), .Z(n50814) );
  NOR U63640 ( .A(n52271), .B(n50814), .Z(n52268) );
  NOR U63641 ( .A(n52277), .B(n52268), .Z(n50812) );
  XOR U63642 ( .A(n52267), .B(n50812), .Z(n52272) );
  IV U63643 ( .A(n50813), .Z(n52276) );
  NOR U63644 ( .A(n52276), .B(n50814), .Z(n50817) );
  IV U63645 ( .A(n50815), .Z(n50816) );
  NOR U63646 ( .A(n50821), .B(n50816), .Z(n52265) );
  NOR U63647 ( .A(n50817), .B(n52265), .Z(n50818) );
  XOR U63648 ( .A(n52272), .B(n50818), .Z(n52257) );
  IV U63649 ( .A(n50819), .Z(n50820) );
  NOR U63650 ( .A(n50821), .B(n50820), .Z(n50822) );
  IV U63651 ( .A(n50822), .Z(n52258) );
  XOR U63652 ( .A(n52257), .B(n52258), .Z(n52261) );
  XOR U63653 ( .A(n52260), .B(n52261), .Z(n52256) );
  XOR U63654 ( .A(n50823), .B(n52256), .Z(n52246) );
  XOR U63655 ( .A(n50824), .B(n52246), .Z(n52245) );
  XOR U63656 ( .A(n52244), .B(n52245), .Z(n50834) );
  IV U63657 ( .A(n50834), .Z(n50832) );
  IV U63658 ( .A(n50825), .Z(n50826) );
  NOR U63659 ( .A(n50827), .B(n50826), .Z(n50828) );
  IV U63660 ( .A(n50828), .Z(n50830) );
  NOR U63661 ( .A(n50830), .B(n50829), .Z(n50833) );
  IV U63662 ( .A(n50833), .Z(n50831) );
  NOR U63663 ( .A(n50832), .B(n50831), .Z(n55808) );
  NOR U63664 ( .A(n50834), .B(n50833), .Z(n52243) );
  NOR U63665 ( .A(n55808), .B(n52243), .Z(n55807) );
  XOR U63666 ( .A(n50835), .B(n55807), .Z(n52234) );
  XOR U63667 ( .A(n50836), .B(n52234), .Z(n52229) );
  XOR U63668 ( .A(n52231), .B(n52229), .Z(n55830) );
  XOR U63669 ( .A(n52228), .B(n55830), .Z(n50837) );
  IV U63670 ( .A(n50837), .Z(n52221) );
  XOR U63671 ( .A(n52220), .B(n52221), .Z(n52224) );
  XOR U63672 ( .A(n52223), .B(n52224), .Z(n52213) );
  XOR U63673 ( .A(n52214), .B(n52213), .Z(n50838) );
  XOR U63674 ( .A(n50839), .B(n50838), .Z(n52208) );
  NOR U63675 ( .A(n50841), .B(n50840), .Z(n50845) );
  IV U63676 ( .A(n50845), .Z(n50842) );
  NOR U63677 ( .A(n52208), .B(n50842), .Z(n52203) );
  IV U63678 ( .A(n50843), .Z(n52207) );
  XOR U63679 ( .A(n52207), .B(n52208), .Z(n50844) );
  NOR U63680 ( .A(n50845), .B(n50844), .Z(n52206) );
  NOR U63681 ( .A(n52203), .B(n52206), .Z(n52199) );
  XOR U63682 ( .A(n50846), .B(n52199), .Z(n52197) );
  XOR U63683 ( .A(n50847), .B(n52197), .Z(n52188) );
  XOR U63684 ( .A(n54409), .B(n52188), .Z(n52186) );
  XOR U63685 ( .A(n50848), .B(n52186), .Z(n52173) );
  XOR U63686 ( .A(n50849), .B(n52173), .Z(n52182) );
  XOR U63687 ( .A(n50850), .B(n52182), .Z(n54421) );
  XOR U63688 ( .A(n50851), .B(n54421), .Z(n54419) );
  XOR U63689 ( .A(n54418), .B(n54419), .Z(n52167) );
  XOR U63690 ( .A(n50852), .B(n52167), .Z(n54434) );
  XOR U63691 ( .A(n50853), .B(n54434), .Z(n54445) );
  XOR U63692 ( .A(n50854), .B(n54445), .Z(n50855) );
  IV U63693 ( .A(n50855), .Z(n52151) );
  XOR U63694 ( .A(n52149), .B(n52151), .Z(n52153) );
  XOR U63695 ( .A(n52152), .B(n52153), .Z(n52159) );
  IV U63696 ( .A(n50856), .Z(n50857) );
  NOR U63697 ( .A(n50858), .B(n50857), .Z(n52157) );
  XOR U63698 ( .A(n52159), .B(n52157), .Z(n52145) );
  IV U63699 ( .A(n50859), .Z(n50861) );
  NOR U63700 ( .A(n50861), .B(n50860), .Z(n52143) );
  XOR U63701 ( .A(n52145), .B(n52143), .Z(n52138) );
  IV U63702 ( .A(n50862), .Z(n52140) );
  NOR U63703 ( .A(n52140), .B(n50863), .Z(n50867) );
  IV U63704 ( .A(n50864), .Z(n50866) );
  NOR U63705 ( .A(n50866), .B(n50865), .Z(n52136) );
  NOR U63706 ( .A(n50867), .B(n52136), .Z(n50868) );
  XOR U63707 ( .A(n52138), .B(n50868), .Z(n50869) );
  IV U63708 ( .A(n50869), .Z(n52135) );
  XOR U63709 ( .A(n52132), .B(n52135), .Z(n52131) );
  NOR U63710 ( .A(n50870), .B(n52128), .Z(n50871) );
  NOR U63711 ( .A(n52133), .B(n50871), .Z(n50872) );
  XOR U63712 ( .A(n52131), .B(n50872), .Z(n54452) );
  IV U63713 ( .A(n50873), .Z(n50874) );
  NOR U63714 ( .A(n50875), .B(n50874), .Z(n54455) );
  IV U63715 ( .A(n50876), .Z(n50878) );
  NOR U63716 ( .A(n50878), .B(n50877), .Z(n54451) );
  NOR U63717 ( .A(n54455), .B(n54451), .Z(n50879) );
  XOR U63718 ( .A(n54452), .B(n50879), .Z(n52124) );
  XOR U63719 ( .A(n52123), .B(n52124), .Z(n54462) );
  XOR U63720 ( .A(n54461), .B(n54462), .Z(n54466) );
  XOR U63721 ( .A(n54464), .B(n54466), .Z(n52120) );
  IV U63722 ( .A(n50880), .Z(n50881) );
  NOR U63723 ( .A(n50882), .B(n50881), .Z(n50887) );
  IV U63724 ( .A(n50883), .Z(n50885) );
  NOR U63725 ( .A(n50885), .B(n50884), .Z(n50886) );
  NOR U63726 ( .A(n50887), .B(n50886), .Z(n52121) );
  XOR U63727 ( .A(n52120), .B(n52121), .Z(n50888) );
  NOR U63728 ( .A(n50889), .B(n50888), .Z(n52117) );
  IV U63729 ( .A(n50889), .Z(n50890) );
  NOR U63730 ( .A(n50890), .B(n52120), .Z(n52119) );
  NOR U63731 ( .A(n52117), .B(n52119), .Z(n54472) );
  XOR U63732 ( .A(n50891), .B(n54472), .Z(n54471) );
  XOR U63733 ( .A(n54469), .B(n54471), .Z(n54480) );
  XOR U63734 ( .A(n54479), .B(n54480), .Z(n50892) );
  XOR U63735 ( .A(n50893), .B(n50892), .Z(n52113) );
  IV U63736 ( .A(n50894), .Z(n50896) );
  NOR U63737 ( .A(n50896), .B(n50895), .Z(n50897) );
  IV U63738 ( .A(n50897), .Z(n52108) );
  XOR U63739 ( .A(n52113), .B(n52108), .Z(n52110) );
  XOR U63740 ( .A(n52111), .B(n52110), .Z(n52099) );
  IV U63741 ( .A(n52099), .Z(n52097) );
  NOR U63742 ( .A(n50899), .B(n50898), .Z(n50900) );
  IV U63743 ( .A(n50900), .Z(n52102) );
  NOR U63744 ( .A(n50901), .B(n52102), .Z(n50905) );
  IV U63745 ( .A(n50902), .Z(n50904) );
  NOR U63746 ( .A(n50904), .B(n50903), .Z(n52098) );
  XOR U63747 ( .A(n50905), .B(n52098), .Z(n50906) );
  XOR U63748 ( .A(n52097), .B(n50906), .Z(n52087) );
  XOR U63749 ( .A(n52086), .B(n52087), .Z(n52090) );
  XOR U63750 ( .A(n52089), .B(n52090), .Z(n52084) );
  XOR U63751 ( .A(n52083), .B(n52084), .Z(n52074) );
  XOR U63752 ( .A(n50907), .B(n52074), .Z(n54487) );
  XOR U63753 ( .A(n50908), .B(n54487), .Z(n54489) );
  IV U63754 ( .A(n54489), .Z(n54492) );
  XOR U63755 ( .A(n54490), .B(n54492), .Z(n54498) );
  IV U63756 ( .A(n50909), .Z(n50910) );
  NOR U63757 ( .A(n50911), .B(n50910), .Z(n54494) );
  NOR U63758 ( .A(n50912), .B(n54499), .Z(n50913) );
  NOR U63759 ( .A(n54494), .B(n50913), .Z(n50914) );
  XOR U63760 ( .A(n54498), .B(n50914), .Z(n50915) );
  IV U63761 ( .A(n50915), .Z(n52066) );
  IV U63762 ( .A(n50916), .Z(n50917) );
  NOR U63763 ( .A(n50918), .B(n50917), .Z(n50919) );
  IV U63764 ( .A(n50919), .Z(n50925) );
  NOR U63765 ( .A(n52066), .B(n50925), .Z(n55646) );
  IV U63766 ( .A(n50920), .Z(n52065) );
  NOR U63767 ( .A(n50921), .B(n52065), .Z(n50922) );
  XOR U63768 ( .A(n50922), .B(n52066), .Z(n54507) );
  IV U63769 ( .A(n50923), .Z(n50924) );
  NOR U63770 ( .A(n50924), .B(n50931), .Z(n50926) );
  IV U63771 ( .A(n50926), .Z(n54506) );
  XOR U63772 ( .A(n54507), .B(n54506), .Z(n50928) );
  NOR U63773 ( .A(n50926), .B(n50925), .Z(n50927) );
  NOR U63774 ( .A(n50928), .B(n50927), .Z(n50929) );
  NOR U63775 ( .A(n55646), .B(n50929), .Z(n54508) );
  IV U63776 ( .A(n50930), .Z(n50932) );
  NOR U63777 ( .A(n50932), .B(n50931), .Z(n54509) );
  XOR U63778 ( .A(n54508), .B(n54509), .Z(n50939) );
  IV U63779 ( .A(n50939), .Z(n50937) );
  IV U63780 ( .A(n50933), .Z(n50934) );
  NOR U63781 ( .A(n50935), .B(n50934), .Z(n50938) );
  IV U63782 ( .A(n50938), .Z(n50936) );
  NOR U63783 ( .A(n50937), .B(n50936), .Z(n55639) );
  NOR U63784 ( .A(n50939), .B(n50938), .Z(n52063) );
  NOR U63785 ( .A(n55639), .B(n52063), .Z(n58215) );
  XOR U63786 ( .A(n58217), .B(n58215), .Z(n52050) );
  XOR U63787 ( .A(n52047), .B(n52050), .Z(n52045) );
  IV U63788 ( .A(n50940), .Z(n52051) );
  NOR U63789 ( .A(n50941), .B(n52051), .Z(n50945) );
  IV U63790 ( .A(n50942), .Z(n50943) );
  NOR U63791 ( .A(n50944), .B(n50943), .Z(n52044) );
  NOR U63792 ( .A(n50945), .B(n52044), .Z(n50946) );
  XOR U63793 ( .A(n52045), .B(n50946), .Z(n52041) );
  IV U63794 ( .A(n50947), .Z(n50948) );
  NOR U63795 ( .A(n50949), .B(n50948), .Z(n50953) );
  IV U63796 ( .A(n50950), .Z(n50951) );
  NOR U63797 ( .A(n50956), .B(n50951), .Z(n50952) );
  NOR U63798 ( .A(n50953), .B(n50952), .Z(n52042) );
  XOR U63799 ( .A(n52041), .B(n52042), .Z(n52031) );
  IV U63800 ( .A(n50954), .Z(n50955) );
  NOR U63801 ( .A(n50956), .B(n50955), .Z(n52029) );
  XOR U63802 ( .A(n52031), .B(n52029), .Z(n52034) );
  IV U63803 ( .A(n50957), .Z(n50958) );
  NOR U63804 ( .A(n50959), .B(n50958), .Z(n52032) );
  XOR U63805 ( .A(n52034), .B(n52032), .Z(n52039) );
  IV U63806 ( .A(n50960), .Z(n50966) );
  IV U63807 ( .A(n50961), .Z(n50962) );
  NOR U63808 ( .A(n50966), .B(n50962), .Z(n52037) );
  XOR U63809 ( .A(n52039), .B(n52037), .Z(n52027) );
  NOR U63810 ( .A(n50963), .B(n52027), .Z(n55672) );
  IV U63811 ( .A(n50964), .Z(n50965) );
  NOR U63812 ( .A(n50966), .B(n50965), .Z(n52025) );
  XOR U63813 ( .A(n52027), .B(n52025), .Z(n50972) );
  IV U63814 ( .A(n50972), .Z(n50967) );
  NOR U63815 ( .A(n50968), .B(n50967), .Z(n50969) );
  NOR U63816 ( .A(n55672), .B(n50969), .Z(n50970) );
  NOR U63817 ( .A(n50971), .B(n50970), .Z(n50974) );
  IV U63818 ( .A(n50971), .Z(n50973) );
  NOR U63819 ( .A(n50973), .B(n50972), .Z(n55677) );
  NOR U63820 ( .A(n50974), .B(n55677), .Z(n52022) );
  XOR U63821 ( .A(n52024), .B(n52022), .Z(n54522) );
  XOR U63822 ( .A(n50975), .B(n54522), .Z(n52017) );
  IV U63823 ( .A(n50976), .Z(n50978) );
  NOR U63824 ( .A(n50978), .B(n50977), .Z(n50979) );
  IV U63825 ( .A(n50979), .Z(n50980) );
  NOR U63826 ( .A(n50981), .B(n50980), .Z(n52018) );
  NOR U63827 ( .A(n54524), .B(n52018), .Z(n50982) );
  XOR U63828 ( .A(n52017), .B(n50982), .Z(n52015) );
  XOR U63829 ( .A(n52007), .B(n52015), .Z(n52005) );
  XOR U63830 ( .A(n50983), .B(n52005), .Z(n50984) );
  IV U63831 ( .A(n50984), .Z(n52000) );
  IV U63832 ( .A(n50985), .Z(n50986) );
  NOR U63833 ( .A(n50987), .B(n50986), .Z(n51998) );
  XOR U63834 ( .A(n52000), .B(n51998), .Z(n51992) );
  IV U63835 ( .A(n51992), .Z(n50994) );
  IV U63836 ( .A(n50988), .Z(n50990) );
  NOR U63837 ( .A(n50990), .B(n50989), .Z(n51993) );
  IV U63838 ( .A(n50991), .Z(n50992) );
  NOR U63839 ( .A(n50992), .B(n50999), .Z(n51990) );
  NOR U63840 ( .A(n51993), .B(n51990), .Z(n50993) );
  XOR U63841 ( .A(n50994), .B(n50993), .Z(n51989) );
  IV U63842 ( .A(n50995), .Z(n51003) );
  NOR U63843 ( .A(n51003), .B(n50996), .Z(n51985) );
  IV U63844 ( .A(n50997), .Z(n50998) );
  NOR U63845 ( .A(n50999), .B(n50998), .Z(n51987) );
  NOR U63846 ( .A(n51985), .B(n51987), .Z(n51000) );
  XOR U63847 ( .A(n51989), .B(n51000), .Z(n51979) );
  IV U63848 ( .A(n51979), .Z(n51976) );
  XOR U63849 ( .A(n51980), .B(n51976), .Z(n51975) );
  IV U63850 ( .A(n51975), .Z(n51007) );
  IV U63851 ( .A(n51001), .Z(n51002) );
  NOR U63852 ( .A(n51003), .B(n51002), .Z(n51978) );
  IV U63853 ( .A(n51004), .Z(n51005) );
  NOR U63854 ( .A(n51005), .B(n51009), .Z(n51973) );
  NOR U63855 ( .A(n51978), .B(n51973), .Z(n51006) );
  XOR U63856 ( .A(n51007), .B(n51006), .Z(n51972) );
  IV U63857 ( .A(n51008), .Z(n51010) );
  NOR U63858 ( .A(n51010), .B(n51009), .Z(n51970) );
  XOR U63859 ( .A(n51972), .B(n51970), .Z(n54529) );
  XOR U63860 ( .A(n51011), .B(n54529), .Z(n51961) );
  XOR U63861 ( .A(n51012), .B(n51961), .Z(n51013) );
  IV U63862 ( .A(n51013), .Z(n54537) );
  XOR U63863 ( .A(n54535), .B(n54537), .Z(n54532) );
  NOR U63864 ( .A(n51014), .B(n54532), .Z(n55547) );
  IV U63865 ( .A(n51015), .Z(n51016) );
  NOR U63866 ( .A(n51017), .B(n51016), .Z(n54531) );
  XOR U63867 ( .A(n54531), .B(n54532), .Z(n51023) );
  IV U63868 ( .A(n51023), .Z(n51018) );
  NOR U63869 ( .A(n51019), .B(n51018), .Z(n51020) );
  NOR U63870 ( .A(n55547), .B(n51020), .Z(n51021) );
  NOR U63871 ( .A(n51022), .B(n51021), .Z(n54546) );
  IV U63872 ( .A(n51022), .Z(n51024) );
  NOR U63873 ( .A(n51024), .B(n51023), .Z(n54544) );
  NOR U63874 ( .A(n54546), .B(n54544), .Z(n51025) );
  IV U63875 ( .A(n51025), .Z(n51956) );
  IV U63876 ( .A(n51026), .Z(n51028) );
  NOR U63877 ( .A(n51028), .B(n51027), .Z(n51955) );
  IV U63878 ( .A(n51029), .Z(n51031) );
  NOR U63879 ( .A(n51031), .B(n51030), .Z(n54543) );
  NOR U63880 ( .A(n51955), .B(n54543), .Z(n51032) );
  XOR U63881 ( .A(n51956), .B(n51032), .Z(n51042) );
  IV U63882 ( .A(n51033), .Z(n51034) );
  NOR U63883 ( .A(n51035), .B(n51034), .Z(n51952) );
  IV U63884 ( .A(n51036), .Z(n51038) );
  NOR U63885 ( .A(n51038), .B(n51037), .Z(n51946) );
  NOR U63886 ( .A(n51952), .B(n51946), .Z(n51039) );
  XOR U63887 ( .A(n51042), .B(n51039), .Z(n51948) );
  XOR U63888 ( .A(n51949), .B(n51948), .Z(n51040) );
  NOR U63889 ( .A(n51041), .B(n51040), .Z(n51045) );
  IV U63890 ( .A(n51041), .Z(n51044) );
  IV U63891 ( .A(n51042), .Z(n51954) );
  XOR U63892 ( .A(n51952), .B(n51954), .Z(n51043) );
  NOR U63893 ( .A(n51044), .B(n51043), .Z(n55521) );
  NOR U63894 ( .A(n51045), .B(n55521), .Z(n51944) );
  XOR U63895 ( .A(n51046), .B(n51944), .Z(n54550) );
  XOR U63896 ( .A(n54548), .B(n54550), .Z(n51941) );
  IV U63897 ( .A(n51047), .Z(n51049) );
  NOR U63898 ( .A(n51049), .B(n51048), .Z(n51940) );
  IV U63899 ( .A(n51050), .Z(n51051) );
  NOR U63900 ( .A(n51051), .B(n51054), .Z(n51938) );
  NOR U63901 ( .A(n51940), .B(n51938), .Z(n51052) );
  XOR U63902 ( .A(n51941), .B(n51052), .Z(n51936) );
  IV U63903 ( .A(n51053), .Z(n51055) );
  NOR U63904 ( .A(n51055), .B(n51054), .Z(n51933) );
  IV U63905 ( .A(n51056), .Z(n54573) );
  NOR U63906 ( .A(n51057), .B(n54573), .Z(n54574) );
  NOR U63907 ( .A(n51933), .B(n54574), .Z(n51058) );
  XOR U63908 ( .A(n51936), .B(n51058), .Z(n51930) );
  IV U63909 ( .A(n51059), .Z(n51060) );
  NOR U63910 ( .A(n51061), .B(n51060), .Z(n51932) );
  IV U63911 ( .A(n51062), .Z(n51064) );
  NOR U63912 ( .A(n51064), .B(n51063), .Z(n51929) );
  NOR U63913 ( .A(n51932), .B(n51929), .Z(n51065) );
  XOR U63914 ( .A(n51930), .B(n51065), .Z(n51926) );
  IV U63915 ( .A(n51066), .Z(n51068) );
  NOR U63916 ( .A(n51068), .B(n51067), .Z(n51069) );
  IV U63917 ( .A(n51069), .Z(n51927) );
  XOR U63918 ( .A(n51926), .B(n51927), .Z(n51915) );
  XOR U63919 ( .A(n51914), .B(n51915), .Z(n51919) );
  XOR U63920 ( .A(n51917), .B(n51919), .Z(n51925) );
  XOR U63921 ( .A(n51923), .B(n51925), .Z(n51076) );
  NOR U63922 ( .A(n51078), .B(n51076), .Z(n58314) );
  IV U63923 ( .A(n51070), .Z(n51072) );
  NOR U63924 ( .A(n51072), .B(n51071), .Z(n51073) );
  IV U63925 ( .A(n51073), .Z(n51906) );
  IV U63926 ( .A(n51074), .Z(n51908) );
  NOR U63927 ( .A(n51908), .B(n51075), .Z(n51077) );
  XOR U63928 ( .A(n51077), .B(n51076), .Z(n51905) );
  XOR U63929 ( .A(n51906), .B(n51905), .Z(n51081) );
  IV U63930 ( .A(n51905), .Z(n51079) );
  NOR U63931 ( .A(n51079), .B(n51078), .Z(n51080) );
  NOR U63932 ( .A(n51081), .B(n51080), .Z(n51082) );
  NOR U63933 ( .A(n58314), .B(n51082), .Z(n51083) );
  IV U63934 ( .A(n51083), .Z(n51898) );
  IV U63935 ( .A(n51084), .Z(n51086) );
  NOR U63936 ( .A(n51086), .B(n51085), .Z(n51897) );
  XOR U63937 ( .A(n51898), .B(n51897), .Z(n51901) );
  XOR U63938 ( .A(n51900), .B(n51901), .Z(n51894) );
  IV U63939 ( .A(n51089), .Z(n51087) );
  NOR U63940 ( .A(n51088), .B(n51087), .Z(n51093) );
  IV U63941 ( .A(n51088), .Z(n51880) );
  NOR U63942 ( .A(n51089), .B(n51880), .Z(n51091) );
  NOR U63943 ( .A(n51091), .B(n51090), .Z(n51092) );
  NOR U63944 ( .A(n51093), .B(n51092), .Z(n51094) );
  XOR U63945 ( .A(n51894), .B(n51094), .Z(n51095) );
  XOR U63946 ( .A(n51096), .B(n51095), .Z(n51876) );
  XOR U63947 ( .A(n51097), .B(n51876), .Z(n51869) );
  XOR U63948 ( .A(n51098), .B(n51869), .Z(n54600) );
  IV U63949 ( .A(n51099), .Z(n51100) );
  NOR U63950 ( .A(n51101), .B(n51100), .Z(n54599) );
  IV U63951 ( .A(n51102), .Z(n51103) );
  NOR U63952 ( .A(n51104), .B(n51103), .Z(n51864) );
  NOR U63953 ( .A(n54599), .B(n51864), .Z(n51105) );
  XOR U63954 ( .A(n54600), .B(n51105), .Z(n54605) );
  IV U63955 ( .A(n51106), .Z(n51108) );
  NOR U63956 ( .A(n51108), .B(n51107), .Z(n54603) );
  XOR U63957 ( .A(n54605), .B(n54603), .Z(n54607) );
  XOR U63958 ( .A(n54606), .B(n54607), .Z(n51115) );
  IV U63959 ( .A(n51115), .Z(n51109) );
  NOR U63960 ( .A(n51110), .B(n51109), .Z(n58364) );
  IV U63961 ( .A(n51111), .Z(n51121) );
  IV U63962 ( .A(n51112), .Z(n51113) );
  NOR U63963 ( .A(n51121), .B(n51113), .Z(n51116) );
  IV U63964 ( .A(n51116), .Z(n51114) );
  NOR U63965 ( .A(n51114), .B(n54607), .Z(n54612) );
  NOR U63966 ( .A(n51116), .B(n51115), .Z(n51117) );
  NOR U63967 ( .A(n54612), .B(n51117), .Z(n51118) );
  IV U63968 ( .A(n51118), .Z(n54610) );
  IV U63969 ( .A(n51119), .Z(n51120) );
  NOR U63970 ( .A(n51121), .B(n51120), .Z(n51122) );
  IV U63971 ( .A(n51122), .Z(n54609) );
  XOR U63972 ( .A(n54610), .B(n54609), .Z(n51123) );
  NOR U63973 ( .A(n51124), .B(n51123), .Z(n51125) );
  NOR U63974 ( .A(n58364), .B(n51125), .Z(n51126) );
  IV U63975 ( .A(n51126), .Z(n54616) );
  XOR U63976 ( .A(n54615), .B(n54616), .Z(n54621) );
  IV U63977 ( .A(n51127), .Z(n51135) );
  IV U63978 ( .A(n51128), .Z(n51129) );
  NOR U63979 ( .A(n51135), .B(n51129), .Z(n54619) );
  XOR U63980 ( .A(n54621), .B(n54619), .Z(n54622) );
  IV U63981 ( .A(n54622), .Z(n51138) );
  IV U63982 ( .A(n51130), .Z(n51132) );
  NOR U63983 ( .A(n51132), .B(n51131), .Z(n51137) );
  IV U63984 ( .A(n51133), .Z(n51134) );
  NOR U63985 ( .A(n51135), .B(n51134), .Z(n51136) );
  NOR U63986 ( .A(n51137), .B(n51136), .Z(n54623) );
  XOR U63987 ( .A(n51138), .B(n54623), .Z(n54628) );
  XOR U63988 ( .A(n54627), .B(n54628), .Z(n54625) );
  XOR U63989 ( .A(n54626), .B(n54625), .Z(n51139) );
  IV U63990 ( .A(n51139), .Z(n54640) );
  XOR U63991 ( .A(n51856), .B(n54640), .Z(n51140) );
  XOR U63992 ( .A(n51141), .B(n51140), .Z(n51850) );
  IV U63993 ( .A(n51142), .Z(n51144) );
  NOR U63994 ( .A(n51144), .B(n51143), .Z(n51848) );
  XOR U63995 ( .A(n51850), .B(n51848), .Z(n51853) );
  XOR U63996 ( .A(n51851), .B(n51853), .Z(n51846) );
  XOR U63997 ( .A(n51145), .B(n51846), .Z(n51835) );
  XOR U63998 ( .A(n51146), .B(n51835), .Z(n54647) );
  XOR U63999 ( .A(n54646), .B(n54647), .Z(n54650) );
  XOR U64000 ( .A(n54651), .B(n54650), .Z(n51148) );
  NOR U64001 ( .A(n51147), .B(n51148), .Z(n54657) );
  IV U64002 ( .A(n51147), .Z(n51150) );
  IV U64003 ( .A(n51148), .Z(n51149) );
  NOR U64004 ( .A(n51150), .B(n51149), .Z(n55439) );
  NOR U64005 ( .A(n54657), .B(n55439), .Z(n51828) );
  XOR U64006 ( .A(n51832), .B(n51828), .Z(n54663) );
  XOR U64007 ( .A(n51151), .B(n54663), .Z(n51826) );
  XOR U64008 ( .A(n51152), .B(n51826), .Z(n51814) );
  IV U64009 ( .A(n51814), .Z(n51816) );
  XOR U64010 ( .A(n51815), .B(n51816), .Z(n51813) );
  IV U64011 ( .A(n51813), .Z(n51160) );
  IV U64012 ( .A(n51153), .Z(n51158) );
  IV U64013 ( .A(n51154), .Z(n51155) );
  NOR U64014 ( .A(n51156), .B(n51155), .Z(n51157) );
  IV U64015 ( .A(n51157), .Z(n51162) );
  NOR U64016 ( .A(n51158), .B(n51162), .Z(n51811) );
  NOR U64017 ( .A(n51819), .B(n51811), .Z(n51159) );
  XOR U64018 ( .A(n51160), .B(n51159), .Z(n51807) );
  IV U64019 ( .A(n51161), .Z(n51163) );
  NOR U64020 ( .A(n51163), .B(n51162), .Z(n51805) );
  XOR U64021 ( .A(n51807), .B(n51805), .Z(n51810) );
  XOR U64022 ( .A(n51808), .B(n51810), .Z(n54690) );
  XOR U64023 ( .A(n51164), .B(n54690), .Z(n51165) );
  IV U64024 ( .A(n51165), .Z(n51797) );
  XOR U64025 ( .A(n51795), .B(n51797), .Z(n54692) );
  XOR U64026 ( .A(n54691), .B(n54692), .Z(n54695) );
  IV U64027 ( .A(n54695), .Z(n51172) );
  IV U64028 ( .A(n51166), .Z(n51167) );
  NOR U64029 ( .A(n51168), .B(n51167), .Z(n54694) );
  NOR U64030 ( .A(n51170), .B(n51169), .Z(n51793) );
  NOR U64031 ( .A(n54694), .B(n51793), .Z(n51171) );
  XOR U64032 ( .A(n51172), .B(n51171), .Z(n54701) );
  XOR U64033 ( .A(n54699), .B(n54701), .Z(n54704) );
  XOR U64034 ( .A(n54702), .B(n54704), .Z(n54709) );
  XOR U64035 ( .A(n51173), .B(n54709), .Z(n51174) );
  IV U64036 ( .A(n51174), .Z(n54715) );
  XOR U64037 ( .A(n54706), .B(n54715), .Z(n55391) );
  IV U64038 ( .A(n54712), .Z(n58402) );
  NOR U64039 ( .A(n58402), .B(n54714), .Z(n51177) );
  NOR U64040 ( .A(n51176), .B(n51175), .Z(n55389) );
  NOR U64041 ( .A(n51177), .B(n55389), .Z(n51178) );
  XOR U64042 ( .A(n55391), .B(n51178), .Z(n51787) );
  IV U64043 ( .A(n51179), .Z(n51180) );
  NOR U64044 ( .A(n51186), .B(n51180), .Z(n54720) );
  IV U64045 ( .A(n51181), .Z(n51183) );
  NOR U64046 ( .A(n51183), .B(n51182), .Z(n51788) );
  NOR U64047 ( .A(n54720), .B(n51788), .Z(n51184) );
  XOR U64048 ( .A(n51787), .B(n51184), .Z(n54729) );
  IV U64049 ( .A(n51185), .Z(n51189) );
  NOR U64050 ( .A(n51187), .B(n51186), .Z(n51188) );
  IV U64051 ( .A(n51188), .Z(n51191) );
  NOR U64052 ( .A(n51189), .B(n51191), .Z(n54727) );
  XOR U64053 ( .A(n54729), .B(n54727), .Z(n54732) );
  IV U64054 ( .A(n51190), .Z(n51192) );
  NOR U64055 ( .A(n51192), .B(n51191), .Z(n54730) );
  XOR U64056 ( .A(n54732), .B(n54730), .Z(n51785) );
  XOR U64057 ( .A(n51786), .B(n51785), .Z(n51780) );
  IV U64058 ( .A(n51193), .Z(n51194) );
  NOR U64059 ( .A(n51195), .B(n51194), .Z(n51783) );
  IV U64060 ( .A(n51196), .Z(n51197) );
  NOR U64061 ( .A(n51198), .B(n51197), .Z(n51779) );
  NOR U64062 ( .A(n51783), .B(n51779), .Z(n51199) );
  XOR U64063 ( .A(n51780), .B(n51199), .Z(n51776) );
  IV U64064 ( .A(n51200), .Z(n51202) );
  NOR U64065 ( .A(n51202), .B(n51201), .Z(n51203) );
  IV U64066 ( .A(n51203), .Z(n51211) );
  NOR U64067 ( .A(n51776), .B(n51211), .Z(n51777) );
  IV U64068 ( .A(n51204), .Z(n51206) );
  NOR U64069 ( .A(n51206), .B(n51205), .Z(n51207) );
  IV U64070 ( .A(n51207), .Z(n51773) );
  IV U64071 ( .A(n51208), .Z(n51210) );
  NOR U64072 ( .A(n51210), .B(n51209), .Z(n51774) );
  XOR U64073 ( .A(n51774), .B(n51776), .Z(n51772) );
  XOR U64074 ( .A(n51773), .B(n51772), .Z(n51214) );
  IV U64075 ( .A(n51772), .Z(n51212) );
  NOR U64076 ( .A(n51212), .B(n51211), .Z(n51213) );
  NOR U64077 ( .A(n51214), .B(n51213), .Z(n51215) );
  NOR U64078 ( .A(n51777), .B(n51215), .Z(n51216) );
  IV U64079 ( .A(n51216), .Z(n54737) );
  XOR U64080 ( .A(n54736), .B(n54737), .Z(n54740) );
  XOR U64081 ( .A(n54739), .B(n54740), .Z(n51765) );
  XOR U64082 ( .A(n51764), .B(n51765), .Z(n51769) );
  IV U64083 ( .A(n51217), .Z(n51221) );
  IV U64084 ( .A(n51218), .Z(n51219) );
  NOR U64085 ( .A(n51221), .B(n51219), .Z(n51767) );
  XOR U64086 ( .A(n51769), .B(n51767), .Z(n51759) );
  IV U64087 ( .A(n51759), .Z(n51757) );
  IV U64088 ( .A(n51220), .Z(n51224) );
  NOR U64089 ( .A(n51222), .B(n51221), .Z(n51223) );
  IV U64090 ( .A(n51223), .Z(n51229) );
  NOR U64091 ( .A(n51224), .B(n51229), .Z(n51756) );
  IV U64092 ( .A(n51756), .Z(n51758) );
  XOR U64093 ( .A(n51757), .B(n51758), .Z(n51754) );
  IV U64094 ( .A(n51225), .Z(n51227) );
  NOR U64095 ( .A(n51227), .B(n51226), .Z(n51753) );
  IV U64096 ( .A(n51228), .Z(n51230) );
  NOR U64097 ( .A(n51230), .B(n51229), .Z(n51760) );
  NOR U64098 ( .A(n51753), .B(n51760), .Z(n51231) );
  XOR U64099 ( .A(n51754), .B(n51231), .Z(n51232) );
  IV U64100 ( .A(n51232), .Z(n51752) );
  IV U64101 ( .A(n51233), .Z(n51235) );
  NOR U64102 ( .A(n51235), .B(n51234), .Z(n51236) );
  IV U64103 ( .A(n51236), .Z(n51751) );
  XOR U64104 ( .A(n51752), .B(n51751), .Z(n51744) );
  XOR U64105 ( .A(n51746), .B(n51744), .Z(n51741) );
  XOR U64106 ( .A(n51237), .B(n51741), .Z(n51737) );
  XOR U64107 ( .A(n51238), .B(n51737), .Z(n51732) );
  NOR U64108 ( .A(n51246), .B(n51732), .Z(n55247) );
  IV U64109 ( .A(n51239), .Z(n51240) );
  NOR U64110 ( .A(n51241), .B(n51240), .Z(n51242) );
  IV U64111 ( .A(n51242), .Z(n51734) );
  IV U64112 ( .A(n51243), .Z(n51245) );
  NOR U64113 ( .A(n51245), .B(n51244), .Z(n51730) );
  XOR U64114 ( .A(n51732), .B(n51730), .Z(n51733) );
  XOR U64115 ( .A(n51734), .B(n51733), .Z(n51249) );
  IV U64116 ( .A(n51733), .Z(n51247) );
  NOR U64117 ( .A(n51247), .B(n51246), .Z(n51248) );
  NOR U64118 ( .A(n51249), .B(n51248), .Z(n51250) );
  NOR U64119 ( .A(n55247), .B(n51250), .Z(n54754) );
  IV U64120 ( .A(n51251), .Z(n51253) );
  NOR U64121 ( .A(n51253), .B(n51252), .Z(n51728) );
  IV U64122 ( .A(n51254), .Z(n51255) );
  NOR U64123 ( .A(n51255), .B(n51258), .Z(n54753) );
  NOR U64124 ( .A(n51728), .B(n54753), .Z(n51256) );
  XOR U64125 ( .A(n54754), .B(n51256), .Z(n54761) );
  IV U64126 ( .A(n51257), .Z(n51259) );
  NOR U64127 ( .A(n51259), .B(n51258), .Z(n54759) );
  IV U64128 ( .A(n51260), .Z(n51262) );
  IV U64129 ( .A(n51261), .Z(n51266) );
  NOR U64130 ( .A(n51262), .B(n51266), .Z(n51726) );
  NOR U64131 ( .A(n54759), .B(n51726), .Z(n51263) );
  XOR U64132 ( .A(n54761), .B(n51263), .Z(n51722) );
  IV U64133 ( .A(n51264), .Z(n51265) );
  NOR U64134 ( .A(n51266), .B(n51265), .Z(n51718) );
  IV U64135 ( .A(n51267), .Z(n51269) );
  NOR U64136 ( .A(n51269), .B(n51268), .Z(n51721) );
  NOR U64137 ( .A(n51718), .B(n51721), .Z(n51270) );
  XOR U64138 ( .A(n51722), .B(n51270), .Z(n51716) );
  XOR U64139 ( .A(n51271), .B(n51716), .Z(n54764) );
  IV U64140 ( .A(n54764), .Z(n54767) );
  XOR U64141 ( .A(n54765), .B(n54767), .Z(n51713) );
  IV U64142 ( .A(n51713), .Z(n51278) );
  IV U64143 ( .A(n51272), .Z(n51273) );
  NOR U64144 ( .A(n51276), .B(n51273), .Z(n54769) );
  IV U64145 ( .A(n51274), .Z(n51275) );
  NOR U64146 ( .A(n51276), .B(n51275), .Z(n51711) );
  NOR U64147 ( .A(n54769), .B(n51711), .Z(n51277) );
  XOR U64148 ( .A(n51278), .B(n51277), .Z(n51710) );
  IV U64149 ( .A(n51279), .Z(n51281) );
  NOR U64150 ( .A(n51281), .B(n51280), .Z(n51708) );
  XOR U64151 ( .A(n51710), .B(n51708), .Z(n51704) );
  XOR U64152 ( .A(n51282), .B(n51704), .Z(n51283) );
  IV U64153 ( .A(n51283), .Z(n51702) );
  XOR U64154 ( .A(n51284), .B(n51702), .Z(n54774) );
  XOR U64155 ( .A(n54773), .B(n54774), .Z(n51696) );
  XOR U64156 ( .A(n51285), .B(n51696), .Z(n51286) );
  IV U64157 ( .A(n51286), .Z(n54787) );
  XOR U64158 ( .A(n54785), .B(n54787), .Z(n54790) );
  IV U64159 ( .A(n54790), .Z(n51295) );
  IV U64160 ( .A(n51287), .Z(n51288) );
  NOR U64161 ( .A(n51289), .B(n51288), .Z(n51294) );
  NOR U64162 ( .A(n51295), .B(n51294), .Z(n51293) );
  IV U64163 ( .A(n51290), .Z(n51291) );
  NOR U64164 ( .A(n51298), .B(n51291), .Z(n51301) );
  IV U64165 ( .A(n51301), .Z(n51292) );
  NOR U64166 ( .A(n51293), .B(n51292), .Z(n54791) );
  IV U64167 ( .A(n51294), .Z(n54789) );
  XOR U64168 ( .A(n51295), .B(n54789), .Z(n51693) );
  IV U64169 ( .A(n51296), .Z(n51297) );
  NOR U64170 ( .A(n51298), .B(n51297), .Z(n51299) );
  IV U64171 ( .A(n51299), .Z(n51692) );
  XOR U64172 ( .A(n51693), .B(n51692), .Z(n51300) );
  NOR U64173 ( .A(n51301), .B(n51300), .Z(n51302) );
  NOR U64174 ( .A(n54791), .B(n51302), .Z(n51688) );
  IV U64175 ( .A(n51303), .Z(n51305) );
  NOR U64176 ( .A(n51305), .B(n51304), .Z(n51306) );
  IV U64177 ( .A(n51306), .Z(n51690) );
  XOR U64178 ( .A(n51688), .B(n51690), .Z(n51685) );
  XOR U64179 ( .A(n51683), .B(n51685), .Z(n51307) );
  XOR U64180 ( .A(n51308), .B(n51307), .Z(n51682) );
  IV U64181 ( .A(n51309), .Z(n51310) );
  NOR U64182 ( .A(n51311), .B(n51310), .Z(n51680) );
  IV U64183 ( .A(n51312), .Z(n51314) );
  NOR U64184 ( .A(n51314), .B(n51313), .Z(n51678) );
  NOR U64185 ( .A(n51680), .B(n51678), .Z(n51315) );
  XOR U64186 ( .A(n51682), .B(n51315), .Z(n51675) );
  XOR U64187 ( .A(n51673), .B(n51675), .Z(n51667) );
  IV U64188 ( .A(n51316), .Z(n51318) );
  NOR U64189 ( .A(n51318), .B(n51317), .Z(n51674) );
  IV U64190 ( .A(n51319), .Z(n51321) );
  NOR U64191 ( .A(n51321), .B(n51320), .Z(n51668) );
  NOR U64192 ( .A(n51674), .B(n51668), .Z(n51322) );
  XOR U64193 ( .A(n51667), .B(n51322), .Z(n51666) );
  XOR U64194 ( .A(n51665), .B(n51666), .Z(n54796) );
  XOR U64195 ( .A(n54793), .B(n54796), .Z(n51664) );
  XOR U64196 ( .A(n51323), .B(n51664), .Z(n51653) );
  XOR U64197 ( .A(n51324), .B(n51653), .Z(n51646) );
  NOR U64198 ( .A(n51325), .B(n51646), .Z(n51644) );
  IV U64199 ( .A(n51326), .Z(n51327) );
  NOR U64200 ( .A(n51327), .B(n51329), .Z(n51648) );
  IV U64201 ( .A(n51328), .Z(n51330) );
  NOR U64202 ( .A(n51330), .B(n51329), .Z(n51645) );
  NOR U64203 ( .A(n51648), .B(n51645), .Z(n51331) );
  XOR U64204 ( .A(n51331), .B(n51646), .Z(n54805) );
  NOR U64205 ( .A(n51332), .B(n54805), .Z(n51333) );
  NOR U64206 ( .A(n51644), .B(n51333), .Z(n51334) );
  IV U64207 ( .A(n51334), .Z(n51641) );
  IV U64208 ( .A(n51335), .Z(n51341) );
  IV U64209 ( .A(n51336), .Z(n51337) );
  NOR U64210 ( .A(n51341), .B(n51337), .Z(n51338) );
  IV U64211 ( .A(n51338), .Z(n54806) );
  IV U64212 ( .A(n51339), .Z(n51340) );
  NOR U64213 ( .A(n51341), .B(n51340), .Z(n51342) );
  IV U64214 ( .A(n51342), .Z(n51642) );
  XOR U64215 ( .A(n54806), .B(n51642), .Z(n51343) );
  XOR U64216 ( .A(n51641), .B(n51343), .Z(n54803) );
  XOR U64217 ( .A(n54802), .B(n54803), .Z(n54811) );
  IV U64218 ( .A(n51344), .Z(n51346) );
  NOR U64219 ( .A(n51346), .B(n51345), .Z(n54809) );
  XOR U64220 ( .A(n54811), .B(n54809), .Z(n54812) );
  IV U64221 ( .A(n54812), .Z(n51354) );
  IV U64222 ( .A(n51347), .Z(n51351) );
  IV U64223 ( .A(n51348), .Z(n51349) );
  NOR U64224 ( .A(n51351), .B(n51349), .Z(n51353) );
  NOR U64225 ( .A(n51351), .B(n51350), .Z(n51352) );
  NOR U64226 ( .A(n51353), .B(n51352), .Z(n54813) );
  XOR U64227 ( .A(n51354), .B(n54813), .Z(n54817) );
  XOR U64228 ( .A(n54815), .B(n54817), .Z(n54820) );
  XOR U64229 ( .A(n54818), .B(n54820), .Z(n54824) );
  XOR U64230 ( .A(n54823), .B(n54824), .Z(n54827) );
  XOR U64231 ( .A(n54826), .B(n54827), .Z(n51635) );
  XOR U64232 ( .A(n51633), .B(n51635), .Z(n51638) );
  XOR U64233 ( .A(n51636), .B(n51638), .Z(n51631) );
  XOR U64234 ( .A(n51629), .B(n51631), .Z(n51628) );
  IV U64235 ( .A(n51355), .Z(n51360) );
  IV U64236 ( .A(n51356), .Z(n51357) );
  NOR U64237 ( .A(n51360), .B(n51357), .Z(n51626) );
  XOR U64238 ( .A(n51628), .B(n51626), .Z(n54832) );
  IV U64239 ( .A(n51358), .Z(n51359) );
  NOR U64240 ( .A(n51360), .B(n51359), .Z(n51361) );
  IV U64241 ( .A(n51361), .Z(n54831) );
  XOR U64242 ( .A(n54832), .B(n54831), .Z(n51362) );
  NOR U64243 ( .A(n51363), .B(n51362), .Z(n51373) );
  IV U64244 ( .A(n51364), .Z(n51367) );
  NOR U64245 ( .A(n51365), .B(n51628), .Z(n51366) );
  IV U64246 ( .A(n51366), .Z(n51369) );
  NOR U64247 ( .A(n51367), .B(n51369), .Z(n51624) );
  IV U64248 ( .A(n51368), .Z(n51370) );
  NOR U64249 ( .A(n51370), .B(n51369), .Z(n51625) );
  NOR U64250 ( .A(n51624), .B(n51625), .Z(n51371) );
  IV U64251 ( .A(n51371), .Z(n51372) );
  NOR U64252 ( .A(n51373), .B(n51372), .Z(n51617) );
  IV U64253 ( .A(n51374), .Z(n51376) );
  IV U64254 ( .A(n51375), .Z(n51380) );
  NOR U64255 ( .A(n51376), .B(n51380), .Z(n51377) );
  IV U64256 ( .A(n51377), .Z(n54846) );
  XOR U64257 ( .A(n51617), .B(n54846), .Z(n54843) );
  IV U64258 ( .A(n54843), .Z(n51384) );
  NOR U64259 ( .A(n51378), .B(n51618), .Z(n51382) );
  IV U64260 ( .A(n51379), .Z(n51381) );
  NOR U64261 ( .A(n51381), .B(n51380), .Z(n54841) );
  NOR U64262 ( .A(n51382), .B(n54841), .Z(n51383) );
  XOR U64263 ( .A(n51384), .B(n51383), .Z(n51615) );
  IV U64264 ( .A(n51385), .Z(n51387) );
  NOR U64265 ( .A(n51387), .B(n51386), .Z(n51613) );
  XOR U64266 ( .A(n51615), .B(n51613), .Z(n51607) );
  XOR U64267 ( .A(n51605), .B(n51607), .Z(n51609) );
  XOR U64268 ( .A(n51608), .B(n51609), .Z(n51603) );
  IV U64269 ( .A(n51388), .Z(n51598) );
  NOR U64270 ( .A(n51389), .B(n51598), .Z(n51592) );
  IV U64271 ( .A(n51390), .Z(n51391) );
  NOR U64272 ( .A(n51392), .B(n51391), .Z(n51602) );
  NOR U64273 ( .A(n51592), .B(n51602), .Z(n51393) );
  XOR U64274 ( .A(n51603), .B(n51393), .Z(n51394) );
  NOR U64275 ( .A(n51395), .B(n51394), .Z(n51398) );
  IV U64276 ( .A(n51395), .Z(n51397) );
  XOR U64277 ( .A(n51602), .B(n51603), .Z(n51396) );
  NOR U64278 ( .A(n51397), .B(n51396), .Z(n58621) );
  NOR U64279 ( .A(n51398), .B(n58621), .Z(n51585) );
  IV U64280 ( .A(n51399), .Z(n51401) );
  IV U64281 ( .A(n51400), .Z(n51405) );
  NOR U64282 ( .A(n51401), .B(n51405), .Z(n51402) );
  IV U64283 ( .A(n51402), .Z(n51586) );
  XOR U64284 ( .A(n51585), .B(n51586), .Z(n51590) );
  IV U64285 ( .A(n51590), .Z(n51409) );
  IV U64286 ( .A(n51403), .Z(n51404) );
  NOR U64287 ( .A(n51405), .B(n51404), .Z(n51588) );
  IV U64288 ( .A(n51406), .Z(n51407) );
  NOR U64289 ( .A(n51412), .B(n51407), .Z(n51581) );
  NOR U64290 ( .A(n51588), .B(n51581), .Z(n51408) );
  XOR U64291 ( .A(n51409), .B(n51408), .Z(n51580) );
  IV U64292 ( .A(n51410), .Z(n51411) );
  NOR U64293 ( .A(n51412), .B(n51411), .Z(n51578) );
  XOR U64294 ( .A(n51580), .B(n51578), .Z(n51572) );
  XOR U64295 ( .A(n51570), .B(n51572), .Z(n51575) );
  XOR U64296 ( .A(n51573), .B(n51575), .Z(n51568) );
  XOR U64297 ( .A(n51413), .B(n51568), .Z(n51414) );
  IV U64298 ( .A(n51414), .Z(n54860) );
  IV U64299 ( .A(n51415), .Z(n51417) );
  NOR U64300 ( .A(n51417), .B(n51416), .Z(n51563) );
  XOR U64301 ( .A(n54860), .B(n51563), .Z(n54866) );
  IV U64302 ( .A(n54866), .Z(n51425) );
  IV U64303 ( .A(n51418), .Z(n51419) );
  NOR U64304 ( .A(n51420), .B(n51419), .Z(n54859) );
  IV U64305 ( .A(n51421), .Z(n51422) );
  NOR U64306 ( .A(n51423), .B(n51422), .Z(n54865) );
  NOR U64307 ( .A(n54859), .B(n54865), .Z(n51424) );
  XOR U64308 ( .A(n51425), .B(n51424), .Z(n54863) );
  IV U64309 ( .A(n51426), .Z(n51429) );
  NOR U64310 ( .A(n51427), .B(n51432), .Z(n51428) );
  IV U64311 ( .A(n51428), .Z(n51435) );
  NOR U64312 ( .A(n51429), .B(n51435), .Z(n51438) );
  IV U64313 ( .A(n51438), .Z(n51430) );
  NOR U64314 ( .A(n54863), .B(n51430), .Z(n51560) );
  IV U64315 ( .A(n51431), .Z(n51433) );
  NOR U64316 ( .A(n51433), .B(n51432), .Z(n54862) );
  IV U64317 ( .A(n51434), .Z(n51436) );
  NOR U64318 ( .A(n51436), .B(n51435), .Z(n51561) );
  NOR U64319 ( .A(n54862), .B(n51561), .Z(n51437) );
  XOR U64320 ( .A(n54863), .B(n51437), .Z(n51554) );
  NOR U64321 ( .A(n51554), .B(n51438), .Z(n51439) );
  NOR U64322 ( .A(n51560), .B(n51439), .Z(n51440) );
  IV U64323 ( .A(n51440), .Z(n51557) );
  NOR U64324 ( .A(n51441), .B(n51557), .Z(n51553) );
  IV U64325 ( .A(n51442), .Z(n51558) );
  IV U64326 ( .A(n51443), .Z(n51446) );
  IV U64327 ( .A(n51444), .Z(n51445) );
  NOR U64328 ( .A(n51446), .B(n51445), .Z(n51447) );
  IV U64329 ( .A(n51447), .Z(n51556) );
  XOR U64330 ( .A(n51558), .B(n51556), .Z(n51448) );
  XOR U64331 ( .A(n51557), .B(n51448), .Z(n51547) );
  IV U64332 ( .A(n51547), .Z(n51449) );
  NOR U64333 ( .A(n51450), .B(n51449), .Z(n51451) );
  NOR U64334 ( .A(n51553), .B(n51451), .Z(n51472) );
  IV U64335 ( .A(n51472), .Z(n51550) );
  IV U64336 ( .A(n51452), .Z(n51453) );
  NOR U64337 ( .A(n51454), .B(n51453), .Z(n51471) );
  IV U64338 ( .A(n51455), .Z(n51457) );
  NOR U64339 ( .A(n51457), .B(n51456), .Z(n51546) );
  NOR U64340 ( .A(n51471), .B(n51546), .Z(n51458) );
  XOR U64341 ( .A(n51550), .B(n51458), .Z(n51475) );
  IV U64342 ( .A(n51475), .Z(n51463) );
  IV U64343 ( .A(n51459), .Z(n51461) );
  NOR U64344 ( .A(n51461), .B(n51460), .Z(n51480) );
  IV U64345 ( .A(n51480), .Z(n51462) );
  NOR U64346 ( .A(n51463), .B(n51462), .Z(n55137) );
  IV U64347 ( .A(n51464), .Z(n51465) );
  NOR U64348 ( .A(n51466), .B(n51465), .Z(n51467) );
  IV U64349 ( .A(n51467), .Z(n51543) );
  IV U64350 ( .A(n51468), .Z(n51469) );
  NOR U64351 ( .A(n51470), .B(n51469), .Z(n51476) );
  IV U64352 ( .A(n51476), .Z(n51474) );
  IV U64353 ( .A(n51471), .Z(n51551) );
  XOR U64354 ( .A(n51551), .B(n51472), .Z(n51473) );
  NOR U64355 ( .A(n51474), .B(n51473), .Z(n51545) );
  NOR U64356 ( .A(n51476), .B(n51475), .Z(n51477) );
  NOR U64357 ( .A(n51545), .B(n51477), .Z(n51478) );
  IV U64358 ( .A(n51478), .Z(n51542) );
  XOR U64359 ( .A(n51543), .B(n51542), .Z(n51479) );
  NOR U64360 ( .A(n51480), .B(n51479), .Z(n51481) );
  NOR U64361 ( .A(n55137), .B(n51481), .Z(n54872) );
  XOR U64362 ( .A(n54874), .B(n54872), .Z(n54885) );
  XOR U64363 ( .A(n51482), .B(n54885), .Z(n51483) );
  IV U64364 ( .A(n51483), .Z(n54877) );
  XOR U64365 ( .A(n54876), .B(n54877), .Z(n51537) );
  IV U64366 ( .A(n51484), .Z(n51486) );
  NOR U64367 ( .A(n51486), .B(n51485), .Z(n51535) );
  XOR U64368 ( .A(n51537), .B(n51535), .Z(n54892) );
  XOR U64369 ( .A(n51538), .B(n54892), .Z(n51531) );
  IV U64370 ( .A(n51531), .Z(n51493) );
  IV U64371 ( .A(n51487), .Z(n54893) );
  NOR U64372 ( .A(n54893), .B(n51488), .Z(n51491) );
  NOR U64373 ( .A(n51489), .B(n51532), .Z(n51490) );
  NOR U64374 ( .A(n51491), .B(n51490), .Z(n51492) );
  XOR U64375 ( .A(n51493), .B(n51492), .Z(n51529) );
  IV U64376 ( .A(n51494), .Z(n51495) );
  NOR U64377 ( .A(n51495), .B(n51532), .Z(n51527) );
  XOR U64378 ( .A(n51529), .B(n51527), .Z(n54903) );
  XOR U64379 ( .A(n54902), .B(n54903), .Z(n54907) );
  XOR U64380 ( .A(n54905), .B(n54907), .Z(n51525) );
  XOR U64381 ( .A(n51524), .B(n51525), .Z(n51523) );
  IV U64382 ( .A(n51496), .Z(n51497) );
  NOR U64383 ( .A(n51506), .B(n51497), .Z(n51512) );
  IV U64384 ( .A(n51512), .Z(n51498) );
  NOR U64385 ( .A(n51523), .B(n51498), .Z(n51499) );
  NOR U64386 ( .A(n51514), .B(n51499), .Z(n51520) );
  IV U64387 ( .A(n51520), .Z(n51513) );
  IV U64388 ( .A(n51500), .Z(n51502) );
  NOR U64389 ( .A(n51502), .B(n51501), .Z(n51503) );
  IV U64390 ( .A(n51503), .Z(n51507) );
  NOR U64391 ( .A(n51507), .B(n51525), .Z(n55094) );
  IV U64392 ( .A(n51504), .Z(n51505) );
  NOR U64393 ( .A(n51506), .B(n51505), .Z(n51508) );
  IV U64394 ( .A(n51508), .Z(n51522) );
  XOR U64395 ( .A(n51523), .B(n51522), .Z(n51510) );
  NOR U64396 ( .A(n51508), .B(n51507), .Z(n51509) );
  NOR U64397 ( .A(n51510), .B(n51509), .Z(n51511) );
  NOR U64398 ( .A(n55094), .B(n51511), .Z(n51516) );
  NOR U64399 ( .A(n51516), .B(n51512), .Z(n51521) );
  NOR U64400 ( .A(n51513), .B(n51521), .Z(n51518) );
  IV U64401 ( .A(n51514), .Z(n51515) );
  NOR U64402 ( .A(n51516), .B(n51515), .Z(n51517) );
  NOR U64403 ( .A(n51518), .B(n51517), .Z(n54911) );
  NOR U64404 ( .A(n54912), .B(n54911), .Z(n51519) );
  IV U64405 ( .A(n51519), .Z(n55046) );
  NOR U64406 ( .A(n51521), .B(n51520), .Z(n58668) );
  NOR U64407 ( .A(n51523), .B(n51522), .Z(n58665) );
  IV U64408 ( .A(n51524), .Z(n51526) );
  NOR U64409 ( .A(n51526), .B(n51525), .Z(n58675) );
  IV U64410 ( .A(n51527), .Z(n51528) );
  NOR U64411 ( .A(n51529), .B(n51528), .Z(n55116) );
  IV U64412 ( .A(n51530), .Z(n51534) );
  NOR U64413 ( .A(n51532), .B(n51531), .Z(n51533) );
  IV U64414 ( .A(n51533), .Z(n54900) );
  NOR U64415 ( .A(n51534), .B(n54900), .Z(n55124) );
  IV U64416 ( .A(n51535), .Z(n51536) );
  NOR U64417 ( .A(n51537), .B(n51536), .Z(n51541) );
  IV U64418 ( .A(n51538), .Z(n51539) );
  NOR U64419 ( .A(n51539), .B(n54892), .Z(n51540) );
  NOR U64420 ( .A(n51541), .B(n51540), .Z(n58651) );
  NOR U64421 ( .A(n51543), .B(n51542), .Z(n51544) );
  NOR U64422 ( .A(n51545), .B(n51544), .Z(n58638) );
  IV U64423 ( .A(n51546), .Z(n51548) );
  NOR U64424 ( .A(n51548), .B(n51547), .Z(n51549) );
  IV U64425 ( .A(n51549), .Z(n58636) );
  NOR U64426 ( .A(n51551), .B(n51550), .Z(n51552) );
  NOR U64427 ( .A(n51553), .B(n51552), .Z(n55144) );
  IV U64428 ( .A(n51554), .Z(n51555) );
  NOR U64429 ( .A(n51556), .B(n51555), .Z(n55140) );
  NOR U64430 ( .A(n51558), .B(n51557), .Z(n51559) );
  NOR U64431 ( .A(n51560), .B(n51559), .Z(n55151) );
  IV U64432 ( .A(n51561), .Z(n51562) );
  NOR U64433 ( .A(n54863), .B(n51562), .Z(n55147) );
  IV U64434 ( .A(n51563), .Z(n51564) );
  NOR U64435 ( .A(n54860), .B(n51564), .Z(n55156) );
  IV U64436 ( .A(n51565), .Z(n51566) );
  NOR U64437 ( .A(n51566), .B(n51568), .Z(n58583) );
  IV U64438 ( .A(n51567), .Z(n51569) );
  NOR U64439 ( .A(n51569), .B(n51568), .Z(n58580) );
  IV U64440 ( .A(n51570), .Z(n51571) );
  NOR U64441 ( .A(n51572), .B(n51571), .Z(n51577) );
  IV U64442 ( .A(n51573), .Z(n51574) );
  NOR U64443 ( .A(n51575), .B(n51574), .Z(n51576) );
  NOR U64444 ( .A(n51577), .B(n51576), .Z(n58579) );
  IV U64445 ( .A(n51578), .Z(n51579) );
  NOR U64446 ( .A(n51580), .B(n51579), .Z(n51584) );
  IV U64447 ( .A(n51581), .Z(n51582) );
  NOR U64448 ( .A(n51582), .B(n51590), .Z(n51583) );
  NOR U64449 ( .A(n51584), .B(n51583), .Z(n58618) );
  IV U64450 ( .A(n51585), .Z(n51587) );
  NOR U64451 ( .A(n51587), .B(n51586), .Z(n58620) );
  IV U64452 ( .A(n51588), .Z(n51589) );
  NOR U64453 ( .A(n51590), .B(n51589), .Z(n58591) );
  NOR U64454 ( .A(n58620), .B(n58591), .Z(n54858) );
  IV U64455 ( .A(n51591), .Z(n51596) );
  IV U64456 ( .A(n51592), .Z(n51593) );
  NOR U64457 ( .A(n51593), .B(n51603), .Z(n51594) );
  IV U64458 ( .A(n51594), .Z(n51595) );
  NOR U64459 ( .A(n51596), .B(n51595), .Z(n58599) );
  IV U64460 ( .A(n51597), .Z(n51601) );
  NOR U64461 ( .A(n51598), .B(n51609), .Z(n51599) );
  IV U64462 ( .A(n51599), .Z(n51600) );
  NOR U64463 ( .A(n51601), .B(n51600), .Z(n58596) );
  IV U64464 ( .A(n51602), .Z(n51604) );
  NOR U64465 ( .A(n51604), .B(n51603), .Z(n58607) );
  IV U64466 ( .A(n51605), .Z(n51606) );
  NOR U64467 ( .A(n51607), .B(n51606), .Z(n51612) );
  IV U64468 ( .A(n51608), .Z(n51610) );
  NOR U64469 ( .A(n51610), .B(n51609), .Z(n51611) );
  NOR U64470 ( .A(n51612), .B(n51611), .Z(n58605) );
  IV U64471 ( .A(n51613), .Z(n51614) );
  NOR U64472 ( .A(n51615), .B(n51614), .Z(n58550) );
  IV U64473 ( .A(n51616), .Z(n51620) );
  IV U64474 ( .A(n51617), .Z(n54847) );
  NOR U64475 ( .A(n51618), .B(n54847), .Z(n51619) );
  IV U64476 ( .A(n51619), .Z(n51622) );
  NOR U64477 ( .A(n51620), .B(n51622), .Z(n58539) );
  NOR U64478 ( .A(n58550), .B(n58539), .Z(n54856) );
  IV U64479 ( .A(n51621), .Z(n51623) );
  NOR U64480 ( .A(n51623), .B(n51622), .Z(n58541) );
  IV U64481 ( .A(n58541), .Z(n58538) );
  IV U64482 ( .A(n51624), .Z(n58527) );
  IV U64483 ( .A(n51625), .Z(n58529) );
  IV U64484 ( .A(n51626), .Z(n51627) );
  NOR U64485 ( .A(n51628), .B(n51627), .Z(n54833) );
  IV U64486 ( .A(n51629), .Z(n51630) );
  NOR U64487 ( .A(n51631), .B(n51630), .Z(n51632) );
  IV U64488 ( .A(n51632), .Z(n58520) );
  IV U64489 ( .A(n51633), .Z(n51634) );
  NOR U64490 ( .A(n51635), .B(n51634), .Z(n51640) );
  IV U64491 ( .A(n51636), .Z(n51637) );
  NOR U64492 ( .A(n51638), .B(n51637), .Z(n51639) );
  NOR U64493 ( .A(n51640), .B(n51639), .Z(n58518) );
  NOR U64494 ( .A(n51642), .B(n51641), .Z(n51643) );
  NOR U64495 ( .A(n51644), .B(n51643), .Z(n55184) );
  IV U64496 ( .A(n51645), .Z(n51647) );
  NOR U64497 ( .A(n51647), .B(n51646), .Z(n55180) );
  IV U64498 ( .A(n51648), .Z(n51651) );
  IV U64499 ( .A(n51649), .Z(n51660) );
  XOR U64500 ( .A(n51653), .B(n51660), .Z(n51650) );
  NOR U64501 ( .A(n51651), .B(n51650), .Z(n58479) );
  IV U64502 ( .A(n51652), .Z(n51656) );
  IV U64503 ( .A(n51653), .Z(n51661) );
  NOR U64504 ( .A(n51661), .B(n51654), .Z(n51655) );
  IV U64505 ( .A(n51655), .Z(n51658) );
  NOR U64506 ( .A(n51656), .B(n51658), .Z(n58476) );
  IV U64507 ( .A(n51657), .Z(n51659) );
  NOR U64508 ( .A(n51659), .B(n51658), .Z(n58493) );
  NOR U64509 ( .A(n51661), .B(n51660), .Z(n58499) );
  IV U64510 ( .A(n51662), .Z(n51663) );
  NOR U64511 ( .A(n51664), .B(n51663), .Z(n58496) );
  NOR U64512 ( .A(n51666), .B(n51665), .Z(n51672) );
  IV U64513 ( .A(n51667), .Z(n51670) );
  IV U64514 ( .A(n51668), .Z(n51669) );
  NOR U64515 ( .A(n51670), .B(n51669), .Z(n51671) );
  NOR U64516 ( .A(n51672), .B(n51671), .Z(n58485) );
  NOR U64517 ( .A(n51674), .B(n51673), .Z(n51677) );
  IV U64518 ( .A(n51675), .Z(n51676) );
  NOR U64519 ( .A(n51677), .B(n51676), .Z(n55242) );
  IV U64520 ( .A(n51678), .Z(n51679) );
  NOR U64521 ( .A(n51682), .B(n51679), .Z(n55239) );
  IV U64522 ( .A(n51680), .Z(n51681) );
  NOR U64523 ( .A(n51682), .B(n51681), .Z(n58459) );
  NOR U64524 ( .A(n51683), .B(n51685), .Z(n58456) );
  IV U64525 ( .A(n51684), .Z(n51686) );
  NOR U64526 ( .A(n51686), .B(n51685), .Z(n58467) );
  IV U64527 ( .A(n51687), .Z(n51689) );
  IV U64528 ( .A(n51688), .Z(n51691) );
  NOR U64529 ( .A(n51689), .B(n51691), .Z(n58464) );
  NOR U64530 ( .A(n51691), .B(n51690), .Z(n55230) );
  NOR U64531 ( .A(n51693), .B(n51692), .Z(n55227) );
  IV U64532 ( .A(n51694), .Z(n51695) );
  NOR U64533 ( .A(n51696), .B(n51695), .Z(n54784) );
  IV U64534 ( .A(n54784), .Z(n54782) );
  NOR U64535 ( .A(n51698), .B(n51697), .Z(n51699) );
  NOR U64536 ( .A(n51702), .B(n51699), .Z(n55207) );
  IV U64537 ( .A(n51700), .Z(n51701) );
  NOR U64538 ( .A(n51702), .B(n51701), .Z(n55192) );
  IV U64539 ( .A(n51703), .Z(n51705) );
  NOR U64540 ( .A(n51705), .B(n51704), .Z(n55189) );
  IV U64541 ( .A(n51706), .Z(n51707) );
  NOR U64542 ( .A(n51710), .B(n51707), .Z(n55200) );
  IV U64543 ( .A(n51708), .Z(n51709) );
  NOR U64544 ( .A(n51710), .B(n51709), .Z(n55258) );
  IV U64545 ( .A(n51711), .Z(n51712) );
  NOR U64546 ( .A(n51713), .B(n51712), .Z(n55255) );
  IV U64547 ( .A(n51714), .Z(n51715) );
  NOR U64548 ( .A(n51716), .B(n51715), .Z(n55266) );
  IV U64549 ( .A(n51717), .Z(n51720) );
  IV U64550 ( .A(n51718), .Z(n51725) );
  XOR U64551 ( .A(n51725), .B(n51722), .Z(n51719) );
  NOR U64552 ( .A(n51720), .B(n51719), .Z(n55263) );
  IV U64553 ( .A(n51721), .Z(n51723) );
  IV U64554 ( .A(n51722), .Z(n51724) );
  NOR U64555 ( .A(n51723), .B(n51724), .Z(n55274) );
  NOR U64556 ( .A(n51725), .B(n51724), .Z(n55271) );
  IV U64557 ( .A(n51726), .Z(n51727) );
  NOR U64558 ( .A(n54761), .B(n51727), .Z(n55251) );
  NOR U64559 ( .A(n55271), .B(n55251), .Z(n54762) );
  IV U64560 ( .A(n51728), .Z(n51729) );
  NOR U64561 ( .A(n51729), .B(n51733), .Z(n54752) );
  IV U64562 ( .A(n54752), .Z(n54750) );
  IV U64563 ( .A(n51730), .Z(n51731) );
  NOR U64564 ( .A(n51732), .B(n51731), .Z(n51736) );
  NOR U64565 ( .A(n51734), .B(n51733), .Z(n51735) );
  NOR U64566 ( .A(n51736), .B(n51735), .Z(n55285) );
  IV U64567 ( .A(n51737), .Z(n54748) );
  IV U64568 ( .A(n51738), .Z(n51739) );
  NOR U64569 ( .A(n54748), .B(n51739), .Z(n55281) );
  IV U64570 ( .A(n51740), .Z(n51742) );
  NOR U64571 ( .A(n51742), .B(n51741), .Z(n55370) );
  NOR U64572 ( .A(n51743), .B(n51744), .Z(n51750) );
  IV U64573 ( .A(n51744), .Z(n51745) );
  NOR U64574 ( .A(n51746), .B(n51745), .Z(n51748) );
  NOR U64575 ( .A(n51748), .B(n51747), .Z(n51749) );
  NOR U64576 ( .A(n51750), .B(n51749), .Z(n55358) );
  NOR U64577 ( .A(n51752), .B(n51751), .Z(n55361) );
  IV U64578 ( .A(n51753), .Z(n51755) );
  NOR U64579 ( .A(n51755), .B(n51754), .Z(n55332) );
  NOR U64580 ( .A(n55361), .B(n55332), .Z(n54744) );
  NOR U64581 ( .A(n51757), .B(n51756), .Z(n51763) );
  NOR U64582 ( .A(n51759), .B(n51758), .Z(n51761) );
  NOR U64583 ( .A(n51761), .B(n51760), .Z(n51762) );
  NOR U64584 ( .A(n51763), .B(n51762), .Z(n55333) );
  IV U64585 ( .A(n55333), .Z(n55339) );
  IV U64586 ( .A(n51764), .Z(n51766) );
  NOR U64587 ( .A(n51766), .B(n51765), .Z(n51771) );
  IV U64588 ( .A(n51767), .Z(n51768) );
  NOR U64589 ( .A(n51769), .B(n51768), .Z(n51770) );
  NOR U64590 ( .A(n51771), .B(n51770), .Z(n55337) );
  NOR U64591 ( .A(n51773), .B(n51772), .Z(n54734) );
  IV U64592 ( .A(n51774), .Z(n51775) );
  NOR U64593 ( .A(n51776), .B(n51775), .Z(n51778) );
  NOR U64594 ( .A(n51778), .B(n51777), .Z(n55307) );
  IV U64595 ( .A(n51779), .Z(n51782) );
  IV U64596 ( .A(n51780), .Z(n51781) );
  NOR U64597 ( .A(n51782), .B(n51781), .Z(n55311) );
  IV U64598 ( .A(n51783), .Z(n51784) );
  NOR U64599 ( .A(n51784), .B(n51785), .Z(n55308) );
  NOR U64600 ( .A(n51786), .B(n51785), .Z(n55321) );
  IV U64601 ( .A(n51787), .Z(n54722) );
  IV U64602 ( .A(n51788), .Z(n51789) );
  NOR U64603 ( .A(n54722), .B(n51789), .Z(n55301) );
  IV U64604 ( .A(n51790), .Z(n51791) );
  NOR U64605 ( .A(n51791), .B(n54709), .Z(n51792) );
  IV U64606 ( .A(n51792), .Z(n55399) );
  IV U64607 ( .A(n51793), .Z(n51794) );
  NOR U64608 ( .A(n51794), .B(n54695), .Z(n58422) );
  IV U64609 ( .A(n51795), .Z(n51796) );
  NOR U64610 ( .A(n51797), .B(n51796), .Z(n55433) );
  IV U64611 ( .A(n51798), .Z(n51801) );
  NOR U64612 ( .A(n51799), .B(n51810), .Z(n51800) );
  IV U64613 ( .A(n51800), .Z(n51803) );
  NOR U64614 ( .A(n51801), .B(n51803), .Z(n55429) );
  IV U64615 ( .A(n51802), .Z(n51804) );
  NOR U64616 ( .A(n51804), .B(n51803), .Z(n58410) );
  IV U64617 ( .A(n51805), .Z(n51806) );
  NOR U64618 ( .A(n51807), .B(n51806), .Z(n55424) );
  IV U64619 ( .A(n51808), .Z(n51809) );
  NOR U64620 ( .A(n51810), .B(n51809), .Z(n58407) );
  NOR U64621 ( .A(n55424), .B(n58407), .Z(n54686) );
  IV U64622 ( .A(n51811), .Z(n51812) );
  NOR U64623 ( .A(n51813), .B(n51812), .Z(n55423) );
  NOR U64624 ( .A(n51815), .B(n51814), .Z(n51821) );
  IV U64625 ( .A(n51815), .Z(n51817) );
  NOR U64626 ( .A(n51817), .B(n51816), .Z(n51818) );
  NOR U64627 ( .A(n51819), .B(n51818), .Z(n51820) );
  NOR U64628 ( .A(n51821), .B(n51820), .Z(n55408) );
  IV U64629 ( .A(n51822), .Z(n51823) );
  NOR U64630 ( .A(n51823), .B(n51826), .Z(n55405) );
  IV U64631 ( .A(n51824), .Z(n51825) );
  NOR U64632 ( .A(n51826), .B(n51825), .Z(n55416) );
  IV U64633 ( .A(n51827), .Z(n51829) );
  IV U64634 ( .A(n51828), .Z(n51831) );
  NOR U64635 ( .A(n51829), .B(n51831), .Z(n54670) );
  IV U64636 ( .A(n51830), .Z(n51834) );
  NOR U64637 ( .A(n51832), .B(n51831), .Z(n51833) );
  IV U64638 ( .A(n51833), .Z(n55451) );
  NOR U64639 ( .A(n51834), .B(n55451), .Z(n54661) );
  IV U64640 ( .A(n51835), .Z(n51840) );
  IV U64641 ( .A(n51836), .Z(n51837) );
  NOR U64642 ( .A(n51840), .B(n51837), .Z(n54645) );
  IV U64643 ( .A(n54645), .Z(n54643) );
  IV U64644 ( .A(n51838), .Z(n51839) );
  NOR U64645 ( .A(n51840), .B(n51839), .Z(n51841) );
  IV U64646 ( .A(n51841), .Z(n55461) );
  IV U64647 ( .A(n51842), .Z(n51843) );
  NOR U64648 ( .A(n51846), .B(n51843), .Z(n55457) );
  IV U64649 ( .A(n51844), .Z(n51845) );
  NOR U64650 ( .A(n51846), .B(n51845), .Z(n51847) );
  IV U64651 ( .A(n51847), .Z(n55498) );
  IV U64652 ( .A(n51848), .Z(n51849) );
  NOR U64653 ( .A(n51850), .B(n51849), .Z(n51855) );
  IV U64654 ( .A(n51851), .Z(n51852) );
  NOR U64655 ( .A(n51853), .B(n51852), .Z(n51854) );
  NOR U64656 ( .A(n51855), .B(n51854), .Z(n55495) );
  NOR U64657 ( .A(n51856), .B(n54640), .Z(n55501) );
  IV U64658 ( .A(n51857), .Z(n51860) );
  NOR U64659 ( .A(n51858), .B(n54640), .Z(n51859) );
  IV U64660 ( .A(n51859), .Z(n51862) );
  NOR U64661 ( .A(n51860), .B(n51862), .Z(n55469) );
  IV U64662 ( .A(n51861), .Z(n51863) );
  NOR U64663 ( .A(n51863), .B(n51862), .Z(n55466) );
  IV U64664 ( .A(n51864), .Z(n51865) );
  NOR U64665 ( .A(n51865), .B(n51869), .Z(n58348) );
  IV U64666 ( .A(n51866), .Z(n51867) );
  NOR U64667 ( .A(n51869), .B(n51867), .Z(n58354) );
  IV U64668 ( .A(n51868), .Z(n51870) );
  NOR U64669 ( .A(n51870), .B(n51869), .Z(n58351) );
  IV U64670 ( .A(n51876), .Z(n54597) );
  IV U64671 ( .A(n51871), .Z(n51872) );
  NOR U64672 ( .A(n54597), .B(n51872), .Z(n58343) );
  NOR U64673 ( .A(n51874), .B(n51873), .Z(n51875) );
  IV U64674 ( .A(n51875), .Z(n51877) );
  NOR U64675 ( .A(n51877), .B(n51876), .Z(n58344) );
  NOR U64676 ( .A(n58343), .B(n58344), .Z(n54594) );
  IV U64677 ( .A(n51878), .Z(n51882) );
  XOR U64678 ( .A(n51893), .B(n51894), .Z(n51879) );
  NOR U64679 ( .A(n51880), .B(n51879), .Z(n51881) );
  IV U64680 ( .A(n51881), .Z(n51884) );
  NOR U64681 ( .A(n51882), .B(n51884), .Z(n58325) );
  IV U64682 ( .A(n51883), .Z(n51885) );
  NOR U64683 ( .A(n51885), .B(n51884), .Z(n58331) );
  IV U64684 ( .A(n51886), .Z(n51889) );
  NOR U64685 ( .A(n51887), .B(n51894), .Z(n51888) );
  IV U64686 ( .A(n51888), .Z(n51891) );
  NOR U64687 ( .A(n51889), .B(n51891), .Z(n55516) );
  IV U64688 ( .A(n51890), .Z(n51892) );
  NOR U64689 ( .A(n51892), .B(n51891), .Z(n55513) );
  IV U64690 ( .A(n51893), .Z(n51895) );
  NOR U64691 ( .A(n51895), .B(n51894), .Z(n51896) );
  IV U64692 ( .A(n51896), .Z(n58330) );
  IV U64693 ( .A(n51897), .Z(n51899) );
  NOR U64694 ( .A(n51899), .B(n51898), .Z(n51904) );
  IV U64695 ( .A(n51900), .Z(n51902) );
  NOR U64696 ( .A(n51902), .B(n51901), .Z(n51903) );
  NOR U64697 ( .A(n51904), .B(n51903), .Z(n58308) );
  NOR U64698 ( .A(n51906), .B(n51905), .Z(n58304) );
  IV U64699 ( .A(n51907), .Z(n51910) );
  NOR U64700 ( .A(n51908), .B(n51919), .Z(n51909) );
  IV U64701 ( .A(n51909), .Z(n51912) );
  NOR U64702 ( .A(n51910), .B(n51912), .Z(n58311) );
  IV U64703 ( .A(n51911), .Z(n51913) );
  NOR U64704 ( .A(n51913), .B(n51912), .Z(n58289) );
  IV U64705 ( .A(n51914), .Z(n51916) );
  NOR U64706 ( .A(n51916), .B(n51915), .Z(n51921) );
  IV U64707 ( .A(n51917), .Z(n51918) );
  NOR U64708 ( .A(n51919), .B(n51918), .Z(n51920) );
  NOR U64709 ( .A(n51921), .B(n51920), .Z(n51922) );
  IV U64710 ( .A(n51922), .Z(n58273) );
  IV U64711 ( .A(n51923), .Z(n51924) );
  NOR U64712 ( .A(n51925), .B(n51924), .Z(n58292) );
  NOR U64713 ( .A(n58273), .B(n58292), .Z(n54593) );
  IV U64714 ( .A(n51926), .Z(n51928) );
  NOR U64715 ( .A(n51928), .B(n51927), .Z(n54584) );
  IV U64716 ( .A(n51929), .Z(n51931) );
  NOR U64717 ( .A(n51931), .B(n51930), .Z(n54587) );
  IV U64718 ( .A(n51932), .Z(n51935) );
  IV U64719 ( .A(n51933), .Z(n54565) );
  XOR U64720 ( .A(n54565), .B(n51936), .Z(n51934) );
  NOR U64721 ( .A(n51935), .B(n51934), .Z(n58277) );
  IV U64722 ( .A(n51936), .Z(n54576) );
  IV U64723 ( .A(n51937), .Z(n54563) );
  IV U64724 ( .A(n51938), .Z(n51939) );
  NOR U64725 ( .A(n51939), .B(n51941), .Z(n55560) );
  IV U64726 ( .A(n51940), .Z(n51942) );
  NOR U64727 ( .A(n51942), .B(n51941), .Z(n55557) );
  IV U64728 ( .A(n51943), .Z(n51945) );
  IV U64729 ( .A(n51944), .Z(n54552) );
  NOR U64730 ( .A(n51945), .B(n54552), .Z(n55565) );
  NOR U64731 ( .A(n55521), .B(n55565), .Z(n54547) );
  IV U64732 ( .A(n51946), .Z(n51947) );
  NOR U64733 ( .A(n51954), .B(n51947), .Z(n51951) );
  NOR U64734 ( .A(n51949), .B(n51948), .Z(n51950) );
  NOR U64735 ( .A(n51951), .B(n51950), .Z(n55532) );
  IV U64736 ( .A(n51952), .Z(n51953) );
  NOR U64737 ( .A(n51954), .B(n51953), .Z(n51959) );
  IV U64738 ( .A(n51955), .Z(n51957) );
  NOR U64739 ( .A(n51957), .B(n51956), .Z(n51958) );
  NOR U64740 ( .A(n51959), .B(n51958), .Z(n55529) );
  IV U64741 ( .A(n51960), .Z(n51962) );
  NOR U64742 ( .A(n51962), .B(n51961), .Z(n55535) );
  IV U64743 ( .A(n51963), .Z(n51966) );
  NOR U64744 ( .A(n51964), .B(n51972), .Z(n51965) );
  IV U64745 ( .A(n51965), .Z(n51968) );
  NOR U64746 ( .A(n51966), .B(n51968), .Z(n55603) );
  IV U64747 ( .A(n51967), .Z(n51969) );
  NOR U64748 ( .A(n51969), .B(n51968), .Z(n55614) );
  IV U64749 ( .A(n51970), .Z(n51971) );
  NOR U64750 ( .A(n51972), .B(n51971), .Z(n55577) );
  IV U64751 ( .A(n51973), .Z(n51974) );
  NOR U64752 ( .A(n51975), .B(n51974), .Z(n55574) );
  IV U64753 ( .A(n51980), .Z(n51977) );
  NOR U64754 ( .A(n51977), .B(n51976), .Z(n51984) );
  IV U64755 ( .A(n51978), .Z(n51982) );
  NOR U64756 ( .A(n51980), .B(n51979), .Z(n51981) );
  NOR U64757 ( .A(n51982), .B(n51981), .Z(n51983) );
  NOR U64758 ( .A(n51984), .B(n51983), .Z(n55588) );
  IV U64759 ( .A(n51985), .Z(n51986) );
  NOR U64760 ( .A(n51989), .B(n51986), .Z(n55584) );
  IV U64761 ( .A(n51987), .Z(n51988) );
  NOR U64762 ( .A(n51989), .B(n51988), .Z(n55611) );
  IV U64763 ( .A(n51990), .Z(n51991) );
  NOR U64764 ( .A(n51992), .B(n51991), .Z(n55594) );
  IV U64765 ( .A(n51993), .Z(n51994) );
  NOR U64766 ( .A(n51994), .B(n52000), .Z(n51995) );
  IV U64767 ( .A(n51995), .Z(n55592) );
  IV U64768 ( .A(n51996), .Z(n51997) );
  NOR U64769 ( .A(n52005), .B(n51997), .Z(n52002) );
  IV U64770 ( .A(n51998), .Z(n51999) );
  NOR U64771 ( .A(n52000), .B(n51999), .Z(n52001) );
  NOR U64772 ( .A(n52002), .B(n52001), .Z(n55583) );
  IV U64773 ( .A(n52003), .Z(n52004) );
  NOR U64774 ( .A(n52005), .B(n52004), .Z(n58239) );
  IV U64775 ( .A(n52006), .Z(n52011) );
  IV U64776 ( .A(n52007), .Z(n52008) );
  NOR U64777 ( .A(n52015), .B(n52008), .Z(n52009) );
  IV U64778 ( .A(n52009), .Z(n52010) );
  NOR U64779 ( .A(n52011), .B(n52010), .Z(n58245) );
  NOR U64780 ( .A(n52013), .B(n52012), .Z(n52014) );
  IV U64781 ( .A(n52014), .Z(n52016) );
  NOR U64782 ( .A(n52016), .B(n52015), .Z(n58242) );
  IV U64783 ( .A(n52017), .Z(n54526) );
  IV U64784 ( .A(n52018), .Z(n52019) );
  NOR U64785 ( .A(n54526), .B(n52019), .Z(n58255) );
  IV U64786 ( .A(n52020), .Z(n52021) );
  NOR U64787 ( .A(n52021), .B(n54522), .Z(n55626) );
  IV U64788 ( .A(n52022), .Z(n52023) );
  NOR U64789 ( .A(n52024), .B(n52023), .Z(n55623) );
  NOR U64790 ( .A(n55677), .B(n55623), .Z(n54519) );
  IV U64791 ( .A(n55672), .Z(n55675) );
  IV U64792 ( .A(n52025), .Z(n52026) );
  NOR U64793 ( .A(n52027), .B(n52026), .Z(n52028) );
  IV U64794 ( .A(n52028), .Z(n55664) );
  IV U64795 ( .A(n52029), .Z(n52030) );
  NOR U64796 ( .A(n52031), .B(n52030), .Z(n52036) );
  IV U64797 ( .A(n52032), .Z(n52033) );
  NOR U64798 ( .A(n52034), .B(n52033), .Z(n52035) );
  NOR U64799 ( .A(n52036), .B(n52035), .Z(n55657) );
  IV U64800 ( .A(n55657), .Z(n52040) );
  IV U64801 ( .A(n52037), .Z(n52038) );
  NOR U64802 ( .A(n52039), .B(n52038), .Z(n55665) );
  NOR U64803 ( .A(n52040), .B(n55665), .Z(n54518) );
  IV U64804 ( .A(n52041), .Z(n52043) );
  NOR U64805 ( .A(n52043), .B(n52042), .Z(n55658) );
  IV U64806 ( .A(n52044), .Z(n52046) );
  NOR U64807 ( .A(n52046), .B(n52045), .Z(n58210) );
  NOR U64808 ( .A(n55658), .B(n58210), .Z(n54517) );
  IV U64809 ( .A(n52047), .Z(n52048) );
  NOR U64810 ( .A(n52048), .B(n52050), .Z(n52055) );
  IV U64811 ( .A(n52049), .Z(n52053) );
  NOR U64812 ( .A(n52051), .B(n52050), .Z(n52052) );
  IV U64813 ( .A(n52052), .Z(n52057) );
  NOR U64814 ( .A(n52053), .B(n52057), .Z(n52054) );
  NOR U64815 ( .A(n52055), .B(n52054), .Z(n58211) );
  IV U64816 ( .A(n52056), .Z(n52058) );
  NOR U64817 ( .A(n52058), .B(n52057), .Z(n58207) );
  XOR U64818 ( .A(n52060), .B(n52059), .Z(n52061) );
  NOR U64819 ( .A(n55639), .B(n52061), .Z(n52062) );
  NOR U64820 ( .A(n52063), .B(n52062), .Z(n54515) );
  IV U64821 ( .A(n52064), .Z(n52068) );
  NOR U64822 ( .A(n52066), .B(n52065), .Z(n52067) );
  IV U64823 ( .A(n52067), .Z(n52071) );
  NOR U64824 ( .A(n52068), .B(n52071), .Z(n52069) );
  NOR U64825 ( .A(n55646), .B(n52069), .Z(n55649) );
  IV U64826 ( .A(n52070), .Z(n52072) );
  NOR U64827 ( .A(n52072), .B(n52071), .Z(n55651) );
  IV U64828 ( .A(n52073), .Z(n52075) );
  NOR U64829 ( .A(n52075), .B(n52074), .Z(n58226) );
  IV U64830 ( .A(n52076), .Z(n52079) );
  NOR U64831 ( .A(n52077), .B(n52090), .Z(n52078) );
  IV U64832 ( .A(n52078), .Z(n52081) );
  NOR U64833 ( .A(n52079), .B(n52081), .Z(n58144) );
  IV U64834 ( .A(n52080), .Z(n52082) );
  NOR U64835 ( .A(n52082), .B(n52081), .Z(n58141) );
  IV U64836 ( .A(n52083), .Z(n52085) );
  NOR U64837 ( .A(n52085), .B(n52084), .Z(n58191) );
  IV U64838 ( .A(n52086), .Z(n52088) );
  NOR U64839 ( .A(n52088), .B(n52087), .Z(n55686) );
  IV U64840 ( .A(n52089), .Z(n52091) );
  NOR U64841 ( .A(n52091), .B(n52090), .Z(n58138) );
  NOR U64842 ( .A(n55686), .B(n58138), .Z(n54484) );
  IV U64843 ( .A(n52092), .Z(n52095) );
  NOR U64844 ( .A(n52102), .B(n52097), .Z(n52093) );
  IV U64845 ( .A(n52093), .Z(n52094) );
  NOR U64846 ( .A(n52095), .B(n52094), .Z(n55684) );
  IV U64847 ( .A(n55684), .Z(n55682) );
  IV U64848 ( .A(n52098), .Z(n52096) );
  NOR U64849 ( .A(n52097), .B(n52096), .Z(n52107) );
  NOR U64850 ( .A(n52099), .B(n52098), .Z(n52105) );
  IV U64851 ( .A(n52100), .Z(n52101) );
  NOR U64852 ( .A(n52102), .B(n52101), .Z(n52103) );
  IV U64853 ( .A(n52103), .Z(n52104) );
  NOR U64854 ( .A(n52105), .B(n52104), .Z(n52106) );
  NOR U64855 ( .A(n52107), .B(n52106), .Z(n58176) );
  IV U64856 ( .A(n52113), .Z(n52109) );
  NOR U64857 ( .A(n52109), .B(n52108), .Z(n55728) );
  NOR U64858 ( .A(n52111), .B(n52110), .Z(n58178) );
  NOR U64859 ( .A(n55728), .B(n58178), .Z(n54482) );
  IV U64860 ( .A(n52112), .Z(n52114) );
  NOR U64861 ( .A(n52114), .B(n52113), .Z(n55727) );
  IV U64862 ( .A(n52115), .Z(n52116) );
  NOR U64863 ( .A(n52117), .B(n52116), .Z(n52118) );
  NOR U64864 ( .A(n52119), .B(n52118), .Z(n58155) );
  NOR U64865 ( .A(n52121), .B(n52120), .Z(n52122) );
  IV U64866 ( .A(n52122), .Z(n55713) );
  IV U64867 ( .A(n52123), .Z(n52125) );
  NOR U64868 ( .A(n52125), .B(n52124), .Z(n54459) );
  IV U64869 ( .A(n54459), .Z(n54450) );
  IV U64870 ( .A(n52126), .Z(n52127) );
  NOR U64871 ( .A(n52128), .B(n52127), .Z(n52129) );
  IV U64872 ( .A(n52129), .Z(n52130) );
  NOR U64873 ( .A(n52131), .B(n52130), .Z(n55696) );
  NOR U64874 ( .A(n52133), .B(n52132), .Z(n52134) );
  NOR U64875 ( .A(n52135), .B(n52134), .Z(n55707) );
  IV U64876 ( .A(n52136), .Z(n52137) );
  NOR U64877 ( .A(n52138), .B(n52137), .Z(n55705) );
  IV U64878 ( .A(n52139), .Z(n52142) );
  NOR U64879 ( .A(n52140), .B(n52145), .Z(n52141) );
  IV U64880 ( .A(n52141), .Z(n52147) );
  NOR U64881 ( .A(n52142), .B(n52147), .Z(n55774) );
  NOR U64882 ( .A(n55705), .B(n55774), .Z(n54449) );
  IV U64883 ( .A(n52143), .Z(n52144) );
  NOR U64884 ( .A(n52145), .B(n52144), .Z(n55767) );
  IV U64885 ( .A(n52146), .Z(n52148) );
  NOR U64886 ( .A(n52148), .B(n52147), .Z(n55777) );
  NOR U64887 ( .A(n55767), .B(n55777), .Z(n54448) );
  IV U64888 ( .A(n52149), .Z(n52150) );
  NOR U64889 ( .A(n52151), .B(n52150), .Z(n52156) );
  IV U64890 ( .A(n52152), .Z(n52154) );
  NOR U64891 ( .A(n52154), .B(n52153), .Z(n52155) );
  NOR U64892 ( .A(n52156), .B(n52155), .Z(n55766) );
  IV U64893 ( .A(n52157), .Z(n52158) );
  NOR U64894 ( .A(n52159), .B(n52158), .Z(n55768) );
  IV U64895 ( .A(n52160), .Z(n52161) );
  NOR U64896 ( .A(n52161), .B(n54445), .Z(n54441) );
  IV U64897 ( .A(n54441), .Z(n54429) );
  IV U64898 ( .A(n54434), .Z(n54432) );
  NOR U64899 ( .A(n54432), .B(n54435), .Z(n55748) );
  IV U64900 ( .A(n52162), .Z(n52163) );
  NOR U64901 ( .A(n52163), .B(n52167), .Z(n55750) );
  IV U64902 ( .A(n52164), .Z(n52165) );
  NOR U64903 ( .A(n52165), .B(n52167), .Z(n55734) );
  IV U64904 ( .A(n52166), .Z(n52168) );
  NOR U64905 ( .A(n52168), .B(n52167), .Z(n55731) );
  NOR U64906 ( .A(n52170), .B(n52169), .Z(n52171) );
  IV U64907 ( .A(n52171), .Z(n52172) );
  NOR U64908 ( .A(n52172), .B(n52182), .Z(n55739) );
  IV U64909 ( .A(n52173), .Z(n52178) );
  IV U64910 ( .A(n52174), .Z(n52175) );
  NOR U64911 ( .A(n52178), .B(n52175), .Z(n58115) );
  IV U64912 ( .A(n52176), .Z(n52177) );
  NOR U64913 ( .A(n52178), .B(n52177), .Z(n58113) );
  NOR U64914 ( .A(n58115), .B(n58113), .Z(n52179) );
  IV U64915 ( .A(n52179), .Z(n52183) );
  IV U64916 ( .A(n52180), .Z(n52181) );
  NOR U64917 ( .A(n52182), .B(n52181), .Z(n58112) );
  NOR U64918 ( .A(n52183), .B(n58112), .Z(n54416) );
  IV U64919 ( .A(n52184), .Z(n52185) );
  NOR U64920 ( .A(n52186), .B(n52185), .Z(n58108) );
  IV U64921 ( .A(n58108), .Z(n58110) );
  IV U64922 ( .A(n52187), .Z(n52191) );
  IV U64923 ( .A(n52188), .Z(n54408) );
  NOR U64924 ( .A(n52189), .B(n54408), .Z(n52190) );
  IV U64925 ( .A(n52190), .Z(n54413) );
  NOR U64926 ( .A(n52191), .B(n54413), .Z(n52192) );
  IV U64927 ( .A(n52192), .Z(n58125) );
  IV U64928 ( .A(n52193), .Z(n52194) );
  NOR U64929 ( .A(n52197), .B(n52194), .Z(n54407) );
  IV U64930 ( .A(n54407), .Z(n54405) );
  IV U64931 ( .A(n52195), .Z(n52196) );
  NOR U64932 ( .A(n52197), .B(n52196), .Z(n52198) );
  IV U64933 ( .A(n52198), .Z(n58090) );
  IV U64934 ( .A(n52199), .Z(n52202) );
  IV U64935 ( .A(n52200), .Z(n52201) );
  NOR U64936 ( .A(n52202), .B(n52201), .Z(n58094) );
  NOR U64937 ( .A(n52204), .B(n52203), .Z(n52205) );
  NOR U64938 ( .A(n52206), .B(n52205), .Z(n58091) );
  NOR U64939 ( .A(n52208), .B(n52207), .Z(n55801) );
  IV U64940 ( .A(n52209), .Z(n52210) );
  NOR U64941 ( .A(n52210), .B(n52213), .Z(n55798) );
  IV U64942 ( .A(n52213), .Z(n52211) );
  NOR U64943 ( .A(n52212), .B(n52211), .Z(n52218) );
  NOR U64944 ( .A(n52214), .B(n52213), .Z(n52215) );
  NOR U64945 ( .A(n52216), .B(n52215), .Z(n52217) );
  NOR U64946 ( .A(n52218), .B(n52217), .Z(n52219) );
  IV U64947 ( .A(n52219), .Z(n55852) );
  IV U64948 ( .A(n52220), .Z(n52222) );
  NOR U64949 ( .A(n52222), .B(n52221), .Z(n52227) );
  IV U64950 ( .A(n52223), .Z(n52225) );
  NOR U64951 ( .A(n52225), .B(n52224), .Z(n52226) );
  NOR U64952 ( .A(n52227), .B(n52226), .Z(n55837) );
  NOR U64953 ( .A(n52228), .B(n55830), .Z(n55838) );
  IV U64954 ( .A(n52229), .Z(n52230) );
  NOR U64955 ( .A(n52231), .B(n52230), .Z(n52236) );
  IV U64956 ( .A(n52232), .Z(n52233) );
  NOR U64957 ( .A(n52234), .B(n52233), .Z(n52235) );
  NOR U64958 ( .A(n52236), .B(n52235), .Z(n55825) );
  NOR U64959 ( .A(n52238), .B(n52237), .Z(n55809) );
  IV U64960 ( .A(n55809), .Z(n52239) );
  NOR U64961 ( .A(n52239), .B(n55806), .Z(n52240) );
  IV U64962 ( .A(n52240), .Z(n52241) );
  NOR U64963 ( .A(n55808), .B(n52241), .Z(n52242) );
  NOR U64964 ( .A(n52243), .B(n52242), .Z(n54403) );
  NOR U64965 ( .A(n52245), .B(n52244), .Z(n54396) );
  IV U64966 ( .A(n52246), .Z(n52251) );
  IV U64967 ( .A(n52247), .Z(n52248) );
  NOR U64968 ( .A(n52251), .B(n52248), .Z(n54393) );
  IV U64969 ( .A(n52249), .Z(n52250) );
  NOR U64970 ( .A(n52251), .B(n52250), .Z(n55819) );
  IV U64971 ( .A(n52252), .Z(n52253) );
  NOR U64972 ( .A(n52253), .B(n52256), .Z(n55817) );
  IV U64973 ( .A(n52254), .Z(n52255) );
  NOR U64974 ( .A(n52256), .B(n52255), .Z(n55814) );
  NOR U64975 ( .A(n55817), .B(n55814), .Z(n54390) );
  IV U64976 ( .A(n52257), .Z(n52259) );
  NOR U64977 ( .A(n52259), .B(n52258), .Z(n52264) );
  IV U64978 ( .A(n52260), .Z(n52262) );
  NOR U64979 ( .A(n52262), .B(n52261), .Z(n52263) );
  NOR U64980 ( .A(n52264), .B(n52263), .Z(n58063) );
  IV U64981 ( .A(n52265), .Z(n52266) );
  NOR U64982 ( .A(n52266), .B(n52272), .Z(n55854) );
  IV U64983 ( .A(n52267), .Z(n52279) );
  IV U64984 ( .A(n52268), .Z(n52269) );
  NOR U64985 ( .A(n52279), .B(n52269), .Z(n58069) );
  XOR U64986 ( .A(n52271), .B(n52270), .Z(n52273) );
  NOR U64987 ( .A(n52273), .B(n52272), .Z(n52274) );
  IV U64988 ( .A(n52274), .Z(n52275) );
  NOR U64989 ( .A(n52276), .B(n52275), .Z(n55858) );
  NOR U64990 ( .A(n58069), .B(n55858), .Z(n54389) );
  IV U64991 ( .A(n52277), .Z(n52278) );
  NOR U64992 ( .A(n52279), .B(n52278), .Z(n58068) );
  IV U64993 ( .A(n52280), .Z(n52281) );
  NOR U64994 ( .A(n52281), .B(n54385), .Z(n58043) );
  NOR U64995 ( .A(n58068), .B(n58043), .Z(n54388) );
  NOR U64996 ( .A(n52283), .B(n52282), .Z(n54379) );
  IV U64997 ( .A(n54379), .Z(n54369) );
  IV U64998 ( .A(n52284), .Z(n52286) );
  NOR U64999 ( .A(n52286), .B(n52285), .Z(n58017) );
  IV U65000 ( .A(n52287), .Z(n52289) );
  NOR U65001 ( .A(n52289), .B(n52288), .Z(n52294) );
  IV U65002 ( .A(n52290), .Z(n52292) );
  NOR U65003 ( .A(n52292), .B(n52291), .Z(n52293) );
  NOR U65004 ( .A(n52294), .B(n52293), .Z(n58035) );
  IV U65005 ( .A(n52295), .Z(n52296) );
  NOR U65006 ( .A(n52297), .B(n52296), .Z(n58001) );
  IV U65007 ( .A(n52298), .Z(n52300) );
  NOR U65008 ( .A(n52300), .B(n52299), .Z(n52304) );
  NOR U65009 ( .A(n52302), .B(n52301), .Z(n52303) );
  NOR U65010 ( .A(n52304), .B(n52303), .Z(n58010) );
  IV U65011 ( .A(n52305), .Z(n52306) );
  NOR U65012 ( .A(n52307), .B(n52306), .Z(n52312) );
  IV U65013 ( .A(n52308), .Z(n52310) );
  NOR U65014 ( .A(n52310), .B(n52309), .Z(n52311) );
  NOR U65015 ( .A(n52312), .B(n52311), .Z(n58008) );
  IV U65016 ( .A(n52313), .Z(n52314) );
  NOR U65017 ( .A(n52315), .B(n52314), .Z(n52320) );
  IV U65018 ( .A(n52316), .Z(n52317) );
  NOR U65019 ( .A(n52318), .B(n52317), .Z(n52319) );
  NOR U65020 ( .A(n52320), .B(n52319), .Z(n58023) );
  IV U65021 ( .A(n52321), .Z(n52323) );
  NOR U65022 ( .A(n52323), .B(n52322), .Z(n58020) );
  IV U65023 ( .A(n52324), .Z(n52326) );
  NOR U65024 ( .A(n52326), .B(n52325), .Z(n52327) );
  IV U65025 ( .A(n52327), .Z(n52328) );
  NOR U65026 ( .A(n52329), .B(n52328), .Z(n55877) );
  IV U65027 ( .A(n58026), .Z(n58024) );
  IV U65028 ( .A(n52330), .Z(n58028) );
  NOR U65029 ( .A(n58024), .B(n58028), .Z(n54331) );
  IV U65030 ( .A(n52331), .Z(n52332) );
  NOR U65031 ( .A(n54315), .B(n52332), .Z(n54317) );
  IV U65032 ( .A(n52333), .Z(n52334) );
  NOR U65033 ( .A(n52334), .B(n54307), .Z(n54320) );
  NOR U65034 ( .A(n52336), .B(n52335), .Z(n57976) );
  IV U65035 ( .A(n52337), .Z(n52338) );
  NOR U65036 ( .A(n52338), .B(n52342), .Z(n52340) );
  NOR U65037 ( .A(n52340), .B(n52339), .Z(n57961) );
  IV U65038 ( .A(n52341), .Z(n52343) );
  NOR U65039 ( .A(n52343), .B(n52342), .Z(n55892) );
  IV U65040 ( .A(n52344), .Z(n52345) );
  NOR U65041 ( .A(n52345), .B(n54301), .Z(n57965) );
  NOR U65042 ( .A(n52347), .B(n52346), .Z(n57962) );
  IV U65043 ( .A(n52348), .Z(n52349) );
  NOR U65044 ( .A(n52350), .B(n52349), .Z(n57949) );
  IV U65045 ( .A(n52351), .Z(n52352) );
  NOR U65046 ( .A(n52353), .B(n52352), .Z(n57936) );
  NOR U65047 ( .A(n54285), .B(n52354), .Z(n52355) );
  IV U65048 ( .A(n52355), .Z(n55917) );
  IV U65049 ( .A(n52356), .Z(n52357) );
  NOR U65050 ( .A(n52357), .B(n52359), .Z(n55900) );
  IV U65051 ( .A(n52358), .Z(n52360) );
  NOR U65052 ( .A(n52360), .B(n52359), .Z(n55897) );
  IV U65053 ( .A(n52361), .Z(n52363) );
  IV U65054 ( .A(n52362), .Z(n54279) );
  NOR U65055 ( .A(n52363), .B(n54279), .Z(n55905) );
  IV U65056 ( .A(n52364), .Z(n52365) );
  NOR U65057 ( .A(n52365), .B(n54279), .Z(n55941) );
  IV U65058 ( .A(n52366), .Z(n52368) );
  NOR U65059 ( .A(n52368), .B(n52367), .Z(n54239) );
  IV U65060 ( .A(n52369), .Z(n52371) );
  NOR U65061 ( .A(n52371), .B(n52370), .Z(n55918) );
  IV U65062 ( .A(n52372), .Z(n52377) );
  IV U65063 ( .A(n52378), .Z(n54213) );
  IV U65064 ( .A(n52373), .Z(n52374) );
  NOR U65065 ( .A(n54213), .B(n52374), .Z(n52375) );
  IV U65066 ( .A(n52375), .Z(n52376) );
  NOR U65067 ( .A(n52377), .B(n52376), .Z(n55929) );
  NOR U65068 ( .A(n52379), .B(n52378), .Z(n52390) );
  NOR U65069 ( .A(n54213), .B(n52380), .Z(n52388) );
  IV U65070 ( .A(n52381), .Z(n52382) );
  NOR U65071 ( .A(n52383), .B(n52382), .Z(n52384) );
  IV U65072 ( .A(n52384), .Z(n52385) );
  NOR U65073 ( .A(n52386), .B(n52385), .Z(n52387) );
  NOR U65074 ( .A(n52388), .B(n52387), .Z(n52389) );
  NOR U65075 ( .A(n52390), .B(n52389), .Z(n55958) );
  IV U65076 ( .A(n52391), .Z(n52393) );
  NOR U65077 ( .A(n52393), .B(n52392), .Z(n57897) );
  IV U65078 ( .A(n52397), .Z(n52394) );
  NOR U65079 ( .A(n52394), .B(n52395), .Z(n52405) );
  IV U65080 ( .A(n52395), .Z(n52396) );
  NOR U65081 ( .A(n52397), .B(n52396), .Z(n52403) );
  IV U65082 ( .A(n52398), .Z(n52400) );
  NOR U65083 ( .A(n52400), .B(n52399), .Z(n52401) );
  IV U65084 ( .A(n52401), .Z(n52402) );
  NOR U65085 ( .A(n52403), .B(n52402), .Z(n52404) );
  NOR U65086 ( .A(n52405), .B(n52404), .Z(n57903) );
  IV U65087 ( .A(n52406), .Z(n52407) );
  NOR U65088 ( .A(n52407), .B(n54194), .Z(n57884) );
  IV U65089 ( .A(n52408), .Z(n52410) );
  NOR U65090 ( .A(n52410), .B(n52409), .Z(n54188) );
  IV U65091 ( .A(n54188), .Z(n54186) );
  IV U65092 ( .A(n52411), .Z(n55997) );
  NOR U65093 ( .A(n52413), .B(n52412), .Z(n55965) );
  IV U65094 ( .A(n52414), .Z(n52417) );
  IV U65095 ( .A(n52415), .Z(n52416) );
  NOR U65096 ( .A(n52417), .B(n52416), .Z(n55993) );
  NOR U65097 ( .A(n55965), .B(n55993), .Z(n54180) );
  NOR U65098 ( .A(n52419), .B(n52418), .Z(n52420) );
  NOR U65099 ( .A(n52421), .B(n52420), .Z(n55986) );
  IV U65100 ( .A(n55975), .Z(n55972) );
  IV U65101 ( .A(n52422), .Z(n52426) );
  NOR U65102 ( .A(n54170), .B(n52423), .Z(n52424) );
  IV U65103 ( .A(n52424), .Z(n52425) );
  NOR U65104 ( .A(n52426), .B(n52425), .Z(n57865) );
  IV U65105 ( .A(n52427), .Z(n52429) );
  NOR U65106 ( .A(n52429), .B(n52428), .Z(n52434) );
  IV U65107 ( .A(n52430), .Z(n52431) );
  NOR U65108 ( .A(n52432), .B(n52431), .Z(n52433) );
  NOR U65109 ( .A(n52434), .B(n52433), .Z(n57856) );
  IV U65110 ( .A(n52435), .Z(n52436) );
  NOR U65111 ( .A(n52437), .B(n52436), .Z(n52442) );
  IV U65112 ( .A(n52438), .Z(n52440) );
  NOR U65113 ( .A(n52440), .B(n52439), .Z(n52441) );
  NOR U65114 ( .A(n52442), .B(n52441), .Z(n56019) );
  IV U65115 ( .A(n52443), .Z(n52446) );
  IV U65116 ( .A(n52444), .Z(n52445) );
  NOR U65117 ( .A(n52446), .B(n52445), .Z(n56010) );
  IV U65118 ( .A(n52447), .Z(n52448) );
  NOR U65119 ( .A(n52448), .B(n52450), .Z(n56020) );
  IV U65120 ( .A(n52449), .Z(n52451) );
  NOR U65121 ( .A(n52451), .B(n52450), .Z(n56037) );
  IV U65122 ( .A(n52452), .Z(n52454) );
  NOR U65123 ( .A(n52454), .B(n52453), .Z(n52455) );
  NOR U65124 ( .A(n52456), .B(n52455), .Z(n56032) );
  IV U65125 ( .A(n52457), .Z(n52459) );
  NOR U65126 ( .A(n52459), .B(n52458), .Z(n56058) );
  NOR U65127 ( .A(n54141), .B(n52460), .Z(n56066) );
  IV U65128 ( .A(n52464), .Z(n52462) );
  NOR U65129 ( .A(n52462), .B(n52461), .Z(n52469) );
  NOR U65130 ( .A(n52464), .B(n52463), .Z(n52467) );
  IV U65131 ( .A(n52465), .Z(n52466) );
  NOR U65132 ( .A(n52467), .B(n52466), .Z(n52468) );
  NOR U65133 ( .A(n52469), .B(n52468), .Z(n56044) );
  NOR U65134 ( .A(n52471), .B(n52470), .Z(n52478) );
  IV U65135 ( .A(n52472), .Z(n52476) );
  NOR U65136 ( .A(n52474), .B(n52473), .Z(n52475) );
  IV U65137 ( .A(n52475), .Z(n52482) );
  NOR U65138 ( .A(n52476), .B(n52482), .Z(n52477) );
  NOR U65139 ( .A(n52478), .B(n52477), .Z(n56051) );
  IV U65140 ( .A(n52479), .Z(n52480) );
  NOR U65141 ( .A(n52480), .B(n52482), .Z(n56047) );
  IV U65142 ( .A(n52481), .Z(n52485) );
  NOR U65143 ( .A(n52483), .B(n52482), .Z(n52484) );
  IV U65144 ( .A(n52484), .Z(n52487) );
  NOR U65145 ( .A(n52485), .B(n52487), .Z(n56081) );
  IV U65146 ( .A(n52486), .Z(n52488) );
  NOR U65147 ( .A(n52488), .B(n52487), .Z(n56078) );
  IV U65148 ( .A(n52489), .Z(n52494) );
  IV U65149 ( .A(n52490), .Z(n52491) );
  NOR U65150 ( .A(n52492), .B(n52491), .Z(n52493) );
  IV U65151 ( .A(n52493), .Z(n52496) );
  NOR U65152 ( .A(n52494), .B(n52496), .Z(n56089) );
  IV U65153 ( .A(n52495), .Z(n52497) );
  NOR U65154 ( .A(n52497), .B(n52496), .Z(n56086) );
  IV U65155 ( .A(n52498), .Z(n52500) );
  NOR U65156 ( .A(n52500), .B(n52499), .Z(n54130) );
  IV U65157 ( .A(n52501), .Z(n52503) );
  NOR U65158 ( .A(n52503), .B(n52502), .Z(n57796) );
  IV U65159 ( .A(n52504), .Z(n52506) );
  NOR U65160 ( .A(n52506), .B(n52505), .Z(n57809) );
  NOR U65161 ( .A(n57796), .B(n57809), .Z(n54117) );
  IV U65162 ( .A(n52507), .Z(n52509) );
  NOR U65163 ( .A(n52509), .B(n52508), .Z(n54083) );
  IV U65164 ( .A(n52510), .Z(n54078) );
  NOR U65165 ( .A(n52511), .B(n54078), .Z(n54074) );
  IV U65166 ( .A(n54074), .Z(n54070) );
  IV U65167 ( .A(n52512), .Z(n52514) );
  NOR U65168 ( .A(n52514), .B(n52513), .Z(n52515) );
  NOR U65169 ( .A(n52516), .B(n52515), .Z(n57745) );
  IV U65170 ( .A(n52517), .Z(n52519) );
  NOR U65171 ( .A(n52519), .B(n52518), .Z(n54064) );
  IV U65172 ( .A(n54064), .Z(n54058) );
  IV U65173 ( .A(n52520), .Z(n52521) );
  NOR U65174 ( .A(n52522), .B(n52521), .Z(n57759) );
  IV U65175 ( .A(n52523), .Z(n52524) );
  NOR U65176 ( .A(n52524), .B(n52526), .Z(n57763) );
  IV U65177 ( .A(n52525), .Z(n52527) );
  NOR U65178 ( .A(n52527), .B(n52526), .Z(n57756) );
  IV U65179 ( .A(n52528), .Z(n54055) );
  IV U65180 ( .A(n52529), .Z(n52530) );
  NOR U65181 ( .A(n54055), .B(n52530), .Z(n57751) );
  IV U65182 ( .A(n52531), .Z(n52532) );
  NOR U65183 ( .A(n54055), .B(n52532), .Z(n52533) );
  IV U65184 ( .A(n52533), .Z(n57750) );
  IV U65185 ( .A(n52534), .Z(n52536) );
  NOR U65186 ( .A(n52536), .B(n52535), .Z(n54052) );
  IV U65187 ( .A(n54052), .Z(n54050) );
  NOR U65188 ( .A(n52538), .B(n52537), .Z(n52544) );
  IV U65189 ( .A(n52538), .Z(n52540) );
  NOR U65190 ( .A(n52540), .B(n52539), .Z(n52541) );
  NOR U65191 ( .A(n52542), .B(n52541), .Z(n52543) );
  NOR U65192 ( .A(n52544), .B(n52543), .Z(n52545) );
  IV U65193 ( .A(n52545), .Z(n56121) );
  NOR U65194 ( .A(n52547), .B(n52546), .Z(n56124) );
  IV U65195 ( .A(n52548), .Z(n52550) );
  NOR U65196 ( .A(n52550), .B(n52549), .Z(n56118) );
  IV U65197 ( .A(n52551), .Z(n52552) );
  NOR U65198 ( .A(n52555), .B(n52552), .Z(n56107) );
  IV U65199 ( .A(n52553), .Z(n52554) );
  NOR U65200 ( .A(n52555), .B(n52554), .Z(n56113) );
  IV U65201 ( .A(n52556), .Z(n52559) );
  IV U65202 ( .A(n52557), .Z(n52558) );
  NOR U65203 ( .A(n52559), .B(n52558), .Z(n52560) );
  IV U65204 ( .A(n52560), .Z(n56112) );
  IV U65205 ( .A(n52561), .Z(n52562) );
  NOR U65206 ( .A(n52563), .B(n52562), .Z(n52564) );
  NOR U65207 ( .A(n56137), .B(n52564), .Z(n57723) );
  IV U65208 ( .A(n52565), .Z(n52567) );
  NOR U65209 ( .A(n52567), .B(n52566), .Z(n52572) );
  IV U65210 ( .A(n52568), .Z(n52570) );
  NOR U65211 ( .A(n52570), .B(n52569), .Z(n52571) );
  NOR U65212 ( .A(n52572), .B(n52571), .Z(n52573) );
  IV U65213 ( .A(n52573), .Z(n57700) );
  NOR U65214 ( .A(n57700), .B(n57719), .Z(n54048) );
  IV U65215 ( .A(n52574), .Z(n52576) );
  NOR U65216 ( .A(n52576), .B(n52575), .Z(n54044) );
  IV U65217 ( .A(n52577), .Z(n52579) );
  NOR U65218 ( .A(n52579), .B(n52578), .Z(n54041) );
  IV U65219 ( .A(n54041), .Z(n54036) );
  NOR U65220 ( .A(n52581), .B(n52580), .Z(n52589) );
  IV U65221 ( .A(n52582), .Z(n52587) );
  IV U65222 ( .A(n52583), .Z(n52584) );
  NOR U65223 ( .A(n52585), .B(n52584), .Z(n52586) );
  IV U65224 ( .A(n52586), .Z(n52591) );
  NOR U65225 ( .A(n52587), .B(n52591), .Z(n52588) );
  NOR U65226 ( .A(n52589), .B(n52588), .Z(n56144) );
  IV U65227 ( .A(n52590), .Z(n52592) );
  NOR U65228 ( .A(n52592), .B(n52591), .Z(n56140) );
  IV U65229 ( .A(n52593), .Z(n52595) );
  NOR U65230 ( .A(n52595), .B(n52594), .Z(n52596) );
  NOR U65231 ( .A(n52597), .B(n52596), .Z(n57690) );
  IV U65232 ( .A(n52598), .Z(n52599) );
  NOR U65233 ( .A(n52599), .B(n52601), .Z(n57677) );
  IV U65234 ( .A(n57677), .Z(n57674) );
  IV U65235 ( .A(n52600), .Z(n52602) );
  NOR U65236 ( .A(n52602), .B(n52601), .Z(n52603) );
  IV U65237 ( .A(n52603), .Z(n57665) );
  NOR U65238 ( .A(n52604), .B(n54011), .Z(n57661) );
  IV U65239 ( .A(n52605), .Z(n52607) );
  NOR U65240 ( .A(n52607), .B(n52606), .Z(n56154) );
  IV U65241 ( .A(n52608), .Z(n52612) );
  NOR U65242 ( .A(n52609), .B(n53999), .Z(n52610) );
  IV U65243 ( .A(n52610), .Z(n52611) );
  NOR U65244 ( .A(n52612), .B(n52611), .Z(n57637) );
  IV U65245 ( .A(n57637), .Z(n57632) );
  IV U65246 ( .A(n52613), .Z(n53996) );
  IV U65247 ( .A(n52614), .Z(n52615) );
  NOR U65248 ( .A(n53996), .B(n52615), .Z(n57647) );
  IV U65249 ( .A(n52616), .Z(n52618) );
  NOR U65250 ( .A(n52618), .B(n52617), .Z(n56182) );
  IV U65251 ( .A(n52619), .Z(n52621) );
  NOR U65252 ( .A(n52621), .B(n52620), .Z(n52626) );
  IV U65253 ( .A(n52622), .Z(n52624) );
  NOR U65254 ( .A(n52624), .B(n52623), .Z(n52625) );
  NOR U65255 ( .A(n52626), .B(n52625), .Z(n56173) );
  IV U65256 ( .A(n52630), .Z(n52628) );
  IV U65257 ( .A(n52629), .Z(n52627) );
  NOR U65258 ( .A(n52628), .B(n52627), .Z(n52635) );
  NOR U65259 ( .A(n52630), .B(n52629), .Z(n52633) );
  IV U65260 ( .A(n52631), .Z(n52632) );
  NOR U65261 ( .A(n52633), .B(n52632), .Z(n52634) );
  NOR U65262 ( .A(n52635), .B(n52634), .Z(n56189) );
  NOR U65263 ( .A(n52637), .B(n52636), .Z(n52642) );
  IV U65264 ( .A(n52638), .Z(n52639) );
  NOR U65265 ( .A(n52640), .B(n52639), .Z(n52641) );
  NOR U65266 ( .A(n52642), .B(n52641), .Z(n56194) );
  IV U65267 ( .A(n52643), .Z(n52645) );
  NOR U65268 ( .A(n52645), .B(n52644), .Z(n52650) );
  IV U65269 ( .A(n52646), .Z(n52647) );
  NOR U65270 ( .A(n52648), .B(n52647), .Z(n52649) );
  NOR U65271 ( .A(n52650), .B(n52649), .Z(n56198) );
  IV U65272 ( .A(n52651), .Z(n52653) );
  NOR U65273 ( .A(n52653), .B(n52652), .Z(n52658) );
  IV U65274 ( .A(n52654), .Z(n52655) );
  NOR U65275 ( .A(n52656), .B(n52655), .Z(n52657) );
  NOR U65276 ( .A(n52658), .B(n52657), .Z(n57580) );
  IV U65277 ( .A(n52659), .Z(n52660) );
  NOR U65278 ( .A(n52661), .B(n52660), .Z(n56210) );
  IV U65279 ( .A(n52662), .Z(n52665) );
  IV U65280 ( .A(n52663), .Z(n52664) );
  NOR U65281 ( .A(n52665), .B(n52664), .Z(n56207) );
  IV U65282 ( .A(n52666), .Z(n52667) );
  NOR U65283 ( .A(n52667), .B(n53953), .Z(n57589) );
  IV U65284 ( .A(n52668), .Z(n52669) );
  NOR U65285 ( .A(n52669), .B(n53940), .Z(n53943) );
  IV U65286 ( .A(n52670), .Z(n52671) );
  NOR U65287 ( .A(n52671), .B(n53927), .Z(n57552) );
  IV U65288 ( .A(n52672), .Z(n52674) );
  NOR U65289 ( .A(n52674), .B(n52673), .Z(n57549) );
  IV U65290 ( .A(n52675), .Z(n52678) );
  NOR U65291 ( .A(n52676), .B(n52687), .Z(n52677) );
  IV U65292 ( .A(n52677), .Z(n52680) );
  NOR U65293 ( .A(n52678), .B(n52680), .Z(n57557) );
  IV U65294 ( .A(n52679), .Z(n52681) );
  NOR U65295 ( .A(n52681), .B(n52680), .Z(n56251) );
  IV U65296 ( .A(n52682), .Z(n52683) );
  NOR U65297 ( .A(n52684), .B(n52683), .Z(n56254) );
  IV U65298 ( .A(n52685), .Z(n52686) );
  NOR U65299 ( .A(n52687), .B(n52686), .Z(n56248) );
  NOR U65300 ( .A(n56254), .B(n56248), .Z(n53918) );
  IV U65301 ( .A(n52688), .Z(n52693) );
  IV U65302 ( .A(n52689), .Z(n52690) );
  NOR U65303 ( .A(n52693), .B(n52690), .Z(n56243) );
  IV U65304 ( .A(n56243), .Z(n56245) );
  IV U65305 ( .A(n52691), .Z(n52692) );
  NOR U65306 ( .A(n52693), .B(n52692), .Z(n52694) );
  IV U65307 ( .A(n52694), .Z(n56239) );
  IV U65308 ( .A(n52700), .Z(n52699) );
  IV U65309 ( .A(n52695), .Z(n52696) );
  NOR U65310 ( .A(n52699), .B(n52696), .Z(n52697) );
  IV U65311 ( .A(n52697), .Z(n56238) );
  NOR U65312 ( .A(n52699), .B(n52698), .Z(n52706) );
  NOR U65313 ( .A(n52701), .B(n52700), .Z(n52704) );
  IV U65314 ( .A(n52702), .Z(n52703) );
  NOR U65315 ( .A(n52704), .B(n52703), .Z(n52705) );
  NOR U65316 ( .A(n52706), .B(n52705), .Z(n56265) );
  IV U65317 ( .A(n52707), .Z(n52709) );
  NOR U65318 ( .A(n52709), .B(n52708), .Z(n52710) );
  NOR U65319 ( .A(n52711), .B(n52710), .Z(n56277) );
  NOR U65320 ( .A(n52713), .B(n52712), .Z(n56271) );
  IV U65321 ( .A(n52714), .Z(n52715) );
  NOR U65322 ( .A(n53899), .B(n52715), .Z(n56268) );
  IV U65323 ( .A(n52716), .Z(n52719) );
  IV U65324 ( .A(n52717), .Z(n52718) );
  NOR U65325 ( .A(n52719), .B(n52718), .Z(n56280) );
  IV U65326 ( .A(n52720), .Z(n52721) );
  NOR U65327 ( .A(n52722), .B(n52721), .Z(n56301) );
  IV U65328 ( .A(n52723), .Z(n52727) );
  NOR U65329 ( .A(n52725), .B(n52724), .Z(n52726) );
  IV U65330 ( .A(n52726), .Z(n52729) );
  NOR U65331 ( .A(n52727), .B(n52729), .Z(n56304) );
  IV U65332 ( .A(n52728), .Z(n52730) );
  NOR U65333 ( .A(n52730), .B(n52729), .Z(n56285) );
  IV U65334 ( .A(n52731), .Z(n52732) );
  NOR U65335 ( .A(n52732), .B(n53895), .Z(n56291) );
  IV U65336 ( .A(n52733), .Z(n52734) );
  NOR U65337 ( .A(n52734), .B(n53895), .Z(n56288) );
  IV U65338 ( .A(n57530), .Z(n57525) );
  NOR U65339 ( .A(n52736), .B(n52735), .Z(n52737) );
  NOR U65340 ( .A(n52738), .B(n52737), .Z(n56318) );
  IV U65341 ( .A(n52739), .Z(n52740) );
  NOR U65342 ( .A(n52740), .B(n53888), .Z(n56324) );
  IV U65343 ( .A(n52741), .Z(n56343) );
  IV U65344 ( .A(n52742), .Z(n52743) );
  NOR U65345 ( .A(n52747), .B(n52743), .Z(n56341) );
  IV U65346 ( .A(n56341), .Z(n56339) );
  XOR U65347 ( .A(n56343), .B(n56339), .Z(n52744) );
  NOR U65348 ( .A(n56324), .B(n52744), .Z(n53885) );
  IV U65349 ( .A(n52745), .Z(n52746) );
  NOR U65350 ( .A(n52747), .B(n52746), .Z(n56321) );
  IV U65351 ( .A(n52748), .Z(n52750) );
  NOR U65352 ( .A(n52750), .B(n52749), .Z(n56328) );
  NOR U65353 ( .A(n52752), .B(n52751), .Z(n52754) );
  NOR U65354 ( .A(n52754), .B(n52753), .Z(n56331) );
  NOR U65355 ( .A(n52756), .B(n52755), .Z(n53882) );
  IV U65356 ( .A(n53882), .Z(n53868) );
  IV U65357 ( .A(n52757), .Z(n52758) );
  NOR U65358 ( .A(n52758), .B(n53855), .Z(n53853) );
  IV U65359 ( .A(n53853), .Z(n53851) );
  IV U65360 ( .A(n52759), .Z(n52760) );
  NOR U65361 ( .A(n52761), .B(n52760), .Z(n52766) );
  IV U65362 ( .A(n52762), .Z(n52764) );
  NOR U65363 ( .A(n52764), .B(n52763), .Z(n52765) );
  NOR U65364 ( .A(n52766), .B(n52765), .Z(n56347) );
  IV U65365 ( .A(n52767), .Z(n52768) );
  NOR U65366 ( .A(n52768), .B(n52774), .Z(n56352) );
  IV U65367 ( .A(n52769), .Z(n52770) );
  NOR U65368 ( .A(n52771), .B(n52770), .Z(n56361) );
  IV U65369 ( .A(n52772), .Z(n52773) );
  NOR U65370 ( .A(n52774), .B(n52773), .Z(n56348) );
  NOR U65371 ( .A(n56361), .B(n56348), .Z(n53848) );
  IV U65372 ( .A(n52775), .Z(n52779) );
  IV U65373 ( .A(n52776), .Z(n52777) );
  NOR U65374 ( .A(n52779), .B(n52777), .Z(n56360) );
  IV U65375 ( .A(n52778), .Z(n52780) );
  NOR U65376 ( .A(n52780), .B(n52779), .Z(n52785) );
  IV U65377 ( .A(n52781), .Z(n52783) );
  NOR U65378 ( .A(n52783), .B(n52782), .Z(n52784) );
  NOR U65379 ( .A(n52785), .B(n52784), .Z(n56368) );
  IV U65380 ( .A(n52788), .Z(n52787) );
  NOR U65381 ( .A(n52787), .B(n52786), .Z(n52794) );
  NOR U65382 ( .A(n52789), .B(n52788), .Z(n52792) );
  IV U65383 ( .A(n52790), .Z(n52791) );
  NOR U65384 ( .A(n52792), .B(n52791), .Z(n52793) );
  NOR U65385 ( .A(n52794), .B(n52793), .Z(n56365) );
  IV U65386 ( .A(n52795), .Z(n52797) );
  NOR U65387 ( .A(n52797), .B(n52796), .Z(n56384) );
  IV U65388 ( .A(n56372), .Z(n56374) );
  IV U65389 ( .A(n52798), .Z(n52799) );
  NOR U65390 ( .A(n52800), .B(n52799), .Z(n56392) );
  IV U65391 ( .A(n52801), .Z(n52802) );
  NOR U65392 ( .A(n53833), .B(n52802), .Z(n56444) );
  IV U65393 ( .A(n52803), .Z(n52804) );
  NOR U65394 ( .A(n52805), .B(n52804), .Z(n56437) );
  IV U65395 ( .A(n52806), .Z(n52807) );
  NOR U65396 ( .A(n52807), .B(n53823), .Z(n52811) );
  NOR U65397 ( .A(n52809), .B(n52808), .Z(n52810) );
  NOR U65398 ( .A(n52811), .B(n52810), .Z(n56429) );
  IV U65399 ( .A(n56429), .Z(n56426) );
  IV U65400 ( .A(n52812), .Z(n52813) );
  NOR U65401 ( .A(n52813), .B(n52817), .Z(n56416) );
  IV U65402 ( .A(n52814), .Z(n52815) );
  NOR U65403 ( .A(n52815), .B(n52817), .Z(n56409) );
  IV U65404 ( .A(n52816), .Z(n52818) );
  NOR U65405 ( .A(n52818), .B(n52817), .Z(n53804) );
  IV U65406 ( .A(n52819), .Z(n52820) );
  NOR U65407 ( .A(n52821), .B(n52820), .Z(n52822) );
  IV U65408 ( .A(n52822), .Z(n53791) );
  IV U65409 ( .A(n52823), .Z(n52824) );
  NOR U65410 ( .A(n52825), .B(n52824), .Z(n52831) );
  IV U65411 ( .A(n52826), .Z(n52829) );
  IV U65412 ( .A(n52827), .Z(n52828) );
  NOR U65413 ( .A(n52829), .B(n52828), .Z(n52830) );
  NOR U65414 ( .A(n52831), .B(n52830), .Z(n57449) );
  NOR U65415 ( .A(n52833), .B(n52832), .Z(n53771) );
  IV U65416 ( .A(n52834), .Z(n56451) );
  IV U65417 ( .A(n52835), .Z(n52836) );
  NOR U65418 ( .A(n52837), .B(n52836), .Z(n56447) );
  IV U65419 ( .A(n52838), .Z(n52842) );
  IV U65420 ( .A(n52839), .Z(n52840) );
  NOR U65421 ( .A(n52842), .B(n52840), .Z(n57428) );
  IV U65422 ( .A(n52841), .Z(n52843) );
  NOR U65423 ( .A(n52843), .B(n52842), .Z(n57437) );
  IV U65424 ( .A(n52844), .Z(n52847) );
  NOR U65425 ( .A(n52845), .B(n53765), .Z(n52846) );
  IV U65426 ( .A(n52846), .Z(n52849) );
  NOR U65427 ( .A(n52847), .B(n52849), .Z(n57408) );
  IV U65428 ( .A(n52848), .Z(n52850) );
  NOR U65429 ( .A(n52850), .B(n52849), .Z(n52851) );
  IV U65430 ( .A(n52851), .Z(n57421) );
  NOR U65431 ( .A(n52853), .B(n52852), .Z(n57404) );
  NOR U65432 ( .A(n52855), .B(n52854), .Z(n52856) );
  NOR U65433 ( .A(n52857), .B(n52856), .Z(n56472) );
  IV U65434 ( .A(n52858), .Z(n52860) );
  NOR U65435 ( .A(n52860), .B(n52859), .Z(n56469) );
  IV U65436 ( .A(n52864), .Z(n52861) );
  NOR U65437 ( .A(n52862), .B(n52861), .Z(n52868) );
  IV U65438 ( .A(n52862), .Z(n52863) );
  NOR U65439 ( .A(n52864), .B(n52863), .Z(n52865) );
  NOR U65440 ( .A(n52866), .B(n52865), .Z(n52867) );
  NOR U65441 ( .A(n52868), .B(n52867), .Z(n56454) );
  NOR U65442 ( .A(n52870), .B(n52869), .Z(n57431) );
  IV U65443 ( .A(n52871), .Z(n52872) );
  NOR U65444 ( .A(n52873), .B(n52872), .Z(n57433) );
  IV U65445 ( .A(n52877), .Z(n52875) );
  NOR U65446 ( .A(n52875), .B(n52874), .Z(n52882) );
  NOR U65447 ( .A(n52877), .B(n52876), .Z(n52880) );
  IV U65448 ( .A(n52878), .Z(n52879) );
  NOR U65449 ( .A(n52880), .B(n52879), .Z(n52881) );
  NOR U65450 ( .A(n52882), .B(n52881), .Z(n57393) );
  IV U65451 ( .A(n52883), .Z(n52886) );
  IV U65452 ( .A(n52884), .Z(n52885) );
  NOR U65453 ( .A(n52886), .B(n52885), .Z(n57388) );
  NOR U65454 ( .A(n52888), .B(n52887), .Z(n52889) );
  IV U65455 ( .A(n52889), .Z(n57387) );
  IV U65456 ( .A(n57385), .Z(n56480) );
  XOR U65457 ( .A(n57387), .B(n56480), .Z(n52890) );
  NOR U65458 ( .A(n57388), .B(n52890), .Z(n53752) );
  IV U65459 ( .A(n52891), .Z(n52892) );
  NOR U65460 ( .A(n52895), .B(n52892), .Z(n56477) );
  IV U65461 ( .A(n52893), .Z(n52894) );
  NOR U65462 ( .A(n52895), .B(n52894), .Z(n57364) );
  IV U65463 ( .A(n52896), .Z(n52898) );
  NOR U65464 ( .A(n52898), .B(n52897), .Z(n57361) );
  NOR U65465 ( .A(n52900), .B(n52899), .Z(n52906) );
  IV U65466 ( .A(n52900), .Z(n52901) );
  NOR U65467 ( .A(n52902), .B(n52901), .Z(n52903) );
  NOR U65468 ( .A(n52904), .B(n52903), .Z(n52905) );
  NOR U65469 ( .A(n52906), .B(n52905), .Z(n57358) );
  IV U65470 ( .A(n52907), .Z(n52908) );
  NOR U65471 ( .A(n52915), .B(n52908), .Z(n57372) );
  IV U65472 ( .A(n52909), .Z(n52910) );
  NOR U65473 ( .A(n52910), .B(n52915), .Z(n52911) );
  IV U65474 ( .A(n52911), .Z(n57370) );
  NOR U65475 ( .A(n52913), .B(n52912), .Z(n57337) );
  IV U65476 ( .A(n52914), .Z(n52916) );
  NOR U65477 ( .A(n52916), .B(n52915), .Z(n56483) );
  NOR U65478 ( .A(n57337), .B(n56483), .Z(n53751) );
  IV U65479 ( .A(n52917), .Z(n52919) );
  NOR U65480 ( .A(n52919), .B(n52918), .Z(n57336) );
  IV U65481 ( .A(n52920), .Z(n52921) );
  NOR U65482 ( .A(n53734), .B(n52921), .Z(n52922) );
  IV U65483 ( .A(n52922), .Z(n57322) );
  IV U65484 ( .A(n52923), .Z(n52927) );
  NOR U65485 ( .A(n52925), .B(n52924), .Z(n52926) );
  IV U65486 ( .A(n52926), .Z(n53722) );
  NOR U65487 ( .A(n52927), .B(n53722), .Z(n57318) );
  IV U65488 ( .A(n52928), .Z(n52929) );
  NOR U65489 ( .A(n52929), .B(n53719), .Z(n53727) );
  NOR U65490 ( .A(n52931), .B(n52930), .Z(n52936) );
  IV U65491 ( .A(n52932), .Z(n52934) );
  NOR U65492 ( .A(n52934), .B(n52933), .Z(n52935) );
  NOR U65493 ( .A(n52936), .B(n52935), .Z(n57317) );
  IV U65494 ( .A(n52937), .Z(n52941) );
  NOR U65495 ( .A(n52939), .B(n52938), .Z(n52940) );
  IV U65496 ( .A(n52940), .Z(n52943) );
  NOR U65497 ( .A(n52941), .B(n52943), .Z(n56489) );
  IV U65498 ( .A(n52942), .Z(n52944) );
  NOR U65499 ( .A(n52944), .B(n52943), .Z(n56492) );
  IV U65500 ( .A(n52945), .Z(n52946) );
  NOR U65501 ( .A(n52947), .B(n52946), .Z(n52951) );
  NOR U65502 ( .A(n52949), .B(n52948), .Z(n52950) );
  NOR U65503 ( .A(n52951), .B(n52950), .Z(n57305) );
  NOR U65504 ( .A(n52953), .B(n52952), .Z(n52954) );
  NOR U65505 ( .A(n52954), .B(n53704), .Z(n53707) );
  IV U65506 ( .A(n52955), .Z(n52956) );
  NOR U65507 ( .A(n52957), .B(n52956), .Z(n57286) );
  IV U65508 ( .A(n52958), .Z(n52959) );
  NOR U65509 ( .A(n52959), .B(n53704), .Z(n57296) );
  NOR U65510 ( .A(n57286), .B(n57296), .Z(n53702) );
  IV U65511 ( .A(n52960), .Z(n52969) );
  IV U65512 ( .A(n52961), .Z(n52962) );
  NOR U65513 ( .A(n52969), .B(n52962), .Z(n52966) );
  IV U65514 ( .A(n52963), .Z(n52965) );
  NOR U65515 ( .A(n52965), .B(n52964), .Z(n57295) );
  NOR U65516 ( .A(n52966), .B(n57295), .Z(n57289) );
  IV U65517 ( .A(n57289), .Z(n57292) );
  IV U65518 ( .A(n52967), .Z(n52968) );
  NOR U65519 ( .A(n52969), .B(n52968), .Z(n57271) );
  IV U65520 ( .A(n52970), .Z(n52971) );
  NOR U65521 ( .A(n53700), .B(n52971), .Z(n57268) );
  IV U65522 ( .A(n52972), .Z(n52975) );
  NOR U65523 ( .A(n52973), .B(n52981), .Z(n52974) );
  IV U65524 ( .A(n52974), .Z(n52977) );
  NOR U65525 ( .A(n52975), .B(n52977), .Z(n57276) );
  IV U65526 ( .A(n52976), .Z(n52978) );
  NOR U65527 ( .A(n52978), .B(n52977), .Z(n56503) );
  IV U65528 ( .A(n52979), .Z(n52985) );
  IV U65529 ( .A(n52980), .Z(n52982) );
  NOR U65530 ( .A(n52982), .B(n52981), .Z(n52983) );
  IV U65531 ( .A(n52983), .Z(n52984) );
  NOR U65532 ( .A(n52985), .B(n52984), .Z(n56500) );
  IV U65533 ( .A(n52986), .Z(n52987) );
  NOR U65534 ( .A(n52988), .B(n52987), .Z(n57245) );
  IV U65535 ( .A(n52989), .Z(n52991) );
  NOR U65536 ( .A(n52991), .B(n52990), .Z(n52995) );
  IV U65537 ( .A(n52992), .Z(n52993) );
  NOR U65538 ( .A(n53694), .B(n52993), .Z(n52994) );
  NOR U65539 ( .A(n52995), .B(n52994), .Z(n56511) );
  IV U65540 ( .A(n52996), .Z(n52998) );
  NOR U65541 ( .A(n52998), .B(n52997), .Z(n56508) );
  IV U65542 ( .A(n52999), .Z(n57257) );
  IV U65543 ( .A(n57255), .Z(n57253) );
  XOR U65544 ( .A(n57257), .B(n57253), .Z(n53000) );
  NOR U65545 ( .A(n56508), .B(n53000), .Z(n53687) );
  IV U65546 ( .A(n53001), .Z(n53003) );
  NOR U65547 ( .A(n53003), .B(n53002), .Z(n56524) );
  IV U65548 ( .A(n53004), .Z(n53006) );
  IV U65549 ( .A(n53005), .Z(n53683) );
  NOR U65550 ( .A(n53006), .B(n53683), .Z(n53007) );
  IV U65551 ( .A(n53007), .Z(n56523) );
  IV U65552 ( .A(n53008), .Z(n53009) );
  NOR U65553 ( .A(n53009), .B(n53680), .Z(n53010) );
  IV U65554 ( .A(n53010), .Z(n53675) );
  IV U65555 ( .A(n53011), .Z(n53015) );
  IV U65556 ( .A(n53012), .Z(n53663) );
  NOR U65557 ( .A(n53013), .B(n53663), .Z(n53014) );
  IV U65558 ( .A(n53014), .Z(n53660) );
  NOR U65559 ( .A(n53015), .B(n53660), .Z(n57226) );
  IV U65560 ( .A(n53016), .Z(n53019) );
  IV U65561 ( .A(n53017), .Z(n53018) );
  NOR U65562 ( .A(n53019), .B(n53018), .Z(n57216) );
  NOR U65563 ( .A(n53021), .B(n53020), .Z(n57211) );
  IV U65564 ( .A(n53022), .Z(n53026) );
  NOR U65565 ( .A(n53024), .B(n53023), .Z(n53025) );
  IV U65566 ( .A(n53025), .Z(n53644) );
  NOR U65567 ( .A(n53026), .B(n53644), .Z(n57195) );
  IV U65568 ( .A(n53027), .Z(n53031) );
  NOR U65569 ( .A(n53029), .B(n53028), .Z(n53030) );
  IV U65570 ( .A(n53030), .Z(n53036) );
  NOR U65571 ( .A(n53031), .B(n53036), .Z(n57206) );
  IV U65572 ( .A(n53032), .Z(n53040) );
  IV U65573 ( .A(n53033), .Z(n53034) );
  NOR U65574 ( .A(n53040), .B(n53034), .Z(n56553) );
  IV U65575 ( .A(n53035), .Z(n53037) );
  NOR U65576 ( .A(n53037), .B(n53036), .Z(n57171) );
  NOR U65577 ( .A(n56553), .B(n57171), .Z(n53636) );
  IV U65578 ( .A(n53038), .Z(n53039) );
  NOR U65579 ( .A(n53040), .B(n53039), .Z(n57164) );
  IV U65580 ( .A(n53041), .Z(n53043) );
  NOR U65581 ( .A(n53043), .B(n53042), .Z(n57161) );
  IV U65582 ( .A(n53044), .Z(n53046) );
  NOR U65583 ( .A(n53046), .B(n53045), .Z(n56566) );
  IV U65584 ( .A(n53047), .Z(n53049) );
  IV U65585 ( .A(n53048), .Z(n53617) );
  NOR U65586 ( .A(n53049), .B(n53617), .Z(n56571) );
  IV U65587 ( .A(n53050), .Z(n53051) );
  NOR U65588 ( .A(n53052), .B(n53051), .Z(n53611) );
  IV U65589 ( .A(n53053), .Z(n53055) );
  IV U65590 ( .A(n53054), .Z(n53057) );
  NOR U65591 ( .A(n53055), .B(n53057), .Z(n53608) );
  IV U65592 ( .A(n53056), .Z(n53058) );
  NOR U65593 ( .A(n53058), .B(n53057), .Z(n53059) );
  IV U65594 ( .A(n53059), .Z(n56546) );
  NOR U65595 ( .A(n53062), .B(n53060), .Z(n56542) );
  IV U65596 ( .A(n53061), .Z(n53063) );
  NOR U65597 ( .A(n53063), .B(n53062), .Z(n53064) );
  IV U65598 ( .A(n53064), .Z(n53065) );
  NOR U65599 ( .A(n53066), .B(n53065), .Z(n56560) );
  NOR U65600 ( .A(n53068), .B(n53067), .Z(n53069) );
  IV U65601 ( .A(n53069), .Z(n53071) );
  NOR U65602 ( .A(n53071), .B(n53070), .Z(n56557) );
  IV U65603 ( .A(n53072), .Z(n53074) );
  NOR U65604 ( .A(n53074), .B(n53073), .Z(n57137) );
  IV U65605 ( .A(n53075), .Z(n53076) );
  NOR U65606 ( .A(n53077), .B(n53076), .Z(n57128) );
  NOR U65607 ( .A(n57137), .B(n57128), .Z(n53604) );
  IV U65608 ( .A(n53078), .Z(n53079) );
  NOR U65609 ( .A(n53080), .B(n53079), .Z(n57139) );
  IV U65610 ( .A(n57139), .Z(n57136) );
  IV U65611 ( .A(n53081), .Z(n53083) );
  IV U65612 ( .A(n53082), .Z(n53088) );
  NOR U65613 ( .A(n53083), .B(n53088), .Z(n53084) );
  IV U65614 ( .A(n53084), .Z(n57084) );
  IV U65615 ( .A(n53085), .Z(n53086) );
  NOR U65616 ( .A(n53086), .B(n53088), .Z(n57089) );
  IV U65617 ( .A(n53087), .Z(n53089) );
  NOR U65618 ( .A(n53089), .B(n53088), .Z(n57086) );
  IV U65619 ( .A(n53090), .Z(n53091) );
  NOR U65620 ( .A(n53091), .B(n53094), .Z(n57115) );
  IV U65621 ( .A(n53092), .Z(n53093) );
  NOR U65622 ( .A(n53094), .B(n53093), .Z(n57112) );
  IV U65623 ( .A(n53095), .Z(n53096) );
  NOR U65624 ( .A(n53096), .B(n53578), .Z(n53580) );
  IV U65625 ( .A(n53097), .Z(n53099) );
  NOR U65626 ( .A(n53099), .B(n53098), .Z(n57074) );
  IV U65627 ( .A(n53102), .Z(n53100) );
  NOR U65628 ( .A(n53101), .B(n53100), .Z(n53108) );
  NOR U65629 ( .A(n53103), .B(n53102), .Z(n53106) );
  IV U65630 ( .A(n53104), .Z(n53105) );
  NOR U65631 ( .A(n53106), .B(n53105), .Z(n53107) );
  NOR U65632 ( .A(n53108), .B(n53107), .Z(n57057) );
  IV U65633 ( .A(n53109), .Z(n53110) );
  NOR U65634 ( .A(n53111), .B(n53110), .Z(n53115) );
  NOR U65635 ( .A(n53113), .B(n53112), .Z(n53114) );
  NOR U65636 ( .A(n53115), .B(n53114), .Z(n57054) );
  IV U65637 ( .A(n53116), .Z(n53117) );
  NOR U65638 ( .A(n53119), .B(n53117), .Z(n57063) );
  IV U65639 ( .A(n53118), .Z(n53120) );
  NOR U65640 ( .A(n53120), .B(n53119), .Z(n53121) );
  IV U65641 ( .A(n53121), .Z(n57062) );
  IV U65642 ( .A(n53122), .Z(n53124) );
  NOR U65643 ( .A(n53124), .B(n53123), .Z(n53125) );
  NOR U65644 ( .A(n53126), .B(n53125), .Z(n57052) );
  IV U65645 ( .A(n53127), .Z(n53128) );
  NOR U65646 ( .A(n53129), .B(n53128), .Z(n57022) );
  IV U65647 ( .A(n57034), .Z(n53134) );
  NOR U65648 ( .A(n53130), .B(n53134), .Z(n57027) );
  NOR U65649 ( .A(n53132), .B(n53131), .Z(n53136) );
  IV U65650 ( .A(n53133), .Z(n53135) );
  NOR U65651 ( .A(n53135), .B(n53134), .Z(n57038) );
  NOR U65652 ( .A(n53136), .B(n57038), .Z(n53565) );
  IV U65653 ( .A(n53137), .Z(n53140) );
  IV U65654 ( .A(n53138), .Z(n53139) );
  NOR U65655 ( .A(n53140), .B(n53139), .Z(n56595) );
  IV U65656 ( .A(n56595), .Z(n56601) );
  NOR U65657 ( .A(n53142), .B(n53141), .Z(n53143) );
  NOR U65658 ( .A(n53143), .B(n53146), .Z(n53144) );
  IV U65659 ( .A(n53144), .Z(n56599) );
  IV U65660 ( .A(n53145), .Z(n53147) );
  NOR U65661 ( .A(n53147), .B(n53146), .Z(n56590) );
  IV U65662 ( .A(n53148), .Z(n53150) );
  NOR U65663 ( .A(n53150), .B(n53149), .Z(n53557) );
  IV U65664 ( .A(n53151), .Z(n53152) );
  NOR U65665 ( .A(n53153), .B(n53152), .Z(n56581) );
  IV U65666 ( .A(n53154), .Z(n53155) );
  NOR U65667 ( .A(n53156), .B(n53155), .Z(n53558) );
  NOR U65668 ( .A(n56581), .B(n53558), .Z(n53555) );
  NOR U65669 ( .A(n53158), .B(n53157), .Z(n56614) );
  IV U65670 ( .A(n53159), .Z(n53160) );
  NOR U65671 ( .A(n53161), .B(n53160), .Z(n53166) );
  IV U65672 ( .A(n53162), .Z(n53164) );
  NOR U65673 ( .A(n53164), .B(n53163), .Z(n53165) );
  NOR U65674 ( .A(n53166), .B(n53165), .Z(n57005) );
  NOR U65675 ( .A(n53169), .B(n53167), .Z(n53529) );
  IV U65676 ( .A(n53168), .Z(n53170) );
  NOR U65677 ( .A(n53170), .B(n53169), .Z(n53527) );
  IV U65678 ( .A(n53171), .Z(n53173) );
  NOR U65679 ( .A(n53173), .B(n53172), .Z(n56974) );
  NOR U65680 ( .A(n53174), .B(n53175), .Z(n53181) );
  IV U65681 ( .A(n53175), .Z(n53176) );
  NOR U65682 ( .A(n53177), .B(n53176), .Z(n53178) );
  NOR U65683 ( .A(n53179), .B(n53178), .Z(n53180) );
  NOR U65684 ( .A(n53181), .B(n53180), .Z(n56984) );
  IV U65685 ( .A(n53182), .Z(n53183) );
  NOR U65686 ( .A(n53184), .B(n53183), .Z(n53188) );
  NOR U65687 ( .A(n53186), .B(n53185), .Z(n53187) );
  NOR U65688 ( .A(n53188), .B(n53187), .Z(n56982) );
  IV U65689 ( .A(n53189), .Z(n53190) );
  NOR U65690 ( .A(n53190), .B(n53191), .Z(n56955) );
  NOR U65691 ( .A(n53192), .B(n53191), .Z(n56963) );
  IV U65692 ( .A(n53193), .Z(n53194) );
  NOR U65693 ( .A(n53195), .B(n53194), .Z(n53489) );
  IV U65694 ( .A(n53489), .Z(n53484) );
  IV U65695 ( .A(n53196), .Z(n53197) );
  NOR U65696 ( .A(n53198), .B(n53197), .Z(n56642) );
  IV U65697 ( .A(n53199), .Z(n53200) );
  NOR U65698 ( .A(n53207), .B(n53200), .Z(n56658) );
  IV U65699 ( .A(n53201), .Z(n53202) );
  NOR U65700 ( .A(n53202), .B(n53205), .Z(n56655) );
  IV U65701 ( .A(n53203), .Z(n53204) );
  NOR U65702 ( .A(n53205), .B(n53204), .Z(n53210) );
  IV U65703 ( .A(n53206), .Z(n53208) );
  NOR U65704 ( .A(n53208), .B(n53207), .Z(n53209) );
  NOR U65705 ( .A(n53210), .B(n53209), .Z(n56653) );
  IV U65706 ( .A(n53211), .Z(n53212) );
  NOR U65707 ( .A(n53213), .B(n53212), .Z(n56935) );
  IV U65708 ( .A(n53214), .Z(n53216) );
  NOR U65709 ( .A(n53216), .B(n53215), .Z(n56649) );
  NOR U65710 ( .A(n56935), .B(n56649), .Z(n53482) );
  IV U65711 ( .A(n53217), .Z(n53218) );
  NOR U65712 ( .A(n53219), .B(n53218), .Z(n56934) );
  IV U65713 ( .A(n53220), .Z(n53221) );
  NOR U65714 ( .A(n53221), .B(n53223), .Z(n56919) );
  IV U65715 ( .A(n53222), .Z(n53224) );
  NOR U65716 ( .A(n53224), .B(n53223), .Z(n56916) );
  IV U65717 ( .A(n53225), .Z(n53226) );
  NOR U65718 ( .A(n53229), .B(n53226), .Z(n56927) );
  IV U65719 ( .A(n53227), .Z(n53228) );
  NOR U65720 ( .A(n53229), .B(n53228), .Z(n56924) );
  IV U65721 ( .A(n53230), .Z(n53231) );
  NOR U65722 ( .A(n53231), .B(n53479), .Z(n53236) );
  IV U65723 ( .A(n53232), .Z(n53234) );
  NOR U65724 ( .A(n53234), .B(n53233), .Z(n53235) );
  NOR U65725 ( .A(n53236), .B(n53235), .Z(n56667) );
  IV U65726 ( .A(n53237), .Z(n53239) );
  NOR U65727 ( .A(n53239), .B(n53238), .Z(n56907) );
  IV U65728 ( .A(n53240), .Z(n53241) );
  NOR U65729 ( .A(n53241), .B(n53244), .Z(n56888) );
  IV U65730 ( .A(n53242), .Z(n53243) );
  NOR U65731 ( .A(n53244), .B(n53243), .Z(n56885) );
  IV U65732 ( .A(n53245), .Z(n53246) );
  NOR U65733 ( .A(n53246), .B(n53248), .Z(n56669) );
  IV U65734 ( .A(n53247), .Z(n53249) );
  NOR U65735 ( .A(n53249), .B(n53248), .Z(n56685) );
  IV U65736 ( .A(n53250), .Z(n53252) );
  NOR U65737 ( .A(n53252), .B(n53251), .Z(n56840) );
  IV U65738 ( .A(n53253), .Z(n53254) );
  NOR U65739 ( .A(n53257), .B(n53254), .Z(n56846) );
  IV U65740 ( .A(n53255), .Z(n53256) );
  NOR U65741 ( .A(n53257), .B(n53256), .Z(n56843) );
  IV U65742 ( .A(n53258), .Z(n53448) );
  NOR U65743 ( .A(n53259), .B(n53448), .Z(n56833) );
  NOR U65744 ( .A(n53261), .B(n53260), .Z(n56691) );
  IV U65745 ( .A(n53262), .Z(n53263) );
  NOR U65746 ( .A(n53263), .B(n53433), .Z(n53441) );
  IV U65747 ( .A(n53441), .Z(n53439) );
  IV U65748 ( .A(n53264), .Z(n53265) );
  NOR U65749 ( .A(n53265), .B(n53433), .Z(n53266) );
  IV U65750 ( .A(n53266), .Z(n56810) );
  IV U65751 ( .A(n53267), .Z(n53268) );
  NOR U65752 ( .A(n53269), .B(n53268), .Z(n56812) );
  IV U65753 ( .A(n53270), .Z(n53271) );
  NOR U65754 ( .A(n53279), .B(n53271), .Z(n53276) );
  IV U65755 ( .A(n53272), .Z(n53274) );
  IV U65756 ( .A(n53273), .Z(n53427) );
  NOR U65757 ( .A(n53274), .B(n53427), .Z(n53275) );
  NOR U65758 ( .A(n53276), .B(n53275), .Z(n56700) );
  IV U65759 ( .A(n53277), .Z(n53278) );
  NOR U65760 ( .A(n53279), .B(n53278), .Z(n56696) );
  IV U65761 ( .A(n53280), .Z(n53283) );
  IV U65762 ( .A(n53281), .Z(n53282) );
  NOR U65763 ( .A(n53283), .B(n53282), .Z(n56788) );
  IV U65764 ( .A(n53284), .Z(n53288) );
  NOR U65765 ( .A(n53286), .B(n53285), .Z(n53287) );
  IV U65766 ( .A(n53287), .Z(n53421) );
  NOR U65767 ( .A(n53288), .B(n53421), .Z(n56785) );
  IV U65768 ( .A(n53289), .Z(n53291) );
  NOR U65769 ( .A(n53291), .B(n53290), .Z(n53296) );
  IV U65770 ( .A(n53292), .Z(n53294) );
  NOR U65771 ( .A(n53294), .B(n53293), .Z(n53295) );
  NOR U65772 ( .A(n53296), .B(n53295), .Z(n56797) );
  IV U65773 ( .A(n53297), .Z(n53299) );
  IV U65774 ( .A(n53298), .Z(n53405) );
  NOR U65775 ( .A(n53299), .B(n53405), .Z(n53300) );
  IV U65776 ( .A(n53300), .Z(n53415) );
  IV U65777 ( .A(n53301), .Z(n53303) );
  NOR U65778 ( .A(n53303), .B(n53302), .Z(n53396) );
  IV U65779 ( .A(n53304), .Z(n53306) );
  NOR U65780 ( .A(n53306), .B(n53305), .Z(n53307) );
  IV U65781 ( .A(n53307), .Z(n56712) );
  IV U65782 ( .A(n53389), .Z(n53367) );
  IV U65783 ( .A(n53308), .Z(n53309) );
  NOR U65784 ( .A(n53310), .B(n53309), .Z(n53315) );
  IV U65785 ( .A(n53311), .Z(n53313) );
  NOR U65786 ( .A(n53313), .B(n53312), .Z(n53314) );
  NOR U65787 ( .A(n53315), .B(n53314), .Z(n56722) );
  IV U65788 ( .A(n53316), .Z(n53320) );
  NOR U65789 ( .A(n53318), .B(n53317), .Z(n53319) );
  IV U65790 ( .A(n53319), .Z(n53322) );
  NOR U65791 ( .A(n53320), .B(n53322), .Z(n56753) );
  IV U65792 ( .A(n56753), .Z(n56754) );
  IV U65793 ( .A(n53321), .Z(n53323) );
  NOR U65794 ( .A(n53323), .B(n53322), .Z(n56723) );
  NOR U65795 ( .A(n56742), .B(n56723), .Z(n53356) );
  IV U65796 ( .A(n53324), .Z(n53325) );
  NOR U65797 ( .A(n53326), .B(n53325), .Z(n53327) );
  IV U65798 ( .A(n53327), .Z(n53350) );
  IV U65799 ( .A(n53328), .Z(n53329) );
  NOR U65800 ( .A(n53329), .B(n53338), .Z(n56729) );
  IV U65801 ( .A(n53330), .Z(n53331) );
  NOR U65802 ( .A(n53332), .B(n53331), .Z(n53336) );
  NOR U65803 ( .A(n53334), .B(n53333), .Z(n53335) );
  NOR U65804 ( .A(n53336), .B(n53335), .Z(n56728) );
  IV U65805 ( .A(n53337), .Z(n53339) );
  NOR U65806 ( .A(n53339), .B(n53338), .Z(n56726) );
  XOR U65807 ( .A(n56728), .B(n56726), .Z(n56730) );
  XOR U65808 ( .A(n56729), .B(n56730), .Z(n53347) );
  NOR U65809 ( .A(n53350), .B(n53347), .Z(n53345) );
  IV U65810 ( .A(n53340), .Z(n53341) );
  NOR U65811 ( .A(n53342), .B(n53341), .Z(n53348) );
  IV U65812 ( .A(n53348), .Z(n53343) );
  NOR U65813 ( .A(n56730), .B(n53343), .Z(n53344) );
  NOR U65814 ( .A(n53345), .B(n53344), .Z(n53346) );
  IV U65815 ( .A(n53346), .Z(n56738) );
  IV U65816 ( .A(n53347), .Z(n53351) );
  NOR U65817 ( .A(n53348), .B(n53351), .Z(n53349) );
  NOR U65818 ( .A(n56738), .B(n53349), .Z(n53353) );
  NOR U65819 ( .A(n53351), .B(n53350), .Z(n53352) );
  NOR U65820 ( .A(n53353), .B(n53352), .Z(n56736) );
  NOR U65821 ( .A(n53355), .B(n53354), .Z(n56734) );
  XOR U65822 ( .A(n56736), .B(n56734), .Z(n56743) );
  XOR U65823 ( .A(n56744), .B(n56743), .Z(n56724) );
  XOR U65824 ( .A(n53356), .B(n56724), .Z(n56752) );
  IV U65825 ( .A(n56752), .Z(n56755) );
  XOR U65826 ( .A(n56754), .B(n56755), .Z(n53357) );
  XOR U65827 ( .A(n53358), .B(n53357), .Z(n56721) );
  XOR U65828 ( .A(n56722), .B(n56721), .Z(n53378) );
  IV U65829 ( .A(n53378), .Z(n56768) );
  IV U65830 ( .A(n53359), .Z(n53360) );
  NOR U65831 ( .A(n53361), .B(n53360), .Z(n53377) );
  IV U65832 ( .A(n53362), .Z(n53363) );
  NOR U65833 ( .A(n53364), .B(n53363), .Z(n56767) );
  NOR U65834 ( .A(n53377), .B(n56767), .Z(n53365) );
  XOR U65835 ( .A(n56768), .B(n53365), .Z(n53384) );
  IV U65836 ( .A(n53384), .Z(n53366) );
  NOR U65837 ( .A(n53367), .B(n53366), .Z(n56774) );
  IV U65838 ( .A(n53368), .Z(n53375) );
  NOR U65839 ( .A(n53370), .B(n53369), .Z(n53371) );
  IV U65840 ( .A(n53371), .Z(n53372) );
  NOR U65841 ( .A(n53373), .B(n53372), .Z(n53374) );
  IV U65842 ( .A(n53374), .Z(n53380) );
  NOR U65843 ( .A(n53375), .B(n53380), .Z(n53376) );
  IV U65844 ( .A(n53376), .Z(n56718) );
  IV U65845 ( .A(n53377), .Z(n56766) );
  XOR U65846 ( .A(n56766), .B(n53378), .Z(n53383) );
  IV U65847 ( .A(n53379), .Z(n53381) );
  NOR U65848 ( .A(n53381), .B(n53380), .Z(n53385) );
  IV U65849 ( .A(n53385), .Z(n53382) );
  NOR U65850 ( .A(n53383), .B(n53382), .Z(n56720) );
  NOR U65851 ( .A(n53385), .B(n53384), .Z(n53386) );
  NOR U65852 ( .A(n56720), .B(n53386), .Z(n53387) );
  IV U65853 ( .A(n53387), .Z(n56717) );
  XOR U65854 ( .A(n56718), .B(n56717), .Z(n53388) );
  NOR U65855 ( .A(n53389), .B(n53388), .Z(n53390) );
  NOR U65856 ( .A(n56774), .B(n53390), .Z(n53391) );
  IV U65857 ( .A(n53391), .Z(n56709) );
  XOR U65858 ( .A(n56708), .B(n56709), .Z(n56711) );
  XOR U65859 ( .A(n56712), .B(n56711), .Z(n53392) );
  NOR U65860 ( .A(n53396), .B(n53392), .Z(n53411) );
  IV U65861 ( .A(n53393), .Z(n53395) );
  NOR U65862 ( .A(n53395), .B(n53394), .Z(n53401) );
  IV U65863 ( .A(n53396), .Z(n53397) );
  NOR U65864 ( .A(n56711), .B(n53397), .Z(n53398) );
  NOR U65865 ( .A(n53401), .B(n53398), .Z(n53399) );
  NOR U65866 ( .A(n53411), .B(n53399), .Z(n56716) );
  IV U65867 ( .A(n53411), .Z(n53400) );
  NOR U65868 ( .A(n53401), .B(n53400), .Z(n53402) );
  NOR U65869 ( .A(n56716), .B(n53402), .Z(n53412) );
  IV U65870 ( .A(n53412), .Z(n53403) );
  NOR U65871 ( .A(n53415), .B(n53403), .Z(n56782) );
  IV U65872 ( .A(n53404), .Z(n53406) );
  NOR U65873 ( .A(n53406), .B(n53405), .Z(n53407) );
  IV U65874 ( .A(n53407), .Z(n56794) );
  NOR U65875 ( .A(n53409), .B(n53408), .Z(n53413) );
  IV U65876 ( .A(n53413), .Z(n53410) );
  NOR U65877 ( .A(n53411), .B(n53410), .Z(n56715) );
  NOR U65878 ( .A(n53413), .B(n53412), .Z(n53414) );
  NOR U65879 ( .A(n56715), .B(n53414), .Z(n53416) );
  IV U65880 ( .A(n53416), .Z(n56793) );
  XOR U65881 ( .A(n56794), .B(n56793), .Z(n53418) );
  NOR U65882 ( .A(n53416), .B(n53415), .Z(n53417) );
  NOR U65883 ( .A(n53418), .B(n53417), .Z(n53419) );
  NOR U65884 ( .A(n56782), .B(n53419), .Z(n56795) );
  XOR U65885 ( .A(n56797), .B(n56795), .Z(n56706) );
  IV U65886 ( .A(n56706), .Z(n53425) );
  IV U65887 ( .A(n53420), .Z(n53422) );
  NOR U65888 ( .A(n53422), .B(n53421), .Z(n53423) );
  NOR U65889 ( .A(n53424), .B(n53423), .Z(n56707) );
  XOR U65890 ( .A(n53425), .B(n56707), .Z(n56787) );
  XOR U65891 ( .A(n56785), .B(n56787), .Z(n56789) );
  XOR U65892 ( .A(n56788), .B(n56789), .Z(n56697) );
  XOR U65893 ( .A(n56696), .B(n56697), .Z(n56699) );
  XOR U65894 ( .A(n56700), .B(n56699), .Z(n56701) );
  IV U65895 ( .A(n53426), .Z(n53428) );
  NOR U65896 ( .A(n53428), .B(n53427), .Z(n53429) );
  IV U65897 ( .A(n53429), .Z(n56702) );
  XOR U65898 ( .A(n56701), .B(n56702), .Z(n56813) );
  XOR U65899 ( .A(n56812), .B(n56813), .Z(n56815) );
  IV U65900 ( .A(n56815), .Z(n53437) );
  IV U65901 ( .A(n53430), .Z(n53431) );
  NOR U65902 ( .A(n53432), .B(n53431), .Z(n53436) );
  NOR U65903 ( .A(n53434), .B(n53433), .Z(n53435) );
  NOR U65904 ( .A(n53436), .B(n53435), .Z(n56816) );
  XOR U65905 ( .A(n53437), .B(n56816), .Z(n56811) );
  XOR U65906 ( .A(n56810), .B(n56811), .Z(n53440) );
  IV U65907 ( .A(n53440), .Z(n53438) );
  NOR U65908 ( .A(n53439), .B(n53438), .Z(n56832) );
  NOR U65909 ( .A(n53441), .B(n53440), .Z(n56830) );
  IV U65910 ( .A(n53442), .Z(n53443) );
  NOR U65911 ( .A(n53444), .B(n53443), .Z(n56828) );
  XOR U65912 ( .A(n56830), .B(n56828), .Z(n53445) );
  NOR U65913 ( .A(n56832), .B(n53445), .Z(n53446) );
  IV U65914 ( .A(n53446), .Z(n56689) );
  XOR U65915 ( .A(n56688), .B(n56689), .Z(n56692) );
  XOR U65916 ( .A(n56691), .B(n56692), .Z(n56834) );
  XOR U65917 ( .A(n56833), .B(n56834), .Z(n56679) );
  IV U65918 ( .A(n53447), .Z(n53449) );
  NOR U65919 ( .A(n53449), .B(n53448), .Z(n56677) );
  XOR U65920 ( .A(n56679), .B(n56677), .Z(n56682) );
  IV U65921 ( .A(n53450), .Z(n53452) );
  NOR U65922 ( .A(n53452), .B(n53451), .Z(n56680) );
  XOR U65923 ( .A(n56682), .B(n56680), .Z(n56844) );
  XOR U65924 ( .A(n56843), .B(n56844), .Z(n56847) );
  XOR U65925 ( .A(n56846), .B(n56847), .Z(n56841) );
  XOR U65926 ( .A(n56840), .B(n56841), .Z(n56857) );
  XOR U65927 ( .A(n56856), .B(n56857), .Z(n56859) );
  IV U65928 ( .A(n53453), .Z(n53455) );
  NOR U65929 ( .A(n53455), .B(n53454), .Z(n53456) );
  NOR U65930 ( .A(n53457), .B(n53456), .Z(n56860) );
  XOR U65931 ( .A(n56859), .B(n56860), .Z(n53458) );
  IV U65932 ( .A(n53458), .Z(n56876) );
  NOR U65933 ( .A(n56869), .B(n53459), .Z(n53460) );
  NOR U65934 ( .A(n53460), .B(n56870), .Z(n53461) );
  XOR U65935 ( .A(n56876), .B(n53461), .Z(n56879) );
  IV U65936 ( .A(n53462), .Z(n53464) );
  NOR U65937 ( .A(n53464), .B(n53463), .Z(n56878) );
  IV U65938 ( .A(n53465), .Z(n53466) );
  NOR U65939 ( .A(n53466), .B(n56870), .Z(n53467) );
  NOR U65940 ( .A(n56878), .B(n53467), .Z(n53468) );
  XOR U65941 ( .A(n56879), .B(n53468), .Z(n53469) );
  IV U65942 ( .A(n53469), .Z(n56686) );
  XOR U65943 ( .A(n56685), .B(n56686), .Z(n56670) );
  XOR U65944 ( .A(n56669), .B(n56670), .Z(n56673) );
  XOR U65945 ( .A(n56672), .B(n56673), .Z(n56896) );
  IV U65946 ( .A(n56896), .Z(n53474) );
  IV U65947 ( .A(n53470), .Z(n53472) );
  NOR U65948 ( .A(n53472), .B(n53471), .Z(n56895) );
  NOR U65949 ( .A(n56893), .B(n56895), .Z(n53473) );
  XOR U65950 ( .A(n53474), .B(n53473), .Z(n56886) );
  XOR U65951 ( .A(n56885), .B(n56886), .Z(n56889) );
  XOR U65952 ( .A(n56888), .B(n56889), .Z(n56908) );
  XOR U65953 ( .A(n56907), .B(n56908), .Z(n56665) );
  IV U65954 ( .A(n53475), .Z(n53477) );
  NOR U65955 ( .A(n53477), .B(n53476), .Z(n56906) );
  IV U65956 ( .A(n53478), .Z(n53480) );
  NOR U65957 ( .A(n53480), .B(n53479), .Z(n56663) );
  NOR U65958 ( .A(n56906), .B(n56663), .Z(n53481) );
  XOR U65959 ( .A(n56665), .B(n53481), .Z(n56666) );
  XOR U65960 ( .A(n56667), .B(n56666), .Z(n56925) );
  XOR U65961 ( .A(n56924), .B(n56925), .Z(n56928) );
  XOR U65962 ( .A(n56927), .B(n56928), .Z(n56917) );
  XOR U65963 ( .A(n56916), .B(n56917), .Z(n56920) );
  XOR U65964 ( .A(n56919), .B(n56920), .Z(n56936) );
  XOR U65965 ( .A(n56934), .B(n56936), .Z(n56651) );
  XOR U65966 ( .A(n53482), .B(n56651), .Z(n56652) );
  XOR U65967 ( .A(n56653), .B(n56652), .Z(n56656) );
  XOR U65968 ( .A(n56655), .B(n56656), .Z(n56659) );
  XOR U65969 ( .A(n56658), .B(n56659), .Z(n56645) );
  XOR U65970 ( .A(n56642), .B(n56645), .Z(n53483) );
  NOR U65971 ( .A(n53484), .B(n53483), .Z(n56949) );
  IV U65972 ( .A(n53485), .Z(n53486) );
  NOR U65973 ( .A(n53487), .B(n53486), .Z(n56644) );
  NOR U65974 ( .A(n56642), .B(n56644), .Z(n53488) );
  XOR U65975 ( .A(n53488), .B(n56645), .Z(n56638) );
  NOR U65976 ( .A(n53489), .B(n56638), .Z(n53490) );
  NOR U65977 ( .A(n56949), .B(n53490), .Z(n53491) );
  IV U65978 ( .A(n53491), .Z(n56637) );
  IV U65979 ( .A(n53492), .Z(n53494) );
  NOR U65980 ( .A(n53494), .B(n53493), .Z(n56639) );
  IV U65981 ( .A(n53495), .Z(n53497) );
  NOR U65982 ( .A(n53497), .B(n53496), .Z(n56635) );
  NOR U65983 ( .A(n56639), .B(n56635), .Z(n53498) );
  XOR U65984 ( .A(n56637), .B(n53498), .Z(n56960) );
  IV U65985 ( .A(n53499), .Z(n53500) );
  NOR U65986 ( .A(n53501), .B(n53500), .Z(n53505) );
  IV U65987 ( .A(n53502), .Z(n53503) );
  NOR U65988 ( .A(n53503), .B(n53508), .Z(n53504) );
  NOR U65989 ( .A(n53505), .B(n53504), .Z(n56961) );
  XOR U65990 ( .A(n56960), .B(n56961), .Z(n56964) );
  XOR U65991 ( .A(n56963), .B(n56964), .Z(n56954) );
  IV U65992 ( .A(n53506), .Z(n53507) );
  NOR U65993 ( .A(n53508), .B(n53507), .Z(n56952) );
  XOR U65994 ( .A(n56954), .B(n56952), .Z(n56956) );
  XOR U65995 ( .A(n56955), .B(n56956), .Z(n56981) );
  XOR U65996 ( .A(n56982), .B(n56981), .Z(n56983) );
  XOR U65997 ( .A(n56984), .B(n56983), .Z(n56996) );
  IV U65998 ( .A(n53509), .Z(n53511) );
  NOR U65999 ( .A(n53511), .B(n53510), .Z(n56995) );
  IV U66000 ( .A(n56995), .Z(n56998) );
  IV U66001 ( .A(n53512), .Z(n53513) );
  NOR U66002 ( .A(n53514), .B(n53513), .Z(n53518) );
  IV U66003 ( .A(n53515), .Z(n53516) );
  NOR U66004 ( .A(n53516), .B(n53522), .Z(n53517) );
  NOR U66005 ( .A(n53518), .B(n53517), .Z(n53519) );
  IV U66006 ( .A(n53519), .Z(n57000) );
  XOR U66007 ( .A(n56998), .B(n57000), .Z(n53520) );
  XOR U66008 ( .A(n56996), .B(n53520), .Z(n56976) );
  XOR U66009 ( .A(n56974), .B(n56976), .Z(n56978) );
  IV U66010 ( .A(n53521), .Z(n53523) );
  NOR U66011 ( .A(n53523), .B(n53522), .Z(n53524) );
  IV U66012 ( .A(n53524), .Z(n56977) );
  XOR U66013 ( .A(n56978), .B(n56977), .Z(n53525) );
  NOR U66014 ( .A(n53527), .B(n53525), .Z(n53530) );
  IV U66015 ( .A(n53530), .Z(n53526) );
  NOR U66016 ( .A(n53529), .B(n53526), .Z(n57006) );
  IV U66017 ( .A(n53527), .Z(n53528) );
  NOR U66018 ( .A(n53528), .B(n56976), .Z(n53533) );
  IV U66019 ( .A(n53529), .Z(n53531) );
  NOR U66020 ( .A(n53531), .B(n53530), .Z(n53532) );
  NOR U66021 ( .A(n53533), .B(n53532), .Z(n53534) );
  IV U66022 ( .A(n53534), .Z(n57007) );
  NOR U66023 ( .A(n57006), .B(n57007), .Z(n53535) );
  XOR U66024 ( .A(n57005), .B(n53535), .Z(n56616) );
  XOR U66025 ( .A(n56614), .B(n56616), .Z(n56617) );
  NOR U66026 ( .A(n53537), .B(n53536), .Z(n53544) );
  XOR U66027 ( .A(n56617), .B(n56618), .Z(n56621) );
  IV U66028 ( .A(n53543), .Z(n53546) );
  IV U66029 ( .A(n53544), .Z(n53545) );
  NOR U66030 ( .A(n53546), .B(n53545), .Z(n56622) );
  XOR U66031 ( .A(n53548), .B(n53547), .Z(n53549) );
  IV U66032 ( .A(n53549), .Z(n53550) );
  NOR U66033 ( .A(n53551), .B(n53550), .Z(n53552) );
  NOR U66034 ( .A(n56629), .B(n53552), .Z(n53553) );
  XOR U66035 ( .A(n56622), .B(n53553), .Z(n53554) );
  XOR U66036 ( .A(n56621), .B(n53554), .Z(n56583) );
  IV U66037 ( .A(n56583), .Z(n56586) );
  XOR U66038 ( .A(n53555), .B(n56586), .Z(n53556) );
  NOR U66039 ( .A(n53557), .B(n53556), .Z(n53561) );
  IV U66040 ( .A(n53557), .Z(n56587) );
  IV U66041 ( .A(n53558), .Z(n56589) );
  XOR U66042 ( .A(n56589), .B(n56583), .Z(n53559) );
  NOR U66043 ( .A(n56587), .B(n53559), .Z(n53560) );
  NOR U66044 ( .A(n53561), .B(n53560), .Z(n56591) );
  XOR U66045 ( .A(n56590), .B(n56591), .Z(n56598) );
  XOR U66046 ( .A(n56599), .B(n56598), .Z(n56600) );
  XOR U66047 ( .A(n56601), .B(n56600), .Z(n57036) );
  IV U66048 ( .A(n53562), .Z(n53563) );
  NOR U66049 ( .A(n56596), .B(n53563), .Z(n53564) );
  XOR U66050 ( .A(n57036), .B(n53564), .Z(n57039) );
  XOR U66051 ( .A(n53565), .B(n57039), .Z(n53566) );
  IV U66052 ( .A(n53566), .Z(n57029) );
  XOR U66053 ( .A(n57027), .B(n57029), .Z(n57021) );
  IV U66054 ( .A(n53567), .Z(n53568) );
  NOR U66055 ( .A(n53569), .B(n53568), .Z(n57019) );
  XOR U66056 ( .A(n57021), .B(n57019), .Z(n57023) );
  XOR U66057 ( .A(n57022), .B(n57023), .Z(n57051) );
  XOR U66058 ( .A(n57052), .B(n57051), .Z(n57060) );
  XOR U66059 ( .A(n57062), .B(n57060), .Z(n57064) );
  XOR U66060 ( .A(n57063), .B(n57064), .Z(n57053) );
  XOR U66061 ( .A(n57054), .B(n57053), .Z(n57055) );
  XOR U66062 ( .A(n57057), .B(n57055), .Z(n57076) );
  XOR U66063 ( .A(n57074), .B(n57076), .Z(n56580) );
  IV U66064 ( .A(n53570), .Z(n53571) );
  NOR U66065 ( .A(n53572), .B(n53571), .Z(n57075) );
  IV U66066 ( .A(n53573), .Z(n53574) );
  NOR U66067 ( .A(n53574), .B(n53578), .Z(n56578) );
  NOR U66068 ( .A(n57075), .B(n56578), .Z(n53575) );
  XOR U66069 ( .A(n56580), .B(n53575), .Z(n53576) );
  NOR U66070 ( .A(n53580), .B(n53576), .Z(n53584) );
  IV U66071 ( .A(n53577), .Z(n53579) );
  NOR U66072 ( .A(n53579), .B(n53578), .Z(n53585) );
  IV U66073 ( .A(n53580), .Z(n53581) );
  NOR U66074 ( .A(n56580), .B(n53581), .Z(n53582) );
  NOR U66075 ( .A(n53585), .B(n53582), .Z(n53583) );
  NOR U66076 ( .A(n53584), .B(n53583), .Z(n57081) );
  IV U66077 ( .A(n53584), .Z(n53586) );
  NOR U66078 ( .A(n53586), .B(n53585), .Z(n53587) );
  NOR U66079 ( .A(n57081), .B(n53587), .Z(n57100) );
  IV U66080 ( .A(n53588), .Z(n53589) );
  NOR U66081 ( .A(n53590), .B(n53589), .Z(n53595) );
  IV U66082 ( .A(n53591), .Z(n53592) );
  NOR U66083 ( .A(n53593), .B(n53592), .Z(n53594) );
  NOR U66084 ( .A(n53595), .B(n53594), .Z(n57102) );
  XOR U66085 ( .A(n57100), .B(n57102), .Z(n57110) );
  IV U66086 ( .A(n57110), .Z(n53603) );
  IV U66087 ( .A(n53596), .Z(n53597) );
  NOR U66088 ( .A(n53598), .B(n53597), .Z(n57104) );
  IV U66089 ( .A(n53599), .Z(n53601) );
  NOR U66090 ( .A(n53601), .B(n53600), .Z(n57109) );
  NOR U66091 ( .A(n57104), .B(n57109), .Z(n53602) );
  XOR U66092 ( .A(n53603), .B(n53602), .Z(n57114) );
  XOR U66093 ( .A(n57112), .B(n57114), .Z(n57116) );
  XOR U66094 ( .A(n57115), .B(n57116), .Z(n57087) );
  XOR U66095 ( .A(n57086), .B(n57087), .Z(n57091) );
  XOR U66096 ( .A(n57089), .B(n57091), .Z(n57085) );
  XOR U66097 ( .A(n57084), .B(n57085), .Z(n57138) );
  XOR U66098 ( .A(n57136), .B(n57138), .Z(n57130) );
  XOR U66099 ( .A(n53604), .B(n57130), .Z(n53605) );
  IV U66100 ( .A(n53605), .Z(n57127) );
  XOR U66101 ( .A(n57125), .B(n57127), .Z(n56558) );
  XOR U66102 ( .A(n56557), .B(n56558), .Z(n56561) );
  XOR U66103 ( .A(n56560), .B(n56561), .Z(n56543) );
  XOR U66104 ( .A(n56542), .B(n56543), .Z(n56545) );
  XOR U66105 ( .A(n56546), .B(n56545), .Z(n53606) );
  NOR U66106 ( .A(n53608), .B(n53606), .Z(n53613) );
  IV U66107 ( .A(n53613), .Z(n53607) );
  NOR U66108 ( .A(n53611), .B(n53607), .Z(n57151) );
  IV U66109 ( .A(n53608), .Z(n53609) );
  NOR U66110 ( .A(n56545), .B(n53609), .Z(n53610) );
  NOR U66111 ( .A(n53611), .B(n53610), .Z(n53612) );
  NOR U66112 ( .A(n53613), .B(n53612), .Z(n57154) );
  NOR U66113 ( .A(n57151), .B(n57154), .Z(n53620) );
  NOR U66114 ( .A(n53615), .B(n53614), .Z(n57150) );
  IV U66115 ( .A(n53616), .Z(n53618) );
  NOR U66116 ( .A(n53618), .B(n53617), .Z(n56570) );
  NOR U66117 ( .A(n57150), .B(n56570), .Z(n53619) );
  XOR U66118 ( .A(n53620), .B(n53619), .Z(n56573) );
  XOR U66119 ( .A(n56571), .B(n56573), .Z(n56565) );
  XOR U66120 ( .A(n56566), .B(n56565), .Z(n56541) );
  IV U66121 ( .A(n53621), .Z(n53622) );
  NOR U66122 ( .A(n53623), .B(n53622), .Z(n56568) );
  NOR U66123 ( .A(n53625), .B(n53624), .Z(n56539) );
  NOR U66124 ( .A(n56568), .B(n56539), .Z(n53626) );
  XOR U66125 ( .A(n56541), .B(n53626), .Z(n56550) );
  IV U66126 ( .A(n56550), .Z(n56551) );
  IV U66127 ( .A(n53629), .Z(n53627) );
  NOR U66128 ( .A(n53628), .B(n53627), .Z(n53635) );
  NOR U66129 ( .A(n53630), .B(n53629), .Z(n53633) );
  IV U66130 ( .A(n53631), .Z(n53632) );
  NOR U66131 ( .A(n53633), .B(n53632), .Z(n53634) );
  NOR U66132 ( .A(n53635), .B(n53634), .Z(n56552) );
  IV U66133 ( .A(n56552), .Z(n56549) );
  XOR U66134 ( .A(n56551), .B(n56549), .Z(n57163) );
  XOR U66135 ( .A(n57161), .B(n57163), .Z(n57166) );
  XOR U66136 ( .A(n57164), .B(n57166), .Z(n57172) );
  XOR U66137 ( .A(n53636), .B(n57172), .Z(n53637) );
  IV U66138 ( .A(n53637), .Z(n57208) );
  XOR U66139 ( .A(n57206), .B(n57208), .Z(n57176) );
  IV U66140 ( .A(n53638), .Z(n53639) );
  NOR U66141 ( .A(n53639), .B(n53641), .Z(n57174) );
  XOR U66142 ( .A(n57176), .B(n57174), .Z(n57179) );
  IV U66143 ( .A(n53640), .Z(n53642) );
  NOR U66144 ( .A(n53642), .B(n53641), .Z(n57177) );
  XOR U66145 ( .A(n57179), .B(n57177), .Z(n57196) );
  XOR U66146 ( .A(n57195), .B(n57196), .Z(n57198) );
  IV U66147 ( .A(n53643), .Z(n53645) );
  NOR U66148 ( .A(n53645), .B(n53644), .Z(n53647) );
  NOR U66149 ( .A(n53647), .B(n53646), .Z(n57199) );
  XOR U66150 ( .A(n57198), .B(n57199), .Z(n57209) );
  XOR U66151 ( .A(n57211), .B(n57209), .Z(n57189) );
  XOR U66152 ( .A(n57188), .B(n57189), .Z(n57191) );
  IV U66153 ( .A(n53648), .Z(n53650) );
  NOR U66154 ( .A(n53650), .B(n53649), .Z(n53651) );
  NOR U66155 ( .A(n53652), .B(n53651), .Z(n57192) );
  XOR U66156 ( .A(n57191), .B(n57192), .Z(n57217) );
  XOR U66157 ( .A(n57216), .B(n57217), .Z(n57229) );
  IV U66158 ( .A(n53653), .Z(n53654) );
  NOR U66159 ( .A(n53655), .B(n53654), .Z(n57221) );
  NOR U66160 ( .A(n53657), .B(n53656), .Z(n57230) );
  NOR U66161 ( .A(n57221), .B(n57230), .Z(n53658) );
  XOR U66162 ( .A(n57229), .B(n53658), .Z(n57228) );
  XOR U66163 ( .A(n57226), .B(n57228), .Z(n56531) );
  IV U66164 ( .A(n53659), .Z(n53661) );
  NOR U66165 ( .A(n53661), .B(n53660), .Z(n56529) );
  XOR U66166 ( .A(n56531), .B(n56529), .Z(n56534) );
  IV U66167 ( .A(n53662), .Z(n53664) );
  NOR U66168 ( .A(n53664), .B(n53663), .Z(n56532) );
  XOR U66169 ( .A(n56534), .B(n56532), .Z(n53671) );
  NOR U66170 ( .A(n53675), .B(n53671), .Z(n53670) );
  IV U66171 ( .A(n53665), .Z(n53666) );
  NOR U66172 ( .A(n53667), .B(n53666), .Z(n53672) );
  IV U66173 ( .A(n53672), .Z(n53668) );
  NOR U66174 ( .A(n56534), .B(n53668), .Z(n53669) );
  NOR U66175 ( .A(n53670), .B(n53669), .Z(n57242) );
  IV U66176 ( .A(n57242), .Z(n53674) );
  IV U66177 ( .A(n53671), .Z(n53676) );
  NOR U66178 ( .A(n53672), .B(n53676), .Z(n53673) );
  NOR U66179 ( .A(n53674), .B(n53673), .Z(n53678) );
  NOR U66180 ( .A(n53676), .B(n53675), .Z(n53677) );
  NOR U66181 ( .A(n53678), .B(n53677), .Z(n56538) );
  IV U66182 ( .A(n53679), .Z(n53681) );
  NOR U66183 ( .A(n53681), .B(n53680), .Z(n53686) );
  IV U66184 ( .A(n53682), .Z(n53684) );
  NOR U66185 ( .A(n53684), .B(n53683), .Z(n53685) );
  NOR U66186 ( .A(n53686), .B(n53685), .Z(n56537) );
  XOR U66187 ( .A(n56538), .B(n56537), .Z(n56521) );
  XOR U66188 ( .A(n56523), .B(n56521), .Z(n56525) );
  XOR U66189 ( .A(n56524), .B(n56525), .Z(n57254) );
  XOR U66190 ( .A(n53687), .B(n57254), .Z(n53688) );
  IV U66191 ( .A(n53688), .Z(n56514) );
  IV U66192 ( .A(n53689), .Z(n53691) );
  NOR U66193 ( .A(n53691), .B(n53690), .Z(n56513) );
  XOR U66194 ( .A(n56514), .B(n56513), .Z(n56510) );
  XOR U66195 ( .A(n56511), .B(n56510), .Z(n53692) );
  IV U66196 ( .A(n53692), .Z(n57246) );
  XOR U66197 ( .A(n57245), .B(n57246), .Z(n57250) );
  IV U66198 ( .A(n53693), .Z(n53695) );
  NOR U66199 ( .A(n53695), .B(n53694), .Z(n53696) );
  IV U66200 ( .A(n53696), .Z(n53697) );
  NOR U66201 ( .A(n53698), .B(n53697), .Z(n57248) );
  XOR U66202 ( .A(n57250), .B(n57248), .Z(n56501) );
  XOR U66203 ( .A(n56500), .B(n56501), .Z(n56504) );
  XOR U66204 ( .A(n56503), .B(n56504), .Z(n57277) );
  XOR U66205 ( .A(n57276), .B(n57277), .Z(n57281) );
  IV U66206 ( .A(n53699), .Z(n53701) );
  NOR U66207 ( .A(n53701), .B(n53700), .Z(n57279) );
  XOR U66208 ( .A(n57281), .B(n57279), .Z(n57269) );
  XOR U66209 ( .A(n57268), .B(n57269), .Z(n57272) );
  XOR U66210 ( .A(n57271), .B(n57272), .Z(n57291) );
  XOR U66211 ( .A(n57292), .B(n57291), .Z(n57287) );
  XOR U66212 ( .A(n53702), .B(n57287), .Z(n53708) );
  NOR U66213 ( .A(n53707), .B(n53708), .Z(n53712) );
  IV U66214 ( .A(n53712), .Z(n53706) );
  IV U66215 ( .A(n53703), .Z(n53705) );
  NOR U66216 ( .A(n53705), .B(n53704), .Z(n53711) );
  NOR U66217 ( .A(n53706), .B(n53711), .Z(n53717) );
  IV U66218 ( .A(n53707), .Z(n53710) );
  IV U66219 ( .A(n53708), .Z(n53709) );
  NOR U66220 ( .A(n53710), .B(n53709), .Z(n53715) );
  IV U66221 ( .A(n53711), .Z(n53713) );
  NOR U66222 ( .A(n53713), .B(n53712), .Z(n53714) );
  NOR U66223 ( .A(n53715), .B(n53714), .Z(n53716) );
  IV U66224 ( .A(n53716), .Z(n57306) );
  NOR U66225 ( .A(n53717), .B(n57306), .Z(n57303) );
  XOR U66226 ( .A(n57305), .B(n57303), .Z(n56494) );
  XOR U66227 ( .A(n56492), .B(n56494), .Z(n56491) );
  XOR U66228 ( .A(n56489), .B(n56491), .Z(n56487) );
  XOR U66229 ( .A(n56486), .B(n56487), .Z(n57316) );
  XOR U66230 ( .A(n57317), .B(n57316), .Z(n57325) );
  NOR U66231 ( .A(n53727), .B(n57325), .Z(n53726) );
  IV U66232 ( .A(n53718), .Z(n53720) );
  NOR U66233 ( .A(n53720), .B(n53719), .Z(n53725) );
  IV U66234 ( .A(n53721), .Z(n53723) );
  NOR U66235 ( .A(n53723), .B(n53722), .Z(n53724) );
  NOR U66236 ( .A(n53725), .B(n53724), .Z(n53729) );
  NOR U66237 ( .A(n53726), .B(n53729), .Z(n57328) );
  IV U66238 ( .A(n53727), .Z(n57327) );
  XOR U66239 ( .A(n57327), .B(n57325), .Z(n53728) );
  NOR U66240 ( .A(n57328), .B(n53728), .Z(n53731) );
  NOR U66241 ( .A(n57328), .B(n53729), .Z(n53730) );
  NOR U66242 ( .A(n53731), .B(n53730), .Z(n57320) );
  XOR U66243 ( .A(n57318), .B(n57320), .Z(n57321) );
  XOR U66244 ( .A(n57322), .B(n57321), .Z(n57345) );
  IV U66245 ( .A(n53732), .Z(n53733) );
  NOR U66246 ( .A(n53734), .B(n53733), .Z(n53738) );
  NOR U66247 ( .A(n53736), .B(n53735), .Z(n53737) );
  NOR U66248 ( .A(n53738), .B(n53737), .Z(n57347) );
  IV U66249 ( .A(n53739), .Z(n53740) );
  NOR U66250 ( .A(n53740), .B(n53745), .Z(n57338) );
  NOR U66251 ( .A(n57342), .B(n57338), .Z(n53748) );
  IV U66252 ( .A(n53741), .Z(n53743) );
  NOR U66253 ( .A(n53743), .B(n53742), .Z(n57343) );
  IV U66254 ( .A(n53744), .Z(n53746) );
  NOR U66255 ( .A(n53746), .B(n53745), .Z(n57339) );
  NOR U66256 ( .A(n57343), .B(n57339), .Z(n53747) );
  XOR U66257 ( .A(n53748), .B(n53747), .Z(n53749) );
  XOR U66258 ( .A(n57347), .B(n53749), .Z(n53750) );
  XOR U66259 ( .A(n57345), .B(n53750), .Z(n57340) );
  XOR U66260 ( .A(n57336), .B(n57340), .Z(n56484) );
  XOR U66261 ( .A(n53751), .B(n56484), .Z(n57369) );
  XOR U66262 ( .A(n57370), .B(n57369), .Z(n57374) );
  XOR U66263 ( .A(n57372), .B(n57374), .Z(n57359) );
  XOR U66264 ( .A(n57358), .B(n57359), .Z(n57363) );
  XOR U66265 ( .A(n57361), .B(n57363), .Z(n57365) );
  XOR U66266 ( .A(n57364), .B(n57365), .Z(n56478) );
  XOR U66267 ( .A(n56477), .B(n56478), .Z(n57389) );
  XOR U66268 ( .A(n53752), .B(n57389), .Z(n57391) );
  XOR U66269 ( .A(n57393), .B(n57391), .Z(n57434) );
  XOR U66270 ( .A(n57433), .B(n57434), .Z(n57432) );
  XOR U66271 ( .A(n57431), .B(n57432), .Z(n56459) );
  IV U66272 ( .A(n56459), .Z(n53757) );
  IV U66273 ( .A(n53753), .Z(n53755) );
  IV U66274 ( .A(n53754), .Z(n53759) );
  NOR U66275 ( .A(n53755), .B(n53759), .Z(n56457) );
  NOR U66276 ( .A(n57430), .B(n56457), .Z(n53756) );
  XOR U66277 ( .A(n53757), .B(n53756), .Z(n56463) );
  IV U66278 ( .A(n53758), .Z(n53760) );
  NOR U66279 ( .A(n53760), .B(n53759), .Z(n56461) );
  XOR U66280 ( .A(n56463), .B(n56461), .Z(n56456) );
  XOR U66281 ( .A(n56454), .B(n56456), .Z(n56471) );
  XOR U66282 ( .A(n56469), .B(n56471), .Z(n56473) );
  XOR U66283 ( .A(n56472), .B(n56473), .Z(n57406) );
  XOR U66284 ( .A(n57404), .B(n57406), .Z(n57418) );
  XOR U66285 ( .A(n57417), .B(n57418), .Z(n57420) );
  XOR U66286 ( .A(n57421), .B(n57420), .Z(n57407) );
  XOR U66287 ( .A(n57408), .B(n57407), .Z(n57440) );
  NOR U66288 ( .A(n53762), .B(n53761), .Z(n57441) );
  IV U66289 ( .A(n53763), .Z(n53764) );
  NOR U66290 ( .A(n53765), .B(n53764), .Z(n57411) );
  NOR U66291 ( .A(n57441), .B(n57411), .Z(n53766) );
  XOR U66292 ( .A(n57440), .B(n53766), .Z(n57439) );
  XOR U66293 ( .A(n57437), .B(n57439), .Z(n57429) );
  XOR U66294 ( .A(n57428), .B(n57429), .Z(n56448) );
  XOR U66295 ( .A(n56447), .B(n56448), .Z(n56450) );
  XOR U66296 ( .A(n56451), .B(n56450), .Z(n53767) );
  NOR U66297 ( .A(n53771), .B(n53767), .Z(n53775) );
  IV U66298 ( .A(n53768), .Z(n53770) );
  NOR U66299 ( .A(n53770), .B(n53769), .Z(n53777) );
  IV U66300 ( .A(n53771), .Z(n53772) );
  NOR U66301 ( .A(n56450), .B(n53772), .Z(n53773) );
  NOR U66302 ( .A(n53777), .B(n53773), .Z(n53774) );
  NOR U66303 ( .A(n53775), .B(n53774), .Z(n57451) );
  IV U66304 ( .A(n53775), .Z(n53776) );
  NOR U66305 ( .A(n53777), .B(n53776), .Z(n53778) );
  NOR U66306 ( .A(n57451), .B(n53778), .Z(n53779) );
  IV U66307 ( .A(n53779), .Z(n57448) );
  XOR U66308 ( .A(n57449), .B(n57448), .Z(n57469) );
  IV U66309 ( .A(n53780), .Z(n53782) );
  NOR U66310 ( .A(n53782), .B(n53781), .Z(n53784) );
  NOR U66311 ( .A(n53784), .B(n53783), .Z(n57471) );
  XOR U66312 ( .A(n57469), .B(n57471), .Z(n57473) );
  NOR U66313 ( .A(n53791), .B(n57473), .Z(n57479) );
  IV U66314 ( .A(n53785), .Z(n53786) );
  NOR U66315 ( .A(n53787), .B(n53786), .Z(n53788) );
  IV U66316 ( .A(n53788), .Z(n57454) );
  NOR U66317 ( .A(n53790), .B(n53789), .Z(n57472) );
  XOR U66318 ( .A(n57472), .B(n57473), .Z(n57453) );
  XOR U66319 ( .A(n57454), .B(n57453), .Z(n53794) );
  IV U66320 ( .A(n57453), .Z(n53792) );
  NOR U66321 ( .A(n53792), .B(n53791), .Z(n53793) );
  NOR U66322 ( .A(n53794), .B(n53793), .Z(n53795) );
  NOR U66323 ( .A(n57479), .B(n53795), .Z(n53806) );
  IV U66324 ( .A(n53806), .Z(n57456) );
  IV U66325 ( .A(n53796), .Z(n53797) );
  NOR U66326 ( .A(n53798), .B(n53797), .Z(n53805) );
  IV U66327 ( .A(n53799), .Z(n53800) );
  NOR U66328 ( .A(n53801), .B(n53800), .Z(n57455) );
  NOR U66329 ( .A(n53805), .B(n57455), .Z(n53802) );
  XOR U66330 ( .A(n57456), .B(n53802), .Z(n53803) );
  NOR U66331 ( .A(n53804), .B(n53803), .Z(n53809) );
  IV U66332 ( .A(n53804), .Z(n53808) );
  IV U66333 ( .A(n53805), .Z(n57452) );
  XOR U66334 ( .A(n57452), .B(n53806), .Z(n53807) );
  NOR U66335 ( .A(n53808), .B(n53807), .Z(n56413) );
  NOR U66336 ( .A(n53809), .B(n56413), .Z(n53810) );
  IV U66337 ( .A(n53810), .Z(n56410) );
  XOR U66338 ( .A(n56409), .B(n56410), .Z(n56417) );
  XOR U66339 ( .A(n56416), .B(n56417), .Z(n56421) );
  NOR U66340 ( .A(n53812), .B(n53811), .Z(n53813) );
  NOR U66341 ( .A(n53814), .B(n53813), .Z(n56419) );
  XOR U66342 ( .A(n56421), .B(n56419), .Z(n56404) );
  IV U66343 ( .A(n53815), .Z(n53816) );
  NOR U66344 ( .A(n53817), .B(n53816), .Z(n56402) );
  XOR U66345 ( .A(n56404), .B(n56402), .Z(n56405) );
  IV U66346 ( .A(n53818), .Z(n53820) );
  NOR U66347 ( .A(n53820), .B(n53819), .Z(n53825) );
  IV U66348 ( .A(n53821), .Z(n53822) );
  NOR U66349 ( .A(n53823), .B(n53822), .Z(n53824) );
  NOR U66350 ( .A(n53825), .B(n53824), .Z(n56406) );
  XOR U66351 ( .A(n56405), .B(n56406), .Z(n56427) );
  XOR U66352 ( .A(n56426), .B(n56427), .Z(n53830) );
  IV U66353 ( .A(n53826), .Z(n53827) );
  NOR U66354 ( .A(n53828), .B(n53827), .Z(n56431) );
  NOR U66355 ( .A(n56430), .B(n56431), .Z(n53829) );
  XOR U66356 ( .A(n53830), .B(n53829), .Z(n56439) );
  XOR U66357 ( .A(n56437), .B(n56439), .Z(n56398) );
  IV U66358 ( .A(n53831), .Z(n53832) );
  NOR U66359 ( .A(n53833), .B(n53832), .Z(n56436) );
  IV U66360 ( .A(n53834), .Z(n53835) );
  NOR U66361 ( .A(n53835), .B(n53839), .Z(n56397) );
  NOR U66362 ( .A(n56436), .B(n56397), .Z(n53836) );
  XOR U66363 ( .A(n56398), .B(n53836), .Z(n53837) );
  IV U66364 ( .A(n53837), .Z(n56445) );
  XOR U66365 ( .A(n56444), .B(n56445), .Z(n56391) );
  IV U66366 ( .A(n53838), .Z(n53840) );
  NOR U66367 ( .A(n53840), .B(n53839), .Z(n56389) );
  XOR U66368 ( .A(n56391), .B(n56389), .Z(n56393) );
  XOR U66369 ( .A(n56392), .B(n56393), .Z(n56373) );
  XOR U66370 ( .A(n56374), .B(n56373), .Z(n53844) );
  IV U66371 ( .A(n53841), .Z(n53847) );
  NOR U66372 ( .A(n53847), .B(n53842), .Z(n56376) );
  NOR U66373 ( .A(n56375), .B(n56376), .Z(n53843) );
  XOR U66374 ( .A(n53844), .B(n53843), .Z(n56383) );
  IV U66375 ( .A(n53845), .Z(n53846) );
  NOR U66376 ( .A(n53847), .B(n53846), .Z(n56381) );
  XOR U66377 ( .A(n56383), .B(n56381), .Z(n56385) );
  XOR U66378 ( .A(n56384), .B(n56385), .Z(n56364) );
  XOR U66379 ( .A(n56365), .B(n56364), .Z(n56366) );
  XOR U66380 ( .A(n56368), .B(n56366), .Z(n56362) );
  XOR U66381 ( .A(n56360), .B(n56362), .Z(n56349) );
  XOR U66382 ( .A(n53848), .B(n56349), .Z(n53849) );
  IV U66383 ( .A(n53849), .Z(n56354) );
  XOR U66384 ( .A(n56352), .B(n56354), .Z(n56346) );
  XOR U66385 ( .A(n56347), .B(n56346), .Z(n53852) );
  IV U66386 ( .A(n53852), .Z(n53850) );
  NOR U66387 ( .A(n53851), .B(n53850), .Z(n57501) );
  NOR U66388 ( .A(n53853), .B(n53852), .Z(n57499) );
  IV U66389 ( .A(n53854), .Z(n53858) );
  NOR U66390 ( .A(n53856), .B(n53855), .Z(n53857) );
  IV U66391 ( .A(n53857), .Z(n53864) );
  NOR U66392 ( .A(n53858), .B(n53864), .Z(n57498) );
  XOR U66393 ( .A(n57499), .B(n57498), .Z(n53859) );
  NOR U66394 ( .A(n57501), .B(n53859), .Z(n53874) );
  IV U66395 ( .A(n53874), .Z(n57512) );
  IV U66396 ( .A(n53860), .Z(n53861) );
  NOR U66397 ( .A(n53862), .B(n53861), .Z(n57509) );
  IV U66398 ( .A(n53863), .Z(n53865) );
  NOR U66399 ( .A(n53865), .B(n53864), .Z(n53873) );
  NOR U66400 ( .A(n57509), .B(n53873), .Z(n53866) );
  XOR U66401 ( .A(n57512), .B(n53866), .Z(n53877) );
  IV U66402 ( .A(n53877), .Z(n53867) );
  NOR U66403 ( .A(n53868), .B(n53867), .Z(n56334) );
  IV U66404 ( .A(n53869), .Z(n57504) );
  IV U66405 ( .A(n53870), .Z(n53872) );
  NOR U66406 ( .A(n53872), .B(n53871), .Z(n53878) );
  IV U66407 ( .A(n53878), .Z(n53876) );
  IV U66408 ( .A(n53873), .Z(n57511) );
  XOR U66409 ( .A(n57511), .B(n53874), .Z(n53875) );
  NOR U66410 ( .A(n53876), .B(n53875), .Z(n57506) );
  NOR U66411 ( .A(n53878), .B(n53877), .Z(n53879) );
  NOR U66412 ( .A(n57506), .B(n53879), .Z(n53880) );
  IV U66413 ( .A(n53880), .Z(n57503) );
  XOR U66414 ( .A(n57504), .B(n57503), .Z(n53881) );
  NOR U66415 ( .A(n53882), .B(n53881), .Z(n53883) );
  NOR U66416 ( .A(n56334), .B(n53883), .Z(n53884) );
  IV U66417 ( .A(n53884), .Z(n56332) );
  XOR U66418 ( .A(n56331), .B(n56332), .Z(n56329) );
  XOR U66419 ( .A(n56328), .B(n56329), .Z(n56322) );
  XOR U66420 ( .A(n56321), .B(n56322), .Z(n56340) );
  XOR U66421 ( .A(n53885), .B(n56340), .Z(n53886) );
  IV U66422 ( .A(n53886), .Z(n56316) );
  IV U66423 ( .A(n53887), .Z(n53889) );
  NOR U66424 ( .A(n53889), .B(n53888), .Z(n56314) );
  XOR U66425 ( .A(n56316), .B(n56314), .Z(n56317) );
  XOR U66426 ( .A(n56318), .B(n56317), .Z(n53890) );
  IV U66427 ( .A(n53890), .Z(n57531) );
  XOR U66428 ( .A(n57525), .B(n57531), .Z(n53898) );
  IV U66429 ( .A(n53891), .Z(n53893) );
  NOR U66430 ( .A(n53893), .B(n53892), .Z(n57527) );
  IV U66431 ( .A(n53894), .Z(n53896) );
  NOR U66432 ( .A(n53896), .B(n53895), .Z(n57528) );
  NOR U66433 ( .A(n57527), .B(n57528), .Z(n53897) );
  XOR U66434 ( .A(n53898), .B(n53897), .Z(n56290) );
  XOR U66435 ( .A(n56288), .B(n56290), .Z(n56292) );
  XOR U66436 ( .A(n56291), .B(n56292), .Z(n56287) );
  XOR U66437 ( .A(n56285), .B(n56287), .Z(n56306) );
  XOR U66438 ( .A(n56304), .B(n56306), .Z(n56302) );
  XOR U66439 ( .A(n56301), .B(n56302), .Z(n56278) );
  IV U66440 ( .A(n56278), .Z(n53906) );
  NOR U66441 ( .A(n53900), .B(n53899), .Z(n53910) );
  IV U66442 ( .A(n53910), .Z(n56279) );
  NOR U66443 ( .A(n53906), .B(n56279), .Z(n53912) );
  IV U66444 ( .A(n53901), .Z(n53902) );
  NOR U66445 ( .A(n53903), .B(n53902), .Z(n53905) );
  IV U66446 ( .A(n53905), .Z(n53904) );
  NOR U66447 ( .A(n53904), .B(n56302), .Z(n56307) );
  NOR U66448 ( .A(n53906), .B(n53905), .Z(n53907) );
  NOR U66449 ( .A(n56307), .B(n53907), .Z(n53908) );
  IV U66450 ( .A(n53908), .Z(n53909) );
  NOR U66451 ( .A(n53910), .B(n53909), .Z(n53911) );
  NOR U66452 ( .A(n53912), .B(n53911), .Z(n56282) );
  XOR U66453 ( .A(n56280), .B(n56282), .Z(n56269) );
  XOR U66454 ( .A(n56268), .B(n56269), .Z(n56272) );
  XOR U66455 ( .A(n56271), .B(n56272), .Z(n56276) );
  XOR U66456 ( .A(n56277), .B(n56276), .Z(n56261) );
  NOR U66457 ( .A(n53914), .B(n53913), .Z(n53916) );
  NOR U66458 ( .A(n53916), .B(n53915), .Z(n53917) );
  IV U66459 ( .A(n53917), .Z(n56262) );
  XOR U66460 ( .A(n56261), .B(n56262), .Z(n56264) );
  XOR U66461 ( .A(n56265), .B(n56264), .Z(n56236) );
  XOR U66462 ( .A(n56238), .B(n56236), .Z(n56240) );
  XOR U66463 ( .A(n56239), .B(n56240), .Z(n56244) );
  XOR U66464 ( .A(n56245), .B(n56244), .Z(n56256) );
  XOR U66465 ( .A(n53918), .B(n56256), .Z(n53919) );
  IV U66466 ( .A(n53919), .Z(n56253) );
  XOR U66467 ( .A(n56251), .B(n56253), .Z(n57558) );
  XOR U66468 ( .A(n57557), .B(n57558), .Z(n56228) );
  IV U66469 ( .A(n53920), .Z(n53921) );
  NOR U66470 ( .A(n53922), .B(n53921), .Z(n56226) );
  XOR U66471 ( .A(n56228), .B(n56226), .Z(n57561) );
  IV U66472 ( .A(n57561), .Z(n53930) );
  IV U66473 ( .A(n53923), .Z(n53924) );
  NOR U66474 ( .A(n53925), .B(n53924), .Z(n57560) );
  IV U66475 ( .A(n53926), .Z(n53928) );
  NOR U66476 ( .A(n53928), .B(n53927), .Z(n56229) );
  NOR U66477 ( .A(n57560), .B(n56229), .Z(n53929) );
  XOR U66478 ( .A(n53930), .B(n53929), .Z(n57550) );
  XOR U66479 ( .A(n57549), .B(n57550), .Z(n57553) );
  XOR U66480 ( .A(n57552), .B(n57553), .Z(n56220) );
  IV U66481 ( .A(n53931), .Z(n53932) );
  NOR U66482 ( .A(n53933), .B(n53932), .Z(n56219) );
  IV U66483 ( .A(n53934), .Z(n53935) );
  NOR U66484 ( .A(n53936), .B(n53935), .Z(n56217) );
  NOR U66485 ( .A(n56219), .B(n56217), .Z(n53937) );
  XOR U66486 ( .A(n56220), .B(n53937), .Z(n53938) );
  NOR U66487 ( .A(n53943), .B(n53938), .Z(n53946) );
  IV U66488 ( .A(n53939), .Z(n53941) );
  NOR U66489 ( .A(n53941), .B(n53940), .Z(n53948) );
  IV U66490 ( .A(n53948), .Z(n53942) );
  NOR U66491 ( .A(n53946), .B(n53942), .Z(n56215) );
  IV U66492 ( .A(n53943), .Z(n53945) );
  XOR U66493 ( .A(n56219), .B(n56220), .Z(n53944) );
  NOR U66494 ( .A(n53945), .B(n53944), .Z(n56216) );
  NOR U66495 ( .A(n53946), .B(n56216), .Z(n53947) );
  NOR U66496 ( .A(n53948), .B(n53947), .Z(n53949) );
  NOR U66497 ( .A(n56215), .B(n53949), .Z(n56234) );
  IV U66498 ( .A(n53950), .Z(n53951) );
  NOR U66499 ( .A(n53952), .B(n53951), .Z(n56233) );
  NOR U66500 ( .A(n53954), .B(n53953), .Z(n57586) );
  NOR U66501 ( .A(n56233), .B(n57586), .Z(n53955) );
  XOR U66502 ( .A(n56234), .B(n53955), .Z(n57591) );
  XOR U66503 ( .A(n57589), .B(n57591), .Z(n56208) );
  XOR U66504 ( .A(n56207), .B(n56208), .Z(n56211) );
  XOR U66505 ( .A(n56210), .B(n56211), .Z(n57579) );
  XOR U66506 ( .A(n57580), .B(n57579), .Z(n53956) );
  IV U66507 ( .A(n53956), .Z(n57582) );
  XOR U66508 ( .A(n57581), .B(n57582), .Z(n56200) );
  XOR U66509 ( .A(n56199), .B(n56200), .Z(n56204) );
  IV U66510 ( .A(n53957), .Z(n53961) );
  NOR U66511 ( .A(n53959), .B(n53958), .Z(n53960) );
  IV U66512 ( .A(n53960), .Z(n53963) );
  NOR U66513 ( .A(n53961), .B(n53963), .Z(n56202) );
  XOR U66514 ( .A(n56204), .B(n56202), .Z(n57613) );
  IV U66515 ( .A(n57613), .Z(n57611) );
  IV U66516 ( .A(n53962), .Z(n53964) );
  NOR U66517 ( .A(n53964), .B(n53963), .Z(n57610) );
  IV U66518 ( .A(n57610), .Z(n57612) );
  XOR U66519 ( .A(n57611), .B(n57612), .Z(n57605) );
  IV U66520 ( .A(n57605), .Z(n53969) );
  IV U66521 ( .A(n53965), .Z(n53967) );
  NOR U66522 ( .A(n53967), .B(n53966), .Z(n57614) );
  NOR U66523 ( .A(n57603), .B(n57614), .Z(n53968) );
  XOR U66524 ( .A(n53969), .B(n53968), .Z(n57602) );
  XOR U66525 ( .A(n57600), .B(n57602), .Z(n56197) );
  XOR U66526 ( .A(n56198), .B(n56197), .Z(n56190) );
  NOR U66527 ( .A(n53971), .B(n53970), .Z(n53977) );
  NOR U66528 ( .A(n53973), .B(n53972), .Z(n53975) );
  NOR U66529 ( .A(n53975), .B(n53974), .Z(n53976) );
  NOR U66530 ( .A(n53977), .B(n53976), .Z(n53978) );
  IV U66531 ( .A(n53978), .Z(n56191) );
  XOR U66532 ( .A(n56190), .B(n56191), .Z(n56193) );
  XOR U66533 ( .A(n56194), .B(n56193), .Z(n56187) );
  XOR U66534 ( .A(n56189), .B(n56187), .Z(n56164) );
  IV U66535 ( .A(n56164), .Z(n56168) );
  IV U66536 ( .A(n53979), .Z(n53982) );
  IV U66537 ( .A(n53980), .Z(n53981) );
  NOR U66538 ( .A(n53982), .B(n53981), .Z(n56167) );
  IV U66539 ( .A(n56167), .Z(n56163) );
  XOR U66540 ( .A(n56168), .B(n56163), .Z(n56175) );
  IV U66541 ( .A(n53983), .Z(n53984) );
  NOR U66542 ( .A(n53985), .B(n53984), .Z(n56166) );
  IV U66543 ( .A(n53986), .Z(n53988) );
  NOR U66544 ( .A(n53988), .B(n53987), .Z(n56174) );
  NOR U66545 ( .A(n56166), .B(n56174), .Z(n53989) );
  XOR U66546 ( .A(n56175), .B(n53989), .Z(n56171) );
  XOR U66547 ( .A(n56173), .B(n56171), .Z(n56180) );
  NOR U66548 ( .A(n53991), .B(n53990), .Z(n53993) );
  NOR U66549 ( .A(n53993), .B(n53992), .Z(n56179) );
  XOR U66550 ( .A(n56180), .B(n56179), .Z(n56183) );
  XOR U66551 ( .A(n56182), .B(n56183), .Z(n57642) );
  IV U66552 ( .A(n53994), .Z(n53995) );
  NOR U66553 ( .A(n53996), .B(n53995), .Z(n57640) );
  XOR U66554 ( .A(n57642), .B(n57640), .Z(n57648) );
  XOR U66555 ( .A(n57647), .B(n57648), .Z(n57645) );
  NOR U66556 ( .A(n53998), .B(n53997), .Z(n54003) );
  NOR U66557 ( .A(n54000), .B(n53999), .Z(n54001) );
  IV U66558 ( .A(n54001), .Z(n54002) );
  NOR U66559 ( .A(n54003), .B(n54002), .Z(n57643) );
  XOR U66560 ( .A(n57645), .B(n57643), .Z(n57635) );
  XOR U66561 ( .A(n57632), .B(n57635), .Z(n56157) );
  IV U66562 ( .A(n54004), .Z(n54005) );
  NOR U66563 ( .A(n54006), .B(n54005), .Z(n57634) );
  NOR U66564 ( .A(n54008), .B(n54007), .Z(n56158) );
  NOR U66565 ( .A(n57634), .B(n56158), .Z(n54009) );
  XOR U66566 ( .A(n56157), .B(n54009), .Z(n56156) );
  XOR U66567 ( .A(n56154), .B(n56156), .Z(n57668) );
  IV U66568 ( .A(n57668), .Z(n54017) );
  NOR U66569 ( .A(n54011), .B(n54010), .Z(n54021) );
  IV U66570 ( .A(n54021), .Z(n57669) );
  NOR U66571 ( .A(n54017), .B(n57669), .Z(n54023) );
  IV U66572 ( .A(n54012), .Z(n54013) );
  NOR U66573 ( .A(n54014), .B(n54013), .Z(n54016) );
  IV U66574 ( .A(n54016), .Z(n54015) );
  NOR U66575 ( .A(n56156), .B(n54015), .Z(n57670) );
  NOR U66576 ( .A(n54017), .B(n54016), .Z(n54018) );
  NOR U66577 ( .A(n57670), .B(n54018), .Z(n54019) );
  IV U66578 ( .A(n54019), .Z(n54020) );
  NOR U66579 ( .A(n54021), .B(n54020), .Z(n54022) );
  NOR U66580 ( .A(n54023), .B(n54022), .Z(n57663) );
  XOR U66581 ( .A(n57661), .B(n57663), .Z(n57664) );
  XOR U66582 ( .A(n57665), .B(n57664), .Z(n57678) );
  XOR U66583 ( .A(n57674), .B(n57678), .Z(n57694) );
  NOR U66584 ( .A(n54025), .B(n54024), .Z(n57676) );
  NOR U66585 ( .A(n54027), .B(n54026), .Z(n57692) );
  NOR U66586 ( .A(n57676), .B(n57692), .Z(n54028) );
  XOR U66587 ( .A(n57694), .B(n54028), .Z(n57689) );
  XOR U66588 ( .A(n57690), .B(n57689), .Z(n56141) );
  XOR U66589 ( .A(n56140), .B(n56141), .Z(n56143) );
  XOR U66590 ( .A(n56144), .B(n56143), .Z(n54029) );
  IV U66591 ( .A(n54029), .Z(n56148) );
  XOR U66592 ( .A(n56147), .B(n56148), .Z(n56150) );
  IV U66593 ( .A(n56150), .Z(n54034) );
  NOR U66594 ( .A(n54031), .B(n54030), .Z(n54032) );
  NOR U66595 ( .A(n54033), .B(n54032), .Z(n56151) );
  XOR U66596 ( .A(n54034), .B(n56151), .Z(n57708) );
  XOR U66597 ( .A(n57705), .B(n57708), .Z(n54035) );
  NOR U66598 ( .A(n54036), .B(n54035), .Z(n57704) );
  IV U66599 ( .A(n54037), .Z(n54038) );
  NOR U66600 ( .A(n54039), .B(n54038), .Z(n57707) );
  NOR U66601 ( .A(n57705), .B(n57707), .Z(n54040) );
  XOR U66602 ( .A(n54040), .B(n57708), .Z(n54045) );
  NOR U66603 ( .A(n54041), .B(n54045), .Z(n54042) );
  NOR U66604 ( .A(n57704), .B(n54042), .Z(n54043) );
  NOR U66605 ( .A(n54044), .B(n54043), .Z(n57702) );
  IV U66606 ( .A(n54044), .Z(n54047) );
  IV U66607 ( .A(n54045), .Z(n54046) );
  NOR U66608 ( .A(n54047), .B(n54046), .Z(n57699) );
  NOR U66609 ( .A(n57702), .B(n57699), .Z(n57718) );
  XOR U66610 ( .A(n54048), .B(n57718), .Z(n56135) );
  XOR U66611 ( .A(n56133), .B(n56135), .Z(n57722) );
  XOR U66612 ( .A(n57723), .B(n57722), .Z(n56110) );
  XOR U66613 ( .A(n56112), .B(n56110), .Z(n56114) );
  XOR U66614 ( .A(n56113), .B(n56114), .Z(n56108) );
  XOR U66615 ( .A(n56107), .B(n56108), .Z(n56119) );
  XOR U66616 ( .A(n56118), .B(n56119), .Z(n56125) );
  XOR U66617 ( .A(n56124), .B(n56125), .Z(n56122) );
  XOR U66618 ( .A(n56121), .B(n56122), .Z(n54051) );
  IV U66619 ( .A(n54051), .Z(n54049) );
  NOR U66620 ( .A(n54050), .B(n54049), .Z(n56105) );
  NOR U66621 ( .A(n54052), .B(n54051), .Z(n56103) );
  IV U66622 ( .A(n54053), .Z(n54054) );
  NOR U66623 ( .A(n54055), .B(n54054), .Z(n56102) );
  XOR U66624 ( .A(n56103), .B(n56102), .Z(n54056) );
  NOR U66625 ( .A(n56105), .B(n54056), .Z(n57748) );
  XOR U66626 ( .A(n57750), .B(n57748), .Z(n57753) );
  XOR U66627 ( .A(n57751), .B(n57753), .Z(n57757) );
  XOR U66628 ( .A(n57756), .B(n57757), .Z(n57764) );
  XOR U66629 ( .A(n57763), .B(n57764), .Z(n57760) );
  XOR U66630 ( .A(n57759), .B(n57760), .Z(n54057) );
  NOR U66631 ( .A(n54058), .B(n54057), .Z(n57804) );
  IV U66632 ( .A(n54059), .Z(n54061) );
  NOR U66633 ( .A(n54061), .B(n54060), .Z(n57741) );
  NOR U66634 ( .A(n57759), .B(n57741), .Z(n54062) );
  XOR U66635 ( .A(n57760), .B(n54062), .Z(n54063) );
  NOR U66636 ( .A(n54064), .B(n54063), .Z(n54068) );
  NOR U66637 ( .A(n57804), .B(n54068), .Z(n54065) );
  NOR U66638 ( .A(n54066), .B(n54065), .Z(n54069) );
  IV U66639 ( .A(n54066), .Z(n54067) );
  NOR U66640 ( .A(n54068), .B(n54067), .Z(n57803) );
  NOR U66641 ( .A(n54069), .B(n57803), .Z(n57743) );
  XOR U66642 ( .A(n57745), .B(n57743), .Z(n57782) );
  NOR U66643 ( .A(n54070), .B(n57782), .Z(n57784) );
  NOR U66644 ( .A(n54072), .B(n54071), .Z(n57781) );
  XOR U66645 ( .A(n57781), .B(n57782), .Z(n54085) );
  IV U66646 ( .A(n54085), .Z(n54073) );
  NOR U66647 ( .A(n54074), .B(n54073), .Z(n54075) );
  NOR U66648 ( .A(n57784), .B(n54075), .Z(n54076) );
  NOR U66649 ( .A(n54083), .B(n54076), .Z(n54086) );
  IV U66650 ( .A(n54077), .Z(n54081) );
  NOR U66651 ( .A(n54079), .B(n54078), .Z(n54080) );
  IV U66652 ( .A(n54080), .Z(n54092) );
  NOR U66653 ( .A(n54081), .B(n54092), .Z(n54088) );
  IV U66654 ( .A(n54088), .Z(n54082) );
  NOR U66655 ( .A(n54086), .B(n54082), .Z(n57779) );
  IV U66656 ( .A(n54083), .Z(n54084) );
  NOR U66657 ( .A(n54085), .B(n54084), .Z(n57780) );
  NOR U66658 ( .A(n57780), .B(n54086), .Z(n54087) );
  NOR U66659 ( .A(n54088), .B(n54087), .Z(n54089) );
  NOR U66660 ( .A(n57779), .B(n54089), .Z(n56094) );
  IV U66661 ( .A(n54097), .Z(n54104) );
  IV U66662 ( .A(n54090), .Z(n54098) );
  NOR U66663 ( .A(n54104), .B(n54098), .Z(n54095) );
  IV U66664 ( .A(n54091), .Z(n54093) );
  NOR U66665 ( .A(n54093), .B(n54092), .Z(n54094) );
  NOR U66666 ( .A(n54095), .B(n54094), .Z(n57778) );
  IV U66667 ( .A(n54096), .Z(n54100) );
  XOR U66668 ( .A(n54098), .B(n54097), .Z(n54099) );
  NOR U66669 ( .A(n54100), .B(n54099), .Z(n56099) );
  XOR U66670 ( .A(n57778), .B(n56099), .Z(n54101) );
  XOR U66671 ( .A(n56094), .B(n54101), .Z(n54105) );
  IV U66672 ( .A(n54102), .Z(n54103) );
  NOR U66673 ( .A(n54104), .B(n54103), .Z(n56096) );
  NOR U66674 ( .A(n54105), .B(n56096), .Z(n54109) );
  IV U66675 ( .A(n56096), .Z(n56097) );
  NOR U66676 ( .A(n56094), .B(n56099), .Z(n54106) );
  IV U66677 ( .A(n54106), .Z(n54107) );
  NOR U66678 ( .A(n56097), .B(n54107), .Z(n54108) );
  NOR U66679 ( .A(n54109), .B(n54108), .Z(n57794) );
  IV U66680 ( .A(n54110), .Z(n54111) );
  NOR U66681 ( .A(n54112), .B(n54111), .Z(n57797) );
  IV U66682 ( .A(n54113), .Z(n54115) );
  NOR U66683 ( .A(n54115), .B(n54114), .Z(n57793) );
  XOR U66684 ( .A(n57797), .B(n57793), .Z(n54116) );
  XOR U66685 ( .A(n57794), .B(n54116), .Z(n57811) );
  XOR U66686 ( .A(n54117), .B(n57811), .Z(n57821) );
  NOR U66687 ( .A(n54119), .B(n54118), .Z(n54121) );
  NOR U66688 ( .A(n54121), .B(n54120), .Z(n54122) );
  IV U66689 ( .A(n54122), .Z(n57822) );
  XOR U66690 ( .A(n57821), .B(n57822), .Z(n54131) );
  IV U66691 ( .A(n54131), .Z(n54123) );
  NOR U66692 ( .A(n54130), .B(n54123), .Z(n54128) );
  IV U66693 ( .A(n54128), .Z(n54126) );
  NOR U66694 ( .A(n54125), .B(n54124), .Z(n54127) );
  NOR U66695 ( .A(n54126), .B(n54127), .Z(n54136) );
  IV U66696 ( .A(n54127), .Z(n54129) );
  NOR U66697 ( .A(n54129), .B(n54128), .Z(n54134) );
  IV U66698 ( .A(n54130), .Z(n54132) );
  NOR U66699 ( .A(n54132), .B(n54131), .Z(n54133) );
  NOR U66700 ( .A(n54134), .B(n54133), .Z(n54135) );
  IV U66701 ( .A(n54135), .Z(n57824) );
  NOR U66702 ( .A(n54136), .B(n57824), .Z(n57818) );
  NOR U66703 ( .A(n54138), .B(n54137), .Z(n57820) );
  XOR U66704 ( .A(n57818), .B(n57820), .Z(n56087) );
  XOR U66705 ( .A(n56086), .B(n56087), .Z(n56090) );
  XOR U66706 ( .A(n56089), .B(n56090), .Z(n56079) );
  XOR U66707 ( .A(n56078), .B(n56079), .Z(n56082) );
  XOR U66708 ( .A(n56081), .B(n56082), .Z(n56049) );
  XOR U66709 ( .A(n56047), .B(n56049), .Z(n56050) );
  XOR U66710 ( .A(n56051), .B(n56050), .Z(n54139) );
  IV U66711 ( .A(n54139), .Z(n56041) );
  XOR U66712 ( .A(n56041), .B(n56040), .Z(n56043) );
  XOR U66713 ( .A(n56044), .B(n56043), .Z(n56063) );
  IV U66714 ( .A(n54140), .Z(n54142) );
  NOR U66715 ( .A(n54142), .B(n54141), .Z(n54143) );
  IV U66716 ( .A(n54143), .Z(n56064) );
  XOR U66717 ( .A(n56063), .B(n56064), .Z(n56067) );
  XOR U66718 ( .A(n56066), .B(n56067), .Z(n56056) );
  IV U66719 ( .A(n56056), .Z(n54152) );
  IV U66720 ( .A(n54144), .Z(n54145) );
  NOR U66721 ( .A(n54146), .B(n54145), .Z(n54151) );
  IV U66722 ( .A(n54147), .Z(n54148) );
  NOR U66723 ( .A(n54149), .B(n54148), .Z(n54150) );
  NOR U66724 ( .A(n54151), .B(n54150), .Z(n56057) );
  XOR U66725 ( .A(n54152), .B(n56057), .Z(n56059) );
  XOR U66726 ( .A(n56058), .B(n56059), .Z(n56076) );
  XOR U66727 ( .A(n56075), .B(n56076), .Z(n56029) );
  XOR U66728 ( .A(n56028), .B(n56029), .Z(n56031) );
  XOR U66729 ( .A(n56032), .B(n56031), .Z(n54153) );
  IV U66730 ( .A(n54153), .Z(n56038) );
  XOR U66731 ( .A(n56037), .B(n56038), .Z(n56021) );
  XOR U66732 ( .A(n56020), .B(n56021), .Z(n56024) );
  XOR U66733 ( .A(n56023), .B(n56024), .Z(n56008) );
  XOR U66734 ( .A(n56007), .B(n56008), .Z(n56011) );
  XOR U66735 ( .A(n56010), .B(n56011), .Z(n56015) );
  IV U66736 ( .A(n54154), .Z(n54157) );
  IV U66737 ( .A(n54155), .Z(n54156) );
  NOR U66738 ( .A(n54157), .B(n54156), .Z(n56013) );
  XOR U66739 ( .A(n56015), .B(n56013), .Z(n56018) );
  XOR U66740 ( .A(n56019), .B(n56018), .Z(n57858) );
  XOR U66741 ( .A(n57856), .B(n57858), .Z(n57851) );
  IV U66742 ( .A(n54158), .Z(n54159) );
  NOR U66743 ( .A(n54160), .B(n54159), .Z(n57855) );
  NOR U66744 ( .A(n54162), .B(n54161), .Z(n57849) );
  NOR U66745 ( .A(n57855), .B(n57849), .Z(n54163) );
  XOR U66746 ( .A(n57851), .B(n54163), .Z(n57846) );
  IV U66747 ( .A(n54166), .Z(n54164) );
  NOR U66748 ( .A(n54165), .B(n54164), .Z(n54175) );
  NOR U66749 ( .A(n54167), .B(n54166), .Z(n54173) );
  IV U66750 ( .A(n54168), .Z(n54169) );
  NOR U66751 ( .A(n54170), .B(n54169), .Z(n54171) );
  IV U66752 ( .A(n54171), .Z(n54172) );
  NOR U66753 ( .A(n54173), .B(n54172), .Z(n54174) );
  NOR U66754 ( .A(n54175), .B(n54174), .Z(n57847) );
  XOR U66755 ( .A(n57846), .B(n57847), .Z(n57866) );
  XOR U66756 ( .A(n57865), .B(n57866), .Z(n57869) );
  XOR U66757 ( .A(n57868), .B(n57869), .Z(n55973) );
  XOR U66758 ( .A(n55972), .B(n55973), .Z(n54179) );
  NOR U66759 ( .A(n54177), .B(n54176), .Z(n55977) );
  NOR U66760 ( .A(n55976), .B(n55977), .Z(n54178) );
  XOR U66761 ( .A(n54179), .B(n54178), .Z(n55985) );
  XOR U66762 ( .A(n55983), .B(n55985), .Z(n55988) );
  XOR U66763 ( .A(n55986), .B(n55988), .Z(n55995) );
  XOR U66764 ( .A(n54180), .B(n55995), .Z(n54181) );
  IV U66765 ( .A(n54181), .Z(n55968) );
  XOR U66766 ( .A(n55967), .B(n55968), .Z(n55996) );
  XOR U66767 ( .A(n55997), .B(n55996), .Z(n55998) );
  NOR U66768 ( .A(n54183), .B(n54182), .Z(n54184) );
  NOR U66769 ( .A(n54185), .B(n54184), .Z(n56000) );
  XOR U66770 ( .A(n55998), .B(n56000), .Z(n57880) );
  NOR U66771 ( .A(n54186), .B(n57880), .Z(n57883) );
  XOR U66772 ( .A(n57879), .B(n57880), .Z(n57887) );
  IV U66773 ( .A(n57887), .Z(n54187) );
  NOR U66774 ( .A(n54188), .B(n54187), .Z(n54189) );
  NOR U66775 ( .A(n57883), .B(n54189), .Z(n55961) );
  NOR U66776 ( .A(n57884), .B(n55961), .Z(n54192) );
  IV U66777 ( .A(n57884), .Z(n54190) );
  NOR U66778 ( .A(n57887), .B(n54190), .Z(n54191) );
  NOR U66779 ( .A(n54192), .B(n54191), .Z(n54200) );
  IV U66780 ( .A(n54193), .Z(n54195) );
  NOR U66781 ( .A(n54195), .B(n54194), .Z(n57885) );
  IV U66782 ( .A(n54196), .Z(n54198) );
  NOR U66783 ( .A(n54198), .B(n54197), .Z(n55962) );
  NOR U66784 ( .A(n57885), .B(n55962), .Z(n54199) );
  XOR U66785 ( .A(n54200), .B(n54199), .Z(n57902) );
  XOR U66786 ( .A(n57903), .B(n57902), .Z(n57904) );
  IV U66787 ( .A(n54201), .Z(n54206) );
  IV U66788 ( .A(n54202), .Z(n54203) );
  NOR U66789 ( .A(n54203), .B(n54209), .Z(n54204) );
  IV U66790 ( .A(n54204), .Z(n54205) );
  NOR U66791 ( .A(n54206), .B(n54205), .Z(n54207) );
  IV U66792 ( .A(n54207), .Z(n57905) );
  XOR U66793 ( .A(n57904), .B(n57905), .Z(n57896) );
  IV U66794 ( .A(n54208), .Z(n54210) );
  NOR U66795 ( .A(n54210), .B(n54209), .Z(n57894) );
  XOR U66796 ( .A(n57896), .B(n57894), .Z(n57898) );
  XOR U66797 ( .A(n57897), .B(n57898), .Z(n55959) );
  XOR U66798 ( .A(n55958), .B(n55959), .Z(n55930) );
  XOR U66799 ( .A(n55929), .B(n55930), .Z(n55934) );
  IV U66800 ( .A(n54211), .Z(n54212) );
  NOR U66801 ( .A(n54213), .B(n54212), .Z(n55932) );
  XOR U66802 ( .A(n55934), .B(n55932), .Z(n55919) );
  XOR U66803 ( .A(n55918), .B(n55919), .Z(n55923) );
  IV U66804 ( .A(n54214), .Z(n54217) );
  IV U66805 ( .A(n54215), .Z(n54216) );
  NOR U66806 ( .A(n54217), .B(n54216), .Z(n55921) );
  XOR U66807 ( .A(n55923), .B(n55921), .Z(n55926) );
  IV U66808 ( .A(n54218), .Z(n54219) );
  NOR U66809 ( .A(n54236), .B(n54219), .Z(n54220) );
  IV U66810 ( .A(n54220), .Z(n54226) );
  IV U66811 ( .A(n54221), .Z(n54223) );
  NOR U66812 ( .A(n54223), .B(n54222), .Z(n54224) );
  IV U66813 ( .A(n54224), .Z(n54225) );
  NOR U66814 ( .A(n54226), .B(n54225), .Z(n55924) );
  XOR U66815 ( .A(n55926), .B(n55924), .Z(n54244) );
  IV U66816 ( .A(n54244), .Z(n54233) );
  IV U66817 ( .A(n54227), .Z(n54232) );
  IV U66818 ( .A(n54228), .Z(n54229) );
  NOR U66819 ( .A(n54229), .B(n54236), .Z(n54230) );
  IV U66820 ( .A(n54230), .Z(n54231) );
  NOR U66821 ( .A(n54232), .B(n54231), .Z(n54242) );
  NOR U66822 ( .A(n54233), .B(n54242), .Z(n54240) );
  IV U66823 ( .A(n54240), .Z(n54234) );
  NOR U66824 ( .A(n54239), .B(n54234), .Z(n54248) );
  IV U66825 ( .A(n54235), .Z(n54237) );
  NOR U66826 ( .A(n54237), .B(n54236), .Z(n54250) );
  IV U66827 ( .A(n54250), .Z(n54238) );
  NOR U66828 ( .A(n54248), .B(n54238), .Z(n55915) );
  IV U66829 ( .A(n54239), .Z(n54241) );
  NOR U66830 ( .A(n54241), .B(n54240), .Z(n54246) );
  IV U66831 ( .A(n54242), .Z(n54243) );
  NOR U66832 ( .A(n54244), .B(n54243), .Z(n54245) );
  NOR U66833 ( .A(n54246), .B(n54245), .Z(n54247) );
  IV U66834 ( .A(n54247), .Z(n55914) );
  NOR U66835 ( .A(n54248), .B(n55914), .Z(n54249) );
  NOR U66836 ( .A(n54250), .B(n54249), .Z(n54251) );
  NOR U66837 ( .A(n55915), .B(n54251), .Z(n54252) );
  IV U66838 ( .A(n54252), .Z(n55947) );
  XOR U66839 ( .A(n55946), .B(n55947), .Z(n55951) );
  IV U66840 ( .A(n54253), .Z(n54255) );
  NOR U66841 ( .A(n54255), .B(n54254), .Z(n55949) );
  XOR U66842 ( .A(n55951), .B(n55949), .Z(n54265) );
  IV U66843 ( .A(n54265), .Z(n54260) );
  NOR U66844 ( .A(n54257), .B(n54256), .Z(n54259) );
  NOR U66845 ( .A(n54259), .B(n54258), .Z(n54264) );
  NOR U66846 ( .A(n54260), .B(n54264), .Z(n54269) );
  IV U66847 ( .A(n54261), .Z(n54262) );
  NOR U66848 ( .A(n54263), .B(n54262), .Z(n54271) );
  IV U66849 ( .A(n54264), .Z(n54266) );
  NOR U66850 ( .A(n54266), .B(n54265), .Z(n54267) );
  NOR U66851 ( .A(n54271), .B(n54267), .Z(n54268) );
  NOR U66852 ( .A(n54269), .B(n54268), .Z(n55945) );
  IV U66853 ( .A(n54269), .Z(n54270) );
  NOR U66854 ( .A(n54271), .B(n54270), .Z(n54272) );
  NOR U66855 ( .A(n55945), .B(n54272), .Z(n54273) );
  IV U66856 ( .A(n54273), .Z(n55942) );
  XOR U66857 ( .A(n55941), .B(n55942), .Z(n55906) );
  XOR U66858 ( .A(n55905), .B(n55906), .Z(n55908) );
  IV U66859 ( .A(n55908), .Z(n54282) );
  IV U66860 ( .A(n54274), .Z(n54275) );
  NOR U66861 ( .A(n54276), .B(n54275), .Z(n54281) );
  IV U66862 ( .A(n54277), .Z(n54278) );
  NOR U66863 ( .A(n54279), .B(n54278), .Z(n54280) );
  NOR U66864 ( .A(n54281), .B(n54280), .Z(n55909) );
  XOR U66865 ( .A(n54282), .B(n55909), .Z(n55899) );
  XOR U66866 ( .A(n55897), .B(n55899), .Z(n55901) );
  XOR U66867 ( .A(n55900), .B(n55901), .Z(n55916) );
  XOR U66868 ( .A(n55917), .B(n55916), .Z(n54289) );
  IV U66869 ( .A(n54289), .Z(n54287) );
  IV U66870 ( .A(n54283), .Z(n54284) );
  NOR U66871 ( .A(n54285), .B(n54284), .Z(n54288) );
  IV U66872 ( .A(n54288), .Z(n54286) );
  NOR U66873 ( .A(n54287), .B(n54286), .Z(n57928) );
  NOR U66874 ( .A(n54289), .B(n54288), .Z(n57926) );
  IV U66875 ( .A(n54290), .Z(n54293) );
  IV U66876 ( .A(n54291), .Z(n54292) );
  NOR U66877 ( .A(n54293), .B(n54292), .Z(n57925) );
  XOR U66878 ( .A(n57926), .B(n57925), .Z(n54294) );
  NOR U66879 ( .A(n57928), .B(n54294), .Z(n54295) );
  IV U66880 ( .A(n54295), .Z(n57937) );
  XOR U66881 ( .A(n57936), .B(n57937), .Z(n57934) );
  XOR U66882 ( .A(n57933), .B(n57934), .Z(n57931) );
  XOR U66883 ( .A(n57930), .B(n57931), .Z(n57947) );
  XOR U66884 ( .A(n57946), .B(n57947), .Z(n57950) );
  XOR U66885 ( .A(n57949), .B(n57950), .Z(n57963) );
  XOR U66886 ( .A(n57962), .B(n57963), .Z(n57966) );
  XOR U66887 ( .A(n57965), .B(n57966), .Z(n55890) );
  IV U66888 ( .A(n55890), .Z(n54304) );
  IV U66889 ( .A(n54296), .Z(n54297) );
  NOR U66890 ( .A(n54298), .B(n54297), .Z(n54303) );
  IV U66891 ( .A(n54299), .Z(n54300) );
  NOR U66892 ( .A(n54301), .B(n54300), .Z(n54302) );
  NOR U66893 ( .A(n54303), .B(n54302), .Z(n55891) );
  XOR U66894 ( .A(n54304), .B(n55891), .Z(n55893) );
  XOR U66895 ( .A(n55892), .B(n55893), .Z(n57960) );
  XOR U66896 ( .A(n57961), .B(n57960), .Z(n54305) );
  IV U66897 ( .A(n54305), .Z(n55883) );
  XOR U66898 ( .A(n55882), .B(n55883), .Z(n55886) );
  XOR U66899 ( .A(n55885), .B(n55886), .Z(n57977) );
  XOR U66900 ( .A(n57976), .B(n57977), .Z(n57981) );
  IV U66901 ( .A(n54306), .Z(n54308) );
  NOR U66902 ( .A(n54308), .B(n54307), .Z(n57979) );
  XOR U66903 ( .A(n57981), .B(n57979), .Z(n54321) );
  IV U66904 ( .A(n54321), .Z(n54309) );
  NOR U66905 ( .A(n54320), .B(n54309), .Z(n54318) );
  IV U66906 ( .A(n54318), .Z(n54310) );
  NOR U66907 ( .A(n54317), .B(n54310), .Z(n54326) );
  NOR U66908 ( .A(n54312), .B(n54311), .Z(n54313) );
  IV U66909 ( .A(n54313), .Z(n54314) );
  NOR U66910 ( .A(n54315), .B(n54314), .Z(n54328) );
  IV U66911 ( .A(n54328), .Z(n54316) );
  NOR U66912 ( .A(n54326), .B(n54316), .Z(n57984) );
  IV U66913 ( .A(n54317), .Z(n54319) );
  NOR U66914 ( .A(n54319), .B(n54318), .Z(n54324) );
  IV U66915 ( .A(n54320), .Z(n54322) );
  NOR U66916 ( .A(n54322), .B(n54321), .Z(n54323) );
  NOR U66917 ( .A(n54324), .B(n54323), .Z(n54325) );
  IV U66918 ( .A(n54325), .Z(n57985) );
  NOR U66919 ( .A(n54326), .B(n57985), .Z(n54327) );
  NOR U66920 ( .A(n54328), .B(n54327), .Z(n54329) );
  NOR U66921 ( .A(n57984), .B(n54329), .Z(n54330) );
  IV U66922 ( .A(n54330), .Z(n58027) );
  NOR U66923 ( .A(n54331), .B(n58027), .Z(n54334) );
  NOR U66924 ( .A(n58025), .B(n54332), .Z(n54333) );
  XOR U66925 ( .A(n54334), .B(n54333), .Z(n55874) );
  IV U66926 ( .A(n54339), .Z(n54335) );
  NOR U66927 ( .A(n54336), .B(n54335), .Z(n54347) );
  NOR U66928 ( .A(n54338), .B(n54337), .Z(n54345) );
  NOR U66929 ( .A(n54340), .B(n54339), .Z(n54342) );
  NOR U66930 ( .A(n54342), .B(n54341), .Z(n54343) );
  IV U66931 ( .A(n54343), .Z(n54344) );
  NOR U66932 ( .A(n54345), .B(n54344), .Z(n54346) );
  NOR U66933 ( .A(n54347), .B(n54346), .Z(n55876) );
  XOR U66934 ( .A(n55874), .B(n55876), .Z(n55879) );
  XOR U66935 ( .A(n55877), .B(n55879), .Z(n58021) );
  XOR U66936 ( .A(n58020), .B(n58021), .Z(n58022) );
  XOR U66937 ( .A(n58023), .B(n58022), .Z(n58006) );
  XOR U66938 ( .A(n58008), .B(n58006), .Z(n58009) );
  XOR U66939 ( .A(n58010), .B(n58009), .Z(n54348) );
  IV U66940 ( .A(n54348), .Z(n58002) );
  XOR U66941 ( .A(n58001), .B(n58002), .Z(n57996) );
  IV U66942 ( .A(n54349), .Z(n54351) );
  NOR U66943 ( .A(n54351), .B(n54350), .Z(n58000) );
  NOR U66944 ( .A(n54353), .B(n54352), .Z(n57995) );
  NOR U66945 ( .A(n58000), .B(n57995), .Z(n54354) );
  XOR U66946 ( .A(n57996), .B(n54354), .Z(n54355) );
  IV U66947 ( .A(n54355), .Z(n57993) );
  NOR U66948 ( .A(n54356), .B(n57992), .Z(n54357) );
  NOR U66949 ( .A(n54358), .B(n54357), .Z(n54359) );
  XOR U66950 ( .A(n57993), .B(n54359), .Z(n58037) );
  IV U66951 ( .A(n54360), .Z(n54362) );
  NOR U66952 ( .A(n54362), .B(n54361), .Z(n58036) );
  IV U66953 ( .A(n54363), .Z(n55870) );
  IV U66954 ( .A(n54364), .Z(n54365) );
  NOR U66955 ( .A(n55870), .B(n54365), .Z(n54366) );
  NOR U66956 ( .A(n58036), .B(n54366), .Z(n54367) );
  XOR U66957 ( .A(n58037), .B(n54367), .Z(n58033) );
  XOR U66958 ( .A(n58035), .B(n58033), .Z(n58018) );
  XOR U66959 ( .A(n58017), .B(n58018), .Z(n54368) );
  NOR U66960 ( .A(n54369), .B(n54368), .Z(n58055) );
  IV U66961 ( .A(n54370), .Z(n54372) );
  NOR U66962 ( .A(n54372), .B(n54371), .Z(n55865) );
  IV U66963 ( .A(n54373), .Z(n54375) );
  NOR U66964 ( .A(n54375), .B(n54374), .Z(n55863) );
  NOR U66965 ( .A(n58017), .B(n55863), .Z(n54376) );
  XOR U66966 ( .A(n54376), .B(n58018), .Z(n54377) );
  IV U66967 ( .A(n54377), .Z(n55866) );
  XOR U66968 ( .A(n55865), .B(n55866), .Z(n58053) );
  IV U66969 ( .A(n58053), .Z(n54378) );
  NOR U66970 ( .A(n54379), .B(n54378), .Z(n54380) );
  NOR U66971 ( .A(n58055), .B(n54380), .Z(n58045) );
  IV U66972 ( .A(n54381), .Z(n54382) );
  NOR U66973 ( .A(n54383), .B(n54382), .Z(n58051) );
  IV U66974 ( .A(n54384), .Z(n54386) );
  NOR U66975 ( .A(n54386), .B(n54385), .Z(n58046) );
  NOR U66976 ( .A(n58051), .B(n58046), .Z(n54387) );
  XOR U66977 ( .A(n58045), .B(n54387), .Z(n58070) );
  XOR U66978 ( .A(n54388), .B(n58070), .Z(n55857) );
  XOR U66979 ( .A(n54389), .B(n55857), .Z(n55856) );
  XOR U66980 ( .A(n55854), .B(n55856), .Z(n58062) );
  XOR U66981 ( .A(n58063), .B(n58062), .Z(n55815) );
  XOR U66982 ( .A(n54390), .B(n55815), .Z(n55818) );
  XOR U66983 ( .A(n55819), .B(n55818), .Z(n54394) );
  IV U66984 ( .A(n54394), .Z(n54391) );
  NOR U66985 ( .A(n54393), .B(n54391), .Z(n54397) );
  IV U66986 ( .A(n54397), .Z(n54392) );
  NOR U66987 ( .A(n54396), .B(n54392), .Z(n55813) );
  IV U66988 ( .A(n54393), .Z(n54395) );
  NOR U66989 ( .A(n54395), .B(n54394), .Z(n54400) );
  IV U66990 ( .A(n54396), .Z(n54398) );
  NOR U66991 ( .A(n54398), .B(n54397), .Z(n54399) );
  NOR U66992 ( .A(n54400), .B(n54399), .Z(n54401) );
  IV U66993 ( .A(n54401), .Z(n55811) );
  NOR U66994 ( .A(n55813), .B(n55811), .Z(n54402) );
  XOR U66995 ( .A(n54403), .B(n54402), .Z(n55827) );
  XOR U66996 ( .A(n55825), .B(n55827), .Z(n55839) );
  XOR U66997 ( .A(n55838), .B(n55839), .Z(n55836) );
  XOR U66998 ( .A(n55837), .B(n55836), .Z(n55851) );
  XOR U66999 ( .A(n55852), .B(n55851), .Z(n55799) );
  XOR U67000 ( .A(n55798), .B(n55799), .Z(n55802) );
  XOR U67001 ( .A(n55801), .B(n55802), .Z(n58093) );
  XOR U67002 ( .A(n58091), .B(n58093), .Z(n58095) );
  XOR U67003 ( .A(n58094), .B(n58095), .Z(n58089) );
  XOR U67004 ( .A(n58090), .B(n58089), .Z(n54406) );
  IV U67005 ( .A(n54406), .Z(n54404) );
  NOR U67006 ( .A(n54405), .B(n54404), .Z(n58087) );
  NOR U67007 ( .A(n54407), .B(n54406), .Z(n58085) );
  NOR U67008 ( .A(n54409), .B(n54408), .Z(n58084) );
  XOR U67009 ( .A(n58085), .B(n58084), .Z(n54410) );
  NOR U67010 ( .A(n58087), .B(n54410), .Z(n54411) );
  IV U67011 ( .A(n54411), .Z(n58123) );
  IV U67012 ( .A(n54412), .Z(n54414) );
  NOR U67013 ( .A(n54414), .B(n54413), .Z(n58121) );
  XOR U67014 ( .A(n58123), .B(n58121), .Z(n58124) );
  XOR U67015 ( .A(n58125), .B(n58124), .Z(n58109) );
  XOR U67016 ( .A(n58110), .B(n58109), .Z(n54415) );
  XOR U67017 ( .A(n54416), .B(n54415), .Z(n54417) );
  IV U67018 ( .A(n54417), .Z(n55741) );
  XOR U67019 ( .A(n55739), .B(n55741), .Z(n55742) );
  IV U67020 ( .A(n55742), .Z(n54427) );
  IV U67021 ( .A(n54418), .Z(n54420) );
  NOR U67022 ( .A(n54420), .B(n54419), .Z(n54426) );
  IV U67023 ( .A(n54421), .Z(n54424) );
  IV U67024 ( .A(n54422), .Z(n54423) );
  NOR U67025 ( .A(n54424), .B(n54423), .Z(n54425) );
  NOR U67026 ( .A(n54426), .B(n54425), .Z(n55743) );
  XOR U67027 ( .A(n54427), .B(n55743), .Z(n55733) );
  XOR U67028 ( .A(n55731), .B(n55733), .Z(n55735) );
  XOR U67029 ( .A(n55734), .B(n55735), .Z(n55752) );
  XOR U67030 ( .A(n55750), .B(n55752), .Z(n55754) );
  XOR U67031 ( .A(n55748), .B(n55754), .Z(n54428) );
  NOR U67032 ( .A(n54429), .B(n54428), .Z(n55789) );
  IV U67033 ( .A(n54430), .Z(n54431) );
  NOR U67034 ( .A(n54432), .B(n54431), .Z(n54433) );
  IV U67035 ( .A(n54433), .Z(n55788) );
  XOR U67036 ( .A(n54435), .B(n54434), .Z(n54437) );
  NOR U67037 ( .A(n54437), .B(n54436), .Z(n55753) );
  NOR U67038 ( .A(n55748), .B(n55753), .Z(n54438) );
  XOR U67039 ( .A(n54438), .B(n55754), .Z(n54439) );
  IV U67040 ( .A(n54439), .Z(n55787) );
  XOR U67041 ( .A(n55788), .B(n55787), .Z(n54440) );
  NOR U67042 ( .A(n54441), .B(n54440), .Z(n54442) );
  NOR U67043 ( .A(n55789), .B(n54442), .Z(n55784) );
  IV U67044 ( .A(n54443), .Z(n54444) );
  NOR U67045 ( .A(n54445), .B(n54444), .Z(n54446) );
  IV U67046 ( .A(n54446), .Z(n55785) );
  XOR U67047 ( .A(n55784), .B(n55785), .Z(n55765) );
  IV U67048 ( .A(n55765), .Z(n55764) );
  XOR U67049 ( .A(n55768), .B(n55764), .Z(n54447) );
  XOR U67050 ( .A(n55766), .B(n54447), .Z(n55779) );
  XOR U67051 ( .A(n54448), .B(n55779), .Z(n55704) );
  XOR U67052 ( .A(n54449), .B(n55704), .Z(n55709) );
  XOR U67053 ( .A(n55707), .B(n55709), .Z(n55697) );
  XOR U67054 ( .A(n55696), .B(n55697), .Z(n55694) );
  NOR U67055 ( .A(n54450), .B(n55694), .Z(n55714) );
  IV U67056 ( .A(n54451), .Z(n54453) );
  IV U67057 ( .A(n54452), .Z(n54456) );
  NOR U67058 ( .A(n54453), .B(n54456), .Z(n54454) );
  IV U67059 ( .A(n54454), .Z(n55692) );
  IV U67060 ( .A(n54455), .Z(n54457) );
  NOR U67061 ( .A(n54457), .B(n54456), .Z(n55693) );
  XOR U67062 ( .A(n55693), .B(n55694), .Z(n55691) );
  XOR U67063 ( .A(n55692), .B(n55691), .Z(n54458) );
  NOR U67064 ( .A(n54459), .B(n54458), .Z(n54460) );
  NOR U67065 ( .A(n55714), .B(n54460), .Z(n55715) );
  IV U67066 ( .A(n54461), .Z(n54463) );
  NOR U67067 ( .A(n54463), .B(n54462), .Z(n54468) );
  IV U67068 ( .A(n54464), .Z(n54465) );
  NOR U67069 ( .A(n54466), .B(n54465), .Z(n54467) );
  NOR U67070 ( .A(n54468), .B(n54467), .Z(n55717) );
  XOR U67071 ( .A(n55715), .B(n55717), .Z(n55712) );
  XOR U67072 ( .A(n55713), .B(n55712), .Z(n58153) );
  XOR U67073 ( .A(n58155), .B(n58153), .Z(n58165) );
  IV U67074 ( .A(n58165), .Z(n54477) );
  IV U67075 ( .A(n54469), .Z(n54470) );
  NOR U67076 ( .A(n54471), .B(n54470), .Z(n58163) );
  IV U67077 ( .A(n54472), .Z(n54475) );
  IV U67078 ( .A(n54473), .Z(n54474) );
  NOR U67079 ( .A(n54475), .B(n54474), .Z(n58156) );
  NOR U67080 ( .A(n58163), .B(n58156), .Z(n54476) );
  XOR U67081 ( .A(n54477), .B(n54476), .Z(n58162) );
  NOR U67082 ( .A(n54479), .B(n54478), .Z(n54481) );
  NOR U67083 ( .A(n54481), .B(n54480), .Z(n58160) );
  XOR U67084 ( .A(n58162), .B(n58160), .Z(n55729) );
  XOR U67085 ( .A(n55727), .B(n55729), .Z(n58180) );
  XOR U67086 ( .A(n54482), .B(n58180), .Z(n54483) );
  IV U67087 ( .A(n54483), .Z(n58177) );
  XOR U67088 ( .A(n58176), .B(n58177), .Z(n55685) );
  XOR U67089 ( .A(n55682), .B(n55685), .Z(n58140) );
  XOR U67090 ( .A(n54484), .B(n58140), .Z(n54485) );
  IV U67091 ( .A(n54485), .Z(n58193) );
  XOR U67092 ( .A(n58191), .B(n58193), .Z(n58142) );
  XOR U67093 ( .A(n58141), .B(n58142), .Z(n58145) );
  XOR U67094 ( .A(n58144), .B(n58145), .Z(n58225) );
  IV U67095 ( .A(n54486), .Z(n54488) );
  NOR U67096 ( .A(n54488), .B(n54487), .Z(n58223) );
  XOR U67097 ( .A(n58225), .B(n58223), .Z(n58227) );
  XOR U67098 ( .A(n58226), .B(n58227), .Z(n58196) );
  NOR U67099 ( .A(n54490), .B(n54489), .Z(n54496) );
  IV U67100 ( .A(n54490), .Z(n54491) );
  NOR U67101 ( .A(n54492), .B(n54491), .Z(n54493) );
  NOR U67102 ( .A(n54494), .B(n54493), .Z(n54495) );
  NOR U67103 ( .A(n54496), .B(n54495), .Z(n58194) );
  XOR U67104 ( .A(n58196), .B(n58194), .Z(n58185) );
  IV U67105 ( .A(n54497), .Z(n54501) );
  NOR U67106 ( .A(n54499), .B(n54498), .Z(n54500) );
  IV U67107 ( .A(n54500), .Z(n54503) );
  NOR U67108 ( .A(n54501), .B(n54503), .Z(n58183) );
  XOR U67109 ( .A(n58185), .B(n58183), .Z(n58188) );
  IV U67110 ( .A(n54502), .Z(n54504) );
  NOR U67111 ( .A(n54504), .B(n54503), .Z(n58186) );
  XOR U67112 ( .A(n58188), .B(n58186), .Z(n55648) );
  IV U67113 ( .A(n55648), .Z(n55647) );
  XOR U67114 ( .A(n55651), .B(n55647), .Z(n54505) );
  XOR U67115 ( .A(n55649), .B(n54505), .Z(n55643) );
  IV U67116 ( .A(n55643), .Z(n55638) );
  NOR U67117 ( .A(n54507), .B(n54506), .Z(n54513) );
  IV U67118 ( .A(n54508), .Z(n54511) );
  IV U67119 ( .A(n54509), .Z(n54510) );
  NOR U67120 ( .A(n54511), .B(n54510), .Z(n54512) );
  NOR U67121 ( .A(n54513), .B(n54512), .Z(n55642) );
  IV U67122 ( .A(n55642), .Z(n55637) );
  XOR U67123 ( .A(n55638), .B(n55637), .Z(n54514) );
  XOR U67124 ( .A(n54515), .B(n54514), .Z(n58220) );
  XOR U67125 ( .A(n58207), .B(n58220), .Z(n54516) );
  XOR U67126 ( .A(n58211), .B(n54516), .Z(n55659) );
  XOR U67127 ( .A(n54517), .B(n55659), .Z(n55656) );
  XOR U67128 ( .A(n54518), .B(n55656), .Z(n55663) );
  XOR U67129 ( .A(n55664), .B(n55663), .Z(n55673) );
  XOR U67130 ( .A(n55675), .B(n55673), .Z(n55625) );
  XOR U67131 ( .A(n54519), .B(n55625), .Z(n54520) );
  IV U67132 ( .A(n54520), .Z(n55628) );
  XOR U67133 ( .A(n55626), .B(n55628), .Z(n55631) );
  IV U67134 ( .A(n54521), .Z(n54523) );
  NOR U67135 ( .A(n54523), .B(n54522), .Z(n55629) );
  XOR U67136 ( .A(n55631), .B(n55629), .Z(n58256) );
  XOR U67137 ( .A(n58255), .B(n58256), .Z(n58260) );
  IV U67138 ( .A(n54524), .Z(n54525) );
  NOR U67139 ( .A(n54526), .B(n54525), .Z(n58258) );
  XOR U67140 ( .A(n58260), .B(n58258), .Z(n58243) );
  XOR U67141 ( .A(n58242), .B(n58243), .Z(n58246) );
  XOR U67142 ( .A(n58245), .B(n58246), .Z(n58240) );
  XOR U67143 ( .A(n58239), .B(n58240), .Z(n55582) );
  XOR U67144 ( .A(n55583), .B(n55582), .Z(n55591) );
  XOR U67145 ( .A(n55592), .B(n55591), .Z(n55595) );
  XOR U67146 ( .A(n55594), .B(n55595), .Z(n55612) );
  XOR U67147 ( .A(n55611), .B(n55612), .Z(n55585) );
  XOR U67148 ( .A(n55584), .B(n55585), .Z(n55587) );
  XOR U67149 ( .A(n55588), .B(n55587), .Z(n54527) );
  IV U67150 ( .A(n54527), .Z(n55575) );
  XOR U67151 ( .A(n55574), .B(n55575), .Z(n55578) );
  XOR U67152 ( .A(n55577), .B(n55578), .Z(n55615) );
  XOR U67153 ( .A(n55614), .B(n55615), .Z(n55604) );
  XOR U67154 ( .A(n55603), .B(n55604), .Z(n55608) );
  IV U67155 ( .A(n54528), .Z(n54530) );
  NOR U67156 ( .A(n54530), .B(n54529), .Z(n55606) );
  XOR U67157 ( .A(n55608), .B(n55606), .Z(n55536) );
  XOR U67158 ( .A(n55535), .B(n55536), .Z(n55538) );
  IV U67159 ( .A(n54531), .Z(n54533) );
  NOR U67160 ( .A(n54533), .B(n54532), .Z(n54540) );
  IV U67161 ( .A(n54540), .Z(n54534) );
  NOR U67162 ( .A(n55538), .B(n54534), .Z(n55550) );
  IV U67163 ( .A(n54535), .Z(n54536) );
  NOR U67164 ( .A(n54537), .B(n54536), .Z(n54538) );
  IV U67165 ( .A(n54538), .Z(n55539) );
  XOR U67166 ( .A(n55539), .B(n55538), .Z(n54539) );
  NOR U67167 ( .A(n54540), .B(n54539), .Z(n55548) );
  XOR U67168 ( .A(n55548), .B(n55547), .Z(n54541) );
  NOR U67169 ( .A(n55550), .B(n54541), .Z(n54542) );
  IV U67170 ( .A(n54542), .Z(n55546) );
  NOR U67171 ( .A(n54544), .B(n54543), .Z(n54545) );
  NOR U67172 ( .A(n54546), .B(n54545), .Z(n55544) );
  XOR U67173 ( .A(n55546), .B(n55544), .Z(n55528) );
  XOR U67174 ( .A(n55529), .B(n55528), .Z(n55530) );
  XOR U67175 ( .A(n55532), .B(n55530), .Z(n55567) );
  XOR U67176 ( .A(n54547), .B(n55567), .Z(n55523) );
  IV U67177 ( .A(n54548), .Z(n54549) );
  NOR U67178 ( .A(n54550), .B(n54549), .Z(n54560) );
  IV U67179 ( .A(n54560), .Z(n55525) );
  NOR U67180 ( .A(n55523), .B(n55525), .Z(n54562) );
  XOR U67181 ( .A(n55521), .B(n55567), .Z(n54555) );
  IV U67182 ( .A(n54551), .Z(n54553) );
  NOR U67183 ( .A(n54553), .B(n54552), .Z(n54556) );
  IV U67184 ( .A(n54556), .Z(n54554) );
  NOR U67185 ( .A(n54555), .B(n54554), .Z(n55568) );
  NOR U67186 ( .A(n55523), .B(n54556), .Z(n54557) );
  NOR U67187 ( .A(n55568), .B(n54557), .Z(n54558) );
  IV U67188 ( .A(n54558), .Z(n54559) );
  NOR U67189 ( .A(n54560), .B(n54559), .Z(n54561) );
  NOR U67190 ( .A(n54562), .B(n54561), .Z(n55558) );
  XOR U67191 ( .A(n55557), .B(n55558), .Z(n55562) );
  XOR U67192 ( .A(n55560), .B(n55562), .Z(n58280) );
  NOR U67193 ( .A(n54563), .B(n58280), .Z(n54569) );
  IV U67194 ( .A(n54564), .Z(n54567) );
  NOR U67195 ( .A(n54576), .B(n54565), .Z(n54577) );
  XOR U67196 ( .A(n58280), .B(n54577), .Z(n54566) );
  NOR U67197 ( .A(n54567), .B(n54566), .Z(n54568) );
  NOR U67198 ( .A(n54569), .B(n54568), .Z(n54570) );
  NOR U67199 ( .A(n54576), .B(n54570), .Z(n54571) );
  IV U67200 ( .A(n54571), .Z(n54572) );
  NOR U67201 ( .A(n54573), .B(n54572), .Z(n58282) );
  IV U67202 ( .A(n54574), .Z(n54575) );
  NOR U67203 ( .A(n54576), .B(n54575), .Z(n54579) );
  IV U67204 ( .A(n54577), .Z(n58281) );
  XOR U67205 ( .A(n58281), .B(n58280), .Z(n54578) );
  NOR U67206 ( .A(n54579), .B(n54578), .Z(n54580) );
  NOR U67207 ( .A(n58282), .B(n54580), .Z(n54581) );
  IV U67208 ( .A(n54581), .Z(n58278) );
  XOR U67209 ( .A(n58277), .B(n58278), .Z(n54588) );
  IV U67210 ( .A(n54588), .Z(n54582) );
  NOR U67211 ( .A(n54587), .B(n54582), .Z(n54585) );
  IV U67212 ( .A(n54585), .Z(n54583) );
  NOR U67213 ( .A(n54584), .B(n54583), .Z(n58276) );
  IV U67214 ( .A(n54584), .Z(n54586) );
  NOR U67215 ( .A(n54586), .B(n54585), .Z(n54591) );
  IV U67216 ( .A(n54587), .Z(n54589) );
  NOR U67217 ( .A(n54589), .B(n54588), .Z(n54590) );
  NOR U67218 ( .A(n54591), .B(n54590), .Z(n54592) );
  IV U67219 ( .A(n54592), .Z(n58274) );
  NOR U67220 ( .A(n58276), .B(n58274), .Z(n58293) );
  XOR U67221 ( .A(n54593), .B(n58293), .Z(n58291) );
  XOR U67222 ( .A(n58289), .B(n58291), .Z(n58312) );
  XOR U67223 ( .A(n58311), .B(n58312), .Z(n58315) );
  XOR U67224 ( .A(n58314), .B(n58315), .Z(n58305) );
  XOR U67225 ( .A(n58304), .B(n58305), .Z(n58307) );
  XOR U67226 ( .A(n58308), .B(n58307), .Z(n58328) );
  XOR U67227 ( .A(n58330), .B(n58328), .Z(n55514) );
  XOR U67228 ( .A(n55513), .B(n55514), .Z(n55517) );
  XOR U67229 ( .A(n55516), .B(n55517), .Z(n58332) );
  XOR U67230 ( .A(n58331), .B(n58332), .Z(n58327) );
  XOR U67231 ( .A(n58325), .B(n58327), .Z(n58345) );
  XOR U67232 ( .A(n54594), .B(n58345), .Z(n58341) );
  IV U67233 ( .A(n54595), .Z(n54596) );
  NOR U67234 ( .A(n54597), .B(n54596), .Z(n54598) );
  IV U67235 ( .A(n54598), .Z(n58342) );
  XOR U67236 ( .A(n58341), .B(n58342), .Z(n58352) );
  XOR U67237 ( .A(n58351), .B(n58352), .Z(n58355) );
  XOR U67238 ( .A(n58354), .B(n58355), .Z(n58349) );
  XOR U67239 ( .A(n58348), .B(n58349), .Z(n58382) );
  IV U67240 ( .A(n54599), .Z(n54602) );
  IV U67241 ( .A(n54600), .Z(n54601) );
  NOR U67242 ( .A(n54602), .B(n54601), .Z(n58379) );
  IV U67243 ( .A(n58379), .Z(n58381) );
  XOR U67244 ( .A(n58382), .B(n58381), .Z(n58371) );
  IV U67245 ( .A(n54603), .Z(n54604) );
  NOR U67246 ( .A(n54605), .B(n54604), .Z(n58384) );
  NOR U67247 ( .A(n54607), .B(n54606), .Z(n58372) );
  NOR U67248 ( .A(n58384), .B(n58372), .Z(n54608) );
  XOR U67249 ( .A(n58371), .B(n54608), .Z(n58370) );
  NOR U67250 ( .A(n54610), .B(n54609), .Z(n54614) );
  IV U67251 ( .A(n54614), .Z(n54611) );
  NOR U67252 ( .A(n58370), .B(n54611), .Z(n58368) );
  IV U67253 ( .A(n54612), .Z(n58369) );
  XOR U67254 ( .A(n58369), .B(n58370), .Z(n54613) );
  NOR U67255 ( .A(n54614), .B(n54613), .Z(n58366) );
  NOR U67256 ( .A(n58368), .B(n58366), .Z(n55479) );
  IV U67257 ( .A(n54615), .Z(n54617) );
  NOR U67258 ( .A(n54617), .B(n54616), .Z(n55480) );
  NOR U67259 ( .A(n58364), .B(n55480), .Z(n54618) );
  XOR U67260 ( .A(n55479), .B(n54618), .Z(n55489) );
  IV U67261 ( .A(n54619), .Z(n54620) );
  NOR U67262 ( .A(n54621), .B(n54620), .Z(n55477) );
  NOR U67263 ( .A(n54623), .B(n54622), .Z(n55487) );
  NOR U67264 ( .A(n55477), .B(n55487), .Z(n54624) );
  XOR U67265 ( .A(n55489), .B(n54624), .Z(n55474) );
  NOR U67266 ( .A(n54626), .B(n54625), .Z(n54636) );
  IV U67267 ( .A(n54636), .Z(n55476) );
  NOR U67268 ( .A(n55474), .B(n55476), .Z(n54638) );
  IV U67269 ( .A(n54627), .Z(n54629) );
  NOR U67270 ( .A(n54629), .B(n54628), .Z(n54632) );
  IV U67271 ( .A(n54632), .Z(n54631) );
  XOR U67272 ( .A(n55477), .B(n55489), .Z(n54630) );
  NOR U67273 ( .A(n54631), .B(n54630), .Z(n55490) );
  NOR U67274 ( .A(n55474), .B(n54632), .Z(n54633) );
  NOR U67275 ( .A(n55490), .B(n54633), .Z(n54634) );
  IV U67276 ( .A(n54634), .Z(n54635) );
  NOR U67277 ( .A(n54636), .B(n54635), .Z(n54637) );
  NOR U67278 ( .A(n54638), .B(n54637), .Z(n55467) );
  XOR U67279 ( .A(n55466), .B(n55467), .Z(n55470) );
  XOR U67280 ( .A(n55469), .B(n55470), .Z(n55502) );
  XOR U67281 ( .A(n55501), .B(n55502), .Z(n55506) );
  IV U67282 ( .A(n54639), .Z(n54641) );
  NOR U67283 ( .A(n54641), .B(n54640), .Z(n55504) );
  XOR U67284 ( .A(n55506), .B(n55504), .Z(n55494) );
  XOR U67285 ( .A(n55495), .B(n55494), .Z(n55496) );
  XOR U67286 ( .A(n55498), .B(n55496), .Z(n55459) );
  XOR U67287 ( .A(n55457), .B(n55459), .Z(n55460) );
  XOR U67288 ( .A(n55461), .B(n55460), .Z(n54644) );
  IV U67289 ( .A(n54644), .Z(n54642) );
  NOR U67290 ( .A(n54643), .B(n54642), .Z(n55446) );
  NOR U67291 ( .A(n54645), .B(n54644), .Z(n55444) );
  IV U67292 ( .A(n54646), .Z(n54648) );
  NOR U67293 ( .A(n54648), .B(n54647), .Z(n55443) );
  XOR U67294 ( .A(n55444), .B(n55443), .Z(n54649) );
  NOR U67295 ( .A(n55446), .B(n54649), .Z(n55438) );
  NOR U67296 ( .A(n54651), .B(n54650), .Z(n55440) );
  IV U67297 ( .A(n54652), .Z(n54654) );
  NOR U67298 ( .A(n54654), .B(n54653), .Z(n54655) );
  IV U67299 ( .A(n54655), .Z(n54656) );
  NOR U67300 ( .A(n54657), .B(n54656), .Z(n54658) );
  NOR U67301 ( .A(n55439), .B(n54658), .Z(n54659) );
  XOR U67302 ( .A(n55440), .B(n54659), .Z(n54660) );
  XOR U67303 ( .A(n55438), .B(n54660), .Z(n54672) );
  XOR U67304 ( .A(n54661), .B(n54672), .Z(n54662) );
  IV U67305 ( .A(n54662), .Z(n55452) );
  NOR U67306 ( .A(n54670), .B(n55452), .Z(n54675) );
  IV U67307 ( .A(n54685), .Z(n54669) );
  NOR U67308 ( .A(n54664), .B(n54663), .Z(n54665) );
  IV U67309 ( .A(n54665), .Z(n54681) );
  NOR U67310 ( .A(n54666), .B(n54681), .Z(n54667) );
  IV U67311 ( .A(n54667), .Z(n54668) );
  NOR U67312 ( .A(n54669), .B(n54668), .Z(n54677) );
  IV U67313 ( .A(n54670), .Z(n54671) );
  NOR U67314 ( .A(n54672), .B(n54671), .Z(n54673) );
  NOR U67315 ( .A(n54677), .B(n54673), .Z(n54674) );
  NOR U67316 ( .A(n54675), .B(n54674), .Z(n55454) );
  IV U67317 ( .A(n54675), .Z(n54676) );
  NOR U67318 ( .A(n54677), .B(n54676), .Z(n54678) );
  NOR U67319 ( .A(n55454), .B(n54678), .Z(n54679) );
  IV U67320 ( .A(n54679), .Z(n55415) );
  IV U67321 ( .A(n54680), .Z(n54682) );
  NOR U67322 ( .A(n54682), .B(n54681), .Z(n54683) );
  IV U67323 ( .A(n54683), .Z(n54684) );
  NOR U67324 ( .A(n54685), .B(n54684), .Z(n55413) );
  XOR U67325 ( .A(n55415), .B(n55413), .Z(n55417) );
  XOR U67326 ( .A(n55416), .B(n55417), .Z(n55406) );
  XOR U67327 ( .A(n55405), .B(n55406), .Z(n55410) );
  XOR U67328 ( .A(n55408), .B(n55410), .Z(n55425) );
  XOR U67329 ( .A(n55423), .B(n55425), .Z(n58409) );
  XOR U67330 ( .A(n54686), .B(n58409), .Z(n54687) );
  IV U67331 ( .A(n54687), .Z(n58412) );
  XOR U67332 ( .A(n58410), .B(n58412), .Z(n55430) );
  XOR U67333 ( .A(n55429), .B(n55430), .Z(n58415) );
  IV U67334 ( .A(n54688), .Z(n54689) );
  NOR U67335 ( .A(n54690), .B(n54689), .Z(n58413) );
  XOR U67336 ( .A(n58415), .B(n58413), .Z(n55435) );
  XOR U67337 ( .A(n55433), .B(n55435), .Z(n58427) );
  IV U67338 ( .A(n58427), .Z(n54698) );
  IV U67339 ( .A(n54691), .Z(n54693) );
  NOR U67340 ( .A(n54693), .B(n54692), .Z(n55432) );
  IV U67341 ( .A(n54694), .Z(n54696) );
  NOR U67342 ( .A(n54696), .B(n54695), .Z(n58425) );
  NOR U67343 ( .A(n55432), .B(n58425), .Z(n54697) );
  XOR U67344 ( .A(n54698), .B(n54697), .Z(n58424) );
  XOR U67345 ( .A(n58422), .B(n58424), .Z(n55402) );
  IV U67346 ( .A(n54699), .Z(n54700) );
  NOR U67347 ( .A(n54701), .B(n54700), .Z(n58421) );
  IV U67348 ( .A(n54702), .Z(n54703) );
  NOR U67349 ( .A(n54704), .B(n54703), .Z(n55400) );
  NOR U67350 ( .A(n58421), .B(n55400), .Z(n54705) );
  XOR U67351 ( .A(n55402), .B(n54705), .Z(n55397) );
  XOR U67352 ( .A(n55399), .B(n55397), .Z(n55384) );
  IV U67353 ( .A(n55384), .Z(n55381) );
  IV U67354 ( .A(n54706), .Z(n54707) );
  NOR U67355 ( .A(n54715), .B(n54707), .Z(n55386) );
  IV U67356 ( .A(n54708), .Z(n54710) );
  NOR U67357 ( .A(n54710), .B(n54709), .Z(n55382) );
  NOR U67358 ( .A(n55386), .B(n55382), .Z(n54711) );
  XOR U67359 ( .A(n55381), .B(n54711), .Z(n54719) );
  NOR U67360 ( .A(n54713), .B(n54712), .Z(n54717) );
  NOR U67361 ( .A(n54715), .B(n54714), .Z(n54716) );
  IV U67362 ( .A(n54716), .Z(n58401) );
  NOR U67363 ( .A(n54717), .B(n58401), .Z(n54718) );
  XOR U67364 ( .A(n54719), .B(n54718), .Z(n55380) );
  IV U67365 ( .A(n54720), .Z(n54721) );
  NOR U67366 ( .A(n54722), .B(n54721), .Z(n55378) );
  IV U67367 ( .A(n54723), .Z(n54724) );
  NOR U67368 ( .A(n54724), .B(n58401), .Z(n54725) );
  NOR U67369 ( .A(n55378), .B(n54725), .Z(n54726) );
  XOR U67370 ( .A(n55380), .B(n54726), .Z(n55303) );
  XOR U67371 ( .A(n55301), .B(n55303), .Z(n55324) );
  IV U67372 ( .A(n54727), .Z(n54728) );
  NOR U67373 ( .A(n54729), .B(n54728), .Z(n55302) );
  IV U67374 ( .A(n54730), .Z(n54731) );
  NOR U67375 ( .A(n54732), .B(n54731), .Z(n55325) );
  NOR U67376 ( .A(n55302), .B(n55325), .Z(n54733) );
  XOR U67377 ( .A(n55324), .B(n54733), .Z(n55323) );
  XOR U67378 ( .A(n55321), .B(n55323), .Z(n55310) );
  XOR U67379 ( .A(n55308), .B(n55310), .Z(n55312) );
  XOR U67380 ( .A(n55311), .B(n55312), .Z(n55306) );
  XOR U67381 ( .A(n55307), .B(n55306), .Z(n55350) );
  NOR U67382 ( .A(n54734), .B(n55350), .Z(n55349) );
  IV U67383 ( .A(n54734), .Z(n54735) );
  NOR U67384 ( .A(n54735), .B(n55306), .Z(n55346) );
  NOR U67385 ( .A(n55349), .B(n55346), .Z(n54743) );
  IV U67386 ( .A(n54736), .Z(n54738) );
  NOR U67387 ( .A(n54738), .B(n54737), .Z(n55347) );
  IV U67388 ( .A(n54739), .Z(n54741) );
  NOR U67389 ( .A(n54741), .B(n54740), .Z(n55351) );
  NOR U67390 ( .A(n55347), .B(n55351), .Z(n54742) );
  XOR U67391 ( .A(n54743), .B(n54742), .Z(n55336) );
  XOR U67392 ( .A(n55337), .B(n55336), .Z(n55338) );
  XOR U67393 ( .A(n55339), .B(n55338), .Z(n55363) );
  XOR U67394 ( .A(n54744), .B(n55363), .Z(n54745) );
  IV U67395 ( .A(n54745), .Z(n55360) );
  XOR U67396 ( .A(n55358), .B(n55360), .Z(n55371) );
  XOR U67397 ( .A(n55370), .B(n55371), .Z(n55375) );
  IV U67398 ( .A(n54746), .Z(n54747) );
  NOR U67399 ( .A(n54748), .B(n54747), .Z(n55373) );
  XOR U67400 ( .A(n55375), .B(n55373), .Z(n55282) );
  XOR U67401 ( .A(n55281), .B(n55282), .Z(n55284) );
  XOR U67402 ( .A(n55285), .B(n55284), .Z(n55248) );
  XOR U67403 ( .A(n55247), .B(n55248), .Z(n54751) );
  IV U67404 ( .A(n54751), .Z(n54749) );
  NOR U67405 ( .A(n54750), .B(n54749), .Z(n55291) );
  NOR U67406 ( .A(n54752), .B(n54751), .Z(n55289) );
  IV U67407 ( .A(n54753), .Z(n54756) );
  IV U67408 ( .A(n54754), .Z(n54755) );
  NOR U67409 ( .A(n54756), .B(n54755), .Z(n55288) );
  XOR U67410 ( .A(n55289), .B(n55288), .Z(n54757) );
  NOR U67411 ( .A(n55291), .B(n54757), .Z(n54758) );
  IV U67412 ( .A(n54758), .Z(n55296) );
  IV U67413 ( .A(n54759), .Z(n54760) );
  NOR U67414 ( .A(n54761), .B(n54760), .Z(n55294) );
  XOR U67415 ( .A(n55296), .B(n55294), .Z(n55272) );
  XOR U67416 ( .A(n54762), .B(n55272), .Z(n54763) );
  IV U67417 ( .A(n54763), .Z(n55275) );
  XOR U67418 ( .A(n55274), .B(n55275), .Z(n55264) );
  XOR U67419 ( .A(n55263), .B(n55264), .Z(n55267) );
  XOR U67420 ( .A(n55266), .B(n55267), .Z(n55199) );
  NOR U67421 ( .A(n54765), .B(n54764), .Z(n54771) );
  IV U67422 ( .A(n54765), .Z(n54766) );
  NOR U67423 ( .A(n54767), .B(n54766), .Z(n54768) );
  NOR U67424 ( .A(n54769), .B(n54768), .Z(n54770) );
  NOR U67425 ( .A(n54771), .B(n54770), .Z(n55197) );
  XOR U67426 ( .A(n55199), .B(n55197), .Z(n55256) );
  XOR U67427 ( .A(n55255), .B(n55256), .Z(n55259) );
  XOR U67428 ( .A(n55258), .B(n55259), .Z(n55201) );
  XOR U67429 ( .A(n55200), .B(n55201), .Z(n55190) );
  XOR U67430 ( .A(n55189), .B(n55190), .Z(n55193) );
  XOR U67431 ( .A(n55192), .B(n55193), .Z(n55208) );
  XOR U67432 ( .A(n55207), .B(n55208), .Z(n55210) );
  IV U67433 ( .A(n54774), .Z(n54772) );
  NOR U67434 ( .A(n54773), .B(n54772), .Z(n54780) );
  NOR U67435 ( .A(n54775), .B(n54774), .Z(n54778) );
  IV U67436 ( .A(n54776), .Z(n54777) );
  NOR U67437 ( .A(n54778), .B(n54777), .Z(n54779) );
  NOR U67438 ( .A(n54780), .B(n54779), .Z(n55211) );
  XOR U67439 ( .A(n55210), .B(n55211), .Z(n54783) );
  IV U67440 ( .A(n54783), .Z(n54781) );
  NOR U67441 ( .A(n54782), .B(n54781), .Z(n55217) );
  NOR U67442 ( .A(n54784), .B(n54783), .Z(n55215) );
  IV U67443 ( .A(n54785), .Z(n54786) );
  NOR U67444 ( .A(n54787), .B(n54786), .Z(n55214) );
  XOR U67445 ( .A(n55215), .B(n55214), .Z(n54788) );
  NOR U67446 ( .A(n55217), .B(n54788), .Z(n55220) );
  NOR U67447 ( .A(n54790), .B(n54789), .Z(n54792) );
  NOR U67448 ( .A(n54792), .B(n54791), .Z(n55222) );
  XOR U67449 ( .A(n55220), .B(n55222), .Z(n55228) );
  XOR U67450 ( .A(n55227), .B(n55228), .Z(n55231) );
  XOR U67451 ( .A(n55230), .B(n55231), .Z(n58465) );
  XOR U67452 ( .A(n58464), .B(n58465), .Z(n58469) );
  XOR U67453 ( .A(n58467), .B(n58469), .Z(n58457) );
  XOR U67454 ( .A(n58456), .B(n58457), .Z(n58461) );
  XOR U67455 ( .A(n58459), .B(n58461), .Z(n55241) );
  XOR U67456 ( .A(n55239), .B(n55241), .Z(n55243) );
  XOR U67457 ( .A(n55242), .B(n55243), .Z(n58484) );
  XOR U67458 ( .A(n58485), .B(n58484), .Z(n58486) );
  IV U67459 ( .A(n54796), .Z(n54794) );
  NOR U67460 ( .A(n54794), .B(n54793), .Z(n54801) );
  NOR U67461 ( .A(n54796), .B(n54795), .Z(n54799) );
  IV U67462 ( .A(n54797), .Z(n54798) );
  NOR U67463 ( .A(n54799), .B(n54798), .Z(n54800) );
  NOR U67464 ( .A(n54801), .B(n54800), .Z(n58488) );
  XOR U67465 ( .A(n58486), .B(n58488), .Z(n58497) );
  XOR U67466 ( .A(n58496), .B(n58497), .Z(n58500) );
  XOR U67467 ( .A(n58499), .B(n58500), .Z(n58495) );
  XOR U67468 ( .A(n58493), .B(n58495), .Z(n58478) );
  XOR U67469 ( .A(n58476), .B(n58478), .Z(n58480) );
  XOR U67470 ( .A(n58479), .B(n58480), .Z(n55181) );
  XOR U67471 ( .A(n55180), .B(n55181), .Z(n55183) );
  XOR U67472 ( .A(n55184), .B(n55183), .Z(n55169) );
  IV U67473 ( .A(n55169), .Z(n55171) );
  IV U67474 ( .A(n54802), .Z(n54804) );
  NOR U67475 ( .A(n54804), .B(n54803), .Z(n55174) );
  IV U67476 ( .A(n54805), .Z(n54807) );
  NOR U67477 ( .A(n54807), .B(n54806), .Z(n55170) );
  XOR U67478 ( .A(n55174), .B(n55170), .Z(n54808) );
  XOR U67479 ( .A(n55171), .B(n54808), .Z(n58560) );
  IV U67480 ( .A(n54809), .Z(n54810) );
  NOR U67481 ( .A(n54811), .B(n54810), .Z(n55173) );
  NOR U67482 ( .A(n54813), .B(n54812), .Z(n58558) );
  NOR U67483 ( .A(n55173), .B(n58558), .Z(n54814) );
  XOR U67484 ( .A(n58560), .B(n54814), .Z(n58564) );
  IV U67485 ( .A(n58564), .Z(n58562) );
  IV U67486 ( .A(n54815), .Z(n54816) );
  NOR U67487 ( .A(n54817), .B(n54816), .Z(n54822) );
  IV U67488 ( .A(n54818), .Z(n54819) );
  NOR U67489 ( .A(n54820), .B(n54819), .Z(n54821) );
  NOR U67490 ( .A(n54822), .B(n54821), .Z(n58561) );
  IV U67491 ( .A(n58561), .Z(n58563) );
  XOR U67492 ( .A(n58562), .B(n58563), .Z(n58515) );
  IV U67493 ( .A(n54823), .Z(n54825) );
  NOR U67494 ( .A(n54825), .B(n54824), .Z(n58565) );
  IV U67495 ( .A(n54826), .Z(n54828) );
  NOR U67496 ( .A(n54828), .B(n54827), .Z(n58513) );
  NOR U67497 ( .A(n58565), .B(n58513), .Z(n54829) );
  XOR U67498 ( .A(n58515), .B(n54829), .Z(n58516) );
  XOR U67499 ( .A(n58518), .B(n58516), .Z(n58519) );
  XOR U67500 ( .A(n58520), .B(n58519), .Z(n54830) );
  NOR U67501 ( .A(n54833), .B(n54830), .Z(n54837) );
  NOR U67502 ( .A(n54832), .B(n54831), .Z(n54839) );
  IV U67503 ( .A(n54833), .Z(n54834) );
  NOR U67504 ( .A(n58519), .B(n54834), .Z(n54835) );
  NOR U67505 ( .A(n54839), .B(n54835), .Z(n54836) );
  NOR U67506 ( .A(n54837), .B(n54836), .Z(n58531) );
  IV U67507 ( .A(n54837), .Z(n54838) );
  NOR U67508 ( .A(n54839), .B(n54838), .Z(n54840) );
  NOR U67509 ( .A(n58531), .B(n54840), .Z(n54848) );
  XOR U67510 ( .A(n58529), .B(n54848), .Z(n58526) );
  XOR U67511 ( .A(n58527), .B(n58526), .Z(n54850) );
  IV U67512 ( .A(n54850), .Z(n54845) );
  IV U67513 ( .A(n54841), .Z(n54842) );
  NOR U67514 ( .A(n54843), .B(n54842), .Z(n54854) );
  IV U67515 ( .A(n54854), .Z(n54844) );
  NOR U67516 ( .A(n54845), .B(n54844), .Z(n58553) );
  NOR U67517 ( .A(n54847), .B(n54846), .Z(n54851) );
  IV U67518 ( .A(n54851), .Z(n54849) );
  IV U67519 ( .A(n54848), .Z(n58528) );
  NOR U67520 ( .A(n54849), .B(n58528), .Z(n58554) );
  NOR U67521 ( .A(n54851), .B(n54850), .Z(n54852) );
  NOR U67522 ( .A(n58554), .B(n54852), .Z(n54853) );
  NOR U67523 ( .A(n54854), .B(n54853), .Z(n54855) );
  NOR U67524 ( .A(n58553), .B(n54855), .Z(n58540) );
  XOR U67525 ( .A(n58538), .B(n58540), .Z(n58551) );
  XOR U67526 ( .A(n54856), .B(n58551), .Z(n58604) );
  XOR U67527 ( .A(n58605), .B(n58604), .Z(n58608) );
  XOR U67528 ( .A(n58607), .B(n58608), .Z(n58598) );
  XOR U67529 ( .A(n58596), .B(n58598), .Z(n58601) );
  XOR U67530 ( .A(n58599), .B(n58601), .Z(n58622) );
  XOR U67531 ( .A(n58621), .B(n58622), .Z(n54857) );
  IV U67532 ( .A(n54857), .Z(n58589) );
  XOR U67533 ( .A(n54858), .B(n58589), .Z(n58619) );
  XOR U67534 ( .A(n58618), .B(n58619), .Z(n58577) );
  XOR U67535 ( .A(n58579), .B(n58577), .Z(n58581) );
  XOR U67536 ( .A(n58580), .B(n58581), .Z(n58584) );
  XOR U67537 ( .A(n58583), .B(n58584), .Z(n55157) );
  XOR U67538 ( .A(n55156), .B(n55157), .Z(n55161) );
  IV U67539 ( .A(n54859), .Z(n54861) );
  NOR U67540 ( .A(n54861), .B(n54860), .Z(n55159) );
  XOR U67541 ( .A(n55161), .B(n55159), .Z(n55154) );
  IV U67542 ( .A(n55154), .Z(n54870) );
  IV U67543 ( .A(n54862), .Z(n54864) );
  NOR U67544 ( .A(n54864), .B(n54863), .Z(n54869) );
  IV U67545 ( .A(n54865), .Z(n54867) );
  NOR U67546 ( .A(n54867), .B(n54866), .Z(n54868) );
  NOR U67547 ( .A(n54869), .B(n54868), .Z(n55155) );
  XOR U67548 ( .A(n54870), .B(n55155), .Z(n55148) );
  XOR U67549 ( .A(n55147), .B(n55148), .Z(n55150) );
  XOR U67550 ( .A(n55151), .B(n55150), .Z(n54871) );
  IV U67551 ( .A(n54871), .Z(n55141) );
  XOR U67552 ( .A(n55140), .B(n55141), .Z(n55143) );
  XOR U67553 ( .A(n55144), .B(n55143), .Z(n58634) );
  XOR U67554 ( .A(n58636), .B(n58634), .Z(n58637) );
  XOR U67555 ( .A(n58638), .B(n58637), .Z(n55132) );
  IV U67556 ( .A(n54872), .Z(n54873) );
  NOR U67557 ( .A(n54874), .B(n54873), .Z(n55133) );
  NOR U67558 ( .A(n55137), .B(n55133), .Z(n54875) );
  XOR U67559 ( .A(n55132), .B(n54875), .Z(n55131) );
  IV U67560 ( .A(n54876), .Z(n54878) );
  NOR U67561 ( .A(n54878), .B(n54877), .Z(n54879) );
  IV U67562 ( .A(n54879), .Z(n54886) );
  NOR U67563 ( .A(n55131), .B(n54886), .Z(n58658) );
  IV U67564 ( .A(n54880), .Z(n54881) );
  NOR U67565 ( .A(n54881), .B(n54885), .Z(n54882) );
  IV U67566 ( .A(n54882), .Z(n58648) );
  IV U67567 ( .A(n54883), .Z(n54884) );
  NOR U67568 ( .A(n54885), .B(n54884), .Z(n55129) );
  XOR U67569 ( .A(n55129), .B(n55131), .Z(n58647) );
  XOR U67570 ( .A(n58648), .B(n58647), .Z(n54889) );
  IV U67571 ( .A(n58647), .Z(n54887) );
  NOR U67572 ( .A(n54887), .B(n54886), .Z(n54888) );
  NOR U67573 ( .A(n54889), .B(n54888), .Z(n54890) );
  NOR U67574 ( .A(n58658), .B(n54890), .Z(n58649) );
  XOR U67575 ( .A(n58651), .B(n58649), .Z(n58656) );
  IV U67576 ( .A(n54891), .Z(n54895) );
  NOR U67577 ( .A(n54893), .B(n54892), .Z(n54894) );
  IV U67578 ( .A(n54894), .Z(n54897) );
  NOR U67579 ( .A(n54895), .B(n54897), .Z(n58654) );
  XOR U67580 ( .A(n58656), .B(n58654), .Z(n55123) );
  IV U67581 ( .A(n54896), .Z(n54898) );
  NOR U67582 ( .A(n54898), .B(n54897), .Z(n55121) );
  XOR U67583 ( .A(n55123), .B(n55121), .Z(n55125) );
  XOR U67584 ( .A(n55124), .B(n55125), .Z(n55115) );
  IV U67585 ( .A(n54899), .Z(n54901) );
  NOR U67586 ( .A(n54901), .B(n54900), .Z(n55113) );
  XOR U67587 ( .A(n55115), .B(n55113), .Z(n55117) );
  XOR U67588 ( .A(n55116), .B(n55117), .Z(n58673) );
  IV U67589 ( .A(n58673), .Z(n54910) );
  IV U67590 ( .A(n54902), .Z(n54904) );
  NOR U67591 ( .A(n54904), .B(n54903), .Z(n54909) );
  IV U67592 ( .A(n54905), .Z(n54906) );
  NOR U67593 ( .A(n54907), .B(n54906), .Z(n54908) );
  NOR U67594 ( .A(n54909), .B(n54908), .Z(n58674) );
  XOR U67595 ( .A(n54910), .B(n58674), .Z(n58676) );
  XOR U67596 ( .A(n58675), .B(n58676), .Z(n55095) );
  XOR U67597 ( .A(n55094), .B(n55095), .Z(n58666) );
  XOR U67598 ( .A(n58665), .B(n58666), .Z(n58670) );
  XOR U67599 ( .A(n58668), .B(n58670), .Z(n55045) );
  NOR U67600 ( .A(n55046), .B(n55045), .Z(n55093) );
  XOR U67601 ( .A(n54912), .B(n54911), .Z(n55050) );
  NOR U67602 ( .A(n54914), .B(n54913), .Z(n54915) );
  XOR U67603 ( .A(n54916), .B(n54915), .Z(n54917) );
  IV U67604 ( .A(n54917), .Z(n54949) );
  XOR U67605 ( .A(n54919), .B(n54918), .Z(n54975) );
  NOR U67606 ( .A(n54972), .B(n54975), .Z(n54920) );
  IV U67607 ( .A(n54920), .Z(n54963) );
  IV U67608 ( .A(n54921), .Z(n54925) );
  NOR U67609 ( .A(n54923), .B(n54922), .Z(n54924) );
  XOR U67610 ( .A(n54925), .B(n54924), .Z(n54978) );
  XOR U67611 ( .A(n54927), .B(n54926), .Z(n54951) );
  IV U67612 ( .A(n54928), .Z(n54931) );
  NOR U67613 ( .A(n54929), .B(n54944), .Z(n54930) );
  XOR U67614 ( .A(n54931), .B(n54930), .Z(n54981) );
  IV U67615 ( .A(n54932), .Z(n54934) );
  NOR U67616 ( .A(n54934), .B(n54933), .Z(n54980) );
  IV U67617 ( .A(n54980), .Z(n54935) );
  NOR U67618 ( .A(n54981), .B(n54935), .Z(n54936) );
  NOR U67619 ( .A(n54937), .B(n54936), .Z(n54954) );
  NOR U67620 ( .A(n54939), .B(n54938), .Z(n54940) );
  XOR U67621 ( .A(n54941), .B(n54940), .Z(n54953) );
  NOR U67622 ( .A(n54954), .B(n54953), .Z(n54942) );
  IV U67623 ( .A(n54942), .Z(n54943) );
  NOR U67624 ( .A(n54944), .B(n54943), .Z(n54952) );
  IV U67625 ( .A(n54952), .Z(n54945) );
  NOR U67626 ( .A(n54951), .B(n54945), .Z(n54977) );
  IV U67627 ( .A(n54977), .Z(n54946) );
  NOR U67628 ( .A(n54978), .B(n54946), .Z(n54968) );
  IV U67629 ( .A(n54968), .Z(n54947) );
  NOR U67630 ( .A(n54963), .B(n54947), .Z(n54950) );
  IV U67631 ( .A(n54950), .Z(n54948) );
  NOR U67632 ( .A(n54949), .B(n54948), .Z(n55049) );
  IV U67633 ( .A(n55049), .Z(n55047) );
  XOR U67634 ( .A(n55050), .B(n55047), .Z(n55062) );
  XOR U67635 ( .A(n54950), .B(n54949), .Z(n54965) );
  XOR U67636 ( .A(n54952), .B(n54951), .Z(n55016) );
  XOR U67637 ( .A(n54954), .B(n54953), .Z(n55008) );
  IV U67638 ( .A(n55008), .Z(n54988) );
  IV U67639 ( .A(n54955), .Z(n54957) );
  NOR U67640 ( .A(n54957), .B(n54956), .Z(n54979) );
  IV U67641 ( .A(n54979), .Z(n54958) );
  NOR U67642 ( .A(n54981), .B(n54958), .Z(n55006) );
  IV U67643 ( .A(n55006), .Z(n54959) );
  NOR U67644 ( .A(n54988), .B(n54959), .Z(n54960) );
  IV U67645 ( .A(n54960), .Z(n54989) );
  NOR U67646 ( .A(n55016), .B(n54989), .Z(n55001) );
  IV U67647 ( .A(n55001), .Z(n54961) );
  NOR U67648 ( .A(n54978), .B(n54961), .Z(n54967) );
  IV U67649 ( .A(n54967), .Z(n54962) );
  NOR U67650 ( .A(n54963), .B(n54962), .Z(n54966) );
  IV U67651 ( .A(n54966), .Z(n54964) );
  NOR U67652 ( .A(n54965), .B(n54964), .Z(n55051) );
  XOR U67653 ( .A(n54966), .B(n54965), .Z(n55020) );
  NOR U67654 ( .A(n54968), .B(n54967), .Z(n54974) );
  NOR U67655 ( .A(n54974), .B(n54975), .Z(n54969) );
  NOR U67656 ( .A(n54970), .B(n54969), .Z(n54971) );
  XOR U67657 ( .A(n54972), .B(n54971), .Z(n54973) );
  IV U67658 ( .A(n54973), .Z(n55024) );
  XOR U67659 ( .A(n54975), .B(n54974), .Z(n54976) );
  IV U67660 ( .A(n54976), .Z(n54998) );
  XOR U67661 ( .A(n54978), .B(n54977), .Z(n55003) );
  NOR U67662 ( .A(n54980), .B(n54979), .Z(n54982) );
  XOR U67663 ( .A(n54982), .B(n54981), .Z(n55037) );
  IV U67664 ( .A(n55037), .Z(n55013) );
  IV U67665 ( .A(n54983), .Z(n54985) );
  NOR U67666 ( .A(n54985), .B(n54984), .Z(n55035) );
  IV U67667 ( .A(n55035), .Z(n54986) );
  NOR U67668 ( .A(n55013), .B(n54986), .Z(n55005) );
  IV U67669 ( .A(n55005), .Z(n54987) );
  NOR U67670 ( .A(n54988), .B(n54987), .Z(n55026) );
  IV U67671 ( .A(n55026), .Z(n54991) );
  XOR U67672 ( .A(n54989), .B(n55016), .Z(n55028) );
  IV U67673 ( .A(n55028), .Z(n54990) );
  NOR U67674 ( .A(n54991), .B(n54990), .Z(n55000) );
  IV U67675 ( .A(n55000), .Z(n54992) );
  NOR U67676 ( .A(n55003), .B(n54992), .Z(n54999) );
  IV U67677 ( .A(n54999), .Z(n54993) );
  NOR U67678 ( .A(n54998), .B(n54993), .Z(n55023) );
  IV U67679 ( .A(n55023), .Z(n54994) );
  NOR U67680 ( .A(n55024), .B(n54994), .Z(n55021) );
  IV U67681 ( .A(n55021), .Z(n54995) );
  NOR U67682 ( .A(n55020), .B(n54995), .Z(n55060) );
  NOR U67683 ( .A(n55051), .B(n55060), .Z(n54996) );
  XOR U67684 ( .A(n55062), .B(n54996), .Z(n54997) );
  IV U67685 ( .A(n54997), .Z(n58716) );
  XOR U67686 ( .A(n54999), .B(n54998), .Z(n58705) );
  NOR U67687 ( .A(n55001), .B(n55000), .Z(n55002) );
  XOR U67688 ( .A(n55003), .B(n55002), .Z(n55004) );
  IV U67689 ( .A(n55004), .Z(n55030) );
  NOR U67690 ( .A(n55006), .B(n55005), .Z(n55007) );
  XOR U67691 ( .A(n55008), .B(n55007), .Z(n55070) );
  IV U67692 ( .A(n55009), .Z(n55011) );
  NOR U67693 ( .A(n55011), .B(n55010), .Z(n55034) );
  IV U67694 ( .A(n55034), .Z(n55012) );
  NOR U67695 ( .A(n55013), .B(n55012), .Z(n55069) );
  IV U67696 ( .A(n55069), .Z(n55014) );
  NOR U67697 ( .A(n55070), .B(n55014), .Z(n55025) );
  IV U67698 ( .A(n55025), .Z(n55015) );
  NOR U67699 ( .A(n55016), .B(n55015), .Z(n55029) );
  IV U67700 ( .A(n55029), .Z(n55017) );
  NOR U67701 ( .A(n55030), .B(n55017), .Z(n58704) );
  IV U67702 ( .A(n58704), .Z(n55018) );
  NOR U67703 ( .A(n58705), .B(n55018), .Z(n55019) );
  IV U67704 ( .A(n55019), .Z(n55081) );
  NOR U67705 ( .A(n55024), .B(n55081), .Z(n55086) );
  XOR U67706 ( .A(n55021), .B(n55020), .Z(n55066) );
  XOR U67707 ( .A(n55086), .B(n55066), .Z(n58711) );
  NOR U67708 ( .A(n58716), .B(n58711), .Z(n55022) );
  IV U67709 ( .A(n55022), .Z(n55090) );
  XOR U67710 ( .A(n55024), .B(n55023), .Z(n55080) );
  NOR U67711 ( .A(n55026), .B(n55025), .Z(n55027) );
  XOR U67712 ( .A(n55028), .B(n55027), .Z(n58699) );
  XOR U67713 ( .A(n55030), .B(n55029), .Z(n58702) );
  NOR U67714 ( .A(n58699), .B(n58702), .Z(n55031) );
  IV U67715 ( .A(n55031), .Z(n55032) );
  NOR U67716 ( .A(n58705), .B(n55032), .Z(n55033) );
  IV U67717 ( .A(n55033), .Z(n55078) );
  NOR U67718 ( .A(n55035), .B(n55034), .Z(n55036) );
  XOR U67719 ( .A(n55037), .B(n55036), .Z(n58693) );
  IV U67720 ( .A(n55038), .Z(n55040) );
  NOR U67721 ( .A(n55040), .B(n55039), .Z(n58691) );
  IV U67722 ( .A(n58691), .Z(n55041) );
  NOR U67723 ( .A(n58693), .B(n55041), .Z(n55068) );
  IV U67724 ( .A(n55068), .Z(n55042) );
  NOR U67725 ( .A(n55070), .B(n55042), .Z(n58697) );
  IV U67726 ( .A(n58697), .Z(n55043) );
  NOR U67727 ( .A(n55078), .B(n55043), .Z(n55082) );
  IV U67728 ( .A(n55082), .Z(n55079) );
  NOR U67729 ( .A(n55080), .B(n55079), .Z(n58710) );
  IV U67730 ( .A(n58710), .Z(n55044) );
  NOR U67731 ( .A(n55090), .B(n55044), .Z(n55108) );
  XOR U67732 ( .A(n55046), .B(n55045), .Z(n55059) );
  IV U67733 ( .A(n55059), .Z(n55056) );
  IV U67734 ( .A(n55050), .Z(n55048) );
  NOR U67735 ( .A(n55048), .B(n55047), .Z(n55055) );
  NOR U67736 ( .A(n55050), .B(n55049), .Z(n55053) );
  IV U67737 ( .A(n55051), .Z(n55052) );
  NOR U67738 ( .A(n55053), .B(n55052), .Z(n55054) );
  NOR U67739 ( .A(n55055), .B(n55054), .Z(n55057) );
  NOR U67740 ( .A(n55056), .B(n55057), .Z(n55101) );
  IV U67741 ( .A(n55057), .Z(n55058) );
  NOR U67742 ( .A(n55059), .B(n55058), .Z(n55098) );
  IV U67743 ( .A(n55060), .Z(n55061) );
  NOR U67744 ( .A(n55062), .B(n55061), .Z(n55097) );
  XOR U67745 ( .A(n55098), .B(n55097), .Z(n55063) );
  NOR U67746 ( .A(n55101), .B(n55063), .Z(n55064) );
  IV U67747 ( .A(n55064), .Z(n55107) );
  IV U67748 ( .A(n55086), .Z(n55065) );
  NOR U67749 ( .A(n55066), .B(n55065), .Z(n58714) );
  IV U67750 ( .A(n58714), .Z(n55067) );
  NOR U67751 ( .A(n58716), .B(n55067), .Z(n55105) );
  XOR U67752 ( .A(n55107), .B(n55105), .Z(n55110) );
  XOR U67753 ( .A(n55108), .B(n55110), .Z(n58718) );
  NOR U67754 ( .A(n55069), .B(n55068), .Z(n55071) );
  XOR U67755 ( .A(n55071), .B(n55070), .Z(n55072) );
  IV U67756 ( .A(n55072), .Z(n58695) );
  NOR U67757 ( .A(n55074), .B(n55073), .Z(n58690) );
  IV U67758 ( .A(n58690), .Z(n55075) );
  NOR U67759 ( .A(n58693), .B(n55075), .Z(n55076) );
  IV U67760 ( .A(n55076), .Z(n58694) );
  NOR U67761 ( .A(n58695), .B(n58694), .Z(n58696) );
  IV U67762 ( .A(n58696), .Z(n55077) );
  NOR U67763 ( .A(n55078), .B(n55077), .Z(n58708) );
  IV U67764 ( .A(n58708), .Z(n55088) );
  XOR U67765 ( .A(n55080), .B(n55079), .Z(n55084) );
  NOR U67766 ( .A(n55082), .B(n55081), .Z(n55083) );
  NOR U67767 ( .A(n55084), .B(n55083), .Z(n55085) );
  NOR U67768 ( .A(n55086), .B(n55085), .Z(n58707) );
  IV U67769 ( .A(n58707), .Z(n55087) );
  NOR U67770 ( .A(n55088), .B(n55087), .Z(n58709) );
  IV U67771 ( .A(n58709), .Z(n55089) );
  NOR U67772 ( .A(n55090), .B(n55089), .Z(n55091) );
  IV U67773 ( .A(n55091), .Z(n58717) );
  NOR U67774 ( .A(n58718), .B(n58717), .Z(n55092) );
  NOR U67775 ( .A(n55093), .B(n55092), .Z(n58689) );
  IV U67776 ( .A(n55094), .Z(n55096) );
  NOR U67777 ( .A(n55096), .B(n55095), .Z(n55104) );
  IV U67778 ( .A(n55097), .Z(n55099) );
  NOR U67779 ( .A(n55099), .B(n55098), .Z(n55100) );
  NOR U67780 ( .A(n55101), .B(n55100), .Z(n55102) );
  IV U67781 ( .A(n55102), .Z(n55103) );
  NOR U67782 ( .A(n55104), .B(n55103), .Z(n58687) );
  IV U67783 ( .A(n55105), .Z(n55106) );
  NOR U67784 ( .A(n55107), .B(n55106), .Z(n55112) );
  IV U67785 ( .A(n55108), .Z(n55109) );
  NOR U67786 ( .A(n55110), .B(n55109), .Z(n55111) );
  NOR U67787 ( .A(n55112), .B(n55111), .Z(n58685) );
  IV U67788 ( .A(n55113), .Z(n55114) );
  NOR U67789 ( .A(n55115), .B(n55114), .Z(n55120) );
  IV U67790 ( .A(n55116), .Z(n55118) );
  NOR U67791 ( .A(n55118), .B(n55117), .Z(n55119) );
  NOR U67792 ( .A(n55120), .B(n55119), .Z(n58664) );
  IV U67793 ( .A(n55121), .Z(n55122) );
  NOR U67794 ( .A(n55123), .B(n55122), .Z(n55128) );
  IV U67795 ( .A(n55124), .Z(n55126) );
  NOR U67796 ( .A(n55126), .B(n55125), .Z(n55127) );
  NOR U67797 ( .A(n55128), .B(n55127), .Z(n58646) );
  IV U67798 ( .A(n55129), .Z(n55130) );
  NOR U67799 ( .A(n55131), .B(n55130), .Z(n55136) );
  IV U67800 ( .A(n55132), .Z(n55139) );
  IV U67801 ( .A(n55133), .Z(n55134) );
  NOR U67802 ( .A(n55139), .B(n55134), .Z(n55135) );
  NOR U67803 ( .A(n55136), .B(n55135), .Z(n58644) );
  IV U67804 ( .A(n55137), .Z(n55138) );
  NOR U67805 ( .A(n55139), .B(n55138), .Z(n58633) );
  IV U67806 ( .A(n55140), .Z(n55142) );
  NOR U67807 ( .A(n55142), .B(n55141), .Z(n55146) );
  NOR U67808 ( .A(n55144), .B(n55143), .Z(n55145) );
  NOR U67809 ( .A(n55146), .B(n55145), .Z(n58631) );
  IV U67810 ( .A(n55147), .Z(n55149) );
  NOR U67811 ( .A(n55149), .B(n55148), .Z(n55153) );
  NOR U67812 ( .A(n55151), .B(n55150), .Z(n55152) );
  NOR U67813 ( .A(n55153), .B(n55152), .Z(n55168) );
  NOR U67814 ( .A(n55155), .B(n55154), .Z(n55166) );
  IV U67815 ( .A(n55156), .Z(n55158) );
  NOR U67816 ( .A(n55158), .B(n55157), .Z(n55163) );
  IV U67817 ( .A(n55159), .Z(n55160) );
  NOR U67818 ( .A(n55161), .B(n55160), .Z(n55162) );
  NOR U67819 ( .A(n55163), .B(n55162), .Z(n55164) );
  IV U67820 ( .A(n55164), .Z(n55165) );
  NOR U67821 ( .A(n55166), .B(n55165), .Z(n55167) );
  XOR U67822 ( .A(n55168), .B(n55167), .Z(n58629) );
  NOR U67823 ( .A(n55170), .B(n55169), .Z(n55179) );
  IV U67824 ( .A(n55170), .Z(n55172) );
  NOR U67825 ( .A(n55172), .B(n55171), .Z(n55177) );
  NOR U67826 ( .A(n55174), .B(n55173), .Z(n55175) );
  IV U67827 ( .A(n55175), .Z(n55176) );
  NOR U67828 ( .A(n55177), .B(n55176), .Z(n55178) );
  NOR U67829 ( .A(n55179), .B(n55178), .Z(n55188) );
  IV U67830 ( .A(n55180), .Z(n55182) );
  NOR U67831 ( .A(n55182), .B(n55181), .Z(n55186) );
  NOR U67832 ( .A(n55184), .B(n55183), .Z(n55185) );
  NOR U67833 ( .A(n55186), .B(n55185), .Z(n55187) );
  XOR U67834 ( .A(n55188), .B(n55187), .Z(n58512) );
  IV U67835 ( .A(n55189), .Z(n55191) );
  NOR U67836 ( .A(n55191), .B(n55190), .Z(n55196) );
  IV U67837 ( .A(n55192), .Z(n55194) );
  NOR U67838 ( .A(n55194), .B(n55193), .Z(n55195) );
  NOR U67839 ( .A(n55196), .B(n55195), .Z(n55206) );
  IV U67840 ( .A(n55197), .Z(n55198) );
  NOR U67841 ( .A(n55199), .B(n55198), .Z(n55204) );
  IV U67842 ( .A(n55200), .Z(n55202) );
  NOR U67843 ( .A(n55202), .B(n55201), .Z(n55203) );
  NOR U67844 ( .A(n55204), .B(n55203), .Z(n55205) );
  XOR U67845 ( .A(n55206), .B(n55205), .Z(n55238) );
  IV U67846 ( .A(n55207), .Z(n55209) );
  NOR U67847 ( .A(n55209), .B(n55208), .Z(n55213) );
  NOR U67848 ( .A(n55211), .B(n55210), .Z(n55212) );
  NOR U67849 ( .A(n55213), .B(n55212), .Z(n55226) );
  IV U67850 ( .A(n55214), .Z(n55216) );
  NOR U67851 ( .A(n55216), .B(n55215), .Z(n55218) );
  NOR U67852 ( .A(n55218), .B(n55217), .Z(n55219) );
  IV U67853 ( .A(n55219), .Z(n55224) );
  IV U67854 ( .A(n55220), .Z(n55221) );
  NOR U67855 ( .A(n55222), .B(n55221), .Z(n55223) );
  NOR U67856 ( .A(n55224), .B(n55223), .Z(n55225) );
  XOR U67857 ( .A(n55226), .B(n55225), .Z(n55236) );
  IV U67858 ( .A(n55227), .Z(n55229) );
  NOR U67859 ( .A(n55229), .B(n55228), .Z(n55234) );
  IV U67860 ( .A(n55230), .Z(n55232) );
  NOR U67861 ( .A(n55232), .B(n55231), .Z(n55233) );
  NOR U67862 ( .A(n55234), .B(n55233), .Z(n55235) );
  XOR U67863 ( .A(n55236), .B(n55235), .Z(n55237) );
  XOR U67864 ( .A(n55238), .B(n55237), .Z(n58455) );
  IV U67865 ( .A(n55239), .Z(n55240) );
  NOR U67866 ( .A(n55241), .B(n55240), .Z(n55246) );
  IV U67867 ( .A(n55242), .Z(n55244) );
  NOR U67868 ( .A(n55244), .B(n55243), .Z(n55245) );
  NOR U67869 ( .A(n55246), .B(n55245), .Z(n58453) );
  IV U67870 ( .A(n55247), .Z(n55250) );
  IV U67871 ( .A(n55248), .Z(n55249) );
  NOR U67872 ( .A(n55250), .B(n55249), .Z(n55254) );
  IV U67873 ( .A(n55251), .Z(n55252) );
  NOR U67874 ( .A(n55272), .B(n55252), .Z(n55253) );
  NOR U67875 ( .A(n55254), .B(n55253), .Z(n58451) );
  IV U67876 ( .A(n55255), .Z(n55257) );
  NOR U67877 ( .A(n55257), .B(n55256), .Z(n55262) );
  IV U67878 ( .A(n55258), .Z(n55260) );
  NOR U67879 ( .A(n55260), .B(n55259), .Z(n55261) );
  NOR U67880 ( .A(n55262), .B(n55261), .Z(n58449) );
  IV U67881 ( .A(n55263), .Z(n55265) );
  NOR U67882 ( .A(n55265), .B(n55264), .Z(n55270) );
  IV U67883 ( .A(n55266), .Z(n55268) );
  NOR U67884 ( .A(n55268), .B(n55267), .Z(n55269) );
  NOR U67885 ( .A(n55270), .B(n55269), .Z(n55280) );
  IV U67886 ( .A(n55271), .Z(n55273) );
  NOR U67887 ( .A(n55273), .B(n55272), .Z(n55278) );
  IV U67888 ( .A(n55274), .Z(n55276) );
  NOR U67889 ( .A(n55276), .B(n55275), .Z(n55277) );
  NOR U67890 ( .A(n55278), .B(n55277), .Z(n55279) );
  XOR U67891 ( .A(n55280), .B(n55279), .Z(n58447) );
  IV U67892 ( .A(n55281), .Z(n55283) );
  NOR U67893 ( .A(n55283), .B(n55282), .Z(n55287) );
  NOR U67894 ( .A(n55285), .B(n55284), .Z(n55286) );
  NOR U67895 ( .A(n55287), .B(n55286), .Z(n55300) );
  IV U67896 ( .A(n55288), .Z(n55290) );
  NOR U67897 ( .A(n55290), .B(n55289), .Z(n55292) );
  NOR U67898 ( .A(n55292), .B(n55291), .Z(n55293) );
  IV U67899 ( .A(n55293), .Z(n55298) );
  IV U67900 ( .A(n55294), .Z(n55295) );
  NOR U67901 ( .A(n55296), .B(n55295), .Z(n55297) );
  NOR U67902 ( .A(n55298), .B(n55297), .Z(n55299) );
  XOR U67903 ( .A(n55300), .B(n55299), .Z(n58445) );
  NOR U67904 ( .A(n55302), .B(n55301), .Z(n55305) );
  IV U67905 ( .A(n55303), .Z(n55304) );
  NOR U67906 ( .A(n55305), .B(n55304), .Z(n55320) );
  NOR U67907 ( .A(n55307), .B(n55306), .Z(n55318) );
  IV U67908 ( .A(n55308), .Z(n55309) );
  NOR U67909 ( .A(n55310), .B(n55309), .Z(n55315) );
  IV U67910 ( .A(n55311), .Z(n55313) );
  NOR U67911 ( .A(n55313), .B(n55312), .Z(n55314) );
  NOR U67912 ( .A(n55315), .B(n55314), .Z(n55316) );
  IV U67913 ( .A(n55316), .Z(n55317) );
  NOR U67914 ( .A(n55318), .B(n55317), .Z(n55319) );
  XOR U67915 ( .A(n55320), .B(n55319), .Z(n55331) );
  IV U67916 ( .A(n55321), .Z(n55322) );
  NOR U67917 ( .A(n55323), .B(n55322), .Z(n55329) );
  IV U67918 ( .A(n55324), .Z(n55327) );
  IV U67919 ( .A(n55325), .Z(n55326) );
  NOR U67920 ( .A(n55327), .B(n55326), .Z(n55328) );
  NOR U67921 ( .A(n55329), .B(n55328), .Z(n55330) );
  XOR U67922 ( .A(n55331), .B(n55330), .Z(n55369) );
  IV U67923 ( .A(n55332), .Z(n55335) );
  NOR U67924 ( .A(n55338), .B(n55333), .Z(n55334) );
  NOR U67925 ( .A(n55335), .B(n55334), .Z(n55345) );
  NOR U67926 ( .A(n55337), .B(n55336), .Z(n55342) );
  IV U67927 ( .A(n55338), .Z(n55340) );
  NOR U67928 ( .A(n55340), .B(n55339), .Z(n55341) );
  NOR U67929 ( .A(n55342), .B(n55341), .Z(n55343) );
  IV U67930 ( .A(n55343), .Z(n55344) );
  NOR U67931 ( .A(n55345), .B(n55344), .Z(n55357) );
  NOR U67932 ( .A(n55347), .B(n55346), .Z(n55348) );
  NOR U67933 ( .A(n55349), .B(n55348), .Z(n55355) );
  IV U67934 ( .A(n55350), .Z(n55353) );
  IV U67935 ( .A(n55351), .Z(n55352) );
  NOR U67936 ( .A(n55353), .B(n55352), .Z(n55354) );
  NOR U67937 ( .A(n55355), .B(n55354), .Z(n55356) );
  XOR U67938 ( .A(n55357), .B(n55356), .Z(n55367) );
  IV U67939 ( .A(n55358), .Z(n55359) );
  NOR U67940 ( .A(n55360), .B(n55359), .Z(n55365) );
  IV U67941 ( .A(n55361), .Z(n55362) );
  NOR U67942 ( .A(n55363), .B(n55362), .Z(n55364) );
  NOR U67943 ( .A(n55365), .B(n55364), .Z(n55366) );
  XOR U67944 ( .A(n55367), .B(n55366), .Z(n55368) );
  XOR U67945 ( .A(n55369), .B(n55368), .Z(n58443) );
  IV U67946 ( .A(n55370), .Z(n55372) );
  NOR U67947 ( .A(n55372), .B(n55371), .Z(n55377) );
  IV U67948 ( .A(n55373), .Z(n55374) );
  NOR U67949 ( .A(n55375), .B(n55374), .Z(n55376) );
  NOR U67950 ( .A(n55377), .B(n55376), .Z(n58441) );
  IV U67951 ( .A(n55378), .Z(n55379) );
  NOR U67952 ( .A(n55380), .B(n55379), .Z(n55396) );
  NOR U67953 ( .A(n55381), .B(n55382), .Z(n58406) );
  IV U67954 ( .A(n55382), .Z(n55383) );
  NOR U67955 ( .A(n55384), .B(n55383), .Z(n55385) );
  NOR U67956 ( .A(n55386), .B(n55385), .Z(n55387) );
  IV U67957 ( .A(n55387), .Z(n58403) );
  NOR U67958 ( .A(n58406), .B(n58403), .Z(n55388) );
  IV U67959 ( .A(n55388), .Z(n55394) );
  IV U67960 ( .A(n55389), .Z(n55390) );
  NOR U67961 ( .A(n55391), .B(n55390), .Z(n55392) );
  IV U67962 ( .A(n55392), .Z(n55393) );
  NOR U67963 ( .A(n55394), .B(n55393), .Z(n55395) );
  NOR U67964 ( .A(n55396), .B(n55395), .Z(n58439) );
  IV U67965 ( .A(n55397), .Z(n55398) );
  NOR U67966 ( .A(n55399), .B(n55398), .Z(n55404) );
  IV U67967 ( .A(n55400), .Z(n55401) );
  NOR U67968 ( .A(n55402), .B(n55401), .Z(n55403) );
  NOR U67969 ( .A(n55404), .B(n55403), .Z(n58437) );
  IV U67970 ( .A(n55405), .Z(n55407) );
  NOR U67971 ( .A(n55407), .B(n55406), .Z(n55412) );
  IV U67972 ( .A(n55408), .Z(n55409) );
  NOR U67973 ( .A(n55410), .B(n55409), .Z(n55411) );
  NOR U67974 ( .A(n55412), .B(n55411), .Z(n55422) );
  IV U67975 ( .A(n55413), .Z(n55414) );
  NOR U67976 ( .A(n55415), .B(n55414), .Z(n55420) );
  IV U67977 ( .A(n55416), .Z(n55418) );
  NOR U67978 ( .A(n55418), .B(n55417), .Z(n55419) );
  NOR U67979 ( .A(n55420), .B(n55419), .Z(n55421) );
  XOR U67980 ( .A(n55422), .B(n55421), .Z(n55428) );
  NOR U67981 ( .A(n55424), .B(n55423), .Z(n55426) );
  NOR U67982 ( .A(n55426), .B(n55425), .Z(n55427) );
  XOR U67983 ( .A(n55428), .B(n55427), .Z(n58400) );
  IV U67984 ( .A(n55429), .Z(n55431) );
  NOR U67985 ( .A(n55431), .B(n55430), .Z(n55437) );
  NOR U67986 ( .A(n55433), .B(n55432), .Z(n55434) );
  NOR U67987 ( .A(n55435), .B(n55434), .Z(n55436) );
  NOR U67988 ( .A(n55437), .B(n55436), .Z(n58398) );
  IV U67989 ( .A(n55438), .Z(n55442) );
  NOR U67990 ( .A(n55440), .B(n55439), .Z(n55441) );
  NOR U67991 ( .A(n55442), .B(n55441), .Z(n55450) );
  IV U67992 ( .A(n55443), .Z(n55445) );
  NOR U67993 ( .A(n55445), .B(n55444), .Z(n55447) );
  NOR U67994 ( .A(n55447), .B(n55446), .Z(n55448) );
  IV U67995 ( .A(n55448), .Z(n55449) );
  NOR U67996 ( .A(n55450), .B(n55449), .Z(n55456) );
  NOR U67997 ( .A(n55452), .B(n55451), .Z(n55453) );
  NOR U67998 ( .A(n55454), .B(n55453), .Z(n55455) );
  XOR U67999 ( .A(n55456), .B(n55455), .Z(n55465) );
  IV U68000 ( .A(n55457), .Z(n55458) );
  NOR U68001 ( .A(n55459), .B(n55458), .Z(n55463) );
  NOR U68002 ( .A(n55461), .B(n55460), .Z(n55462) );
  NOR U68003 ( .A(n55463), .B(n55462), .Z(n55464) );
  XOR U68004 ( .A(n55465), .B(n55464), .Z(n58396) );
  IV U68005 ( .A(n55466), .Z(n55468) );
  NOR U68006 ( .A(n55468), .B(n55467), .Z(n55473) );
  IV U68007 ( .A(n55469), .Z(n55471) );
  NOR U68008 ( .A(n55471), .B(n55470), .Z(n55472) );
  NOR U68009 ( .A(n55473), .B(n55472), .Z(n58394) );
  IV U68010 ( .A(n55474), .Z(n55475) );
  NOR U68011 ( .A(n55476), .B(n55475), .Z(n55486) );
  IV U68012 ( .A(n55477), .Z(n55478) );
  NOR U68013 ( .A(n55489), .B(n55478), .Z(n55484) );
  IV U68014 ( .A(n55479), .Z(n55482) );
  IV U68015 ( .A(n55480), .Z(n55481) );
  NOR U68016 ( .A(n55482), .B(n55481), .Z(n55483) );
  NOR U68017 ( .A(n55484), .B(n55483), .Z(n55485) );
  XOR U68018 ( .A(n55486), .B(n55485), .Z(n55493) );
  IV U68019 ( .A(n55487), .Z(n55488) );
  NOR U68020 ( .A(n55489), .B(n55488), .Z(n55491) );
  NOR U68021 ( .A(n55491), .B(n55490), .Z(n55492) );
  XOR U68022 ( .A(n55493), .B(n55492), .Z(n55512) );
  NOR U68023 ( .A(n55495), .B(n55494), .Z(n55500) );
  IV U68024 ( .A(n55496), .Z(n55497) );
  NOR U68025 ( .A(n55498), .B(n55497), .Z(n55499) );
  NOR U68026 ( .A(n55500), .B(n55499), .Z(n55510) );
  IV U68027 ( .A(n55501), .Z(n55503) );
  NOR U68028 ( .A(n55503), .B(n55502), .Z(n55508) );
  IV U68029 ( .A(n55504), .Z(n55505) );
  NOR U68030 ( .A(n55506), .B(n55505), .Z(n55507) );
  NOR U68031 ( .A(n55508), .B(n55507), .Z(n55509) );
  XOR U68032 ( .A(n55510), .B(n55509), .Z(n55511) );
  XOR U68033 ( .A(n55512), .B(n55511), .Z(n58392) );
  IV U68034 ( .A(n55513), .Z(n55515) );
  NOR U68035 ( .A(n55515), .B(n55514), .Z(n55520) );
  IV U68036 ( .A(n55516), .Z(n55518) );
  NOR U68037 ( .A(n55518), .B(n55517), .Z(n55519) );
  NOR U68038 ( .A(n55520), .B(n55519), .Z(n58324) );
  IV U68039 ( .A(n55521), .Z(n55522) );
  NOR U68040 ( .A(n55522), .B(n55567), .Z(n55527) );
  IV U68041 ( .A(n55523), .Z(n55524) );
  NOR U68042 ( .A(n55525), .B(n55524), .Z(n55526) );
  NOR U68043 ( .A(n55527), .B(n55526), .Z(n58303) );
  NOR U68044 ( .A(n55529), .B(n55528), .Z(n55534) );
  IV U68045 ( .A(n55530), .Z(n55531) );
  NOR U68046 ( .A(n55532), .B(n55531), .Z(n55533) );
  NOR U68047 ( .A(n55534), .B(n55533), .Z(n55543) );
  IV U68048 ( .A(n55535), .Z(n55537) );
  NOR U68049 ( .A(n55537), .B(n55536), .Z(n55541) );
  NOR U68050 ( .A(n55539), .B(n55538), .Z(n55540) );
  NOR U68051 ( .A(n55541), .B(n55540), .Z(n55542) );
  XOR U68052 ( .A(n55543), .B(n55542), .Z(n55556) );
  IV U68053 ( .A(n55544), .Z(n55545) );
  NOR U68054 ( .A(n55546), .B(n55545), .Z(n55554) );
  IV U68055 ( .A(n55547), .Z(n55549) );
  NOR U68056 ( .A(n55549), .B(n55548), .Z(n55551) );
  NOR U68057 ( .A(n55551), .B(n55550), .Z(n55552) );
  IV U68058 ( .A(n55552), .Z(n55553) );
  NOR U68059 ( .A(n55554), .B(n55553), .Z(n55555) );
  XOR U68060 ( .A(n55556), .B(n55555), .Z(n55573) );
  IV U68061 ( .A(n55557), .Z(n55559) );
  NOR U68062 ( .A(n55559), .B(n55558), .Z(n55564) );
  IV U68063 ( .A(n55560), .Z(n55561) );
  NOR U68064 ( .A(n55562), .B(n55561), .Z(n55563) );
  NOR U68065 ( .A(n55564), .B(n55563), .Z(n55571) );
  IV U68066 ( .A(n55565), .Z(n55566) );
  NOR U68067 ( .A(n55567), .B(n55566), .Z(n55569) );
  NOR U68068 ( .A(n55569), .B(n55568), .Z(n55570) );
  XOR U68069 ( .A(n55571), .B(n55570), .Z(n55572) );
  XOR U68070 ( .A(n55573), .B(n55572), .Z(n58272) );
  IV U68071 ( .A(n55574), .Z(n55576) );
  NOR U68072 ( .A(n55576), .B(n55575), .Z(n55581) );
  IV U68073 ( .A(n55577), .Z(n55579) );
  NOR U68074 ( .A(n55579), .B(n55578), .Z(n55580) );
  NOR U68075 ( .A(n55581), .B(n55580), .Z(n58270) );
  NOR U68076 ( .A(n55583), .B(n55582), .Z(n55602) );
  IV U68077 ( .A(n55584), .Z(n55586) );
  NOR U68078 ( .A(n55586), .B(n55585), .Z(n55590) );
  NOR U68079 ( .A(n55588), .B(n55587), .Z(n55589) );
  NOR U68080 ( .A(n55590), .B(n55589), .Z(n55600) );
  IV U68081 ( .A(n55591), .Z(n55593) );
  NOR U68082 ( .A(n55593), .B(n55592), .Z(n55598) );
  IV U68083 ( .A(n55594), .Z(n55596) );
  NOR U68084 ( .A(n55596), .B(n55595), .Z(n55597) );
  NOR U68085 ( .A(n55598), .B(n55597), .Z(n55599) );
  XOR U68086 ( .A(n55600), .B(n55599), .Z(n55601) );
  XOR U68087 ( .A(n55602), .B(n55601), .Z(n55622) );
  IV U68088 ( .A(n55603), .Z(n55605) );
  NOR U68089 ( .A(n55605), .B(n55604), .Z(n55610) );
  IV U68090 ( .A(n55606), .Z(n55607) );
  NOR U68091 ( .A(n55608), .B(n55607), .Z(n55609) );
  NOR U68092 ( .A(n55610), .B(n55609), .Z(n55620) );
  IV U68093 ( .A(n55611), .Z(n55613) );
  NOR U68094 ( .A(n55613), .B(n55612), .Z(n55618) );
  IV U68095 ( .A(n55614), .Z(n55616) );
  NOR U68096 ( .A(n55616), .B(n55615), .Z(n55617) );
  NOR U68097 ( .A(n55618), .B(n55617), .Z(n55619) );
  XOR U68098 ( .A(n55620), .B(n55619), .Z(n55621) );
  XOR U68099 ( .A(n55622), .B(n55621), .Z(n58268) );
  IV U68100 ( .A(n55623), .Z(n55624) );
  NOR U68101 ( .A(n55625), .B(n55624), .Z(n55636) );
  IV U68102 ( .A(n55626), .Z(n55627) );
  NOR U68103 ( .A(n55628), .B(n55627), .Z(n55633) );
  IV U68104 ( .A(n55629), .Z(n55630) );
  NOR U68105 ( .A(n55631), .B(n55630), .Z(n55632) );
  NOR U68106 ( .A(n55633), .B(n55632), .Z(n55634) );
  IV U68107 ( .A(n55634), .Z(n55635) );
  NOR U68108 ( .A(n55636), .B(n55635), .Z(n58266) );
  NOR U68109 ( .A(n55638), .B(n55637), .Z(n55641) );
  IV U68110 ( .A(n55639), .Z(n55640) );
  NOR U68111 ( .A(n55641), .B(n55640), .Z(n55645) );
  NOR U68112 ( .A(n55643), .B(n55642), .Z(n55644) );
  NOR U68113 ( .A(n55645), .B(n55644), .Z(n55655) );
  NOR U68114 ( .A(n55647), .B(n55646), .Z(n55653) );
  NOR U68115 ( .A(n55649), .B(n55648), .Z(n55650) );
  NOR U68116 ( .A(n55651), .B(n55650), .Z(n55652) );
  NOR U68117 ( .A(n55653), .B(n55652), .Z(n55654) );
  XOR U68118 ( .A(n55655), .B(n55654), .Z(n58238) );
  IV U68119 ( .A(n55656), .Z(n55666) );
  NOR U68120 ( .A(n55657), .B(n55666), .Z(n55662) );
  IV U68121 ( .A(n55658), .Z(n55660) );
  NOR U68122 ( .A(n55660), .B(n55659), .Z(n55661) );
  NOR U68123 ( .A(n55662), .B(n55661), .Z(n55671) );
  NOR U68124 ( .A(n55664), .B(n55663), .Z(n55669) );
  IV U68125 ( .A(n55665), .Z(n55667) );
  NOR U68126 ( .A(n55667), .B(n55666), .Z(n55668) );
  NOR U68127 ( .A(n55669), .B(n55668), .Z(n55670) );
  XOR U68128 ( .A(n55671), .B(n55670), .Z(n55681) );
  NOR U68129 ( .A(n55672), .B(n55673), .Z(n55679) );
  IV U68130 ( .A(n55673), .Z(n55674) );
  NOR U68131 ( .A(n55675), .B(n55674), .Z(n55676) );
  NOR U68132 ( .A(n55677), .B(n55676), .Z(n55678) );
  NOR U68133 ( .A(n55679), .B(n55678), .Z(n55680) );
  XOR U68134 ( .A(n55681), .B(n55680), .Z(n58236) );
  IV U68135 ( .A(n55685), .Z(n55683) );
  NOR U68136 ( .A(n55683), .B(n55682), .Z(n55690) );
  NOR U68137 ( .A(n55685), .B(n55684), .Z(n55688) );
  IV U68138 ( .A(n55686), .Z(n55687) );
  NOR U68139 ( .A(n55688), .B(n55687), .Z(n55689) );
  NOR U68140 ( .A(n55690), .B(n55689), .Z(n58175) );
  NOR U68141 ( .A(n55692), .B(n55691), .Z(n55703) );
  IV U68142 ( .A(n55693), .Z(n55695) );
  NOR U68143 ( .A(n55695), .B(n55694), .Z(n55700) );
  IV U68144 ( .A(n55696), .Z(n55698) );
  NOR U68145 ( .A(n55698), .B(n55697), .Z(n55699) );
  NOR U68146 ( .A(n55700), .B(n55699), .Z(n55701) );
  IV U68147 ( .A(n55701), .Z(n55702) );
  NOR U68148 ( .A(n55703), .B(n55702), .Z(n55726) );
  IV U68149 ( .A(n55704), .Z(n55776) );
  IV U68150 ( .A(n55705), .Z(n55706) );
  NOR U68151 ( .A(n55776), .B(n55706), .Z(n55711) );
  IV U68152 ( .A(n55707), .Z(n55708) );
  NOR U68153 ( .A(n55709), .B(n55708), .Z(n55710) );
  NOR U68154 ( .A(n55711), .B(n55710), .Z(n55724) );
  NOR U68155 ( .A(n55713), .B(n55712), .Z(n55720) );
  XOR U68156 ( .A(n55714), .B(n55720), .Z(n55722) );
  IV U68157 ( .A(n55715), .Z(n55716) );
  NOR U68158 ( .A(n55717), .B(n55716), .Z(n55718) );
  IV U68159 ( .A(n55718), .Z(n55719) );
  NOR U68160 ( .A(n55720), .B(n55719), .Z(n55721) );
  NOR U68161 ( .A(n55722), .B(n55721), .Z(n55723) );
  XOR U68162 ( .A(n55724), .B(n55723), .Z(n55725) );
  XOR U68163 ( .A(n55726), .B(n55725), .Z(n58137) );
  NOR U68164 ( .A(n55728), .B(n55727), .Z(n55730) );
  NOR U68165 ( .A(n55730), .B(n55729), .Z(n58135) );
  IV U68166 ( .A(n55731), .Z(n55732) );
  NOR U68167 ( .A(n55733), .B(n55732), .Z(n55738) );
  IV U68168 ( .A(n55734), .Z(n55736) );
  NOR U68169 ( .A(n55736), .B(n55735), .Z(n55737) );
  NOR U68170 ( .A(n55738), .B(n55737), .Z(n55747) );
  IV U68171 ( .A(n55739), .Z(n55740) );
  NOR U68172 ( .A(n55741), .B(n55740), .Z(n55745) );
  NOR U68173 ( .A(n55743), .B(n55742), .Z(n55744) );
  NOR U68174 ( .A(n55745), .B(n55744), .Z(n55746) );
  XOR U68175 ( .A(n55747), .B(n55746), .Z(n55762) );
  IV U68176 ( .A(n55748), .Z(n55749) );
  NOR U68177 ( .A(n55749), .B(n55754), .Z(n55760) );
  IV U68178 ( .A(n55750), .Z(n55751) );
  NOR U68179 ( .A(n55752), .B(n55751), .Z(n55757) );
  IV U68180 ( .A(n55753), .Z(n55755) );
  NOR U68181 ( .A(n55755), .B(n55754), .Z(n55756) );
  NOR U68182 ( .A(n55757), .B(n55756), .Z(n55758) );
  IV U68183 ( .A(n55758), .Z(n55759) );
  NOR U68184 ( .A(n55760), .B(n55759), .Z(n55761) );
  XOR U68185 ( .A(n55762), .B(n55761), .Z(n55797) );
  IV U68186 ( .A(n55766), .Z(n55763) );
  NOR U68187 ( .A(n55764), .B(n55763), .Z(n55773) );
  NOR U68188 ( .A(n55766), .B(n55765), .Z(n55771) );
  NOR U68189 ( .A(n55768), .B(n55767), .Z(n55769) );
  IV U68190 ( .A(n55769), .Z(n55770) );
  NOR U68191 ( .A(n55771), .B(n55770), .Z(n55772) );
  NOR U68192 ( .A(n55773), .B(n55772), .Z(n55783) );
  IV U68193 ( .A(n55774), .Z(n55775) );
  NOR U68194 ( .A(n55776), .B(n55775), .Z(n55781) );
  IV U68195 ( .A(n55777), .Z(n55778) );
  NOR U68196 ( .A(n55779), .B(n55778), .Z(n55780) );
  NOR U68197 ( .A(n55781), .B(n55780), .Z(n55782) );
  XOR U68198 ( .A(n55783), .B(n55782), .Z(n55795) );
  IV U68199 ( .A(n55784), .Z(n55786) );
  NOR U68200 ( .A(n55786), .B(n55785), .Z(n55793) );
  NOR U68201 ( .A(n55788), .B(n55787), .Z(n55790) );
  NOR U68202 ( .A(n55790), .B(n55789), .Z(n55791) );
  IV U68203 ( .A(n55791), .Z(n55792) );
  NOR U68204 ( .A(n55793), .B(n55792), .Z(n55794) );
  XOR U68205 ( .A(n55795), .B(n55794), .Z(n55796) );
  XOR U68206 ( .A(n55797), .B(n55796), .Z(n58133) );
  IV U68207 ( .A(n55798), .Z(n55800) );
  NOR U68208 ( .A(n55800), .B(n55799), .Z(n55805) );
  IV U68209 ( .A(n55801), .Z(n55803) );
  NOR U68210 ( .A(n55803), .B(n55802), .Z(n55804) );
  NOR U68211 ( .A(n55805), .B(n55804), .Z(n58107) );
  NOR U68212 ( .A(n55811), .B(n55810), .Z(n55812) );
  NOR U68213 ( .A(n55813), .B(n55812), .Z(n55823) );
  IV U68214 ( .A(n55814), .Z(n58065) );
  IV U68215 ( .A(n55815), .Z(n58064) );
  XOR U68216 ( .A(n58065), .B(n58064), .Z(n55816) );
  NOR U68217 ( .A(n55817), .B(n55816), .Z(n55821) );
  NOR U68218 ( .A(n55819), .B(n55818), .Z(n55820) );
  NOR U68219 ( .A(n55821), .B(n55820), .Z(n55822) );
  XOR U68220 ( .A(n55823), .B(n55822), .Z(n55850) );
  IV U68221 ( .A(n55827), .Z(n55824) );
  NOR U68222 ( .A(n55825), .B(n55824), .Z(n55835) );
  IV U68223 ( .A(n55825), .Z(n55826) );
  NOR U68224 ( .A(n55827), .B(n55826), .Z(n55833) );
  IV U68225 ( .A(n55828), .Z(n55829) );
  NOR U68226 ( .A(n55830), .B(n55829), .Z(n55831) );
  IV U68227 ( .A(n55831), .Z(n55832) );
  NOR U68228 ( .A(n55833), .B(n55832), .Z(n55834) );
  NOR U68229 ( .A(n55835), .B(n55834), .Z(n55848) );
  NOR U68230 ( .A(n55837), .B(n55836), .Z(n55846) );
  IV U68231 ( .A(n55838), .Z(n55840) );
  NOR U68232 ( .A(n55840), .B(n55839), .Z(n55841) );
  IV U68233 ( .A(n55841), .Z(n55844) );
  IV U68234 ( .A(n55842), .Z(n55843) );
  NOR U68235 ( .A(n55844), .B(n55843), .Z(n55845) );
  NOR U68236 ( .A(n55846), .B(n55845), .Z(n55847) );
  XOR U68237 ( .A(n55848), .B(n55847), .Z(n55849) );
  XOR U68238 ( .A(n55850), .B(n55849), .Z(n58083) );
  IV U68239 ( .A(n55851), .Z(n55853) );
  NOR U68240 ( .A(n55853), .B(n55852), .Z(n58081) );
  IV U68241 ( .A(n55854), .Z(n55855) );
  NOR U68242 ( .A(n55856), .B(n55855), .Z(n55862) );
  IV U68243 ( .A(n55857), .Z(n55860) );
  IV U68244 ( .A(n55858), .Z(n55859) );
  NOR U68245 ( .A(n55860), .B(n55859), .Z(n55861) );
  NOR U68246 ( .A(n55862), .B(n55861), .Z(n58079) );
  IV U68247 ( .A(n55863), .Z(n55864) );
  NOR U68248 ( .A(n55864), .B(n58018), .Z(n55869) );
  IV U68249 ( .A(n55865), .Z(n55867) );
  NOR U68250 ( .A(n55867), .B(n55866), .Z(n55868) );
  NOR U68251 ( .A(n55869), .B(n55868), .Z(n58077) );
  NOR U68252 ( .A(n55871), .B(n55870), .Z(n55872) );
  IV U68253 ( .A(n55872), .Z(n55873) );
  NOR U68254 ( .A(n57993), .B(n55873), .Z(n58061) );
  IV U68255 ( .A(n55874), .Z(n55875) );
  NOR U68256 ( .A(n55876), .B(n55875), .Z(n55881) );
  IV U68257 ( .A(n55877), .Z(n55878) );
  NOR U68258 ( .A(n55879), .B(n55878), .Z(n55880) );
  NOR U68259 ( .A(n55881), .B(n55880), .Z(n57991) );
  IV U68260 ( .A(n55882), .Z(n55884) );
  NOR U68261 ( .A(n55884), .B(n55883), .Z(n55889) );
  IV U68262 ( .A(n55885), .Z(n55887) );
  NOR U68263 ( .A(n55887), .B(n55886), .Z(n55888) );
  NOR U68264 ( .A(n55889), .B(n55888), .Z(n57975) );
  NOR U68265 ( .A(n55891), .B(n55890), .Z(n55896) );
  IV U68266 ( .A(n55892), .Z(n55894) );
  NOR U68267 ( .A(n55894), .B(n55893), .Z(n55895) );
  NOR U68268 ( .A(n55896), .B(n55895), .Z(n57959) );
  IV U68269 ( .A(n55897), .Z(n55898) );
  NOR U68270 ( .A(n55899), .B(n55898), .Z(n55904) );
  IV U68271 ( .A(n55900), .Z(n55902) );
  NOR U68272 ( .A(n55902), .B(n55901), .Z(n55903) );
  NOR U68273 ( .A(n55904), .B(n55903), .Z(n55913) );
  IV U68274 ( .A(n55905), .Z(n55907) );
  NOR U68275 ( .A(n55907), .B(n55906), .Z(n55911) );
  NOR U68276 ( .A(n55909), .B(n55908), .Z(n55910) );
  NOR U68277 ( .A(n55911), .B(n55910), .Z(n55912) );
  XOR U68278 ( .A(n55913), .B(n55912), .Z(n57924) );
  NOR U68279 ( .A(n55915), .B(n55914), .Z(n57922) );
  NOR U68280 ( .A(n55917), .B(n55916), .Z(n57920) );
  IV U68281 ( .A(n55918), .Z(n55920) );
  NOR U68282 ( .A(n55920), .B(n55919), .Z(n55940) );
  IV U68283 ( .A(n55921), .Z(n55922) );
  NOR U68284 ( .A(n55923), .B(n55922), .Z(n55928) );
  IV U68285 ( .A(n55924), .Z(n55925) );
  NOR U68286 ( .A(n55926), .B(n55925), .Z(n55927) );
  NOR U68287 ( .A(n55928), .B(n55927), .Z(n55938) );
  IV U68288 ( .A(n55929), .Z(n55931) );
  NOR U68289 ( .A(n55931), .B(n55930), .Z(n55936) );
  IV U68290 ( .A(n55932), .Z(n55933) );
  NOR U68291 ( .A(n55934), .B(n55933), .Z(n55935) );
  NOR U68292 ( .A(n55936), .B(n55935), .Z(n55937) );
  XOR U68293 ( .A(n55938), .B(n55937), .Z(n55939) );
  XOR U68294 ( .A(n55940), .B(n55939), .Z(n55957) );
  IV U68295 ( .A(n55941), .Z(n55943) );
  NOR U68296 ( .A(n55943), .B(n55942), .Z(n55944) );
  NOR U68297 ( .A(n55945), .B(n55944), .Z(n55955) );
  IV U68298 ( .A(n55946), .Z(n55948) );
  NOR U68299 ( .A(n55948), .B(n55947), .Z(n55953) );
  IV U68300 ( .A(n55949), .Z(n55950) );
  NOR U68301 ( .A(n55951), .B(n55950), .Z(n55952) );
  NOR U68302 ( .A(n55953), .B(n55952), .Z(n55954) );
  XOR U68303 ( .A(n55955), .B(n55954), .Z(n55956) );
  XOR U68304 ( .A(n55957), .B(n55956), .Z(n57918) );
  IV U68305 ( .A(n55958), .Z(n55960) );
  NOR U68306 ( .A(n55960), .B(n55959), .Z(n57916) );
  IV U68307 ( .A(n55961), .Z(n55964) );
  IV U68308 ( .A(n55962), .Z(n55963) );
  NOR U68309 ( .A(n55964), .B(n55963), .Z(n57914) );
  IV U68310 ( .A(n55965), .Z(n55966) );
  NOR U68311 ( .A(n55966), .B(n55995), .Z(n55971) );
  IV U68312 ( .A(n55967), .Z(n55969) );
  NOR U68313 ( .A(n55969), .B(n55968), .Z(n55970) );
  NOR U68314 ( .A(n55971), .B(n55970), .Z(n57893) );
  NOR U68315 ( .A(n55972), .B(n55973), .Z(n55982) );
  IV U68316 ( .A(n55973), .Z(n55974) );
  NOR U68317 ( .A(n55975), .B(n55974), .Z(n55980) );
  XOR U68318 ( .A(n55977), .B(n55976), .Z(n55978) );
  IV U68319 ( .A(n55978), .Z(n55979) );
  NOR U68320 ( .A(n55980), .B(n55979), .Z(n55981) );
  NOR U68321 ( .A(n55982), .B(n55981), .Z(n55992) );
  IV U68322 ( .A(n55983), .Z(n55984) );
  NOR U68323 ( .A(n55985), .B(n55984), .Z(n55990) );
  IV U68324 ( .A(n55986), .Z(n55987) );
  NOR U68325 ( .A(n55988), .B(n55987), .Z(n55989) );
  NOR U68326 ( .A(n55990), .B(n55989), .Z(n55991) );
  XOR U68327 ( .A(n55992), .B(n55991), .Z(n56006) );
  IV U68328 ( .A(n55993), .Z(n55994) );
  NOR U68329 ( .A(n55995), .B(n55994), .Z(n56004) );
  NOR U68330 ( .A(n55997), .B(n55996), .Z(n56002) );
  IV U68331 ( .A(n55998), .Z(n55999) );
  NOR U68332 ( .A(n56000), .B(n55999), .Z(n56001) );
  NOR U68333 ( .A(n56002), .B(n56001), .Z(n56003) );
  XOR U68334 ( .A(n56004), .B(n56003), .Z(n56005) );
  XOR U68335 ( .A(n56006), .B(n56005), .Z(n57878) );
  IV U68336 ( .A(n56007), .Z(n56009) );
  NOR U68337 ( .A(n56009), .B(n56008), .Z(n57845) );
  IV U68338 ( .A(n56010), .Z(n56012) );
  NOR U68339 ( .A(n56012), .B(n56011), .Z(n56017) );
  IV U68340 ( .A(n56013), .Z(n56014) );
  NOR U68341 ( .A(n56015), .B(n56014), .Z(n56016) );
  NOR U68342 ( .A(n56017), .B(n56016), .Z(n57843) );
  NOR U68343 ( .A(n56019), .B(n56018), .Z(n57841) );
  IV U68344 ( .A(n56020), .Z(n56022) );
  NOR U68345 ( .A(n56022), .B(n56021), .Z(n56027) );
  IV U68346 ( .A(n56023), .Z(n56025) );
  NOR U68347 ( .A(n56025), .B(n56024), .Z(n56026) );
  NOR U68348 ( .A(n56027), .B(n56026), .Z(n56036) );
  IV U68349 ( .A(n56028), .Z(n56030) );
  NOR U68350 ( .A(n56030), .B(n56029), .Z(n56034) );
  NOR U68351 ( .A(n56032), .B(n56031), .Z(n56033) );
  NOR U68352 ( .A(n56034), .B(n56033), .Z(n56035) );
  XOR U68353 ( .A(n56036), .B(n56035), .Z(n57839) );
  IV U68354 ( .A(n56037), .Z(n56039) );
  NOR U68355 ( .A(n56039), .B(n56038), .Z(n57837) );
  IV U68356 ( .A(n56040), .Z(n56042) );
  NOR U68357 ( .A(n56042), .B(n56041), .Z(n56046) );
  NOR U68358 ( .A(n56044), .B(n56043), .Z(n56045) );
  NOR U68359 ( .A(n56046), .B(n56045), .Z(n56055) );
  IV U68360 ( .A(n56047), .Z(n56048) );
  NOR U68361 ( .A(n56049), .B(n56048), .Z(n56053) );
  NOR U68362 ( .A(n56051), .B(n56050), .Z(n56052) );
  NOR U68363 ( .A(n56053), .B(n56052), .Z(n56054) );
  XOR U68364 ( .A(n56055), .B(n56054), .Z(n56074) );
  NOR U68365 ( .A(n56057), .B(n56056), .Z(n56062) );
  IV U68366 ( .A(n56058), .Z(n56060) );
  NOR U68367 ( .A(n56060), .B(n56059), .Z(n56061) );
  NOR U68368 ( .A(n56062), .B(n56061), .Z(n56072) );
  IV U68369 ( .A(n56063), .Z(n56065) );
  NOR U68370 ( .A(n56065), .B(n56064), .Z(n56070) );
  IV U68371 ( .A(n56066), .Z(n56068) );
  NOR U68372 ( .A(n56068), .B(n56067), .Z(n56069) );
  NOR U68373 ( .A(n56070), .B(n56069), .Z(n56071) );
  XOR U68374 ( .A(n56072), .B(n56071), .Z(n56073) );
  XOR U68375 ( .A(n56074), .B(n56073), .Z(n57835) );
  IV U68376 ( .A(n56075), .Z(n56077) );
  NOR U68377 ( .A(n56077), .B(n56076), .Z(n57833) );
  IV U68378 ( .A(n56078), .Z(n56080) );
  NOR U68379 ( .A(n56080), .B(n56079), .Z(n56085) );
  IV U68380 ( .A(n56081), .Z(n56083) );
  NOR U68381 ( .A(n56083), .B(n56082), .Z(n56084) );
  NOR U68382 ( .A(n56085), .B(n56084), .Z(n57831) );
  IV U68383 ( .A(n56086), .Z(n56088) );
  NOR U68384 ( .A(n56088), .B(n56087), .Z(n56093) );
  IV U68385 ( .A(n56089), .Z(n56091) );
  NOR U68386 ( .A(n56091), .B(n56090), .Z(n56092) );
  NOR U68387 ( .A(n56093), .B(n56092), .Z(n57817) );
  IV U68388 ( .A(n56094), .Z(n57777) );
  XOR U68389 ( .A(n57777), .B(n57778), .Z(n56095) );
  NOR U68390 ( .A(n56096), .B(n56095), .Z(n56101) );
  NOR U68391 ( .A(n57777), .B(n56097), .Z(n56098) );
  NOR U68392 ( .A(n56099), .B(n56098), .Z(n56100) );
  NOR U68393 ( .A(n56101), .B(n56100), .Z(n57815) );
  IV U68394 ( .A(n56102), .Z(n56104) );
  NOR U68395 ( .A(n56104), .B(n56103), .Z(n56106) );
  NOR U68396 ( .A(n56106), .B(n56105), .Z(n57740) );
  IV U68397 ( .A(n56107), .Z(n56109) );
  NOR U68398 ( .A(n56109), .B(n56108), .Z(n57738) );
  IV U68399 ( .A(n56110), .Z(n56111) );
  NOR U68400 ( .A(n56112), .B(n56111), .Z(n56117) );
  IV U68401 ( .A(n56113), .Z(n56115) );
  NOR U68402 ( .A(n56115), .B(n56114), .Z(n56116) );
  NOR U68403 ( .A(n56117), .B(n56116), .Z(n57736) );
  IV U68404 ( .A(n56118), .Z(n56120) );
  NOR U68405 ( .A(n56120), .B(n56119), .Z(n56123) );
  NOR U68406 ( .A(n56122), .B(n56121), .Z(n56129) );
  XOR U68407 ( .A(n56123), .B(n56129), .Z(n56131) );
  IV U68408 ( .A(n56124), .Z(n56126) );
  NOR U68409 ( .A(n56126), .B(n56125), .Z(n56127) );
  IV U68410 ( .A(n56127), .Z(n56128) );
  NOR U68411 ( .A(n56129), .B(n56128), .Z(n56130) );
  NOR U68412 ( .A(n56131), .B(n56130), .Z(n57734) );
  IV U68413 ( .A(n56135), .Z(n56132) );
  NOR U68414 ( .A(n56133), .B(n56132), .Z(n56139) );
  IV U68415 ( .A(n56133), .Z(n56134) );
  NOR U68416 ( .A(n56135), .B(n56134), .Z(n56136) );
  NOR U68417 ( .A(n56137), .B(n56136), .Z(n56138) );
  NOR U68418 ( .A(n56139), .B(n56138), .Z(n57732) );
  IV U68419 ( .A(n56140), .Z(n56142) );
  NOR U68420 ( .A(n56142), .B(n56141), .Z(n56146) );
  NOR U68421 ( .A(n56144), .B(n56143), .Z(n56145) );
  NOR U68422 ( .A(n56146), .B(n56145), .Z(n57717) );
  IV U68423 ( .A(n56147), .Z(n56149) );
  NOR U68424 ( .A(n56149), .B(n56148), .Z(n56153) );
  NOR U68425 ( .A(n56151), .B(n56150), .Z(n56152) );
  NOR U68426 ( .A(n56153), .B(n56152), .Z(n57688) );
  IV U68427 ( .A(n56154), .Z(n56155) );
  NOR U68428 ( .A(n56156), .B(n56155), .Z(n56162) );
  IV U68429 ( .A(n56157), .Z(n56160) );
  IV U68430 ( .A(n56158), .Z(n56159) );
  NOR U68431 ( .A(n56160), .B(n56159), .Z(n56161) );
  NOR U68432 ( .A(n56162), .B(n56161), .Z(n57660) );
  NOR U68433 ( .A(n56164), .B(n56163), .Z(n56165) );
  NOR U68434 ( .A(n56166), .B(n56165), .Z(n56170) );
  NOR U68435 ( .A(n56168), .B(n56167), .Z(n56169) );
  NOR U68436 ( .A(n56170), .B(n56169), .Z(n57631) );
  IV U68437 ( .A(n56171), .Z(n56172) );
  NOR U68438 ( .A(n56173), .B(n56172), .Z(n56178) );
  IV U68439 ( .A(n56174), .Z(n56176) );
  NOR U68440 ( .A(n56176), .B(n56175), .Z(n56177) );
  NOR U68441 ( .A(n56178), .B(n56177), .Z(n57629) );
  IV U68442 ( .A(n56179), .Z(n56181) );
  NOR U68443 ( .A(n56181), .B(n56180), .Z(n56186) );
  IV U68444 ( .A(n56182), .Z(n56184) );
  NOR U68445 ( .A(n56184), .B(n56183), .Z(n56185) );
  NOR U68446 ( .A(n56186), .B(n56185), .Z(n57627) );
  IV U68447 ( .A(n56187), .Z(n56188) );
  NOR U68448 ( .A(n56189), .B(n56188), .Z(n57625) );
  IV U68449 ( .A(n56190), .Z(n56192) );
  NOR U68450 ( .A(n56192), .B(n56191), .Z(n56196) );
  NOR U68451 ( .A(n56194), .B(n56193), .Z(n56195) );
  NOR U68452 ( .A(n56196), .B(n56195), .Z(n57623) );
  NOR U68453 ( .A(n56198), .B(n56197), .Z(n57621) );
  IV U68454 ( .A(n56199), .Z(n56201) );
  NOR U68455 ( .A(n56201), .B(n56200), .Z(n56206) );
  IV U68456 ( .A(n56202), .Z(n56203) );
  NOR U68457 ( .A(n56204), .B(n56203), .Z(n56205) );
  NOR U68458 ( .A(n56206), .B(n56205), .Z(n57599) );
  IV U68459 ( .A(n56207), .Z(n56209) );
  NOR U68460 ( .A(n56209), .B(n56208), .Z(n56214) );
  IV U68461 ( .A(n56210), .Z(n56212) );
  NOR U68462 ( .A(n56212), .B(n56211), .Z(n56213) );
  NOR U68463 ( .A(n56214), .B(n56213), .Z(n57578) );
  NOR U68464 ( .A(n56216), .B(n56215), .Z(n56225) );
  IV U68465 ( .A(n56217), .Z(n56218) );
  NOR U68466 ( .A(n56218), .B(n56220), .Z(n56223) );
  IV U68467 ( .A(n56219), .Z(n56221) );
  NOR U68468 ( .A(n56221), .B(n56220), .Z(n56222) );
  NOR U68469 ( .A(n56223), .B(n56222), .Z(n56224) );
  XOR U68470 ( .A(n56225), .B(n56224), .Z(n57576) );
  IV U68471 ( .A(n56226), .Z(n56227) );
  NOR U68472 ( .A(n56228), .B(n56227), .Z(n56232) );
  IV U68473 ( .A(n56229), .Z(n56230) );
  NOR U68474 ( .A(n56230), .B(n57561), .Z(n56231) );
  NOR U68475 ( .A(n56232), .B(n56231), .Z(n57574) );
  IV U68476 ( .A(n56233), .Z(n56235) );
  IV U68477 ( .A(n56234), .Z(n57587) );
  NOR U68478 ( .A(n56235), .B(n57587), .Z(n57572) );
  IV U68479 ( .A(n56236), .Z(n56237) );
  NOR U68480 ( .A(n56238), .B(n56237), .Z(n56242) );
  NOR U68481 ( .A(n56240), .B(n56239), .Z(n56241) );
  NOR U68482 ( .A(n56242), .B(n56241), .Z(n57570) );
  NOR U68483 ( .A(n56244), .B(n56243), .Z(n56250) );
  IV U68484 ( .A(n56244), .Z(n56246) );
  NOR U68485 ( .A(n56246), .B(n56245), .Z(n56247) );
  NOR U68486 ( .A(n56248), .B(n56247), .Z(n56249) );
  NOR U68487 ( .A(n56250), .B(n56249), .Z(n56260) );
  IV U68488 ( .A(n56251), .Z(n56252) );
  NOR U68489 ( .A(n56253), .B(n56252), .Z(n56258) );
  IV U68490 ( .A(n56254), .Z(n56255) );
  NOR U68491 ( .A(n56256), .B(n56255), .Z(n56257) );
  NOR U68492 ( .A(n56258), .B(n56257), .Z(n56259) );
  XOR U68493 ( .A(n56260), .B(n56259), .Z(n57548) );
  IV U68494 ( .A(n56261), .Z(n56263) );
  NOR U68495 ( .A(n56263), .B(n56262), .Z(n56267) );
  NOR U68496 ( .A(n56265), .B(n56264), .Z(n56266) );
  NOR U68497 ( .A(n56267), .B(n56266), .Z(n57546) );
  IV U68498 ( .A(n56268), .Z(n56270) );
  NOR U68499 ( .A(n56270), .B(n56269), .Z(n56275) );
  IV U68500 ( .A(n56271), .Z(n56273) );
  NOR U68501 ( .A(n56273), .B(n56272), .Z(n56274) );
  NOR U68502 ( .A(n56275), .B(n56274), .Z(n57544) );
  NOR U68503 ( .A(n56277), .B(n56276), .Z(n57542) );
  NOR U68504 ( .A(n56279), .B(n56278), .Z(n56284) );
  IV U68505 ( .A(n56280), .Z(n56281) );
  NOR U68506 ( .A(n56282), .B(n56281), .Z(n56283) );
  NOR U68507 ( .A(n56284), .B(n56283), .Z(n56300) );
  IV U68508 ( .A(n56285), .Z(n56286) );
  NOR U68509 ( .A(n56287), .B(n56286), .Z(n56298) );
  IV U68510 ( .A(n56288), .Z(n56289) );
  NOR U68511 ( .A(n56290), .B(n56289), .Z(n56295) );
  IV U68512 ( .A(n56291), .Z(n56293) );
  NOR U68513 ( .A(n56293), .B(n56292), .Z(n56294) );
  NOR U68514 ( .A(n56295), .B(n56294), .Z(n56296) );
  IV U68515 ( .A(n56296), .Z(n56297) );
  NOR U68516 ( .A(n56298), .B(n56297), .Z(n56299) );
  XOR U68517 ( .A(n56300), .B(n56299), .Z(n56313) );
  IV U68518 ( .A(n56301), .Z(n56303) );
  NOR U68519 ( .A(n56303), .B(n56302), .Z(n56311) );
  IV U68520 ( .A(n56304), .Z(n56305) );
  NOR U68521 ( .A(n56306), .B(n56305), .Z(n56308) );
  NOR U68522 ( .A(n56308), .B(n56307), .Z(n56309) );
  IV U68523 ( .A(n56309), .Z(n56310) );
  NOR U68524 ( .A(n56311), .B(n56310), .Z(n56312) );
  XOR U68525 ( .A(n56313), .B(n56312), .Z(n57540) );
  IV U68526 ( .A(n56314), .Z(n56315) );
  NOR U68527 ( .A(n56316), .B(n56315), .Z(n56320) );
  NOR U68528 ( .A(n56318), .B(n56317), .Z(n56319) );
  NOR U68529 ( .A(n56320), .B(n56319), .Z(n57538) );
  IV U68530 ( .A(n56321), .Z(n56323) );
  NOR U68531 ( .A(n56323), .B(n56322), .Z(n56327) );
  IV U68532 ( .A(n56324), .Z(n56325) );
  NOR U68533 ( .A(n56325), .B(n56340), .Z(n56326) );
  NOR U68534 ( .A(n56327), .B(n56326), .Z(n57524) );
  IV U68535 ( .A(n56328), .Z(n56330) );
  NOR U68536 ( .A(n56330), .B(n56329), .Z(n56338) );
  IV U68537 ( .A(n56331), .Z(n56333) );
  NOR U68538 ( .A(n56333), .B(n56332), .Z(n56335) );
  NOR U68539 ( .A(n56335), .B(n56334), .Z(n56336) );
  IV U68540 ( .A(n56336), .Z(n56337) );
  NOR U68541 ( .A(n56338), .B(n56337), .Z(n57522) );
  NOR U68542 ( .A(n56339), .B(n56340), .Z(n56345) );
  XOR U68543 ( .A(n56341), .B(n56340), .Z(n56342) );
  NOR U68544 ( .A(n56343), .B(n56342), .Z(n56344) );
  NOR U68545 ( .A(n56345), .B(n56344), .Z(n57520) );
  NOR U68546 ( .A(n56347), .B(n56346), .Z(n56351) );
  IV U68547 ( .A(n56348), .Z(n56350) );
  NOR U68548 ( .A(n56350), .B(n56349), .Z(n56357) );
  XOR U68549 ( .A(n56351), .B(n56357), .Z(n56359) );
  IV U68550 ( .A(n56352), .Z(n56353) );
  NOR U68551 ( .A(n56354), .B(n56353), .Z(n56355) );
  IV U68552 ( .A(n56355), .Z(n56356) );
  NOR U68553 ( .A(n56357), .B(n56356), .Z(n56358) );
  NOR U68554 ( .A(n56359), .B(n56358), .Z(n57497) );
  NOR U68555 ( .A(n56361), .B(n56360), .Z(n56363) );
  NOR U68556 ( .A(n56363), .B(n56362), .Z(n57495) );
  NOR U68557 ( .A(n56365), .B(n56364), .Z(n56370) );
  IV U68558 ( .A(n56366), .Z(n56367) );
  NOR U68559 ( .A(n56368), .B(n56367), .Z(n56369) );
  NOR U68560 ( .A(n56370), .B(n56369), .Z(n57493) );
  IV U68561 ( .A(n56373), .Z(n56371) );
  NOR U68562 ( .A(n56372), .B(n56371), .Z(n56380) );
  NOR U68563 ( .A(n56374), .B(n56373), .Z(n56378) );
  XOR U68564 ( .A(n56376), .B(n56375), .Z(n56377) );
  NOR U68565 ( .A(n56378), .B(n56377), .Z(n56379) );
  NOR U68566 ( .A(n56380), .B(n56379), .Z(n57491) );
  IV U68567 ( .A(n56381), .Z(n56382) );
  NOR U68568 ( .A(n56383), .B(n56382), .Z(n56388) );
  IV U68569 ( .A(n56384), .Z(n56386) );
  NOR U68570 ( .A(n56386), .B(n56385), .Z(n56387) );
  NOR U68571 ( .A(n56388), .B(n56387), .Z(n57489) );
  IV U68572 ( .A(n56389), .Z(n56390) );
  NOR U68573 ( .A(n56391), .B(n56390), .Z(n56396) );
  IV U68574 ( .A(n56392), .Z(n56394) );
  NOR U68575 ( .A(n56394), .B(n56393), .Z(n56395) );
  NOR U68576 ( .A(n56396), .B(n56395), .Z(n56401) );
  IV U68577 ( .A(n56397), .Z(n56399) );
  NOR U68578 ( .A(n56399), .B(n56398), .Z(n56400) );
  XOR U68579 ( .A(n56401), .B(n56400), .Z(n57487) );
  IV U68580 ( .A(n56402), .Z(n56403) );
  NOR U68581 ( .A(n56404), .B(n56403), .Z(n56408) );
  NOR U68582 ( .A(n56406), .B(n56405), .Z(n56407) );
  NOR U68583 ( .A(n56408), .B(n56407), .Z(n56415) );
  IV U68584 ( .A(n56409), .Z(n56411) );
  NOR U68585 ( .A(n56411), .B(n56410), .Z(n56412) );
  NOR U68586 ( .A(n56413), .B(n56412), .Z(n56414) );
  XOR U68587 ( .A(n56415), .B(n56414), .Z(n56425) );
  IV U68588 ( .A(n56416), .Z(n56418) );
  NOR U68589 ( .A(n56418), .B(n56417), .Z(n56423) );
  IV U68590 ( .A(n56419), .Z(n56420) );
  NOR U68591 ( .A(n56421), .B(n56420), .Z(n56422) );
  NOR U68592 ( .A(n56423), .B(n56422), .Z(n56424) );
  XOR U68593 ( .A(n56425), .B(n56424), .Z(n56443) );
  NOR U68594 ( .A(n56427), .B(n56426), .Z(n56435) );
  IV U68595 ( .A(n56427), .Z(n56428) );
  NOR U68596 ( .A(n56429), .B(n56428), .Z(n56433) );
  XOR U68597 ( .A(n56431), .B(n56430), .Z(n56432) );
  NOR U68598 ( .A(n56433), .B(n56432), .Z(n56434) );
  NOR U68599 ( .A(n56435), .B(n56434), .Z(n56441) );
  NOR U68600 ( .A(n56437), .B(n56436), .Z(n56438) );
  NOR U68601 ( .A(n56439), .B(n56438), .Z(n56440) );
  XOR U68602 ( .A(n56441), .B(n56440), .Z(n56442) );
  XOR U68603 ( .A(n56443), .B(n56442), .Z(n57485) );
  IV U68604 ( .A(n56444), .Z(n56446) );
  NOR U68605 ( .A(n56446), .B(n56445), .Z(n57483) );
  IV U68606 ( .A(n56447), .Z(n56449) );
  NOR U68607 ( .A(n56449), .B(n56448), .Z(n56453) );
  NOR U68608 ( .A(n56451), .B(n56450), .Z(n56452) );
  NOR U68609 ( .A(n56453), .B(n56452), .Z(n57468) );
  IV U68610 ( .A(n56454), .Z(n56455) );
  NOR U68611 ( .A(n56456), .B(n56455), .Z(n56460) );
  IV U68612 ( .A(n56457), .Z(n56458) );
  NOR U68613 ( .A(n56459), .B(n56458), .Z(n56466) );
  XOR U68614 ( .A(n56460), .B(n56466), .Z(n56468) );
  IV U68615 ( .A(n56461), .Z(n56462) );
  NOR U68616 ( .A(n56463), .B(n56462), .Z(n56464) );
  IV U68617 ( .A(n56464), .Z(n56465) );
  NOR U68618 ( .A(n56466), .B(n56465), .Z(n56467) );
  NOR U68619 ( .A(n56468), .B(n56467), .Z(n57403) );
  IV U68620 ( .A(n56469), .Z(n56470) );
  NOR U68621 ( .A(n56471), .B(n56470), .Z(n56476) );
  IV U68622 ( .A(n56472), .Z(n56474) );
  NOR U68623 ( .A(n56474), .B(n56473), .Z(n56475) );
  NOR U68624 ( .A(n56476), .B(n56475), .Z(n57401) );
  IV U68625 ( .A(n56477), .Z(n56479) );
  NOR U68626 ( .A(n56479), .B(n56478), .Z(n56482) );
  NOR U68627 ( .A(n56480), .B(n57389), .Z(n56481) );
  NOR U68628 ( .A(n56482), .B(n56481), .Z(n57384) );
  IV U68629 ( .A(n56483), .Z(n56485) );
  NOR U68630 ( .A(n56485), .B(n56484), .Z(n57357) );
  IV U68631 ( .A(n56486), .Z(n56488) );
  NOR U68632 ( .A(n56488), .B(n56487), .Z(n56499) );
  IV U68633 ( .A(n56489), .Z(n56490) );
  NOR U68634 ( .A(n56491), .B(n56490), .Z(n56496) );
  IV U68635 ( .A(n56492), .Z(n56493) );
  NOR U68636 ( .A(n56494), .B(n56493), .Z(n56495) );
  NOR U68637 ( .A(n56496), .B(n56495), .Z(n56497) );
  IV U68638 ( .A(n56497), .Z(n56498) );
  NOR U68639 ( .A(n56499), .B(n56498), .Z(n57315) );
  IV U68640 ( .A(n56500), .Z(n56502) );
  NOR U68641 ( .A(n56502), .B(n56501), .Z(n56507) );
  IV U68642 ( .A(n56503), .Z(n56505) );
  NOR U68643 ( .A(n56505), .B(n56504), .Z(n56506) );
  NOR U68644 ( .A(n56507), .B(n56506), .Z(n57267) );
  IV U68645 ( .A(n56508), .Z(n56509) );
  NOR U68646 ( .A(n56509), .B(n57254), .Z(n56512) );
  NOR U68647 ( .A(n56511), .B(n56510), .Z(n56518) );
  XOR U68648 ( .A(n56512), .B(n56518), .Z(n56520) );
  IV U68649 ( .A(n56513), .Z(n56515) );
  NOR U68650 ( .A(n56515), .B(n56514), .Z(n56516) );
  IV U68651 ( .A(n56516), .Z(n56517) );
  NOR U68652 ( .A(n56518), .B(n56517), .Z(n56519) );
  NOR U68653 ( .A(n56520), .B(n56519), .Z(n57265) );
  IV U68654 ( .A(n56521), .Z(n56522) );
  NOR U68655 ( .A(n56523), .B(n56522), .Z(n56528) );
  IV U68656 ( .A(n56524), .Z(n56526) );
  NOR U68657 ( .A(n56526), .B(n56525), .Z(n56527) );
  NOR U68658 ( .A(n56528), .B(n56527), .Z(n57244) );
  IV U68659 ( .A(n56529), .Z(n56530) );
  NOR U68660 ( .A(n56531), .B(n56530), .Z(n56536) );
  IV U68661 ( .A(n56532), .Z(n56533) );
  NOR U68662 ( .A(n56534), .B(n56533), .Z(n56535) );
  NOR U68663 ( .A(n56536), .B(n56535), .Z(n57240) );
  NOR U68664 ( .A(n56538), .B(n56537), .Z(n57238) );
  IV U68665 ( .A(n56539), .Z(n56540) );
  NOR U68666 ( .A(n56541), .B(n56540), .Z(n57187) );
  IV U68667 ( .A(n56542), .Z(n56544) );
  NOR U68668 ( .A(n56544), .B(n56543), .Z(n56548) );
  NOR U68669 ( .A(n56546), .B(n56545), .Z(n56547) );
  NOR U68670 ( .A(n56548), .B(n56547), .Z(n57160) );
  NOR U68671 ( .A(n56550), .B(n56549), .Z(n56556) );
  NOR U68672 ( .A(n56552), .B(n56551), .Z(n56554) );
  NOR U68673 ( .A(n56554), .B(n56553), .Z(n56555) );
  NOR U68674 ( .A(n56556), .B(n56555), .Z(n57158) );
  IV U68675 ( .A(n56557), .Z(n56559) );
  NOR U68676 ( .A(n56559), .B(n56558), .Z(n56564) );
  IV U68677 ( .A(n56560), .Z(n56562) );
  NOR U68678 ( .A(n56562), .B(n56561), .Z(n56563) );
  NOR U68679 ( .A(n56564), .B(n56563), .Z(n57149) );
  NOR U68680 ( .A(n56566), .B(n56565), .Z(n56567) );
  IV U68681 ( .A(n56567), .Z(n56569) );
  NOR U68682 ( .A(n56569), .B(n56568), .Z(n56577) );
  NOR U68683 ( .A(n56571), .B(n56570), .Z(n56572) );
  IV U68684 ( .A(n56572), .Z(n56575) );
  IV U68685 ( .A(n56573), .Z(n56574) );
  NOR U68686 ( .A(n56575), .B(n56574), .Z(n56576) );
  NOR U68687 ( .A(n56577), .B(n56576), .Z(n57147) );
  IV U68688 ( .A(n56578), .Z(n56579) );
  NOR U68689 ( .A(n56580), .B(n56579), .Z(n57083) );
  NOR U68690 ( .A(n56583), .B(n56587), .Z(n56585) );
  IV U68691 ( .A(n56581), .Z(n56582) );
  NOR U68692 ( .A(n56583), .B(n56582), .Z(n56584) );
  NOR U68693 ( .A(n56585), .B(n56584), .Z(n57050) );
  XOR U68694 ( .A(n56587), .B(n56586), .Z(n56588) );
  NOR U68695 ( .A(n56589), .B(n56588), .Z(n56594) );
  IV U68696 ( .A(n56590), .Z(n56592) );
  NOR U68697 ( .A(n56592), .B(n56591), .Z(n56593) );
  NOR U68698 ( .A(n56594), .B(n56593), .Z(n57018) );
  NOR U68699 ( .A(n56600), .B(n56595), .Z(n56597) );
  NOR U68700 ( .A(n56597), .B(n56596), .Z(n56606) );
  NOR U68701 ( .A(n56599), .B(n56598), .Z(n56604) );
  IV U68702 ( .A(n56600), .Z(n56602) );
  NOR U68703 ( .A(n56602), .B(n56601), .Z(n56603) );
  NOR U68704 ( .A(n56604), .B(n56603), .Z(n56605) );
  IV U68705 ( .A(n56605), .Z(n56610) );
  NOR U68706 ( .A(n56606), .B(n56610), .Z(n56613) );
  IV U68707 ( .A(n56607), .Z(n56609) );
  NOR U68708 ( .A(n56609), .B(n56608), .Z(n56611) );
  NOR U68709 ( .A(n56611), .B(n56610), .Z(n56612) );
  NOR U68710 ( .A(n56613), .B(n56612), .Z(n57016) );
  IV U68711 ( .A(n56614), .Z(n56615) );
  NOR U68712 ( .A(n56616), .B(n56615), .Z(n56620) );
  NOR U68713 ( .A(n56618), .B(n56617), .Z(n56619) );
  NOR U68714 ( .A(n56620), .B(n56619), .Z(n57014) );
  NOR U68715 ( .A(n56621), .B(n56622), .Z(n56634) );
  IV U68716 ( .A(n56621), .Z(n56624) );
  IV U68717 ( .A(n56622), .Z(n56623) );
  NOR U68718 ( .A(n56624), .B(n56623), .Z(n56632) );
  IV U68719 ( .A(n56625), .Z(n56626) );
  NOR U68720 ( .A(n56627), .B(n56626), .Z(n56628) );
  NOR U68721 ( .A(n56629), .B(n56628), .Z(n56630) );
  IV U68722 ( .A(n56630), .Z(n56631) );
  NOR U68723 ( .A(n56632), .B(n56631), .Z(n56633) );
  NOR U68724 ( .A(n56634), .B(n56633), .Z(n57012) );
  IV U68725 ( .A(n56635), .Z(n56636) );
  NOR U68726 ( .A(n56637), .B(n56636), .Z(n56994) );
  IV U68727 ( .A(n56638), .Z(n56641) );
  IV U68728 ( .A(n56639), .Z(n56640) );
  NOR U68729 ( .A(n56641), .B(n56640), .Z(n56973) );
  IV U68730 ( .A(n56642), .Z(n56643) );
  NOR U68731 ( .A(n56643), .B(n56645), .Z(n56648) );
  IV U68732 ( .A(n56644), .Z(n56646) );
  NOR U68733 ( .A(n56646), .B(n56645), .Z(n56647) );
  NOR U68734 ( .A(n56648), .B(n56647), .Z(n56951) );
  IV U68735 ( .A(n56649), .Z(n56650) );
  NOR U68736 ( .A(n56651), .B(n56650), .Z(n56947) );
  IV U68737 ( .A(n56652), .Z(n56654) );
  NOR U68738 ( .A(n56654), .B(n56653), .Z(n56945) );
  IV U68739 ( .A(n56655), .Z(n56657) );
  NOR U68740 ( .A(n56657), .B(n56656), .Z(n56662) );
  IV U68741 ( .A(n56658), .Z(n56660) );
  NOR U68742 ( .A(n56660), .B(n56659), .Z(n56661) );
  NOR U68743 ( .A(n56662), .B(n56661), .Z(n56943) );
  IV U68744 ( .A(n56663), .Z(n56664) );
  NOR U68745 ( .A(n56665), .B(n56664), .Z(n56915) );
  IV U68746 ( .A(n56666), .Z(n56668) );
  NOR U68747 ( .A(n56668), .B(n56667), .Z(n56913) );
  IV U68748 ( .A(n56669), .Z(n56671) );
  NOR U68749 ( .A(n56671), .B(n56670), .Z(n56676) );
  IV U68750 ( .A(n56672), .Z(n56674) );
  NOR U68751 ( .A(n56674), .B(n56673), .Z(n56675) );
  NOR U68752 ( .A(n56676), .B(n56675), .Z(n56905) );
  IV U68753 ( .A(n56677), .Z(n56678) );
  NOR U68754 ( .A(n56679), .B(n56678), .Z(n56684) );
  IV U68755 ( .A(n56680), .Z(n56681) );
  NOR U68756 ( .A(n56682), .B(n56681), .Z(n56683) );
  NOR U68757 ( .A(n56684), .B(n56683), .Z(n56868) );
  IV U68758 ( .A(n56685), .Z(n56687) );
  NOR U68759 ( .A(n56687), .B(n56686), .Z(n56866) );
  IV U68760 ( .A(n56688), .Z(n56690) );
  NOR U68761 ( .A(n56690), .B(n56689), .Z(n56695) );
  IV U68762 ( .A(n56691), .Z(n56693) );
  NOR U68763 ( .A(n56693), .B(n56692), .Z(n56694) );
  NOR U68764 ( .A(n56695), .B(n56694), .Z(n56827) );
  IV U68765 ( .A(n56696), .Z(n56698) );
  NOR U68766 ( .A(n56698), .B(n56697), .Z(n56825) );
  NOR U68767 ( .A(n56700), .B(n56699), .Z(n56705) );
  IV U68768 ( .A(n56701), .Z(n56703) );
  NOR U68769 ( .A(n56703), .B(n56702), .Z(n56704) );
  NOR U68770 ( .A(n56705), .B(n56704), .Z(n56809) );
  NOR U68771 ( .A(n56707), .B(n56706), .Z(n56807) );
  IV U68772 ( .A(n56708), .Z(n56710) );
  NOR U68773 ( .A(n56710), .B(n56709), .Z(n56714) );
  NOR U68774 ( .A(n56712), .B(n56711), .Z(n56713) );
  NOR U68775 ( .A(n56714), .B(n56713), .Z(n56805) );
  NOR U68776 ( .A(n56716), .B(n56715), .Z(n56784) );
  NOR U68777 ( .A(n56718), .B(n56717), .Z(n56719) );
  NOR U68778 ( .A(n56720), .B(n56719), .Z(n56780) );
  NOR U68779 ( .A(n56722), .B(n56721), .Z(n56778) );
  IV U68780 ( .A(n56723), .Z(n56725) );
  NOR U68781 ( .A(n56725), .B(n56724), .Z(n56765) );
  IV U68782 ( .A(n56726), .Z(n56727) );
  NOR U68783 ( .A(n56728), .B(n56727), .Z(n56733) );
  IV U68784 ( .A(n56729), .Z(n56731) );
  NOR U68785 ( .A(n56731), .B(n56730), .Z(n56732) );
  NOR U68786 ( .A(n56733), .B(n56732), .Z(n56740) );
  IV U68787 ( .A(n56734), .Z(n56735) );
  NOR U68788 ( .A(n56736), .B(n56735), .Z(n56737) );
  NOR U68789 ( .A(n56738), .B(n56737), .Z(n56739) );
  XOR U68790 ( .A(n56740), .B(n56739), .Z(n56751) );
  NOR U68791 ( .A(n56741), .B(n56743), .Z(n56749) );
  IV U68792 ( .A(n56742), .Z(n56747) );
  IV U68793 ( .A(n56743), .Z(n56745) );
  NOR U68794 ( .A(n56745), .B(n56744), .Z(n56746) );
  NOR U68795 ( .A(n56747), .B(n56746), .Z(n56748) );
  NOR U68796 ( .A(n56749), .B(n56748), .Z(n56750) );
  XOR U68797 ( .A(n56751), .B(n56750), .Z(n56763) );
  NOR U68798 ( .A(n56753), .B(n56752), .Z(n56761) );
  NOR U68799 ( .A(n56755), .B(n56754), .Z(n56759) );
  XOR U68800 ( .A(n56757), .B(n56756), .Z(n56758) );
  NOR U68801 ( .A(n56759), .B(n56758), .Z(n56760) );
  NOR U68802 ( .A(n56761), .B(n56760), .Z(n56762) );
  XOR U68803 ( .A(n56763), .B(n56762), .Z(n56764) );
  XOR U68804 ( .A(n56765), .B(n56764), .Z(n56776) );
  NOR U68805 ( .A(n56766), .B(n56768), .Z(n56771) );
  IV U68806 ( .A(n56767), .Z(n56769) );
  NOR U68807 ( .A(n56769), .B(n56768), .Z(n56770) );
  NOR U68808 ( .A(n56771), .B(n56770), .Z(n56772) );
  IV U68809 ( .A(n56772), .Z(n56773) );
  NOR U68810 ( .A(n56774), .B(n56773), .Z(n56775) );
  XOR U68811 ( .A(n56776), .B(n56775), .Z(n56777) );
  XOR U68812 ( .A(n56778), .B(n56777), .Z(n56779) );
  XOR U68813 ( .A(n56780), .B(n56779), .Z(n56781) );
  XOR U68814 ( .A(n56782), .B(n56781), .Z(n56783) );
  XOR U68815 ( .A(n56784), .B(n56783), .Z(n56803) );
  IV U68816 ( .A(n56785), .Z(n56786) );
  NOR U68817 ( .A(n56787), .B(n56786), .Z(n56792) );
  IV U68818 ( .A(n56788), .Z(n56790) );
  NOR U68819 ( .A(n56790), .B(n56789), .Z(n56791) );
  NOR U68820 ( .A(n56792), .B(n56791), .Z(n56801) );
  NOR U68821 ( .A(n56794), .B(n56793), .Z(n56799) );
  IV U68822 ( .A(n56795), .Z(n56796) );
  NOR U68823 ( .A(n56797), .B(n56796), .Z(n56798) );
  NOR U68824 ( .A(n56799), .B(n56798), .Z(n56800) );
  XOR U68825 ( .A(n56801), .B(n56800), .Z(n56802) );
  XOR U68826 ( .A(n56803), .B(n56802), .Z(n56804) );
  XOR U68827 ( .A(n56805), .B(n56804), .Z(n56806) );
  XOR U68828 ( .A(n56807), .B(n56806), .Z(n56808) );
  XOR U68829 ( .A(n56809), .B(n56808), .Z(n56823) );
  NOR U68830 ( .A(n56811), .B(n56810), .Z(n56821) );
  IV U68831 ( .A(n56812), .Z(n56814) );
  NOR U68832 ( .A(n56814), .B(n56813), .Z(n56818) );
  NOR U68833 ( .A(n56816), .B(n56815), .Z(n56817) );
  NOR U68834 ( .A(n56818), .B(n56817), .Z(n56819) );
  IV U68835 ( .A(n56819), .Z(n56820) );
  NOR U68836 ( .A(n56821), .B(n56820), .Z(n56822) );
  XOR U68837 ( .A(n56823), .B(n56822), .Z(n56824) );
  XOR U68838 ( .A(n56825), .B(n56824), .Z(n56826) );
  XOR U68839 ( .A(n56827), .B(n56826), .Z(n56839) );
  IV U68840 ( .A(n56828), .Z(n56829) );
  NOR U68841 ( .A(n56830), .B(n56829), .Z(n56831) );
  NOR U68842 ( .A(n56832), .B(n56831), .Z(n56837) );
  IV U68843 ( .A(n56833), .Z(n56835) );
  NOR U68844 ( .A(n56835), .B(n56834), .Z(n56836) );
  XOR U68845 ( .A(n56837), .B(n56836), .Z(n56838) );
  XOR U68846 ( .A(n56839), .B(n56838), .Z(n56855) );
  IV U68847 ( .A(n56840), .Z(n56842) );
  NOR U68848 ( .A(n56842), .B(n56841), .Z(n56853) );
  IV U68849 ( .A(n56843), .Z(n56845) );
  NOR U68850 ( .A(n56845), .B(n56844), .Z(n56850) );
  IV U68851 ( .A(n56846), .Z(n56848) );
  NOR U68852 ( .A(n56848), .B(n56847), .Z(n56849) );
  NOR U68853 ( .A(n56850), .B(n56849), .Z(n56851) );
  IV U68854 ( .A(n56851), .Z(n56852) );
  NOR U68855 ( .A(n56853), .B(n56852), .Z(n56854) );
  XOR U68856 ( .A(n56855), .B(n56854), .Z(n56864) );
  IV U68857 ( .A(n56856), .Z(n56858) );
  NOR U68858 ( .A(n56858), .B(n56857), .Z(n56862) );
  NOR U68859 ( .A(n56860), .B(n56859), .Z(n56861) );
  NOR U68860 ( .A(n56862), .B(n56861), .Z(n56863) );
  XOR U68861 ( .A(n56864), .B(n56863), .Z(n56865) );
  XOR U68862 ( .A(n56866), .B(n56865), .Z(n56867) );
  XOR U68863 ( .A(n56868), .B(n56867), .Z(n56884) );
  IV U68864 ( .A(n56869), .Z(n56871) );
  NOR U68865 ( .A(n56871), .B(n56870), .Z(n56875) );
  NOR U68866 ( .A(n56873), .B(n56872), .Z(n56874) );
  NOR U68867 ( .A(n56875), .B(n56874), .Z(n56877) );
  NOR U68868 ( .A(n56877), .B(n56876), .Z(n56882) );
  IV U68869 ( .A(n56878), .Z(n56880) );
  NOR U68870 ( .A(n56880), .B(n56879), .Z(n56881) );
  NOR U68871 ( .A(n56882), .B(n56881), .Z(n56883) );
  XOR U68872 ( .A(n56884), .B(n56883), .Z(n56903) );
  IV U68873 ( .A(n56885), .Z(n56887) );
  NOR U68874 ( .A(n56887), .B(n56886), .Z(n56892) );
  IV U68875 ( .A(n56888), .Z(n56890) );
  NOR U68876 ( .A(n56890), .B(n56889), .Z(n56891) );
  NOR U68877 ( .A(n56892), .B(n56891), .Z(n56901) );
  IV U68878 ( .A(n56893), .Z(n56894) );
  NOR U68879 ( .A(n56894), .B(n56896), .Z(n56899) );
  IV U68880 ( .A(n56895), .Z(n56897) );
  NOR U68881 ( .A(n56897), .B(n56896), .Z(n56898) );
  XOR U68882 ( .A(n56899), .B(n56898), .Z(n56900) );
  XOR U68883 ( .A(n56901), .B(n56900), .Z(n56902) );
  XOR U68884 ( .A(n56903), .B(n56902), .Z(n56904) );
  XOR U68885 ( .A(n56905), .B(n56904), .Z(n56911) );
  NOR U68886 ( .A(n56907), .B(n56906), .Z(n56909) );
  NOR U68887 ( .A(n56909), .B(n56908), .Z(n56910) );
  XOR U68888 ( .A(n56911), .B(n56910), .Z(n56912) );
  XOR U68889 ( .A(n56913), .B(n56912), .Z(n56914) );
  XOR U68890 ( .A(n56915), .B(n56914), .Z(n56941) );
  IV U68891 ( .A(n56916), .Z(n56918) );
  NOR U68892 ( .A(n56918), .B(n56917), .Z(n56923) );
  IV U68893 ( .A(n56919), .Z(n56921) );
  NOR U68894 ( .A(n56921), .B(n56920), .Z(n56922) );
  NOR U68895 ( .A(n56923), .B(n56922), .Z(n56933) );
  IV U68896 ( .A(n56924), .Z(n56926) );
  NOR U68897 ( .A(n56926), .B(n56925), .Z(n56931) );
  IV U68898 ( .A(n56927), .Z(n56929) );
  NOR U68899 ( .A(n56929), .B(n56928), .Z(n56930) );
  NOR U68900 ( .A(n56931), .B(n56930), .Z(n56932) );
  XOR U68901 ( .A(n56933), .B(n56932), .Z(n56939) );
  NOR U68902 ( .A(n56935), .B(n56934), .Z(n56937) );
  NOR U68903 ( .A(n56937), .B(n56936), .Z(n56938) );
  XOR U68904 ( .A(n56939), .B(n56938), .Z(n56940) );
  XOR U68905 ( .A(n56941), .B(n56940), .Z(n56942) );
  XOR U68906 ( .A(n56943), .B(n56942), .Z(n56944) );
  XOR U68907 ( .A(n56945), .B(n56944), .Z(n56946) );
  XOR U68908 ( .A(n56947), .B(n56946), .Z(n56948) );
  XOR U68909 ( .A(n56949), .B(n56948), .Z(n56950) );
  XOR U68910 ( .A(n56951), .B(n56950), .Z(n56971) );
  IV U68911 ( .A(n56952), .Z(n56953) );
  NOR U68912 ( .A(n56954), .B(n56953), .Z(n56959) );
  IV U68913 ( .A(n56955), .Z(n56957) );
  NOR U68914 ( .A(n56957), .B(n56956), .Z(n56958) );
  NOR U68915 ( .A(n56959), .B(n56958), .Z(n56969) );
  IV U68916 ( .A(n56960), .Z(n56962) );
  NOR U68917 ( .A(n56962), .B(n56961), .Z(n56967) );
  IV U68918 ( .A(n56963), .Z(n56965) );
  NOR U68919 ( .A(n56965), .B(n56964), .Z(n56966) );
  NOR U68920 ( .A(n56967), .B(n56966), .Z(n56968) );
  XOR U68921 ( .A(n56969), .B(n56968), .Z(n56970) );
  XOR U68922 ( .A(n56971), .B(n56970), .Z(n56972) );
  XOR U68923 ( .A(n56973), .B(n56972), .Z(n56992) );
  IV U68924 ( .A(n56974), .Z(n56975) );
  NOR U68925 ( .A(n56976), .B(n56975), .Z(n56980) );
  NOR U68926 ( .A(n56978), .B(n56977), .Z(n56979) );
  NOR U68927 ( .A(n56980), .B(n56979), .Z(n56990) );
  NOR U68928 ( .A(n56982), .B(n56981), .Z(n56988) );
  IV U68929 ( .A(n56983), .Z(n56986) );
  IV U68930 ( .A(n56984), .Z(n56985) );
  NOR U68931 ( .A(n56986), .B(n56985), .Z(n56987) );
  NOR U68932 ( .A(n56988), .B(n56987), .Z(n56989) );
  XOR U68933 ( .A(n56990), .B(n56989), .Z(n56991) );
  XOR U68934 ( .A(n56992), .B(n56991), .Z(n56993) );
  XOR U68935 ( .A(n56994), .B(n56993), .Z(n57004) );
  NOR U68936 ( .A(n56995), .B(n56996), .Z(n57002) );
  IV U68937 ( .A(n56996), .Z(n56997) );
  NOR U68938 ( .A(n56998), .B(n56997), .Z(n56999) );
  NOR U68939 ( .A(n57000), .B(n56999), .Z(n57001) );
  NOR U68940 ( .A(n57002), .B(n57001), .Z(n57003) );
  XOR U68941 ( .A(n57004), .B(n57003), .Z(n57010) );
  NOR U68942 ( .A(n57006), .B(n57005), .Z(n57008) );
  NOR U68943 ( .A(n57008), .B(n57007), .Z(n57009) );
  XOR U68944 ( .A(n57010), .B(n57009), .Z(n57011) );
  XOR U68945 ( .A(n57012), .B(n57011), .Z(n57013) );
  XOR U68946 ( .A(n57014), .B(n57013), .Z(n57015) );
  XOR U68947 ( .A(n57016), .B(n57015), .Z(n57017) );
  XOR U68948 ( .A(n57018), .B(n57017), .Z(n57048) );
  IV U68949 ( .A(n57019), .Z(n57020) );
  NOR U68950 ( .A(n57021), .B(n57020), .Z(n57026) );
  IV U68951 ( .A(n57022), .Z(n57024) );
  NOR U68952 ( .A(n57024), .B(n57023), .Z(n57025) );
  NOR U68953 ( .A(n57026), .B(n57025), .Z(n57046) );
  IV U68954 ( .A(n57027), .Z(n57028) );
  NOR U68955 ( .A(n57029), .B(n57028), .Z(n57044) );
  NOR U68956 ( .A(n57031), .B(n57030), .Z(n57032) );
  IV U68957 ( .A(n57032), .Z(n57033) );
  NOR U68958 ( .A(n57034), .B(n57033), .Z(n57035) );
  IV U68959 ( .A(n57035), .Z(n57037) );
  NOR U68960 ( .A(n57037), .B(n57036), .Z(n57042) );
  IV U68961 ( .A(n57038), .Z(n57040) );
  NOR U68962 ( .A(n57040), .B(n57039), .Z(n57041) );
  NOR U68963 ( .A(n57042), .B(n57041), .Z(n57043) );
  XOR U68964 ( .A(n57044), .B(n57043), .Z(n57045) );
  XOR U68965 ( .A(n57046), .B(n57045), .Z(n57047) );
  XOR U68966 ( .A(n57048), .B(n57047), .Z(n57049) );
  XOR U68967 ( .A(n57050), .B(n57049), .Z(n57073) );
  NOR U68968 ( .A(n57052), .B(n57051), .Z(n57071) );
  NOR U68969 ( .A(n57054), .B(n57053), .Z(n57059) );
  IV U68970 ( .A(n57055), .Z(n57056) );
  NOR U68971 ( .A(n57057), .B(n57056), .Z(n57058) );
  NOR U68972 ( .A(n57059), .B(n57058), .Z(n57069) );
  IV U68973 ( .A(n57060), .Z(n57061) );
  NOR U68974 ( .A(n57062), .B(n57061), .Z(n57067) );
  IV U68975 ( .A(n57063), .Z(n57065) );
  NOR U68976 ( .A(n57065), .B(n57064), .Z(n57066) );
  NOR U68977 ( .A(n57067), .B(n57066), .Z(n57068) );
  XOR U68978 ( .A(n57069), .B(n57068), .Z(n57070) );
  XOR U68979 ( .A(n57071), .B(n57070), .Z(n57072) );
  XOR U68980 ( .A(n57073), .B(n57072), .Z(n57079) );
  NOR U68981 ( .A(n57075), .B(n57074), .Z(n57077) );
  NOR U68982 ( .A(n57077), .B(n57076), .Z(n57078) );
  XOR U68983 ( .A(n57079), .B(n57078), .Z(n57080) );
  XOR U68984 ( .A(n57081), .B(n57080), .Z(n57082) );
  XOR U68985 ( .A(n57083), .B(n57082), .Z(n57098) );
  NOR U68986 ( .A(n57085), .B(n57084), .Z(n57096) );
  IV U68987 ( .A(n57086), .Z(n57088) );
  NOR U68988 ( .A(n57088), .B(n57087), .Z(n57093) );
  IV U68989 ( .A(n57089), .Z(n57090) );
  NOR U68990 ( .A(n57091), .B(n57090), .Z(n57092) );
  NOR U68991 ( .A(n57093), .B(n57092), .Z(n57094) );
  IV U68992 ( .A(n57094), .Z(n57095) );
  NOR U68993 ( .A(n57096), .B(n57095), .Z(n57097) );
  XOR U68994 ( .A(n57098), .B(n57097), .Z(n57108) );
  IV U68995 ( .A(n57102), .Z(n57099) );
  NOR U68996 ( .A(n57100), .B(n57099), .Z(n57106) );
  IV U68997 ( .A(n57100), .Z(n57101) );
  NOR U68998 ( .A(n57102), .B(n57101), .Z(n57103) );
  NOR U68999 ( .A(n57104), .B(n57103), .Z(n57105) );
  NOR U69000 ( .A(n57106), .B(n57105), .Z(n57107) );
  XOR U69001 ( .A(n57108), .B(n57107), .Z(n57124) );
  IV U69002 ( .A(n57109), .Z(n57111) );
  NOR U69003 ( .A(n57111), .B(n57110), .Z(n57122) );
  IV U69004 ( .A(n57112), .Z(n57113) );
  NOR U69005 ( .A(n57114), .B(n57113), .Z(n57119) );
  IV U69006 ( .A(n57115), .Z(n57117) );
  NOR U69007 ( .A(n57117), .B(n57116), .Z(n57118) );
  NOR U69008 ( .A(n57119), .B(n57118), .Z(n57120) );
  IV U69009 ( .A(n57120), .Z(n57121) );
  NOR U69010 ( .A(n57122), .B(n57121), .Z(n57123) );
  XOR U69011 ( .A(n57124), .B(n57123), .Z(n57134) );
  IV U69012 ( .A(n57125), .Z(n57126) );
  NOR U69013 ( .A(n57127), .B(n57126), .Z(n57132) );
  IV U69014 ( .A(n57128), .Z(n57129) );
  NOR U69015 ( .A(n57130), .B(n57129), .Z(n57131) );
  NOR U69016 ( .A(n57132), .B(n57131), .Z(n57133) );
  XOR U69017 ( .A(n57134), .B(n57133), .Z(n57145) );
  IV U69018 ( .A(n57138), .Z(n57135) );
  NOR U69019 ( .A(n57136), .B(n57135), .Z(n57143) );
  IV U69020 ( .A(n57137), .Z(n57141) );
  NOR U69021 ( .A(n57139), .B(n57138), .Z(n57140) );
  NOR U69022 ( .A(n57141), .B(n57140), .Z(n57142) );
  NOR U69023 ( .A(n57143), .B(n57142), .Z(n57144) );
  XOR U69024 ( .A(n57145), .B(n57144), .Z(n57146) );
  XOR U69025 ( .A(n57147), .B(n57146), .Z(n57148) );
  XOR U69026 ( .A(n57149), .B(n57148), .Z(n57156) );
  IV U69027 ( .A(n57150), .Z(n57152) );
  NOR U69028 ( .A(n57152), .B(n57151), .Z(n57153) );
  NOR U69029 ( .A(n57154), .B(n57153), .Z(n57155) );
  XOR U69030 ( .A(n57156), .B(n57155), .Z(n57157) );
  XOR U69031 ( .A(n57158), .B(n57157), .Z(n57159) );
  XOR U69032 ( .A(n57160), .B(n57159), .Z(n57170) );
  IV U69033 ( .A(n57161), .Z(n57162) );
  NOR U69034 ( .A(n57163), .B(n57162), .Z(n57168) );
  IV U69035 ( .A(n57164), .Z(n57165) );
  NOR U69036 ( .A(n57166), .B(n57165), .Z(n57167) );
  NOR U69037 ( .A(n57168), .B(n57167), .Z(n57169) );
  XOR U69038 ( .A(n57170), .B(n57169), .Z(n57185) );
  IV U69039 ( .A(n57171), .Z(n57173) );
  NOR U69040 ( .A(n57173), .B(n57172), .Z(n57183) );
  IV U69041 ( .A(n57174), .Z(n57175) );
  NOR U69042 ( .A(n57176), .B(n57175), .Z(n57181) );
  IV U69043 ( .A(n57177), .Z(n57178) );
  NOR U69044 ( .A(n57179), .B(n57178), .Z(n57180) );
  NOR U69045 ( .A(n57181), .B(n57180), .Z(n57182) );
  XOR U69046 ( .A(n57183), .B(n57182), .Z(n57184) );
  XOR U69047 ( .A(n57185), .B(n57184), .Z(n57186) );
  XOR U69048 ( .A(n57187), .B(n57186), .Z(n57205) );
  IV U69049 ( .A(n57188), .Z(n57190) );
  NOR U69050 ( .A(n57190), .B(n57189), .Z(n57194) );
  NOR U69051 ( .A(n57192), .B(n57191), .Z(n57193) );
  NOR U69052 ( .A(n57194), .B(n57193), .Z(n57203) );
  IV U69053 ( .A(n57195), .Z(n57197) );
  NOR U69054 ( .A(n57197), .B(n57196), .Z(n57201) );
  NOR U69055 ( .A(n57199), .B(n57198), .Z(n57200) );
  NOR U69056 ( .A(n57201), .B(n57200), .Z(n57202) );
  XOR U69057 ( .A(n57203), .B(n57202), .Z(n57204) );
  XOR U69058 ( .A(n57205), .B(n57204), .Z(n57215) );
  IV U69059 ( .A(n57206), .Z(n57207) );
  NOR U69060 ( .A(n57208), .B(n57207), .Z(n57213) );
  IV U69061 ( .A(n57209), .Z(n57210) );
  NOR U69062 ( .A(n57211), .B(n57210), .Z(n57212) );
  XOR U69063 ( .A(n57213), .B(n57212), .Z(n57214) );
  XOR U69064 ( .A(n57215), .B(n57214), .Z(n57225) );
  NOR U69065 ( .A(n57216), .B(n57217), .Z(n57223) );
  IV U69066 ( .A(n57216), .Z(n57219) );
  IV U69067 ( .A(n57217), .Z(n57218) );
  NOR U69068 ( .A(n57219), .B(n57218), .Z(n57220) );
  NOR U69069 ( .A(n57221), .B(n57220), .Z(n57222) );
  NOR U69070 ( .A(n57223), .B(n57222), .Z(n57224) );
  XOR U69071 ( .A(n57225), .B(n57224), .Z(n57236) );
  IV U69072 ( .A(n57226), .Z(n57227) );
  NOR U69073 ( .A(n57228), .B(n57227), .Z(n57234) );
  IV U69074 ( .A(n57229), .Z(n57232) );
  IV U69075 ( .A(n57230), .Z(n57231) );
  NOR U69076 ( .A(n57232), .B(n57231), .Z(n57233) );
  NOR U69077 ( .A(n57234), .B(n57233), .Z(n57235) );
  XOR U69078 ( .A(n57236), .B(n57235), .Z(n57237) );
  XOR U69079 ( .A(n57238), .B(n57237), .Z(n57239) );
  XOR U69080 ( .A(n57240), .B(n57239), .Z(n57241) );
  XOR U69081 ( .A(n57242), .B(n57241), .Z(n57243) );
  XOR U69082 ( .A(n57244), .B(n57243), .Z(n57263) );
  IV U69083 ( .A(n57245), .Z(n57247) );
  NOR U69084 ( .A(n57247), .B(n57246), .Z(n57252) );
  IV U69085 ( .A(n57248), .Z(n57249) );
  NOR U69086 ( .A(n57250), .B(n57249), .Z(n57251) );
  NOR U69087 ( .A(n57252), .B(n57251), .Z(n57261) );
  NOR U69088 ( .A(n57253), .B(n57254), .Z(n57259) );
  XOR U69089 ( .A(n57255), .B(n57254), .Z(n57256) );
  NOR U69090 ( .A(n57257), .B(n57256), .Z(n57258) );
  NOR U69091 ( .A(n57259), .B(n57258), .Z(n57260) );
  XOR U69092 ( .A(n57261), .B(n57260), .Z(n57262) );
  XOR U69093 ( .A(n57263), .B(n57262), .Z(n57264) );
  XOR U69094 ( .A(n57265), .B(n57264), .Z(n57266) );
  XOR U69095 ( .A(n57267), .B(n57266), .Z(n57313) );
  IV U69096 ( .A(n57268), .Z(n57270) );
  NOR U69097 ( .A(n57270), .B(n57269), .Z(n57275) );
  IV U69098 ( .A(n57271), .Z(n57273) );
  NOR U69099 ( .A(n57273), .B(n57272), .Z(n57274) );
  NOR U69100 ( .A(n57275), .B(n57274), .Z(n57285) );
  IV U69101 ( .A(n57276), .Z(n57278) );
  NOR U69102 ( .A(n57278), .B(n57277), .Z(n57283) );
  IV U69103 ( .A(n57279), .Z(n57280) );
  NOR U69104 ( .A(n57281), .B(n57280), .Z(n57282) );
  NOR U69105 ( .A(n57283), .B(n57282), .Z(n57284) );
  XOR U69106 ( .A(n57285), .B(n57284), .Z(n57311) );
  IV U69107 ( .A(n57286), .Z(n57288) );
  NOR U69108 ( .A(n57288), .B(n57287), .Z(n57302) );
  NOR U69109 ( .A(n57289), .B(n57291), .Z(n57290) );
  NOR U69110 ( .A(n57290), .B(n57296), .Z(n57300) );
  IV U69111 ( .A(n57291), .Z(n57293) );
  NOR U69112 ( .A(n57293), .B(n57292), .Z(n57294) );
  NOR U69113 ( .A(n57295), .B(n57294), .Z(n57298) );
  IV U69114 ( .A(n57296), .Z(n57297) );
  NOR U69115 ( .A(n57298), .B(n57297), .Z(n57299) );
  NOR U69116 ( .A(n57300), .B(n57299), .Z(n57301) );
  NOR U69117 ( .A(n57302), .B(n57301), .Z(n57309) );
  IV U69118 ( .A(n57303), .Z(n57304) );
  NOR U69119 ( .A(n57305), .B(n57304), .Z(n57307) );
  NOR U69120 ( .A(n57307), .B(n57306), .Z(n57308) );
  XOR U69121 ( .A(n57309), .B(n57308), .Z(n57310) );
  XOR U69122 ( .A(n57311), .B(n57310), .Z(n57312) );
  XOR U69123 ( .A(n57313), .B(n57312), .Z(n57314) );
  XOR U69124 ( .A(n57315), .B(n57314), .Z(n57335) );
  NOR U69125 ( .A(n57317), .B(n57316), .Z(n57333) );
  IV U69126 ( .A(n57318), .Z(n57319) );
  NOR U69127 ( .A(n57320), .B(n57319), .Z(n57324) );
  NOR U69128 ( .A(n57322), .B(n57321), .Z(n57323) );
  NOR U69129 ( .A(n57324), .B(n57323), .Z(n57331) );
  IV U69130 ( .A(n57325), .Z(n57326) );
  NOR U69131 ( .A(n57327), .B(n57326), .Z(n57329) );
  NOR U69132 ( .A(n57329), .B(n57328), .Z(n57330) );
  XOR U69133 ( .A(n57331), .B(n57330), .Z(n57332) );
  XOR U69134 ( .A(n57333), .B(n57332), .Z(n57334) );
  XOR U69135 ( .A(n57335), .B(n57334), .Z(n57355) );
  IV U69136 ( .A(n57347), .Z(n57341) );
  NOR U69137 ( .A(n57345), .B(n57341), .Z(n57351) );
  NOR U69138 ( .A(n57343), .B(n57342), .Z(n57344) );
  IV U69139 ( .A(n57344), .Z(n57349) );
  IV U69140 ( .A(n57345), .Z(n57346) );
  NOR U69141 ( .A(n57347), .B(n57346), .Z(n57348) );
  NOR U69142 ( .A(n57349), .B(n57348), .Z(n57350) );
  NOR U69143 ( .A(n57351), .B(n57350), .Z(n57352) );
  XOR U69144 ( .A(n57353), .B(n57352), .Z(n57354) );
  XOR U69145 ( .A(n57355), .B(n57354), .Z(n57356) );
  XOR U69146 ( .A(n57357), .B(n57356), .Z(n57382) );
  IV U69147 ( .A(n57358), .Z(n57360) );
  NOR U69148 ( .A(n57360), .B(n57359), .Z(n57380) );
  IV U69149 ( .A(n57361), .Z(n57362) );
  NOR U69150 ( .A(n57363), .B(n57362), .Z(n57368) );
  IV U69151 ( .A(n57364), .Z(n57366) );
  NOR U69152 ( .A(n57366), .B(n57365), .Z(n57367) );
  NOR U69153 ( .A(n57368), .B(n57367), .Z(n57378) );
  IV U69154 ( .A(n57369), .Z(n57371) );
  NOR U69155 ( .A(n57371), .B(n57370), .Z(n57376) );
  IV U69156 ( .A(n57372), .Z(n57373) );
  NOR U69157 ( .A(n57374), .B(n57373), .Z(n57375) );
  NOR U69158 ( .A(n57376), .B(n57375), .Z(n57377) );
  XOR U69159 ( .A(n57378), .B(n57377), .Z(n57379) );
  XOR U69160 ( .A(n57380), .B(n57379), .Z(n57381) );
  XOR U69161 ( .A(n57382), .B(n57381), .Z(n57383) );
  XOR U69162 ( .A(n57384), .B(n57383), .Z(n57399) );
  XOR U69163 ( .A(n57385), .B(n57389), .Z(n57386) );
  NOR U69164 ( .A(n57387), .B(n57386), .Z(n57397) );
  IV U69165 ( .A(n57388), .Z(n57390) );
  NOR U69166 ( .A(n57390), .B(n57389), .Z(n57395) );
  IV U69167 ( .A(n57391), .Z(n57392) );
  NOR U69168 ( .A(n57393), .B(n57392), .Z(n57394) );
  NOR U69169 ( .A(n57395), .B(n57394), .Z(n57396) );
  XOR U69170 ( .A(n57397), .B(n57396), .Z(n57398) );
  XOR U69171 ( .A(n57399), .B(n57398), .Z(n57400) );
  XOR U69172 ( .A(n57401), .B(n57400), .Z(n57402) );
  XOR U69173 ( .A(n57403), .B(n57402), .Z(n57427) );
  IV U69174 ( .A(n57404), .Z(n57405) );
  NOR U69175 ( .A(n57406), .B(n57405), .Z(n57416) );
  NOR U69176 ( .A(n57407), .B(n57408), .Z(n57414) );
  IV U69177 ( .A(n57407), .Z(n57410) );
  IV U69178 ( .A(n57408), .Z(n57409) );
  NOR U69179 ( .A(n57410), .B(n57409), .Z(n57412) );
  NOR U69180 ( .A(n57412), .B(n57411), .Z(n57413) );
  NOR U69181 ( .A(n57414), .B(n57413), .Z(n57415) );
  XOR U69182 ( .A(n57416), .B(n57415), .Z(n57425) );
  IV U69183 ( .A(n57417), .Z(n57419) );
  NOR U69184 ( .A(n57419), .B(n57418), .Z(n57423) );
  NOR U69185 ( .A(n57421), .B(n57420), .Z(n57422) );
  NOR U69186 ( .A(n57423), .B(n57422), .Z(n57424) );
  XOR U69187 ( .A(n57425), .B(n57424), .Z(n57426) );
  XOR U69188 ( .A(n57427), .B(n57426), .Z(n57436) );
  XOR U69189 ( .A(n57436), .B(n57435), .Z(n57447) );
  IV U69190 ( .A(n57437), .Z(n57438) );
  NOR U69191 ( .A(n57439), .B(n57438), .Z(n57445) );
  IV U69192 ( .A(n57440), .Z(n57443) );
  IV U69193 ( .A(n57441), .Z(n57442) );
  NOR U69194 ( .A(n57443), .B(n57442), .Z(n57444) );
  NOR U69195 ( .A(n57445), .B(n57444), .Z(n57446) );
  XOR U69196 ( .A(n57447), .B(n57446), .Z(n57466) );
  NOR U69197 ( .A(n57449), .B(n57448), .Z(n57450) );
  NOR U69198 ( .A(n57451), .B(n57450), .Z(n57464) );
  NOR U69199 ( .A(n57452), .B(n57456), .Z(n57462) );
  NOR U69200 ( .A(n57454), .B(n57453), .Z(n57459) );
  IV U69201 ( .A(n57455), .Z(n57457) );
  NOR U69202 ( .A(n57457), .B(n57456), .Z(n57458) );
  NOR U69203 ( .A(n57459), .B(n57458), .Z(n57460) );
  IV U69204 ( .A(n57460), .Z(n57461) );
  NOR U69205 ( .A(n57462), .B(n57461), .Z(n57463) );
  XOR U69206 ( .A(n57464), .B(n57463), .Z(n57465) );
  XOR U69207 ( .A(n57466), .B(n57465), .Z(n57467) );
  XOR U69208 ( .A(n57468), .B(n57467), .Z(n57481) );
  IV U69209 ( .A(n57469), .Z(n57470) );
  NOR U69210 ( .A(n57471), .B(n57470), .Z(n57476) );
  IV U69211 ( .A(n57472), .Z(n57474) );
  NOR U69212 ( .A(n57474), .B(n57473), .Z(n57475) );
  NOR U69213 ( .A(n57476), .B(n57475), .Z(n57477) );
  IV U69214 ( .A(n57477), .Z(n57478) );
  NOR U69215 ( .A(n57479), .B(n57478), .Z(n57480) );
  XOR U69216 ( .A(n57481), .B(n57480), .Z(n57482) );
  XOR U69217 ( .A(n57483), .B(n57482), .Z(n57484) );
  XOR U69218 ( .A(n57485), .B(n57484), .Z(n57486) );
  XOR U69219 ( .A(n57487), .B(n57486), .Z(n57488) );
  XOR U69220 ( .A(n57489), .B(n57488), .Z(n57490) );
  XOR U69221 ( .A(n57491), .B(n57490), .Z(n57492) );
  XOR U69222 ( .A(n57493), .B(n57492), .Z(n57494) );
  XOR U69223 ( .A(n57495), .B(n57494), .Z(n57496) );
  XOR U69224 ( .A(n57497), .B(n57496), .Z(n57518) );
  IV U69225 ( .A(n57498), .Z(n57500) );
  NOR U69226 ( .A(n57500), .B(n57499), .Z(n57502) );
  NOR U69227 ( .A(n57502), .B(n57501), .Z(n57508) );
  NOR U69228 ( .A(n57504), .B(n57503), .Z(n57505) );
  NOR U69229 ( .A(n57506), .B(n57505), .Z(n57507) );
  XOR U69230 ( .A(n57508), .B(n57507), .Z(n57516) );
  IV U69231 ( .A(n57509), .Z(n57510) );
  NOR U69232 ( .A(n57510), .B(n57512), .Z(n57514) );
  NOR U69233 ( .A(n57512), .B(n57511), .Z(n57513) );
  NOR U69234 ( .A(n57514), .B(n57513), .Z(n57515) );
  XOR U69235 ( .A(n57516), .B(n57515), .Z(n57517) );
  XOR U69236 ( .A(n57518), .B(n57517), .Z(n57519) );
  XOR U69237 ( .A(n57520), .B(n57519), .Z(n57521) );
  XOR U69238 ( .A(n57522), .B(n57521), .Z(n57523) );
  XOR U69239 ( .A(n57524), .B(n57523), .Z(n57536) );
  IV U69240 ( .A(n57528), .Z(n57526) );
  NOR U69241 ( .A(n57526), .B(n57525), .Z(n57534) );
  XOR U69242 ( .A(n57528), .B(n57527), .Z(n57529) );
  NOR U69243 ( .A(n57530), .B(n57529), .Z(n57532) );
  NOR U69244 ( .A(n57532), .B(n57531), .Z(n57533) );
  NOR U69245 ( .A(n57534), .B(n57533), .Z(n57535) );
  XOR U69246 ( .A(n57536), .B(n57535), .Z(n57537) );
  XOR U69247 ( .A(n57538), .B(n57537), .Z(n57539) );
  XOR U69248 ( .A(n57540), .B(n57539), .Z(n57541) );
  XOR U69249 ( .A(n57542), .B(n57541), .Z(n57543) );
  XOR U69250 ( .A(n57544), .B(n57543), .Z(n57545) );
  XOR U69251 ( .A(n57546), .B(n57545), .Z(n57547) );
  XOR U69252 ( .A(n57548), .B(n57547), .Z(n57568) );
  IV U69253 ( .A(n57549), .Z(n57551) );
  NOR U69254 ( .A(n57551), .B(n57550), .Z(n57556) );
  IV U69255 ( .A(n57552), .Z(n57554) );
  NOR U69256 ( .A(n57554), .B(n57553), .Z(n57555) );
  NOR U69257 ( .A(n57556), .B(n57555), .Z(n57566) );
  IV U69258 ( .A(n57557), .Z(n57559) );
  NOR U69259 ( .A(n57559), .B(n57558), .Z(n57564) );
  IV U69260 ( .A(n57560), .Z(n57562) );
  NOR U69261 ( .A(n57562), .B(n57561), .Z(n57563) );
  NOR U69262 ( .A(n57564), .B(n57563), .Z(n57565) );
  XOR U69263 ( .A(n57566), .B(n57565), .Z(n57567) );
  XOR U69264 ( .A(n57568), .B(n57567), .Z(n57569) );
  XOR U69265 ( .A(n57570), .B(n57569), .Z(n57571) );
  XOR U69266 ( .A(n57572), .B(n57571), .Z(n57573) );
  XOR U69267 ( .A(n57574), .B(n57573), .Z(n57575) );
  XOR U69268 ( .A(n57576), .B(n57575), .Z(n57577) );
  XOR U69269 ( .A(n57578), .B(n57577), .Z(n57597) );
  NOR U69270 ( .A(n57580), .B(n57579), .Z(n57585) );
  IV U69271 ( .A(n57581), .Z(n57583) );
  NOR U69272 ( .A(n57583), .B(n57582), .Z(n57584) );
  NOR U69273 ( .A(n57585), .B(n57584), .Z(n57595) );
  IV U69274 ( .A(n57586), .Z(n57588) );
  NOR U69275 ( .A(n57588), .B(n57587), .Z(n57593) );
  IV U69276 ( .A(n57589), .Z(n57590) );
  NOR U69277 ( .A(n57591), .B(n57590), .Z(n57592) );
  NOR U69278 ( .A(n57593), .B(n57592), .Z(n57594) );
  XOR U69279 ( .A(n57595), .B(n57594), .Z(n57596) );
  XOR U69280 ( .A(n57597), .B(n57596), .Z(n57598) );
  XOR U69281 ( .A(n57599), .B(n57598), .Z(n57609) );
  IV U69282 ( .A(n57600), .Z(n57601) );
  NOR U69283 ( .A(n57602), .B(n57601), .Z(n57607) );
  IV U69284 ( .A(n57603), .Z(n57604) );
  NOR U69285 ( .A(n57605), .B(n57604), .Z(n57606) );
  NOR U69286 ( .A(n57607), .B(n57606), .Z(n57608) );
  XOR U69287 ( .A(n57609), .B(n57608), .Z(n57619) );
  NOR U69288 ( .A(n57611), .B(n57610), .Z(n57617) );
  NOR U69289 ( .A(n57613), .B(n57612), .Z(n57615) );
  NOR U69290 ( .A(n57615), .B(n57614), .Z(n57616) );
  NOR U69291 ( .A(n57617), .B(n57616), .Z(n57618) );
  XOR U69292 ( .A(n57619), .B(n57618), .Z(n57620) );
  XOR U69293 ( .A(n57621), .B(n57620), .Z(n57622) );
  XOR U69294 ( .A(n57623), .B(n57622), .Z(n57624) );
  XOR U69295 ( .A(n57625), .B(n57624), .Z(n57626) );
  XOR U69296 ( .A(n57627), .B(n57626), .Z(n57628) );
  XOR U69297 ( .A(n57629), .B(n57628), .Z(n57630) );
  XOR U69298 ( .A(n57631), .B(n57630), .Z(n57658) );
  NOR U69299 ( .A(n57632), .B(n57635), .Z(n57633) );
  NOR U69300 ( .A(n57634), .B(n57633), .Z(n57639) );
  IV U69301 ( .A(n57635), .Z(n57636) );
  NOR U69302 ( .A(n57637), .B(n57636), .Z(n57638) );
  NOR U69303 ( .A(n57639), .B(n57638), .Z(n57656) );
  IV U69304 ( .A(n57640), .Z(n57641) );
  NOR U69305 ( .A(n57642), .B(n57641), .Z(n57646) );
  IV U69306 ( .A(n57643), .Z(n57644) );
  NOR U69307 ( .A(n57645), .B(n57644), .Z(n57652) );
  XOR U69308 ( .A(n57646), .B(n57652), .Z(n57654) );
  IV U69309 ( .A(n57647), .Z(n57649) );
  NOR U69310 ( .A(n57649), .B(n57648), .Z(n57650) );
  IV U69311 ( .A(n57650), .Z(n57651) );
  NOR U69312 ( .A(n57652), .B(n57651), .Z(n57653) );
  NOR U69313 ( .A(n57654), .B(n57653), .Z(n57655) );
  XOR U69314 ( .A(n57656), .B(n57655), .Z(n57657) );
  XOR U69315 ( .A(n57658), .B(n57657), .Z(n57659) );
  XOR U69316 ( .A(n57660), .B(n57659), .Z(n57686) );
  IV U69317 ( .A(n57661), .Z(n57662) );
  NOR U69318 ( .A(n57663), .B(n57662), .Z(n57667) );
  NOR U69319 ( .A(n57665), .B(n57664), .Z(n57666) );
  NOR U69320 ( .A(n57667), .B(n57666), .Z(n57673) );
  NOR U69321 ( .A(n57669), .B(n57668), .Z(n57671) );
  NOR U69322 ( .A(n57671), .B(n57670), .Z(n57672) );
  XOR U69323 ( .A(n57673), .B(n57672), .Z(n57684) );
  IV U69324 ( .A(n57678), .Z(n57675) );
  NOR U69325 ( .A(n57675), .B(n57674), .Z(n57682) );
  IV U69326 ( .A(n57676), .Z(n57680) );
  NOR U69327 ( .A(n57678), .B(n57677), .Z(n57679) );
  NOR U69328 ( .A(n57680), .B(n57679), .Z(n57681) );
  NOR U69329 ( .A(n57682), .B(n57681), .Z(n57683) );
  XOR U69330 ( .A(n57684), .B(n57683), .Z(n57685) );
  XOR U69331 ( .A(n57686), .B(n57685), .Z(n57687) );
  XOR U69332 ( .A(n57688), .B(n57687), .Z(n57698) );
  IV U69333 ( .A(n57689), .Z(n57691) );
  NOR U69334 ( .A(n57691), .B(n57690), .Z(n57696) );
  IV U69335 ( .A(n57692), .Z(n57693) );
  NOR U69336 ( .A(n57694), .B(n57693), .Z(n57695) );
  NOR U69337 ( .A(n57696), .B(n57695), .Z(n57697) );
  XOR U69338 ( .A(n57698), .B(n57697), .Z(n57715) );
  NOR U69339 ( .A(n57700), .B(n57699), .Z(n57701) );
  NOR U69340 ( .A(n57702), .B(n57701), .Z(n57703) );
  XOR U69341 ( .A(n57704), .B(n57703), .Z(n57713) );
  IV U69342 ( .A(n57705), .Z(n57706) );
  NOR U69343 ( .A(n57706), .B(n57708), .Z(n57711) );
  IV U69344 ( .A(n57707), .Z(n57709) );
  NOR U69345 ( .A(n57709), .B(n57708), .Z(n57710) );
  NOR U69346 ( .A(n57711), .B(n57710), .Z(n57712) );
  XOR U69347 ( .A(n57713), .B(n57712), .Z(n57714) );
  XOR U69348 ( .A(n57715), .B(n57714), .Z(n57716) );
  XOR U69349 ( .A(n57717), .B(n57716), .Z(n57730) );
  IV U69350 ( .A(n57718), .Z(n57721) );
  IV U69351 ( .A(n57719), .Z(n57720) );
  NOR U69352 ( .A(n57721), .B(n57720), .Z(n57728) );
  NOR U69353 ( .A(n57723), .B(n57722), .Z(n57724) );
  IV U69354 ( .A(n57724), .Z(n57726) );
  NOR U69355 ( .A(n57726), .B(n57725), .Z(n57727) );
  XOR U69356 ( .A(n57728), .B(n57727), .Z(n57729) );
  XOR U69357 ( .A(n57730), .B(n57729), .Z(n57731) );
  XOR U69358 ( .A(n57732), .B(n57731), .Z(n57733) );
  XOR U69359 ( .A(n57734), .B(n57733), .Z(n57735) );
  XOR U69360 ( .A(n57736), .B(n57735), .Z(n57737) );
  XOR U69361 ( .A(n57738), .B(n57737), .Z(n57739) );
  XOR U69362 ( .A(n57740), .B(n57739), .Z(n57776) );
  IV U69363 ( .A(n57741), .Z(n57742) );
  NOR U69364 ( .A(n57742), .B(n57760), .Z(n57747) );
  IV U69365 ( .A(n57743), .Z(n57744) );
  NOR U69366 ( .A(n57745), .B(n57744), .Z(n57746) );
  XOR U69367 ( .A(n57747), .B(n57746), .Z(n57774) );
  IV U69368 ( .A(n57748), .Z(n57749) );
  NOR U69369 ( .A(n57750), .B(n57749), .Z(n57755) );
  IV U69370 ( .A(n57751), .Z(n57752) );
  NOR U69371 ( .A(n57753), .B(n57752), .Z(n57754) );
  NOR U69372 ( .A(n57755), .B(n57754), .Z(n57772) );
  IV U69373 ( .A(n57756), .Z(n57758) );
  NOR U69374 ( .A(n57758), .B(n57757), .Z(n57762) );
  IV U69375 ( .A(n57759), .Z(n57761) );
  NOR U69376 ( .A(n57761), .B(n57760), .Z(n57768) );
  XOR U69377 ( .A(n57762), .B(n57768), .Z(n57770) );
  IV U69378 ( .A(n57763), .Z(n57765) );
  NOR U69379 ( .A(n57765), .B(n57764), .Z(n57766) );
  IV U69380 ( .A(n57766), .Z(n57767) );
  NOR U69381 ( .A(n57768), .B(n57767), .Z(n57769) );
  NOR U69382 ( .A(n57770), .B(n57769), .Z(n57771) );
  XOR U69383 ( .A(n57772), .B(n57771), .Z(n57773) );
  XOR U69384 ( .A(n57774), .B(n57773), .Z(n57775) );
  XOR U69385 ( .A(n57776), .B(n57775), .Z(n57791) );
  NOR U69386 ( .A(n57778), .B(n57777), .Z(n57789) );
  NOR U69387 ( .A(n57780), .B(n57779), .Z(n57787) );
  IV U69388 ( .A(n57781), .Z(n57783) );
  NOR U69389 ( .A(n57783), .B(n57782), .Z(n57785) );
  NOR U69390 ( .A(n57785), .B(n57784), .Z(n57786) );
  XOR U69391 ( .A(n57787), .B(n57786), .Z(n57788) );
  XOR U69392 ( .A(n57789), .B(n57788), .Z(n57790) );
  XOR U69393 ( .A(n57791), .B(n57790), .Z(n57808) );
  IV U69394 ( .A(n57794), .Z(n57792) );
  NOR U69395 ( .A(n57793), .B(n57792), .Z(n57802) );
  IV U69396 ( .A(n57793), .Z(n57795) );
  NOR U69397 ( .A(n57795), .B(n57794), .Z(n57800) );
  NOR U69398 ( .A(n57797), .B(n57796), .Z(n57798) );
  IV U69399 ( .A(n57798), .Z(n57799) );
  NOR U69400 ( .A(n57800), .B(n57799), .Z(n57801) );
  NOR U69401 ( .A(n57802), .B(n57801), .Z(n57806) );
  NOR U69402 ( .A(n57804), .B(n57803), .Z(n57805) );
  XOR U69403 ( .A(n57806), .B(n57805), .Z(n57807) );
  XOR U69404 ( .A(n57808), .B(n57807), .Z(n57813) );
  IV U69405 ( .A(n57809), .Z(n57810) );
  NOR U69406 ( .A(n57811), .B(n57810), .Z(n57812) );
  XOR U69407 ( .A(n57813), .B(n57812), .Z(n57814) );
  XOR U69408 ( .A(n57815), .B(n57814), .Z(n57816) );
  XOR U69409 ( .A(n57817), .B(n57816), .Z(n57829) );
  IV U69410 ( .A(n57818), .Z(n57819) );
  NOR U69411 ( .A(n57820), .B(n57819), .Z(n57827) );
  IV U69412 ( .A(n57821), .Z(n57823) );
  NOR U69413 ( .A(n57823), .B(n57822), .Z(n57825) );
  NOR U69414 ( .A(n57825), .B(n57824), .Z(n57826) );
  XOR U69415 ( .A(n57827), .B(n57826), .Z(n57828) );
  XOR U69416 ( .A(n57829), .B(n57828), .Z(n57830) );
  XOR U69417 ( .A(n57831), .B(n57830), .Z(n57832) );
  XOR U69418 ( .A(n57833), .B(n57832), .Z(n57834) );
  XOR U69419 ( .A(n57835), .B(n57834), .Z(n57836) );
  XOR U69420 ( .A(n57837), .B(n57836), .Z(n57838) );
  XOR U69421 ( .A(n57839), .B(n57838), .Z(n57840) );
  XOR U69422 ( .A(n57841), .B(n57840), .Z(n57842) );
  XOR U69423 ( .A(n57843), .B(n57842), .Z(n57844) );
  XOR U69424 ( .A(n57845), .B(n57844), .Z(n57876) );
  IV U69425 ( .A(n57846), .Z(n57848) );
  NOR U69426 ( .A(n57848), .B(n57847), .Z(n57853) );
  IV U69427 ( .A(n57849), .Z(n57850) );
  NOR U69428 ( .A(n57851), .B(n57850), .Z(n57852) );
  NOR U69429 ( .A(n57853), .B(n57852), .Z(n57864) );
  IV U69430 ( .A(n57858), .Z(n57854) );
  NOR U69431 ( .A(n57856), .B(n57854), .Z(n57862) );
  IV U69432 ( .A(n57855), .Z(n57860) );
  IV U69433 ( .A(n57856), .Z(n57857) );
  NOR U69434 ( .A(n57858), .B(n57857), .Z(n57859) );
  NOR U69435 ( .A(n57860), .B(n57859), .Z(n57861) );
  NOR U69436 ( .A(n57862), .B(n57861), .Z(n57863) );
  XOR U69437 ( .A(n57864), .B(n57863), .Z(n57874) );
  IV U69438 ( .A(n57865), .Z(n57867) );
  NOR U69439 ( .A(n57867), .B(n57866), .Z(n57872) );
  IV U69440 ( .A(n57868), .Z(n57870) );
  NOR U69441 ( .A(n57870), .B(n57869), .Z(n57871) );
  NOR U69442 ( .A(n57872), .B(n57871), .Z(n57873) );
  XOR U69443 ( .A(n57874), .B(n57873), .Z(n57875) );
  XOR U69444 ( .A(n57876), .B(n57875), .Z(n57877) );
  XOR U69445 ( .A(n57878), .B(n57877), .Z(n57891) );
  IV U69446 ( .A(n57879), .Z(n57881) );
  NOR U69447 ( .A(n57881), .B(n57880), .Z(n57882) );
  NOR U69448 ( .A(n57883), .B(n57882), .Z(n57889) );
  NOR U69449 ( .A(n57885), .B(n57884), .Z(n57886) );
  NOR U69450 ( .A(n57887), .B(n57886), .Z(n57888) );
  XOR U69451 ( .A(n57889), .B(n57888), .Z(n57890) );
  XOR U69452 ( .A(n57891), .B(n57890), .Z(n57892) );
  XOR U69453 ( .A(n57893), .B(n57892), .Z(n57912) );
  IV U69454 ( .A(n57894), .Z(n57895) );
  NOR U69455 ( .A(n57896), .B(n57895), .Z(n57901) );
  IV U69456 ( .A(n57897), .Z(n57899) );
  NOR U69457 ( .A(n57899), .B(n57898), .Z(n57900) );
  NOR U69458 ( .A(n57901), .B(n57900), .Z(n57910) );
  NOR U69459 ( .A(n57903), .B(n57902), .Z(n57908) );
  IV U69460 ( .A(n57904), .Z(n57906) );
  NOR U69461 ( .A(n57906), .B(n57905), .Z(n57907) );
  NOR U69462 ( .A(n57908), .B(n57907), .Z(n57909) );
  XOR U69463 ( .A(n57910), .B(n57909), .Z(n57911) );
  XOR U69464 ( .A(n57912), .B(n57911), .Z(n57913) );
  XOR U69465 ( .A(n57914), .B(n57913), .Z(n57915) );
  XOR U69466 ( .A(n57916), .B(n57915), .Z(n57917) );
  XOR U69467 ( .A(n57918), .B(n57917), .Z(n57919) );
  XOR U69468 ( .A(n57920), .B(n57919), .Z(n57921) );
  XOR U69469 ( .A(n57922), .B(n57921), .Z(n57923) );
  XOR U69470 ( .A(n57924), .B(n57923), .Z(n57957) );
  IV U69471 ( .A(n57925), .Z(n57927) );
  NOR U69472 ( .A(n57927), .B(n57926), .Z(n57929) );
  NOR U69473 ( .A(n57929), .B(n57928), .Z(n57945) );
  IV U69474 ( .A(n57930), .Z(n57932) );
  NOR U69475 ( .A(n57932), .B(n57931), .Z(n57943) );
  IV U69476 ( .A(n57933), .Z(n57935) );
  NOR U69477 ( .A(n57935), .B(n57934), .Z(n57940) );
  IV U69478 ( .A(n57936), .Z(n57938) );
  NOR U69479 ( .A(n57938), .B(n57937), .Z(n57939) );
  NOR U69480 ( .A(n57940), .B(n57939), .Z(n57941) );
  IV U69481 ( .A(n57941), .Z(n57942) );
  NOR U69482 ( .A(n57943), .B(n57942), .Z(n57944) );
  XOR U69483 ( .A(n57945), .B(n57944), .Z(n57955) );
  IV U69484 ( .A(n57946), .Z(n57948) );
  NOR U69485 ( .A(n57948), .B(n57947), .Z(n57953) );
  IV U69486 ( .A(n57949), .Z(n57951) );
  NOR U69487 ( .A(n57951), .B(n57950), .Z(n57952) );
  NOR U69488 ( .A(n57953), .B(n57952), .Z(n57954) );
  XOR U69489 ( .A(n57955), .B(n57954), .Z(n57956) );
  XOR U69490 ( .A(n57957), .B(n57956), .Z(n57958) );
  XOR U69491 ( .A(n57959), .B(n57958), .Z(n57973) );
  NOR U69492 ( .A(n57961), .B(n57960), .Z(n57971) );
  IV U69493 ( .A(n57962), .Z(n57964) );
  NOR U69494 ( .A(n57964), .B(n57963), .Z(n57969) );
  IV U69495 ( .A(n57965), .Z(n57967) );
  NOR U69496 ( .A(n57967), .B(n57966), .Z(n57968) );
  NOR U69497 ( .A(n57969), .B(n57968), .Z(n57970) );
  XOR U69498 ( .A(n57971), .B(n57970), .Z(n57972) );
  XOR U69499 ( .A(n57973), .B(n57972), .Z(n57974) );
  XOR U69500 ( .A(n57975), .B(n57974), .Z(n57989) );
  IV U69501 ( .A(n57976), .Z(n57978) );
  NOR U69502 ( .A(n57978), .B(n57977), .Z(n57983) );
  IV U69503 ( .A(n57979), .Z(n57980) );
  NOR U69504 ( .A(n57981), .B(n57980), .Z(n57982) );
  NOR U69505 ( .A(n57983), .B(n57982), .Z(n57987) );
  NOR U69506 ( .A(n57985), .B(n57984), .Z(n57986) );
  XOR U69507 ( .A(n57987), .B(n57986), .Z(n57988) );
  XOR U69508 ( .A(n57989), .B(n57988), .Z(n57990) );
  XOR U69509 ( .A(n57991), .B(n57990), .Z(n58016) );
  IV U69510 ( .A(n57992), .Z(n57994) );
  NOR U69511 ( .A(n57994), .B(n57993), .Z(n57999) );
  IV U69512 ( .A(n57995), .Z(n57997) );
  NOR U69513 ( .A(n57997), .B(n57996), .Z(n57998) );
  NOR U69514 ( .A(n57999), .B(n57998), .Z(n58005) );
  NOR U69515 ( .A(n58001), .B(n58000), .Z(n58003) );
  NOR U69516 ( .A(n58003), .B(n58002), .Z(n58004) );
  XOR U69517 ( .A(n58005), .B(n58004), .Z(n58014) );
  IV U69518 ( .A(n58006), .Z(n58007) );
  NOR U69519 ( .A(n58008), .B(n58007), .Z(n58012) );
  NOR U69520 ( .A(n58010), .B(n58009), .Z(n58011) );
  NOR U69521 ( .A(n58012), .B(n58011), .Z(n58013) );
  XOR U69522 ( .A(n58014), .B(n58013), .Z(n58015) );
  XOR U69523 ( .A(n58016), .B(n58015), .Z(n58032) );
  IV U69524 ( .A(n58017), .Z(n58019) );
  NOR U69525 ( .A(n58019), .B(n58018), .Z(n58030) );
  XOR U69526 ( .A(n58030), .B(n58029), .Z(n58031) );
  XOR U69527 ( .A(n58032), .B(n58031), .Z(n58042) );
  IV U69528 ( .A(n58033), .Z(n58034) );
  NOR U69529 ( .A(n58035), .B(n58034), .Z(n58040) );
  IV U69530 ( .A(n58036), .Z(n58038) );
  NOR U69531 ( .A(n58038), .B(n58037), .Z(n58039) );
  NOR U69532 ( .A(n58040), .B(n58039), .Z(n58041) );
  XOR U69533 ( .A(n58042), .B(n58041), .Z(n58059) );
  IV U69534 ( .A(n58043), .Z(n58044) );
  NOR U69535 ( .A(n58044), .B(n58070), .Z(n58050) );
  IV U69536 ( .A(n58045), .Z(n58048) );
  IV U69537 ( .A(n58046), .Z(n58047) );
  NOR U69538 ( .A(n58048), .B(n58047), .Z(n58049) );
  NOR U69539 ( .A(n58050), .B(n58049), .Z(n58057) );
  IV U69540 ( .A(n58051), .Z(n58052) );
  NOR U69541 ( .A(n58053), .B(n58052), .Z(n58054) );
  NOR U69542 ( .A(n58055), .B(n58054), .Z(n58056) );
  XOR U69543 ( .A(n58057), .B(n58056), .Z(n58058) );
  XOR U69544 ( .A(n58059), .B(n58058), .Z(n58060) );
  XOR U69545 ( .A(n58061), .B(n58060), .Z(n58075) );
  NOR U69546 ( .A(n58063), .B(n58062), .Z(n58067) );
  NOR U69547 ( .A(n58065), .B(n58064), .Z(n58066) );
  NOR U69548 ( .A(n58067), .B(n58066), .Z(n58073) );
  NOR U69549 ( .A(n58069), .B(n58068), .Z(n58071) );
  NOR U69550 ( .A(n58071), .B(n58070), .Z(n58072) );
  XOR U69551 ( .A(n58073), .B(n58072), .Z(n58074) );
  XOR U69552 ( .A(n58075), .B(n58074), .Z(n58076) );
  XOR U69553 ( .A(n58077), .B(n58076), .Z(n58078) );
  XOR U69554 ( .A(n58079), .B(n58078), .Z(n58080) );
  XOR U69555 ( .A(n58081), .B(n58080), .Z(n58082) );
  XOR U69556 ( .A(n58083), .B(n58082), .Z(n58105) );
  IV U69557 ( .A(n58084), .Z(n58086) );
  NOR U69558 ( .A(n58086), .B(n58085), .Z(n58088) );
  NOR U69559 ( .A(n58088), .B(n58087), .Z(n58103) );
  NOR U69560 ( .A(n58090), .B(n58089), .Z(n58101) );
  IV U69561 ( .A(n58091), .Z(n58092) );
  NOR U69562 ( .A(n58093), .B(n58092), .Z(n58098) );
  IV U69563 ( .A(n58094), .Z(n58096) );
  NOR U69564 ( .A(n58096), .B(n58095), .Z(n58097) );
  NOR U69565 ( .A(n58098), .B(n58097), .Z(n58099) );
  IV U69566 ( .A(n58099), .Z(n58100) );
  NOR U69567 ( .A(n58101), .B(n58100), .Z(n58102) );
  XOR U69568 ( .A(n58103), .B(n58102), .Z(n58104) );
  XOR U69569 ( .A(n58105), .B(n58104), .Z(n58106) );
  XOR U69570 ( .A(n58107), .B(n58106), .Z(n58131) );
  NOR U69571 ( .A(n58109), .B(n58108), .Z(n58120) );
  IV U69572 ( .A(n58109), .Z(n58111) );
  NOR U69573 ( .A(n58111), .B(n58110), .Z(n58118) );
  NOR U69574 ( .A(n58113), .B(n58112), .Z(n58114) );
  XOR U69575 ( .A(n58115), .B(n58114), .Z(n58116) );
  IV U69576 ( .A(n58116), .Z(n58117) );
  NOR U69577 ( .A(n58118), .B(n58117), .Z(n58119) );
  NOR U69578 ( .A(n58120), .B(n58119), .Z(n58129) );
  IV U69579 ( .A(n58121), .Z(n58122) );
  NOR U69580 ( .A(n58123), .B(n58122), .Z(n58127) );
  NOR U69581 ( .A(n58125), .B(n58124), .Z(n58126) );
  NOR U69582 ( .A(n58127), .B(n58126), .Z(n58128) );
  XOR U69583 ( .A(n58129), .B(n58128), .Z(n58130) );
  XOR U69584 ( .A(n58131), .B(n58130), .Z(n58132) );
  XOR U69585 ( .A(n58133), .B(n58132), .Z(n58134) );
  XOR U69586 ( .A(n58135), .B(n58134), .Z(n58136) );
  XOR U69587 ( .A(n58137), .B(n58136), .Z(n58173) );
  IV U69588 ( .A(n58138), .Z(n58139) );
  NOR U69589 ( .A(n58140), .B(n58139), .Z(n58151) );
  IV U69590 ( .A(n58141), .Z(n58143) );
  NOR U69591 ( .A(n58143), .B(n58142), .Z(n58148) );
  IV U69592 ( .A(n58144), .Z(n58146) );
  NOR U69593 ( .A(n58146), .B(n58145), .Z(n58147) );
  NOR U69594 ( .A(n58148), .B(n58147), .Z(n58149) );
  IV U69595 ( .A(n58149), .Z(n58150) );
  NOR U69596 ( .A(n58151), .B(n58150), .Z(n58171) );
  IV U69597 ( .A(n58155), .Z(n58152) );
  NOR U69598 ( .A(n58153), .B(n58152), .Z(n58159) );
  IV U69599 ( .A(n58153), .Z(n58154) );
  NOR U69600 ( .A(n58155), .B(n58154), .Z(n58157) );
  NOR U69601 ( .A(n58157), .B(n58156), .Z(n58158) );
  NOR U69602 ( .A(n58159), .B(n58158), .Z(n58169) );
  IV U69603 ( .A(n58160), .Z(n58161) );
  NOR U69604 ( .A(n58162), .B(n58161), .Z(n58167) );
  IV U69605 ( .A(n58163), .Z(n58164) );
  NOR U69606 ( .A(n58165), .B(n58164), .Z(n58166) );
  NOR U69607 ( .A(n58167), .B(n58166), .Z(n58168) );
  XOR U69608 ( .A(n58169), .B(n58168), .Z(n58170) );
  XOR U69609 ( .A(n58171), .B(n58170), .Z(n58172) );
  XOR U69610 ( .A(n58173), .B(n58172), .Z(n58174) );
  XOR U69611 ( .A(n58175), .B(n58174), .Z(n58204) );
  NOR U69612 ( .A(n58177), .B(n58176), .Z(n58182) );
  IV U69613 ( .A(n58178), .Z(n58179) );
  NOR U69614 ( .A(n58180), .B(n58179), .Z(n58181) );
  NOR U69615 ( .A(n58182), .B(n58181), .Z(n58202) );
  IV U69616 ( .A(n58183), .Z(n58184) );
  NOR U69617 ( .A(n58185), .B(n58184), .Z(n58190) );
  IV U69618 ( .A(n58186), .Z(n58187) );
  NOR U69619 ( .A(n58188), .B(n58187), .Z(n58189) );
  NOR U69620 ( .A(n58190), .B(n58189), .Z(n58200) );
  IV U69621 ( .A(n58191), .Z(n58192) );
  NOR U69622 ( .A(n58193), .B(n58192), .Z(n58198) );
  IV U69623 ( .A(n58194), .Z(n58195) );
  NOR U69624 ( .A(n58196), .B(n58195), .Z(n58197) );
  NOR U69625 ( .A(n58198), .B(n58197), .Z(n58199) );
  XOR U69626 ( .A(n58200), .B(n58199), .Z(n58201) );
  XOR U69627 ( .A(n58202), .B(n58201), .Z(n58203) );
  XOR U69628 ( .A(n58204), .B(n58203), .Z(n58234) );
  IV U69629 ( .A(n58220), .Z(n58205) );
  NOR U69630 ( .A(n58211), .B(n58205), .Z(n58206) );
  NOR U69631 ( .A(n58207), .B(n58206), .Z(n58208) );
  IV U69632 ( .A(n58208), .Z(n58209) );
  NOR U69633 ( .A(n58210), .B(n58209), .Z(n58214) );
  IV U69634 ( .A(n58211), .Z(n58212) );
  NOR U69635 ( .A(n58220), .B(n58212), .Z(n58213) );
  NOR U69636 ( .A(n58214), .B(n58213), .Z(n58222) );
  IV U69637 ( .A(n58215), .Z(n58216) );
  NOR U69638 ( .A(n58217), .B(n58216), .Z(n58218) );
  IV U69639 ( .A(n58218), .Z(n58219) );
  NOR U69640 ( .A(n58220), .B(n58219), .Z(n58221) );
  NOR U69641 ( .A(n58222), .B(n58221), .Z(n58232) );
  IV U69642 ( .A(n58223), .Z(n58224) );
  NOR U69643 ( .A(n58225), .B(n58224), .Z(n58230) );
  IV U69644 ( .A(n58226), .Z(n58228) );
  NOR U69645 ( .A(n58228), .B(n58227), .Z(n58229) );
  NOR U69646 ( .A(n58230), .B(n58229), .Z(n58231) );
  XOR U69647 ( .A(n58232), .B(n58231), .Z(n58233) );
  XOR U69648 ( .A(n58234), .B(n58233), .Z(n58235) );
  XOR U69649 ( .A(n58236), .B(n58235), .Z(n58237) );
  XOR U69650 ( .A(n58238), .B(n58237), .Z(n58254) );
  IV U69651 ( .A(n58239), .Z(n58241) );
  NOR U69652 ( .A(n58241), .B(n58240), .Z(n58252) );
  IV U69653 ( .A(n58242), .Z(n58244) );
  NOR U69654 ( .A(n58244), .B(n58243), .Z(n58249) );
  IV U69655 ( .A(n58245), .Z(n58247) );
  NOR U69656 ( .A(n58247), .B(n58246), .Z(n58248) );
  NOR U69657 ( .A(n58249), .B(n58248), .Z(n58250) );
  IV U69658 ( .A(n58250), .Z(n58251) );
  NOR U69659 ( .A(n58252), .B(n58251), .Z(n58253) );
  XOR U69660 ( .A(n58254), .B(n58253), .Z(n58264) );
  IV U69661 ( .A(n58255), .Z(n58257) );
  NOR U69662 ( .A(n58257), .B(n58256), .Z(n58262) );
  IV U69663 ( .A(n58258), .Z(n58259) );
  NOR U69664 ( .A(n58260), .B(n58259), .Z(n58261) );
  NOR U69665 ( .A(n58262), .B(n58261), .Z(n58263) );
  XOR U69666 ( .A(n58264), .B(n58263), .Z(n58265) );
  XOR U69667 ( .A(n58266), .B(n58265), .Z(n58267) );
  XOR U69668 ( .A(n58268), .B(n58267), .Z(n58269) );
  XOR U69669 ( .A(n58270), .B(n58269), .Z(n58271) );
  XOR U69670 ( .A(n58272), .B(n58271), .Z(n58301) );
  NOR U69671 ( .A(n58274), .B(n58273), .Z(n58275) );
  NOR U69672 ( .A(n58276), .B(n58275), .Z(n58288) );
  IV U69673 ( .A(n58277), .Z(n58279) );
  NOR U69674 ( .A(n58279), .B(n58278), .Z(n58286) );
  NOR U69675 ( .A(n58281), .B(n58280), .Z(n58283) );
  NOR U69676 ( .A(n58283), .B(n58282), .Z(n58284) );
  IV U69677 ( .A(n58284), .Z(n58285) );
  NOR U69678 ( .A(n58286), .B(n58285), .Z(n58287) );
  XOR U69679 ( .A(n58288), .B(n58287), .Z(n58299) );
  IV U69680 ( .A(n58289), .Z(n58290) );
  NOR U69681 ( .A(n58291), .B(n58290), .Z(n58297) );
  IV U69682 ( .A(n58292), .Z(n58295) );
  IV U69683 ( .A(n58293), .Z(n58294) );
  NOR U69684 ( .A(n58295), .B(n58294), .Z(n58296) );
  NOR U69685 ( .A(n58297), .B(n58296), .Z(n58298) );
  XOR U69686 ( .A(n58299), .B(n58298), .Z(n58300) );
  XOR U69687 ( .A(n58301), .B(n58300), .Z(n58302) );
  XOR U69688 ( .A(n58303), .B(n58302), .Z(n58322) );
  IV U69689 ( .A(n58304), .Z(n58306) );
  NOR U69690 ( .A(n58306), .B(n58305), .Z(n58310) );
  NOR U69691 ( .A(n58308), .B(n58307), .Z(n58309) );
  NOR U69692 ( .A(n58310), .B(n58309), .Z(n58320) );
  IV U69693 ( .A(n58311), .Z(n58313) );
  NOR U69694 ( .A(n58313), .B(n58312), .Z(n58318) );
  IV U69695 ( .A(n58314), .Z(n58316) );
  NOR U69696 ( .A(n58316), .B(n58315), .Z(n58317) );
  NOR U69697 ( .A(n58318), .B(n58317), .Z(n58319) );
  XOR U69698 ( .A(n58320), .B(n58319), .Z(n58321) );
  XOR U69699 ( .A(n58322), .B(n58321), .Z(n58323) );
  XOR U69700 ( .A(n58324), .B(n58323), .Z(n58340) );
  IV U69701 ( .A(n58325), .Z(n58326) );
  NOR U69702 ( .A(n58327), .B(n58326), .Z(n58338) );
  IV U69703 ( .A(n58328), .Z(n58329) );
  NOR U69704 ( .A(n58330), .B(n58329), .Z(n58335) );
  IV U69705 ( .A(n58331), .Z(n58333) );
  NOR U69706 ( .A(n58333), .B(n58332), .Z(n58334) );
  NOR U69707 ( .A(n58335), .B(n58334), .Z(n58336) );
  IV U69708 ( .A(n58336), .Z(n58337) );
  NOR U69709 ( .A(n58338), .B(n58337), .Z(n58339) );
  XOR U69710 ( .A(n58340), .B(n58339), .Z(n58347) );
  XOR U69711 ( .A(n58347), .B(n58346), .Z(n58363) );
  IV U69712 ( .A(n58348), .Z(n58350) );
  NOR U69713 ( .A(n58350), .B(n58349), .Z(n58361) );
  IV U69714 ( .A(n58351), .Z(n58353) );
  NOR U69715 ( .A(n58353), .B(n58352), .Z(n58358) );
  IV U69716 ( .A(n58354), .Z(n58356) );
  NOR U69717 ( .A(n58356), .B(n58355), .Z(n58357) );
  NOR U69718 ( .A(n58358), .B(n58357), .Z(n58359) );
  IV U69719 ( .A(n58359), .Z(n58360) );
  NOR U69720 ( .A(n58361), .B(n58360), .Z(n58362) );
  XOR U69721 ( .A(n58363), .B(n58362), .Z(n58390) );
  IV U69722 ( .A(n58364), .Z(n58365) );
  NOR U69723 ( .A(n58366), .B(n58365), .Z(n58367) );
  NOR U69724 ( .A(n58368), .B(n58367), .Z(n58378) );
  NOR U69725 ( .A(n58370), .B(n58369), .Z(n58376) );
  IV U69726 ( .A(n58371), .Z(n58374) );
  IV U69727 ( .A(n58372), .Z(n58373) );
  NOR U69728 ( .A(n58374), .B(n58373), .Z(n58375) );
  NOR U69729 ( .A(n58376), .B(n58375), .Z(n58377) );
  XOR U69730 ( .A(n58378), .B(n58377), .Z(n58388) );
  IV U69731 ( .A(n58382), .Z(n58380) );
  NOR U69732 ( .A(n58380), .B(n58379), .Z(n58386) );
  NOR U69733 ( .A(n58382), .B(n58381), .Z(n58383) );
  NOR U69734 ( .A(n58384), .B(n58383), .Z(n58385) );
  NOR U69735 ( .A(n58386), .B(n58385), .Z(n58387) );
  XOR U69736 ( .A(n58388), .B(n58387), .Z(n58389) );
  XOR U69737 ( .A(n58390), .B(n58389), .Z(n58391) );
  XOR U69738 ( .A(n58392), .B(n58391), .Z(n58393) );
  XOR U69739 ( .A(n58394), .B(n58393), .Z(n58395) );
  XOR U69740 ( .A(n58396), .B(n58395), .Z(n58397) );
  XOR U69741 ( .A(n58398), .B(n58397), .Z(n58399) );
  XOR U69742 ( .A(n58400), .B(n58399), .Z(n58435) );
  NOR U69743 ( .A(n58402), .B(n58401), .Z(n58404) );
  NOR U69744 ( .A(n58404), .B(n58403), .Z(n58405) );
  NOR U69745 ( .A(n58406), .B(n58405), .Z(n58433) );
  IV U69746 ( .A(n58407), .Z(n58408) );
  NOR U69747 ( .A(n58409), .B(n58408), .Z(n58420) );
  IV U69748 ( .A(n58410), .Z(n58411) );
  NOR U69749 ( .A(n58412), .B(n58411), .Z(n58417) );
  IV U69750 ( .A(n58413), .Z(n58414) );
  NOR U69751 ( .A(n58415), .B(n58414), .Z(n58416) );
  NOR U69752 ( .A(n58417), .B(n58416), .Z(n58418) );
  IV U69753 ( .A(n58418), .Z(n58419) );
  NOR U69754 ( .A(n58420), .B(n58419), .Z(n58431) );
  NOR U69755 ( .A(n58422), .B(n58421), .Z(n58423) );
  NOR U69756 ( .A(n58424), .B(n58423), .Z(n58429) );
  IV U69757 ( .A(n58425), .Z(n58426) );
  NOR U69758 ( .A(n58427), .B(n58426), .Z(n58428) );
  NOR U69759 ( .A(n58429), .B(n58428), .Z(n58430) );
  XOR U69760 ( .A(n58431), .B(n58430), .Z(n58432) );
  XOR U69761 ( .A(n58433), .B(n58432), .Z(n58434) );
  XOR U69762 ( .A(n58435), .B(n58434), .Z(n58436) );
  XOR U69763 ( .A(n58437), .B(n58436), .Z(n58438) );
  XOR U69764 ( .A(n58439), .B(n58438), .Z(n58440) );
  XOR U69765 ( .A(n58441), .B(n58440), .Z(n58442) );
  XOR U69766 ( .A(n58443), .B(n58442), .Z(n58444) );
  XOR U69767 ( .A(n58445), .B(n58444), .Z(n58446) );
  XOR U69768 ( .A(n58447), .B(n58446), .Z(n58448) );
  XOR U69769 ( .A(n58449), .B(n58448), .Z(n58450) );
  XOR U69770 ( .A(n58451), .B(n58450), .Z(n58452) );
  XOR U69771 ( .A(n58453), .B(n58452), .Z(n58454) );
  XOR U69772 ( .A(n58455), .B(n58454), .Z(n58475) );
  IV U69773 ( .A(n58456), .Z(n58458) );
  NOR U69774 ( .A(n58458), .B(n58457), .Z(n58463) );
  IV U69775 ( .A(n58459), .Z(n58460) );
  NOR U69776 ( .A(n58461), .B(n58460), .Z(n58462) );
  NOR U69777 ( .A(n58463), .B(n58462), .Z(n58473) );
  IV U69778 ( .A(n58464), .Z(n58466) );
  NOR U69779 ( .A(n58466), .B(n58465), .Z(n58471) );
  IV U69780 ( .A(n58467), .Z(n58468) );
  NOR U69781 ( .A(n58469), .B(n58468), .Z(n58470) );
  NOR U69782 ( .A(n58471), .B(n58470), .Z(n58472) );
  XOR U69783 ( .A(n58473), .B(n58472), .Z(n58474) );
  XOR U69784 ( .A(n58475), .B(n58474), .Z(n58510) );
  IV U69785 ( .A(n58476), .Z(n58477) );
  NOR U69786 ( .A(n58478), .B(n58477), .Z(n58483) );
  IV U69787 ( .A(n58479), .Z(n58481) );
  NOR U69788 ( .A(n58481), .B(n58480), .Z(n58482) );
  NOR U69789 ( .A(n58483), .B(n58482), .Z(n58492) );
  NOR U69790 ( .A(n58485), .B(n58484), .Z(n58490) );
  IV U69791 ( .A(n58486), .Z(n58487) );
  NOR U69792 ( .A(n58488), .B(n58487), .Z(n58489) );
  NOR U69793 ( .A(n58490), .B(n58489), .Z(n58491) );
  XOR U69794 ( .A(n58492), .B(n58491), .Z(n58508) );
  IV U69795 ( .A(n58493), .Z(n58494) );
  NOR U69796 ( .A(n58495), .B(n58494), .Z(n58506) );
  IV U69797 ( .A(n58496), .Z(n58498) );
  NOR U69798 ( .A(n58498), .B(n58497), .Z(n58503) );
  IV U69799 ( .A(n58499), .Z(n58501) );
  NOR U69800 ( .A(n58501), .B(n58500), .Z(n58502) );
  NOR U69801 ( .A(n58503), .B(n58502), .Z(n58504) );
  IV U69802 ( .A(n58504), .Z(n58505) );
  NOR U69803 ( .A(n58506), .B(n58505), .Z(n58507) );
  XOR U69804 ( .A(n58508), .B(n58507), .Z(n58509) );
  XOR U69805 ( .A(n58510), .B(n58509), .Z(n58511) );
  XOR U69806 ( .A(n58512), .B(n58511), .Z(n58549) );
  IV U69807 ( .A(n58513), .Z(n58514) );
  NOR U69808 ( .A(n58515), .B(n58514), .Z(n58525) );
  IV U69809 ( .A(n58516), .Z(n58517) );
  NOR U69810 ( .A(n58518), .B(n58517), .Z(n58522) );
  NOR U69811 ( .A(n58520), .B(n58519), .Z(n58521) );
  NOR U69812 ( .A(n58522), .B(n58521), .Z(n58523) );
  IV U69813 ( .A(n58523), .Z(n58524) );
  NOR U69814 ( .A(n58525), .B(n58524), .Z(n58536) );
  NOR U69815 ( .A(n58527), .B(n58526), .Z(n58534) );
  NOR U69816 ( .A(n58529), .B(n58528), .Z(n58530) );
  NOR U69817 ( .A(n58531), .B(n58530), .Z(n58532) );
  IV U69818 ( .A(n58532), .Z(n58533) );
  NOR U69819 ( .A(n58534), .B(n58533), .Z(n58535) );
  XOR U69820 ( .A(n58536), .B(n58535), .Z(n58547) );
  IV U69821 ( .A(n58540), .Z(n58537) );
  NOR U69822 ( .A(n58538), .B(n58537), .Z(n58545) );
  IV U69823 ( .A(n58539), .Z(n58543) );
  NOR U69824 ( .A(n58541), .B(n58540), .Z(n58542) );
  NOR U69825 ( .A(n58543), .B(n58542), .Z(n58544) );
  NOR U69826 ( .A(n58545), .B(n58544), .Z(n58546) );
  XOR U69827 ( .A(n58547), .B(n58546), .Z(n58548) );
  XOR U69828 ( .A(n58549), .B(n58548), .Z(n58576) );
  IV U69829 ( .A(n58550), .Z(n58552) );
  NOR U69830 ( .A(n58552), .B(n58551), .Z(n58557) );
  NOR U69831 ( .A(n58554), .B(n58553), .Z(n58555) );
  IV U69832 ( .A(n58555), .Z(n58556) );
  NOR U69833 ( .A(n58557), .B(n58556), .Z(n58574) );
  IV U69834 ( .A(n58558), .Z(n58559) );
  NOR U69835 ( .A(n58560), .B(n58559), .Z(n58572) );
  NOR U69836 ( .A(n58562), .B(n58561), .Z(n58569) );
  NOR U69837 ( .A(n58564), .B(n58563), .Z(n58567) );
  IV U69838 ( .A(n58565), .Z(n58566) );
  NOR U69839 ( .A(n58567), .B(n58566), .Z(n58568) );
  NOR U69840 ( .A(n58569), .B(n58568), .Z(n58570) );
  IV U69841 ( .A(n58570), .Z(n58571) );
  NOR U69842 ( .A(n58572), .B(n58571), .Z(n58573) );
  XOR U69843 ( .A(n58574), .B(n58573), .Z(n58575) );
  XOR U69844 ( .A(n58576), .B(n58575), .Z(n58617) );
  IV U69845 ( .A(n58577), .Z(n58578) );
  NOR U69846 ( .A(n58579), .B(n58578), .Z(n58595) );
  IV U69847 ( .A(n58580), .Z(n58582) );
  NOR U69848 ( .A(n58582), .B(n58581), .Z(n58587) );
  IV U69849 ( .A(n58583), .Z(n58585) );
  NOR U69850 ( .A(n58585), .B(n58584), .Z(n58586) );
  NOR U69851 ( .A(n58587), .B(n58586), .Z(n58588) );
  IV U69852 ( .A(n58588), .Z(n58590) );
  NOR U69853 ( .A(n58589), .B(n58590), .Z(n58593) );
  NOR U69854 ( .A(n58591), .B(n58590), .Z(n58592) );
  NOR U69855 ( .A(n58593), .B(n58592), .Z(n58594) );
  NOR U69856 ( .A(n58595), .B(n58594), .Z(n58615) );
  IV U69857 ( .A(n58596), .Z(n58597) );
  NOR U69858 ( .A(n58598), .B(n58597), .Z(n58603) );
  IV U69859 ( .A(n58599), .Z(n58600) );
  NOR U69860 ( .A(n58601), .B(n58600), .Z(n58602) );
  NOR U69861 ( .A(n58603), .B(n58602), .Z(n58613) );
  IV U69862 ( .A(n58604), .Z(n58606) );
  NOR U69863 ( .A(n58606), .B(n58605), .Z(n58611) );
  IV U69864 ( .A(n58607), .Z(n58609) );
  NOR U69865 ( .A(n58609), .B(n58608), .Z(n58610) );
  NOR U69866 ( .A(n58611), .B(n58610), .Z(n58612) );
  XOR U69867 ( .A(n58613), .B(n58612), .Z(n58614) );
  XOR U69868 ( .A(n58615), .B(n58614), .Z(n58616) );
  XOR U69869 ( .A(n58617), .B(n58616), .Z(n58627) );
  NOR U69870 ( .A(n58619), .B(n58618), .Z(n58625) );
  NOR U69871 ( .A(n58621), .B(n58620), .Z(n58623) );
  NOR U69872 ( .A(n58623), .B(n58622), .Z(n58624) );
  XOR U69873 ( .A(n58625), .B(n58624), .Z(n58626) );
  XOR U69874 ( .A(n58627), .B(n58626), .Z(n58628) );
  XOR U69875 ( .A(n58629), .B(n58628), .Z(n58630) );
  XOR U69876 ( .A(n58631), .B(n58630), .Z(n58632) );
  XOR U69877 ( .A(n58633), .B(n58632), .Z(n58642) );
  IV U69878 ( .A(n58634), .Z(n58635) );
  NOR U69879 ( .A(n58636), .B(n58635), .Z(n58640) );
  NOR U69880 ( .A(n58638), .B(n58637), .Z(n58639) );
  NOR U69881 ( .A(n58640), .B(n58639), .Z(n58641) );
  XOR U69882 ( .A(n58642), .B(n58641), .Z(n58643) );
  XOR U69883 ( .A(n58644), .B(n58643), .Z(n58645) );
  XOR U69884 ( .A(n58646), .B(n58645), .Z(n58662) );
  NOR U69885 ( .A(n58648), .B(n58647), .Z(n58653) );
  IV U69886 ( .A(n58649), .Z(n58650) );
  NOR U69887 ( .A(n58651), .B(n58650), .Z(n58652) );
  NOR U69888 ( .A(n58653), .B(n58652), .Z(n58660) );
  IV U69889 ( .A(n58654), .Z(n58655) );
  NOR U69890 ( .A(n58656), .B(n58655), .Z(n58657) );
  NOR U69891 ( .A(n58658), .B(n58657), .Z(n58659) );
  XOR U69892 ( .A(n58660), .B(n58659), .Z(n58661) );
  XOR U69893 ( .A(n58662), .B(n58661), .Z(n58663) );
  XOR U69894 ( .A(n58664), .B(n58663), .Z(n58683) );
  IV U69895 ( .A(n58665), .Z(n58667) );
  NOR U69896 ( .A(n58667), .B(n58666), .Z(n58672) );
  IV U69897 ( .A(n58668), .Z(n58669) );
  NOR U69898 ( .A(n58670), .B(n58669), .Z(n58671) );
  NOR U69899 ( .A(n58672), .B(n58671), .Z(n58681) );
  NOR U69900 ( .A(n58674), .B(n58673), .Z(n58679) );
  IV U69901 ( .A(n58675), .Z(n58677) );
  NOR U69902 ( .A(n58677), .B(n58676), .Z(n58678) );
  NOR U69903 ( .A(n58679), .B(n58678), .Z(n58680) );
  XOR U69904 ( .A(n58681), .B(n58680), .Z(n58682) );
  XOR U69905 ( .A(n58683), .B(n58682), .Z(n58684) );
  XOR U69906 ( .A(n58685), .B(n58684), .Z(n58686) );
  XOR U69907 ( .A(n58687), .B(n58686), .Z(n58688) );
  XOR U69908 ( .A(n58689), .B(n58688), .Z(o[10]) );
  NOR U69909 ( .A(n58691), .B(n58690), .Z(n58692) );
  XOR U69910 ( .A(n58693), .B(n58692), .Z(o[1]) );
  XOR U69911 ( .A(n58695), .B(n58694), .Z(o[2]) );
  NOR U69912 ( .A(n58697), .B(n58696), .Z(n58698) );
  XOR U69913 ( .A(n58699), .B(n58698), .Z(o[3]) );
  NOR U69914 ( .A(n58699), .B(n58698), .Z(n58700) );
  IV U69915 ( .A(n58700), .Z(n58701) );
  XOR U69916 ( .A(n58702), .B(n58701), .Z(o[4]) );
  NOR U69917 ( .A(n58702), .B(n58701), .Z(n58703) );
  NOR U69918 ( .A(n58704), .B(n58703), .Z(n58706) );
  XOR U69919 ( .A(n58706), .B(n58705), .Z(o[5]) );
  XOR U69920 ( .A(n58708), .B(n58707), .Z(o[6]) );
  NOR U69921 ( .A(n58710), .B(n58709), .Z(n58712) );
  XOR U69922 ( .A(n58712), .B(n58711), .Z(o[7]) );
  NOR U69923 ( .A(n58712), .B(n58711), .Z(n58713) );
  NOR U69924 ( .A(n58714), .B(n58713), .Z(n58715) );
  XOR U69925 ( .A(n58716), .B(n58715), .Z(o[8]) );
  XOR U69926 ( .A(n58718), .B(n58717), .Z(o[9]) );
endmodule

