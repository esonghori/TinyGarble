
module hamming_N1600_CC4 ( clk, rst, x, y, o );
  input [399:0] x;
  input [399:0] y;
  output [10:0] o;
  input clk, rst;
  wire   n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050;
  wire   [10:0] oglobal;

  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[0]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[1]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[2]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[3]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[4]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[5]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[6]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[7]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[8]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[9]) );
  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[10]) );
  XNOR U414 ( .A(n404), .B(n789), .Z(n410) );
  XNOR U415 ( .A(n470), .B(n471), .Z(n483) );
  XNOR U416 ( .A(n548), .B(n1017), .Z(n554) );
  XNOR U417 ( .A(n184), .B(n356), .Z(n186) );
  XNOR U418 ( .A(n262), .B(n508), .Z(n268) );
  XNOR U419 ( .A(n286), .B(n556), .Z(n292) );
  XNOR U420 ( .A(n335), .B(n652), .Z(n341) );
  XNOR U421 ( .A(n118), .B(n221), .Z(n124) );
  XNOR U422 ( .A(n168), .B(n319), .Z(n174) );
  XNOR U423 ( .A(n148), .B(n245), .Z(n131) );
  XNOR U424 ( .A(n373), .B(n676), .Z(n348) );
  XNOR U425 ( .A(n524), .B(n979), .Z(n530) );
  XNOR U426 ( .A(n494), .B(n495), .Z(n507) );
  XNOR U427 ( .A(n614), .B(n615), .Z(n627) );
  XNOR U428 ( .A(n662), .B(n663), .Z(n675) );
  XNOR U429 ( .A(n717), .B(n1283), .Z(n723) );
  XNOR U430 ( .A(n686), .B(n687), .Z(n699) );
  XNOR U431 ( .A(n237), .B(n460), .Z(n243) );
  XNOR U432 ( .A(n602), .B(n603), .Z(n610) );
  XNOR U433 ( .A(n650), .B(n651), .Z(n658) );
  XNOR U434 ( .A(n747), .B(n748), .Z(n755) );
  XNOR U435 ( .A(n1020), .B(n1022), .Z(n1041) );
  XNOR U436 ( .A(n1096), .B(n1098), .Z(n1117) );
  XNOR U437 ( .A(n192), .B(n368), .Z(n198) );
  XNOR U438 ( .A(n219), .B(n220), .Z(n227) );
  XNOR U439 ( .A(n417), .B(n418), .Z(n442) );
  XNOR U440 ( .A(n561), .B(n998), .Z(n537) );
  XNOR U441 ( .A(n811), .B(n813), .Z(n851) );
  XNOR U442 ( .A(n97), .B(n176), .Z(n103) );
  XNOR U443 ( .A(n275), .B(n484), .Z(n250) );
  XNOR U444 ( .A(n52), .B(n81), .Z(n58) );
  XNOR U445 ( .A(n348), .B(n580), .Z(n299) );
  XNOR U446 ( .A(n452), .B(n865), .Z(n458) );
  XNOR U447 ( .A(n500), .B(n941), .Z(n506) );
  XNOR U448 ( .A(n596), .B(n1093), .Z(n602) );
  XNOR U449 ( .A(n620), .B(n1131), .Z(n626) );
  XNOR U450 ( .A(n644), .B(n1169), .Z(n650) );
  XNOR U451 ( .A(n668), .B(n1207), .Z(n674) );
  XNOR U452 ( .A(n692), .B(n1245), .Z(n698) );
  XNOR U453 ( .A(n741), .B(n1321), .Z(n747) );
  XNOR U454 ( .A(n759), .B(n760), .Z(n772) );
  XNOR U455 ( .A(n213), .B(n412), .Z(n219) );
  XNOR U456 ( .A(n311), .B(n604), .Z(n317) );
  XNOR U457 ( .A(n530), .B(n960), .Z(n513) );
  XNOR U458 ( .A(n723), .B(n1264), .Z(n706) );
  XNOR U459 ( .A(n1058), .B(n1672), .Z(n1039) );
  XNOR U460 ( .A(n1324), .B(n1326), .Z(n1345) );
  XNOR U461 ( .A(n111), .B(n113), .Z(n125) );
  XNOR U462 ( .A(n142), .B(n270), .Z(n148) );
  XNOR U463 ( .A(n243), .B(n436), .Z(n226) );
  XNOR U464 ( .A(n341), .B(n628), .Z(n324) );
  XNOR U465 ( .A(n963), .B(n965), .Z(n1003) );
  XNOR U466 ( .A(n1267), .B(n1269), .Z(n1307) );
  XNOR U467 ( .A(n73), .B(n126), .Z(n79) );
  XNOR U468 ( .A(n198), .B(n343), .Z(n181) );
  XNOR U469 ( .A(n441), .B(n442), .Z(n490) );
  XNOR U470 ( .A(n849), .B(n851), .Z(n927) );
  XNOR U471 ( .A(n1153), .B(n1155), .Z(n1231) );
  XNOR U472 ( .A(n103), .B(n150), .Z(n86) );
  XNOR U473 ( .A(n681), .B(n1074), .Z(n585) );
  XOR U474 ( .A(oglobal[7]), .B(n40), .Z(n14) );
  XOR U475 ( .A(oglobal[4]), .B(n201), .Z(n20) );
  ANDN U476 ( .B(n1816), .A(n1175), .Z(n1177) );
  ANDN U477 ( .B(n2030), .A(n1365), .Z(n1367) );
  XNOR U478 ( .A(n229), .B(n448), .Z(n231) );
  XNOR U479 ( .A(n376), .B(n737), .Z(n378) );
  XNOR U480 ( .A(n542), .B(n543), .Z(n555) );
  XNOR U481 ( .A(n572), .B(n1055), .Z(n578) );
  XNOR U482 ( .A(n638), .B(n639), .Z(n651) );
  XNOR U483 ( .A(n711), .B(n712), .Z(n724) );
  XNOR U484 ( .A(n2018), .B(n2017), .Z(n2037) );
  XNOR U485 ( .A(n1997), .B(n1996), .Z(n1994) );
  XNOR U486 ( .A(n1955), .B(n1954), .Z(n1952) );
  XNOR U487 ( .A(n1913), .B(n1912), .Z(n1910) );
  XNOR U488 ( .A(n1871), .B(n1870), .Z(n1868) );
  XNOR U489 ( .A(n1806), .B(n1805), .Z(n1823) );
  XNOR U490 ( .A(n1764), .B(n1763), .Z(n1783) );
  XNOR U491 ( .A(n1745), .B(n1744), .Z(n1742) );
  XNOR U492 ( .A(n1619), .B(n1618), .Z(n1616) );
  XNOR U493 ( .A(n1577), .B(n1576), .Z(n1574) );
  XNOR U494 ( .A(n1537), .B(n1536), .Z(n1534) );
  XNOR U495 ( .A(n1493), .B(n1492), .Z(n1490) );
  XNOR U496 ( .A(n1453), .B(n1452), .Z(n1450) );
  XNOR U497 ( .A(n1411), .B(n1410), .Z(n1408) );
  XNOR U498 ( .A(n134), .B(n258), .Z(n136) );
  XNOR U499 ( .A(n304), .B(n306), .Z(n318) );
  XNOR U500 ( .A(n384), .B(n749), .Z(n390) );
  XNOR U501 ( .A(n434), .B(n808), .Z(n417) );
  XNOR U502 ( .A(n698), .B(n699), .Z(n707) );
  XNOR U503 ( .A(n868), .B(n870), .Z(n889) );
  XNOR U504 ( .A(n944), .B(n946), .Z(n965) );
  XNOR U505 ( .A(n1172), .B(n1174), .Z(n1193) );
  XNOR U506 ( .A(n292), .B(n532), .Z(n275) );
  XNOR U507 ( .A(n465), .B(n846), .Z(n441) );
  XNOR U508 ( .A(n754), .B(n1302), .Z(n730) );
  XNOR U509 ( .A(n1115), .B(n1117), .Z(n1155) );
  XNOR U510 ( .A(n66), .B(n68), .Z(n80) );
  XNOR U511 ( .A(n124), .B(n125), .Z(n132) );
  XNOR U512 ( .A(n226), .B(n227), .Z(n251) );
  XNOR U513 ( .A(n537), .B(n922), .Z(n489) );
  XNOR U514 ( .A(n633), .B(n634), .Z(n682) );
  XNOR U515 ( .A(n1305), .B(n1882), .Z(n1229) );
  XNOR U516 ( .A(n35), .B(n48), .Z(n37) );
  XNOR U517 ( .A(n181), .B(n294), .Z(n155) );
  XNOR U518 ( .A(n925), .B(n927), .Z(n1079) );
  XOR U519 ( .A(oglobal[6]), .B(n61), .Z(n16) );
  XOR U520 ( .A(oglobal[3]), .B(n393), .Z(n22) );
  ANDN U521 ( .B(n1442), .A(n833), .Z(n835) );
  ANDN U522 ( .B(n1526), .A(n909), .Z(n911) );
  XNOR U523 ( .A(n278), .B(n544), .Z(n280) );
  XNOR U524 ( .A(n327), .B(n640), .Z(n329) );
  XNOR U525 ( .A(n398), .B(n399), .Z(n411) );
  XNOR U526 ( .A(n422), .B(n423), .Z(n435) );
  XNOR U527 ( .A(n446), .B(n447), .Z(n459) );
  XNOR U528 ( .A(n518), .B(n519), .Z(n531) );
  XNOR U529 ( .A(n566), .B(n567), .Z(n579) );
  XNOR U530 ( .A(n590), .B(n591), .Z(n603) );
  XNOR U531 ( .A(n735), .B(n736), .Z(n748) );
  XNOR U532 ( .A(n765), .B(n1359), .Z(n771) );
  XNOR U533 ( .A(n1932), .B(n1931), .Z(n1951) );
  XNOR U534 ( .A(n1892), .B(n1891), .Z(n1909) );
  XNOR U535 ( .A(n1787), .B(n1786), .Z(n1784) );
  XNOR U536 ( .A(n1724), .B(n1723), .Z(n1741) );
  XNOR U537 ( .A(n1705), .B(n1704), .Z(n1702) );
  XNOR U538 ( .A(n1661), .B(n1660), .Z(n1658) );
  XNOR U539 ( .A(n1596), .B(n1595), .Z(n1615) );
  XNOR U540 ( .A(n1556), .B(n1555), .Z(n1573) );
  XNOR U541 ( .A(n1514), .B(n1513), .Z(n1533) );
  XNOR U542 ( .A(n1472), .B(n1471), .Z(n1489) );
  XNOR U543 ( .A(n1430), .B(n1429), .Z(n1449) );
  XNOR U544 ( .A(n1390), .B(n1389), .Z(n1407) );
  XNOR U545 ( .A(n255), .B(n257), .Z(n269) );
  XNOR U546 ( .A(n353), .B(n355), .Z(n367) );
  XNOR U547 ( .A(n482), .B(n884), .Z(n465) );
  XNOR U548 ( .A(n506), .B(n507), .Z(n514) );
  XNOR U549 ( .A(n554), .B(n555), .Z(n562) );
  XNOR U550 ( .A(n626), .B(n1112), .Z(n609) );
  XNOR U551 ( .A(n792), .B(n794), .Z(n813) );
  XNOR U552 ( .A(n1210), .B(n1838), .Z(n1191) );
  XNOR U553 ( .A(n1248), .B(n1250), .Z(n1269) );
  XNOR U554 ( .A(n1362), .B(n2008), .Z(n1343) );
  XNOR U555 ( .A(n390), .B(n725), .Z(n373) );
  XNOR U556 ( .A(n657), .B(n1150), .Z(n633) );
  XNOR U557 ( .A(n887), .B(n1462), .Z(n849) );
  XNOR U558 ( .A(n91), .B(n92), .Z(n104) );
  XNOR U559 ( .A(n174), .B(n175), .Z(n182) );
  XNOR U560 ( .A(n324), .B(n325), .Z(n349) );
  XNOR U561 ( .A(n730), .B(n1226), .Z(n681) );
  XNOR U562 ( .A(n1001), .B(n1546), .Z(n925) );
  XNOR U563 ( .A(n45), .B(n47), .Z(n59) );
  XNOR U564 ( .A(n79), .B(n80), .Z(n87) );
  XNOR U565 ( .A(n131), .B(n132), .Z(n156) );
  XNOR U566 ( .A(n250), .B(n251), .Z(n300) );
  XNOR U567 ( .A(n489), .B(n490), .Z(n586) );
  XNOR U568 ( .A(n1229), .B(n1714), .Z(n1077) );
  XOR U569 ( .A(oglobal[8]), .B(n32), .Z(n12) );
  XOR U570 ( .A(oglobal[5]), .B(n106), .Z(n18) );
  XOR U571 ( .A(oglobal[2]), .B(n774), .Z(n24) );
  ANDN U572 ( .B(n1400), .A(n795), .Z(n797) );
  ANDN U573 ( .B(n1482), .A(n871), .Z(n873) );
  ANDN U574 ( .B(n1566), .A(n947), .Z(n949) );
  ANDN U575 ( .B(n1608), .A(n985), .Z(n987) );
  ANDN U576 ( .B(n1650), .A(n1023), .Z(n1025) );
  ANDN U577 ( .B(n1694), .A(n1061), .Z(n1063) );
  ANDN U578 ( .B(n1734), .A(n1099), .Z(n1101) );
  ANDN U579 ( .B(n1776), .A(n1137), .Z(n1139) );
  ANDN U580 ( .B(n1860), .A(n1213), .Z(n1215) );
  ANDN U581 ( .B(n1902), .A(n1251), .Z(n1253) );
  ANDN U582 ( .B(n1944), .A(n1289), .Z(n1291) );
  ANDN U583 ( .B(n1986), .A(n1327), .Z(n1329) );
  XNOR U584 ( .A(n428), .B(n827), .Z(n434) );
  XNOR U585 ( .A(n476), .B(n903), .Z(n482) );
  XNOR U586 ( .A(n2041), .B(n2040), .Z(n2038) );
  XNOR U587 ( .A(n1976), .B(n1975), .Z(n1993) );
  XNOR U588 ( .A(n1848), .B(n1847), .Z(n1867) );
  XNOR U589 ( .A(n1827), .B(n1826), .Z(n1824) );
  XNOR U590 ( .A(n1682), .B(n1681), .Z(n1701) );
  XNOR U591 ( .A(n1640), .B(n1639), .Z(n1657) );
  XNOR U592 ( .A(n206), .B(n208), .Z(n220) );
  XNOR U593 ( .A(n231), .B(n232), .Z(n244) );
  XNOR U594 ( .A(n280), .B(n281), .Z(n293) );
  XNOR U595 ( .A(n329), .B(n330), .Z(n342) );
  XNOR U596 ( .A(n378), .B(n379), .Z(n391) );
  XNOR U597 ( .A(n410), .B(n411), .Z(n418) );
  XNOR U598 ( .A(n458), .B(n459), .Z(n466) );
  XNOR U599 ( .A(n578), .B(n1036), .Z(n561) );
  XNOR U600 ( .A(n674), .B(n1188), .Z(n657) );
  XNOR U601 ( .A(n771), .B(n1340), .Z(n754) );
  XNOR U602 ( .A(n830), .B(n1420), .Z(n811) );
  XNOR U603 ( .A(n906), .B(n1504), .Z(n887) );
  XNOR U604 ( .A(n982), .B(n1586), .Z(n963) );
  XNOR U605 ( .A(n1134), .B(n1754), .Z(n1115) );
  XNOR U606 ( .A(n1286), .B(n1922), .Z(n1267) );
  XNOR U607 ( .A(n136), .B(n137), .Z(n149) );
  XNOR U608 ( .A(n160), .B(n162), .Z(n175) );
  XNOR U609 ( .A(n186), .B(n187), .Z(n199) );
  XNOR U610 ( .A(n268), .B(n269), .Z(n276) );
  XNOR U611 ( .A(n317), .B(n318), .Z(n325) );
  XNOR U612 ( .A(n366), .B(n367), .Z(n374) );
  XNOR U613 ( .A(n513), .B(n514), .Z(n538) );
  XNOR U614 ( .A(n609), .B(n610), .Z(n634) );
  XNOR U615 ( .A(n706), .B(n707), .Z(n731) );
  XNOR U616 ( .A(n1039), .B(n1630), .Z(n1001) );
  XNOR U617 ( .A(n1191), .B(n1796), .Z(n1153) );
  XNOR U618 ( .A(n1343), .B(n1966), .Z(n1305) );
  XNOR U619 ( .A(n37), .B(n38), .Z(n15) );
  XNOR U620 ( .A(n58), .B(n59), .Z(n17) );
  XNOR U621 ( .A(n86), .B(n87), .Z(n19) );
  XNOR U622 ( .A(n155), .B(n156), .Z(n21) );
  XNOR U623 ( .A(n299), .B(n300), .Z(n23) );
  XNOR U624 ( .A(n585), .B(n586), .Z(n25) );
  XNOR U625 ( .A(n1077), .B(n1079), .Z(n27) );
  XNOR U626 ( .A(n12), .B(n13), .Z(o[8]) );
  XOR U627 ( .A(n14), .B(n15), .Z(o[7]) );
  XOR U628 ( .A(n16), .B(n17), .Z(o[6]) );
  XOR U629 ( .A(n18), .B(n19), .Z(o[5]) );
  XOR U630 ( .A(n20), .B(n21), .Z(o[4]) );
  XOR U631 ( .A(n22), .B(n23), .Z(o[3]) );
  XOR U632 ( .A(n24), .B(n25), .Z(o[2]) );
  XOR U633 ( .A(n26), .B(n27), .Z(o[1]) );
  XOR U634 ( .A(n28), .B(n29), .Z(o[10]) );
  XOR U635 ( .A(oglobal[10]), .B(n30), .Z(n29) );
  AND U636 ( .A(n28), .B(o[9]), .Z(n30) );
  XOR U637 ( .A(oglobal[9]), .B(n28), .Z(o[9]) );
  XNOR U638 ( .A(n31), .B(n32), .Z(n28) );
  ANDN U639 ( .B(n33), .A(n12), .Z(n31) );
  XNOR U640 ( .A(n32), .B(n13), .Z(n33) );
  XNOR U641 ( .A(n34), .B(n35), .Z(n13) );
  ANDN U642 ( .B(n36), .A(n37), .Z(n34) );
  XOR U643 ( .A(n35), .B(n38), .Z(n36) );
  XOR U644 ( .A(n39), .B(n40), .Z(n32) );
  ANDN U645 ( .B(n41), .A(n14), .Z(n39) );
  XOR U646 ( .A(n40), .B(n15), .Z(n41) );
  XNOR U647 ( .A(n42), .B(n43), .Z(n38) );
  ANDN U648 ( .B(n44), .A(n45), .Z(n42) );
  XOR U649 ( .A(n46), .B(n47), .Z(n44) );
  XNOR U650 ( .A(n49), .B(n50), .Z(n48) );
  ANDN U651 ( .B(n51), .A(n52), .Z(n49) );
  XNOR U652 ( .A(n53), .B(n54), .Z(n51) );
  XOR U653 ( .A(n55), .B(n56), .Z(n35) );
  ANDN U654 ( .B(n57), .A(n58), .Z(n55) );
  XOR U655 ( .A(n56), .B(n59), .Z(n57) );
  XOR U656 ( .A(n60), .B(n61), .Z(n40) );
  ANDN U657 ( .B(n62), .A(n16), .Z(n60) );
  XOR U658 ( .A(n61), .B(n17), .Z(n62) );
  XNOR U659 ( .A(n63), .B(n64), .Z(n47) );
  ANDN U660 ( .B(n65), .A(n66), .Z(n63) );
  XOR U661 ( .A(n67), .B(n68), .Z(n65) );
  XOR U662 ( .A(n43), .B(n69), .Z(n45) );
  XNOR U663 ( .A(n70), .B(n71), .Z(n69) );
  ANDN U664 ( .B(n72), .A(n73), .Z(n70) );
  XNOR U665 ( .A(n74), .B(n75), .Z(n72) );
  IV U666 ( .A(n46), .Z(n43) );
  XOR U667 ( .A(n76), .B(n77), .Z(n46) );
  ANDN U668 ( .B(n78), .A(n79), .Z(n76) );
  XOR U669 ( .A(n77), .B(n80), .Z(n78) );
  XNOR U670 ( .A(n53), .B(n82), .Z(n81) );
  IV U671 ( .A(n56), .Z(n82) );
  XOR U672 ( .A(n83), .B(n84), .Z(n56) );
  ANDN U673 ( .B(n85), .A(n86), .Z(n83) );
  XOR U674 ( .A(n84), .B(n87), .Z(n85) );
  XNOR U675 ( .A(n88), .B(n89), .Z(n53) );
  ANDN U676 ( .B(n90), .A(n91), .Z(n88) );
  XOR U677 ( .A(n89), .B(n92), .Z(n90) );
  XOR U678 ( .A(n50), .B(n93), .Z(n52) );
  XNOR U679 ( .A(n94), .B(n95), .Z(n93) );
  ANDN U680 ( .B(n96), .A(n97), .Z(n94) );
  XNOR U681 ( .A(n98), .B(n99), .Z(n96) );
  IV U682 ( .A(n54), .Z(n50) );
  XOR U683 ( .A(n100), .B(n101), .Z(n54) );
  ANDN U684 ( .B(n102), .A(n103), .Z(n100) );
  XOR U685 ( .A(n104), .B(n101), .Z(n102) );
  XOR U686 ( .A(n105), .B(n106), .Z(n61) );
  ANDN U687 ( .B(n107), .A(n18), .Z(n105) );
  XOR U688 ( .A(n106), .B(n19), .Z(n107) );
  XNOR U689 ( .A(n108), .B(n109), .Z(n68) );
  ANDN U690 ( .B(n110), .A(n111), .Z(n108) );
  XOR U691 ( .A(n112), .B(n113), .Z(n110) );
  XOR U692 ( .A(n64), .B(n114), .Z(n66) );
  XNOR U693 ( .A(n115), .B(n116), .Z(n114) );
  ANDN U694 ( .B(n117), .A(n118), .Z(n115) );
  XNOR U695 ( .A(n119), .B(n120), .Z(n117) );
  IV U696 ( .A(n67), .Z(n64) );
  XOR U697 ( .A(n121), .B(n122), .Z(n67) );
  ANDN U698 ( .B(n123), .A(n124), .Z(n121) );
  XOR U699 ( .A(n122), .B(n125), .Z(n123) );
  XNOR U700 ( .A(n74), .B(n127), .Z(n126) );
  IV U701 ( .A(n77), .Z(n127) );
  XOR U702 ( .A(n128), .B(n129), .Z(n77) );
  ANDN U703 ( .B(n130), .A(n131), .Z(n128) );
  XOR U704 ( .A(n129), .B(n132), .Z(n130) );
  XNOR U705 ( .A(n133), .B(n134), .Z(n74) );
  ANDN U706 ( .B(n135), .A(n136), .Z(n133) );
  XOR U707 ( .A(n134), .B(n137), .Z(n135) );
  XOR U708 ( .A(n71), .B(n138), .Z(n73) );
  XNOR U709 ( .A(n139), .B(n140), .Z(n138) );
  ANDN U710 ( .B(n141), .A(n142), .Z(n139) );
  XNOR U711 ( .A(n143), .B(n144), .Z(n141) );
  IV U712 ( .A(n75), .Z(n71) );
  XOR U713 ( .A(n145), .B(n146), .Z(n75) );
  ANDN U714 ( .B(n147), .A(n148), .Z(n145) );
  XOR U715 ( .A(n149), .B(n146), .Z(n147) );
  XOR U716 ( .A(n104), .B(n151), .Z(n150) );
  IV U717 ( .A(n84), .Z(n151) );
  XOR U718 ( .A(n152), .B(n153), .Z(n84) );
  ANDN U719 ( .B(n154), .A(n155), .Z(n152) );
  XOR U720 ( .A(n153), .B(n156), .Z(n154) );
  XNOR U721 ( .A(n157), .B(n158), .Z(n92) );
  ANDN U722 ( .B(n159), .A(n160), .Z(n157) );
  XOR U723 ( .A(n161), .B(n162), .Z(n159) );
  XOR U724 ( .A(n163), .B(n164), .Z(n91) );
  XNOR U725 ( .A(n165), .B(n166), .Z(n164) );
  ANDN U726 ( .B(n167), .A(n168), .Z(n165) );
  XNOR U727 ( .A(n169), .B(n170), .Z(n167) );
  IV U728 ( .A(n89), .Z(n163) );
  XOR U729 ( .A(n171), .B(n172), .Z(n89) );
  ANDN U730 ( .B(n173), .A(n174), .Z(n171) );
  XOR U731 ( .A(n172), .B(n175), .Z(n173) );
  XNOR U732 ( .A(n98), .B(n177), .Z(n176) );
  IV U733 ( .A(n101), .Z(n177) );
  XOR U734 ( .A(n178), .B(n179), .Z(n101) );
  ANDN U735 ( .B(n180), .A(n181), .Z(n178) );
  XOR U736 ( .A(n182), .B(n179), .Z(n180) );
  XNOR U737 ( .A(n183), .B(n184), .Z(n98) );
  ANDN U738 ( .B(n185), .A(n186), .Z(n183) );
  XOR U739 ( .A(n184), .B(n187), .Z(n185) );
  XOR U740 ( .A(n95), .B(n188), .Z(n97) );
  XNOR U741 ( .A(n189), .B(n190), .Z(n188) );
  ANDN U742 ( .B(n191), .A(n192), .Z(n189) );
  XNOR U743 ( .A(n193), .B(n194), .Z(n191) );
  IV U744 ( .A(n99), .Z(n95) );
  XOR U745 ( .A(n195), .B(n196), .Z(n99) );
  ANDN U746 ( .B(n197), .A(n198), .Z(n195) );
  XOR U747 ( .A(n199), .B(n196), .Z(n197) );
  XOR U748 ( .A(n200), .B(n201), .Z(n106) );
  ANDN U749 ( .B(n202), .A(n20), .Z(n200) );
  XOR U750 ( .A(n201), .B(n21), .Z(n202) );
  XNOR U751 ( .A(n203), .B(n204), .Z(n113) );
  ANDN U752 ( .B(n205), .A(n206), .Z(n203) );
  XOR U753 ( .A(n207), .B(n208), .Z(n205) );
  XOR U754 ( .A(n109), .B(n209), .Z(n111) );
  XNOR U755 ( .A(n210), .B(n211), .Z(n209) );
  ANDN U756 ( .B(n212), .A(n213), .Z(n210) );
  XNOR U757 ( .A(n214), .B(n215), .Z(n212) );
  IV U758 ( .A(n112), .Z(n109) );
  XOR U759 ( .A(n216), .B(n217), .Z(n112) );
  ANDN U760 ( .B(n218), .A(n219), .Z(n216) );
  XOR U761 ( .A(n217), .B(n220), .Z(n218) );
  XNOR U762 ( .A(n119), .B(n222), .Z(n221) );
  IV U763 ( .A(n122), .Z(n222) );
  XOR U764 ( .A(n223), .B(n224), .Z(n122) );
  ANDN U765 ( .B(n225), .A(n226), .Z(n223) );
  XOR U766 ( .A(n224), .B(n227), .Z(n225) );
  XNOR U767 ( .A(n228), .B(n229), .Z(n119) );
  ANDN U768 ( .B(n230), .A(n231), .Z(n228) );
  XOR U769 ( .A(n229), .B(n232), .Z(n230) );
  XOR U770 ( .A(n116), .B(n233), .Z(n118) );
  XNOR U771 ( .A(n234), .B(n235), .Z(n233) );
  ANDN U772 ( .B(n236), .A(n237), .Z(n234) );
  XNOR U773 ( .A(n238), .B(n239), .Z(n236) );
  IV U774 ( .A(n120), .Z(n116) );
  XOR U775 ( .A(n240), .B(n241), .Z(n120) );
  ANDN U776 ( .B(n242), .A(n243), .Z(n240) );
  XOR U777 ( .A(n244), .B(n241), .Z(n242) );
  XOR U778 ( .A(n149), .B(n246), .Z(n245) );
  IV U779 ( .A(n129), .Z(n246) );
  XOR U780 ( .A(n247), .B(n248), .Z(n129) );
  ANDN U781 ( .B(n249), .A(n250), .Z(n247) );
  XOR U782 ( .A(n248), .B(n251), .Z(n249) );
  XNOR U783 ( .A(n252), .B(n253), .Z(n137) );
  ANDN U784 ( .B(n254), .A(n255), .Z(n252) );
  XOR U785 ( .A(n256), .B(n257), .Z(n254) );
  XNOR U786 ( .A(n259), .B(n260), .Z(n258) );
  ANDN U787 ( .B(n261), .A(n262), .Z(n259) );
  XNOR U788 ( .A(n263), .B(n264), .Z(n261) );
  XOR U789 ( .A(n265), .B(n266), .Z(n134) );
  ANDN U790 ( .B(n267), .A(n268), .Z(n265) );
  XOR U791 ( .A(n266), .B(n269), .Z(n267) );
  XNOR U792 ( .A(n143), .B(n271), .Z(n270) );
  IV U793 ( .A(n146), .Z(n271) );
  XOR U794 ( .A(n272), .B(n273), .Z(n146) );
  ANDN U795 ( .B(n274), .A(n275), .Z(n272) );
  XOR U796 ( .A(n276), .B(n273), .Z(n274) );
  XNOR U797 ( .A(n277), .B(n278), .Z(n143) );
  ANDN U798 ( .B(n279), .A(n280), .Z(n277) );
  XOR U799 ( .A(n278), .B(n281), .Z(n279) );
  XOR U800 ( .A(n140), .B(n282), .Z(n142) );
  XNOR U801 ( .A(n283), .B(n284), .Z(n282) );
  ANDN U802 ( .B(n285), .A(n286), .Z(n283) );
  XNOR U803 ( .A(n287), .B(n288), .Z(n285) );
  IV U804 ( .A(n144), .Z(n140) );
  XOR U805 ( .A(n289), .B(n290), .Z(n144) );
  ANDN U806 ( .B(n291), .A(n292), .Z(n289) );
  XOR U807 ( .A(n293), .B(n290), .Z(n291) );
  XOR U808 ( .A(n182), .B(n295), .Z(n294) );
  IV U809 ( .A(n153), .Z(n295) );
  XOR U810 ( .A(n296), .B(n297), .Z(n153) );
  ANDN U811 ( .B(n298), .A(n299), .Z(n296) );
  XOR U812 ( .A(n297), .B(n300), .Z(n298) );
  XNOR U813 ( .A(n301), .B(n302), .Z(n162) );
  ANDN U814 ( .B(n303), .A(n304), .Z(n301) );
  XOR U815 ( .A(n305), .B(n306), .Z(n303) );
  XOR U816 ( .A(n158), .B(n307), .Z(n160) );
  XNOR U817 ( .A(n308), .B(n309), .Z(n307) );
  ANDN U818 ( .B(n310), .A(n311), .Z(n308) );
  XNOR U819 ( .A(n312), .B(n313), .Z(n310) );
  IV U820 ( .A(n161), .Z(n158) );
  XOR U821 ( .A(n314), .B(n315), .Z(n161) );
  ANDN U822 ( .B(n316), .A(n317), .Z(n314) );
  XOR U823 ( .A(n315), .B(n318), .Z(n316) );
  XNOR U824 ( .A(n169), .B(n320), .Z(n319) );
  IV U825 ( .A(n172), .Z(n320) );
  XOR U826 ( .A(n321), .B(n322), .Z(n172) );
  ANDN U827 ( .B(n323), .A(n324), .Z(n321) );
  XOR U828 ( .A(n322), .B(n325), .Z(n323) );
  XNOR U829 ( .A(n326), .B(n327), .Z(n169) );
  ANDN U830 ( .B(n328), .A(n329), .Z(n326) );
  XOR U831 ( .A(n327), .B(n330), .Z(n328) );
  XOR U832 ( .A(n166), .B(n331), .Z(n168) );
  XNOR U833 ( .A(n332), .B(n333), .Z(n331) );
  ANDN U834 ( .B(n334), .A(n335), .Z(n332) );
  XNOR U835 ( .A(n336), .B(n337), .Z(n334) );
  IV U836 ( .A(n170), .Z(n166) );
  XOR U837 ( .A(n338), .B(n339), .Z(n170) );
  ANDN U838 ( .B(n340), .A(n341), .Z(n338) );
  XOR U839 ( .A(n342), .B(n339), .Z(n340) );
  XOR U840 ( .A(n199), .B(n344), .Z(n343) );
  IV U841 ( .A(n179), .Z(n344) );
  XOR U842 ( .A(n345), .B(n346), .Z(n179) );
  ANDN U843 ( .B(n347), .A(n348), .Z(n345) );
  XOR U844 ( .A(n349), .B(n346), .Z(n347) );
  XNOR U845 ( .A(n350), .B(n351), .Z(n187) );
  ANDN U846 ( .B(n352), .A(n353), .Z(n350) );
  XOR U847 ( .A(n354), .B(n355), .Z(n352) );
  XNOR U848 ( .A(n357), .B(n358), .Z(n356) );
  ANDN U849 ( .B(n359), .A(n360), .Z(n357) );
  XNOR U850 ( .A(n361), .B(n362), .Z(n359) );
  XOR U851 ( .A(n363), .B(n364), .Z(n184) );
  ANDN U852 ( .B(n365), .A(n366), .Z(n363) );
  XOR U853 ( .A(n364), .B(n367), .Z(n365) );
  XNOR U854 ( .A(n193), .B(n369), .Z(n368) );
  IV U855 ( .A(n196), .Z(n369) );
  XOR U856 ( .A(n370), .B(n371), .Z(n196) );
  ANDN U857 ( .B(n372), .A(n373), .Z(n370) );
  XOR U858 ( .A(n374), .B(n371), .Z(n372) );
  XNOR U859 ( .A(n375), .B(n376), .Z(n193) );
  ANDN U860 ( .B(n377), .A(n378), .Z(n375) );
  XOR U861 ( .A(n376), .B(n379), .Z(n377) );
  XOR U862 ( .A(n190), .B(n380), .Z(n192) );
  XNOR U863 ( .A(n381), .B(n382), .Z(n380) );
  ANDN U864 ( .B(n383), .A(n384), .Z(n381) );
  XNOR U865 ( .A(n385), .B(n386), .Z(n383) );
  IV U866 ( .A(n194), .Z(n190) );
  XOR U867 ( .A(n387), .B(n388), .Z(n194) );
  ANDN U868 ( .B(n389), .A(n390), .Z(n387) );
  XOR U869 ( .A(n391), .B(n388), .Z(n389) );
  XOR U870 ( .A(n392), .B(n393), .Z(n201) );
  ANDN U871 ( .B(n394), .A(n22), .Z(n392) );
  XOR U872 ( .A(n393), .B(n23), .Z(n394) );
  XNOR U873 ( .A(n395), .B(n396), .Z(n208) );
  ANDN U874 ( .B(n397), .A(n398), .Z(n395) );
  XNOR U875 ( .A(n396), .B(n399), .Z(n397) );
  XOR U876 ( .A(n204), .B(n400), .Z(n206) );
  XNOR U877 ( .A(n401), .B(n402), .Z(n400) );
  ANDN U878 ( .B(n403), .A(n404), .Z(n401) );
  XNOR U879 ( .A(n405), .B(n406), .Z(n403) );
  IV U880 ( .A(n207), .Z(n204) );
  XOR U881 ( .A(n407), .B(n408), .Z(n207) );
  ANDN U882 ( .B(n409), .A(n410), .Z(n407) );
  XOR U883 ( .A(n408), .B(n411), .Z(n409) );
  XNOR U884 ( .A(n214), .B(n413), .Z(n412) );
  IV U885 ( .A(n217), .Z(n413) );
  XOR U886 ( .A(n414), .B(n415), .Z(n217) );
  ANDN U887 ( .B(n416), .A(n417), .Z(n414) );
  XOR U888 ( .A(n415), .B(n418), .Z(n416) );
  XOR U889 ( .A(n419), .B(n420), .Z(n214) );
  ANDN U890 ( .B(n421), .A(n422), .Z(n419) );
  XNOR U891 ( .A(n420), .B(n423), .Z(n421) );
  XOR U892 ( .A(n211), .B(n424), .Z(n213) );
  XNOR U893 ( .A(n425), .B(n426), .Z(n424) );
  ANDN U894 ( .B(n427), .A(n428), .Z(n425) );
  XNOR U895 ( .A(n429), .B(n430), .Z(n427) );
  IV U896 ( .A(n215), .Z(n211) );
  XOR U897 ( .A(n431), .B(n432), .Z(n215) );
  ANDN U898 ( .B(n433), .A(n434), .Z(n431) );
  XOR U899 ( .A(n435), .B(n432), .Z(n433) );
  XOR U900 ( .A(n244), .B(n437), .Z(n436) );
  IV U901 ( .A(n224), .Z(n437) );
  XOR U902 ( .A(n438), .B(n439), .Z(n224) );
  ANDN U903 ( .B(n440), .A(n441), .Z(n438) );
  XOR U904 ( .A(n439), .B(n442), .Z(n440) );
  XNOR U905 ( .A(n443), .B(n444), .Z(n232) );
  ANDN U906 ( .B(n445), .A(n446), .Z(n443) );
  XNOR U907 ( .A(n444), .B(n447), .Z(n445) );
  XNOR U908 ( .A(n449), .B(n450), .Z(n448) );
  ANDN U909 ( .B(n451), .A(n452), .Z(n449) );
  XNOR U910 ( .A(n453), .B(n454), .Z(n451) );
  XOR U911 ( .A(n455), .B(n456), .Z(n229) );
  ANDN U912 ( .B(n457), .A(n458), .Z(n455) );
  XOR U913 ( .A(n456), .B(n459), .Z(n457) );
  XNOR U914 ( .A(n238), .B(n461), .Z(n460) );
  IV U915 ( .A(n241), .Z(n461) );
  XOR U916 ( .A(n462), .B(n463), .Z(n241) );
  ANDN U917 ( .B(n464), .A(n465), .Z(n462) );
  XOR U918 ( .A(n466), .B(n463), .Z(n464) );
  XOR U919 ( .A(n467), .B(n468), .Z(n238) );
  ANDN U920 ( .B(n469), .A(n470), .Z(n467) );
  XNOR U921 ( .A(n468), .B(n471), .Z(n469) );
  XOR U922 ( .A(n235), .B(n472), .Z(n237) );
  XNOR U923 ( .A(n473), .B(n474), .Z(n472) );
  ANDN U924 ( .B(n475), .A(n476), .Z(n473) );
  XNOR U925 ( .A(n477), .B(n478), .Z(n475) );
  IV U926 ( .A(n239), .Z(n235) );
  XOR U927 ( .A(n479), .B(n480), .Z(n239) );
  ANDN U928 ( .B(n481), .A(n482), .Z(n479) );
  XOR U929 ( .A(n483), .B(n480), .Z(n481) );
  XOR U930 ( .A(n276), .B(n485), .Z(n484) );
  IV U931 ( .A(n248), .Z(n485) );
  XOR U932 ( .A(n486), .B(n487), .Z(n248) );
  ANDN U933 ( .B(n488), .A(n489), .Z(n486) );
  XOR U934 ( .A(n487), .B(n490), .Z(n488) );
  XNOR U935 ( .A(n491), .B(n492), .Z(n257) );
  ANDN U936 ( .B(n493), .A(n494), .Z(n491) );
  XNOR U937 ( .A(n492), .B(n495), .Z(n493) );
  XOR U938 ( .A(n253), .B(n496), .Z(n255) );
  XNOR U939 ( .A(n497), .B(n498), .Z(n496) );
  ANDN U940 ( .B(n499), .A(n500), .Z(n497) );
  XNOR U941 ( .A(n501), .B(n502), .Z(n499) );
  IV U942 ( .A(n256), .Z(n253) );
  XOR U943 ( .A(n503), .B(n504), .Z(n256) );
  ANDN U944 ( .B(n505), .A(n506), .Z(n503) );
  XOR U945 ( .A(n504), .B(n507), .Z(n505) );
  XNOR U946 ( .A(n263), .B(n509), .Z(n508) );
  IV U947 ( .A(n266), .Z(n509) );
  XOR U948 ( .A(n510), .B(n511), .Z(n266) );
  ANDN U949 ( .B(n512), .A(n513), .Z(n510) );
  XOR U950 ( .A(n511), .B(n514), .Z(n512) );
  XOR U951 ( .A(n515), .B(n516), .Z(n263) );
  ANDN U952 ( .B(n517), .A(n518), .Z(n515) );
  XNOR U953 ( .A(n516), .B(n519), .Z(n517) );
  XOR U954 ( .A(n260), .B(n520), .Z(n262) );
  XNOR U955 ( .A(n521), .B(n522), .Z(n520) );
  ANDN U956 ( .B(n523), .A(n524), .Z(n521) );
  XNOR U957 ( .A(n525), .B(n526), .Z(n523) );
  IV U958 ( .A(n264), .Z(n260) );
  XOR U959 ( .A(n527), .B(n528), .Z(n264) );
  ANDN U960 ( .B(n529), .A(n530), .Z(n527) );
  XOR U961 ( .A(n531), .B(n528), .Z(n529) );
  XOR U962 ( .A(n293), .B(n533), .Z(n532) );
  IV U963 ( .A(n273), .Z(n533) );
  XOR U964 ( .A(n534), .B(n535), .Z(n273) );
  ANDN U965 ( .B(n536), .A(n537), .Z(n534) );
  XOR U966 ( .A(n538), .B(n535), .Z(n536) );
  XNOR U967 ( .A(n539), .B(n540), .Z(n281) );
  ANDN U968 ( .B(n541), .A(n542), .Z(n539) );
  XNOR U969 ( .A(n540), .B(n543), .Z(n541) );
  XNOR U970 ( .A(n545), .B(n546), .Z(n544) );
  ANDN U971 ( .B(n547), .A(n548), .Z(n545) );
  XNOR U972 ( .A(n549), .B(n550), .Z(n547) );
  XOR U973 ( .A(n551), .B(n552), .Z(n278) );
  ANDN U974 ( .B(n553), .A(n554), .Z(n551) );
  XOR U975 ( .A(n552), .B(n555), .Z(n553) );
  XNOR U976 ( .A(n287), .B(n557), .Z(n556) );
  IV U977 ( .A(n290), .Z(n557) );
  XOR U978 ( .A(n558), .B(n559), .Z(n290) );
  ANDN U979 ( .B(n560), .A(n561), .Z(n558) );
  XOR U980 ( .A(n562), .B(n559), .Z(n560) );
  XOR U981 ( .A(n563), .B(n564), .Z(n287) );
  ANDN U982 ( .B(n565), .A(n566), .Z(n563) );
  XNOR U983 ( .A(n564), .B(n567), .Z(n565) );
  XOR U984 ( .A(n284), .B(n568), .Z(n286) );
  XNOR U985 ( .A(n569), .B(n570), .Z(n568) );
  ANDN U986 ( .B(n571), .A(n572), .Z(n569) );
  XNOR U987 ( .A(n573), .B(n574), .Z(n571) );
  IV U988 ( .A(n288), .Z(n284) );
  XOR U989 ( .A(n575), .B(n576), .Z(n288) );
  ANDN U990 ( .B(n577), .A(n578), .Z(n575) );
  XOR U991 ( .A(n579), .B(n576), .Z(n577) );
  XOR U992 ( .A(n349), .B(n581), .Z(n580) );
  IV U993 ( .A(n297), .Z(n581) );
  XOR U994 ( .A(n582), .B(n583), .Z(n297) );
  ANDN U995 ( .B(n584), .A(n585), .Z(n582) );
  XOR U996 ( .A(n583), .B(n586), .Z(n584) );
  XNOR U997 ( .A(n587), .B(n588), .Z(n306) );
  ANDN U998 ( .B(n589), .A(n590), .Z(n587) );
  XNOR U999 ( .A(n588), .B(n591), .Z(n589) );
  XOR U1000 ( .A(n302), .B(n592), .Z(n304) );
  XNOR U1001 ( .A(n593), .B(n594), .Z(n592) );
  ANDN U1002 ( .B(n595), .A(n596), .Z(n593) );
  XNOR U1003 ( .A(n597), .B(n598), .Z(n595) );
  IV U1004 ( .A(n305), .Z(n302) );
  XOR U1005 ( .A(n599), .B(n600), .Z(n305) );
  ANDN U1006 ( .B(n601), .A(n602), .Z(n599) );
  XOR U1007 ( .A(n600), .B(n603), .Z(n601) );
  XNOR U1008 ( .A(n312), .B(n605), .Z(n604) );
  IV U1009 ( .A(n315), .Z(n605) );
  XOR U1010 ( .A(n606), .B(n607), .Z(n315) );
  ANDN U1011 ( .B(n608), .A(n609), .Z(n606) );
  XOR U1012 ( .A(n607), .B(n610), .Z(n608) );
  XOR U1013 ( .A(n611), .B(n612), .Z(n312) );
  ANDN U1014 ( .B(n613), .A(n614), .Z(n611) );
  XNOR U1015 ( .A(n612), .B(n615), .Z(n613) );
  XOR U1016 ( .A(n309), .B(n616), .Z(n311) );
  XNOR U1017 ( .A(n617), .B(n618), .Z(n616) );
  ANDN U1018 ( .B(n619), .A(n620), .Z(n617) );
  XNOR U1019 ( .A(n621), .B(n622), .Z(n619) );
  IV U1020 ( .A(n313), .Z(n309) );
  XOR U1021 ( .A(n623), .B(n624), .Z(n313) );
  ANDN U1022 ( .B(n625), .A(n626), .Z(n623) );
  XOR U1023 ( .A(n627), .B(n624), .Z(n625) );
  XOR U1024 ( .A(n342), .B(n629), .Z(n628) );
  IV U1025 ( .A(n322), .Z(n629) );
  XOR U1026 ( .A(n630), .B(n631), .Z(n322) );
  ANDN U1027 ( .B(n632), .A(n633), .Z(n630) );
  XOR U1028 ( .A(n631), .B(n634), .Z(n632) );
  XNOR U1029 ( .A(n635), .B(n636), .Z(n330) );
  ANDN U1030 ( .B(n637), .A(n638), .Z(n635) );
  XNOR U1031 ( .A(n636), .B(n639), .Z(n637) );
  XNOR U1032 ( .A(n641), .B(n642), .Z(n640) );
  ANDN U1033 ( .B(n643), .A(n644), .Z(n641) );
  XNOR U1034 ( .A(n645), .B(n646), .Z(n643) );
  XOR U1035 ( .A(n647), .B(n648), .Z(n327) );
  ANDN U1036 ( .B(n649), .A(n650), .Z(n647) );
  XOR U1037 ( .A(n648), .B(n651), .Z(n649) );
  XNOR U1038 ( .A(n336), .B(n653), .Z(n652) );
  IV U1039 ( .A(n339), .Z(n653) );
  XOR U1040 ( .A(n654), .B(n655), .Z(n339) );
  ANDN U1041 ( .B(n656), .A(n657), .Z(n654) );
  XOR U1042 ( .A(n658), .B(n655), .Z(n656) );
  XOR U1043 ( .A(n659), .B(n660), .Z(n336) );
  ANDN U1044 ( .B(n661), .A(n662), .Z(n659) );
  XNOR U1045 ( .A(n660), .B(n663), .Z(n661) );
  XOR U1046 ( .A(n333), .B(n664), .Z(n335) );
  XNOR U1047 ( .A(n665), .B(n666), .Z(n664) );
  ANDN U1048 ( .B(n667), .A(n668), .Z(n665) );
  XNOR U1049 ( .A(n669), .B(n670), .Z(n667) );
  IV U1050 ( .A(n337), .Z(n333) );
  XOR U1051 ( .A(n671), .B(n672), .Z(n337) );
  ANDN U1052 ( .B(n673), .A(n674), .Z(n671) );
  XOR U1053 ( .A(n675), .B(n672), .Z(n673) );
  XOR U1054 ( .A(n374), .B(n677), .Z(n676) );
  IV U1055 ( .A(n346), .Z(n677) );
  XOR U1056 ( .A(n678), .B(n679), .Z(n346) );
  ANDN U1057 ( .B(n680), .A(n681), .Z(n678) );
  XOR U1058 ( .A(n682), .B(n679), .Z(n680) );
  XNOR U1059 ( .A(n683), .B(n684), .Z(n355) );
  ANDN U1060 ( .B(n685), .A(n686), .Z(n683) );
  XNOR U1061 ( .A(n684), .B(n687), .Z(n685) );
  XOR U1062 ( .A(n351), .B(n688), .Z(n353) );
  XNOR U1063 ( .A(n689), .B(n690), .Z(n688) );
  ANDN U1064 ( .B(n691), .A(n692), .Z(n689) );
  XNOR U1065 ( .A(n693), .B(n694), .Z(n691) );
  IV U1066 ( .A(n354), .Z(n351) );
  XOR U1067 ( .A(n695), .B(n696), .Z(n354) );
  ANDN U1068 ( .B(n697), .A(n698), .Z(n695) );
  XOR U1069 ( .A(n696), .B(n699), .Z(n697) );
  XOR U1070 ( .A(n700), .B(n701), .Z(n366) );
  XNOR U1071 ( .A(n361), .B(n702), .Z(n701) );
  IV U1072 ( .A(n364), .Z(n702) );
  XOR U1073 ( .A(n703), .B(n704), .Z(n364) );
  ANDN U1074 ( .B(n705), .A(n706), .Z(n703) );
  XOR U1075 ( .A(n704), .B(n707), .Z(n705) );
  XOR U1076 ( .A(n708), .B(n709), .Z(n361) );
  ANDN U1077 ( .B(n710), .A(n711), .Z(n708) );
  XNOR U1078 ( .A(n709), .B(n712), .Z(n710) );
  IV U1079 ( .A(n360), .Z(n700) );
  XOR U1080 ( .A(n358), .B(n713), .Z(n360) );
  XNOR U1081 ( .A(n714), .B(n715), .Z(n713) );
  ANDN U1082 ( .B(n716), .A(n717), .Z(n714) );
  XNOR U1083 ( .A(n718), .B(n719), .Z(n716) );
  IV U1084 ( .A(n362), .Z(n358) );
  XOR U1085 ( .A(n720), .B(n721), .Z(n362) );
  ANDN U1086 ( .B(n722), .A(n723), .Z(n720) );
  XOR U1087 ( .A(n724), .B(n721), .Z(n722) );
  XOR U1088 ( .A(n391), .B(n726), .Z(n725) );
  IV U1089 ( .A(n371), .Z(n726) );
  XOR U1090 ( .A(n727), .B(n728), .Z(n371) );
  ANDN U1091 ( .B(n729), .A(n730), .Z(n727) );
  XOR U1092 ( .A(n731), .B(n728), .Z(n729) );
  XNOR U1093 ( .A(n732), .B(n733), .Z(n379) );
  ANDN U1094 ( .B(n734), .A(n735), .Z(n732) );
  XNOR U1095 ( .A(n733), .B(n736), .Z(n734) );
  XNOR U1096 ( .A(n738), .B(n739), .Z(n737) );
  ANDN U1097 ( .B(n740), .A(n741), .Z(n738) );
  XNOR U1098 ( .A(n742), .B(n743), .Z(n740) );
  XOR U1099 ( .A(n744), .B(n745), .Z(n376) );
  ANDN U1100 ( .B(n746), .A(n747), .Z(n744) );
  XOR U1101 ( .A(n745), .B(n748), .Z(n746) );
  XNOR U1102 ( .A(n385), .B(n750), .Z(n749) );
  IV U1103 ( .A(n388), .Z(n750) );
  XOR U1104 ( .A(n751), .B(n752), .Z(n388) );
  ANDN U1105 ( .B(n753), .A(n754), .Z(n751) );
  XOR U1106 ( .A(n755), .B(n752), .Z(n753) );
  XOR U1107 ( .A(n756), .B(n757), .Z(n385) );
  ANDN U1108 ( .B(n758), .A(n759), .Z(n756) );
  XNOR U1109 ( .A(n757), .B(n760), .Z(n758) );
  XOR U1110 ( .A(n382), .B(n761), .Z(n384) );
  XNOR U1111 ( .A(n762), .B(n763), .Z(n761) );
  ANDN U1112 ( .B(n764), .A(n765), .Z(n762) );
  XNOR U1113 ( .A(n766), .B(n767), .Z(n764) );
  IV U1114 ( .A(n386), .Z(n382) );
  XOR U1115 ( .A(n768), .B(n769), .Z(n386) );
  ANDN U1116 ( .B(n770), .A(n771), .Z(n768) );
  XOR U1117 ( .A(n772), .B(n769), .Z(n770) );
  XOR U1118 ( .A(n773), .B(n774), .Z(n393) );
  ANDN U1119 ( .B(n775), .A(n24), .Z(n773) );
  XOR U1120 ( .A(n774), .B(n25), .Z(n775) );
  XNOR U1121 ( .A(n776), .B(n777), .Z(n399) );
  NANDN U1122 ( .A(n778), .B(n779), .Z(n777) );
  NANDN U1123 ( .A(n780), .B(n776), .Z(n779) );
  XNOR U1124 ( .A(n781), .B(n396), .Z(n398) );
  XNOR U1125 ( .A(n782), .B(n783), .Z(n396) );
  NAND U1126 ( .A(n784), .B(n785), .Z(n783) );
  XNOR U1127 ( .A(n782), .B(n786), .Z(n784) );
  NOR U1128 ( .A(n787), .B(n788), .Z(n781) );
  XOR U1129 ( .A(n405), .B(n408), .Z(n789) );
  XNOR U1130 ( .A(n790), .B(n791), .Z(n408) );
  NANDN U1131 ( .A(n792), .B(n793), .Z(n791) );
  XOR U1132 ( .A(n790), .B(n794), .Z(n793) );
  XNOR U1133 ( .A(n795), .B(n796), .Z(n405) );
  NANDN U1134 ( .A(n797), .B(n798), .Z(n796) );
  NANDN U1135 ( .A(n795), .B(n799), .Z(n798) );
  XOR U1136 ( .A(n800), .B(n406), .Z(n404) );
  IV U1137 ( .A(n402), .Z(n406) );
  XNOR U1138 ( .A(n801), .B(n802), .Z(n402) );
  NAND U1139 ( .A(n803), .B(n804), .Z(n802) );
  XOR U1140 ( .A(n801), .B(n805), .Z(n803) );
  NOR U1141 ( .A(n806), .B(n807), .Z(n800) );
  XNOR U1142 ( .A(n435), .B(n415), .Z(n808) );
  XNOR U1143 ( .A(n809), .B(n810), .Z(n415) );
  NANDN U1144 ( .A(n811), .B(n812), .Z(n810) );
  XOR U1145 ( .A(n809), .B(n813), .Z(n812) );
  XNOR U1146 ( .A(n814), .B(n815), .Z(n423) );
  NANDN U1147 ( .A(n816), .B(n817), .Z(n815) );
  NANDN U1148 ( .A(n818), .B(n814), .Z(n817) );
  XNOR U1149 ( .A(n819), .B(n420), .Z(n422) );
  XNOR U1150 ( .A(n820), .B(n821), .Z(n420) );
  NAND U1151 ( .A(n822), .B(n823), .Z(n821) );
  XNOR U1152 ( .A(n820), .B(n824), .Z(n822) );
  NOR U1153 ( .A(n825), .B(n826), .Z(n819) );
  XOR U1154 ( .A(n429), .B(n432), .Z(n827) );
  XNOR U1155 ( .A(n828), .B(n829), .Z(n432) );
  NANDN U1156 ( .A(n830), .B(n831), .Z(n829) );
  XNOR U1157 ( .A(n828), .B(n832), .Z(n831) );
  XNOR U1158 ( .A(n833), .B(n834), .Z(n429) );
  NANDN U1159 ( .A(n835), .B(n836), .Z(n834) );
  NANDN U1160 ( .A(n833), .B(n837), .Z(n836) );
  XOR U1161 ( .A(n838), .B(n430), .Z(n428) );
  IV U1162 ( .A(n426), .Z(n430) );
  XNOR U1163 ( .A(n839), .B(n840), .Z(n426) );
  NAND U1164 ( .A(n841), .B(n842), .Z(n840) );
  XOR U1165 ( .A(n839), .B(n843), .Z(n841) );
  NOR U1166 ( .A(n844), .B(n845), .Z(n838) );
  XNOR U1167 ( .A(n466), .B(n439), .Z(n846) );
  XNOR U1168 ( .A(n847), .B(n848), .Z(n439) );
  NANDN U1169 ( .A(n849), .B(n850), .Z(n848) );
  XOR U1170 ( .A(n847), .B(n851), .Z(n850) );
  XNOR U1171 ( .A(n852), .B(n853), .Z(n447) );
  NANDN U1172 ( .A(n854), .B(n855), .Z(n853) );
  NANDN U1173 ( .A(n856), .B(n852), .Z(n855) );
  XNOR U1174 ( .A(n857), .B(n444), .Z(n446) );
  XNOR U1175 ( .A(n858), .B(n859), .Z(n444) );
  NAND U1176 ( .A(n860), .B(n861), .Z(n859) );
  XNOR U1177 ( .A(n858), .B(n862), .Z(n860) );
  NOR U1178 ( .A(n863), .B(n864), .Z(n857) );
  XOR U1179 ( .A(n453), .B(n456), .Z(n865) );
  XNOR U1180 ( .A(n866), .B(n867), .Z(n456) );
  NANDN U1181 ( .A(n868), .B(n869), .Z(n867) );
  XOR U1182 ( .A(n866), .B(n870), .Z(n869) );
  XNOR U1183 ( .A(n871), .B(n872), .Z(n453) );
  NANDN U1184 ( .A(n873), .B(n874), .Z(n872) );
  NANDN U1185 ( .A(n871), .B(n875), .Z(n874) );
  XOR U1186 ( .A(n876), .B(n454), .Z(n452) );
  IV U1187 ( .A(n450), .Z(n454) );
  XNOR U1188 ( .A(n877), .B(n878), .Z(n450) );
  NAND U1189 ( .A(n879), .B(n880), .Z(n878) );
  XOR U1190 ( .A(n877), .B(n881), .Z(n879) );
  NOR U1191 ( .A(n882), .B(n883), .Z(n876) );
  XNOR U1192 ( .A(n483), .B(n463), .Z(n884) );
  XNOR U1193 ( .A(n885), .B(n886), .Z(n463) );
  NANDN U1194 ( .A(n887), .B(n888), .Z(n886) );
  XOR U1195 ( .A(n885), .B(n889), .Z(n888) );
  XNOR U1196 ( .A(n890), .B(n891), .Z(n471) );
  NANDN U1197 ( .A(n892), .B(n893), .Z(n891) );
  NANDN U1198 ( .A(n894), .B(n890), .Z(n893) );
  XNOR U1199 ( .A(n895), .B(n468), .Z(n470) );
  XNOR U1200 ( .A(n896), .B(n897), .Z(n468) );
  NAND U1201 ( .A(n898), .B(n899), .Z(n897) );
  XNOR U1202 ( .A(n896), .B(n900), .Z(n898) );
  NOR U1203 ( .A(n901), .B(n902), .Z(n895) );
  XOR U1204 ( .A(n477), .B(n480), .Z(n903) );
  XNOR U1205 ( .A(n904), .B(n905), .Z(n480) );
  NANDN U1206 ( .A(n906), .B(n907), .Z(n905) );
  XNOR U1207 ( .A(n904), .B(n908), .Z(n907) );
  XNOR U1208 ( .A(n909), .B(n910), .Z(n477) );
  NANDN U1209 ( .A(n911), .B(n912), .Z(n910) );
  NANDN U1210 ( .A(n909), .B(n913), .Z(n912) );
  XOR U1211 ( .A(n914), .B(n478), .Z(n476) );
  IV U1212 ( .A(n474), .Z(n478) );
  XNOR U1213 ( .A(n915), .B(n916), .Z(n474) );
  NAND U1214 ( .A(n917), .B(n918), .Z(n916) );
  XOR U1215 ( .A(n915), .B(n919), .Z(n917) );
  NOR U1216 ( .A(n920), .B(n921), .Z(n914) );
  XNOR U1217 ( .A(n538), .B(n487), .Z(n922) );
  XNOR U1218 ( .A(n923), .B(n924), .Z(n487) );
  NANDN U1219 ( .A(n925), .B(n926), .Z(n924) );
  XOR U1220 ( .A(n923), .B(n927), .Z(n926) );
  XNOR U1221 ( .A(n928), .B(n929), .Z(n495) );
  NANDN U1222 ( .A(n930), .B(n931), .Z(n929) );
  NANDN U1223 ( .A(n932), .B(n928), .Z(n931) );
  XNOR U1224 ( .A(n933), .B(n492), .Z(n494) );
  XNOR U1225 ( .A(n934), .B(n935), .Z(n492) );
  NAND U1226 ( .A(n936), .B(n937), .Z(n935) );
  XNOR U1227 ( .A(n934), .B(n938), .Z(n936) );
  NOR U1228 ( .A(n939), .B(n940), .Z(n933) );
  XOR U1229 ( .A(n501), .B(n504), .Z(n941) );
  XNOR U1230 ( .A(n942), .B(n943), .Z(n504) );
  NANDN U1231 ( .A(n944), .B(n945), .Z(n943) );
  XOR U1232 ( .A(n942), .B(n946), .Z(n945) );
  XNOR U1233 ( .A(n947), .B(n948), .Z(n501) );
  NANDN U1234 ( .A(n949), .B(n950), .Z(n948) );
  NANDN U1235 ( .A(n947), .B(n951), .Z(n950) );
  XOR U1236 ( .A(n952), .B(n502), .Z(n500) );
  IV U1237 ( .A(n498), .Z(n502) );
  XNOR U1238 ( .A(n953), .B(n954), .Z(n498) );
  NAND U1239 ( .A(n955), .B(n956), .Z(n954) );
  XOR U1240 ( .A(n953), .B(n957), .Z(n955) );
  NOR U1241 ( .A(n958), .B(n959), .Z(n952) );
  XNOR U1242 ( .A(n531), .B(n511), .Z(n960) );
  XNOR U1243 ( .A(n961), .B(n962), .Z(n511) );
  NANDN U1244 ( .A(n963), .B(n964), .Z(n962) );
  XOR U1245 ( .A(n961), .B(n965), .Z(n964) );
  XNOR U1246 ( .A(n966), .B(n967), .Z(n519) );
  NANDN U1247 ( .A(n968), .B(n969), .Z(n967) );
  NANDN U1248 ( .A(n970), .B(n966), .Z(n969) );
  XNOR U1249 ( .A(n971), .B(n516), .Z(n518) );
  XNOR U1250 ( .A(n972), .B(n973), .Z(n516) );
  NAND U1251 ( .A(n974), .B(n975), .Z(n973) );
  XNOR U1252 ( .A(n972), .B(n976), .Z(n974) );
  NOR U1253 ( .A(n977), .B(n978), .Z(n971) );
  XOR U1254 ( .A(n525), .B(n528), .Z(n979) );
  XNOR U1255 ( .A(n980), .B(n981), .Z(n528) );
  NANDN U1256 ( .A(n982), .B(n983), .Z(n981) );
  XNOR U1257 ( .A(n980), .B(n984), .Z(n983) );
  XNOR U1258 ( .A(n985), .B(n986), .Z(n525) );
  NANDN U1259 ( .A(n987), .B(n988), .Z(n986) );
  NANDN U1260 ( .A(n985), .B(n989), .Z(n988) );
  XOR U1261 ( .A(n990), .B(n526), .Z(n524) );
  IV U1262 ( .A(n522), .Z(n526) );
  XNOR U1263 ( .A(n991), .B(n992), .Z(n522) );
  NAND U1264 ( .A(n993), .B(n994), .Z(n992) );
  XOR U1265 ( .A(n991), .B(n995), .Z(n993) );
  NOR U1266 ( .A(n996), .B(n997), .Z(n990) );
  XNOR U1267 ( .A(n562), .B(n535), .Z(n998) );
  XNOR U1268 ( .A(n999), .B(n1000), .Z(n535) );
  NANDN U1269 ( .A(n1001), .B(n1002), .Z(n1000) );
  XOR U1270 ( .A(n999), .B(n1003), .Z(n1002) );
  XNOR U1271 ( .A(n1004), .B(n1005), .Z(n543) );
  NANDN U1272 ( .A(n1006), .B(n1007), .Z(n1005) );
  NANDN U1273 ( .A(n1008), .B(n1004), .Z(n1007) );
  XNOR U1274 ( .A(n1009), .B(n540), .Z(n542) );
  XNOR U1275 ( .A(n1010), .B(n1011), .Z(n540) );
  NAND U1276 ( .A(n1012), .B(n1013), .Z(n1011) );
  XNOR U1277 ( .A(n1010), .B(n1014), .Z(n1012) );
  NOR U1278 ( .A(n1015), .B(n1016), .Z(n1009) );
  XOR U1279 ( .A(n549), .B(n552), .Z(n1017) );
  XNOR U1280 ( .A(n1018), .B(n1019), .Z(n552) );
  NANDN U1281 ( .A(n1020), .B(n1021), .Z(n1019) );
  XOR U1282 ( .A(n1018), .B(n1022), .Z(n1021) );
  XNOR U1283 ( .A(n1023), .B(n1024), .Z(n549) );
  NANDN U1284 ( .A(n1025), .B(n1026), .Z(n1024) );
  NANDN U1285 ( .A(n1023), .B(n1027), .Z(n1026) );
  XOR U1286 ( .A(n1028), .B(n550), .Z(n548) );
  IV U1287 ( .A(n546), .Z(n550) );
  XNOR U1288 ( .A(n1029), .B(n1030), .Z(n546) );
  NAND U1289 ( .A(n1031), .B(n1032), .Z(n1030) );
  XOR U1290 ( .A(n1029), .B(n1033), .Z(n1031) );
  NOR U1291 ( .A(n1034), .B(n1035), .Z(n1028) );
  XNOR U1292 ( .A(n579), .B(n559), .Z(n1036) );
  XNOR U1293 ( .A(n1037), .B(n1038), .Z(n559) );
  NANDN U1294 ( .A(n1039), .B(n1040), .Z(n1038) );
  XOR U1295 ( .A(n1037), .B(n1041), .Z(n1040) );
  XNOR U1296 ( .A(n1042), .B(n1043), .Z(n567) );
  NANDN U1297 ( .A(n1044), .B(n1045), .Z(n1043) );
  NANDN U1298 ( .A(n1046), .B(n1042), .Z(n1045) );
  XNOR U1299 ( .A(n1047), .B(n564), .Z(n566) );
  XNOR U1300 ( .A(n1048), .B(n1049), .Z(n564) );
  NAND U1301 ( .A(n1050), .B(n1051), .Z(n1049) );
  XNOR U1302 ( .A(n1048), .B(n1052), .Z(n1050) );
  NOR U1303 ( .A(n1053), .B(n1054), .Z(n1047) );
  XOR U1304 ( .A(n573), .B(n576), .Z(n1055) );
  XNOR U1305 ( .A(n1056), .B(n1057), .Z(n576) );
  NANDN U1306 ( .A(n1058), .B(n1059), .Z(n1057) );
  XNOR U1307 ( .A(n1056), .B(n1060), .Z(n1059) );
  XNOR U1308 ( .A(n1061), .B(n1062), .Z(n573) );
  NANDN U1309 ( .A(n1063), .B(n1064), .Z(n1062) );
  NANDN U1310 ( .A(n1061), .B(n1065), .Z(n1064) );
  XOR U1311 ( .A(n1066), .B(n574), .Z(n572) );
  IV U1312 ( .A(n570), .Z(n574) );
  XNOR U1313 ( .A(n1067), .B(n1068), .Z(n570) );
  NAND U1314 ( .A(n1069), .B(n1070), .Z(n1068) );
  XOR U1315 ( .A(n1067), .B(n1071), .Z(n1069) );
  NOR U1316 ( .A(n1072), .B(n1073), .Z(n1066) );
  XNOR U1317 ( .A(n682), .B(n583), .Z(n1074) );
  XNOR U1318 ( .A(n1075), .B(n1076), .Z(n583) );
  NANDN U1319 ( .A(n1077), .B(n1078), .Z(n1076) );
  XOR U1320 ( .A(n1075), .B(n1079), .Z(n1078) );
  XNOR U1321 ( .A(n1080), .B(n1081), .Z(n591) );
  NANDN U1322 ( .A(n1082), .B(n1083), .Z(n1081) );
  NANDN U1323 ( .A(n1084), .B(n1080), .Z(n1083) );
  XNOR U1324 ( .A(n1085), .B(n588), .Z(n590) );
  XNOR U1325 ( .A(n1086), .B(n1087), .Z(n588) );
  NAND U1326 ( .A(n1088), .B(n1089), .Z(n1087) );
  XNOR U1327 ( .A(n1086), .B(n1090), .Z(n1088) );
  NOR U1328 ( .A(n1091), .B(n1092), .Z(n1085) );
  XOR U1329 ( .A(n597), .B(n600), .Z(n1093) );
  XNOR U1330 ( .A(n1094), .B(n1095), .Z(n600) );
  NANDN U1331 ( .A(n1096), .B(n1097), .Z(n1095) );
  XOR U1332 ( .A(n1094), .B(n1098), .Z(n1097) );
  XNOR U1333 ( .A(n1099), .B(n1100), .Z(n597) );
  NANDN U1334 ( .A(n1101), .B(n1102), .Z(n1100) );
  NANDN U1335 ( .A(n1099), .B(n1103), .Z(n1102) );
  XOR U1336 ( .A(n1104), .B(n598), .Z(n596) );
  IV U1337 ( .A(n594), .Z(n598) );
  XNOR U1338 ( .A(n1105), .B(n1106), .Z(n594) );
  NAND U1339 ( .A(n1107), .B(n1108), .Z(n1106) );
  XOR U1340 ( .A(n1105), .B(n1109), .Z(n1107) );
  NOR U1341 ( .A(n1110), .B(n1111), .Z(n1104) );
  XNOR U1342 ( .A(n627), .B(n607), .Z(n1112) );
  XNOR U1343 ( .A(n1113), .B(n1114), .Z(n607) );
  NANDN U1344 ( .A(n1115), .B(n1116), .Z(n1114) );
  XOR U1345 ( .A(n1113), .B(n1117), .Z(n1116) );
  XNOR U1346 ( .A(n1118), .B(n1119), .Z(n615) );
  NANDN U1347 ( .A(n1120), .B(n1121), .Z(n1119) );
  NANDN U1348 ( .A(n1122), .B(n1118), .Z(n1121) );
  XNOR U1349 ( .A(n1123), .B(n612), .Z(n614) );
  XNOR U1350 ( .A(n1124), .B(n1125), .Z(n612) );
  NAND U1351 ( .A(n1126), .B(n1127), .Z(n1125) );
  XNOR U1352 ( .A(n1124), .B(n1128), .Z(n1126) );
  NOR U1353 ( .A(n1129), .B(n1130), .Z(n1123) );
  XOR U1354 ( .A(n621), .B(n624), .Z(n1131) );
  XNOR U1355 ( .A(n1132), .B(n1133), .Z(n624) );
  NANDN U1356 ( .A(n1134), .B(n1135), .Z(n1133) );
  XNOR U1357 ( .A(n1132), .B(n1136), .Z(n1135) );
  XNOR U1358 ( .A(n1137), .B(n1138), .Z(n621) );
  NANDN U1359 ( .A(n1139), .B(n1140), .Z(n1138) );
  NANDN U1360 ( .A(n1137), .B(n1141), .Z(n1140) );
  XOR U1361 ( .A(n1142), .B(n622), .Z(n620) );
  IV U1362 ( .A(n618), .Z(n622) );
  XNOR U1363 ( .A(n1143), .B(n1144), .Z(n618) );
  NAND U1364 ( .A(n1145), .B(n1146), .Z(n1144) );
  XOR U1365 ( .A(n1143), .B(n1147), .Z(n1145) );
  NOR U1366 ( .A(n1148), .B(n1149), .Z(n1142) );
  XNOR U1367 ( .A(n658), .B(n631), .Z(n1150) );
  XNOR U1368 ( .A(n1151), .B(n1152), .Z(n631) );
  NANDN U1369 ( .A(n1153), .B(n1154), .Z(n1152) );
  XOR U1370 ( .A(n1151), .B(n1155), .Z(n1154) );
  XNOR U1371 ( .A(n1156), .B(n1157), .Z(n639) );
  NANDN U1372 ( .A(n1158), .B(n1159), .Z(n1157) );
  NANDN U1373 ( .A(n1160), .B(n1156), .Z(n1159) );
  XNOR U1374 ( .A(n1161), .B(n636), .Z(n638) );
  XNOR U1375 ( .A(n1162), .B(n1163), .Z(n636) );
  NAND U1376 ( .A(n1164), .B(n1165), .Z(n1163) );
  XNOR U1377 ( .A(n1162), .B(n1166), .Z(n1164) );
  NOR U1378 ( .A(n1167), .B(n1168), .Z(n1161) );
  XOR U1379 ( .A(n645), .B(n648), .Z(n1169) );
  XNOR U1380 ( .A(n1170), .B(n1171), .Z(n648) );
  NANDN U1381 ( .A(n1172), .B(n1173), .Z(n1171) );
  XOR U1382 ( .A(n1170), .B(n1174), .Z(n1173) );
  XNOR U1383 ( .A(n1175), .B(n1176), .Z(n645) );
  NANDN U1384 ( .A(n1177), .B(n1178), .Z(n1176) );
  NANDN U1385 ( .A(n1175), .B(n1179), .Z(n1178) );
  XOR U1386 ( .A(n1180), .B(n646), .Z(n644) );
  IV U1387 ( .A(n642), .Z(n646) );
  XNOR U1388 ( .A(n1181), .B(n1182), .Z(n642) );
  NAND U1389 ( .A(n1183), .B(n1184), .Z(n1182) );
  XOR U1390 ( .A(n1181), .B(n1185), .Z(n1183) );
  NOR U1391 ( .A(n1186), .B(n1187), .Z(n1180) );
  XNOR U1392 ( .A(n675), .B(n655), .Z(n1188) );
  XNOR U1393 ( .A(n1189), .B(n1190), .Z(n655) );
  NANDN U1394 ( .A(n1191), .B(n1192), .Z(n1190) );
  XOR U1395 ( .A(n1189), .B(n1193), .Z(n1192) );
  XNOR U1396 ( .A(n1194), .B(n1195), .Z(n663) );
  NANDN U1397 ( .A(n1196), .B(n1197), .Z(n1195) );
  NANDN U1398 ( .A(n1198), .B(n1194), .Z(n1197) );
  XNOR U1399 ( .A(n1199), .B(n660), .Z(n662) );
  XNOR U1400 ( .A(n1200), .B(n1201), .Z(n660) );
  NAND U1401 ( .A(n1202), .B(n1203), .Z(n1201) );
  XNOR U1402 ( .A(n1200), .B(n1204), .Z(n1202) );
  NOR U1403 ( .A(n1205), .B(n1206), .Z(n1199) );
  XOR U1404 ( .A(n669), .B(n672), .Z(n1207) );
  XNOR U1405 ( .A(n1208), .B(n1209), .Z(n672) );
  NANDN U1406 ( .A(n1210), .B(n1211), .Z(n1209) );
  XNOR U1407 ( .A(n1208), .B(n1212), .Z(n1211) );
  XNOR U1408 ( .A(n1213), .B(n1214), .Z(n669) );
  NANDN U1409 ( .A(n1215), .B(n1216), .Z(n1214) );
  NANDN U1410 ( .A(n1213), .B(n1217), .Z(n1216) );
  XOR U1411 ( .A(n1218), .B(n670), .Z(n668) );
  IV U1412 ( .A(n666), .Z(n670) );
  XNOR U1413 ( .A(n1219), .B(n1220), .Z(n666) );
  NAND U1414 ( .A(n1221), .B(n1222), .Z(n1220) );
  XOR U1415 ( .A(n1219), .B(n1223), .Z(n1221) );
  NOR U1416 ( .A(n1224), .B(n1225), .Z(n1218) );
  XNOR U1417 ( .A(n731), .B(n679), .Z(n1226) );
  XNOR U1418 ( .A(n1227), .B(n1228), .Z(n679) );
  NANDN U1419 ( .A(n1229), .B(n1230), .Z(n1228) );
  XOR U1420 ( .A(n1227), .B(n1231), .Z(n1230) );
  XNOR U1421 ( .A(n1232), .B(n1233), .Z(n687) );
  NANDN U1422 ( .A(n1234), .B(n1235), .Z(n1233) );
  NANDN U1423 ( .A(n1236), .B(n1232), .Z(n1235) );
  XNOR U1424 ( .A(n1237), .B(n684), .Z(n686) );
  XNOR U1425 ( .A(n1238), .B(n1239), .Z(n684) );
  NAND U1426 ( .A(n1240), .B(n1241), .Z(n1239) );
  XNOR U1427 ( .A(n1238), .B(n1242), .Z(n1240) );
  NOR U1428 ( .A(n1243), .B(n1244), .Z(n1237) );
  XOR U1429 ( .A(n693), .B(n696), .Z(n1245) );
  XNOR U1430 ( .A(n1246), .B(n1247), .Z(n696) );
  NANDN U1431 ( .A(n1248), .B(n1249), .Z(n1247) );
  XOR U1432 ( .A(n1246), .B(n1250), .Z(n1249) );
  XNOR U1433 ( .A(n1251), .B(n1252), .Z(n693) );
  NANDN U1434 ( .A(n1253), .B(n1254), .Z(n1252) );
  NANDN U1435 ( .A(n1251), .B(n1255), .Z(n1254) );
  XOR U1436 ( .A(n1256), .B(n694), .Z(n692) );
  IV U1437 ( .A(n690), .Z(n694) );
  XNOR U1438 ( .A(n1257), .B(n1258), .Z(n690) );
  NAND U1439 ( .A(n1259), .B(n1260), .Z(n1258) );
  XOR U1440 ( .A(n1257), .B(n1261), .Z(n1259) );
  NOR U1441 ( .A(n1262), .B(n1263), .Z(n1256) );
  XNOR U1442 ( .A(n724), .B(n704), .Z(n1264) );
  XNOR U1443 ( .A(n1265), .B(n1266), .Z(n704) );
  NANDN U1444 ( .A(n1267), .B(n1268), .Z(n1266) );
  XOR U1445 ( .A(n1265), .B(n1269), .Z(n1268) );
  XNOR U1446 ( .A(n1270), .B(n1271), .Z(n712) );
  NANDN U1447 ( .A(n1272), .B(n1273), .Z(n1271) );
  NANDN U1448 ( .A(n1274), .B(n1270), .Z(n1273) );
  XNOR U1449 ( .A(n1275), .B(n709), .Z(n711) );
  XNOR U1450 ( .A(n1276), .B(n1277), .Z(n709) );
  NAND U1451 ( .A(n1278), .B(n1279), .Z(n1277) );
  XNOR U1452 ( .A(n1276), .B(n1280), .Z(n1278) );
  NOR U1453 ( .A(n1281), .B(n1282), .Z(n1275) );
  XOR U1454 ( .A(n718), .B(n721), .Z(n1283) );
  XNOR U1455 ( .A(n1284), .B(n1285), .Z(n721) );
  NANDN U1456 ( .A(n1286), .B(n1287), .Z(n1285) );
  XNOR U1457 ( .A(n1284), .B(n1288), .Z(n1287) );
  XNOR U1458 ( .A(n1289), .B(n1290), .Z(n718) );
  NANDN U1459 ( .A(n1291), .B(n1292), .Z(n1290) );
  NANDN U1460 ( .A(n1289), .B(n1293), .Z(n1292) );
  XOR U1461 ( .A(n1294), .B(n719), .Z(n717) );
  IV U1462 ( .A(n715), .Z(n719) );
  XNOR U1463 ( .A(n1295), .B(n1296), .Z(n715) );
  NAND U1464 ( .A(n1297), .B(n1298), .Z(n1296) );
  XOR U1465 ( .A(n1295), .B(n1299), .Z(n1297) );
  NOR U1466 ( .A(n1300), .B(n1301), .Z(n1294) );
  XNOR U1467 ( .A(n755), .B(n728), .Z(n1302) );
  XNOR U1468 ( .A(n1303), .B(n1304), .Z(n728) );
  NANDN U1469 ( .A(n1305), .B(n1306), .Z(n1304) );
  XOR U1470 ( .A(n1303), .B(n1307), .Z(n1306) );
  XNOR U1471 ( .A(n1308), .B(n1309), .Z(n736) );
  NANDN U1472 ( .A(n1310), .B(n1311), .Z(n1309) );
  NANDN U1473 ( .A(n1312), .B(n1308), .Z(n1311) );
  XNOR U1474 ( .A(n1313), .B(n733), .Z(n735) );
  XNOR U1475 ( .A(n1314), .B(n1315), .Z(n733) );
  NAND U1476 ( .A(n1316), .B(n1317), .Z(n1315) );
  XNOR U1477 ( .A(n1314), .B(n1318), .Z(n1316) );
  NOR U1478 ( .A(n1319), .B(n1320), .Z(n1313) );
  XOR U1479 ( .A(n742), .B(n745), .Z(n1321) );
  XNOR U1480 ( .A(n1322), .B(n1323), .Z(n745) );
  NANDN U1481 ( .A(n1324), .B(n1325), .Z(n1323) );
  XOR U1482 ( .A(n1322), .B(n1326), .Z(n1325) );
  XNOR U1483 ( .A(n1327), .B(n1328), .Z(n742) );
  NANDN U1484 ( .A(n1329), .B(n1330), .Z(n1328) );
  NANDN U1485 ( .A(n1327), .B(n1331), .Z(n1330) );
  XOR U1486 ( .A(n1332), .B(n743), .Z(n741) );
  IV U1487 ( .A(n739), .Z(n743) );
  XNOR U1488 ( .A(n1333), .B(n1334), .Z(n739) );
  NAND U1489 ( .A(n1335), .B(n1336), .Z(n1334) );
  XOR U1490 ( .A(n1333), .B(n1337), .Z(n1335) );
  NOR U1491 ( .A(n1338), .B(n1339), .Z(n1332) );
  XNOR U1492 ( .A(n772), .B(n752), .Z(n1340) );
  XNOR U1493 ( .A(n1341), .B(n1342), .Z(n752) );
  NANDN U1494 ( .A(n1343), .B(n1344), .Z(n1342) );
  XOR U1495 ( .A(n1341), .B(n1345), .Z(n1344) );
  XNOR U1496 ( .A(n1346), .B(n1347), .Z(n760) );
  NANDN U1497 ( .A(n1348), .B(n1349), .Z(n1347) );
  NANDN U1498 ( .A(n1350), .B(n1346), .Z(n1349) );
  XNOR U1499 ( .A(n1351), .B(n757), .Z(n759) );
  XNOR U1500 ( .A(n1352), .B(n1353), .Z(n757) );
  NAND U1501 ( .A(n1354), .B(n1355), .Z(n1353) );
  XNOR U1502 ( .A(n1352), .B(n1356), .Z(n1354) );
  NOR U1503 ( .A(n1357), .B(n1358), .Z(n1351) );
  XOR U1504 ( .A(n766), .B(n769), .Z(n1359) );
  XNOR U1505 ( .A(n1360), .B(n1361), .Z(n769) );
  NANDN U1506 ( .A(n1362), .B(n1363), .Z(n1361) );
  XNOR U1507 ( .A(n1360), .B(n1364), .Z(n1363) );
  XNOR U1508 ( .A(n1365), .B(n1366), .Z(n766) );
  NANDN U1509 ( .A(n1367), .B(n1368), .Z(n1366) );
  NANDN U1510 ( .A(n1365), .B(n1369), .Z(n1368) );
  XOR U1511 ( .A(n1370), .B(n767), .Z(n765) );
  IV U1512 ( .A(n763), .Z(n767) );
  XNOR U1513 ( .A(n1371), .B(n1372), .Z(n763) );
  NAND U1514 ( .A(n1373), .B(n1374), .Z(n1372) );
  XOR U1515 ( .A(n1371), .B(n1375), .Z(n1373) );
  NOR U1516 ( .A(n1376), .B(n1377), .Z(n1370) );
  XOR U1517 ( .A(n1378), .B(n1379), .Z(n774) );
  NANDN U1518 ( .A(n26), .B(n1380), .Z(n1379) );
  XNOR U1519 ( .A(n1378), .B(n27), .Z(n1380) );
  XOR U1520 ( .A(n785), .B(n786), .Z(n794) );
  XOR U1521 ( .A(n780), .B(n778), .Z(n786) );
  AND U1522 ( .A(n1381), .B(n776), .Z(n778) );
  OR U1523 ( .A(n1382), .B(n1383), .Z(n776) );
  OR U1524 ( .A(n1384), .B(n1385), .Z(n1381) );
  NOR U1525 ( .A(n1386), .B(n1387), .Z(n780) );
  XOR U1526 ( .A(n787), .B(n1388), .Z(n785) );
  XOR U1527 ( .A(n788), .B(n782), .Z(n1388) );
  NOR U1528 ( .A(n1389), .B(n1390), .Z(n782) );
  OR U1529 ( .A(n1391), .B(n1392), .Z(n788) );
  AND U1530 ( .A(n1393), .B(n1394), .Z(n787) );
  OR U1531 ( .A(n1395), .B(n1396), .Z(n1394) );
  OR U1532 ( .A(n1397), .B(n1398), .Z(n1393) );
  XNOR U1533 ( .A(n804), .B(n1399), .Z(n792) );
  XNOR U1534 ( .A(n790), .B(n805), .Z(n1399) );
  XOR U1535 ( .A(n799), .B(n797), .Z(n805) );
  NOR U1536 ( .A(n1401), .B(n1402), .Z(n795) );
  OR U1537 ( .A(n1403), .B(n1404), .Z(n1400) );
  OR U1538 ( .A(n1405), .B(n1406), .Z(n799) );
  OR U1539 ( .A(n1407), .B(n1408), .Z(n790) );
  XOR U1540 ( .A(n806), .B(n1409), .Z(n804) );
  XOR U1541 ( .A(n807), .B(n801), .Z(n1409) );
  NOR U1542 ( .A(n1410), .B(n1411), .Z(n801) );
  OR U1543 ( .A(n1412), .B(n1413), .Z(n807) );
  AND U1544 ( .A(n1414), .B(n1415), .Z(n806) );
  OR U1545 ( .A(n1416), .B(n1417), .Z(n1415) );
  OR U1546 ( .A(n1418), .B(n1419), .Z(n1414) );
  XOR U1547 ( .A(n809), .B(n832), .Z(n1420) );
  XNOR U1548 ( .A(n823), .B(n824), .Z(n832) );
  XOR U1549 ( .A(n818), .B(n816), .Z(n824) );
  AND U1550 ( .A(n1421), .B(n814), .Z(n816) );
  OR U1551 ( .A(n1422), .B(n1423), .Z(n814) );
  OR U1552 ( .A(n1424), .B(n1425), .Z(n1421) );
  NOR U1553 ( .A(n1426), .B(n1427), .Z(n818) );
  XOR U1554 ( .A(n825), .B(n1428), .Z(n823) );
  XOR U1555 ( .A(n826), .B(n820), .Z(n1428) );
  NOR U1556 ( .A(n1429), .B(n1430), .Z(n820) );
  OR U1557 ( .A(n1431), .B(n1432), .Z(n826) );
  AND U1558 ( .A(n1433), .B(n1434), .Z(n825) );
  OR U1559 ( .A(n1435), .B(n1436), .Z(n1434) );
  OR U1560 ( .A(n1437), .B(n1438), .Z(n1433) );
  OR U1561 ( .A(n1439), .B(n1440), .Z(n809) );
  XNOR U1562 ( .A(n842), .B(n1441), .Z(n830) );
  XNOR U1563 ( .A(n828), .B(n843), .Z(n1441) );
  XOR U1564 ( .A(n837), .B(n835), .Z(n843) );
  NOR U1565 ( .A(n1443), .B(n1444), .Z(n833) );
  OR U1566 ( .A(n1445), .B(n1446), .Z(n1442) );
  OR U1567 ( .A(n1447), .B(n1448), .Z(n837) );
  OR U1568 ( .A(n1449), .B(n1450), .Z(n828) );
  XOR U1569 ( .A(n844), .B(n1451), .Z(n842) );
  XOR U1570 ( .A(n845), .B(n839), .Z(n1451) );
  NOR U1571 ( .A(n1452), .B(n1453), .Z(n839) );
  OR U1572 ( .A(n1454), .B(n1455), .Z(n845) );
  AND U1573 ( .A(n1456), .B(n1457), .Z(n844) );
  OR U1574 ( .A(n1458), .B(n1459), .Z(n1457) );
  OR U1575 ( .A(n1460), .B(n1461), .Z(n1456) );
  XNOR U1576 ( .A(n847), .B(n889), .Z(n1462) );
  XOR U1577 ( .A(n861), .B(n862), .Z(n870) );
  XOR U1578 ( .A(n856), .B(n854), .Z(n862) );
  AND U1579 ( .A(n1463), .B(n852), .Z(n854) );
  OR U1580 ( .A(n1464), .B(n1465), .Z(n852) );
  OR U1581 ( .A(n1466), .B(n1467), .Z(n1463) );
  NOR U1582 ( .A(n1468), .B(n1469), .Z(n856) );
  XOR U1583 ( .A(n863), .B(n1470), .Z(n861) );
  XOR U1584 ( .A(n864), .B(n858), .Z(n1470) );
  NOR U1585 ( .A(n1471), .B(n1472), .Z(n858) );
  OR U1586 ( .A(n1473), .B(n1474), .Z(n864) );
  AND U1587 ( .A(n1475), .B(n1476), .Z(n863) );
  OR U1588 ( .A(n1477), .B(n1478), .Z(n1476) );
  OR U1589 ( .A(n1479), .B(n1480), .Z(n1475) );
  XNOR U1590 ( .A(n880), .B(n1481), .Z(n868) );
  XNOR U1591 ( .A(n866), .B(n881), .Z(n1481) );
  XOR U1592 ( .A(n875), .B(n873), .Z(n881) );
  NOR U1593 ( .A(n1483), .B(n1484), .Z(n871) );
  OR U1594 ( .A(n1485), .B(n1486), .Z(n1482) );
  OR U1595 ( .A(n1487), .B(n1488), .Z(n875) );
  OR U1596 ( .A(n1489), .B(n1490), .Z(n866) );
  XOR U1597 ( .A(n882), .B(n1491), .Z(n880) );
  XOR U1598 ( .A(n883), .B(n877), .Z(n1491) );
  NOR U1599 ( .A(n1492), .B(n1493), .Z(n877) );
  OR U1600 ( .A(n1494), .B(n1495), .Z(n883) );
  AND U1601 ( .A(n1496), .B(n1497), .Z(n882) );
  OR U1602 ( .A(n1498), .B(n1499), .Z(n1497) );
  OR U1603 ( .A(n1500), .B(n1501), .Z(n1496) );
  OR U1604 ( .A(n1502), .B(n1503), .Z(n847) );
  XOR U1605 ( .A(n885), .B(n908), .Z(n1504) );
  XNOR U1606 ( .A(n899), .B(n900), .Z(n908) );
  XOR U1607 ( .A(n894), .B(n892), .Z(n900) );
  AND U1608 ( .A(n1505), .B(n890), .Z(n892) );
  OR U1609 ( .A(n1506), .B(n1507), .Z(n890) );
  OR U1610 ( .A(n1508), .B(n1509), .Z(n1505) );
  NOR U1611 ( .A(n1510), .B(n1511), .Z(n894) );
  XOR U1612 ( .A(n901), .B(n1512), .Z(n899) );
  XOR U1613 ( .A(n902), .B(n896), .Z(n1512) );
  NOR U1614 ( .A(n1513), .B(n1514), .Z(n896) );
  OR U1615 ( .A(n1515), .B(n1516), .Z(n902) );
  AND U1616 ( .A(n1517), .B(n1518), .Z(n901) );
  OR U1617 ( .A(n1519), .B(n1520), .Z(n1518) );
  OR U1618 ( .A(n1521), .B(n1522), .Z(n1517) );
  OR U1619 ( .A(n1523), .B(n1524), .Z(n885) );
  XNOR U1620 ( .A(n918), .B(n1525), .Z(n906) );
  XNOR U1621 ( .A(n904), .B(n919), .Z(n1525) );
  XOR U1622 ( .A(n913), .B(n911), .Z(n919) );
  NOR U1623 ( .A(n1527), .B(n1528), .Z(n909) );
  OR U1624 ( .A(n1529), .B(n1530), .Z(n1526) );
  OR U1625 ( .A(n1531), .B(n1532), .Z(n913) );
  OR U1626 ( .A(n1533), .B(n1534), .Z(n904) );
  XOR U1627 ( .A(n920), .B(n1535), .Z(n918) );
  XOR U1628 ( .A(n921), .B(n915), .Z(n1535) );
  NOR U1629 ( .A(n1536), .B(n1537), .Z(n915) );
  OR U1630 ( .A(n1538), .B(n1539), .Z(n921) );
  AND U1631 ( .A(n1540), .B(n1541), .Z(n920) );
  OR U1632 ( .A(n1542), .B(n1543), .Z(n1541) );
  OR U1633 ( .A(n1544), .B(n1545), .Z(n1540) );
  XNOR U1634 ( .A(n923), .B(n1003), .Z(n1546) );
  XOR U1635 ( .A(n937), .B(n938), .Z(n946) );
  XOR U1636 ( .A(n932), .B(n930), .Z(n938) );
  AND U1637 ( .A(n1547), .B(n928), .Z(n930) );
  OR U1638 ( .A(n1548), .B(n1549), .Z(n928) );
  OR U1639 ( .A(n1550), .B(n1551), .Z(n1547) );
  NOR U1640 ( .A(n1552), .B(n1553), .Z(n932) );
  XOR U1641 ( .A(n939), .B(n1554), .Z(n937) );
  XOR U1642 ( .A(n940), .B(n934), .Z(n1554) );
  NOR U1643 ( .A(n1555), .B(n1556), .Z(n934) );
  OR U1644 ( .A(n1557), .B(n1558), .Z(n940) );
  AND U1645 ( .A(n1559), .B(n1560), .Z(n939) );
  OR U1646 ( .A(n1561), .B(n1562), .Z(n1560) );
  OR U1647 ( .A(n1563), .B(n1564), .Z(n1559) );
  XNOR U1648 ( .A(n956), .B(n1565), .Z(n944) );
  XNOR U1649 ( .A(n942), .B(n957), .Z(n1565) );
  XOR U1650 ( .A(n951), .B(n949), .Z(n957) );
  NOR U1651 ( .A(n1567), .B(n1568), .Z(n947) );
  OR U1652 ( .A(n1569), .B(n1570), .Z(n1566) );
  OR U1653 ( .A(n1571), .B(n1572), .Z(n951) );
  OR U1654 ( .A(n1573), .B(n1574), .Z(n942) );
  XOR U1655 ( .A(n958), .B(n1575), .Z(n956) );
  XOR U1656 ( .A(n959), .B(n953), .Z(n1575) );
  NOR U1657 ( .A(n1576), .B(n1577), .Z(n953) );
  OR U1658 ( .A(n1578), .B(n1579), .Z(n959) );
  AND U1659 ( .A(n1580), .B(n1581), .Z(n958) );
  OR U1660 ( .A(n1582), .B(n1583), .Z(n1581) );
  OR U1661 ( .A(n1584), .B(n1585), .Z(n1580) );
  XOR U1662 ( .A(n961), .B(n984), .Z(n1586) );
  XNOR U1663 ( .A(n975), .B(n976), .Z(n984) );
  XOR U1664 ( .A(n970), .B(n968), .Z(n976) );
  AND U1665 ( .A(n1587), .B(n966), .Z(n968) );
  OR U1666 ( .A(n1588), .B(n1589), .Z(n966) );
  OR U1667 ( .A(n1590), .B(n1591), .Z(n1587) );
  NOR U1668 ( .A(n1592), .B(n1593), .Z(n970) );
  XOR U1669 ( .A(n977), .B(n1594), .Z(n975) );
  XOR U1670 ( .A(n978), .B(n972), .Z(n1594) );
  NOR U1671 ( .A(n1595), .B(n1596), .Z(n972) );
  OR U1672 ( .A(n1597), .B(n1598), .Z(n978) );
  AND U1673 ( .A(n1599), .B(n1600), .Z(n977) );
  OR U1674 ( .A(n1601), .B(n1602), .Z(n1600) );
  OR U1675 ( .A(n1603), .B(n1604), .Z(n1599) );
  OR U1676 ( .A(n1605), .B(n1606), .Z(n961) );
  XNOR U1677 ( .A(n994), .B(n1607), .Z(n982) );
  XNOR U1678 ( .A(n980), .B(n995), .Z(n1607) );
  XOR U1679 ( .A(n989), .B(n987), .Z(n995) );
  NOR U1680 ( .A(n1609), .B(n1610), .Z(n985) );
  OR U1681 ( .A(n1611), .B(n1612), .Z(n1608) );
  OR U1682 ( .A(n1613), .B(n1614), .Z(n989) );
  OR U1683 ( .A(n1615), .B(n1616), .Z(n980) );
  XOR U1684 ( .A(n996), .B(n1617), .Z(n994) );
  XOR U1685 ( .A(n997), .B(n991), .Z(n1617) );
  NOR U1686 ( .A(n1618), .B(n1619), .Z(n991) );
  OR U1687 ( .A(n1620), .B(n1621), .Z(n997) );
  AND U1688 ( .A(n1622), .B(n1623), .Z(n996) );
  OR U1689 ( .A(n1624), .B(n1625), .Z(n1623) );
  OR U1690 ( .A(n1626), .B(n1627), .Z(n1622) );
  OR U1691 ( .A(n1628), .B(n1629), .Z(n923) );
  XNOR U1692 ( .A(n999), .B(n1041), .Z(n1630) );
  XOR U1693 ( .A(n1013), .B(n1014), .Z(n1022) );
  XOR U1694 ( .A(n1008), .B(n1006), .Z(n1014) );
  AND U1695 ( .A(n1631), .B(n1004), .Z(n1006) );
  OR U1696 ( .A(n1632), .B(n1633), .Z(n1004) );
  OR U1697 ( .A(n1634), .B(n1635), .Z(n1631) );
  NOR U1698 ( .A(n1636), .B(n1637), .Z(n1008) );
  XOR U1699 ( .A(n1015), .B(n1638), .Z(n1013) );
  XOR U1700 ( .A(n1016), .B(n1010), .Z(n1638) );
  NOR U1701 ( .A(n1639), .B(n1640), .Z(n1010) );
  OR U1702 ( .A(n1641), .B(n1642), .Z(n1016) );
  AND U1703 ( .A(n1643), .B(n1644), .Z(n1015) );
  OR U1704 ( .A(n1645), .B(n1646), .Z(n1644) );
  OR U1705 ( .A(n1647), .B(n1648), .Z(n1643) );
  XNOR U1706 ( .A(n1032), .B(n1649), .Z(n1020) );
  XNOR U1707 ( .A(n1018), .B(n1033), .Z(n1649) );
  XOR U1708 ( .A(n1027), .B(n1025), .Z(n1033) );
  NOR U1709 ( .A(n1651), .B(n1652), .Z(n1023) );
  OR U1710 ( .A(n1653), .B(n1654), .Z(n1650) );
  OR U1711 ( .A(n1655), .B(n1656), .Z(n1027) );
  OR U1712 ( .A(n1657), .B(n1658), .Z(n1018) );
  XOR U1713 ( .A(n1034), .B(n1659), .Z(n1032) );
  XOR U1714 ( .A(n1035), .B(n1029), .Z(n1659) );
  NOR U1715 ( .A(n1660), .B(n1661), .Z(n1029) );
  OR U1716 ( .A(n1662), .B(n1663), .Z(n1035) );
  AND U1717 ( .A(n1664), .B(n1665), .Z(n1034) );
  OR U1718 ( .A(n1666), .B(n1667), .Z(n1665) );
  OR U1719 ( .A(n1668), .B(n1669), .Z(n1664) );
  OR U1720 ( .A(n1670), .B(n1671), .Z(n999) );
  XOR U1721 ( .A(n1037), .B(n1060), .Z(n1672) );
  XNOR U1722 ( .A(n1051), .B(n1052), .Z(n1060) );
  XOR U1723 ( .A(n1046), .B(n1044), .Z(n1052) );
  AND U1724 ( .A(n1673), .B(n1042), .Z(n1044) );
  OR U1725 ( .A(n1674), .B(n1675), .Z(n1042) );
  OR U1726 ( .A(n1676), .B(n1677), .Z(n1673) );
  NOR U1727 ( .A(n1678), .B(n1679), .Z(n1046) );
  XOR U1728 ( .A(n1053), .B(n1680), .Z(n1051) );
  XOR U1729 ( .A(n1054), .B(n1048), .Z(n1680) );
  NOR U1730 ( .A(n1681), .B(n1682), .Z(n1048) );
  OR U1731 ( .A(n1683), .B(n1684), .Z(n1054) );
  AND U1732 ( .A(n1685), .B(n1686), .Z(n1053) );
  OR U1733 ( .A(n1687), .B(n1688), .Z(n1686) );
  OR U1734 ( .A(n1689), .B(n1690), .Z(n1685) );
  OR U1735 ( .A(n1691), .B(n1692), .Z(n1037) );
  XNOR U1736 ( .A(n1070), .B(n1693), .Z(n1058) );
  XNOR U1737 ( .A(n1056), .B(n1071), .Z(n1693) );
  XOR U1738 ( .A(n1065), .B(n1063), .Z(n1071) );
  NOR U1739 ( .A(n1695), .B(n1696), .Z(n1061) );
  OR U1740 ( .A(n1697), .B(n1698), .Z(n1694) );
  OR U1741 ( .A(n1699), .B(n1700), .Z(n1065) );
  OR U1742 ( .A(n1701), .B(n1702), .Z(n1056) );
  XOR U1743 ( .A(n1072), .B(n1703), .Z(n1070) );
  XOR U1744 ( .A(n1073), .B(n1067), .Z(n1703) );
  NOR U1745 ( .A(n1704), .B(n1705), .Z(n1067) );
  OR U1746 ( .A(n1706), .B(n1707), .Z(n1073) );
  AND U1747 ( .A(n1708), .B(n1709), .Z(n1072) );
  OR U1748 ( .A(n1710), .B(n1711), .Z(n1709) );
  OR U1749 ( .A(n1712), .B(n1713), .Z(n1708) );
  XNOR U1750 ( .A(n1075), .B(n1231), .Z(n1714) );
  XOR U1751 ( .A(n1089), .B(n1090), .Z(n1098) );
  XOR U1752 ( .A(n1084), .B(n1082), .Z(n1090) );
  AND U1753 ( .A(n1715), .B(n1080), .Z(n1082) );
  OR U1754 ( .A(n1716), .B(n1717), .Z(n1080) );
  OR U1755 ( .A(n1718), .B(n1719), .Z(n1715) );
  NOR U1756 ( .A(n1720), .B(n1721), .Z(n1084) );
  XOR U1757 ( .A(n1091), .B(n1722), .Z(n1089) );
  XOR U1758 ( .A(n1092), .B(n1086), .Z(n1722) );
  NOR U1759 ( .A(n1723), .B(n1724), .Z(n1086) );
  OR U1760 ( .A(n1725), .B(n1726), .Z(n1092) );
  AND U1761 ( .A(n1727), .B(n1728), .Z(n1091) );
  OR U1762 ( .A(n1729), .B(n1730), .Z(n1728) );
  OR U1763 ( .A(n1731), .B(n1732), .Z(n1727) );
  XNOR U1764 ( .A(n1108), .B(n1733), .Z(n1096) );
  XNOR U1765 ( .A(n1094), .B(n1109), .Z(n1733) );
  XOR U1766 ( .A(n1103), .B(n1101), .Z(n1109) );
  NOR U1767 ( .A(n1735), .B(n1736), .Z(n1099) );
  OR U1768 ( .A(n1737), .B(n1738), .Z(n1734) );
  OR U1769 ( .A(n1739), .B(n1740), .Z(n1103) );
  OR U1770 ( .A(n1741), .B(n1742), .Z(n1094) );
  XOR U1771 ( .A(n1110), .B(n1743), .Z(n1108) );
  XOR U1772 ( .A(n1111), .B(n1105), .Z(n1743) );
  NOR U1773 ( .A(n1744), .B(n1745), .Z(n1105) );
  OR U1774 ( .A(n1746), .B(n1747), .Z(n1111) );
  AND U1775 ( .A(n1748), .B(n1749), .Z(n1110) );
  OR U1776 ( .A(n1750), .B(n1751), .Z(n1749) );
  OR U1777 ( .A(n1752), .B(n1753), .Z(n1748) );
  XOR U1778 ( .A(n1113), .B(n1136), .Z(n1754) );
  XNOR U1779 ( .A(n1127), .B(n1128), .Z(n1136) );
  XOR U1780 ( .A(n1122), .B(n1120), .Z(n1128) );
  AND U1781 ( .A(n1755), .B(n1118), .Z(n1120) );
  OR U1782 ( .A(n1756), .B(n1757), .Z(n1118) );
  OR U1783 ( .A(n1758), .B(n1759), .Z(n1755) );
  NOR U1784 ( .A(n1760), .B(n1761), .Z(n1122) );
  XOR U1785 ( .A(n1129), .B(n1762), .Z(n1127) );
  XOR U1786 ( .A(n1130), .B(n1124), .Z(n1762) );
  NOR U1787 ( .A(n1763), .B(n1764), .Z(n1124) );
  OR U1788 ( .A(n1765), .B(n1766), .Z(n1130) );
  AND U1789 ( .A(n1767), .B(n1768), .Z(n1129) );
  OR U1790 ( .A(n1769), .B(n1770), .Z(n1768) );
  OR U1791 ( .A(n1771), .B(n1772), .Z(n1767) );
  OR U1792 ( .A(n1773), .B(n1774), .Z(n1113) );
  XNOR U1793 ( .A(n1146), .B(n1775), .Z(n1134) );
  XNOR U1794 ( .A(n1132), .B(n1147), .Z(n1775) );
  XOR U1795 ( .A(n1141), .B(n1139), .Z(n1147) );
  NOR U1796 ( .A(n1777), .B(n1778), .Z(n1137) );
  OR U1797 ( .A(n1779), .B(n1780), .Z(n1776) );
  OR U1798 ( .A(n1781), .B(n1782), .Z(n1141) );
  OR U1799 ( .A(n1783), .B(n1784), .Z(n1132) );
  XOR U1800 ( .A(n1148), .B(n1785), .Z(n1146) );
  XOR U1801 ( .A(n1149), .B(n1143), .Z(n1785) );
  NOR U1802 ( .A(n1786), .B(n1787), .Z(n1143) );
  OR U1803 ( .A(n1788), .B(n1789), .Z(n1149) );
  AND U1804 ( .A(n1790), .B(n1791), .Z(n1148) );
  OR U1805 ( .A(n1792), .B(n1793), .Z(n1791) );
  OR U1806 ( .A(n1794), .B(n1795), .Z(n1790) );
  XNOR U1807 ( .A(n1151), .B(n1193), .Z(n1796) );
  XOR U1808 ( .A(n1165), .B(n1166), .Z(n1174) );
  XOR U1809 ( .A(n1160), .B(n1158), .Z(n1166) );
  AND U1810 ( .A(n1797), .B(n1156), .Z(n1158) );
  OR U1811 ( .A(n1798), .B(n1799), .Z(n1156) );
  OR U1812 ( .A(n1800), .B(n1801), .Z(n1797) );
  NOR U1813 ( .A(n1802), .B(n1803), .Z(n1160) );
  XOR U1814 ( .A(n1167), .B(n1804), .Z(n1165) );
  XOR U1815 ( .A(n1168), .B(n1162), .Z(n1804) );
  NOR U1816 ( .A(n1805), .B(n1806), .Z(n1162) );
  OR U1817 ( .A(n1807), .B(n1808), .Z(n1168) );
  AND U1818 ( .A(n1809), .B(n1810), .Z(n1167) );
  OR U1819 ( .A(n1811), .B(n1812), .Z(n1810) );
  OR U1820 ( .A(n1813), .B(n1814), .Z(n1809) );
  XNOR U1821 ( .A(n1184), .B(n1815), .Z(n1172) );
  XNOR U1822 ( .A(n1170), .B(n1185), .Z(n1815) );
  XOR U1823 ( .A(n1179), .B(n1177), .Z(n1185) );
  NOR U1824 ( .A(n1817), .B(n1818), .Z(n1175) );
  OR U1825 ( .A(n1819), .B(n1820), .Z(n1816) );
  OR U1826 ( .A(n1821), .B(n1822), .Z(n1179) );
  OR U1827 ( .A(n1823), .B(n1824), .Z(n1170) );
  XOR U1828 ( .A(n1186), .B(n1825), .Z(n1184) );
  XOR U1829 ( .A(n1187), .B(n1181), .Z(n1825) );
  NOR U1830 ( .A(n1826), .B(n1827), .Z(n1181) );
  OR U1831 ( .A(n1828), .B(n1829), .Z(n1187) );
  AND U1832 ( .A(n1830), .B(n1831), .Z(n1186) );
  OR U1833 ( .A(n1832), .B(n1833), .Z(n1831) );
  OR U1834 ( .A(n1834), .B(n1835), .Z(n1830) );
  OR U1835 ( .A(n1836), .B(n1837), .Z(n1151) );
  XOR U1836 ( .A(n1189), .B(n1212), .Z(n1838) );
  XNOR U1837 ( .A(n1203), .B(n1204), .Z(n1212) );
  XOR U1838 ( .A(n1198), .B(n1196), .Z(n1204) );
  AND U1839 ( .A(n1839), .B(n1194), .Z(n1196) );
  OR U1840 ( .A(n1840), .B(n1841), .Z(n1194) );
  OR U1841 ( .A(n1842), .B(n1843), .Z(n1839) );
  NOR U1842 ( .A(n1844), .B(n1845), .Z(n1198) );
  XOR U1843 ( .A(n1205), .B(n1846), .Z(n1203) );
  XOR U1844 ( .A(n1206), .B(n1200), .Z(n1846) );
  NOR U1845 ( .A(n1847), .B(n1848), .Z(n1200) );
  OR U1846 ( .A(n1849), .B(n1850), .Z(n1206) );
  AND U1847 ( .A(n1851), .B(n1852), .Z(n1205) );
  OR U1848 ( .A(n1853), .B(n1854), .Z(n1852) );
  OR U1849 ( .A(n1855), .B(n1856), .Z(n1851) );
  OR U1850 ( .A(n1857), .B(n1858), .Z(n1189) );
  XNOR U1851 ( .A(n1222), .B(n1859), .Z(n1210) );
  XNOR U1852 ( .A(n1208), .B(n1223), .Z(n1859) );
  XOR U1853 ( .A(n1217), .B(n1215), .Z(n1223) );
  NOR U1854 ( .A(n1861), .B(n1862), .Z(n1213) );
  OR U1855 ( .A(n1863), .B(n1864), .Z(n1860) );
  OR U1856 ( .A(n1865), .B(n1866), .Z(n1217) );
  OR U1857 ( .A(n1867), .B(n1868), .Z(n1208) );
  XOR U1858 ( .A(n1224), .B(n1869), .Z(n1222) );
  XOR U1859 ( .A(n1225), .B(n1219), .Z(n1869) );
  NOR U1860 ( .A(n1870), .B(n1871), .Z(n1219) );
  OR U1861 ( .A(n1872), .B(n1873), .Z(n1225) );
  AND U1862 ( .A(n1874), .B(n1875), .Z(n1224) );
  OR U1863 ( .A(n1876), .B(n1877), .Z(n1875) );
  OR U1864 ( .A(n1878), .B(n1879), .Z(n1874) );
  OR U1865 ( .A(n1880), .B(n1881), .Z(n1075) );
  XNOR U1866 ( .A(n1227), .B(n1307), .Z(n1882) );
  XOR U1867 ( .A(n1241), .B(n1242), .Z(n1250) );
  XOR U1868 ( .A(n1236), .B(n1234), .Z(n1242) );
  AND U1869 ( .A(n1883), .B(n1232), .Z(n1234) );
  OR U1870 ( .A(n1884), .B(n1885), .Z(n1232) );
  OR U1871 ( .A(n1886), .B(n1887), .Z(n1883) );
  NOR U1872 ( .A(n1888), .B(n1889), .Z(n1236) );
  XOR U1873 ( .A(n1243), .B(n1890), .Z(n1241) );
  XOR U1874 ( .A(n1244), .B(n1238), .Z(n1890) );
  NOR U1875 ( .A(n1891), .B(n1892), .Z(n1238) );
  OR U1876 ( .A(n1893), .B(n1894), .Z(n1244) );
  AND U1877 ( .A(n1895), .B(n1896), .Z(n1243) );
  OR U1878 ( .A(n1897), .B(n1898), .Z(n1896) );
  OR U1879 ( .A(n1899), .B(n1900), .Z(n1895) );
  XNOR U1880 ( .A(n1260), .B(n1901), .Z(n1248) );
  XNOR U1881 ( .A(n1246), .B(n1261), .Z(n1901) );
  XOR U1882 ( .A(n1255), .B(n1253), .Z(n1261) );
  NOR U1883 ( .A(n1903), .B(n1904), .Z(n1251) );
  OR U1884 ( .A(n1905), .B(n1906), .Z(n1902) );
  OR U1885 ( .A(n1907), .B(n1908), .Z(n1255) );
  OR U1886 ( .A(n1909), .B(n1910), .Z(n1246) );
  XOR U1887 ( .A(n1262), .B(n1911), .Z(n1260) );
  XOR U1888 ( .A(n1263), .B(n1257), .Z(n1911) );
  NOR U1889 ( .A(n1912), .B(n1913), .Z(n1257) );
  OR U1890 ( .A(n1914), .B(n1915), .Z(n1263) );
  AND U1891 ( .A(n1916), .B(n1917), .Z(n1262) );
  OR U1892 ( .A(n1918), .B(n1919), .Z(n1917) );
  OR U1893 ( .A(n1920), .B(n1921), .Z(n1916) );
  XOR U1894 ( .A(n1265), .B(n1288), .Z(n1922) );
  XNOR U1895 ( .A(n1279), .B(n1280), .Z(n1288) );
  XOR U1896 ( .A(n1274), .B(n1272), .Z(n1280) );
  AND U1897 ( .A(n1923), .B(n1270), .Z(n1272) );
  OR U1898 ( .A(n1924), .B(n1925), .Z(n1270) );
  OR U1899 ( .A(n1926), .B(n1927), .Z(n1923) );
  NOR U1900 ( .A(n1928), .B(n1929), .Z(n1274) );
  XOR U1901 ( .A(n1281), .B(n1930), .Z(n1279) );
  XOR U1902 ( .A(n1282), .B(n1276), .Z(n1930) );
  NOR U1903 ( .A(n1931), .B(n1932), .Z(n1276) );
  OR U1904 ( .A(n1933), .B(n1934), .Z(n1282) );
  AND U1905 ( .A(n1935), .B(n1936), .Z(n1281) );
  OR U1906 ( .A(n1937), .B(n1938), .Z(n1936) );
  OR U1907 ( .A(n1939), .B(n1940), .Z(n1935) );
  OR U1908 ( .A(n1941), .B(n1942), .Z(n1265) );
  XNOR U1909 ( .A(n1298), .B(n1943), .Z(n1286) );
  XNOR U1910 ( .A(n1284), .B(n1299), .Z(n1943) );
  XOR U1911 ( .A(n1293), .B(n1291), .Z(n1299) );
  NOR U1912 ( .A(n1945), .B(n1946), .Z(n1289) );
  OR U1913 ( .A(n1947), .B(n1948), .Z(n1944) );
  OR U1914 ( .A(n1949), .B(n1950), .Z(n1293) );
  OR U1915 ( .A(n1951), .B(n1952), .Z(n1284) );
  XOR U1916 ( .A(n1300), .B(n1953), .Z(n1298) );
  XOR U1917 ( .A(n1301), .B(n1295), .Z(n1953) );
  NOR U1918 ( .A(n1954), .B(n1955), .Z(n1295) );
  OR U1919 ( .A(n1956), .B(n1957), .Z(n1301) );
  AND U1920 ( .A(n1958), .B(n1959), .Z(n1300) );
  OR U1921 ( .A(n1960), .B(n1961), .Z(n1959) );
  OR U1922 ( .A(n1962), .B(n1963), .Z(n1958) );
  OR U1923 ( .A(n1964), .B(n1965), .Z(n1227) );
  XNOR U1924 ( .A(n1303), .B(n1345), .Z(n1966) );
  XOR U1925 ( .A(n1317), .B(n1318), .Z(n1326) );
  XOR U1926 ( .A(n1312), .B(n1310), .Z(n1318) );
  AND U1927 ( .A(n1967), .B(n1308), .Z(n1310) );
  OR U1928 ( .A(n1968), .B(n1969), .Z(n1308) );
  OR U1929 ( .A(n1970), .B(n1971), .Z(n1967) );
  NOR U1930 ( .A(n1972), .B(n1973), .Z(n1312) );
  XOR U1931 ( .A(n1319), .B(n1974), .Z(n1317) );
  XOR U1932 ( .A(n1320), .B(n1314), .Z(n1974) );
  NOR U1933 ( .A(n1975), .B(n1976), .Z(n1314) );
  OR U1934 ( .A(n1977), .B(n1978), .Z(n1320) );
  AND U1935 ( .A(n1979), .B(n1980), .Z(n1319) );
  OR U1936 ( .A(n1981), .B(n1982), .Z(n1980) );
  OR U1937 ( .A(n1983), .B(n1984), .Z(n1979) );
  XNOR U1938 ( .A(n1336), .B(n1985), .Z(n1324) );
  XNOR U1939 ( .A(n1322), .B(n1337), .Z(n1985) );
  XOR U1940 ( .A(n1331), .B(n1329), .Z(n1337) );
  NOR U1941 ( .A(n1987), .B(n1988), .Z(n1327) );
  OR U1942 ( .A(n1989), .B(n1990), .Z(n1986) );
  OR U1943 ( .A(n1991), .B(n1992), .Z(n1331) );
  OR U1944 ( .A(n1993), .B(n1994), .Z(n1322) );
  XOR U1945 ( .A(n1338), .B(n1995), .Z(n1336) );
  XOR U1946 ( .A(n1339), .B(n1333), .Z(n1995) );
  NOR U1947 ( .A(n1996), .B(n1997), .Z(n1333) );
  OR U1948 ( .A(n1998), .B(n1999), .Z(n1339) );
  AND U1949 ( .A(n2000), .B(n2001), .Z(n1338) );
  OR U1950 ( .A(n2002), .B(n2003), .Z(n2001) );
  OR U1951 ( .A(n2004), .B(n2005), .Z(n2000) );
  OR U1952 ( .A(n2006), .B(n2007), .Z(n1303) );
  XOR U1953 ( .A(n1341), .B(n1364), .Z(n2008) );
  XNOR U1954 ( .A(n1355), .B(n1356), .Z(n1364) );
  XOR U1955 ( .A(n1350), .B(n1348), .Z(n1356) );
  AND U1956 ( .A(n2009), .B(n1346), .Z(n1348) );
  OR U1957 ( .A(n2010), .B(n2011), .Z(n1346) );
  OR U1958 ( .A(n2012), .B(n2013), .Z(n2009) );
  NOR U1959 ( .A(n2014), .B(n2015), .Z(n1350) );
  XOR U1960 ( .A(n1357), .B(n2016), .Z(n1355) );
  XOR U1961 ( .A(n1358), .B(n1352), .Z(n2016) );
  NOR U1962 ( .A(n2017), .B(n2018), .Z(n1352) );
  OR U1963 ( .A(n2019), .B(n2020), .Z(n1358) );
  AND U1964 ( .A(n2021), .B(n2022), .Z(n1357) );
  OR U1965 ( .A(n2023), .B(n2024), .Z(n2022) );
  OR U1966 ( .A(n2025), .B(n2026), .Z(n2021) );
  OR U1967 ( .A(n2027), .B(n2028), .Z(n1341) );
  XNOR U1968 ( .A(n1374), .B(n2029), .Z(n1362) );
  XNOR U1969 ( .A(n1360), .B(n1375), .Z(n2029) );
  XOR U1970 ( .A(n1369), .B(n1367), .Z(n1375) );
  NOR U1971 ( .A(n2031), .B(n2032), .Z(n1365) );
  OR U1972 ( .A(n2033), .B(n2034), .Z(n2030) );
  OR U1973 ( .A(n2035), .B(n2036), .Z(n1369) );
  OR U1974 ( .A(n2037), .B(n2038), .Z(n1360) );
  XOR U1975 ( .A(n1376), .B(n2039), .Z(n1374) );
  XOR U1976 ( .A(n1377), .B(n1371), .Z(n2039) );
  NOR U1977 ( .A(n2040), .B(n2041), .Z(n1371) );
  OR U1978 ( .A(n2042), .B(n2043), .Z(n1377) );
  AND U1979 ( .A(n2044), .B(n2045), .Z(n1376) );
  OR U1980 ( .A(n2046), .B(n2047), .Z(n2045) );
  OR U1981 ( .A(n2048), .B(n2049), .Z(n2044) );
  XNOR U1982 ( .A(oglobal[1]), .B(n1378), .Z(n26) );
  ANDN U1983 ( .B(oglobal[0]), .A(n2050), .Z(n1378) );
  XNOR U1984 ( .A(oglobal[0]), .B(n2050), .Z(o[0]) );
  XNOR U1985 ( .A(n1881), .B(n1880), .Z(n2050) );
  XNOR U1986 ( .A(n1629), .B(n1628), .Z(n1880) );
  XNOR U1987 ( .A(n1503), .B(n1502), .Z(n1628) );
  XNOR U1988 ( .A(n1440), .B(n1439), .Z(n1502) );
  XNOR U1989 ( .A(n1408), .B(n1407), .Z(n1439) );
  XNOR U1990 ( .A(n1382), .B(n1383), .Z(n1389) );
  XNOR U1991 ( .A(n1386), .B(n1387), .Z(n1383) );
  XNOR U1992 ( .A(y[255]), .B(x[255]), .Z(n1387) );
  XNOR U1993 ( .A(y[254]), .B(x[254]), .Z(n1386) );
  XNOR U1994 ( .A(n1384), .B(n1385), .Z(n1382) );
  XNOR U1995 ( .A(y[253]), .B(x[253]), .Z(n1385) );
  XNOR U1996 ( .A(y[252]), .B(x[252]), .Z(n1384) );
  XNOR U1997 ( .A(n1397), .B(n1398), .Z(n1390) );
  XNOR U1998 ( .A(n1392), .B(n1391), .Z(n1398) );
  XNOR U1999 ( .A(y[251]), .B(x[251]), .Z(n1391) );
  XNOR U2000 ( .A(y[250]), .B(x[250]), .Z(n1392) );
  XNOR U2001 ( .A(n1395), .B(n1396), .Z(n1397) );
  XNOR U2002 ( .A(y[249]), .B(x[249]), .Z(n1396) );
  XNOR U2003 ( .A(y[248]), .B(x[248]), .Z(n1395) );
  XNOR U2004 ( .A(n1401), .B(n1402), .Z(n1410) );
  XNOR U2005 ( .A(n1405), .B(n1406), .Z(n1402) );
  XNOR U2006 ( .A(y[247]), .B(x[247]), .Z(n1406) );
  XNOR U2007 ( .A(y[246]), .B(x[246]), .Z(n1405) );
  XNOR U2008 ( .A(n1403), .B(n1404), .Z(n1401) );
  XNOR U2009 ( .A(y[245]), .B(x[245]), .Z(n1404) );
  XNOR U2010 ( .A(y[244]), .B(x[244]), .Z(n1403) );
  XNOR U2011 ( .A(n1418), .B(n1419), .Z(n1411) );
  XNOR U2012 ( .A(n1413), .B(n1412), .Z(n1419) );
  XNOR U2013 ( .A(y[243]), .B(x[243]), .Z(n1412) );
  XNOR U2014 ( .A(y[242]), .B(x[242]), .Z(n1413) );
  XNOR U2015 ( .A(n1416), .B(n1417), .Z(n1418) );
  XNOR U2016 ( .A(y[241]), .B(x[241]), .Z(n1417) );
  XNOR U2017 ( .A(y[240]), .B(x[240]), .Z(n1416) );
  XNOR U2018 ( .A(n1450), .B(n1449), .Z(n1440) );
  XNOR U2019 ( .A(n1422), .B(n1423), .Z(n1429) );
  XNOR U2020 ( .A(n1426), .B(n1427), .Z(n1423) );
  XNOR U2021 ( .A(y[239]), .B(x[239]), .Z(n1427) );
  XNOR U2022 ( .A(y[238]), .B(x[238]), .Z(n1426) );
  XNOR U2023 ( .A(n1424), .B(n1425), .Z(n1422) );
  XNOR U2024 ( .A(y[237]), .B(x[237]), .Z(n1425) );
  XNOR U2025 ( .A(y[236]), .B(x[236]), .Z(n1424) );
  XNOR U2026 ( .A(n1437), .B(n1438), .Z(n1430) );
  XNOR U2027 ( .A(n1432), .B(n1431), .Z(n1438) );
  XNOR U2028 ( .A(y[235]), .B(x[235]), .Z(n1431) );
  XNOR U2029 ( .A(y[234]), .B(x[234]), .Z(n1432) );
  XNOR U2030 ( .A(n1435), .B(n1436), .Z(n1437) );
  XNOR U2031 ( .A(y[233]), .B(x[233]), .Z(n1436) );
  XNOR U2032 ( .A(y[232]), .B(x[232]), .Z(n1435) );
  XNOR U2033 ( .A(n1443), .B(n1444), .Z(n1452) );
  XNOR U2034 ( .A(n1447), .B(n1448), .Z(n1444) );
  XNOR U2035 ( .A(y[231]), .B(x[231]), .Z(n1448) );
  XNOR U2036 ( .A(y[230]), .B(x[230]), .Z(n1447) );
  XNOR U2037 ( .A(n1445), .B(n1446), .Z(n1443) );
  XNOR U2038 ( .A(y[229]), .B(x[229]), .Z(n1446) );
  XNOR U2039 ( .A(y[228]), .B(x[228]), .Z(n1445) );
  XNOR U2040 ( .A(n1460), .B(n1461), .Z(n1453) );
  XNOR U2041 ( .A(n1455), .B(n1454), .Z(n1461) );
  XNOR U2042 ( .A(y[227]), .B(x[227]), .Z(n1454) );
  XNOR U2043 ( .A(y[226]), .B(x[226]), .Z(n1455) );
  XNOR U2044 ( .A(n1458), .B(n1459), .Z(n1460) );
  XNOR U2045 ( .A(y[225]), .B(x[225]), .Z(n1459) );
  XNOR U2046 ( .A(y[224]), .B(x[224]), .Z(n1458) );
  XNOR U2047 ( .A(n1524), .B(n1523), .Z(n1503) );
  XNOR U2048 ( .A(n1490), .B(n1489), .Z(n1523) );
  XNOR U2049 ( .A(n1464), .B(n1465), .Z(n1471) );
  XNOR U2050 ( .A(n1468), .B(n1469), .Z(n1465) );
  XNOR U2051 ( .A(y[223]), .B(x[223]), .Z(n1469) );
  XNOR U2052 ( .A(y[222]), .B(x[222]), .Z(n1468) );
  XNOR U2053 ( .A(n1466), .B(n1467), .Z(n1464) );
  XNOR U2054 ( .A(y[221]), .B(x[221]), .Z(n1467) );
  XNOR U2055 ( .A(y[220]), .B(x[220]), .Z(n1466) );
  XNOR U2056 ( .A(n1479), .B(n1480), .Z(n1472) );
  XNOR U2057 ( .A(n1474), .B(n1473), .Z(n1480) );
  XNOR U2058 ( .A(y[219]), .B(x[219]), .Z(n1473) );
  XNOR U2059 ( .A(y[218]), .B(x[218]), .Z(n1474) );
  XNOR U2060 ( .A(n1477), .B(n1478), .Z(n1479) );
  XNOR U2061 ( .A(y[217]), .B(x[217]), .Z(n1478) );
  XNOR U2062 ( .A(y[216]), .B(x[216]), .Z(n1477) );
  XNOR U2063 ( .A(n1483), .B(n1484), .Z(n1492) );
  XNOR U2064 ( .A(n1487), .B(n1488), .Z(n1484) );
  XNOR U2065 ( .A(y[215]), .B(x[215]), .Z(n1488) );
  XNOR U2066 ( .A(y[214]), .B(x[214]), .Z(n1487) );
  XNOR U2067 ( .A(n1485), .B(n1486), .Z(n1483) );
  XNOR U2068 ( .A(y[213]), .B(x[213]), .Z(n1486) );
  XNOR U2069 ( .A(y[212]), .B(x[212]), .Z(n1485) );
  XNOR U2070 ( .A(n1500), .B(n1501), .Z(n1493) );
  XNOR U2071 ( .A(n1495), .B(n1494), .Z(n1501) );
  XNOR U2072 ( .A(y[211]), .B(x[211]), .Z(n1494) );
  XNOR U2073 ( .A(y[210]), .B(x[210]), .Z(n1495) );
  XNOR U2074 ( .A(n1498), .B(n1499), .Z(n1500) );
  XNOR U2075 ( .A(y[209]), .B(x[209]), .Z(n1499) );
  XNOR U2076 ( .A(y[208]), .B(x[208]), .Z(n1498) );
  XNOR U2077 ( .A(n1534), .B(n1533), .Z(n1524) );
  XNOR U2078 ( .A(n1506), .B(n1507), .Z(n1513) );
  XNOR U2079 ( .A(n1510), .B(n1511), .Z(n1507) );
  XNOR U2080 ( .A(y[207]), .B(x[207]), .Z(n1511) );
  XNOR U2081 ( .A(y[206]), .B(x[206]), .Z(n1510) );
  XNOR U2082 ( .A(n1508), .B(n1509), .Z(n1506) );
  XNOR U2083 ( .A(y[205]), .B(x[205]), .Z(n1509) );
  XNOR U2084 ( .A(y[204]), .B(x[204]), .Z(n1508) );
  XNOR U2085 ( .A(n1521), .B(n1522), .Z(n1514) );
  XNOR U2086 ( .A(n1516), .B(n1515), .Z(n1522) );
  XNOR U2087 ( .A(y[203]), .B(x[203]), .Z(n1515) );
  XNOR U2088 ( .A(y[202]), .B(x[202]), .Z(n1516) );
  XNOR U2089 ( .A(n1519), .B(n1520), .Z(n1521) );
  XNOR U2090 ( .A(y[201]), .B(x[201]), .Z(n1520) );
  XNOR U2091 ( .A(y[200]), .B(x[200]), .Z(n1519) );
  XNOR U2092 ( .A(n1527), .B(n1528), .Z(n1536) );
  XNOR U2093 ( .A(n1531), .B(n1532), .Z(n1528) );
  XNOR U2094 ( .A(y[199]), .B(x[199]), .Z(n1532) );
  XNOR U2095 ( .A(y[198]), .B(x[198]), .Z(n1531) );
  XNOR U2096 ( .A(n1529), .B(n1530), .Z(n1527) );
  XNOR U2097 ( .A(y[197]), .B(x[197]), .Z(n1530) );
  XNOR U2098 ( .A(y[196]), .B(x[196]), .Z(n1529) );
  XNOR U2099 ( .A(n1544), .B(n1545), .Z(n1537) );
  XNOR U2100 ( .A(n1539), .B(n1538), .Z(n1545) );
  XNOR U2101 ( .A(y[195]), .B(x[195]), .Z(n1538) );
  XNOR U2102 ( .A(y[194]), .B(x[194]), .Z(n1539) );
  XNOR U2103 ( .A(n1542), .B(n1543), .Z(n1544) );
  XNOR U2104 ( .A(y[193]), .B(x[193]), .Z(n1543) );
  XNOR U2105 ( .A(y[192]), .B(x[192]), .Z(n1542) );
  XNOR U2106 ( .A(n1671), .B(n1670), .Z(n1629) );
  XNOR U2107 ( .A(n1606), .B(n1605), .Z(n1670) );
  XNOR U2108 ( .A(n1574), .B(n1573), .Z(n1605) );
  XNOR U2109 ( .A(n1548), .B(n1549), .Z(n1555) );
  XNOR U2110 ( .A(n1552), .B(n1553), .Z(n1549) );
  XNOR U2111 ( .A(y[191]), .B(x[191]), .Z(n1553) );
  XNOR U2112 ( .A(y[190]), .B(x[190]), .Z(n1552) );
  XNOR U2113 ( .A(n1550), .B(n1551), .Z(n1548) );
  XNOR U2114 ( .A(y[189]), .B(x[189]), .Z(n1551) );
  XNOR U2115 ( .A(y[188]), .B(x[188]), .Z(n1550) );
  XNOR U2116 ( .A(n1563), .B(n1564), .Z(n1556) );
  XNOR U2117 ( .A(n1558), .B(n1557), .Z(n1564) );
  XNOR U2118 ( .A(y[187]), .B(x[187]), .Z(n1557) );
  XNOR U2119 ( .A(y[186]), .B(x[186]), .Z(n1558) );
  XNOR U2120 ( .A(n1561), .B(n1562), .Z(n1563) );
  XNOR U2121 ( .A(y[185]), .B(x[185]), .Z(n1562) );
  XNOR U2122 ( .A(y[184]), .B(x[184]), .Z(n1561) );
  XNOR U2123 ( .A(n1567), .B(n1568), .Z(n1576) );
  XNOR U2124 ( .A(n1571), .B(n1572), .Z(n1568) );
  XNOR U2125 ( .A(y[183]), .B(x[183]), .Z(n1572) );
  XNOR U2126 ( .A(y[182]), .B(x[182]), .Z(n1571) );
  XNOR U2127 ( .A(n1569), .B(n1570), .Z(n1567) );
  XNOR U2128 ( .A(y[181]), .B(x[181]), .Z(n1570) );
  XNOR U2129 ( .A(y[180]), .B(x[180]), .Z(n1569) );
  XNOR U2130 ( .A(n1584), .B(n1585), .Z(n1577) );
  XNOR U2131 ( .A(n1579), .B(n1578), .Z(n1585) );
  XNOR U2132 ( .A(y[179]), .B(x[179]), .Z(n1578) );
  XNOR U2133 ( .A(y[178]), .B(x[178]), .Z(n1579) );
  XNOR U2134 ( .A(n1582), .B(n1583), .Z(n1584) );
  XNOR U2135 ( .A(y[177]), .B(x[177]), .Z(n1583) );
  XNOR U2136 ( .A(y[176]), .B(x[176]), .Z(n1582) );
  XNOR U2137 ( .A(n1616), .B(n1615), .Z(n1606) );
  XNOR U2138 ( .A(n1588), .B(n1589), .Z(n1595) );
  XNOR U2139 ( .A(n1592), .B(n1593), .Z(n1589) );
  XNOR U2140 ( .A(y[175]), .B(x[175]), .Z(n1593) );
  XNOR U2141 ( .A(y[174]), .B(x[174]), .Z(n1592) );
  XNOR U2142 ( .A(n1590), .B(n1591), .Z(n1588) );
  XNOR U2143 ( .A(y[173]), .B(x[173]), .Z(n1591) );
  XNOR U2144 ( .A(y[172]), .B(x[172]), .Z(n1590) );
  XNOR U2145 ( .A(n1603), .B(n1604), .Z(n1596) );
  XNOR U2146 ( .A(n1598), .B(n1597), .Z(n1604) );
  XNOR U2147 ( .A(y[171]), .B(x[171]), .Z(n1597) );
  XNOR U2148 ( .A(y[170]), .B(x[170]), .Z(n1598) );
  XNOR U2149 ( .A(n1601), .B(n1602), .Z(n1603) );
  XNOR U2150 ( .A(y[169]), .B(x[169]), .Z(n1602) );
  XNOR U2151 ( .A(y[168]), .B(x[168]), .Z(n1601) );
  XNOR U2152 ( .A(n1609), .B(n1610), .Z(n1618) );
  XNOR U2153 ( .A(n1613), .B(n1614), .Z(n1610) );
  XNOR U2154 ( .A(y[167]), .B(x[167]), .Z(n1614) );
  XNOR U2155 ( .A(y[166]), .B(x[166]), .Z(n1613) );
  XNOR U2156 ( .A(n1611), .B(n1612), .Z(n1609) );
  XNOR U2157 ( .A(y[165]), .B(x[165]), .Z(n1612) );
  XNOR U2158 ( .A(y[164]), .B(x[164]), .Z(n1611) );
  XNOR U2159 ( .A(n1626), .B(n1627), .Z(n1619) );
  XNOR U2160 ( .A(n1621), .B(n1620), .Z(n1627) );
  XNOR U2161 ( .A(y[163]), .B(x[163]), .Z(n1620) );
  XNOR U2162 ( .A(y[162]), .B(x[162]), .Z(n1621) );
  XNOR U2163 ( .A(n1624), .B(n1625), .Z(n1626) );
  XNOR U2164 ( .A(y[161]), .B(x[161]), .Z(n1625) );
  XNOR U2165 ( .A(y[160]), .B(x[160]), .Z(n1624) );
  XNOR U2166 ( .A(n1692), .B(n1691), .Z(n1671) );
  XNOR U2167 ( .A(n1658), .B(n1657), .Z(n1691) );
  XNOR U2168 ( .A(n1632), .B(n1633), .Z(n1639) );
  XNOR U2169 ( .A(n1636), .B(n1637), .Z(n1633) );
  XNOR U2170 ( .A(y[159]), .B(x[159]), .Z(n1637) );
  XNOR U2171 ( .A(y[158]), .B(x[158]), .Z(n1636) );
  XNOR U2172 ( .A(n1634), .B(n1635), .Z(n1632) );
  XNOR U2173 ( .A(y[157]), .B(x[157]), .Z(n1635) );
  XNOR U2174 ( .A(y[156]), .B(x[156]), .Z(n1634) );
  XNOR U2175 ( .A(n1647), .B(n1648), .Z(n1640) );
  XNOR U2176 ( .A(n1642), .B(n1641), .Z(n1648) );
  XNOR U2177 ( .A(y[155]), .B(x[155]), .Z(n1641) );
  XNOR U2178 ( .A(y[154]), .B(x[154]), .Z(n1642) );
  XNOR U2179 ( .A(n1645), .B(n1646), .Z(n1647) );
  XNOR U2180 ( .A(y[153]), .B(x[153]), .Z(n1646) );
  XNOR U2181 ( .A(y[152]), .B(x[152]), .Z(n1645) );
  XNOR U2182 ( .A(n1651), .B(n1652), .Z(n1660) );
  XNOR U2183 ( .A(n1655), .B(n1656), .Z(n1652) );
  XNOR U2184 ( .A(y[151]), .B(x[151]), .Z(n1656) );
  XNOR U2185 ( .A(y[150]), .B(x[150]), .Z(n1655) );
  XNOR U2186 ( .A(n1653), .B(n1654), .Z(n1651) );
  XNOR U2187 ( .A(y[149]), .B(x[149]), .Z(n1654) );
  XNOR U2188 ( .A(y[148]), .B(x[148]), .Z(n1653) );
  XNOR U2189 ( .A(n1668), .B(n1669), .Z(n1661) );
  XNOR U2190 ( .A(n1663), .B(n1662), .Z(n1669) );
  XNOR U2191 ( .A(y[147]), .B(x[147]), .Z(n1662) );
  XNOR U2192 ( .A(y[146]), .B(x[146]), .Z(n1663) );
  XNOR U2193 ( .A(n1666), .B(n1667), .Z(n1668) );
  XNOR U2194 ( .A(y[145]), .B(x[145]), .Z(n1667) );
  XNOR U2195 ( .A(y[144]), .B(x[144]), .Z(n1666) );
  XNOR U2196 ( .A(n1702), .B(n1701), .Z(n1692) );
  XNOR U2197 ( .A(n1674), .B(n1675), .Z(n1681) );
  XNOR U2198 ( .A(n1678), .B(n1679), .Z(n1675) );
  XNOR U2199 ( .A(y[143]), .B(x[143]), .Z(n1679) );
  XNOR U2200 ( .A(y[142]), .B(x[142]), .Z(n1678) );
  XNOR U2201 ( .A(n1676), .B(n1677), .Z(n1674) );
  XNOR U2202 ( .A(y[141]), .B(x[141]), .Z(n1677) );
  XNOR U2203 ( .A(y[140]), .B(x[140]), .Z(n1676) );
  XNOR U2204 ( .A(n1689), .B(n1690), .Z(n1682) );
  XNOR U2205 ( .A(n1684), .B(n1683), .Z(n1690) );
  XNOR U2206 ( .A(y[139]), .B(x[139]), .Z(n1683) );
  XNOR U2207 ( .A(y[138]), .B(x[138]), .Z(n1684) );
  XNOR U2208 ( .A(n1687), .B(n1688), .Z(n1689) );
  XNOR U2209 ( .A(y[137]), .B(x[137]), .Z(n1688) );
  XNOR U2210 ( .A(y[136]), .B(x[136]), .Z(n1687) );
  XNOR U2211 ( .A(n1695), .B(n1696), .Z(n1704) );
  XNOR U2212 ( .A(n1699), .B(n1700), .Z(n1696) );
  XNOR U2213 ( .A(y[135]), .B(x[135]), .Z(n1700) );
  XNOR U2214 ( .A(y[134]), .B(x[134]), .Z(n1699) );
  XNOR U2215 ( .A(n1697), .B(n1698), .Z(n1695) );
  XNOR U2216 ( .A(y[133]), .B(x[133]), .Z(n1698) );
  XNOR U2217 ( .A(y[132]), .B(x[132]), .Z(n1697) );
  XNOR U2218 ( .A(n1712), .B(n1713), .Z(n1705) );
  XNOR U2219 ( .A(n1707), .B(n1706), .Z(n1713) );
  XNOR U2220 ( .A(y[131]), .B(x[131]), .Z(n1706) );
  XNOR U2221 ( .A(y[130]), .B(x[130]), .Z(n1707) );
  XNOR U2222 ( .A(n1710), .B(n1711), .Z(n1712) );
  XNOR U2223 ( .A(y[129]), .B(x[129]), .Z(n1711) );
  XNOR U2224 ( .A(y[128]), .B(x[128]), .Z(n1710) );
  XNOR U2225 ( .A(n1965), .B(n1964), .Z(n1881) );
  XNOR U2226 ( .A(n1837), .B(n1836), .Z(n1964) );
  XNOR U2227 ( .A(n1774), .B(n1773), .Z(n1836) );
  XNOR U2228 ( .A(n1742), .B(n1741), .Z(n1773) );
  XNOR U2229 ( .A(n1716), .B(n1717), .Z(n1723) );
  XNOR U2230 ( .A(n1720), .B(n1721), .Z(n1717) );
  XNOR U2231 ( .A(y[127]), .B(x[127]), .Z(n1721) );
  XNOR U2232 ( .A(y[126]), .B(x[126]), .Z(n1720) );
  XNOR U2233 ( .A(n1718), .B(n1719), .Z(n1716) );
  XNOR U2234 ( .A(y[125]), .B(x[125]), .Z(n1719) );
  XNOR U2235 ( .A(y[124]), .B(x[124]), .Z(n1718) );
  XNOR U2236 ( .A(n1731), .B(n1732), .Z(n1724) );
  XNOR U2237 ( .A(n1726), .B(n1725), .Z(n1732) );
  XNOR U2238 ( .A(y[123]), .B(x[123]), .Z(n1725) );
  XNOR U2239 ( .A(y[122]), .B(x[122]), .Z(n1726) );
  XNOR U2240 ( .A(n1729), .B(n1730), .Z(n1731) );
  XNOR U2241 ( .A(y[121]), .B(x[121]), .Z(n1730) );
  XNOR U2242 ( .A(y[120]), .B(x[120]), .Z(n1729) );
  XNOR U2243 ( .A(n1735), .B(n1736), .Z(n1744) );
  XNOR U2244 ( .A(n1739), .B(n1740), .Z(n1736) );
  XNOR U2245 ( .A(y[119]), .B(x[119]), .Z(n1740) );
  XNOR U2246 ( .A(y[118]), .B(x[118]), .Z(n1739) );
  XNOR U2247 ( .A(n1737), .B(n1738), .Z(n1735) );
  XNOR U2248 ( .A(y[117]), .B(x[117]), .Z(n1738) );
  XNOR U2249 ( .A(y[116]), .B(x[116]), .Z(n1737) );
  XNOR U2250 ( .A(n1752), .B(n1753), .Z(n1745) );
  XNOR U2251 ( .A(n1747), .B(n1746), .Z(n1753) );
  XNOR U2252 ( .A(y[115]), .B(x[115]), .Z(n1746) );
  XNOR U2253 ( .A(y[114]), .B(x[114]), .Z(n1747) );
  XNOR U2254 ( .A(n1750), .B(n1751), .Z(n1752) );
  XNOR U2255 ( .A(y[113]), .B(x[113]), .Z(n1751) );
  XNOR U2256 ( .A(y[112]), .B(x[112]), .Z(n1750) );
  XNOR U2257 ( .A(n1784), .B(n1783), .Z(n1774) );
  XNOR U2258 ( .A(n1756), .B(n1757), .Z(n1763) );
  XNOR U2259 ( .A(n1760), .B(n1761), .Z(n1757) );
  XNOR U2260 ( .A(y[111]), .B(x[111]), .Z(n1761) );
  XNOR U2261 ( .A(y[110]), .B(x[110]), .Z(n1760) );
  XNOR U2262 ( .A(n1758), .B(n1759), .Z(n1756) );
  XNOR U2263 ( .A(y[109]), .B(x[109]), .Z(n1759) );
  XNOR U2264 ( .A(y[108]), .B(x[108]), .Z(n1758) );
  XNOR U2265 ( .A(n1771), .B(n1772), .Z(n1764) );
  XNOR U2266 ( .A(n1766), .B(n1765), .Z(n1772) );
  XNOR U2267 ( .A(y[107]), .B(x[107]), .Z(n1765) );
  XNOR U2268 ( .A(y[106]), .B(x[106]), .Z(n1766) );
  XNOR U2269 ( .A(n1769), .B(n1770), .Z(n1771) );
  XNOR U2270 ( .A(y[105]), .B(x[105]), .Z(n1770) );
  XNOR U2271 ( .A(y[104]), .B(x[104]), .Z(n1769) );
  XNOR U2272 ( .A(n1777), .B(n1778), .Z(n1786) );
  XNOR U2273 ( .A(n1781), .B(n1782), .Z(n1778) );
  XNOR U2274 ( .A(y[103]), .B(x[103]), .Z(n1782) );
  XNOR U2275 ( .A(y[102]), .B(x[102]), .Z(n1781) );
  XNOR U2276 ( .A(n1779), .B(n1780), .Z(n1777) );
  XNOR U2277 ( .A(y[101]), .B(x[101]), .Z(n1780) );
  XNOR U2278 ( .A(y[100]), .B(x[100]), .Z(n1779) );
  XNOR U2279 ( .A(n1794), .B(n1795), .Z(n1787) );
  XNOR U2280 ( .A(n1789), .B(n1788), .Z(n1795) );
  XNOR U2281 ( .A(y[99]), .B(x[99]), .Z(n1788) );
  XNOR U2282 ( .A(y[98]), .B(x[98]), .Z(n1789) );
  XNOR U2283 ( .A(n1792), .B(n1793), .Z(n1794) );
  XNOR U2284 ( .A(y[97]), .B(x[97]), .Z(n1793) );
  XNOR U2285 ( .A(y[96]), .B(x[96]), .Z(n1792) );
  XNOR U2286 ( .A(n1858), .B(n1857), .Z(n1837) );
  XNOR U2287 ( .A(n1824), .B(n1823), .Z(n1857) );
  XNOR U2288 ( .A(n1798), .B(n1799), .Z(n1805) );
  XNOR U2289 ( .A(n1802), .B(n1803), .Z(n1799) );
  XNOR U2290 ( .A(y[95]), .B(x[95]), .Z(n1803) );
  XNOR U2291 ( .A(y[94]), .B(x[94]), .Z(n1802) );
  XNOR U2292 ( .A(n1800), .B(n1801), .Z(n1798) );
  XNOR U2293 ( .A(y[93]), .B(x[93]), .Z(n1801) );
  XNOR U2294 ( .A(y[92]), .B(x[92]), .Z(n1800) );
  XNOR U2295 ( .A(n1813), .B(n1814), .Z(n1806) );
  XNOR U2296 ( .A(n1808), .B(n1807), .Z(n1814) );
  XNOR U2297 ( .A(y[91]), .B(x[91]), .Z(n1807) );
  XNOR U2298 ( .A(y[90]), .B(x[90]), .Z(n1808) );
  XNOR U2299 ( .A(n1811), .B(n1812), .Z(n1813) );
  XNOR U2300 ( .A(y[89]), .B(x[89]), .Z(n1812) );
  XNOR U2301 ( .A(y[88]), .B(x[88]), .Z(n1811) );
  XNOR U2302 ( .A(n1817), .B(n1818), .Z(n1826) );
  XNOR U2303 ( .A(n1821), .B(n1822), .Z(n1818) );
  XNOR U2304 ( .A(y[87]), .B(x[87]), .Z(n1822) );
  XNOR U2305 ( .A(y[86]), .B(x[86]), .Z(n1821) );
  XNOR U2306 ( .A(n1819), .B(n1820), .Z(n1817) );
  XNOR U2307 ( .A(y[85]), .B(x[85]), .Z(n1820) );
  XNOR U2308 ( .A(y[84]), .B(x[84]), .Z(n1819) );
  XNOR U2309 ( .A(n1834), .B(n1835), .Z(n1827) );
  XNOR U2310 ( .A(n1829), .B(n1828), .Z(n1835) );
  XNOR U2311 ( .A(y[83]), .B(x[83]), .Z(n1828) );
  XNOR U2312 ( .A(y[82]), .B(x[82]), .Z(n1829) );
  XNOR U2313 ( .A(n1832), .B(n1833), .Z(n1834) );
  XNOR U2314 ( .A(y[81]), .B(x[81]), .Z(n1833) );
  XNOR U2315 ( .A(y[80]), .B(x[80]), .Z(n1832) );
  XNOR U2316 ( .A(n1868), .B(n1867), .Z(n1858) );
  XNOR U2317 ( .A(n1840), .B(n1841), .Z(n1847) );
  XNOR U2318 ( .A(n1844), .B(n1845), .Z(n1841) );
  XNOR U2319 ( .A(y[79]), .B(x[79]), .Z(n1845) );
  XNOR U2320 ( .A(y[78]), .B(x[78]), .Z(n1844) );
  XNOR U2321 ( .A(n1842), .B(n1843), .Z(n1840) );
  XNOR U2322 ( .A(y[77]), .B(x[77]), .Z(n1843) );
  XNOR U2323 ( .A(y[76]), .B(x[76]), .Z(n1842) );
  XNOR U2324 ( .A(n1855), .B(n1856), .Z(n1848) );
  XNOR U2325 ( .A(n1850), .B(n1849), .Z(n1856) );
  XNOR U2326 ( .A(y[75]), .B(x[75]), .Z(n1849) );
  XNOR U2327 ( .A(y[74]), .B(x[74]), .Z(n1850) );
  XNOR U2328 ( .A(n1853), .B(n1854), .Z(n1855) );
  XNOR U2329 ( .A(y[73]), .B(x[73]), .Z(n1854) );
  XNOR U2330 ( .A(y[72]), .B(x[72]), .Z(n1853) );
  XNOR U2331 ( .A(n1861), .B(n1862), .Z(n1870) );
  XNOR U2332 ( .A(n1865), .B(n1866), .Z(n1862) );
  XNOR U2333 ( .A(y[71]), .B(x[71]), .Z(n1866) );
  XNOR U2334 ( .A(y[70]), .B(x[70]), .Z(n1865) );
  XNOR U2335 ( .A(n1863), .B(n1864), .Z(n1861) );
  XNOR U2336 ( .A(y[69]), .B(x[69]), .Z(n1864) );
  XNOR U2337 ( .A(y[68]), .B(x[68]), .Z(n1863) );
  XNOR U2338 ( .A(n1878), .B(n1879), .Z(n1871) );
  XNOR U2339 ( .A(n1873), .B(n1872), .Z(n1879) );
  XNOR U2340 ( .A(y[67]), .B(x[67]), .Z(n1872) );
  XNOR U2341 ( .A(y[66]), .B(x[66]), .Z(n1873) );
  XNOR U2342 ( .A(n1876), .B(n1877), .Z(n1878) );
  XNOR U2343 ( .A(y[65]), .B(x[65]), .Z(n1877) );
  XNOR U2344 ( .A(y[64]), .B(x[64]), .Z(n1876) );
  XNOR U2345 ( .A(n2007), .B(n2006), .Z(n1965) );
  XNOR U2346 ( .A(n1942), .B(n1941), .Z(n2006) );
  XNOR U2347 ( .A(n1910), .B(n1909), .Z(n1941) );
  XNOR U2348 ( .A(n1884), .B(n1885), .Z(n1891) );
  XNOR U2349 ( .A(n1888), .B(n1889), .Z(n1885) );
  XNOR U2350 ( .A(y[63]), .B(x[63]), .Z(n1889) );
  XNOR U2351 ( .A(y[62]), .B(x[62]), .Z(n1888) );
  XNOR U2352 ( .A(n1886), .B(n1887), .Z(n1884) );
  XNOR U2353 ( .A(y[61]), .B(x[61]), .Z(n1887) );
  XNOR U2354 ( .A(y[60]), .B(x[60]), .Z(n1886) );
  XNOR U2355 ( .A(n1899), .B(n1900), .Z(n1892) );
  XNOR U2356 ( .A(n1894), .B(n1893), .Z(n1900) );
  XNOR U2357 ( .A(y[59]), .B(x[59]), .Z(n1893) );
  XNOR U2358 ( .A(y[58]), .B(x[58]), .Z(n1894) );
  XNOR U2359 ( .A(n1897), .B(n1898), .Z(n1899) );
  XNOR U2360 ( .A(y[57]), .B(x[57]), .Z(n1898) );
  XNOR U2361 ( .A(y[56]), .B(x[56]), .Z(n1897) );
  XNOR U2362 ( .A(n1903), .B(n1904), .Z(n1912) );
  XNOR U2363 ( .A(n1907), .B(n1908), .Z(n1904) );
  XNOR U2364 ( .A(y[55]), .B(x[55]), .Z(n1908) );
  XNOR U2365 ( .A(y[54]), .B(x[54]), .Z(n1907) );
  XNOR U2366 ( .A(n1905), .B(n1906), .Z(n1903) );
  XNOR U2367 ( .A(y[53]), .B(x[53]), .Z(n1906) );
  XNOR U2368 ( .A(y[52]), .B(x[52]), .Z(n1905) );
  XNOR U2369 ( .A(n1920), .B(n1921), .Z(n1913) );
  XNOR U2370 ( .A(n1915), .B(n1914), .Z(n1921) );
  XNOR U2371 ( .A(y[51]), .B(x[51]), .Z(n1914) );
  XNOR U2372 ( .A(y[50]), .B(x[50]), .Z(n1915) );
  XNOR U2373 ( .A(n1918), .B(n1919), .Z(n1920) );
  XNOR U2374 ( .A(y[49]), .B(x[49]), .Z(n1919) );
  XNOR U2375 ( .A(y[48]), .B(x[48]), .Z(n1918) );
  XNOR U2376 ( .A(n1952), .B(n1951), .Z(n1942) );
  XNOR U2377 ( .A(n1924), .B(n1925), .Z(n1931) );
  XNOR U2378 ( .A(n1928), .B(n1929), .Z(n1925) );
  XNOR U2379 ( .A(y[47]), .B(x[47]), .Z(n1929) );
  XNOR U2380 ( .A(y[46]), .B(x[46]), .Z(n1928) );
  XNOR U2381 ( .A(n1926), .B(n1927), .Z(n1924) );
  XNOR U2382 ( .A(y[45]), .B(x[45]), .Z(n1927) );
  XNOR U2383 ( .A(y[44]), .B(x[44]), .Z(n1926) );
  XNOR U2384 ( .A(n1939), .B(n1940), .Z(n1932) );
  XNOR U2385 ( .A(n1934), .B(n1933), .Z(n1940) );
  XNOR U2386 ( .A(y[43]), .B(x[43]), .Z(n1933) );
  XNOR U2387 ( .A(y[42]), .B(x[42]), .Z(n1934) );
  XNOR U2388 ( .A(n1937), .B(n1938), .Z(n1939) );
  XNOR U2389 ( .A(y[41]), .B(x[41]), .Z(n1938) );
  XNOR U2390 ( .A(y[40]), .B(x[40]), .Z(n1937) );
  XNOR U2391 ( .A(n1945), .B(n1946), .Z(n1954) );
  XNOR U2392 ( .A(n1949), .B(n1950), .Z(n1946) );
  XNOR U2393 ( .A(y[39]), .B(x[39]), .Z(n1950) );
  XNOR U2394 ( .A(y[38]), .B(x[38]), .Z(n1949) );
  XNOR U2395 ( .A(n1947), .B(n1948), .Z(n1945) );
  XNOR U2396 ( .A(y[37]), .B(x[37]), .Z(n1948) );
  XNOR U2397 ( .A(y[36]), .B(x[36]), .Z(n1947) );
  XNOR U2398 ( .A(n1962), .B(n1963), .Z(n1955) );
  XNOR U2399 ( .A(n1957), .B(n1956), .Z(n1963) );
  XNOR U2400 ( .A(y[35]), .B(x[35]), .Z(n1956) );
  XNOR U2401 ( .A(y[34]), .B(x[34]), .Z(n1957) );
  XNOR U2402 ( .A(n1960), .B(n1961), .Z(n1962) );
  XNOR U2403 ( .A(y[33]), .B(x[33]), .Z(n1961) );
  XNOR U2404 ( .A(y[32]), .B(x[32]), .Z(n1960) );
  XNOR U2405 ( .A(n2028), .B(n2027), .Z(n2007) );
  XNOR U2406 ( .A(n1994), .B(n1993), .Z(n2027) );
  XNOR U2407 ( .A(n1968), .B(n1969), .Z(n1975) );
  XNOR U2408 ( .A(n1972), .B(n1973), .Z(n1969) );
  XNOR U2409 ( .A(y[31]), .B(x[31]), .Z(n1973) );
  XNOR U2410 ( .A(y[30]), .B(x[30]), .Z(n1972) );
  XNOR U2411 ( .A(n1970), .B(n1971), .Z(n1968) );
  XNOR U2412 ( .A(y[29]), .B(x[29]), .Z(n1971) );
  XNOR U2413 ( .A(y[28]), .B(x[28]), .Z(n1970) );
  XNOR U2414 ( .A(n1983), .B(n1984), .Z(n1976) );
  XNOR U2415 ( .A(n1978), .B(n1977), .Z(n1984) );
  XNOR U2416 ( .A(y[27]), .B(x[27]), .Z(n1977) );
  XNOR U2417 ( .A(y[26]), .B(x[26]), .Z(n1978) );
  XNOR U2418 ( .A(n1981), .B(n1982), .Z(n1983) );
  XNOR U2419 ( .A(y[25]), .B(x[25]), .Z(n1982) );
  XNOR U2420 ( .A(y[24]), .B(x[24]), .Z(n1981) );
  XNOR U2421 ( .A(n1987), .B(n1988), .Z(n1996) );
  XNOR U2422 ( .A(n1991), .B(n1992), .Z(n1988) );
  XNOR U2423 ( .A(y[23]), .B(x[23]), .Z(n1992) );
  XNOR U2424 ( .A(y[22]), .B(x[22]), .Z(n1991) );
  XNOR U2425 ( .A(n1989), .B(n1990), .Z(n1987) );
  XNOR U2426 ( .A(y[21]), .B(x[21]), .Z(n1990) );
  XNOR U2427 ( .A(y[20]), .B(x[20]), .Z(n1989) );
  XNOR U2428 ( .A(n2004), .B(n2005), .Z(n1997) );
  XNOR U2429 ( .A(n1999), .B(n1998), .Z(n2005) );
  XNOR U2430 ( .A(y[19]), .B(x[19]), .Z(n1998) );
  XNOR U2431 ( .A(y[18]), .B(x[18]), .Z(n1999) );
  XNOR U2432 ( .A(n2002), .B(n2003), .Z(n2004) );
  XNOR U2433 ( .A(y[17]), .B(x[17]), .Z(n2003) );
  XNOR U2434 ( .A(y[16]), .B(x[16]), .Z(n2002) );
  XNOR U2435 ( .A(n2038), .B(n2037), .Z(n2028) );
  XNOR U2436 ( .A(n2010), .B(n2011), .Z(n2017) );
  XNOR U2437 ( .A(n2014), .B(n2015), .Z(n2011) );
  XNOR U2438 ( .A(y[15]), .B(x[15]), .Z(n2015) );
  XNOR U2439 ( .A(y[14]), .B(x[14]), .Z(n2014) );
  XNOR U2440 ( .A(n2012), .B(n2013), .Z(n2010) );
  XNOR U2441 ( .A(y[13]), .B(x[13]), .Z(n2013) );
  XNOR U2442 ( .A(y[12]), .B(x[12]), .Z(n2012) );
  XNOR U2443 ( .A(n2025), .B(n2026), .Z(n2018) );
  XNOR U2444 ( .A(n2020), .B(n2019), .Z(n2026) );
  XNOR U2445 ( .A(y[11]), .B(x[11]), .Z(n2019) );
  XNOR U2446 ( .A(y[10]), .B(x[10]), .Z(n2020) );
  XNOR U2447 ( .A(n2023), .B(n2024), .Z(n2025) );
  XNOR U2448 ( .A(y[9]), .B(x[9]), .Z(n2024) );
  XNOR U2449 ( .A(y[8]), .B(x[8]), .Z(n2023) );
  XNOR U2450 ( .A(n2031), .B(n2032), .Z(n2040) );
  XNOR U2451 ( .A(n2035), .B(n2036), .Z(n2032) );
  XNOR U2452 ( .A(y[7]), .B(x[7]), .Z(n2036) );
  XNOR U2453 ( .A(y[6]), .B(x[6]), .Z(n2035) );
  XNOR U2454 ( .A(n2033), .B(n2034), .Z(n2031) );
  XNOR U2455 ( .A(y[5]), .B(x[5]), .Z(n2034) );
  XNOR U2456 ( .A(y[4]), .B(x[4]), .Z(n2033) );
  XNOR U2457 ( .A(n2048), .B(n2049), .Z(n2041) );
  XNOR U2458 ( .A(n2043), .B(n2042), .Z(n2049) );
  XNOR U2459 ( .A(y[3]), .B(x[3]), .Z(n2042) );
  XNOR U2460 ( .A(y[2]), .B(x[2]), .Z(n2043) );
  XNOR U2461 ( .A(n2046), .B(n2047), .Z(n2048) );
  XNOR U2462 ( .A(y[1]), .B(x[1]), .Z(n2047) );
  XNOR U2463 ( .A(y[0]), .B(x[0]), .Z(n2046) );
endmodule

