
module hamming_N1600_CC1 ( clk, rst, x, y, o );
  input [1599:0] x;
  input [1599:0] y;
  output [10:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686;

  MUX U1601 ( .IN0(n5970), .IN1(n5968), .SEL(n5969), .F(n1) );
  IV U1602 ( .A(n1), .Z(n4523) );
  MUX U1603 ( .IN0(n5507), .IN1(n5505), .SEL(n5506), .F(n2) );
  IV U1604 ( .A(n2), .Z(n4262) );
  MUX U1605 ( .IN0(n6761), .IN1(n6759), .SEL(n6760), .F(n6755) );
  MUX U1606 ( .IN0(n6546), .IN1(n6544), .SEL(n6545), .F(n3) );
  IV U1607 ( .A(n3), .Z(n4844) );
  MUX U1608 ( .IN0(n205), .IN1(n4896), .SEL(n4895), .F(n4) );
  IV U1609 ( .A(n4), .Z(n3928) );
  MUX U1610 ( .IN0(n6120), .IN1(n6118), .SEL(n6119), .F(n6114) );
  MUX U1611 ( .IN0(n302), .IN1(n4669), .SEL(n4668), .F(n5) );
  IV U1612 ( .A(n5), .Z(n3820) );
  MUX U1613 ( .IN0(n5170), .IN1(n5168), .SEL(n5169), .F(n5164) );
  MUX U1614 ( .IN0(n5177), .IN1(n5175), .SEL(n5176), .F(n5171) );
  MUX U1615 ( .IN0(n5262), .IN1(n5260), .SEL(n5261), .F(n5256) );
  MUX U1616 ( .IN0(n5420), .IN1(n5418), .SEL(n5419), .F(n6) );
  IV U1617 ( .A(n6), .Z(n4210) );
  MUX U1618 ( .IN0(n5277), .IN1(n5275), .SEL(n5276), .F(n7) );
  IV U1619 ( .A(n7), .Z(n4131) );
  MUX U1620 ( .IN0(n637), .IN1(n4180), .SEL(n4179), .F(n8) );
  IV U1621 ( .A(n8), .Z(n3577) );
  MUX U1622 ( .IN0(n5657), .IN1(n5655), .SEL(n5656), .F(n5651) );
  MUX U1623 ( .IN0(n5606), .IN1(n5604), .SEL(n5605), .F(n5600) );
  MUX U1624 ( .IN0(n5775), .IN1(n5773), .SEL(n5774), .F(n5769) );
  MUX U1625 ( .IN0(n5782), .IN1(n5780), .SEL(n5781), .F(n5776) );
  XOR U1626 ( .A(n1486), .B(n1484), .Z(n1478) );
  MUX U1627 ( .IN0(n79), .IN1(n1752), .SEL(n1751), .F(n9) );
  IV U1628 ( .A(n9), .Z(n1288) );
  MUX U1629 ( .IN0(n2764), .IN1(n2762), .SEL(n2763), .F(n10) );
  IV U1630 ( .A(n10), .Z(n1845) );
  MUX U1631 ( .IN0(n147), .IN1(n1937), .SEL(n1936), .F(n11) );
  IV U1632 ( .A(n11), .Z(n1373) );
  MUX U1633 ( .IN0(n2793), .IN1(n2791), .SEL(n2792), .F(n12) );
  IV U1634 ( .A(n12), .Z(n1864) );
  MUX U1635 ( .IN0(n674), .IN1(n1546), .SEL(n1545), .F(n13) );
  IV U1636 ( .A(n13), .Z(n1184) );
  MUX U1637 ( .IN0(n146), .IN1(n1513), .SEL(n1512), .F(n14) );
  IV U1638 ( .A(n14), .Z(n1168) );
  MUX U1639 ( .IN0(n295), .IN1(n1639), .SEL(n1638), .F(n15) );
  IV U1640 ( .A(n15), .Z(n1234) );
  MUX U1641 ( .IN0(n89), .IN1(n1705), .SEL(n1704), .F(n16) );
  IV U1642 ( .A(n16), .Z(n1263) );
  MUX U1643 ( .IN0(n598), .IN1(n4955), .SEL(n4953), .F(n4949) );
  MUX U1644 ( .IN0(n486), .IN1(n4581), .SEL(n4579), .F(n3773) );
  MUX U1645 ( .IN0(n627), .IN1(n4772), .SEL(n4770), .F(n4763) );
  MUX U1646 ( .IN0(n581), .IN1(n4120), .SEL(n4118), .F(n4113) );
  MUX U1647 ( .IN0(n499), .IN1(n4316), .SEL(n4314), .F(n4307) );
  MUX U1648 ( .IN0(n506), .IN1(n4518), .SEL(n4516), .F(n3741) );
  MUX U1649 ( .IN0(n584), .IN1(n1748), .SEL(n1746), .F(n1741) );
  MUX U1650 ( .IN0(n70), .IN1(n1316), .SEL(n1315), .F(n17) );
  IV U1651 ( .A(n17), .Z(n1068) );
  MUX U1652 ( .IN0(n427), .IN1(n1609), .SEL(n1608), .F(n18) );
  IV U1653 ( .A(n18), .Z(n1216) );
  MUX U1654 ( .IN0(n3905), .IN1(n19), .SEL(n3906), .F(n3439) );
  IV U1655 ( .A(n3907), .Z(n19) );
  MUX U1656 ( .IN0(n3758), .IN1(n3761), .SEL(n3759), .F(n3754) );
  MUX U1657 ( .IN0(n3766), .IN1(n3769), .SEL(n3767), .F(n3762) );
  MUX U1658 ( .IN0(n3862), .IN1(n3865), .SEL(n3863), .F(n3856) );
  MUX U1659 ( .IN0(n3540), .IN1(n3543), .SEL(n3541), .F(n3534) );
  MUX U1660 ( .IN0(n2058), .IN1(n2056), .SEL(n2057), .F(n20) );
  IV U1661 ( .A(n20), .Z(n1441) );
  MUX U1662 ( .IN0(n263), .IN1(n4680), .SEL(n4679), .F(n21) );
  IV U1663 ( .A(n21), .Z(n3822) );
  XOR U1664 ( .A(n1045), .B(n1043), .Z(n1037) );
  XOR U1665 ( .A(n1095), .B(n1094), .Z(n1088) );
  MUX U1666 ( .IN0(n2038), .IN1(n2036), .SEL(n2037), .F(n2032) );
  MUX U1667 ( .IN0(n2045), .IN1(n2043), .SEL(n2044), .F(n2039) );
  MUX U1668 ( .IN0(n987), .IN1(n22), .SEL(n988), .F(n905) );
  IV U1669 ( .A(n989), .Z(n22) );
  MUX U1670 ( .IN0(n3414), .IN1(n3417), .SEL(n3415), .F(n3410) );
  MUX U1671 ( .IN0(n3154), .IN1(n23), .SEL(n3155), .F(n3077) );
  IV U1672 ( .A(n3156), .Z(n23) );
  MUX U1673 ( .IN0(n934), .IN1(n24), .SEL(n935), .F(n877) );
  IV U1674 ( .A(n936), .Z(n24) );
  MUX U1675 ( .IN0(n907), .IN1(n25), .SEL(n908), .F(n860) );
  IV U1676 ( .A(n909), .Z(n25) );
  MUX U1677 ( .IN0(n3198), .IN1(n3201), .SEL(n3199), .F(n3194) );
  MUX U1678 ( .IN0(n3169), .IN1(n3172), .SEL(n3170), .F(n3165) );
  MUX U1679 ( .IN0(n2964), .IN1(n2962), .SEL(n2963), .F(n26) );
  IV U1680 ( .A(n26), .Z(n1965) );
  MUX U1681 ( .IN0(n2539), .IN1(n2537), .SEL(n2538), .F(n27) );
  IV U1682 ( .A(n27), .Z(n1716) );
  MUX U1683 ( .IN0(n6847), .IN1(n6845), .SEL(n6846), .F(n6839) );
  MUX U1684 ( .IN0(n6803), .IN1(n6801), .SEL(n6802), .F(n28) );
  IV U1685 ( .A(n28), .Z(n4991) );
  MUX U1686 ( .IN0(n6669), .IN1(n6667), .SEL(n6668), .F(n6663) );
  MUX U1687 ( .IN0(n6676), .IN1(n6674), .SEL(n6675), .F(n6670) );
  MUX U1688 ( .IN0(n6486), .IN1(n6484), .SEL(n6485), .F(n29) );
  IV U1689 ( .A(n29), .Z(n4812) );
  MUX U1690 ( .IN0(n6472), .IN1(n6470), .SEL(n6471), .F(n6464) );
  MUX U1691 ( .IN0(n6553), .IN1(n6551), .SEL(n6552), .F(n6547) );
  XOR U1692 ( .A(n6640), .B(n6641), .Z(n4901) );
  MUX U1693 ( .IN0(n6108), .IN1(n6106), .SEL(n6107), .F(n4611) );
  MUX U1694 ( .IN0(n6331), .IN1(n6329), .SEL(n6330), .F(n6325) );
  MUX U1695 ( .IN0(n5103), .IN1(n5101), .SEL(n5102), .F(n30) );
  IV U1696 ( .A(n30), .Z(n4036) );
  MUX U1697 ( .IN0(n5427), .IN1(n5425), .SEL(n5426), .F(n5421) );
  MUX U1698 ( .IN0(n5284), .IN1(n5282), .SEL(n5283), .F(n5278) );
  MUX U1699 ( .IN0(n5378), .IN1(n5376), .SEL(n5377), .F(n5372) );
  XOR U1700 ( .A(n5659), .B(n5660), .Z(n4353) );
  MUX U1701 ( .IN0(n4262), .IN1(n31), .SEL(n4263), .F(n3618) );
  IV U1702 ( .A(n4264), .Z(n31) );
  MUX U1703 ( .IN0(n5599), .IN1(n5597), .SEL(n5598), .F(n5593) );
  MUX U1704 ( .IN0(n32), .IN1(n5607), .SEL(n5608), .F(n4320) );
  IV U1705 ( .A(n5609), .Z(n32) );
  MUX U1706 ( .IN0(n5803), .IN1(n5801), .SEL(n5802), .F(n5797) );
  MUX U1707 ( .IN0(n5812), .IN1(n5810), .SEL(n5811), .F(n5804) );
  MUX U1708 ( .IN0(n5916), .IN1(n5914), .SEL(n5915), .F(n5910) );
  MUX U1709 ( .IN0(n5957), .IN1(n5955), .SEL(n5956), .F(n5951) );
  XOR U1710 ( .A(n1807), .B(n1806), .Z(n1800) );
  XOR U1711 ( .A(n4533), .B(n4531), .Z(n4525) );
  XOR U1712 ( .A(n4614), .B(n4613), .Z(n4607) );
  MUX U1713 ( .IN0(n6433), .IN1(n6435), .SEL(n6434), .F(n33) );
  IV U1714 ( .A(n33), .Z(n4783) );
  XOR U1715 ( .A(n4222), .B(n4220), .Z(n4214) );
  MUX U1716 ( .IN0(n148), .IN1(n4657), .SEL(n4656), .F(n34) );
  IV U1717 ( .A(n34), .Z(n3811) );
  MUX U1718 ( .IN0(n2771), .IN1(n2769), .SEL(n2770), .F(n2765) );
  MUX U1719 ( .IN0(n2778), .IN1(n2776), .SEL(n2777), .F(n2772) );
  MUX U1720 ( .IN0(n2800), .IN1(n2798), .SEL(n2799), .F(n2794) );
  MUX U1721 ( .IN0(n216), .IN1(n1574), .SEL(n1573), .F(n35) );
  IV U1722 ( .A(n35), .Z(n1201) );
  MUX U1723 ( .IN0(n2271), .IN1(n2269), .SEL(n2270), .F(n2265) );
  MUX U1724 ( .IN0(n2132), .IN1(n2130), .SEL(n2131), .F(n2126) );
  MUX U1725 ( .IN0(n2412), .IN1(n2410), .SEL(n2411), .F(n2406) );
  MUX U1726 ( .IN0(n2369), .IN1(n2367), .SEL(n2368), .F(n36) );
  IV U1727 ( .A(n36), .Z(n1619) );
  XNOR U1728 ( .A(n4795), .B(n4796), .Z(n3880) );
  MUX U1729 ( .IN0(n606), .IN1(n4892), .SEL(n4890), .F(n4885) );
  MUX U1730 ( .IN0(n620), .IN1(n4673), .SEL(n4671), .F(n4666) );
  MUX U1731 ( .IN0(n239), .IN1(n4754), .SEL(n4753), .F(n37) );
  IV U1732 ( .A(n37), .Z(n3857) );
  MUX U1733 ( .IN0(n628), .IN1(n4776), .SEL(n4774), .F(n3869) );
  MUX U1734 ( .IN0(n493), .IN1(n4184), .SEL(n4182), .F(n4177) );
  MUX U1735 ( .IN0(n91), .IN1(n4334), .SEL(n4333), .F(n38) );
  IV U1736 ( .A(n38), .Z(n3650) );
  MUX U1737 ( .IN0(n241), .IN1(n4399), .SEL(n4398), .F(n39) );
  IV U1738 ( .A(n39), .Z(n3682) );
  XOR U1739 ( .A(n1752), .B(n1751), .Z(n1740) );
  MUX U1740 ( .IN0(n5876), .IN1(n5878), .SEL(n5877), .F(n40) );
  IV U1741 ( .A(n40), .Z(n4469) );
  XOR U1742 ( .A(n1382), .B(n1381), .Z(n1375) );
  XOR U1743 ( .A(n1250), .B(n1249), .Z(n1257) );
  XOR U1744 ( .A(n3962), .B(n3961), .Z(n3955) );
  MUX U1745 ( .IN0(n106), .IN1(n3622), .SEL(n3621), .F(n41) );
  IV U1746 ( .A(n41), .Z(n3304) );
  MUX U1747 ( .IN0(n585), .IN1(n1735), .SEL(n1733), .F(n1285) );
  MUX U1748 ( .IN0(n156), .IN1(n1903), .SEL(n1902), .F(n42) );
  IV U1749 ( .A(n42), .Z(n1356) );
  MUX U1750 ( .IN0(n675), .IN1(n1554), .SEL(n1552), .F(n1547) );
  MUX U1751 ( .IN0(n677), .IN1(n1562), .SEL(n1560), .F(n1555) );
  MUX U1752 ( .IN0(n680), .IN1(n1482), .SEL(n1480), .F(n1475) );
  MUX U1753 ( .IN0(n522), .IN1(n1534), .SEL(n1532), .F(n1178) );
  MUX U1754 ( .IN0(n172), .IN1(n3458), .SEL(n3457), .F(n43) );
  IV U1755 ( .A(n43), .Z(n3226) );
  MUX U1756 ( .IN0(n3770), .IN1(n3773), .SEL(n3771), .F(n3375) );
  MUX U1757 ( .IN0(n3544), .IN1(n3547), .SEL(n3545), .F(n3267) );
  MUX U1758 ( .IN0(n3571), .IN1(n3574), .SEL(n3572), .F(n3567) );
  XOR U1759 ( .A(n1265), .B(n1264), .Z(n1253) );
  XOR U1760 ( .A(n1220), .B(n1219), .Z(n1238) );
  MUX U1761 ( .IN0(n3399), .IN1(n44), .SEL(n3400), .F(n3195) );
  IV U1762 ( .A(n3401), .Z(n44) );
  MUX U1763 ( .IN0(n1441), .IN1(n45), .SEL(n1442), .F(n1137) );
  IV U1764 ( .A(n1443), .Z(n45) );
  MUX U1765 ( .IN0(n1329), .IN1(n1332), .SEL(n1330), .F(n1325) );
  MUX U1766 ( .IN0(n1163), .IN1(n1166), .SEL(n1164), .F(n1159) );
  MUX U1767 ( .IN0(n541), .IN1(n1174), .SEL(n1172), .F(n1167) );
  MUX U1768 ( .IN0(n3427), .IN1(n46), .SEL(n3428), .F(n3208) );
  IV U1769 ( .A(n3429), .Z(n46) );
  XNOR U1770 ( .A(n3439), .B(n3440), .Z(n3217) );
  MUX U1771 ( .IN0(n3368), .IN1(n3371), .SEL(n3369), .F(n3364) );
  MUX U1772 ( .IN0(n3260), .IN1(n3263), .SEL(n3261), .F(n3256) );
  XOR U1773 ( .A(n1037), .B(n1036), .Z(n1025) );
  XOR U1774 ( .A(n1088), .B(n1087), .Z(n1106) );
  MUX U1775 ( .IN0(n3645), .IN1(n47), .SEL(n3646), .F(n3315) );
  IV U1776 ( .A(n3647), .Z(n47) );
  MUX U1777 ( .IN0(n367), .IN1(n1414), .SEL(n1413), .F(n48) );
  IV U1778 ( .A(n48), .Z(n1122) );
  XNOR U1779 ( .A(n1424), .B(n1425), .Z(n1129) );
  MUX U1780 ( .IN0(n1063), .IN1(n1066), .SEL(n1064), .F(n1059) );
  MUX U1781 ( .IN0(n1071), .IN1(n1074), .SEL(n1072), .F(n1067) );
  MUX U1782 ( .IN0(n3190), .IN1(n3193), .SEL(n3191), .F(n3186) );
  MUX U1783 ( .IN0(n3122), .IN1(n3125), .SEL(n3123), .F(n3118) );
  MUX U1784 ( .IN0(n3173), .IN1(n3176), .SEL(n3174), .F(n3087) );
  XOR U1785 ( .A(n870), .B(n868), .Z(n862) );
  XOR U1786 ( .A(n3100), .B(n3098), .Z(n3092) );
  MUX U1787 ( .IN0(n3080), .IN1(n3083), .SEL(n3081), .F(n3076) );
  MUX U1788 ( .IN0(n6286), .IN1(n6284), .SEL(n6285), .F(n49) );
  IV U1789 ( .A(n49), .Z(n4702) );
  MUX U1790 ( .IN0(n6400), .IN1(n6398), .SEL(n6399), .F(n50) );
  IV U1791 ( .A(n50), .Z(n4764) );
  MUX U1792 ( .IN0(n5048), .IN1(n5046), .SEL(n5047), .F(n5042) );
  MUX U1793 ( .IN0(n51), .IN1(n5178), .SEL(n5179), .F(n4078) );
  IV U1794 ( .A(n5180), .Z(n51) );
  MUX U1795 ( .IN0(n52), .IN1(n5263), .SEL(n5264), .F(n4124) );
  IV U1796 ( .A(n5265), .Z(n52) );
  MUX U1797 ( .IN0(n2648), .IN1(n2646), .SEL(n2647), .F(n53) );
  IV U1798 ( .A(n53), .Z(n1783) );
  MUX U1799 ( .IN0(n2706), .IN1(n2704), .SEL(n2705), .F(n54) );
  IV U1800 ( .A(n54), .Z(n1814) );
  MUX U1801 ( .IN0(n2310), .IN1(n2308), .SEL(n2309), .F(n55) );
  IV U1802 ( .A(n55), .Z(n1589) );
  MUX U1803 ( .IN0(n2201), .IN1(n2199), .SEL(n2200), .F(n56) );
  IV U1804 ( .A(n56), .Z(n1522) );
  MUX U1805 ( .IN0(n2423), .IN1(n2421), .SEL(n2422), .F(n57) );
  IV U1806 ( .A(n57), .Z(n1654) );
  MUX U1807 ( .IN0(n6863), .IN1(n6861), .SEL(n6862), .F(n6855) );
  MUX U1808 ( .IN0(n6838), .IN1(n6836), .SEL(n6837), .F(n6832) );
  MUX U1809 ( .IN0(n58), .IN1(n6848), .SEL(n6849), .F(n5020) );
  IV U1810 ( .A(n6850), .Z(n58) );
  MUX U1811 ( .IN0(n6776), .IN1(n6774), .SEL(n6775), .F(n6770) );
  MUX U1812 ( .IN0(n6817), .IN1(n6815), .SEL(n6816), .F(n6811) );
  MUX U1813 ( .IN0(n59), .IN1(n6762), .SEL(n6763), .F(n4969) );
  IV U1814 ( .A(n6764), .Z(n59) );
  MUX U1815 ( .IN0(n6493), .IN1(n6491), .SEL(n6492), .F(n6487) );
  MUX U1816 ( .IN0(n6502), .IN1(n6500), .SEL(n6501), .F(n6494) );
  XOR U1817 ( .A(n6422), .B(n6423), .Z(n4780) );
  XOR U1818 ( .A(n6465), .B(n6466), .Z(n4804) );
  MUX U1819 ( .IN0(n6647), .IN1(n6645), .SEL(n6646), .F(n6639) );
  MUX U1820 ( .IN0(n6150), .IN1(n6148), .SEL(n6149), .F(n6144) );
  MUX U1821 ( .IN0(n6159), .IN1(n6157), .SEL(n6158), .F(n6151) );
  XOR U1822 ( .A(n6122), .B(n6123), .Z(n4612) );
  MUX U1823 ( .IN0(n5984), .IN1(n5982), .SEL(n5983), .F(n5978) );
  MUX U1824 ( .IN0(n6062), .IN1(n6060), .SEL(n6061), .F(n6056) );
  MUX U1825 ( .IN0(n6069), .IN1(n6067), .SEL(n6068), .F(n6063) );
  MUX U1826 ( .IN0(n6268), .IN1(n6266), .SEL(n6267), .F(n6262) );
  MUX U1827 ( .IN0(n6275), .IN1(n6273), .SEL(n6274), .F(n6269) );
  XOR U1828 ( .A(n6199), .B(n6200), .Z(n4652) );
  MUX U1829 ( .IN0(n6324), .IN1(n6322), .SEL(n6323), .F(n6318) );
  MUX U1830 ( .IN0(n6414), .IN1(n6412), .SEL(n6413), .F(n6408) );
  MUX U1831 ( .IN0(n5455), .IN1(n5453), .SEL(n5454), .F(n5449) );
  MUX U1832 ( .IN0(n5462), .IN1(n5460), .SEL(n5461), .F(n5456) );
  MUX U1833 ( .IN0(n5393), .IN1(n5391), .SEL(n5392), .F(n5387) );
  MUX U1834 ( .IN0(n5687), .IN1(n5685), .SEL(n5686), .F(n5681) );
  MUX U1835 ( .IN0(n5696), .IN1(n5694), .SEL(n5695), .F(n5688) );
  MUX U1836 ( .IN0(n5645), .IN1(n5643), .SEL(n5644), .F(n4352) );
  MUX U1837 ( .IN0(n5514), .IN1(n5512), .SEL(n5513), .F(n5508) );
  MUX U1838 ( .IN0(n5521), .IN1(n5519), .SEL(n5520), .F(n5515) );
  MUX U1839 ( .IN0(n5589), .IN1(n5587), .SEL(n5588), .F(n4316) );
  MUX U1840 ( .IN0(n60), .IN1(n5813), .SEL(n5814), .F(n4436) );
  IV U1841 ( .A(n5815), .Z(n60) );
  MUX U1842 ( .IN0(n5856), .IN1(n5854), .SEL(n5855), .F(n61) );
  IV U1843 ( .A(n61), .Z(n4457) );
  MUX U1844 ( .IN0(n5950), .IN1(n5948), .SEL(n5949), .F(n5944) );
  XOR U1845 ( .A(n1679), .B(n1678), .Z(n1672) );
  XOR U1846 ( .A(n1884), .B(n1882), .Z(n1891) );
  XOR U1847 ( .A(n4727), .B(n4725), .Z(n4719) );
  XOR U1848 ( .A(n4518), .B(n4516), .Z(n4508) );
  MUX U1849 ( .IN0(n5920), .IN1(n5922), .SEL(n5921), .F(n62) );
  IV U1850 ( .A(n62), .Z(n4492) );
  XOR U1851 ( .A(n4419), .B(n4417), .Z(n4411) );
  MUX U1852 ( .IN0(n5569), .IN1(n5571), .SEL(n5570), .F(n63) );
  IV U1853 ( .A(n63), .Z(n4296) );
  XOR U1854 ( .A(n4355), .B(n4354), .Z(n4348) );
  XOR U1855 ( .A(n4142), .B(n4141), .Z(n4135) );
  MUX U1856 ( .IN0(n242), .IN1(n4168), .SEL(n4167), .F(n64) );
  IV U1857 ( .A(n64), .Z(n3568) );
  MUX U1858 ( .IN0(n4783), .IN1(n65), .SEL(n4784), .F(n3873) );
  IV U1859 ( .A(n4785), .Z(n65) );
  MUX U1860 ( .IN0(n574), .IN1(n4016), .SEL(n4014), .F(n4009) );
  MUX U1861 ( .IN0(n578), .IN1(n4074), .SEL(n4072), .F(n4067) );
  MUX U1862 ( .IN0(n2637), .IN1(n2635), .SEL(n2636), .F(n2631) );
  MUX U1863 ( .IN0(n2971), .IN1(n2969), .SEL(n2970), .F(n2965) );
  MUX U1864 ( .IN0(n2980), .IN1(n2978), .SEL(n2979), .F(n2972) );
  MUX U1865 ( .IN0(n2936), .IN1(n2934), .SEL(n2935), .F(n66) );
  IV U1866 ( .A(n66), .Z(n1947) );
  MUX U1867 ( .IN0(n2950), .IN1(n2948), .SEL(n2949), .F(n2944) );
  MUX U1868 ( .IN0(n2873), .IN1(n2871), .SEL(n2872), .F(n1921) );
  MUX U1869 ( .IN0(n2894), .IN1(n2892), .SEL(n2893), .F(n2888) );
  MUX U1870 ( .IN0(n2299), .IN1(n2297), .SEL(n2298), .F(n2293) );
  MUX U1871 ( .IN0(n67), .IN1(n2133), .SEL(n2134), .F(n1486) );
  IV U1872 ( .A(n2135), .Z(n67) );
  MUX U1873 ( .IN0(n2484), .IN1(n2482), .SEL(n2483), .F(n2478) );
  MUX U1874 ( .IN0(n594), .IN1(n4989), .SEL(n4987), .F(n4982) );
  MUX U1875 ( .IN0(n397), .IN1(n4999), .SEL(n4997), .F(n4990) );
  MUX U1876 ( .IN0(n599), .IN1(n4965), .SEL(n4963), .F(n4956) );
  MUX U1877 ( .IN0(n608), .IN1(n4900), .SEL(n4898), .F(n4893) );
  MUX U1878 ( .IN0(n90), .IN1(n4593), .SEL(n4592), .F(n68) );
  IV U1879 ( .A(n68), .Z(n3779) );
  MUX U1880 ( .IN0(n614), .IN1(n4529), .SEL(n4527), .F(n4522) );
  MUX U1881 ( .IN0(n619), .IN1(n4665), .SEL(n4663), .F(n4658) );
  MUX U1882 ( .IN0(n631), .IN1(n4208), .SEL(n4206), .F(n4201) );
  MUX U1883 ( .IN0(n408), .IN1(n4218), .SEL(n4216), .F(n4209) );
  MUX U1884 ( .IN0(n500), .IN1(n4320), .SEL(n4318), .F(n3644) );
  MUX U1885 ( .IN0(n648), .IN1(n4433), .SEL(n4431), .F(n4424) );
  MUX U1886 ( .IN0(n501), .IN1(n4415), .SEL(n4413), .F(n4408) );
  XOR U1887 ( .A(n1639), .B(n1638), .Z(n1658) );
  XOR U1888 ( .A(n1868), .B(n1867), .Z(n1887) );
  MUX U1889 ( .IN0(n6335), .IN1(n6337), .SEL(n6336), .F(n69) );
  IV U1890 ( .A(n69), .Z(n4728) );
  MUX U1891 ( .IN0(n342), .IN1(n1810), .SEL(n1809), .F(n70) );
  IV U1892 ( .A(n70), .Z(n1314) );
  XOR U1893 ( .A(n1289), .B(n1287), .Z(n1281) );
  XOR U1894 ( .A(n1227), .B(n1226), .Z(n1220) );
  XOR U1895 ( .A(n1178), .B(n1176), .Z(n1170) );
  XOR U1896 ( .A(n3499), .B(n3498), .Z(n3492) );
  XOR U1897 ( .A(n3938), .B(n3936), .Z(n3945) );
  XOR U1898 ( .A(n3821), .B(n3819), .Z(n3813) );
  MUX U1899 ( .IN0(n3530), .IN1(n3533), .SEL(n3531), .F(n3526) );
  MUX U1900 ( .IN0(n346), .IN1(n1393), .SEL(n1392), .F(n71) );
  IV U1901 ( .A(n71), .Z(n1108) );
  MUX U1902 ( .IN0(n678), .IN1(n1566), .SEL(n1564), .F(n1194) );
  MUX U1903 ( .IN0(n692), .IN1(n1722), .SEL(n1720), .F(n1715) );
  MUX U1904 ( .IN0(n430), .IN1(n3959), .SEL(n3957), .F(n3950) );
  XNOR U1905 ( .A(n3917), .B(n3918), .Z(n3448) );
  MUX U1906 ( .IN0(n3575), .IN1(n3578), .SEL(n3576), .F(n3283) );
  MUX U1907 ( .IN0(n3627), .IN1(n3630), .SEL(n3628), .F(n3623) );
  MUX U1908 ( .IN0(n3637), .IN1(n3640), .SEL(n3638), .F(n3631) );
  MUX U1909 ( .IN0(n3687), .IN1(n3690), .SEL(n3688), .F(n3681) );
  MUX U1910 ( .IN0(n3717), .IN1(n72), .SEL(n3718), .F(n3349) );
  IV U1911 ( .A(n3719), .Z(n72) );
  MUX U1912 ( .IN0(n3734), .IN1(n3737), .SEL(n3735), .F(n3728) );
  MUX U1913 ( .IN0(n2388), .IN1(n2390), .SEL(n2389), .F(n73) );
  IV U1914 ( .A(n73), .Z(n1632) );
  MUX U1915 ( .IN0(n5786), .IN1(n5788), .SEL(n5787), .F(n74) );
  IV U1916 ( .A(n74), .Z(n4420) );
  XOR U1917 ( .A(n3375), .B(n3373), .Z(n3367) );
  MUX U1918 ( .IN0(n2072), .IN1(n2070), .SEL(n2071), .F(n2066) );
  MUX U1919 ( .IN0(n2004), .IN1(n2002), .SEL(n2003), .F(n1998) );
  MUX U1920 ( .IN0(n75), .IN1(n2046), .SEL(n2047), .F(n1436) );
  IV U1921 ( .A(n2048), .Z(n75) );
  MUX U1922 ( .IN0(n3252), .IN1(n3255), .SEL(n3253), .F(n3248) );
  MUX U1923 ( .IN0(n3264), .IN1(n3267), .SEL(n3265), .F(n3129) );
  MUX U1924 ( .IN0(n1187), .IN1(n1190), .SEL(n1188), .F(n1183) );
  MUX U1925 ( .IN0(n1266), .IN1(n1269), .SEL(n1267), .F(n1262) );
  MUX U1926 ( .IN0(n354), .IN1(n3447), .SEL(n3445), .F(n3438) );
  MUX U1927 ( .IN0(n3276), .IN1(n3279), .SEL(n3277), .F(n3272) );
  MUX U1928 ( .IN0(n368), .IN1(n4584), .SEL(n4583), .F(n76) );
  IV U1929 ( .A(n76), .Z(n3774) );
  XOR U1930 ( .A(n989), .B(n988), .Z(n1008) );
  XOR U1931 ( .A(n951), .B(n950), .Z(n960) );
  MUX U1932 ( .IN0(n3315), .IN1(n77), .SEL(n3316), .F(n3154) );
  IV U1933 ( .A(n3317), .Z(n77) );
  MUX U1934 ( .IN0(n763), .IN1(n1447), .SEL(n1445), .F(n1440) );
  MUX U1935 ( .IN0(n765), .IN1(n1422), .SEL(n1420), .F(n1415) );
  MUX U1936 ( .IN0(n766), .IN1(n1432), .SEL(n1430), .F(n1423) );
  MUX U1937 ( .IN0(n1075), .IN1(n1078), .SEL(n1076), .F(n944) );
  MUX U1938 ( .IN0(n1038), .IN1(n1041), .SEL(n1039), .F(n1034) );
  MUX U1939 ( .IN0(n3213), .IN1(n3216), .SEL(n3214), .F(n3207) );
  MUX U1940 ( .IN0(n3202), .IN1(n3205), .SEL(n3203), .F(n3100) );
  MUX U1941 ( .IN0(n3161), .IN1(n3164), .SEL(n3162), .F(n3157) );
  MUX U1942 ( .IN0(n937), .IN1(n940), .SEL(n938), .F(n933) );
  MUX U1943 ( .IN0(n922), .IN1(n925), .SEL(n923), .F(n918) );
  MUX U1944 ( .IN0(n3093), .IN1(n3096), .SEL(n3094), .F(n3089) );
  MUX U1945 ( .IN0(n3084), .IN1(n3087), .SEL(n3085), .F(n3045) );
  MUX U1946 ( .IN0(n3038), .IN1(n3041), .SEL(n3039), .F(n3033) );
  MUX U1947 ( .IN0(n6662), .IN1(n6660), .SEL(n6661), .F(n78) );
  IV U1948 ( .A(n78), .Z(n4910) );
  MUX U1949 ( .IN0(n5135), .IN1(n5133), .SEL(n5134), .F(n5127) );
  MUX U1950 ( .IN0(n5110), .IN1(n5108), .SEL(n5109), .F(n5104) );
  MUX U1951 ( .IN0(n5119), .IN1(n5117), .SEL(n5118), .F(n5111) );
  MUX U1952 ( .IN0(n5089), .IN1(n5087), .SEL(n5088), .F(n5083) );
  MUX U1953 ( .IN0(n2595), .IN1(n2593), .SEL(n2594), .F(n79) );
  IV U1954 ( .A(n79), .Z(n1750) );
  MUX U1955 ( .IN0(n2143), .IN1(n2141), .SEL(n2142), .F(n80) );
  IV U1956 ( .A(n80), .Z(n1493) );
  MUX U1957 ( .IN0(n81), .IN1(n6777), .SEL(n6778), .F(n4978) );
  IV U1958 ( .A(n6779), .Z(n81) );
  MUX U1959 ( .IN0(n82), .IN1(n6818), .SEL(n6819), .F(n5003) );
  IV U1960 ( .A(n6820), .Z(n82) );
  MUX U1961 ( .IN0(n6692), .IN1(n6690), .SEL(n6691), .F(n6684) );
  MUX U1962 ( .IN0(n6747), .IN1(n6745), .SEL(n6746), .F(n83) );
  IV U1963 ( .A(n83), .Z(n4957) );
  MUX U1964 ( .IN0(n6518), .IN1(n6516), .SEL(n6517), .F(n6510) );
  MUX U1965 ( .IN0(n84), .IN1(n6503), .SEL(n6504), .F(n4823) );
  IV U1966 ( .A(n6505), .Z(n84) );
  MUX U1967 ( .IN0(n6429), .IN1(n6427), .SEL(n6428), .F(n6421) );
  MUX U1968 ( .IN0(n85), .IN1(n6473), .SEL(n6474), .F(n4806) );
  IV U1969 ( .A(n6475), .Z(n85) );
  MUX U1970 ( .IN0(n6576), .IN1(n6574), .SEL(n6575), .F(n6570) );
  MUX U1971 ( .IN0(n6543), .IN1(n6541), .SEL(n6542), .F(n4852) );
  XOR U1972 ( .A(n6555), .B(n6556), .Z(n4853) );
  XOR U1973 ( .A(n6168), .B(n6169), .Z(n4636) );
  XOR U1974 ( .A(n6152), .B(n6153), .Z(n4629) );
  MUX U1975 ( .IN0(n6084), .IN1(n6082), .SEL(n6083), .F(n6078) );
  MUX U1976 ( .IN0(n6129), .IN1(n6127), .SEL(n6128), .F(n6121) );
  MUX U1977 ( .IN0(n5977), .IN1(n5975), .SEL(n5976), .F(n5971) );
  MUX U1978 ( .IN0(n6289), .IN1(n6287), .SEL(n6288), .F(n6283) );
  MUX U1979 ( .IN0(n86), .IN1(n6276), .SEL(n6277), .F(n4695) );
  IV U1980 ( .A(n6278), .Z(n86) );
  MUX U1981 ( .IN0(n6345), .IN1(n6343), .SEL(n6344), .F(n6339) );
  MUX U1982 ( .IN0(n87), .IN1(n6332), .SEL(n6333), .F(n4727) );
  IV U1983 ( .A(n6334), .Z(n87) );
  MUX U1984 ( .IN0(n6373), .IN1(n6371), .SEL(n6372), .F(n6367) );
  MUX U1985 ( .IN0(n5478), .IN1(n5476), .SEL(n5477), .F(n5470) );
  MUX U1986 ( .IN0(n88), .IN1(n5463), .SEL(n5464), .F(n4240) );
  IV U1987 ( .A(n5465), .Z(n88) );
  MUX U1988 ( .IN0(n5417), .IN1(n5415), .SEL(n5416), .F(n4218) );
  MUX U1989 ( .IN0(n5309), .IN1(n5307), .SEL(n5308), .F(n5301) );
  MUX U1990 ( .IN0(n5274), .IN1(n5272), .SEL(n5273), .F(n4139) );
  XOR U1991 ( .A(n5286), .B(n5287), .Z(n4140) );
  MUX U1992 ( .IN0(n5337), .IN1(n5335), .SEL(n5336), .F(n5331) );
  MUX U1993 ( .IN0(n5371), .IN1(n5369), .SEL(n5370), .F(n5365) );
  XOR U1994 ( .A(n5705), .B(n5706), .Z(n4377) );
  XOR U1995 ( .A(n5689), .B(n5690), .Z(n4370) );
  MUX U1996 ( .IN0(n5621), .IN1(n5619), .SEL(n5620), .F(n5615) );
  MUX U1997 ( .IN0(n5666), .IN1(n5664), .SEL(n5665), .F(n5658) );
  MUX U1998 ( .IN0(n5565), .IN1(n5563), .SEL(n5564), .F(n5559) );
  MUX U1999 ( .IN0(n5828), .IN1(n5826), .SEL(n5827), .F(n5820) );
  XOR U2000 ( .A(n5865), .B(n5866), .Z(n4466) );
  MUX U2001 ( .IN0(n2516), .IN1(n2518), .SEL(n2517), .F(n89) );
  IV U2002 ( .A(n89), .Z(n1703) );
  XOR U2003 ( .A(n1980), .B(n1979), .Z(n1987) );
  XOR U2004 ( .A(n1815), .B(n1813), .Z(n1822) );
  XOR U2005 ( .A(n1784), .B(n1782), .Z(n1791) );
  MUX U2006 ( .IN0(n6088), .IN1(n6090), .SEL(n6089), .F(n90) );
  IV U2007 ( .A(n90), .Z(n4591) );
  XOR U2008 ( .A(n4491), .B(n4489), .Z(n4498) );
  MUX U2009 ( .IN0(n5625), .IN1(n5627), .SEL(n5626), .F(n91) );
  IV U2010 ( .A(n91), .Z(n4332) );
  XOR U2011 ( .A(n4197), .B(n4195), .Z(n4204) );
  MUX U2012 ( .IN0(n5052), .IN1(n5054), .SEL(n5053), .F(n92) );
  IV U2013 ( .A(n92), .Z(n4006) );
  MUX U2014 ( .IN0(n319), .IN1(n4382), .SEL(n4381), .F(n93) );
  IV U2015 ( .A(n93), .Z(n3673) );
  MUX U2016 ( .IN0(n240), .IN1(n5029), .SEL(n5028), .F(n94) );
  IV U2017 ( .A(n94), .Z(n3991) );
  MUX U2018 ( .IN0(n317), .IN1(n4641), .SEL(n4640), .F(n95) );
  IV U2019 ( .A(n95), .Z(n3802) );
  MUX U2020 ( .IN0(n657), .IN1(n4559), .SEL(n4558), .F(n96) );
  IV U2021 ( .A(n96), .Z(n3763) );
  MUX U2022 ( .IN0(n575), .IN1(n4005), .SEL(n4003), .F(n3496) );
  XNOR U2023 ( .A(n4018), .B(n4019), .Z(n3497) );
  MUX U2024 ( .IN0(n509), .IN1(n4104), .SEL(n4103), .F(n97) );
  IV U2025 ( .A(n97), .Z(n3535) );
  MUX U2026 ( .IN0(n98), .IN1(n2638), .SEL(n2639), .F(n1776) );
  IV U2027 ( .A(n2640), .Z(n98) );
  MUX U2028 ( .IN0(n2568), .IN1(n2566), .SEL(n2567), .F(n2562) );
  MUX U2029 ( .IN0(n2695), .IN1(n2693), .SEL(n2694), .F(n2687) );
  MUX U2030 ( .IN0(n2961), .IN1(n2959), .SEL(n2960), .F(n1971) );
  MUX U2031 ( .IN0(n99), .IN1(n2981), .SEL(n2982), .F(n1974) );
  IV U2032 ( .A(n2983), .Z(n99) );
  MUX U2033 ( .IN0(n2909), .IN1(n2907), .SEL(n2908), .F(n2903) );
  MUX U2034 ( .IN0(n2821), .IN1(n2819), .SEL(n2820), .F(n2815) );
  MUX U2035 ( .IN0(n2790), .IN1(n2788), .SEL(n2789), .F(n1872) );
  MUX U2036 ( .IN0(n2807), .IN1(n2805), .SEL(n2806), .F(n2801) );
  MUX U2037 ( .IN0(n2849), .IN1(n2847), .SEL(n2848), .F(n2843) );
  MUX U2038 ( .IN0(n2333), .IN1(n2331), .SEL(n2332), .F(n2327) );
  MUX U2039 ( .IN0(n2313), .IN1(n2311), .SEL(n2312), .F(n2307) );
  MUX U2040 ( .IN0(n2174), .IN1(n2172), .SEL(n2173), .F(n2168) );
  MUX U2041 ( .IN0(n2426), .IN1(n2424), .SEL(n2425), .F(n2420) );
  XOR U2042 ( .A(n1663), .B(n683), .Z(n2433) );
  MUX U2043 ( .IN0(n2504), .IN1(n2502), .SEL(n2503), .F(n2498) );
  MUX U2044 ( .IN0(n100), .IN1(n2485), .SEL(n2486), .F(n1687) );
  IV U2045 ( .A(n2487), .Z(n100) );
  MUX U2046 ( .IN0(n2454), .IN1(n2452), .SEL(n2453), .F(n101) );
  IV U2047 ( .A(n101), .Z(n1668) );
  MUX U2048 ( .IN0(n2553), .IN1(n2551), .SEL(n2552), .F(n2547) );
  XNOR U2049 ( .A(n5009), .B(n5010), .Z(n3984) );
  XNOR U2050 ( .A(n4991), .B(n4992), .Z(n3977) );
  MUX U2051 ( .IN0(n476), .IN1(n4969), .SEL(n4967), .F(n3962) );
  MUX U2052 ( .IN0(n601), .IN1(n4820), .SEL(n4818), .F(n4811) );
  MUX U2053 ( .IN0(n602), .IN1(n4793), .SEL(n4791), .F(n4786) );
  MUX U2054 ( .IN0(n603), .IN1(n4803), .SEL(n4801), .F(n4794) );
  MUX U2055 ( .IN0(n4901), .IN1(n4903), .SEL(n4902), .F(n3929) );
  MUX U2056 ( .IN0(n610), .IN1(n4628), .SEL(n4626), .F(n4619) );
  MUX U2057 ( .IN0(n611), .IN1(n4601), .SEL(n4599), .F(n4594) );
  MUX U2058 ( .IN0(n138), .IN1(n4611), .SEL(n4609), .F(n4602) );
  MUX U2059 ( .IN0(n299), .IN1(n4533), .SEL(n4531), .F(n3748) );
  MUX U2060 ( .IN0(n618), .IN1(n4691), .SEL(n4689), .F(n4682) );
  MUX U2061 ( .IN0(n231), .IN1(n4677), .SEL(n4675), .F(n3821) );
  MUX U2062 ( .IN0(n623), .IN1(n4723), .SEL(n4721), .F(n4716) );
  MUX U2063 ( .IN0(n625), .IN1(n4762), .SEL(n4760), .F(n4755) );
  MUX U2064 ( .IN0(n630), .IN1(n4236), .SEL(n4234), .F(n4227) );
  MUX U2065 ( .IN0(n305), .IN1(n4222), .SEL(n4220), .F(n3595) );
  MUX U2066 ( .IN0(n635), .IN1(n4176), .SEL(n4174), .F(n4169) );
  MUX U2067 ( .IN0(n494), .IN1(n4188), .SEL(n4186), .F(n3578) );
  MUX U2068 ( .IN0(n639), .IN1(n4369), .SEL(n4367), .F(n4360) );
  MUX U2069 ( .IN0(n640), .IN1(n4342), .SEL(n4340), .F(n4335) );
  MUX U2070 ( .IN0(n142), .IN1(n4352), .SEL(n4350), .F(n4343) );
  MUX U2071 ( .IN0(n649), .IN1(n4407), .SEL(n4405), .F(n4400) );
  XNOR U2072 ( .A(n4457), .B(n4458), .Z(n3714) );
  XOR U2073 ( .A(n1558), .B(n1557), .Z(n1546) );
  XOR U2074 ( .A(n1917), .B(n1916), .Z(n1903) );
  XOR U2075 ( .A(n1951), .B(n1950), .Z(n1937) );
  MUX U2076 ( .IN0(n5988), .IN1(n5990), .SEL(n5989), .F(n102) );
  IV U2077 ( .A(n102), .Z(n4534) );
  MUX U2078 ( .IN0(n6506), .IN1(n6508), .SEL(n6507), .F(n103) );
  IV U2079 ( .A(n103), .Z(n4824) );
  XOR U2080 ( .A(n4429), .B(n4428), .Z(n4446) );
  MUX U2081 ( .IN0(n5181), .IN1(n5183), .SEL(n5182), .F(n104) );
  IV U2082 ( .A(n104), .Z(n4079) );
  XOR U2083 ( .A(n1235), .B(n1233), .Z(n1242) );
  XOR U2084 ( .A(n1194), .B(n1192), .Z(n1186) );
  XOR U2085 ( .A(n1202), .B(n1200), .Z(n1209) );
  MUX U2086 ( .IN0(n535), .IN1(n1489), .SEL(n1488), .F(n105) );
  IV U2087 ( .A(n105), .Z(n1156) );
  MUX U2088 ( .IN0(n167), .IN1(n4275), .SEL(n4274), .F(n106) );
  IV U2089 ( .A(n106), .Z(n3620) );
  MUX U2090 ( .IN0(n168), .IN1(n4145), .SEL(n4144), .F(n107) );
  IV U2091 ( .A(n107), .Z(n3556) );
  MUX U2092 ( .IN0(n4728), .IN1(n108), .SEL(n4729), .F(n3845) );
  IV U2093 ( .A(n4730), .Z(n108) );
  MUX U2094 ( .IN0(n348), .IN1(n3989), .SEL(n3988), .F(n109) );
  IV U2095 ( .A(n109), .Z(n3477) );
  MUX U2096 ( .IN0(n3519), .IN1(n3522), .SEL(n3520), .F(n3263) );
  MUX U2097 ( .IN0(n583), .IN1(n1772), .SEL(n1770), .F(n1765) );
  MUX U2098 ( .IN0(n588), .IN1(n1804), .SEL(n1802), .F(n1797) );
  MUX U2099 ( .IN0(n655), .IN1(n1834), .SEL(n1833), .F(n110) );
  IV U2100 ( .A(n110), .Z(n1326) );
  XNOR U2101 ( .A(n1845), .B(n1846), .Z(n1333) );
  MUX U2102 ( .IN0(n665), .IN1(n1945), .SEL(n1943), .F(n1938) );
  XNOR U2103 ( .A(n1947), .B(n1948), .Z(n1380) );
  MUX U2104 ( .IN0(n667), .IN1(n1895), .SEL(n1893), .F(n1888) );
  MUX U2105 ( .IN0(n520), .IN1(n1520), .SEL(n1518), .F(n1514) );
  XNOR U2106 ( .A(n1619), .B(n1620), .Z(n1225) );
  XNOR U2107 ( .A(n3968), .B(n3969), .Z(n3470) );
  XNOR U2108 ( .A(n3951), .B(n3952), .Z(n3463) );
  MUX U2109 ( .IN0(n3922), .IN1(n3925), .SEL(n3923), .F(n3916) );
  MUX U2110 ( .IN0(n3814), .IN1(n3817), .SEL(n3815), .F(n3810) );
  MUX U2111 ( .IN0(n3866), .IN1(n3869), .SEL(n3867), .F(n3420) );
  XNOR U2112 ( .A(n3584), .B(n3585), .Z(n3288) );
  MUX U2113 ( .IN0(n3616), .IN1(n3619), .SEL(n3617), .F(n3310) );
  MUX U2114 ( .IN0(n164), .IN1(n3694), .SEL(n3692), .F(n3336) );
  MUX U2115 ( .IN0(n3724), .IN1(n3727), .SEL(n3725), .F(n3720) );
  MUX U2116 ( .IN0(n3738), .IN1(n3741), .SEL(n3739), .F(n3361) );
  MUX U2117 ( .IN0(n2275), .IN1(n2277), .SEL(n2276), .F(n111) );
  IV U2118 ( .A(n111), .Z(n1567) );
  MUX U2119 ( .IN0(n2613), .IN1(n2615), .SEL(n2614), .F(n112) );
  IV U2120 ( .A(n112), .Z(n1761) );
  MUX U2121 ( .IN0(n4420), .IN1(n113), .SEL(n4421), .F(n3695) );
  IV U2122 ( .A(n4422), .Z(n113) );
  MUX U2123 ( .IN0(n2065), .IN1(n2063), .SEL(n2064), .F(n2059) );
  MUX U2124 ( .IN0(n114), .IN1(n2073), .SEL(n2074), .F(n1451) );
  IV U2125 ( .A(n2075), .Z(n114) );
  MUX U2126 ( .IN0(n1228), .IN1(n115), .SEL(n1229), .F(n1021) );
  IV U2127 ( .A(n1230), .Z(n115) );
  MUX U2128 ( .IN0(n3883), .IN1(n116), .SEL(n3884), .F(n3427) );
  IV U2129 ( .A(n3885), .Z(n116) );
  XOR U2130 ( .A(n3314), .B(n3312), .Z(n3306) );
  XOR U2131 ( .A(n3267), .B(n3265), .Z(n3259) );
  MUX U2132 ( .IN0(n3500), .IN1(n117), .SEL(n3501), .F(n3245) );
  IV U2133 ( .A(n3502), .Z(n117) );
  MUX U2134 ( .IN0(n3291), .IN1(n118), .SEL(n3292), .F(n3142) );
  IV U2135 ( .A(n3293), .Z(n118) );
  MUX U2136 ( .IN0(n3473), .IN1(n119), .SEL(n3474), .F(n3232) );
  IV U2137 ( .A(n3475), .Z(n119) );
  MUX U2138 ( .IN0(n2101), .IN1(n2099), .SEL(n2100), .F(n120) );
  IV U2139 ( .A(n120), .Z(n1463) );
  MUX U2140 ( .IN0(n1344), .IN1(n121), .SEL(n1345), .F(n1084) );
  IV U2141 ( .A(n1346), .Z(n121) );
  MUX U2142 ( .IN0(n1175), .IN1(n1178), .SEL(n1176), .F(n997) );
  MUX U2143 ( .IN0(n1221), .IN1(n1224), .SEL(n1222), .F(n1215) );
  MUX U2144 ( .IN0(n3459), .IN1(n3462), .SEL(n3460), .F(n3455) );
  XOR U2145 ( .A(n1436), .B(n1434), .Z(n1428) );
  MUX U2146 ( .IN0(n3774), .IN1(n122), .SEL(n3775), .F(n3376) );
  IV U2147 ( .A(n3776), .Z(n122) );
  MUX U2148 ( .IN0(n3138), .IN1(n123), .SEL(n3139), .F(n3069) );
  IV U2149 ( .A(n3140), .Z(n123) );
  MUX U2150 ( .IN0(n1050), .IN1(n1053), .SEL(n1051), .F(n940) );
  MUX U2151 ( .IN0(n1104), .IN1(n124), .SEL(n1105), .F(n956) );
  IV U2152 ( .A(n1106), .Z(n124) );
  MUX U2153 ( .IN0(n990), .IN1(n993), .SEL(n991), .F(n986) );
  MUX U2154 ( .IN0(n3179), .IN1(n3182), .SEL(n3180), .F(n3096) );
  MUX U2155 ( .IN0(n3077), .IN1(n125), .SEL(n3078), .F(n3044) );
  IV U2156 ( .A(n3079), .Z(n125) );
  MUX U2157 ( .IN0(n375), .IN1(n4127), .SEL(n4126), .F(n126) );
  IV U2158 ( .A(n126), .Z(n3548) );
  MUX U2159 ( .IN0(n1336), .IN1(n127), .SEL(n1337), .F(n1079) );
  IV U2160 ( .A(n1338), .Z(n127) );
  MUX U2161 ( .IN0(n1122), .IN1(n128), .SEL(n1123), .F(n970) );
  IV U2162 ( .A(n1124), .Z(n128) );
  MUX U2163 ( .IN0(n3220), .IN1(n129), .SEL(n3221), .F(n3105) );
  IV U2164 ( .A(n3222), .Z(n129) );
  MUX U2165 ( .IN0(n941), .IN1(n944), .SEL(n942), .F(n878) );
  MUX U2166 ( .IN0(n914), .IN1(n917), .SEL(n915), .F(n910) );
  MUX U2167 ( .IN0(n926), .IN1(n929), .SEL(n927), .F(n870) );
  MUX U2168 ( .IN0(n3097), .IN1(n3100), .SEL(n3098), .F(n3050) );
  MUX U2169 ( .IN0(n3484), .IN1(n130), .SEL(n1118), .F(n3239) );
  IV U2170 ( .A(n1117), .Z(n130) );
  MUX U2171 ( .IN0(n280), .IN1(n983), .SEL(n981), .F(n975) );
  MUX U2172 ( .IN0(n3055), .IN1(n3058), .SEL(n3056), .F(n3051) );
  MUX U2173 ( .IN0(n3035), .IN1(n131), .SEL(n3036), .F(n3024) );
  IV U2174 ( .A(n3037), .Z(n131) );
  MUX U2175 ( .IN0(n804), .IN1(n831), .SEL(n803), .F(n820) );
  MUX U2176 ( .IN0(n5841), .IN1(n5839), .SEL(n5840), .F(n132) );
  IV U2177 ( .A(n132), .Z(n4448) );
  MUX U2178 ( .IN0(n5155), .IN1(n5153), .SEL(n5154), .F(n5149) );
  MUX U2179 ( .IN0(n133), .IN1(n5120), .SEL(n5121), .F(n4047) );
  IV U2180 ( .A(n5122), .Z(n133) );
  MUX U2181 ( .IN0(n134), .IN1(n5090), .SEL(n5091), .F(n4030) );
  IV U2182 ( .A(n5092), .Z(n134) );
  XOR U2183 ( .A(n5186), .B(n5187), .Z(n4083) );
  MUX U2184 ( .IN0(n5221), .IN1(n5219), .SEL(n5220), .F(n5215) );
  MUX U2185 ( .IN0(n2623), .IN1(n2621), .SEL(n2622), .F(n135) );
  IV U2186 ( .A(n135), .Z(n1766) );
  MUX U2187 ( .IN0(n2118), .IN1(n2116), .SEL(n2117), .F(n136) );
  IV U2188 ( .A(n136), .Z(n1476) );
  MUX U2189 ( .IN0(n6883), .IN1(n6881), .SEL(n6882), .F(n6877) );
  XOR U2190 ( .A(n6856), .B(n6857), .Z(n5024) );
  XOR U2191 ( .A(n6840), .B(n6841), .Z(n5018) );
  MUX U2192 ( .IN0(n6810), .IN1(n6808), .SEL(n6809), .F(n6804) );
  MUX U2193 ( .IN0(n6712), .IN1(n6710), .SEL(n6711), .F(n6706) );
  MUX U2194 ( .IN0(n6659), .IN1(n6657), .SEL(n6658), .F(n4916) );
  MUX U2195 ( .IN0(n6740), .IN1(n6738), .SEL(n6739), .F(n6734) );
  MUX U2196 ( .IN0(n6720), .IN1(n6718), .SEL(n6719), .F(n6714) );
  MUX U2197 ( .IN0(n6754), .IN1(n6752), .SEL(n6753), .F(n6748) );
  MUX U2198 ( .IN0(n6538), .IN1(n6536), .SEL(n6537), .F(n6532) );
  MUX U2199 ( .IN0(n6463), .IN1(n6461), .SEL(n6462), .F(n6457) );
  MUX U2200 ( .IN0(n137), .IN1(n6577), .SEL(n6578), .F(n4863) );
  IV U2201 ( .A(n6579), .Z(n137) );
  MUX U2202 ( .IN0(n6562), .IN1(n6560), .SEL(n6561), .F(n6554) );
  MUX U2203 ( .IN0(n6604), .IN1(n6602), .SEL(n6603), .F(n6598) );
  MUX U2204 ( .IN0(n6195), .IN1(n6193), .SEL(n6194), .F(n6189) );
  MUX U2205 ( .IN0(n6175), .IN1(n6173), .SEL(n6174), .F(n6167) );
  MUX U2206 ( .IN0(n6117), .IN1(n6115), .SEL(n6116), .F(n138) );
  IV U2207 ( .A(n138), .Z(n4610) );
  XOR U2208 ( .A(n5993), .B(n5994), .Z(n4538) );
  MUX U2209 ( .IN0(n6028), .IN1(n6026), .SEL(n6027), .F(n6022) );
  MUX U2210 ( .IN0(n139), .IN1(n6290), .SEL(n6291), .F(n4703) );
  IV U2211 ( .A(n6292), .Z(n139) );
  MUX U2212 ( .IN0(n6314), .IN1(n6312), .SEL(n6313), .F(n4723) );
  MUX U2213 ( .IN0(n140), .IN1(n6374), .SEL(n6375), .F(n4751) );
  IV U2214 ( .A(n6376), .Z(n140) );
  MUX U2215 ( .IN0(n141), .IN1(n6415), .SEL(n6416), .F(n4776) );
  IV U2216 ( .A(n6417), .Z(n141) );
  MUX U2217 ( .IN0(n5498), .IN1(n5496), .SEL(n5497), .F(n5492) );
  XOR U2218 ( .A(n5471), .B(n5472), .Z(n4245) );
  MUX U2219 ( .IN0(n5434), .IN1(n5432), .SEL(n5433), .F(n5428) );
  MUX U2220 ( .IN0(n5329), .IN1(n5327), .SEL(n5328), .F(n5323) );
  MUX U2221 ( .IN0(n5732), .IN1(n5730), .SEL(n5731), .F(n5726) );
  MUX U2222 ( .IN0(n5712), .IN1(n5710), .SEL(n5711), .F(n5704) );
  MUX U2223 ( .IN0(n5654), .IN1(n5652), .SEL(n5653), .F(n142) );
  IV U2224 ( .A(n142), .Z(n4351) );
  MUX U2225 ( .IN0(n5537), .IN1(n5535), .SEL(n5536), .F(n5529) );
  MUX U2226 ( .IN0(n5504), .IN1(n5502), .SEL(n5503), .F(n4268) );
  MUX U2227 ( .IN0(n143), .IN1(n5566), .SEL(n5567), .F(n4295) );
  IV U2228 ( .A(n5568), .Z(n143) );
  XOR U2229 ( .A(n5821), .B(n5822), .Z(n4441) );
  XOR U2230 ( .A(n5805), .B(n5806), .Z(n4434) );
  MUX U2231 ( .IN0(n5741), .IN1(n5739), .SEL(n5740), .F(n5735) );
  MUX U2232 ( .IN0(n5888), .IN1(n5886), .SEL(n5887), .F(n5880) );
  MUX U2233 ( .IN0(n5872), .IN1(n5870), .SEL(n5871), .F(n5864) );
  MUX U2234 ( .IN0(n144), .IN1(n5917), .SEL(n5918), .F(n4491) );
  IV U2235 ( .A(n5919), .Z(n144) );
  MUX U2236 ( .IN0(n5940), .IN1(n5938), .SEL(n5939), .F(n4514) );
  MUX U2237 ( .IN0(n145), .IN1(n5958), .SEL(n5959), .F(n4518) );
  IV U2238 ( .A(n5960), .Z(n145) );
  XOR U2239 ( .A(n1726), .B(n1724), .Z(n1718) );
  MUX U2240 ( .IN0(n2178), .IN1(n2180), .SEL(n2179), .F(n146) );
  IV U2241 ( .A(n146), .Z(n1511) );
  XOR U2242 ( .A(n1974), .B(n1973), .Z(n1967) );
  MUX U2243 ( .IN0(n2913), .IN1(n2915), .SEL(n2914), .F(n147) );
  IV U2244 ( .A(n147), .Z(n1935) );
  XOR U2245 ( .A(n1857), .B(n1855), .Z(n1849) );
  MUX U2246 ( .IN0(n6210), .IN1(n6212), .SEL(n6211), .F(n148) );
  IV U2247 ( .A(n148), .Z(n4655) );
  XOR U2248 ( .A(n4969), .B(n4967), .Z(n4961) );
  MUX U2249 ( .IN0(n6724), .IN1(n6726), .SEL(n6725), .F(n149) );
  IV U2250 ( .A(n149), .Z(n4944) );
  XOR U2251 ( .A(n4920), .B(n4918), .Z(n4912) );
  XOR U2252 ( .A(n4927), .B(n4926), .Z(n4934) );
  MUX U2253 ( .IN0(n6780), .IN1(n6782), .SEL(n6781), .F(n150) );
  IV U2254 ( .A(n150), .Z(n4979) );
  XOR U2255 ( .A(n4830), .B(n4829), .Z(n4837) );
  XOR U2256 ( .A(n4272), .B(n4270), .Z(n4264) );
  XOR U2257 ( .A(n4149), .B(n4148), .Z(n4156) );
  XOR U2258 ( .A(n4054), .B(n4053), .Z(n4061) );
  MUX U2259 ( .IN0(n508), .IN1(n4446), .SEL(n4445), .F(n151) );
  IV U2260 ( .A(n151), .Z(n3706) );
  MUX U2261 ( .IN0(n420), .IN1(n4250), .SEL(n4249), .F(n152) );
  IV U2262 ( .A(n152), .Z(n3607) );
  MUX U2263 ( .IN0(n573), .IN1(n4044), .SEL(n4042), .F(n4035) );
  MUX U2264 ( .IN0(n576), .IN1(n4026), .SEL(n4024), .F(n4017) );
  MUX U2265 ( .IN0(n510), .IN1(n4088), .SEL(n4087), .F(n153) );
  IV U2266 ( .A(n153), .Z(n3527) );
  MUX U2267 ( .IN0(n2671), .IN1(n2669), .SEL(n2670), .F(n2665) );
  MUX U2268 ( .IN0(n2651), .IN1(n2649), .SEL(n2650), .F(n2645) );
  MUX U2269 ( .IN0(n2609), .IN1(n2607), .SEL(n2608), .F(n2603) );
  MUX U2270 ( .IN0(n2729), .IN1(n2727), .SEL(n2728), .F(n2723) );
  MUX U2271 ( .IN0(n2709), .IN1(n2707), .SEL(n2708), .F(n2703) );
  MUX U2272 ( .IN0(n2686), .IN1(n2684), .SEL(n2685), .F(n2680) );
  MUX U2273 ( .IN0(n154), .IN1(n2696), .SEL(n2697), .F(n1807) );
  IV U2274 ( .A(n2698), .Z(n154) );
  MUX U2275 ( .IN0(n2761), .IN1(n2759), .SEL(n2760), .F(n1853) );
  MUX U2276 ( .IN0(n3016), .IN1(n3014), .SEL(n3015), .F(n3010) );
  MUX U2277 ( .IN0(n2996), .IN1(n2994), .SEL(n2995), .F(n2988) );
  MUX U2278 ( .IN0(n155), .IN1(n2951), .SEL(n2952), .F(n1959) );
  IV U2279 ( .A(n2953), .Z(n155) );
  MUX U2280 ( .IN0(n2853), .IN1(n2855), .SEL(n2854), .F(n156) );
  IV U2281 ( .A(n156), .Z(n1901) );
  MUX U2282 ( .IN0(n157), .IN1(n2850), .SEL(n2851), .F(n1900) );
  IV U2283 ( .A(n2852), .Z(n157) );
  MUX U2284 ( .IN0(n158), .IN1(n2314), .SEL(n2315), .F(n1590) );
  IV U2285 ( .A(n2316), .Z(n158) );
  MUX U2286 ( .IN0(n159), .IN1(n2300), .SEL(n2301), .F(n1582) );
  IV U2287 ( .A(n2302), .Z(n159) );
  MUX U2288 ( .IN0(n2230), .IN1(n2228), .SEL(n2229), .F(n2224) );
  MUX U2289 ( .IN0(n2146), .IN1(n2144), .SEL(n2145), .F(n2140) );
  XOR U2290 ( .A(n1534), .B(n1532), .Z(n1524) );
  MUX U2291 ( .IN0(n160), .IN1(n2427), .SEL(n2428), .F(n1655) );
  IV U2292 ( .A(n2429), .Z(n160) );
  MUX U2293 ( .IN0(n161), .IN1(n2413), .SEL(n2414), .F(n1647) );
  IV U2294 ( .A(n2415), .Z(n161) );
  XOR U2295 ( .A(n1687), .B(n1685), .Z(n1693) );
  MUX U2296 ( .IN0(n2461), .IN1(n2459), .SEL(n2460), .F(n2455) );
  MUX U2297 ( .IN0(n2470), .IN1(n2468), .SEL(n2469), .F(n2462) );
  XOR U2298 ( .A(n1702), .B(n1700), .Z(n1709) );
  MUX U2299 ( .IN0(n593), .IN1(n5017), .SEL(n5015), .F(n5008) );
  MUX U2300 ( .IN0(n398), .IN1(n5003), .SEL(n5001), .F(n3979) );
  MUX U2301 ( .IN0(n4804), .IN1(n4806), .SEL(n4805), .F(n3882) );
  MUX U2302 ( .IN0(n604), .IN1(n4874), .SEL(n4872), .F(n4867) );
  XNOR U2303 ( .A(n4844), .B(n4845), .Z(n3902) );
  MUX U2304 ( .IN0(n4612), .IN1(n4614), .SEL(n4613), .F(n3790) );
  MUX U2305 ( .IN0(n416), .IN1(n4543), .SEL(n4542), .F(n162) );
  IV U2306 ( .A(n162), .Z(n3755) );
  MUX U2307 ( .IN0(n615), .IN1(n4567), .SEL(n4565), .F(n4560) );
  MUX U2308 ( .IN0(n617), .IN1(n4714), .SEL(n4712), .F(n4707) );
  MUX U2309 ( .IN0(n4652), .IN1(n4654), .SEL(n4653), .F(n3817) );
  MUX U2310 ( .IN0(n624), .IN1(n4727), .SEL(n4725), .F(n3844) );
  XNOR U2311 ( .A(n4228), .B(n4229), .Z(n3600) );
  XNOR U2312 ( .A(n4210), .B(n4211), .Z(n3593) );
  MUX U2313 ( .IN0(n3568), .IN1(n163), .SEL(n3569), .F(n3282) );
  IV U2314 ( .A(n3570), .Z(n163) );
  MUX U2315 ( .IN0(n4353), .IN1(n4355), .SEL(n4354), .F(n3661) );
  MUX U2316 ( .IN0(n644), .IN1(n4306), .SEL(n4304), .F(n4299) );
  XNOR U2317 ( .A(n4425), .B(n4426), .Z(n3699) );
  MUX U2318 ( .IN0(n412), .IN1(n4411), .SEL(n4410), .F(n164) );
  IV U2319 ( .A(n164), .Z(n3693) );
  MUX U2320 ( .IN0(n652), .IN1(n4465), .SEL(n4463), .F(n4456) );
  MUX U2321 ( .IN0(n2641), .IN1(n2643), .SEL(n2642), .F(n165) );
  IV U2322 ( .A(n165), .Z(n1777) );
  XOR U2323 ( .A(n4571), .B(n4570), .Z(n4559) );
  XOR U2324 ( .A(n4896), .B(n4895), .Z(n4884) );
  MUX U2325 ( .IN0(n6566), .IN1(n6568), .SEL(n6567), .F(n166) );
  IV U2326 ( .A(n166), .Z(n4856) );
  MUX U2327 ( .IN0(n5525), .IN1(n5527), .SEL(n5526), .F(n167) );
  IV U2328 ( .A(n167), .Z(n4273) );
  MUX U2329 ( .IN0(n5297), .IN1(n5299), .SEL(n5298), .F(n168) );
  IV U2330 ( .A(n168), .Z(n4143) );
  XOR U2331 ( .A(n4116), .B(n4115), .Z(n4104) );
  XOR U2332 ( .A(n1367), .B(n1366), .Z(n1360) );
  XOR U2333 ( .A(n1343), .B(n1342), .Z(n1350) );
  MUX U2334 ( .IN0(n4469), .IN1(n169), .SEL(n4470), .F(n3717) );
  IV U2335 ( .A(n4471), .Z(n169) );
  XOR U2336 ( .A(n3668), .B(n3667), .Z(n3675) );
  MUX U2337 ( .IN0(n253), .IN1(n4050), .SEL(n4049), .F(n170) );
  IV U2338 ( .A(n170), .Z(n3507) );
  XOR U2339 ( .A(n3555), .B(n3554), .Z(n3562) );
  XOR U2340 ( .A(n3929), .B(n3927), .Z(n3921) );
  MUX U2341 ( .IN0(n4824), .IN1(n171), .SEL(n4825), .F(n3890) );
  IV U2342 ( .A(n4826), .Z(n171) );
  XOR U2343 ( .A(n3828), .B(n3827), .Z(n3835) );
  XOR U2344 ( .A(n3797), .B(n3796), .Z(n3804) );
  MUX U2345 ( .IN0(n257), .IN1(n3941), .SEL(n3940), .F(n172) );
  IV U2346 ( .A(n172), .Z(n3456) );
  MUX U2347 ( .IN0(n3603), .IN1(n173), .SEL(n3604), .F(n3295) );
  IV U2348 ( .A(n3605), .Z(n173) );
  MUX U2349 ( .IN0(n3523), .IN1(n174), .SEL(n3524), .F(n3257) );
  IV U2350 ( .A(n3525), .Z(n174) );
  MUX U2351 ( .IN0(n3493), .IN1(n3496), .SEL(n3494), .F(n3487) );
  XOR U2352 ( .A(n1297), .B(n1295), .Z(n1304) );
  MUX U2353 ( .IN0(n586), .IN1(n1756), .SEL(n1754), .F(n1749) );
  MUX U2354 ( .IN0(n666), .IN1(n1955), .SEL(n1953), .F(n1946) );
  MUX U2355 ( .IN0(n668), .IN1(n1884), .SEL(n1882), .F(n1354) );
  MUX U2356 ( .IN0(n669), .IN1(n1911), .SEL(n1909), .F(n1904) );
  MUX U2357 ( .IN0(n517), .IN1(n1600), .SEL(n1598), .F(n1594) );
  MUX U2358 ( .IN0(n672), .IN1(n1578), .SEL(n1576), .F(n1571) );
  XOR U2359 ( .A(n1155), .B(n1153), .Z(n1162) );
  MUX U2360 ( .IN0(n523), .IN1(n1665), .SEL(n1663), .F(n1659) );
  MUX U2361 ( .IN0(n684), .IN1(n1643), .SEL(n1641), .F(n1636) );
  MUX U2362 ( .IN0(n686), .IN1(n1617), .SEL(n1615), .F(n1610) );
  MUX U2363 ( .IN0(n687), .IN1(n1627), .SEL(n1625), .F(n1618) );
  MUX U2364 ( .IN0(n525), .IN1(n1697), .SEL(n1695), .F(n1691) );
  MUX U2365 ( .IN0(n1263), .IN1(n175), .SEL(n1264), .F(n1044) );
  IV U2366 ( .A(n1265), .Z(n175) );
  MUX U2367 ( .IN0(n3973), .IN1(n3976), .SEL(n3974), .F(n3967) );
  MUX U2368 ( .IN0(n3876), .IN1(n3879), .SEL(n3877), .F(n3872) );
  MUX U2369 ( .IN0(n3784), .IN1(n3787), .SEL(n3785), .F(n3778) );
  MUX U2370 ( .IN0(n3818), .IN1(n3821), .SEL(n3819), .F(n3398) );
  MUX U2371 ( .IN0(n3852), .IN1(n3855), .SEL(n3853), .F(n3848) );
  MUX U2372 ( .IN0(n3589), .IN1(n3592), .SEL(n3590), .F(n3583) );
  MUX U2373 ( .IN0(n3655), .IN1(n3658), .SEL(n3656), .F(n3649) );
  MUX U2374 ( .IN0(n3641), .IN1(n3644), .SEL(n3642), .F(n3314) );
  MUX U2375 ( .IN0(n3702), .IN1(n176), .SEL(n3703), .F(n3341) );
  IV U2376 ( .A(n3704), .Z(n176) );
  XOR U2377 ( .A(n6379), .B(n6378), .Z(n6337) );
  MUX U2378 ( .IN0(n2017), .IN1(n2015), .SEL(n2016), .F(n177) );
  IV U2379 ( .A(n177), .Z(n1416) );
  XOR U2380 ( .A(n5028), .B(n436), .Z(n6824) );
  MUX U2381 ( .IN0(n1761), .IN1(n178), .SEL(n1762), .F(n1290) );
  IV U2382 ( .A(n1763), .Z(n178) );
  MUX U2383 ( .IN0(n1632), .IN1(n179), .SEL(n1633), .F(n1228) );
  IV U2384 ( .A(n1634), .Z(n179) );
  MUX U2385 ( .IN0(n1567), .IN1(n180), .SEL(n1568), .F(n1195) );
  IV U2386 ( .A(n1569), .Z(n180) );
  XOR U2387 ( .A(n1170), .B(n1169), .Z(n1158) );
  MUX U2388 ( .IN0(n2055), .IN1(n2053), .SEL(n2054), .F(n1447) );
  XOR U2389 ( .A(n997), .B(n995), .Z(n989) );
  XOR U2390 ( .A(n3420), .B(n3419), .Z(n3413) );
  MUX U2391 ( .IN0(n3822), .IN1(n181), .SEL(n3823), .F(n3399) );
  IV U2392 ( .A(n3824), .Z(n181) );
  MUX U2393 ( .IN0(n3791), .IN1(n182), .SEL(n3792), .F(n3383) );
  IV U2394 ( .A(n3793), .Z(n182) );
  MUX U2395 ( .IN0(n3662), .IN1(n183), .SEL(n3663), .F(n3322) );
  IV U2396 ( .A(n3664), .Z(n183) );
  MUX U2397 ( .IN0(n2108), .IN1(n2106), .SEL(n2107), .F(n2102) );
  MUX U2398 ( .IN0(n2088), .IN1(n2086), .SEL(n2087), .F(n2080) );
  MUX U2399 ( .IN0(n184), .IN1(n2005), .SEL(n2006), .F(n1411) );
  IV U2400 ( .A(n2007), .Z(n184) );
  MUX U2401 ( .IN0(n1282), .IN1(n1285), .SEL(n1283), .F(n1278) );
  MUX U2402 ( .IN0(n1326), .IN1(n185), .SEL(n1327), .F(n1077) );
  IV U2403 ( .A(n1328), .Z(n185) );
  MUX U2404 ( .IN0(n1376), .IN1(n1379), .SEL(n1377), .F(n1372) );
  XOR U2405 ( .A(n1005), .B(n1003), .Z(n1012) );
  MUX U2406 ( .IN0(n3434), .IN1(n3437), .SEL(n3435), .F(n3430) );
  MUX U2407 ( .IN0(n3365), .IN1(n186), .SEL(n3366), .F(n3181) );
  IV U2408 ( .A(n3367), .Z(n186) );
  MUX U2409 ( .IN0(n3307), .IN1(n3310), .SEL(n3308), .F(n3303) );
  MUX U2410 ( .IN0(n3337), .IN1(n187), .SEL(n3338), .F(n3166) );
  IV U2411 ( .A(n3339), .Z(n187) );
  MUX U2412 ( .IN0(n3358), .IN1(n3361), .SEL(n3359), .F(n3176) );
  MUX U2413 ( .IN0(n5610), .IN1(n5612), .SEL(n5611), .F(n188) );
  IV U2414 ( .A(n188), .Z(n4321) );
  MUX U2415 ( .IN0(n556), .IN1(n4191), .SEL(n4190), .F(n189) );
  IV U2416 ( .A(n189), .Z(n3579) );
  MUX U2417 ( .IN0(n555), .IN1(n4972), .SEL(n4971), .F(n190) );
  IV U2418 ( .A(n190), .Z(n3963) );
  MUX U2419 ( .IN0(n764), .IN1(n1451), .SEL(n1449), .F(n1138) );
  XOR U2420 ( .A(n3275), .B(n3274), .Z(n3293) );
  XOR U2421 ( .A(n3129), .B(n3127), .Z(n3121) );
  XOR U2422 ( .A(n3227), .B(n3225), .Z(n3234) );
  MUX U2423 ( .IN0(n3183), .IN1(n191), .SEL(n3184), .F(n3090) );
  IV U2424 ( .A(n3185), .Z(n191) );
  MUX U2425 ( .IN0(n1068), .IN1(n192), .SEL(n1069), .F(n943) );
  IV U2426 ( .A(n1070), .Z(n192) );
  MUX U2427 ( .IN0(n952), .IN1(n193), .SEL(n953), .F(n883) );
  IV U2428 ( .A(n954), .Z(n193) );
  MUX U2429 ( .IN0(n1111), .IN1(n1114), .SEL(n1112), .F(n1107) );
  XNOR U2430 ( .A(n1084), .B(n1085), .Z(n949) );
  MUX U2431 ( .IN0(n1035), .IN1(n194), .SEL(n1036), .F(n928) );
  IV U2432 ( .A(n1037), .Z(n194) );
  MUX U2433 ( .IN0(n3217), .IN1(n3219), .SEL(n3218), .F(n3104) );
  MUX U2434 ( .IN0(n3069), .IN1(n195), .SEL(n3070), .F(n3040) );
  IV U2435 ( .A(n3071), .Z(n195) );
  MUX U2436 ( .IN0(n282), .IN1(n1454), .SEL(n1453), .F(n196) );
  IV U2437 ( .A(n196), .Z(n1139) );
  MUX U2438 ( .IN0(n3548), .IN1(n197), .SEL(n3549), .F(n3268) );
  IV U2439 ( .A(n3550), .Z(n197) );
  XOR U2440 ( .A(n921), .B(n920), .Z(n909) );
  MUX U2441 ( .IN0(n565), .IN1(n1994), .SEL(n1995), .F(n198) );
  IV U2442 ( .A(n198), .Z(n3998) );
  MUX U2443 ( .IN0(n1046), .IN1(n973), .SEL(n1047), .F(n930) );
  MUX U2444 ( .IN0(n970), .IN1(n199), .SEL(n971), .F(n898) );
  IV U2445 ( .A(n972), .Z(n199) );
  MUX U2446 ( .IN0(n3116), .IN1(n200), .SEL(n892), .F(n3059) );
  IV U2447 ( .A(n891), .Z(n200) );
  MUX U2448 ( .IN0(n863), .IN1(n866), .SEL(n864), .F(n859) );
  MUX U2449 ( .IN0(n879), .IN1(n201), .SEL(n880), .F(n845) );
  IV U2450 ( .A(n881), .Z(n201) );
  MUX U2451 ( .IN0(n3042), .IN1(n3045), .SEL(n3043), .F(n3026) );
  MUX U2452 ( .IN0(n3028), .IN1(n3031), .SEL(n3029), .F(n3027) );
  MUX U2453 ( .IN0(n2634), .IN1(n2632), .SEL(n2633), .F(n202) );
  IV U2454 ( .A(n202), .Z(n1775) );
  MUX U2455 ( .IN0(n6272), .IN1(n6270), .SEL(n6271), .F(n203) );
  IV U2456 ( .A(n203), .Z(n4694) );
  MUX U2457 ( .IN0(n5459), .IN1(n5457), .SEL(n5458), .F(n204) );
  IV U2458 ( .A(n204), .Z(n4239) );
  MUX U2459 ( .IN0(n6631), .IN1(n6629), .SEL(n6630), .F(n205) );
  IV U2460 ( .A(n205), .Z(n4894) );
  MUX U2461 ( .IN0(n6456), .IN1(n6454), .SEL(n6455), .F(n206) );
  IV U2462 ( .A(n206), .Z(n4795) );
  MUX U2463 ( .IN0(n5075), .IN1(n5073), .SEL(n5074), .F(n207) );
  IV U2464 ( .A(n207), .Z(n4018) );
  MUX U2465 ( .IN0(n208), .IN1(n5136), .SEL(n5137), .F(n4054) );
  IV U2466 ( .A(n5138), .Z(n208) );
  MUX U2467 ( .IN0(n209), .IN1(n5049), .SEL(n5050), .F(n4005) );
  IV U2468 ( .A(n5051), .Z(n209) );
  MUX U2469 ( .IN0(n5193), .IN1(n5191), .SEL(n5192), .F(n5185) );
  MUX U2470 ( .IN0(n5206), .IN1(n5204), .SEL(n5205), .F(n210) );
  IV U2471 ( .A(n210), .Z(n4090) );
  MUX U2472 ( .IN0(n5160), .IN1(n5158), .SEL(n5159), .F(n4074) );
  MUX U2473 ( .IN0(n211), .IN1(n5222), .SEL(n5223), .F(n4101) );
  IV U2474 ( .A(n5224), .Z(n211) );
  MUX U2475 ( .IN0(n5234), .IN1(n5232), .SEL(n5233), .F(n212) );
  IV U2476 ( .A(n212), .Z(n4106) );
  MUX U2477 ( .IN0(n5255), .IN1(n5253), .SEL(n5254), .F(n5249) );
  MUX U2478 ( .IN0(n2947), .IN1(n2945), .SEL(n2946), .F(n213) );
  IV U2479 ( .A(n213), .Z(n1958) );
  MUX U2480 ( .IN0(n2862), .IN1(n2860), .SEL(n2861), .F(n214) );
  IV U2481 ( .A(n214), .Z(n1905) );
  MUX U2482 ( .IN0(n2891), .IN1(n2889), .SEL(n2890), .F(n215) );
  IV U2483 ( .A(n215), .Z(n1924) );
  MUX U2484 ( .IN0(n2285), .IN1(n2283), .SEL(n2284), .F(n216) );
  IV U2485 ( .A(n216), .Z(n1572) );
  MUX U2486 ( .IN0(n2381), .IN1(n2379), .SEL(n2380), .F(n217) );
  IV U2487 ( .A(n217), .Z(n1630) );
  MUX U2488 ( .IN0(n218), .IN1(n2652), .SEL(n2653), .F(n1784) );
  IV U2489 ( .A(n2654), .Z(n218) );
  MUX U2490 ( .IN0(n219), .IN1(n2710), .SEL(n2711), .F(n1815) );
  IV U2491 ( .A(n2712), .Z(n219) );
  XOR U2492 ( .A(n2688), .B(n2689), .Z(n1805) );
  MUX U2493 ( .IN0(n2737), .IN1(n2735), .SEL(n2736), .F(n2731) );
  MUX U2494 ( .IN0(n220), .IN1(n2779), .SEL(n2780), .F(n1857) );
  IV U2495 ( .A(n2781), .Z(n220) );
  MUX U2496 ( .IN0(n221), .IN1(n6864), .SEL(n6865), .F(n5026) );
  IV U2497 ( .A(n6866), .Z(n221) );
  MUX U2498 ( .IN0(n6800), .IN1(n6798), .SEL(n6799), .F(n4999) );
  MUX U2499 ( .IN0(n222), .IN1(n6677), .SEL(n6678), .F(n4920) );
  IV U2500 ( .A(n6679), .Z(n222) );
  MUX U2501 ( .IN0(n6730), .IN1(n6728), .SEL(n6729), .F(n4955) );
  MUX U2502 ( .IN0(n223), .IN1(n6721), .SEL(n6722), .F(n4943) );
  IV U2503 ( .A(n6723), .Z(n223) );
  MUX U2504 ( .IN0(n224), .IN1(n6519), .SEL(n6520), .F(n4830) );
  IV U2505 ( .A(n6521), .Z(n224) );
  MUX U2506 ( .IN0(n225), .IN1(n6430), .SEL(n6431), .F(n4782) );
  IV U2507 ( .A(n6432), .Z(n225) );
  MUX U2508 ( .IN0(n226), .IN1(n6563), .SEL(n6564), .F(n4855) );
  IV U2509 ( .A(n6565), .Z(n226) );
  MUX U2510 ( .IN0(n227), .IN1(n6605), .SEL(n6606), .F(n4879) );
  IV U2511 ( .A(n6607), .Z(n227) );
  MUX U2512 ( .IN0(n6140), .IN1(n6138), .SEL(n6139), .F(n4628) );
  MUX U2513 ( .IN0(n228), .IN1(n6085), .SEL(n6086), .F(n4590) );
  IV U2514 ( .A(n6087), .Z(n228) );
  MUX U2515 ( .IN0(n6020), .IN1(n6018), .SEL(n6019), .F(n6014) );
  MUX U2516 ( .IN0(n6000), .IN1(n5998), .SEL(n5999), .F(n5992) );
  MUX U2517 ( .IN0(n229), .IN1(n6029), .SEL(n6030), .F(n4556) );
  IV U2518 ( .A(n6031), .Z(n229) );
  MUX U2519 ( .IN0(n6052), .IN1(n6050), .SEL(n6051), .F(n4577) );
  MUX U2520 ( .IN0(n230), .IN1(n6070), .SEL(n6071), .F(n4581) );
  IV U2521 ( .A(n6072), .Z(n230) );
  MUX U2522 ( .IN0(n6309), .IN1(n6307), .SEL(n6308), .F(n6303) );
  MUX U2523 ( .IN0(n6206), .IN1(n6204), .SEL(n6205), .F(n6198) );
  MUX U2524 ( .IN0(n6244), .IN1(n6242), .SEL(n6243), .F(n231) );
  IV U2525 ( .A(n231), .Z(n4676) );
  MUX U2526 ( .IN0(n6358), .IN1(n6356), .SEL(n6357), .F(n232) );
  IV U2527 ( .A(n232), .Z(n4740) );
  MUX U2528 ( .IN0(n5488), .IN1(n5486), .SEL(n5487), .F(n4258) );
  MUX U2529 ( .IN0(n233), .IN1(n5310), .SEL(n5311), .F(n4149) );
  IV U2530 ( .A(n5312), .Z(n233) );
  MUX U2531 ( .IN0(n5293), .IN1(n5291), .SEL(n5292), .F(n5285) );
  MUX U2532 ( .IN0(n234), .IN1(n5338), .SEL(n5339), .F(n4165) );
  IV U2533 ( .A(n5340), .Z(n234) );
  MUX U2534 ( .IN0(n5361), .IN1(n5359), .SEL(n5360), .F(n4184) );
  MUX U2535 ( .IN0(n235), .IN1(n5379), .SEL(n5380), .F(n4188) );
  IV U2536 ( .A(n5381), .Z(n235) );
  MUX U2537 ( .IN0(n5677), .IN1(n5675), .SEL(n5676), .F(n4369) );
  MUX U2538 ( .IN0(n236), .IN1(n5622), .SEL(n5623), .F(n4331) );
  IV U2539 ( .A(n5624), .Z(n236) );
  MUX U2540 ( .IN0(n5557), .IN1(n5555), .SEL(n5556), .F(n5551) );
  MUX U2541 ( .IN0(n237), .IN1(n5522), .SEL(n5523), .F(n4272) );
  IV U2542 ( .A(n5524), .Z(n237) );
  MUX U2543 ( .IN0(n238), .IN1(n5829), .SEL(n5830), .F(n4443) );
  IV U2544 ( .A(n5831), .Z(n238) );
  MUX U2545 ( .IN0(n5765), .IN1(n5763), .SEL(n5764), .F(n4415) );
  MUX U2546 ( .IN0(n5908), .IN1(n5906), .SEL(n5907), .F(n5902) );
  MUX U2547 ( .IN0(n5863), .IN1(n5861), .SEL(n5862), .F(n5857) );
  MUX U2548 ( .IN0(n5936), .IN1(n5934), .SEL(n5935), .F(n5930) );
  XOR U2549 ( .A(n1876), .B(n1874), .Z(n1868) );
  XOR U2550 ( .A(n1760), .B(n1758), .Z(n1752) );
  MUX U2551 ( .IN0(n6377), .IN1(n6379), .SEL(n6378), .F(n239) );
  IV U2552 ( .A(n239), .Z(n4752) );
  MUX U2553 ( .IN0(n6867), .IN1(n6869), .SEL(n6868), .F(n240) );
  IV U2554 ( .A(n240), .Z(n5027) );
  XOR U2555 ( .A(n5003), .B(n5001), .Z(n4995) );
  XOR U2556 ( .A(n4978), .B(n4976), .Z(n4985) );
  XOR U2557 ( .A(n4475), .B(n4474), .Z(n4482) );
  MUX U2558 ( .IN0(n5745), .IN1(n5747), .SEL(n5746), .F(n241) );
  IV U2559 ( .A(n241), .Z(n4397) );
  XOR U2560 ( .A(n4279), .B(n4278), .Z(n4286) );
  MUX U2561 ( .IN0(n5341), .IN1(n5343), .SEL(n5342), .F(n242) );
  IV U2562 ( .A(n242), .Z(n4166) );
  XOR U2563 ( .A(n4247), .B(n4246), .Z(n4254) );
  MUX U2564 ( .IN0(n5397), .IN1(n5399), .SEL(n5398), .F(n243) );
  IV U2565 ( .A(n243), .Z(n4198) );
  MUX U2566 ( .IN0(n4296), .IN1(n244), .SEL(n4297), .F(n3632) );
  IV U2567 ( .A(n4298), .Z(n244) );
  MUX U2568 ( .IN0(n572), .IN1(n4065), .SEL(n4063), .F(n4058) );
  MUX U2569 ( .IN0(n389), .IN1(n4030), .SEL(n4028), .F(n3499) );
  MUX U2570 ( .IN0(n466), .IN1(n4078), .SEL(n4076), .F(n3522) );
  MUX U2571 ( .IN0(n467), .IN1(n4124), .SEL(n4122), .F(n3547) );
  XOR U2572 ( .A(n2973), .B(n2974), .Z(n1972) );
  MUX U2573 ( .IN0(n2929), .IN1(n2927), .SEL(n2928), .F(n2923) );
  MUX U2574 ( .IN0(n245), .IN1(n2910), .SEL(n2911), .F(n1934) );
  IV U2575 ( .A(n2912), .Z(n245) );
  MUX U2576 ( .IN0(n2841), .IN1(n2839), .SEL(n2840), .F(n2835) );
  MUX U2577 ( .IN0(n246), .IN1(n2822), .SEL(n2823), .F(n1884) );
  IV U2578 ( .A(n2824), .Z(n246) );
  MUX U2579 ( .IN0(n2323), .IN1(n2321), .SEL(n2322), .F(n1600) );
  XOR U2580 ( .A(n1590), .B(n1588), .Z(n1596) );
  MUX U2581 ( .IN0(n2166), .IN1(n2164), .SEL(n2165), .F(n2160) );
  XOR U2582 ( .A(n1494), .B(n1492), .Z(n1501) );
  MUX U2583 ( .IN0(n2125), .IN1(n2123), .SEL(n2124), .F(n2119) );
  MUX U2584 ( .IN0(n2194), .IN1(n2192), .SEL(n2193), .F(n2188) );
  XOR U2585 ( .A(n1510), .B(n1508), .Z(n1516) );
  MUX U2586 ( .IN0(n2208), .IN1(n2206), .SEL(n2207), .F(n2202) );
  MUX U2587 ( .IN0(n2215), .IN1(n2213), .SEL(n2214), .F(n2209) );
  MUX U2588 ( .IN0(n2405), .IN1(n2403), .SEL(n2404), .F(n2399) );
  MUX U2589 ( .IN0(n2362), .IN1(n2360), .SEL(n2361), .F(n2356) );
  MUX U2590 ( .IN0(n2342), .IN1(n2340), .SEL(n2341), .F(n2336) );
  MUX U2591 ( .IN0(n247), .IN1(n2471), .SEL(n2472), .F(n1679) );
  IV U2592 ( .A(n2473), .Z(n247) );
  MUX U2593 ( .IN0(n2532), .IN1(n2530), .SEL(n2531), .F(n2526) );
  MUX U2594 ( .IN0(n582), .IN1(n1795), .SEL(n1793), .F(n1788) );
  MUX U2595 ( .IN0(n587), .IN1(n1826), .SEL(n1824), .F(n1819) );
  MUX U2596 ( .IN0(n589), .IN1(n1842), .SEL(n1840), .F(n1835) );
  MUX U2597 ( .IN0(n591), .IN1(n1853), .SEL(n1851), .F(n1844) );
  MUX U2598 ( .IN0(n592), .IN1(n5037), .SEL(n5035), .F(n5030) );
  MUX U2599 ( .IN0(n597), .IN1(n4916), .SEL(n4914), .F(n4909) );
  MUX U2600 ( .IN0(n600), .IN1(n4841), .SEL(n4839), .F(n4834) );
  MUX U2601 ( .IN0(n402), .IN1(n4852), .SEL(n4850), .F(n4843) );
  MUX U2602 ( .IN0(n4629), .IN1(n4631), .SEL(n4630), .F(n3797) );
  MUX U2603 ( .IN0(n4700), .IN1(n4703), .SEL(n4701), .F(n3839) );
  XNOR U2604 ( .A(n4683), .B(n4684), .Z(n3826) );
  MUX U2605 ( .IN0(n415), .IN1(n4738), .SEL(n4737), .F(n248) );
  IV U2606 ( .A(n248), .Z(n3849) );
  MUX U2607 ( .IN0(n626), .IN1(n4751), .SEL(n4749), .F(n3865) );
  MUX U2608 ( .IN0(n632), .IN1(n4197), .SEL(n4195), .F(n3592) );
  MUX U2609 ( .IN0(n633), .IN1(n4160), .SEL(n4158), .F(n4153) );
  XNOR U2610 ( .A(n4131), .B(n4132), .Z(n3553) );
  MUX U2611 ( .IN0(n4370), .IN1(n4372), .SEL(n4371), .F(n3668) );
  MUX U2612 ( .IN0(n643), .IN1(n4268), .SEL(n4266), .F(n4261) );
  MUX U2613 ( .IN0(n647), .IN1(n4454), .SEL(n4452), .F(n4447) );
  MUX U2614 ( .IN0(n650), .IN1(n4396), .SEL(n4394), .F(n3690) );
  MUX U2615 ( .IN0(n312), .IN1(n4419), .SEL(n4417), .F(n3694) );
  MUX U2616 ( .IN0(n4466), .IN1(n4468), .SEL(n4467), .F(n3716) );
  MUX U2617 ( .IN0(n4492), .IN1(n249), .SEL(n4493), .F(n3729) );
  IV U2618 ( .A(n4494), .Z(n249) );
  MUX U2619 ( .IN0(n2416), .IN1(n2418), .SEL(n2417), .F(n250) );
  IV U2620 ( .A(n250), .Z(n1648) );
  XOR U2621 ( .A(n1623), .B(n1622), .Z(n1609) );
  MUX U2622 ( .IN0(n2303), .IN1(n2305), .SEL(n2304), .F(n251) );
  IV U2623 ( .A(n251), .Z(n1583) );
  MUX U2624 ( .IN0(n2811), .IN1(n2813), .SEL(n2812), .F(n252) );
  IV U2625 ( .A(n252), .Z(n1877) );
  XOR U2626 ( .A(n1800), .B(n1799), .Z(n1818) );
  XOR U2627 ( .A(n1768), .B(n1767), .Z(n1787) );
  XOR U2628 ( .A(n4687), .B(n4686), .Z(n4706) );
  XOR U2629 ( .A(n4669), .B(n4668), .Z(n4657) );
  MUX U2630 ( .IN0(n5123), .IN1(n5125), .SEL(n5124), .F(n253) );
  IV U2631 ( .A(n253), .Z(n4048) );
  XOR U2632 ( .A(n3701), .B(n3700), .Z(n3708) );
  MUX U2633 ( .IN0(n437), .IN1(n4375), .SEL(n4374), .F(n254) );
  IV U2634 ( .A(n254), .Z(n3669) );
  MUX U2635 ( .IN0(n4079), .IN1(n255), .SEL(n4080), .F(n3523) );
  IV U2636 ( .A(n4081), .Z(n255) );
  XOR U2637 ( .A(n3506), .B(n3505), .Z(n3513) );
  MUX U2638 ( .IN0(n4856), .IN1(n256), .SEL(n4857), .F(n3905) );
  IV U2639 ( .A(n4858), .Z(n256) );
  XOR U2640 ( .A(n3889), .B(n3888), .Z(n3896) );
  XOR U2641 ( .A(n3986), .B(n3985), .Z(n3993) );
  MUX U2642 ( .IN0(n343), .IN1(n4923), .SEL(n4922), .F(n257) );
  IV U2643 ( .A(n257), .Z(n3939) );
  XOR U2644 ( .A(n3869), .B(n3867), .Z(n3861) );
  MUX U2645 ( .IN0(n435), .IN1(n4634), .SEL(n4633), .F(n258) );
  IV U2646 ( .A(n258), .Z(n3798) );
  MUX U2647 ( .IN0(n3556), .IN1(n259), .SEL(n3557), .F(n3273) );
  IV U2648 ( .A(n3558), .Z(n259) );
  XNOR U2649 ( .A(n3488), .B(n3489), .Z(n3242) );
  MUX U2650 ( .IN0(n664), .IN1(n1971), .SEL(n1969), .F(n1964) );
  XNOR U2651 ( .A(n1913), .B(n1914), .Z(n1365) );
  MUX U2652 ( .IN0(n676), .IN1(n1543), .SEL(n1541), .F(n1190) );
  MUX U2653 ( .IN0(n519), .IN1(n1486), .SEL(n1484), .F(n1155) );
  MUX U2654 ( .IN0(n685), .IN1(n1647), .SEL(n1645), .F(n1235) );
  MUX U2655 ( .IN0(n729), .IN1(n1682), .SEL(n1681), .F(n260) );
  IV U2656 ( .A(n260), .Z(n1251) );
  MUX U2657 ( .IN0(n527), .IN1(n1676), .SEL(n1674), .F(n1667) );
  MUX U2658 ( .IN0(n1279), .IN1(n261), .SEL(n1280), .F(n1052) );
  IV U2659 ( .A(n1281), .Z(n261) );
  MUX U2660 ( .IN0(n3946), .IN1(n3949), .SEL(n3947), .F(n3942) );
  MUX U2661 ( .IN0(n3912), .IN1(n3915), .SEL(n3913), .F(n3908) );
  MUX U2662 ( .IN0(n3805), .IN1(n3808), .SEL(n3806), .F(n3801) );
  MUX U2663 ( .IN0(n3745), .IN1(n3748), .SEL(n3746), .F(n3371) );
  MUX U2664 ( .IN0(n349), .IN1(n3831), .SEL(n3830), .F(n262) );
  IV U2665 ( .A(n262), .Z(n3403) );
  MUX U2666 ( .IN0(n3593), .IN1(n3595), .SEL(n3594), .F(n3290) );
  MUX U2667 ( .IN0(n3676), .IN1(n3679), .SEL(n3677), .F(n3672) );
  XOR U2668 ( .A(n1982), .B(n434), .Z(n2957) );
  MUX U2669 ( .IN0(n6251), .IN1(n6253), .SEL(n6252), .F(n263) );
  IV U2670 ( .A(n263), .Z(n4678) );
  MUX U2671 ( .IN0(n6133), .IN1(n6135), .SEL(n6134), .F(n264) );
  IV U2672 ( .A(n264), .Z(n4615) );
  MUX U2673 ( .IN0(n6821), .IN1(n6823), .SEL(n6822), .F(n265) );
  IV U2674 ( .A(n265), .Z(n5004) );
  MUX U2675 ( .IN0(n6476), .IN1(n6478), .SEL(n6477), .F(n266) );
  IV U2676 ( .A(n266), .Z(n4807) );
  MUX U2677 ( .IN0(n5670), .IN1(n5672), .SEL(n5671), .F(n267) );
  IV U2678 ( .A(n267), .Z(n4356) );
  MUX U2679 ( .IN0(n5438), .IN1(n5440), .SEL(n5439), .F(n268) );
  IV U2680 ( .A(n268), .Z(n4223) );
  XOR U2681 ( .A(n1360), .B(n1359), .Z(n1346) );
  MUX U2682 ( .IN0(n1290), .IN1(n269), .SEL(n1291), .F(n1054) );
  IV U2683 ( .A(n1292), .Z(n269) );
  XOR U2684 ( .A(n3382), .B(n3381), .Z(n3389) );
  XOR U2685 ( .A(n3361), .B(n3359), .Z(n3351) );
  MUX U2686 ( .IN0(n3695), .IN1(n270), .SEL(n3696), .F(n3337) );
  IV U2687 ( .A(n3697), .Z(n270) );
  XOR U2688 ( .A(n3321), .B(n3320), .Z(n3328) );
  MUX U2689 ( .IN0(n3245), .IN1(n271), .SEL(n3246), .F(n3119) );
  IV U2690 ( .A(n3247), .Z(n271) );
  MUX U2691 ( .IN0(n2098), .IN1(n2096), .SEL(n2097), .F(n1471) );
  MUX U2692 ( .IN0(n2028), .IN1(n2026), .SEL(n2027), .F(n1432) );
  MUX U2693 ( .IN0(n1398), .IN1(n1401), .SEL(n1399), .F(n1394) );
  XNOR U2694 ( .A(n1356), .B(n1357), .Z(n1093) );
  MUX U2695 ( .IN0(n1191), .IN1(n1194), .SEL(n1192), .F(n1005) );
  MUX U2696 ( .IN0(n1195), .IN1(n272), .SEL(n1196), .F(n1006) );
  IV U2697 ( .A(n1197), .Z(n272) );
  MUX U2698 ( .IN0(n543), .IN1(n1246), .SEL(n1244), .F(n1239) );
  XOR U2699 ( .A(n1020), .B(n1019), .Z(n1029) );
  MUX U2700 ( .IN0(n544), .IN1(n1261), .SEL(n1259), .F(n1254) );
  MUX U2701 ( .IN0(n1270), .IN1(n1273), .SEL(n1271), .F(n1045) );
  MUX U2702 ( .IN0(n1060), .IN1(n273), .SEL(n1061), .F(n939) );
  IV U2703 ( .A(n1062), .Z(n273) );
  MUX U2704 ( .IN0(n3463), .IN1(n3465), .SEL(n3464), .F(n3227) );
  MUX U2705 ( .IN0(n3423), .IN1(n3426), .SEL(n3424), .F(n3216) );
  MUX U2706 ( .IN0(n3448), .IN1(n3450), .SEL(n3449), .F(n3219) );
  MUX U2707 ( .IN0(n3372), .IN1(n3375), .SEL(n3373), .F(n3182) );
  MUX U2708 ( .IN0(n3411), .IN1(n274), .SEL(n3412), .F(n3204) );
  IV U2709 ( .A(n3413), .Z(n274) );
  MUX U2710 ( .IN0(n3298), .IN1(n3301), .SEL(n3299), .F(n3294) );
  XOR U2711 ( .A(n2476), .B(n2475), .Z(n2390) );
  XOR U2712 ( .A(n5183), .B(n5182), .Z(n5095) );
  XOR U2713 ( .A(n1451), .B(n1449), .Z(n1443) );
  XOR U2714 ( .A(n1458), .B(n1457), .Z(n1467) );
  MUX U2715 ( .IN0(n2898), .IN1(n2900), .SEL(n2899), .F(n275) );
  IV U2716 ( .A(n275), .Z(n1926) );
  MUX U2717 ( .IN0(n554), .IN1(n1537), .SEL(n1536), .F(n276) );
  IV U2718 ( .A(n276), .Z(n1179) );
  MUX U2719 ( .IN0(n3963), .IN1(n277), .SEL(n3964), .F(n3466) );
  IV U2720 ( .A(n3965), .Z(n277) );
  MUX U2721 ( .IN0(n3579), .IN1(n278), .SEL(n3580), .F(n3284) );
  IV U2722 ( .A(n3581), .Z(n278) );
  XOR U2723 ( .A(n944), .B(n942), .Z(n936) );
  XOR U2724 ( .A(n3137), .B(n3135), .Z(n3144) );
  MUX U2725 ( .IN0(n3376), .IN1(n279), .SEL(n3377), .F(n3183) );
  IV U2726 ( .A(n3378), .Z(n279) );
  MUX U2727 ( .IN0(n370), .IN1(n1145), .SEL(n1144), .F(n280) );
  IV U2728 ( .A(n280), .Z(n982) );
  MUX U2729 ( .IN0(n767), .IN1(n1436), .SEL(n1434), .F(n1131) );
  MUX U2730 ( .IN0(n1100), .IN1(n1103), .SEL(n1101), .F(n964) );
  MUX U2731 ( .IN0(n1089), .IN1(n1092), .SEL(n1090), .F(n1083) );
  MUX U2732 ( .IN0(n1013), .IN1(n1016), .SEL(n1014), .F(n1009) );
  MUX U2733 ( .IN0(n3235), .IN1(n3238), .SEL(n3236), .F(n3231) );
  MUX U2734 ( .IN0(n3195), .IN1(n281), .SEL(n3196), .F(n3099) );
  IV U2735 ( .A(n3197), .Z(n281) );
  MUX U2736 ( .IN0(n3150), .IN1(n3153), .SEL(n3151), .F(n3083) );
  XOR U2737 ( .A(n5788), .B(n5787), .Z(n5612) );
  MUX U2738 ( .IN0(n2076), .IN1(n2078), .SEL(n2077), .F(n282) );
  IV U2739 ( .A(n282), .Z(n1452) );
  MUX U2740 ( .IN0(n6651), .IN1(n6653), .SEL(n6652), .F(n283) );
  IV U2741 ( .A(n283), .Z(n4904) );
  MUX U2742 ( .IN0(n1079), .IN1(n284), .SEL(n1080), .F(n945) );
  IV U2743 ( .A(n1081), .Z(n284) );
  XOR U2744 ( .A(n3168), .B(n3167), .Z(n3156) );
  MUX U2745 ( .IN0(n3268), .IN1(n285), .SEL(n3269), .F(n3130) );
  IV U2746 ( .A(n3270), .Z(n285) );
  MUX U2747 ( .IN0(n1125), .IN1(n1128), .SEL(n1126), .F(n1120) );
  XOR U2748 ( .A(n3087), .B(n3085), .Z(n3079) );
  XOR U2749 ( .A(n3064), .B(n3062), .Z(n3071) );
  MUX U2750 ( .IN0(n903), .IN1(n906), .SEL(n904), .F(n866) );
  MUX U2751 ( .IN0(n3105), .IN1(n286), .SEL(n3106), .F(n3052) );
  IV U2752 ( .A(n3107), .Z(n286) );
  MUX U2753 ( .IN0(n1727), .IN1(n1437), .SEL(n1728), .F(n1274) );
  MUX U2754 ( .IN0(n3998), .IN1(n287), .SEL(n1405), .F(n3484) );
  IV U2755 ( .A(n1404), .Z(n287) );
  MUX U2756 ( .IN0(n871), .IN1(n873), .SEL(n872), .F(n840) );
  MUX U2757 ( .IN0(n867), .IN1(n870), .SEL(n868), .F(n839) );
  MUX U2758 ( .IN0(n3059), .IN1(n288), .SEL(n855), .F(n3032) );
  IV U2759 ( .A(n854), .Z(n288) );
  MUX U2760 ( .IN0(n848), .IN1(n851), .SEL(n849), .F(n843) );
  MUX U2761 ( .IN0(n3024), .IN1(n289), .SEL(n3025), .F(n822) );
  IV U2762 ( .A(n3026), .Z(n289) );
  MUX U2763 ( .IN0(n2679), .IN1(n2677), .SEL(n2678), .F(n290) );
  IV U2764 ( .A(n290), .Z(n1798) );
  MUX U2765 ( .IN0(n6317), .IN1(n6315), .SEL(n6316), .F(n291) );
  IV U2766 ( .A(n291), .Z(n4717) );
  MUX U2767 ( .IN0(n6831), .IN1(n6829), .SEL(n6830), .F(n292) );
  IV U2768 ( .A(n292), .Z(n5009) );
  MUX U2769 ( .IN0(n5448), .IN1(n5446), .SEL(n5447), .F(n293) );
  IV U2770 ( .A(n293), .Z(n4228) );
  MUX U2771 ( .IN0(n5145), .IN1(n5143), .SEL(n5144), .F(n4065) );
  XOR U2772 ( .A(n5128), .B(n5129), .Z(n4052) );
  XOR U2773 ( .A(n5112), .B(n5113), .Z(n4045) );
  MUX U2774 ( .IN0(n5068), .IN1(n5066), .SEL(n5067), .F(n5062) );
  MUX U2775 ( .IN0(n5213), .IN1(n5211), .SEL(n5212), .F(n5207) );
  MUX U2776 ( .IN0(n5248), .IN1(n5246), .SEL(n5247), .F(n294) );
  IV U2777 ( .A(n294), .Z(n4114) );
  MUX U2778 ( .IN0(n2398), .IN1(n2396), .SEL(n2397), .F(n295) );
  IV U2779 ( .A(n295), .Z(n1637) );
  MUX U2780 ( .IN0(n2661), .IN1(n2659), .SEL(n2660), .F(n1795) );
  MUX U2781 ( .IN0(n2630), .IN1(n2628), .SEL(n2629), .F(n2624) );
  MUX U2782 ( .IN0(n2588), .IN1(n2586), .SEL(n2587), .F(n2582) );
  MUX U2783 ( .IN0(n2719), .IN1(n2717), .SEL(n2718), .F(n1826) );
  MUX U2784 ( .IN0(n2757), .IN1(n2755), .SEL(n2756), .F(n2751) );
  MUX U2785 ( .IN0(n6873), .IN1(n6871), .SEL(n6872), .F(n5037) );
  MUX U2786 ( .IN0(n6796), .IN1(n6794), .SEL(n6795), .F(n6790) );
  MUX U2787 ( .IN0(n6702), .IN1(n6700), .SEL(n6701), .F(n4938) );
  XOR U2788 ( .A(n6685), .B(n6686), .Z(n4925) );
  MUX U2789 ( .IN0(n6528), .IN1(n6526), .SEL(n6527), .F(n4841) );
  XOR U2790 ( .A(n6511), .B(n6512), .Z(n4828) );
  XOR U2791 ( .A(n6495), .B(n6496), .Z(n4821) );
  MUX U2792 ( .IN0(n6449), .IN1(n6447), .SEL(n6448), .F(n6443) );
  MUX U2793 ( .IN0(n6596), .IN1(n6594), .SEL(n6595), .F(n6590) );
  MUX U2794 ( .IN0(n6624), .IN1(n6622), .SEL(n6623), .F(n6618) );
  MUX U2795 ( .IN0(n296), .IN1(n6176), .SEL(n6177), .F(n4638) );
  IV U2796 ( .A(n6178), .Z(n296) );
  MUX U2797 ( .IN0(n297), .IN1(n6160), .SEL(n6161), .F(n4631) );
  IV U2798 ( .A(n6162), .Z(n297) );
  MUX U2799 ( .IN0(n6104), .IN1(n6102), .SEL(n6103), .F(n6098) );
  MUX U2800 ( .IN0(n298), .IN1(n6130), .SEL(n6131), .F(n4614) );
  IV U2801 ( .A(n6132), .Z(n298) );
  MUX U2802 ( .IN0(n6010), .IN1(n6008), .SEL(n6009), .F(n4551) );
  MUX U2803 ( .IN0(n5981), .IN1(n5979), .SEL(n5980), .F(n299) );
  IV U2804 ( .A(n299), .Z(n4532) );
  MUX U2805 ( .IN0(n6048), .IN1(n6046), .SEL(n6047), .F(n6042) );
  MUX U2806 ( .IN0(n6055), .IN1(n6053), .SEL(n6054), .F(n300) );
  IV U2807 ( .A(n300), .Z(n4569) );
  MUX U2808 ( .IN0(n6258), .IN1(n6256), .SEL(n6257), .F(n4691) );
  MUX U2809 ( .IN0(n6226), .IN1(n6224), .SEL(n6225), .F(n6220) );
  MUX U2810 ( .IN0(n301), .IN1(n6207), .SEL(n6208), .F(n4654) );
  IV U2811 ( .A(n6209), .Z(n301) );
  MUX U2812 ( .IN0(n6233), .IN1(n6231), .SEL(n6232), .F(n302) );
  IV U2813 ( .A(n302), .Z(n4667) );
  MUX U2814 ( .IN0(n6247), .IN1(n6245), .SEL(n6246), .F(n6241) );
  MUX U2815 ( .IN0(n303), .IN1(n6346), .SEL(n6347), .F(n4735) );
  IV U2816 ( .A(n6348), .Z(n303) );
  MUX U2817 ( .IN0(n6393), .IN1(n6391), .SEL(n6392), .F(n6387) );
  MUX U2818 ( .IN0(n6407), .IN1(n6405), .SEL(n6406), .F(n6401) );
  MUX U2819 ( .IN0(n304), .IN1(n5479), .SEL(n5480), .F(n4247) );
  IV U2820 ( .A(n5481), .Z(n304) );
  MUX U2821 ( .IN0(n5413), .IN1(n5411), .SEL(n5412), .F(n5407) );
  MUX U2822 ( .IN0(n5431), .IN1(n5429), .SEL(n5430), .F(n305) );
  IV U2823 ( .A(n305), .Z(n4221) );
  MUX U2824 ( .IN0(n306), .IN1(n5294), .SEL(n5295), .F(n4142) );
  IV U2825 ( .A(n5296), .Z(n306) );
  MUX U2826 ( .IN0(n5357), .IN1(n5355), .SEL(n5356), .F(n5351) );
  MUX U2827 ( .IN0(n307), .IN1(n5713), .SEL(n5714), .F(n4379) );
  IV U2828 ( .A(n5715), .Z(n307) );
  MUX U2829 ( .IN0(n308), .IN1(n5697), .SEL(n5698), .F(n4372) );
  IV U2830 ( .A(n5699), .Z(n308) );
  MUX U2831 ( .IN0(n5641), .IN1(n5639), .SEL(n5640), .F(n5635) );
  MUX U2832 ( .IN0(n309), .IN1(n5667), .SEL(n5668), .F(n4355) );
  IV U2833 ( .A(n5669), .Z(n309) );
  MUX U2834 ( .IN0(n5547), .IN1(n5545), .SEL(n5546), .F(n4290) );
  XOR U2835 ( .A(n5530), .B(n5531), .Z(n4277) );
  MUX U2836 ( .IN0(n5578), .IN1(n5576), .SEL(n5577), .F(n310) );
  IV U2837 ( .A(n310), .Z(n4300) );
  MUX U2838 ( .IN0(n5793), .IN1(n5791), .SEL(n5792), .F(n4433) );
  MUX U2839 ( .IN0(n5761), .IN1(n5759), .SEL(n5760), .F(n5755) );
  MUX U2840 ( .IN0(n311), .IN1(n5742), .SEL(n5743), .F(n4396) );
  IV U2841 ( .A(n5744), .Z(n311) );
  MUX U2842 ( .IN0(n5779), .IN1(n5777), .SEL(n5778), .F(n312) );
  IV U2843 ( .A(n312), .Z(n4418) );
  MUX U2844 ( .IN0(n313), .IN1(n5889), .SEL(n5890), .F(n4475) );
  IV U2845 ( .A(n5891), .Z(n313) );
  MUX U2846 ( .IN0(n5853), .IN1(n5851), .SEL(n5852), .F(n4465) );
  MUX U2847 ( .IN0(n314), .IN1(n5873), .SEL(n5874), .F(n4468) );
  IV U2848 ( .A(n5875), .Z(n314) );
  MUX U2849 ( .IN0(n5926), .IN1(n5924), .SEL(n5925), .F(n4502) );
  MUX U2850 ( .IN0(n5943), .IN1(n5941), .SEL(n5942), .F(n315) );
  IV U2851 ( .A(n315), .Z(n4504) );
  XOR U2852 ( .A(n1831), .B(n1829), .Z(n1838) );
  XOR U2853 ( .A(n1776), .B(n1774), .Z(n1768) );
  XOR U2854 ( .A(n1735), .B(n1733), .Z(n1744) );
  MUX U2855 ( .IN0(n6293), .IN1(n6295), .SEL(n6294), .F(n316) );
  IV U2856 ( .A(n316), .Z(n4704) );
  XOR U2857 ( .A(n4540), .B(n4539), .Z(n4547) );
  MUX U2858 ( .IN0(n6179), .IN1(n6181), .SEL(n6180), .F(n317) );
  IV U2859 ( .A(n317), .Z(n4639) );
  XOR U2860 ( .A(n4590), .B(n4588), .Z(n4597) );
  XOR U2861 ( .A(n4953), .B(n475), .Z(n6727) );
  XOR U2862 ( .A(n5026), .B(n5025), .Z(n5033) );
  XOR U2863 ( .A(n4855), .B(n4854), .Z(n4848) );
  XOR U2864 ( .A(n4863), .B(n4861), .Z(n4870) );
  XOR U2865 ( .A(n4782), .B(n4781), .Z(n4789) );
  MUX U2866 ( .IN0(n5892), .IN1(n5894), .SEL(n5893), .F(n318) );
  IV U2867 ( .A(n318), .Z(n4476) );
  MUX U2868 ( .IN0(n5716), .IN1(n5718), .SEL(n5717), .F(n319) );
  IV U2869 ( .A(n319), .Z(n4380) );
  XOR U2870 ( .A(n4331), .B(n4329), .Z(n4338) );
  XOR U2871 ( .A(n4188), .B(n4186), .Z(n4180) );
  XOR U2872 ( .A(n4165), .B(n4163), .Z(n4172) );
  MUX U2873 ( .IN0(n5313), .IN1(n5315), .SEL(n5314), .F(n320) );
  IV U2874 ( .A(n320), .Z(n4150) );
  XOR U2875 ( .A(n4085), .B(n4084), .Z(n4092) );
  XOR U2876 ( .A(n4005), .B(n4003), .Z(n4012) );
  MUX U2877 ( .IN0(n4198), .IN1(n321), .SEL(n4199), .F(n3584) );
  IV U2878 ( .A(n4200), .Z(n321) );
  XNOR U2879 ( .A(n4036), .B(n4037), .Z(n3504) );
  MUX U2880 ( .IN0(n421), .IN1(n4057), .SEL(n4056), .F(n322) );
  IV U2881 ( .A(n322), .Z(n3511) );
  MUX U2882 ( .IN0(n579), .IN1(n4112), .SEL(n4110), .F(n4105) );
  MUX U2883 ( .IN0(n323), .IN1(n2997), .SEL(n2998), .F(n1980) );
  IV U2884 ( .A(n2999), .Z(n323) );
  MUX U2885 ( .IN0(n3000), .IN1(n3002), .SEL(n3001), .F(n324) );
  IV U2886 ( .A(n324), .Z(n1981) );
  MUX U2887 ( .IN0(n2922), .IN1(n2920), .SEL(n2921), .F(n325) );
  IV U2888 ( .A(n325), .Z(n1939) );
  MUX U2889 ( .IN0(n326), .IN1(n2808), .SEL(n2809), .F(n1876) );
  IV U2890 ( .A(n2810), .Z(n326) );
  MUX U2891 ( .IN0(n2825), .IN1(n2827), .SEL(n2826), .F(n327) );
  IV U2892 ( .A(n327), .Z(n1885) );
  MUX U2893 ( .IN0(n328), .IN1(n2895), .SEL(n2896), .F(n1925) );
  IV U2894 ( .A(n2897), .Z(n328) );
  MUX U2895 ( .IN0(n2292), .IN1(n2290), .SEL(n2291), .F(n2286) );
  MUX U2896 ( .IN0(n2317), .IN1(n2319), .SEL(n2318), .F(n329) );
  IV U2897 ( .A(n329), .Z(n1591) );
  MUX U2898 ( .IN0(n2250), .IN1(n2248), .SEL(n2249), .F(n2244) );
  MUX U2899 ( .IN0(n330), .IN1(n2231), .SEL(n2232), .F(n1543) );
  IV U2900 ( .A(n2233), .Z(n330) );
  MUX U2901 ( .IN0(n2257), .IN1(n2255), .SEL(n2256), .F(n331) );
  IV U2902 ( .A(n331), .Z(n1556) );
  MUX U2903 ( .IN0(n332), .IN1(n2272), .SEL(n2273), .F(n1566) );
  IV U2904 ( .A(n2274), .Z(n332) );
  MUX U2905 ( .IN0(n333), .IN1(n2147), .SEL(n2148), .F(n1494) );
  IV U2906 ( .A(n2149), .Z(n333) );
  MUX U2907 ( .IN0(n2150), .IN1(n2152), .SEL(n2151), .F(n334) );
  IV U2908 ( .A(n334), .Z(n1495) );
  MUX U2909 ( .IN0(n2184), .IN1(n2182), .SEL(n2183), .F(n1520) );
  MUX U2910 ( .IN0(n335), .IN1(n2175), .SEL(n2176), .F(n1510) );
  IV U2911 ( .A(n2177), .Z(n335) );
  MUX U2912 ( .IN0(n2198), .IN1(n2196), .SEL(n2197), .F(n1530) );
  MUX U2913 ( .IN0(n336), .IN1(n2216), .SEL(n2217), .F(n1534) );
  IV U2914 ( .A(n2218), .Z(n336) );
  MUX U2915 ( .IN0(n2446), .IN1(n2444), .SEL(n2445), .F(n2440) );
  XOR U2916 ( .A(n1655), .B(n1653), .Z(n1661) );
  MUX U2917 ( .IN0(n2355), .IN1(n2353), .SEL(n2354), .F(n337) );
  IV U2918 ( .A(n337), .Z(n1611) );
  MUX U2919 ( .IN0(n2494), .IN1(n2492), .SEL(n2493), .F(n1697) );
  MUX U2920 ( .IN0(n2451), .IN1(n2449), .SEL(n2450), .F(n1676) );
  MUX U2921 ( .IN0(n2522), .IN1(n2520), .SEL(n2521), .F(n1713) );
  MUX U2922 ( .IN0(n2512), .IN1(n2510), .SEL(n2511), .F(n2506) );
  MUX U2923 ( .IN0(n2546), .IN1(n2544), .SEL(n2545), .F(n2540) );
  MUX U2924 ( .IN0(n338), .IN1(n2554), .SEL(n2555), .F(n1726) );
  IV U2925 ( .A(n2556), .Z(n338) );
  MUX U2926 ( .IN0(n1781), .IN1(n1784), .SEL(n1782), .F(n1308) );
  MUX U2927 ( .IN0(n1812), .IN1(n1815), .SEL(n1813), .F(n1324) );
  MUX U2928 ( .IN0(n595), .IN1(n4978), .SEL(n4976), .F(n3976) );
  MUX U2929 ( .IN0(n474), .IN1(n4920), .SEL(n4918), .F(n3938) );
  MUX U2930 ( .IN0(n417), .IN1(n4930), .SEL(n4929), .F(n339) );
  IV U2931 ( .A(n339), .Z(n3943) );
  MUX U2932 ( .IN0(n400), .IN1(n4943), .SEL(n4941), .F(n3959) );
  XNOR U2933 ( .A(n4957), .B(n4958), .Z(n3960) );
  XNOR U2934 ( .A(n4812), .B(n4813), .Z(n3887) );
  MUX U2935 ( .IN0(n418), .IN1(n4833), .SEL(n4832), .F(n340) );
  IV U2936 ( .A(n340), .Z(n3894) );
  MUX U2937 ( .IN0(n607), .IN1(n4879), .SEL(n4877), .F(n3925) );
  MUX U2938 ( .IN0(n609), .IN1(n4649), .SEL(n4647), .F(n4642) );
  XNOR U2939 ( .A(n4620), .B(n4621), .Z(n3795) );
  XNOR U2940 ( .A(n4603), .B(n4604), .Z(n3788) );
  MUX U2941 ( .IN0(n4692), .IN1(n4695), .SEL(n4693), .F(n3828) );
  MUX U2942 ( .IN0(n621), .IN1(n4746), .SEL(n4744), .F(n4739) );
  MUX U2943 ( .IN0(n629), .IN1(n4258), .SEL(n4256), .F(n4251) );
  MUX U2944 ( .IN0(n634), .IN1(n4139), .SEL(n4137), .F(n4130) );
  MUX U2945 ( .IN0(n638), .IN1(n4390), .SEL(n4388), .F(n4383) );
  XNOR U2946 ( .A(n4361), .B(n4362), .Z(n3666) );
  XNOR U2947 ( .A(n4344), .B(n4345), .Z(n3659) );
  MUX U2948 ( .IN0(n498), .IN1(n4272), .SEL(n4270), .F(n3619) );
  MUX U2949 ( .IN0(n419), .IN1(n4282), .SEL(n4281), .F(n341) );
  IV U2950 ( .A(n341), .Z(n3624) );
  MUX U2951 ( .IN0(n4434), .IN1(n4436), .SEL(n4435), .F(n3701) );
  MUX U2952 ( .IN0(n651), .IN1(n4486), .SEL(n4484), .F(n4479) );
  XOR U2953 ( .A(n1849), .B(n1848), .Z(n1834) );
  MUX U2954 ( .IN0(n2699), .IN1(n2701), .SEL(n2700), .F(n342) );
  IV U2955 ( .A(n342), .Z(n1808) );
  XOR U2956 ( .A(n4525), .B(n4524), .Z(n4543) );
  XOR U2957 ( .A(n4961), .B(n4960), .Z(n4948) );
  MUX U2958 ( .IN0(n6680), .IN1(n6682), .SEL(n6681), .F(n343) );
  IV U2959 ( .A(n343), .Z(n4921) );
  MUX U2960 ( .IN0(n5816), .IN1(n5818), .SEL(n5817), .F(n344) );
  IV U2961 ( .A(n344), .Z(n4437) );
  XOR U2962 ( .A(n4411), .B(n4410), .Z(n4399) );
  MUX U2963 ( .IN0(n5466), .IN1(n5468), .SEL(n5467), .F(n345) );
  IV U2964 ( .A(n345), .Z(n4241) );
  XOR U2965 ( .A(n4070), .B(n4069), .Z(n4088) );
  XOR U2966 ( .A(n4022), .B(n4021), .Z(n4008) );
  XOR U2967 ( .A(n1313), .B(n1311), .Z(n1320) );
  MUX U2968 ( .IN0(n434), .IN1(n1976), .SEL(n1975), .F(n346) );
  IV U2969 ( .A(n346), .Z(n1391) );
  MUX U2970 ( .IN0(n1877), .IN1(n347), .SEL(n1878), .F(n1344) );
  IV U2971 ( .A(n1879), .Z(n347) );
  XOR U2972 ( .A(n3547), .B(n3545), .Z(n3539) );
  XOR U2973 ( .A(n3602), .B(n3601), .Z(n3609) );
  MUX U2974 ( .IN0(n436), .IN1(n5022), .SEL(n5021), .F(n348) );
  IV U2975 ( .A(n348), .Z(n3987) );
  XOR U2976 ( .A(n3844), .B(n3842), .Z(n3851) );
  MUX U2977 ( .IN0(n536), .IN1(n4698), .SEL(n4697), .F(n349) );
  IV U2978 ( .A(n349), .Z(n3829) );
  MUX U2979 ( .IN0(n3497), .IN1(n3499), .SEL(n3498), .F(n3244) );
  MUX U2980 ( .IN0(n3507), .IN1(n350), .SEL(n3508), .F(n3249) );
  IV U2981 ( .A(n3509), .Z(n350) );
  MUX U2982 ( .IN0(n663), .IN1(n1991), .SEL(n1989), .F(n1984) );
  MUX U2983 ( .IN0(n424), .IN1(n1934), .SEL(n1932), .F(n1379) );
  MUX U2984 ( .IN0(n515), .IN1(n1872), .SEL(n1870), .F(n1863) );
  MUX U2985 ( .IN0(n516), .IN1(n1921), .SEL(n1919), .F(n1912) );
  MUX U2986 ( .IN0(n673), .IN1(n1582), .SEL(n1580), .F(n1202) );
  MUX U2987 ( .IN0(n1583), .IN1(n351), .SEL(n1584), .F(n1203) );
  IV U2988 ( .A(n1585), .Z(n351) );
  MUX U2989 ( .IN0(n679), .IN1(n1505), .SEL(n1503), .F(n1498) );
  MUX U2990 ( .IN0(n428), .IN1(n1606), .SEL(n1604), .F(n1224) );
  MUX U2991 ( .IN0(n1286), .IN1(n1289), .SEL(n1287), .F(n1053) );
  MUX U2992 ( .IN0(n1298), .IN1(n352), .SEL(n1299), .F(n1060) );
  IV U2993 ( .A(n1300), .Z(n352) );
  MUX U2994 ( .IN0(n3977), .IN1(n3979), .SEL(n3978), .F(n3472) );
  MUX U2995 ( .IN0(n3880), .IN1(n3882), .SEL(n3881), .F(n3426) );
  MUX U2996 ( .IN0(n3890), .IN1(n353), .SEL(n3891), .F(n3431) );
  IV U2997 ( .A(n3892), .Z(n353) );
  MUX U2998 ( .IN0(n431), .IN1(n3911), .SEL(n3910), .F(n354) );
  IV U2999 ( .A(n354), .Z(n3446) );
  MUX U3000 ( .IN0(n3926), .IN1(n3929), .SEL(n3927), .F(n3450) );
  XNOR U3001 ( .A(n3779), .B(n3780), .Z(n3380) );
  MUX U3002 ( .IN0(n3798), .IN1(n355), .SEL(n3799), .F(n3387) );
  IV U3003 ( .A(n3800), .Z(n355) );
  MUX U3004 ( .IN0(n3763), .IN1(n356), .SEL(n3764), .F(n3374) );
  IV U3005 ( .A(n3765), .Z(n356) );
  MUX U3006 ( .IN0(n3836), .IN1(n3839), .SEL(n3837), .F(n3832) );
  MUX U3007 ( .IN0(n3563), .IN1(n3566), .SEL(n3564), .F(n3559) );
  XNOR U3008 ( .A(n3650), .B(n3651), .Z(n3319) );
  MUX U3009 ( .IN0(n3669), .IN1(n357), .SEL(n3670), .F(n3326) );
  IV U3010 ( .A(n3671), .Z(n357) );
  MUX U3011 ( .IN0(n3709), .IN1(n3712), .SEL(n3710), .F(n3705) );
  XOR U3012 ( .A(n2518), .B(n2517), .Z(n2476) );
  XOR U3013 ( .A(n2180), .B(n2179), .Z(n2138) );
  XOR U3014 ( .A(n6610), .B(n6609), .Z(n6568) );
  XOR U3015 ( .A(n1609), .B(n1608), .Z(n1650) );
  MUX U3016 ( .IN0(n2954), .IN1(n2956), .SEL(n2955), .F(n358) );
  IV U3017 ( .A(n358), .Z(n1960) );
  XOR U3018 ( .A(n4559), .B(n4558), .Z(n4536) );
  XOR U3019 ( .A(n4298), .B(n4297), .Z(n4275) );
  XOR U3020 ( .A(n4104), .B(n4103), .Z(n4081) );
  MUX U3021 ( .IN0(n5093), .IN1(n5095), .SEL(n5094), .F(n359) );
  IV U3022 ( .A(n359), .Z(n4031) );
  XOR U3023 ( .A(n1328), .B(n1327), .Z(n1316) );
  XOR U3024 ( .A(n3733), .B(n3732), .Z(n3719) );
  MUX U3025 ( .IN0(n4223), .IN1(n360), .SEL(n4224), .F(n3596) );
  IV U3026 ( .A(n4225), .Z(n360) );
  XOR U3027 ( .A(n3570), .B(n3569), .Z(n3558) );
  MUX U3028 ( .IN0(n4807), .IN1(n361), .SEL(n4808), .F(n3883) );
  IV U3029 ( .A(n4809), .Z(n361) );
  XOR U3030 ( .A(n3861), .B(n3860), .Z(n3847) );
  XOR U3031 ( .A(n3398), .B(n3396), .Z(n3405) );
  MUX U3032 ( .IN0(n3980), .IN1(n362), .SEL(n3981), .F(n3473) );
  IV U3033 ( .A(n3982), .Z(n362) );
  XOR U3034 ( .A(n3336), .B(n3335), .Z(n3343) );
  XOR U3035 ( .A(n2081), .B(n2082), .Z(n1456) );
  MUX U3036 ( .IN0(n1416), .IN1(n363), .SEL(n1417), .F(n1127) );
  IV U3037 ( .A(n1418), .Z(n363) );
  MUX U3038 ( .IN0(n1387), .IN1(n1390), .SEL(n1388), .F(n1114) );
  MUX U3039 ( .IN0(n1380), .IN1(n1382), .SEL(n1381), .F(n1103) );
  MUX U3040 ( .IN0(n1351), .IN1(n1354), .SEL(n1352), .F(n1347) );
  MUX U3041 ( .IN0(n1361), .IN1(n1364), .SEL(n1362), .F(n1355) );
  MUX U3042 ( .IN0(n539), .IN1(n1213), .SEL(n1211), .F(n1206) );
  MUX U3043 ( .IN0(n1152), .IN1(n1155), .SEL(n1153), .F(n993) );
  MUX U3044 ( .IN0(n1225), .IN1(n1227), .SEL(n1226), .F(n1020) );
  MUX U3045 ( .IN0(n1255), .IN1(n364), .SEL(n1256), .F(n1040) );
  IV U3046 ( .A(n1257), .Z(n364) );
  MUX U3047 ( .IN0(n3480), .IN1(n3483), .SEL(n3481), .F(n3476) );
  MUX U3048 ( .IN0(n3383), .IN1(n365), .SEL(n3384), .F(n3187) );
  IV U3049 ( .A(n3385), .Z(n365) );
  MUX U3050 ( .IN0(n3280), .IN1(n3283), .SEL(n3281), .F(n3137) );
  MUX U3051 ( .IN0(n3311), .IN1(n3314), .SEL(n3312), .F(n3153) );
  MUX U3052 ( .IN0(n3322), .IN1(n366), .SEL(n3323), .F(n3158) );
  IV U3053 ( .A(n3324), .Z(n366) );
  MUX U3054 ( .IN0(n2008), .IN1(n2010), .SEL(n2009), .F(n367) );
  IV U3055 ( .A(n367), .Z(n1412) );
  XOR U3056 ( .A(n1682), .B(n1681), .Z(n1634) );
  XOR U3057 ( .A(n1489), .B(n1488), .Z(n1569) );
  XOR U3058 ( .A(n4730), .B(n4729), .Z(n4680) );
  MUX U3059 ( .IN0(n6073), .IN1(n6075), .SEL(n6074), .F(n368) );
  IV U3060 ( .A(n368), .Z(n4582) );
  XOR U3061 ( .A(n4471), .B(n4470), .Z(n4422) );
  MUX U3062 ( .IN0(n1926), .IN1(n369), .SEL(n1927), .F(n1368) );
  IV U3063 ( .A(n1928), .Z(n369) );
  MUX U3064 ( .IN0(n553), .IN1(n1461), .SEL(n1460), .F(n370) );
  IV U3065 ( .A(n370), .Z(n1143) );
  MUX U3066 ( .IN0(n1179), .IN1(n371), .SEL(n1180), .F(n998) );
  IV U3067 ( .A(n1181), .Z(n371) );
  XOR U3068 ( .A(n1070), .B(n1069), .Z(n1058) );
  XOR U3069 ( .A(n3413), .B(n3412), .Z(n3401) );
  XOR U3070 ( .A(n3351), .B(n3350), .Z(n3339) );
  MUX U3071 ( .IN0(n3284), .IN1(n372), .SEL(n3285), .F(n3138) );
  IV U3072 ( .A(n3286), .Z(n372) );
  MUX U3073 ( .IN0(n3466), .IN1(n373), .SEL(n3467), .F(n3228) );
  IV U3074 ( .A(n3468), .Z(n373) );
  XNOR U3075 ( .A(n1463), .B(n1464), .Z(n1146) );
  MUX U3076 ( .IN0(n1002), .IN1(n1005), .SEL(n1003), .F(n917) );
  MUX U3077 ( .IN0(n994), .IN1(n997), .SEL(n995), .F(n906) );
  MUX U3078 ( .IN0(n1030), .IN1(n1033), .SEL(n1031), .F(n1026) );
  MUX U3079 ( .IN0(n1042), .IN1(n1045), .SEL(n1043), .F(n929) );
  MUX U3080 ( .IN0(n3224), .IN1(n3227), .SEL(n3225), .F(n3115) );
  MUX U3081 ( .IN0(n3145), .IN1(n3148), .SEL(n3146), .F(n3141) );
  MUX U3082 ( .IN0(n2782), .IN1(n2784), .SEL(n2783), .F(n374) );
  IV U3083 ( .A(n374), .Z(n1858) );
  MUX U3084 ( .IN0(n5266), .IN1(n5268), .SEL(n5267), .F(n375) );
  IV U3085 ( .A(n375), .Z(n4125) );
  MUX U3086 ( .IN0(n3930), .IN1(n376), .SEL(n3931), .F(n3451) );
  IV U3087 ( .A(n3932), .Z(n376) );
  XOR U3088 ( .A(n3197), .B(n3196), .Z(n3185) );
  MUX U3089 ( .IN0(n1139), .IN1(n377), .SEL(n1140), .F(n977) );
  IV U3090 ( .A(n1141), .Z(n377) );
  MUX U3091 ( .IN0(n1129), .IN1(n1131), .SEL(n1130), .F(n972) );
  XOR U3092 ( .A(n3104), .B(n3103), .Z(n3111) );
  MUX U3093 ( .IN0(n3130), .IN1(n378), .SEL(n3131), .F(n3065) );
  IV U3094 ( .A(n3132), .Z(n378) );
  MUX U3095 ( .IN0(n3061), .IN1(n3064), .SEL(n3062), .F(n3041) );
  MUX U3096 ( .IN0(n883), .IN1(n379), .SEL(n884), .F(n850) );
  IV U3097 ( .A(n885), .Z(n379) );
  XNOR U3098 ( .A(n956), .B(n957), .Z(n886) );
  MUX U3099 ( .IN0(n945), .IN1(n380), .SEL(n946), .F(n879) );
  IV U3100 ( .A(n947), .Z(n380) );
  XOR U3101 ( .A(n3092), .B(n3091), .Z(n3107) );
  XOR U3102 ( .A(n3045), .B(n3043), .Z(n3037) );
  MUX U3103 ( .IN0(n3019), .IN1(n3017), .SEL(n3018), .F(n381) );
  IV U3104 ( .A(n381), .Z(n1992) );
  XOR U3105 ( .A(n3550), .B(n3549), .Z(n1404) );
  MUX U3106 ( .IN0(n382), .IN1(n965), .SEL(n809), .F(n889) );
  IV U3107 ( .A(n810), .Z(n382) );
  MUX U3108 ( .IN0(n836), .IN1(n839), .SEL(n837), .F(n829) );
  MUX U3109 ( .IN0(n3032), .IN1(n383), .SEL(n834), .F(n3023) );
  IV U3110 ( .A(n833), .Z(n383) );
  MUX U3111 ( .IN0(n2775), .IN1(n2773), .SEL(n2774), .F(n384) );
  IV U3112 ( .A(n384), .Z(n1856) );
  MUX U3113 ( .IN0(n6261), .IN1(n6259), .SEL(n6260), .F(n385) );
  IV U3114 ( .A(n385), .Z(n4683) );
  MUX U3115 ( .IN0(n6143), .IN1(n6141), .SEL(n6142), .F(n386) );
  IV U3116 ( .A(n386), .Z(n4620) );
  MUX U3117 ( .IN0(n5796), .IN1(n5794), .SEL(n5795), .F(n387) );
  IV U3118 ( .A(n387), .Z(n4425) );
  MUX U3119 ( .IN0(n5680), .IN1(n5678), .SEL(n5679), .F(n388) );
  IV U3120 ( .A(n388), .Z(n4361) );
  MUX U3121 ( .IN0(n5100), .IN1(n5098), .SEL(n5099), .F(n4044) );
  MUX U3122 ( .IN0(n5058), .IN1(n5056), .SEL(n5057), .F(n4016) );
  MUX U3123 ( .IN0(n5082), .IN1(n5080), .SEL(n5081), .F(n5076) );
  MUX U3124 ( .IN0(n5086), .IN1(n5084), .SEL(n5085), .F(n389) );
  IV U3125 ( .A(n389), .Z(n4029) );
  MUX U3126 ( .IN0(n390), .IN1(n5194), .SEL(n5195), .F(n4085) );
  IV U3127 ( .A(n5196), .Z(n390) );
  MUX U3128 ( .IN0(n5163), .IN1(n5161), .SEL(n5162), .F(n391) );
  IV U3129 ( .A(n391), .Z(n4068) );
  MUX U3130 ( .IN0(n5241), .IN1(n5239), .SEL(n5240), .F(n5235) );
  MUX U3131 ( .IN0(n5245), .IN1(n5243), .SEL(n5244), .F(n4120) );
  MUX U3132 ( .IN0(n2804), .IN1(n2802), .SEL(n2803), .F(n392) );
  IV U3133 ( .A(n392), .Z(n1875) );
  MUX U3134 ( .IN0(n2620), .IN1(n2618), .SEL(n2619), .F(n1772) );
  MUX U3135 ( .IN0(n393), .IN1(n2569), .SEL(n2570), .F(n1735) );
  IV U3136 ( .A(n2571), .Z(n393) );
  MUX U3137 ( .IN0(n2581), .IN1(n2579), .SEL(n2580), .F(n394) );
  IV U3138 ( .A(n394), .Z(n1742) );
  MUX U3139 ( .IN0(n2602), .IN1(n2600), .SEL(n2601), .F(n2596) );
  MUX U3140 ( .IN0(n395), .IN1(n2610), .SEL(n2611), .F(n1760) );
  IV U3141 ( .A(n2612), .Z(n395) );
  MUX U3142 ( .IN0(n2676), .IN1(n2674), .SEL(n2675), .F(n1804) );
  MUX U3143 ( .IN0(n2747), .IN1(n2745), .SEL(n2746), .F(n1842) );
  MUX U3144 ( .IN0(n396), .IN1(n2738), .SEL(n2739), .F(n1831) );
  IV U3145 ( .A(n2740), .Z(n396) );
  MUX U3146 ( .IN0(n6828), .IN1(n6826), .SEL(n6827), .F(n5017) );
  MUX U3147 ( .IN0(n6786), .IN1(n6784), .SEL(n6785), .F(n4989) );
  MUX U3148 ( .IN0(n6807), .IN1(n6805), .SEL(n6806), .F(n397) );
  IV U3149 ( .A(n397), .Z(n4998) );
  MUX U3150 ( .IN0(n6814), .IN1(n6812), .SEL(n6813), .F(n398) );
  IV U3151 ( .A(n398), .Z(n5002) );
  MUX U3152 ( .IN0(n399), .IN1(n6693), .SEL(n6694), .F(n4927) );
  IV U3153 ( .A(n6695), .Z(n399) );
  MUX U3154 ( .IN0(n6717), .IN1(n6715), .SEL(n6716), .F(n400) );
  IV U3155 ( .A(n400), .Z(n4942) );
  MUX U3156 ( .IN0(n6483), .IN1(n6481), .SEL(n6482), .F(n4820) );
  MUX U3157 ( .IN0(n6439), .IN1(n6437), .SEL(n6438), .F(n4793) );
  MUX U3158 ( .IN0(n6589), .IN1(n6587), .SEL(n6588), .F(n401) );
  IV U3159 ( .A(n401), .Z(n4868) );
  MUX U3160 ( .IN0(n6550), .IN1(n6548), .SEL(n6549), .F(n402) );
  IV U3161 ( .A(n402), .Z(n4851) );
  MUX U3162 ( .IN0(n6617), .IN1(n6615), .SEL(n6616), .F(n403) );
  IV U3163 ( .A(n403), .Z(n4886) );
  MUX U3164 ( .IN0(n6638), .IN1(n6636), .SEL(n6637), .F(n6632) );
  MUX U3165 ( .IN0(n6185), .IN1(n6183), .SEL(n6184), .F(n4649) );
  MUX U3166 ( .IN0(n6094), .IN1(n6092), .SEL(n6093), .F(n4601) );
  MUX U3167 ( .IN0(n404), .IN1(n6001), .SEL(n6002), .F(n4540) );
  IV U3168 ( .A(n6003), .Z(n404) );
  MUX U3169 ( .IN0(n6038), .IN1(n6036), .SEL(n6037), .F(n4567) );
  MUX U3170 ( .IN0(n6299), .IN1(n6297), .SEL(n6298), .F(n4714) );
  MUX U3171 ( .IN0(n6219), .IN1(n6217), .SEL(n6218), .F(n405) );
  IV U3172 ( .A(n405), .Z(n4659) );
  MUX U3173 ( .IN0(n6240), .IN1(n6238), .SEL(n6239), .F(n6234) );
  MUX U3174 ( .IN0(n6365), .IN1(n6363), .SEL(n6364), .F(n6359) );
  MUX U3175 ( .IN0(n6386), .IN1(n6384), .SEL(n6385), .F(n406) );
  IV U3176 ( .A(n406), .Z(n4756) );
  MUX U3177 ( .IN0(n5445), .IN1(n5443), .SEL(n5444), .F(n4236) );
  MUX U3178 ( .IN0(n5403), .IN1(n5401), .SEL(n5402), .F(n4208) );
  MUX U3179 ( .IN0(n407), .IN1(n5394), .SEL(n5395), .F(n4197) );
  IV U3180 ( .A(n5396), .Z(n407) );
  MUX U3181 ( .IN0(n5424), .IN1(n5422), .SEL(n5423), .F(n408) );
  IV U3182 ( .A(n408), .Z(n4217) );
  MUX U3183 ( .IN0(n409), .IN1(n5435), .SEL(n5436), .F(n4222) );
  IV U3184 ( .A(n5437), .Z(n409) );
  MUX U3185 ( .IN0(n5319), .IN1(n5317), .SEL(n5318), .F(n4160) );
  XOR U3186 ( .A(n5302), .B(n5303), .Z(n4147) );
  MUX U3187 ( .IN0(n5347), .IN1(n5345), .SEL(n5346), .F(n4176) );
  MUX U3188 ( .IN0(n5722), .IN1(n5720), .SEL(n5721), .F(n4390) );
  MUX U3189 ( .IN0(n5631), .IN1(n5629), .SEL(n5630), .F(n4342) );
  MUX U3190 ( .IN0(n410), .IN1(n5538), .SEL(n5539), .F(n4279) );
  IV U3191 ( .A(n5540), .Z(n410) );
  MUX U3192 ( .IN0(n5585), .IN1(n5583), .SEL(n5584), .F(n5579) );
  MUX U3193 ( .IN0(n5848), .IN1(n5846), .SEL(n5847), .F(n5842) );
  MUX U3194 ( .IN0(n5754), .IN1(n5752), .SEL(n5753), .F(n411) );
  IV U3195 ( .A(n411), .Z(n4401) );
  MUX U3196 ( .IN0(n5768), .IN1(n5766), .SEL(n5767), .F(n412) );
  IV U3197 ( .A(n412), .Z(n4409) );
  MUX U3198 ( .IN0(n5898), .IN1(n5896), .SEL(n5897), .F(n4486) );
  XOR U3199 ( .A(n5881), .B(n5882), .Z(n4473) );
  XOR U3200 ( .A(n1925), .B(n1923), .Z(n1917) );
  MUX U3201 ( .IN0(n2713), .IN1(n2715), .SEL(n2714), .F(n413) );
  IV U3202 ( .A(n413), .Z(n1816) );
  MUX U3203 ( .IN0(n2655), .IN1(n2657), .SEL(n2656), .F(n414) );
  IV U3204 ( .A(n414), .Z(n1785) );
  MUX U3205 ( .IN0(n6349), .IN1(n6351), .SEL(n6350), .F(n415) );
  IV U3206 ( .A(n415), .Z(n4736) );
  XOR U3207 ( .A(n4703), .B(n4701), .Z(n4710) );
  XOR U3208 ( .A(n4581), .B(n4579), .Z(n4571) );
  XOR U3209 ( .A(n4556), .B(n4554), .Z(n4563) );
  MUX U3210 ( .IN0(n6004), .IN1(n6006), .SEL(n6005), .F(n416) );
  IV U3211 ( .A(n416), .Z(n4541) );
  XOR U3212 ( .A(n4638), .B(n4637), .Z(n4645) );
  MUX U3213 ( .IN0(n6696), .IN1(n6698), .SEL(n6697), .F(n417) );
  IV U3214 ( .A(n417), .Z(n4928) );
  MUX U3215 ( .IN0(n6522), .IN1(n6524), .SEL(n6523), .F(n418) );
  IV U3216 ( .A(n418), .Z(n4831) );
  XOR U3217 ( .A(n4443), .B(n4442), .Z(n4450) );
  XOR U3218 ( .A(n4320), .B(n4318), .Z(n4312) );
  XOR U3219 ( .A(n4295), .B(n4293), .Z(n4302) );
  MUX U3220 ( .IN0(n5541), .IN1(n5543), .SEL(n5542), .F(n419) );
  IV U3221 ( .A(n419), .Z(n4280) );
  XOR U3222 ( .A(n4379), .B(n4378), .Z(n4386) );
  MUX U3223 ( .IN0(n5482), .IN1(n5484), .SEL(n5483), .F(n420) );
  IV U3224 ( .A(n420), .Z(n4248) );
  XOR U3225 ( .A(n4101), .B(n4099), .Z(n4108) );
  MUX U3226 ( .IN0(n5139), .IN1(n5141), .SEL(n5140), .F(n421) );
  IV U3227 ( .A(n421), .Z(n4055) );
  MUX U3228 ( .IN0(n4006), .IN1(n422), .SEL(n4007), .F(n3488) );
  IV U3229 ( .A(n4008), .Z(n422) );
  MUX U3230 ( .IN0(n4979), .IN1(n423), .SEL(n4980), .F(n3968) );
  IV U3231 ( .A(n4981), .Z(n423) );
  MUX U3232 ( .IN0(n4045), .IN1(n4047), .SEL(n4046), .F(n3506) );
  MUX U3233 ( .IN0(n577), .IN1(n4096), .SEL(n4094), .F(n4089) );
  MUX U3234 ( .IN0(n3006), .IN1(n3004), .SEL(n3005), .F(n1991) );
  XOR U3235 ( .A(n2989), .B(n2990), .Z(n1978) );
  MUX U3236 ( .IN0(n2906), .IN1(n2904), .SEL(n2905), .F(n424) );
  IV U3237 ( .A(n424), .Z(n1933) );
  MUX U3238 ( .IN0(n2943), .IN1(n2941), .SEL(n2942), .F(n2937) );
  MUX U3239 ( .IN0(n2831), .IN1(n2829), .SEL(n2830), .F(n1895) );
  MUX U3240 ( .IN0(n2869), .IN1(n2867), .SEL(n2868), .F(n2863) );
  XOR U3241 ( .A(n1900), .B(n1898), .Z(n1907) );
  XOR U3242 ( .A(n1598), .B(n671), .Z(n2320) );
  MUX U3243 ( .IN0(n2243), .IN1(n2241), .SEL(n2242), .F(n425) );
  IV U3244 ( .A(n425), .Z(n1548) );
  MUX U3245 ( .IN0(n2264), .IN1(n2262), .SEL(n2263), .F(n2258) );
  MUX U3246 ( .IN0(n2156), .IN1(n2154), .SEL(n2155), .F(n1505) );
  XOR U3247 ( .A(n1518), .B(n681), .Z(n2181) );
  MUX U3248 ( .IN0(n2436), .IN1(n2434), .SEL(n2435), .F(n1665) );
  MUX U3249 ( .IN0(n2430), .IN1(n2432), .SEL(n2431), .F(n426) );
  IV U3250 ( .A(n426), .Z(n1656) );
  MUX U3251 ( .IN0(n2346), .IN1(n2348), .SEL(n2347), .F(n427) );
  IV U3252 ( .A(n427), .Z(n1607) );
  MUX U3253 ( .IN0(n2339), .IN1(n2337), .SEL(n2338), .F(n428) );
  IV U3254 ( .A(n428), .Z(n1605) );
  MUX U3255 ( .IN0(n2376), .IN1(n2374), .SEL(n2375), .F(n2370) );
  XOR U3256 ( .A(n1695), .B(n689), .Z(n2491) );
  XOR U3257 ( .A(n2463), .B(n2464), .Z(n1677) );
  MUX U3258 ( .IN0(n429), .IN1(n2513), .SEL(n2514), .F(n1702) );
  IV U3259 ( .A(n2515), .Z(n429) );
  MUX U3260 ( .IN0(n1773), .IN1(n1776), .SEL(n1774), .F(n1297) );
  MUX U3261 ( .IN0(n1805), .IN1(n1807), .SEL(n1806), .F(n1313) );
  MUX U3262 ( .IN0(n5018), .IN1(n5020), .SEL(n5019), .F(n3986) );
  MUX U3263 ( .IN0(n596), .IN1(n4938), .SEL(n4936), .F(n4931) );
  MUX U3264 ( .IN0(n475), .IN1(n4951), .SEL(n4950), .F(n430) );
  IV U3265 ( .A(n430), .Z(n3958) );
  MUX U3266 ( .IN0(n4821), .IN1(n4823), .SEL(n4822), .F(n3889) );
  MUX U3267 ( .IN0(n4780), .IN1(n4782), .SEL(n4781), .F(n3879) );
  MUX U3268 ( .IN0(n4853), .IN1(n4855), .SEL(n4854), .F(n3904) );
  MUX U3269 ( .IN0(n507), .IN1(n4866), .SEL(n4865), .F(n431) );
  IV U3270 ( .A(n431), .Z(n3909) );
  MUX U3271 ( .IN0(n612), .IN1(n4590), .SEL(n4588), .F(n3787) );
  MUX U3272 ( .IN0(n613), .IN1(n4551), .SEL(n4549), .F(n4544) );
  MUX U3273 ( .IN0(n622), .IN1(n4735), .SEL(n4733), .F(n3855) );
  MUX U3274 ( .IN0(n4237), .IN1(n4240), .SEL(n4238), .F(n3602) );
  MUX U3275 ( .IN0(n4140), .IN1(n4142), .SEL(n4141), .F(n3555) );
  MUX U3276 ( .IN0(n4150), .IN1(n432), .SEL(n4151), .F(n3560) );
  IV U3277 ( .A(n4152), .Z(n432) );
  MUX U3278 ( .IN0(n636), .IN1(n4165), .SEL(n4163), .F(n3574) );
  MUX U3279 ( .IN0(n641), .IN1(n4331), .SEL(n4329), .F(n3658) );
  MUX U3280 ( .IN0(n642), .IN1(n4290), .SEL(n4288), .F(n4283) );
  MUX U3281 ( .IN0(n4476), .IN1(n433), .SEL(n4477), .F(n3721) );
  IV U3282 ( .A(n4478), .Z(n433) );
  MUX U3283 ( .IN0(n653), .IN1(n4502), .SEL(n4500), .F(n4495) );
  XOR U3284 ( .A(n1718), .B(n1717), .Z(n1705) );
  XOR U3285 ( .A(n1672), .B(n1671), .Z(n1690) );
  XOR U3286 ( .A(n1524), .B(n1523), .Z(n1513) );
  XOR U3287 ( .A(n1478), .B(n1477), .Z(n1497) );
  XOR U3288 ( .A(n1574), .B(n1573), .Z(n1593) );
  MUX U3289 ( .IN0(n2984), .IN1(n2986), .SEL(n2985), .F(n434) );
  MUX U3290 ( .IN0(n6163), .IN1(n6165), .SEL(n6164), .F(n435) );
  IV U3291 ( .A(n435), .Z(n4632) );
  MUX U3292 ( .IN0(n6851), .IN1(n6853), .SEL(n6852), .F(n436) );
  XOR U3293 ( .A(n4799), .B(n4798), .Z(n4785) );
  MUX U3294 ( .IN0(n5700), .IN1(n5702), .SEL(n5701), .F(n437) );
  IV U3295 ( .A(n437), .Z(n4373) );
  XOR U3296 ( .A(n4180), .B(n4179), .Z(n4168) );
  MUX U3297 ( .IN0(n1777), .IN1(n438), .SEL(n1778), .F(n1298) );
  IV U3298 ( .A(n1779), .Z(n438) );
  MUX U3299 ( .IN0(n2001), .IN1(n1999), .SEL(n2000), .F(n439) );
  IV U3300 ( .A(n439), .Z(n1410) );
  XOR U3301 ( .A(n3619), .B(n3617), .Z(n3626) );
  XOR U3302 ( .A(n3522), .B(n3520), .Z(n3529) );
  MUX U3303 ( .IN0(n4241), .IN1(n440), .SEL(n4242), .F(n3603) );
  IV U3304 ( .A(n4243), .Z(n440) );
  XOR U3305 ( .A(n3882), .B(n3881), .Z(n3875) );
  XOR U3306 ( .A(n3748), .B(n3746), .Z(n3757) );
  MUX U3307 ( .IN0(n3514), .IN1(n3517), .SEL(n3515), .F(n3510) );
  MUX U3308 ( .IN0(n1972), .IN1(n1974), .SEL(n1973), .F(n1390) );
  MUX U3309 ( .IN0(n1981), .IN1(n441), .SEL(n1982), .F(n1395) );
  IV U3310 ( .A(n1983), .Z(n441) );
  MUX U3311 ( .IN0(n1939), .IN1(n442), .SEL(n1940), .F(n1378) );
  IV U3312 ( .A(n1941), .Z(n442) );
  MUX U3313 ( .IN0(n1956), .IN1(n1959), .SEL(n1957), .F(n1382) );
  XNOR U3314 ( .A(n1864), .B(n1865), .Z(n1341) );
  MUX U3315 ( .IN0(n1587), .IN1(n1590), .SEL(n1588), .F(n1213) );
  MUX U3316 ( .IN0(n1491), .IN1(n1494), .SEL(n1492), .F(n1166) );
  MUX U3317 ( .IN0(n521), .IN1(n1510), .SEL(n1508), .F(n1174) );
  MUX U3318 ( .IN0(n1652), .IN1(n1655), .SEL(n1653), .F(n1246) );
  MUX U3319 ( .IN0(n1611), .IN1(n443), .SEL(n1612), .F(n1223) );
  IV U3320 ( .A(n1613), .Z(n443) );
  MUX U3321 ( .IN0(n1628), .IN1(n1631), .SEL(n1629), .F(n1227) );
  MUX U3322 ( .IN0(n1648), .IN1(n444), .SEL(n1649), .F(n1236) );
  IV U3323 ( .A(n1650), .Z(n444) );
  MUX U3324 ( .IN0(n526), .IN1(n1687), .SEL(n1685), .F(n1261) );
  XNOR U3325 ( .A(n1668), .B(n1669), .Z(n1248) );
  MUX U3326 ( .IN0(n690), .IN1(n1713), .SEL(n1711), .F(n1706) );
  MUX U3327 ( .IN0(n1305), .IN1(n1308), .SEL(n1306), .F(n1301) );
  MUX U3328 ( .IN0(n1321), .IN1(n1324), .SEL(n1322), .F(n1317) );
  MUX U3329 ( .IN0(n3994), .IN1(n3997), .SEL(n3995), .F(n3990) );
  MUX U3330 ( .IN0(n3935), .IN1(n3938), .SEL(n3936), .F(n3462) );
  MUX U3331 ( .IN0(n3960), .IN1(n3962), .SEL(n3961), .F(n3465) );
  MUX U3332 ( .IN0(n3897), .IN1(n3900), .SEL(n3898), .F(n3893) );
  MUX U3333 ( .IN0(n3788), .IN1(n3790), .SEL(n3789), .F(n3382) );
  MUX U3334 ( .IN0(n3841), .IN1(n3844), .SEL(n3842), .F(n3417) );
  XNOR U3335 ( .A(n3857), .B(n3858), .Z(n3418) );
  MUX U3336 ( .IN0(n3610), .IN1(n3613), .SEL(n3611), .F(n3606) );
  MUX U3337 ( .IN0(n3659), .IN1(n3661), .SEL(n3660), .F(n3321) );
  XNOR U3338 ( .A(n3682), .B(n3683), .Z(n3334) );
  MUX U3339 ( .IN0(n3714), .IN1(n3716), .SEL(n3715), .F(n3357) );
  XOR U3340 ( .A(n2743), .B(n2742), .Z(n2701) );
  XOR U3341 ( .A(n5343), .B(n5342), .Z(n5299) );
  XOR U3342 ( .A(n6435), .B(n6434), .Z(n6508) );
  XOR U3343 ( .A(n6726), .B(n6725), .Z(n6682) );
  XOR U3344 ( .A(n6034), .B(n6033), .Z(n5990) );
  XOR U3345 ( .A(n1546), .B(n1545), .Z(n1585) );
  XOR U3346 ( .A(n4754), .B(n4753), .Z(n4730) );
  XOR U3347 ( .A(n4657), .B(n4656), .Z(n4698) );
  XOR U3348 ( .A(n4884), .B(n4883), .Z(n4858) );
  XOR U3349 ( .A(n4494), .B(n4493), .Z(n4471) );
  XOR U3350 ( .A(n4399), .B(n4398), .Z(n4439) );
  MUX U3351 ( .IN0(n1960), .IN1(n445), .SEL(n1961), .F(n1383) );
  IV U3352 ( .A(n1962), .Z(n445) );
  XOR U3353 ( .A(n1186), .B(n1185), .Z(n1205) );
  XOR U3354 ( .A(n3686), .B(n3685), .Z(n3704) );
  MUX U3355 ( .IN0(n4356), .IN1(n446), .SEL(n4357), .F(n3662) );
  IV U3356 ( .A(n4358), .Z(n446) );
  XOR U3357 ( .A(n3636), .B(n3635), .Z(n3622) );
  XOR U3358 ( .A(n3539), .B(n3538), .Z(n3525) );
  MUX U3359 ( .IN0(n4031), .IN1(n447), .SEL(n4032), .F(n3500) );
  IV U3360 ( .A(n4033), .Z(n447) );
  XOR U3361 ( .A(n3921), .B(n3920), .Z(n3907) );
  MUX U3362 ( .IN0(n5004), .IN1(n448), .SEL(n5005), .F(n3980) );
  IV U3363 ( .A(n5006), .Z(n448) );
  XOR U3364 ( .A(n3813), .B(n3812), .Z(n3831) );
  MUX U3365 ( .IN0(n4615), .IN1(n449), .SEL(n4616), .F(n3791) );
  IV U3366 ( .A(n4617), .Z(n449) );
  XOR U3367 ( .A(n3765), .B(n3764), .Z(n3753) );
  XOR U3368 ( .A(n1078), .B(n1076), .Z(n1070) );
  XOR U3369 ( .A(n1053), .B(n1051), .Z(n1062) );
  XOR U3370 ( .A(n3472), .B(n3471), .Z(n3479) );
  MUX U3371 ( .IN0(n3596), .IN1(n450), .SEL(n3597), .F(n3291) );
  IV U3372 ( .A(n3598), .Z(n450) );
  XOR U3373 ( .A(n3244), .B(n3243), .Z(n3251) );
  MUX U3374 ( .IN0(n451), .IN1(n2089), .SEL(n2090), .F(n1458) );
  IV U3375 ( .A(n2091), .Z(n451) );
  MUX U3376 ( .IN0(n2024), .IN1(n2022), .SEL(n2023), .F(n2018) );
  MUX U3377 ( .IN0(n1348), .IN1(n452), .SEL(n1349), .F(n1091) );
  IV U3378 ( .A(n1350), .Z(n452) );
  MUX U3379 ( .IN0(n1199), .IN1(n1202), .SEL(n1200), .F(n1016) );
  MUX U3380 ( .IN0(n1156), .IN1(n453), .SEL(n1157), .F(n987) );
  IV U3381 ( .A(n1158), .Z(n453) );
  MUX U3382 ( .IN0(n1232), .IN1(n1235), .SEL(n1233), .F(n1033) );
  MUX U3383 ( .IN0(n1251), .IN1(n454), .SEL(n1252), .F(n1035) );
  IV U3384 ( .A(n1253), .Z(n454) );
  MUX U3385 ( .IN0(n3390), .IN1(n3393), .SEL(n3391), .F(n3386) );
  MUX U3386 ( .IN0(n3406), .IN1(n3409), .SEL(n3407), .F(n3402) );
  MUX U3387 ( .IN0(n3288), .IN1(n3290), .SEL(n3289), .F(n3148) );
  MUX U3388 ( .IN0(n3329), .IN1(n3332), .SEL(n3330), .F(n3325) );
  MUX U3389 ( .IN0(n3344), .IN1(n3347), .SEL(n3345), .F(n3340) );
  XOR U3390 ( .A(n2138), .B(n2137), .Z(n2277) );
  XOR U3391 ( .A(n6568), .B(n6567), .Z(n6478) );
  XOR U3392 ( .A(n1810), .B(n1809), .Z(n1763) );
  XOR U3393 ( .A(n3719), .B(n3718), .Z(n3697) );
  XOR U3394 ( .A(n3847), .B(n3846), .Z(n3824) );
  MUX U3395 ( .IN0(n1368), .IN1(n455), .SEL(n1369), .F(n1096) );
  IV U3396 ( .A(n1370), .Z(n455) );
  XOR U3397 ( .A(n3367), .B(n3366), .Z(n3385) );
  XOR U3398 ( .A(n3306), .B(n3305), .Z(n3324) );
  XOR U3399 ( .A(n3259), .B(n3258), .Z(n3247) );
  MUX U3400 ( .IN0(n547), .IN1(n1471), .SEL(n1469), .F(n1462) );
  MUX U3401 ( .IN0(n1093), .IN1(n1095), .SEL(n1094), .F(n951) );
  MUX U3402 ( .IN0(n998), .IN1(n456), .SEL(n999), .F(n907) );
  IV U3403 ( .A(n1000), .Z(n456) );
  XNOR U3404 ( .A(n3208), .B(n3209), .Z(n3102) );
  MUX U3405 ( .IN0(n3134), .IN1(n3137), .SEL(n3135), .F(n3075) );
  XOR U3406 ( .A(n2390), .B(n2389), .Z(n2221) );
  XOR U3407 ( .A(n5095), .B(n5094), .Z(n5384) );
  XOR U3408 ( .A(n6253), .B(n6252), .Z(n6075) );
  MUX U3409 ( .IN0(n4904), .IN1(n457), .SEL(n4905), .F(n3930) );
  IV U3410 ( .A(n4906), .Z(n457) );
  MUX U3411 ( .IN0(n1135), .IN1(n1138), .SEL(n1136), .F(n983) );
  XOR U3412 ( .A(n3401), .B(n3400), .Z(n3378) );
  XOR U3413 ( .A(n3429), .B(n3428), .Z(n3468) );
  XOR U3414 ( .A(n3339), .B(n3338), .Z(n3317) );
  XOR U3415 ( .A(n3121), .B(n3120), .Z(n3140) );
  XOR U3416 ( .A(n3212), .B(n3211), .Z(n3230) );
  MUX U3417 ( .IN0(n961), .IN1(n964), .SEL(n962), .F(n955) );
  MUX U3418 ( .IN0(n911), .IN1(n458), .SEL(n912), .F(n865) );
  IV U3419 ( .A(n913), .Z(n458) );
  MUX U3420 ( .IN0(n919), .IN1(n459), .SEL(n920), .F(n869) );
  IV U3421 ( .A(n921), .Z(n459) );
  MUX U3422 ( .IN0(n875), .IN1(n878), .SEL(n876), .F(n851) );
  MUX U3423 ( .IN0(n3112), .IN1(n3115), .SEL(n3113), .F(n3108) );
  XOR U3424 ( .A(n5612), .B(n5611), .Z(n5268) );
  XOR U3425 ( .A(n1414), .B(n1413), .Z(n1454) );
  XOR U3426 ( .A(n1537), .B(n1536), .Z(n1860) );
  XOR U3427 ( .A(n1181), .B(n1180), .Z(n1338) );
  XOR U3428 ( .A(n1124), .B(n1123), .Z(n1141) );
  XOR U3429 ( .A(n3156), .B(n3155), .Z(n3132) );
  XOR U3430 ( .A(n3185), .B(n3184), .Z(n3222) );
  XOR U3431 ( .A(n862), .B(n861), .Z(n881) );
  MUX U3432 ( .IN0(n3047), .IN1(n3050), .SEL(n3048), .F(n3031) );
  XOR U3433 ( .A(n4127), .B(n4126), .Z(n1994) );
  MUX U3434 ( .IN0(n460), .IN1(n1115), .SEL(n811), .F(n965) );
  IV U3435 ( .A(n812), .Z(n460) );
  XOR U3436 ( .A(n3067), .B(n3066), .Z(n891) );
  XOR U3437 ( .A(n3037), .B(n3036), .Z(n854) );
  MUX U3438 ( .IN0(n840), .IN1(n461), .SEL(n841), .F(n830) );
  IV U3439 ( .A(n842), .Z(n461) );
  MUX U3440 ( .IN0(n462), .IN1(n820), .SEL(n801), .F(n817) );
  IV U3441 ( .A(n802), .Z(n462) );
  MUX U3442 ( .IN0(n2606), .IN1(n2604), .SEL(n2605), .F(n463) );
  IV U3443 ( .A(n463), .Z(n1759) );
  MUX U3444 ( .IN0(n5148), .IN1(n5146), .SEL(n5147), .F(n464) );
  IV U3445 ( .A(n464), .Z(n4059) );
  MUX U3446 ( .IN0(n5061), .IN1(n5059), .SEL(n5060), .F(n465) );
  IV U3447 ( .A(n465), .Z(n4010) );
  MUX U3448 ( .IN0(n5072), .IN1(n5070), .SEL(n5071), .F(n4026) );
  MUX U3449 ( .IN0(n5203), .IN1(n5201), .SEL(n5202), .F(n4096) );
  MUX U3450 ( .IN0(n5174), .IN1(n5172), .SEL(n5173), .F(n466) );
  IV U3451 ( .A(n466), .Z(n4077) );
  MUX U3452 ( .IN0(n5231), .IN1(n5229), .SEL(n5230), .F(n4112) );
  MUX U3453 ( .IN0(n5259), .IN1(n5257), .SEL(n5258), .F(n467) );
  IV U3454 ( .A(n467), .Z(n4123) );
  MUX U3455 ( .IN0(n2664), .IN1(n2662), .SEL(n2663), .F(n468) );
  IV U3456 ( .A(n468), .Z(n1789) );
  MUX U3457 ( .IN0(n2578), .IN1(n2576), .SEL(n2577), .F(n1748) );
  MUX U3458 ( .IN0(n2592), .IN1(n2590), .SEL(n2591), .F(n1756) );
  MUX U3459 ( .IN0(n2722), .IN1(n2720), .SEL(n2721), .F(n469) );
  IV U3460 ( .A(n469), .Z(n1820) );
  MUX U3461 ( .IN0(n2750), .IN1(n2748), .SEL(n2749), .F(n470) );
  IV U3462 ( .A(n470), .Z(n1836) );
  MUX U3463 ( .IN0(n6876), .IN1(n6874), .SEL(n6875), .F(n471) );
  IV U3464 ( .A(n471), .Z(n5031) );
  MUX U3465 ( .IN0(n6789), .IN1(n6787), .SEL(n6788), .F(n472) );
  IV U3466 ( .A(n472), .Z(n4983) );
  MUX U3467 ( .IN0(n6705), .IN1(n6703), .SEL(n6704), .F(n473) );
  IV U3468 ( .A(n473), .Z(n4932) );
  MUX U3469 ( .IN0(n6673), .IN1(n6671), .SEL(n6672), .F(n474) );
  IV U3470 ( .A(n474), .Z(n4919) );
  MUX U3471 ( .IN0(n6733), .IN1(n6731), .SEL(n6732), .F(n475) );
  MUX U3472 ( .IN0(n6744), .IN1(n6742), .SEL(n6743), .F(n4965) );
  MUX U3473 ( .IN0(n6758), .IN1(n6756), .SEL(n6757), .F(n476) );
  IV U3474 ( .A(n476), .Z(n4968) );
  MUX U3475 ( .IN0(n6531), .IN1(n6529), .SEL(n6530), .F(n477) );
  IV U3476 ( .A(n477), .Z(n4835) );
  MUX U3477 ( .IN0(n6442), .IN1(n6440), .SEL(n6441), .F(n478) );
  IV U3478 ( .A(n478), .Z(n4787) );
  MUX U3479 ( .IN0(n6453), .IN1(n6451), .SEL(n6452), .F(n4803) );
  MUX U3480 ( .IN0(n6586), .IN1(n6584), .SEL(n6585), .F(n4874) );
  MUX U3481 ( .IN0(n6614), .IN1(n6612), .SEL(n6613), .F(n4892) );
  MUX U3482 ( .IN0(n6628), .IN1(n6626), .SEL(n6627), .F(n4900) );
  MUX U3483 ( .IN0(n479), .IN1(n6648), .SEL(n6649), .F(n4903) );
  IV U3484 ( .A(n6650), .Z(n479) );
  MUX U3485 ( .IN0(n6188), .IN1(n6186), .SEL(n6187), .F(n480) );
  IV U3486 ( .A(n480), .Z(n4643) );
  MUX U3487 ( .IN0(n6097), .IN1(n6095), .SEL(n6096), .F(n481) );
  IV U3488 ( .A(n481), .Z(n4595) );
  MUX U3489 ( .IN0(n6013), .IN1(n6011), .SEL(n6012), .F(n482) );
  IV U3490 ( .A(n482), .Z(n4545) );
  MUX U3491 ( .IN0(n5967), .IN1(n5965), .SEL(n5966), .F(n4529) );
  MUX U3492 ( .IN0(n483), .IN1(n5985), .SEL(n5986), .F(n4533) );
  IV U3493 ( .A(n5987), .Z(n483) );
  MUX U3494 ( .IN0(n6041), .IN1(n6039), .SEL(n6040), .F(n484) );
  IV U3495 ( .A(n484), .Z(n4561) );
  MUX U3496 ( .IN0(n6059), .IN1(n6057), .SEL(n6058), .F(n485) );
  IV U3497 ( .A(n485), .Z(n4576) );
  MUX U3498 ( .IN0(n6066), .IN1(n6064), .SEL(n6065), .F(n486) );
  IV U3499 ( .A(n486), .Z(n4580) );
  MUX U3500 ( .IN0(n6302), .IN1(n6300), .SEL(n6301), .F(n487) );
  IV U3501 ( .A(n487), .Z(n4708) );
  MUX U3502 ( .IN0(n6216), .IN1(n6214), .SEL(n6215), .F(n4665) );
  MUX U3503 ( .IN0(n6230), .IN1(n6228), .SEL(n6229), .F(n4673) );
  MUX U3504 ( .IN0(n488), .IN1(n6248), .SEL(n6249), .F(n4677) );
  IV U3505 ( .A(n6250), .Z(n488) );
  MUX U3506 ( .IN0(n6355), .IN1(n6353), .SEL(n6354), .F(n4746) );
  MUX U3507 ( .IN0(n6383), .IN1(n6381), .SEL(n6382), .F(n4762) );
  MUX U3508 ( .IN0(n6397), .IN1(n6395), .SEL(n6396), .F(n4772) );
  MUX U3509 ( .IN0(n5491), .IN1(n5489), .SEL(n5490), .F(n489) );
  IV U3510 ( .A(n489), .Z(n4252) );
  MUX U3511 ( .IN0(n5406), .IN1(n5404), .SEL(n5405), .F(n490) );
  IV U3512 ( .A(n490), .Z(n4202) );
  MUX U3513 ( .IN0(n5322), .IN1(n5320), .SEL(n5321), .F(n491) );
  IV U3514 ( .A(n491), .Z(n4154) );
  MUX U3515 ( .IN0(n5350), .IN1(n5348), .SEL(n5349), .F(n492) );
  IV U3516 ( .A(n492), .Z(n4170) );
  MUX U3517 ( .IN0(n5368), .IN1(n5366), .SEL(n5367), .F(n493) );
  IV U3518 ( .A(n493), .Z(n4183) );
  MUX U3519 ( .IN0(n5375), .IN1(n5373), .SEL(n5374), .F(n494) );
  IV U3520 ( .A(n494), .Z(n4187) );
  MUX U3521 ( .IN0(n5725), .IN1(n5723), .SEL(n5724), .F(n495) );
  IV U3522 ( .A(n495), .Z(n4384) );
  MUX U3523 ( .IN0(n5634), .IN1(n5632), .SEL(n5633), .F(n496) );
  IV U3524 ( .A(n496), .Z(n4336) );
  MUX U3525 ( .IN0(n5550), .IN1(n5548), .SEL(n5549), .F(n497) );
  IV U3526 ( .A(n497), .Z(n4284) );
  MUX U3527 ( .IN0(n5518), .IN1(n5516), .SEL(n5517), .F(n498) );
  IV U3528 ( .A(n498), .Z(n4271) );
  MUX U3529 ( .IN0(n5575), .IN1(n5573), .SEL(n5574), .F(n4306) );
  MUX U3530 ( .IN0(n5596), .IN1(n5594), .SEL(n5595), .F(n499) );
  IV U3531 ( .A(n499), .Z(n4315) );
  MUX U3532 ( .IN0(n5603), .IN1(n5601), .SEL(n5602), .F(n500) );
  IV U3533 ( .A(n500), .Z(n4319) );
  MUX U3534 ( .IN0(n5838), .IN1(n5836), .SEL(n5837), .F(n4454) );
  MUX U3535 ( .IN0(n5751), .IN1(n5749), .SEL(n5750), .F(n4407) );
  MUX U3536 ( .IN0(n5772), .IN1(n5770), .SEL(n5771), .F(n501) );
  IV U3537 ( .A(n501), .Z(n4414) );
  MUX U3538 ( .IN0(n502), .IN1(n5783), .SEL(n5784), .F(n4419) );
  IV U3539 ( .A(n5785), .Z(n502) );
  MUX U3540 ( .IN0(n5901), .IN1(n5899), .SEL(n5900), .F(n503) );
  IV U3541 ( .A(n503), .Z(n4480) );
  MUX U3542 ( .IN0(n5929), .IN1(n5927), .SEL(n5928), .F(n504) );
  IV U3543 ( .A(n504), .Z(n4496) );
  MUX U3544 ( .IN0(n5947), .IN1(n5945), .SEL(n5946), .F(n505) );
  IV U3545 ( .A(n505), .Z(n4513) );
  MUX U3546 ( .IN0(n5954), .IN1(n5952), .SEL(n5953), .F(n506) );
  IV U3547 ( .A(n506), .Z(n4517) );
  XOR U3548 ( .A(n4776), .B(n4774), .Z(n4768) );
  XOR U3549 ( .A(n4751), .B(n4749), .Z(n4758) );
  XOR U3550 ( .A(n4735), .B(n4733), .Z(n4742) );
  XOR U3551 ( .A(n4654), .B(n4653), .Z(n4661) );
  XOR U3552 ( .A(n4879), .B(n4877), .Z(n4888) );
  MUX U3553 ( .IN0(n6580), .IN1(n6582), .SEL(n6581), .F(n507) );
  IV U3554 ( .A(n507), .Z(n4864) );
  MUX U3555 ( .IN0(n5832), .IN1(n5834), .SEL(n5833), .F(n508) );
  IV U3556 ( .A(n508), .Z(n4444) );
  XOR U3557 ( .A(n4396), .B(n4394), .Z(n4403) );
  MUX U3558 ( .IN0(n5225), .IN1(n5227), .SEL(n5226), .F(n509) );
  IV U3559 ( .A(n509), .Z(n4102) );
  MUX U3560 ( .IN0(n5197), .IN1(n5199), .SEL(n5198), .F(n510) );
  IV U3561 ( .A(n510), .Z(n4086) );
  MUX U3562 ( .IN0(n4052), .IN1(n4054), .SEL(n4053), .F(n3517) );
  MUX U3563 ( .IN0(n4083), .IN1(n4085), .SEL(n4084), .F(n3533) );
  MUX U3564 ( .IN0(n4068), .IN1(n511), .SEL(n4069), .F(n3521) );
  IV U3565 ( .A(n4070), .Z(n511) );
  MUX U3566 ( .IN0(n580), .IN1(n4101), .SEL(n4099), .F(n3543) );
  MUX U3567 ( .IN0(n4114), .IN1(n512), .SEL(n4115), .F(n3546) );
  IV U3568 ( .A(n4116), .Z(n512) );
  MUX U3569 ( .IN0(n3009), .IN1(n3007), .SEL(n3008), .F(n513) );
  IV U3570 ( .A(n513), .Z(n1985) );
  MUX U3571 ( .IN0(n2919), .IN1(n2917), .SEL(n2918), .F(n1945) );
  XOR U3572 ( .A(n1934), .B(n1932), .Z(n1941) );
  XOR U3573 ( .A(n1959), .B(n1957), .Z(n1951) );
  MUX U3574 ( .IN0(n2933), .IN1(n2931), .SEL(n2932), .F(n1955) );
  MUX U3575 ( .IN0(n2834), .IN1(n2832), .SEL(n2833), .F(n514) );
  IV U3576 ( .A(n514), .Z(n1889) );
  MUX U3577 ( .IN0(n2797), .IN1(n2795), .SEL(n2796), .F(n515) );
  IV U3578 ( .A(n515), .Z(n1871) );
  MUX U3579 ( .IN0(n2859), .IN1(n2857), .SEL(n2858), .F(n1911) );
  MUX U3580 ( .IN0(n2882), .IN1(n2880), .SEL(n2881), .F(n516) );
  IV U3581 ( .A(n516), .Z(n1920) );
  MUX U3582 ( .IN0(n2330), .IN1(n2328), .SEL(n2329), .F(n517) );
  IV U3583 ( .A(n517), .Z(n1599) );
  XOR U3584 ( .A(n1582), .B(n1580), .Z(n1574) );
  MUX U3585 ( .IN0(n2282), .IN1(n2280), .SEL(n2281), .F(n1578) );
  MUX U3586 ( .IN0(n2240), .IN1(n2238), .SEL(n2239), .F(n1554) );
  XOR U3587 ( .A(n1543), .B(n1541), .Z(n1550) );
  XOR U3588 ( .A(n1566), .B(n1564), .Z(n1558) );
  MUX U3589 ( .IN0(n2254), .IN1(n2252), .SEL(n2253), .F(n1562) );
  MUX U3590 ( .IN0(n2159), .IN1(n2157), .SEL(n2158), .F(n518) );
  IV U3591 ( .A(n518), .Z(n1499) );
  MUX U3592 ( .IN0(n2115), .IN1(n2113), .SEL(n2114), .F(n1482) );
  MUX U3593 ( .IN0(n2129), .IN1(n2127), .SEL(n2128), .F(n519) );
  IV U3594 ( .A(n519), .Z(n1485) );
  MUX U3595 ( .IN0(n2191), .IN1(n2189), .SEL(n2190), .F(n520) );
  IV U3596 ( .A(n520), .Z(n1519) );
  MUX U3597 ( .IN0(n2171), .IN1(n2169), .SEL(n2170), .F(n521) );
  IV U3598 ( .A(n521), .Z(n1509) );
  MUX U3599 ( .IN0(n2212), .IN1(n2210), .SEL(n2211), .F(n522) );
  IV U3600 ( .A(n522), .Z(n1533) );
  MUX U3601 ( .IN0(n2443), .IN1(n2441), .SEL(n2442), .F(n523) );
  IV U3602 ( .A(n523), .Z(n1664) );
  XOR U3603 ( .A(n1647), .B(n1645), .Z(n1639) );
  MUX U3604 ( .IN0(n2395), .IN1(n2393), .SEL(n2394), .F(n1643) );
  MUX U3605 ( .IN0(n2352), .IN1(n2350), .SEL(n2351), .F(n1617) );
  MUX U3606 ( .IN0(n524), .IN1(n2343), .SEL(n2344), .F(n1606) );
  IV U3607 ( .A(n2345), .Z(n524) );
  MUX U3608 ( .IN0(n2366), .IN1(n2364), .SEL(n2365), .F(n1627) );
  MUX U3609 ( .IN0(n2384), .IN1(n2382), .SEL(n2383), .F(n2378) );
  MUX U3610 ( .IN0(n2501), .IN1(n2499), .SEL(n2500), .F(n525) );
  IV U3611 ( .A(n525), .Z(n1696) );
  MUX U3612 ( .IN0(n2481), .IN1(n2479), .SEL(n2480), .F(n526) );
  IV U3613 ( .A(n526), .Z(n1686) );
  MUX U3614 ( .IN0(n2458), .IN1(n2456), .SEL(n2457), .F(n527) );
  IV U3615 ( .A(n527), .Z(n1675) );
  MUX U3616 ( .IN0(n2488), .IN1(n2490), .SEL(n2489), .F(n528) );
  IV U3617 ( .A(n528), .Z(n1688) );
  MUX U3618 ( .IN0(n2525), .IN1(n2523), .SEL(n2524), .F(n529) );
  IV U3619 ( .A(n529), .Z(n1707) );
  MUX U3620 ( .IN0(n2536), .IN1(n2534), .SEL(n2535), .F(n1722) );
  MUX U3621 ( .IN0(n1785), .IN1(n530), .SEL(n1786), .F(n1302) );
  IV U3622 ( .A(n1787), .Z(n530) );
  MUX U3623 ( .IN0(n1816), .IN1(n531), .SEL(n1817), .F(n1318) );
  IV U3624 ( .A(n1818), .Z(n531) );
  MUX U3625 ( .IN0(n590), .IN1(n1831), .SEL(n1829), .F(n1332) );
  MUX U3626 ( .IN0(n5024), .IN1(n5026), .SEL(n5025), .F(n3997) );
  MUX U3627 ( .IN0(n4925), .IN1(n4927), .SEL(n4926), .F(n3949) );
  MUX U3628 ( .IN0(n4828), .IN1(n4830), .SEL(n4829), .F(n3900) );
  MUX U3629 ( .IN0(n605), .IN1(n4863), .SEL(n4861), .F(n3915) );
  MUX U3630 ( .IN0(n4636), .IN1(n4638), .SEL(n4637), .F(n3808) );
  MUX U3631 ( .IN0(n4538), .IN1(n4540), .SEL(n4539), .F(n3761) );
  MUX U3632 ( .IN0(n616), .IN1(n4556), .SEL(n4554), .F(n3769) );
  MUX U3633 ( .IN0(n4569), .IN1(n532), .SEL(n4570), .F(n3772) );
  IV U3634 ( .A(n4571), .Z(n532) );
  MUX U3635 ( .IN0(n4704), .IN1(n533), .SEL(n4705), .F(n3833) );
  IV U3636 ( .A(n4706), .Z(n533) );
  MUX U3637 ( .IN0(n4717), .IN1(n534), .SEL(n4718), .F(n3843) );
  IV U3638 ( .A(n4719), .Z(n534) );
  MUX U3639 ( .IN0(n4245), .IN1(n4247), .SEL(n4246), .F(n3613) );
  MUX U3640 ( .IN0(n4147), .IN1(n4149), .SEL(n4148), .F(n3566) );
  MUX U3641 ( .IN0(n4377), .IN1(n4379), .SEL(n4378), .F(n3679) );
  MUX U3642 ( .IN0(n4277), .IN1(n4279), .SEL(n4278), .F(n3630) );
  MUX U3643 ( .IN0(n645), .IN1(n4295), .SEL(n4293), .F(n3640) );
  MUX U3644 ( .IN0(n4441), .IN1(n4443), .SEL(n4442), .F(n3712) );
  MUX U3645 ( .IN0(n4473), .IN1(n4475), .SEL(n4474), .F(n3727) );
  MUX U3646 ( .IN0(n654), .IN1(n4491), .SEL(n4489), .F(n3737) );
  MUX U3647 ( .IN0(n2136), .IN1(n2138), .SEL(n2137), .F(n535) );
  IV U3648 ( .A(n535), .Z(n1487) );
  XOR U3649 ( .A(n1967), .B(n1966), .Z(n1983) );
  MUX U3650 ( .IN0(n6279), .IN1(n6281), .SEL(n6280), .F(n536) );
  IV U3651 ( .A(n536), .Z(n4696) );
  XOR U3652 ( .A(n4624), .B(n4623), .Z(n4641) );
  XOR U3653 ( .A(n4912), .B(n4911), .Z(n4930) );
  XOR U3654 ( .A(n5013), .B(n5012), .Z(n5029) );
  XOR U3655 ( .A(n4816), .B(n4815), .Z(n4833) );
  XOR U3656 ( .A(n4508), .B(n4507), .Z(n4494) );
  XOR U3657 ( .A(n4461), .B(n4460), .Z(n4478) );
  XOR U3658 ( .A(n4312), .B(n4311), .Z(n4298) );
  XOR U3659 ( .A(n4264), .B(n4263), .Z(n4282) );
  XOR U3660 ( .A(n4365), .B(n4364), .Z(n4382) );
  XOR U3661 ( .A(n4135), .B(n4134), .Z(n4152) );
  XOR U3662 ( .A(n4232), .B(n4231), .Z(n4250) );
  XOR U3663 ( .A(n4040), .B(n4039), .Z(n4057) );
  XOR U3664 ( .A(n3716), .B(n3715), .Z(n3723) );
  MUX U3665 ( .IN0(n4437), .IN1(n537), .SEL(n4438), .F(n3702) );
  IV U3666 ( .A(n4439), .Z(n537) );
  MUX U3667 ( .IN0(n3504), .IN1(n3506), .SEL(n3505), .F(n3255) );
  MUX U3668 ( .IN0(n1978), .IN1(n1980), .SEL(n1979), .F(n1401) );
  XOR U3669 ( .A(n1390), .B(n1388), .Z(n1397) );
  MUX U3670 ( .IN0(n1873), .IN1(n1876), .SEL(n1874), .F(n1343) );
  MUX U3671 ( .IN0(n1885), .IN1(n538), .SEL(n1886), .F(n1348) );
  IV U3672 ( .A(n1887), .Z(n538) );
  MUX U3673 ( .IN0(n670), .IN1(n1900), .SEL(n1898), .F(n1364) );
  MUX U3674 ( .IN0(n1922), .IN1(n1925), .SEL(n1923), .F(n1367) );
  MUX U3675 ( .IN0(n671), .IN1(n1596), .SEL(n1595), .F(n539) );
  IV U3676 ( .A(n539), .Z(n1212) );
  MUX U3677 ( .IN0(n1495), .IN1(n540), .SEL(n1496), .F(n1160) );
  IV U3678 ( .A(n1497), .Z(n540) );
  MUX U3679 ( .IN0(n681), .IN1(n1516), .SEL(n1515), .F(n541) );
  IV U3680 ( .A(n541), .Z(n1173) );
  MUX U3681 ( .IN0(n1522), .IN1(n542), .SEL(n1523), .F(n1177) );
  IV U3682 ( .A(n1524), .Z(n542) );
  MUX U3683 ( .IN0(n683), .IN1(n1661), .SEL(n1660), .F(n543) );
  IV U3684 ( .A(n543), .Z(n1245) );
  MUX U3685 ( .IN0(n689), .IN1(n1693), .SEL(n1692), .F(n544) );
  IV U3686 ( .A(n544), .Z(n1260) );
  MUX U3687 ( .IN0(n1677), .IN1(n1679), .SEL(n1678), .F(n1250) );
  MUX U3688 ( .IN0(n691), .IN1(n1702), .SEL(n1700), .F(n1269) );
  MUX U3689 ( .IN0(n693), .IN1(n1726), .SEL(n1724), .F(n1273) );
  MUX U3690 ( .IN0(n1294), .IN1(n1297), .SEL(n1295), .F(n1066) );
  MUX U3691 ( .IN0(n1310), .IN1(n1313), .SEL(n1311), .F(n1074) );
  MUX U3692 ( .IN0(n1333), .IN1(n1335), .SEL(n1334), .F(n1078) );
  MUX U3693 ( .IN0(n3984), .IN1(n3986), .SEL(n3985), .F(n3483) );
  MUX U3694 ( .IN0(n3887), .IN1(n3889), .SEL(n3888), .F(n3437) );
  MUX U3695 ( .IN0(n3902), .IN1(n3904), .SEL(n3903), .F(n3447) );
  MUX U3696 ( .IN0(n3795), .IN1(n3797), .SEL(n3796), .F(n3393) );
  MUX U3697 ( .IN0(n3826), .IN1(n3828), .SEL(n3827), .F(n3409) );
  MUX U3698 ( .IN0(n3849), .IN1(n545), .SEL(n3850), .F(n3416) );
  IV U3699 ( .A(n3851), .Z(n545) );
  MUX U3700 ( .IN0(n3600), .IN1(n3602), .SEL(n3601), .F(n3301) );
  MUX U3701 ( .IN0(n3553), .IN1(n3555), .SEL(n3554), .F(n3279) );
  MUX U3702 ( .IN0(n3666), .IN1(n3668), .SEL(n3667), .F(n3332) );
  MUX U3703 ( .IN0(n3699), .IN1(n3701), .SEL(n3700), .F(n3347) );
  XOR U3704 ( .A(n2574), .B(n2573), .Z(n2643) );
  XOR U3705 ( .A(n2855), .B(n2854), .Z(n2813) );
  XOR U3706 ( .A(n2348), .B(n2347), .Z(n2418) );
  XOR U3707 ( .A(n2236), .B(n2235), .Z(n2305) );
  XOR U3708 ( .A(n5571), .B(n5570), .Z(n5527) );
  XOR U3709 ( .A(n1705), .B(n1704), .Z(n1682) );
  XOR U3710 ( .A(n1903), .B(n1902), .Z(n1879) );
  XOR U3711 ( .A(n1834), .B(n1833), .Z(n1810) );
  XOR U3712 ( .A(n1740), .B(n1739), .Z(n1779) );
  XOR U3713 ( .A(n4593), .B(n4592), .Z(n4634) );
  XOR U3714 ( .A(n4948), .B(n4947), .Z(n4923) );
  XOR U3715 ( .A(n4981), .B(n4980), .Z(n5022) );
  XOR U3716 ( .A(n4785), .B(n4784), .Z(n4826) );
  XOR U3717 ( .A(n4334), .B(n4333), .Z(n4375) );
  XOR U3718 ( .A(n4168), .B(n4167), .Z(n4145) );
  XOR U3719 ( .A(n4200), .B(n4199), .Z(n4243) );
  XOR U3720 ( .A(n4008), .B(n4007), .Z(n4050) );
  XOR U3721 ( .A(n1281), .B(n1280), .Z(n1300) );
  XOR U3722 ( .A(n3654), .B(n3653), .Z(n3671) );
  XOR U3723 ( .A(n3492), .B(n3491), .Z(n3509) );
  XOR U3724 ( .A(n3588), .B(n3587), .Z(n3605) );
  XOR U3725 ( .A(n3875), .B(n3874), .Z(n3892) );
  XOR U3726 ( .A(n3972), .B(n3971), .Z(n3989) );
  XOR U3727 ( .A(n3783), .B(n3782), .Z(n3800) );
  MUX U3728 ( .IN0(n1383), .IN1(n546), .SEL(n1384), .F(n1104) );
  IV U3729 ( .A(n1385), .Z(n546) );
  XOR U3730 ( .A(n3450), .B(n3449), .Z(n3443) );
  XOR U3731 ( .A(n3426), .B(n3424), .Z(n3433) );
  XOR U3732 ( .A(n3283), .B(n3281), .Z(n3275) );
  XOR U3733 ( .A(n3290), .B(n3289), .Z(n3297) );
  MUX U3734 ( .IN0(n2105), .IN1(n2103), .SEL(n2104), .F(n547) );
  IV U3735 ( .A(n547), .Z(n1470) );
  MUX U3736 ( .IN0(n2014), .IN1(n2012), .SEL(n2013), .F(n1422) );
  MUX U3737 ( .IN0(n2031), .IN1(n2029), .SEL(n2030), .F(n548) );
  IV U3738 ( .A(n548), .Z(n1424) );
  MUX U3739 ( .IN0(n3242), .IN1(n3244), .SEL(n3243), .F(n3125) );
  MUX U3740 ( .IN0(n1373), .IN1(n549), .SEL(n1374), .F(n1102) );
  IV U3741 ( .A(n1375), .Z(n549) );
  MUX U3742 ( .IN0(n1207), .IN1(n550), .SEL(n1208), .F(n1015) );
  IV U3743 ( .A(n1209), .Z(n550) );
  MUX U3744 ( .IN0(n1184), .IN1(n551), .SEL(n1185), .F(n1004) );
  IV U3745 ( .A(n1186), .Z(n551) );
  MUX U3746 ( .IN0(n1240), .IN1(n552), .SEL(n1241), .F(n1032) );
  IV U3747 ( .A(n1242), .Z(n552) );
  XNOR U3748 ( .A(n1216), .B(n1217), .Z(n1018) );
  MUX U3749 ( .IN0(n3470), .IN1(n3472), .SEL(n3471), .F(n3238) );
  MUX U3750 ( .IN0(n3380), .IN1(n3382), .SEL(n3381), .F(n3193) );
  MUX U3751 ( .IN0(n3395), .IN1(n3398), .SEL(n3396), .F(n3201) );
  MUX U3752 ( .IN0(n3418), .IN1(n3420), .SEL(n3419), .F(n3205) );
  MUX U3753 ( .IN0(n3319), .IN1(n3321), .SEL(n3320), .F(n3164) );
  MUX U3754 ( .IN0(n3334), .IN1(n3336), .SEL(n3335), .F(n3172) );
  XOR U3755 ( .A(n2701), .B(n2700), .Z(n2615) );
  XOR U3756 ( .A(n5878), .B(n5877), .Z(n5788) );
  XOR U3757 ( .A(n6337), .B(n6336), .Z(n6253) );
  XOR U3758 ( .A(n5990), .B(n5989), .Z(n6135) );
  MUX U3759 ( .IN0(n2092), .IN1(n2094), .SEL(n2093), .F(n553) );
  IV U3760 ( .A(n553), .Z(n1459) );
  XOR U3761 ( .A(n1411), .B(n1409), .Z(n1418) );
  MUX U3762 ( .IN0(n2219), .IN1(n2221), .SEL(n2220), .F(n554) );
  IV U3763 ( .A(n554), .Z(n1535) );
  XOR U3764 ( .A(n4536), .B(n4535), .Z(n4617) );
  MUX U3765 ( .IN0(n6765), .IN1(n6767), .SEL(n6766), .F(n555) );
  IV U3766 ( .A(n555), .Z(n4970) );
  XOR U3767 ( .A(n4858), .B(n4857), .Z(n4809) );
  MUX U3768 ( .IN0(n5382), .IN1(n5384), .SEL(n5383), .F(n556) );
  IV U3769 ( .A(n556), .Z(n4189) );
  XOR U3770 ( .A(n4081), .B(n4080), .Z(n4033) );
  XOR U3771 ( .A(n1316), .B(n1315), .Z(n1292) );
  XOR U3772 ( .A(n1158), .B(n1157), .Z(n1197) );
  XOR U3773 ( .A(n3622), .B(n3621), .Z(n3664) );
  XOR U3774 ( .A(n3525), .B(n3524), .Z(n3502) );
  XOR U3775 ( .A(n3558), .B(n3557), .Z(n3598) );
  XOR U3776 ( .A(n3907), .B(n3906), .Z(n3885) );
  XOR U3777 ( .A(n3941), .B(n3940), .Z(n3982) );
  XOR U3778 ( .A(n3753), .B(n3752), .Z(n3793) );
  XOR U3779 ( .A(n3458), .B(n3457), .Z(n3475) );
  MUX U3780 ( .IN0(n1096), .IN1(n557), .SEL(n1097), .F(n952) );
  IV U3781 ( .A(n1098), .Z(n557) );
  XOR U3782 ( .A(n3176), .B(n3174), .Z(n3168) );
  XOR U3783 ( .A(n3153), .B(n3151), .Z(n3160) );
  XOR U3784 ( .A(n3182), .B(n3180), .Z(n3189) );
  MUX U3785 ( .IN0(n1456), .IN1(n1458), .SEL(n1457), .F(n1148) );
  MUX U3786 ( .IN0(n3126), .IN1(n3129), .SEL(n3127), .F(n3064) );
  MUX U3787 ( .IN0(n1108), .IN1(n558), .SEL(n1109), .F(n963) );
  IV U3788 ( .A(n1110), .Z(n558) );
  MUX U3789 ( .IN0(n1010), .IN1(n559), .SEL(n1011), .F(n916) );
  IV U3790 ( .A(n1012), .Z(n559) );
  XOR U3791 ( .A(n906), .B(n904), .Z(n913) );
  XOR U3792 ( .A(n929), .B(n927), .Z(n921) );
  MUX U3793 ( .IN0(n1027), .IN1(n560), .SEL(n1028), .F(n924) );
  IV U3794 ( .A(n1029), .Z(n560) );
  MUX U3795 ( .IN0(n3228), .IN1(n561), .SEL(n3229), .F(n3109) );
  IV U3796 ( .A(n3230), .Z(n561) );
  XOR U3797 ( .A(n4680), .B(n4679), .Z(n4584) );
  MUX U3798 ( .IN0(n1858), .IN1(n562), .SEL(n1859), .F(n1336) );
  IV U3799 ( .A(n1860), .Z(n562) );
  XOR U3800 ( .A(n1230), .B(n1229), .Z(n1181) );
  XOR U3801 ( .A(n1131), .B(n1130), .Z(n1124) );
  XOR U3802 ( .A(n1138), .B(n1136), .Z(n1145) );
  XOR U3803 ( .A(n3697), .B(n3696), .Z(n3647) );
  XOR U3804 ( .A(n3824), .B(n3823), .Z(n3776) );
  XOR U3805 ( .A(n3247), .B(n3246), .Z(n3286) );
  MUX U3806 ( .IN0(n3451), .IN1(n563), .SEL(n3452), .F(n3220) );
  IV U3807 ( .A(n3453), .Z(n563) );
  XOR U3808 ( .A(n878), .B(n876), .Z(n885) );
  MUX U3809 ( .IN0(n949), .IN1(n951), .SEL(n950), .F(n888) );
  MUX U3810 ( .IN0(n3102), .IN1(n3104), .SEL(n3103), .F(n3058) );
  MUX U3811 ( .IN0(n3072), .IN1(n3075), .SEL(n3073), .F(n3068) );
  MUX U3812 ( .IN0(n564), .IN1(n2049), .SEL(n2558), .F(n1727) );
  IV U3813 ( .A(n2557), .Z(n564) );
  MUX U3814 ( .IN0(n6884), .IN1(n6886), .SEL(n6885), .F(n565) );
  IV U3815 ( .A(n565), .Z(n5038) );
  XOR U3816 ( .A(n4325), .B(n4324), .Z(n4127) );
  XOR U3817 ( .A(n1000), .B(n999), .Z(n1081) );
  XOR U3818 ( .A(n3317), .B(n3316), .Z(n3270) );
  MUX U3819 ( .IN0(n977), .IN1(n566), .SEL(n978), .F(n894) );
  IV U3820 ( .A(n979), .Z(n566) );
  MUX U3821 ( .IN0(n930), .IN1(n900), .SEL(n931), .F(n871) );
  MUX U3822 ( .IN0(n3239), .IN1(n567), .SEL(n968), .F(n3116) );
  IV U3823 ( .A(n967), .Z(n567) );
  XOR U3824 ( .A(n3079), .B(n3078), .Z(n3067) );
  XOR U3825 ( .A(n3050), .B(n3048), .Z(n3054) );
  MUX U3826 ( .IN0(n860), .IN1(n568), .SEL(n861), .F(n838) );
  IV U3827 ( .A(n862), .Z(n568) );
  MUX U3828 ( .IN0(n569), .IN1(n1402), .SEL(n813), .F(n1115) );
  IV U3829 ( .A(n814), .Z(n569) );
  MUX U3830 ( .IN0(n570), .IN1(n852), .SEL(n805), .F(n831) );
  IV U3831 ( .A(n806), .Z(n570) );
  MUX U3832 ( .IN0(n845), .IN1(n571), .SEL(n846), .F(n825) );
  IV U3833 ( .A(n847), .Z(n571) );
  XNOR U3834 ( .A(n819), .B(n817), .Z(n800) );
  MUX U3835 ( .IN0(n5152), .IN1(n5150), .SEL(n5151), .F(n572) );
  IV U3836 ( .A(n572), .Z(n4064) );
  MUX U3837 ( .IN0(n5107), .IN1(n5105), .SEL(n5106), .F(n573) );
  IV U3838 ( .A(n573), .Z(n4043) );
  MUX U3839 ( .IN0(n5065), .IN1(n5063), .SEL(n5064), .F(n574) );
  IV U3840 ( .A(n574), .Z(n4015) );
  MUX U3841 ( .IN0(n5045), .IN1(n5043), .SEL(n5044), .F(n575) );
  IV U3842 ( .A(n575), .Z(n4004) );
  MUX U3843 ( .IN0(n5079), .IN1(n5077), .SEL(n5078), .F(n576) );
  IV U3844 ( .A(n576), .Z(n4025) );
  MUX U3845 ( .IN0(n5210), .IN1(n5208), .SEL(n5209), .F(n577) );
  IV U3846 ( .A(n577), .Z(n4095) );
  MUX U3847 ( .IN0(n5167), .IN1(n5165), .SEL(n5166), .F(n578) );
  IV U3848 ( .A(n578), .Z(n4073) );
  MUX U3849 ( .IN0(n5238), .IN1(n5236), .SEL(n5237), .F(n579) );
  IV U3850 ( .A(n579), .Z(n4111) );
  MUX U3851 ( .IN0(n5218), .IN1(n5216), .SEL(n5217), .F(n580) );
  IV U3852 ( .A(n580), .Z(n4100) );
  MUX U3853 ( .IN0(n5252), .IN1(n5250), .SEL(n5251), .F(n581) );
  IV U3854 ( .A(n581), .Z(n4119) );
  MUX U3855 ( .IN0(n2668), .IN1(n2666), .SEL(n2667), .F(n582) );
  IV U3856 ( .A(n582), .Z(n1794) );
  MUX U3857 ( .IN0(n2627), .IN1(n2625), .SEL(n2626), .F(n583) );
  IV U3858 ( .A(n583), .Z(n1771) );
  MUX U3859 ( .IN0(n2585), .IN1(n2583), .SEL(n2584), .F(n584) );
  IV U3860 ( .A(n584), .Z(n1747) );
  MUX U3861 ( .IN0(n2565), .IN1(n2563), .SEL(n2564), .F(n585) );
  IV U3862 ( .A(n585), .Z(n1734) );
  MUX U3863 ( .IN0(n2599), .IN1(n2597), .SEL(n2598), .F(n586) );
  IV U3864 ( .A(n586), .Z(n1755) );
  MUX U3865 ( .IN0(n2726), .IN1(n2724), .SEL(n2725), .F(n587) );
  IV U3866 ( .A(n587), .Z(n1825) );
  MUX U3867 ( .IN0(n2683), .IN1(n2681), .SEL(n2682), .F(n588) );
  IV U3868 ( .A(n588), .Z(n1803) );
  MUX U3869 ( .IN0(n2754), .IN1(n2752), .SEL(n2753), .F(n589) );
  IV U3870 ( .A(n589), .Z(n1841) );
  MUX U3871 ( .IN0(n2734), .IN1(n2732), .SEL(n2733), .F(n590) );
  IV U3872 ( .A(n590), .Z(n1830) );
  MUX U3873 ( .IN0(n2768), .IN1(n2766), .SEL(n2767), .F(n591) );
  IV U3874 ( .A(n591), .Z(n1852) );
  MUX U3875 ( .IN0(n6880), .IN1(n6878), .SEL(n6879), .F(n592) );
  IV U3876 ( .A(n592), .Z(n5036) );
  MUX U3877 ( .IN0(n6835), .IN1(n6833), .SEL(n6834), .F(n593) );
  IV U3878 ( .A(n593), .Z(n5016) );
  MUX U3879 ( .IN0(n6793), .IN1(n6791), .SEL(n6792), .F(n594) );
  IV U3880 ( .A(n594), .Z(n4988) );
  MUX U3881 ( .IN0(n6773), .IN1(n6771), .SEL(n6772), .F(n595) );
  IV U3882 ( .A(n595), .Z(n4977) );
  MUX U3883 ( .IN0(n6709), .IN1(n6707), .SEL(n6708), .F(n596) );
  IV U3884 ( .A(n596), .Z(n4937) );
  MUX U3885 ( .IN0(n6666), .IN1(n6664), .SEL(n6665), .F(n597) );
  IV U3886 ( .A(n597), .Z(n4915) );
  MUX U3887 ( .IN0(n6737), .IN1(n6735), .SEL(n6736), .F(n598) );
  IV U3888 ( .A(n598), .Z(n4954) );
  MUX U3889 ( .IN0(n6751), .IN1(n6749), .SEL(n6750), .F(n599) );
  IV U3890 ( .A(n599), .Z(n4964) );
  MUX U3891 ( .IN0(n6535), .IN1(n6533), .SEL(n6534), .F(n600) );
  IV U3892 ( .A(n600), .Z(n4840) );
  MUX U3893 ( .IN0(n6490), .IN1(n6488), .SEL(n6489), .F(n601) );
  IV U3894 ( .A(n601), .Z(n4819) );
  MUX U3895 ( .IN0(n6446), .IN1(n6444), .SEL(n6445), .F(n602) );
  IV U3896 ( .A(n602), .Z(n4792) );
  MUX U3897 ( .IN0(n6460), .IN1(n6458), .SEL(n6459), .F(n603) );
  IV U3898 ( .A(n603), .Z(n4802) );
  MUX U3899 ( .IN0(n6593), .IN1(n6591), .SEL(n6592), .F(n604) );
  IV U3900 ( .A(n604), .Z(n4873) );
  MUX U3901 ( .IN0(n6573), .IN1(n6571), .SEL(n6572), .F(n605) );
  IV U3902 ( .A(n605), .Z(n4862) );
  MUX U3903 ( .IN0(n6621), .IN1(n6619), .SEL(n6620), .F(n606) );
  IV U3904 ( .A(n606), .Z(n4891) );
  MUX U3905 ( .IN0(n6601), .IN1(n6599), .SEL(n6600), .F(n607) );
  IV U3906 ( .A(n607), .Z(n4878) );
  MUX U3907 ( .IN0(n6635), .IN1(n6633), .SEL(n6634), .F(n608) );
  IV U3908 ( .A(n608), .Z(n4899) );
  MUX U3909 ( .IN0(n6192), .IN1(n6190), .SEL(n6191), .F(n609) );
  IV U3910 ( .A(n609), .Z(n4648) );
  MUX U3911 ( .IN0(n6147), .IN1(n6145), .SEL(n6146), .F(n610) );
  IV U3912 ( .A(n610), .Z(n4627) );
  MUX U3913 ( .IN0(n6101), .IN1(n6099), .SEL(n6100), .F(n611) );
  IV U3914 ( .A(n611), .Z(n4600) );
  MUX U3915 ( .IN0(n6081), .IN1(n6079), .SEL(n6080), .F(n612) );
  IV U3916 ( .A(n612), .Z(n4589) );
  MUX U3917 ( .IN0(n6017), .IN1(n6015), .SEL(n6016), .F(n613) );
  IV U3918 ( .A(n613), .Z(n4550) );
  MUX U3919 ( .IN0(n5974), .IN1(n5972), .SEL(n5973), .F(n614) );
  IV U3920 ( .A(n614), .Z(n4528) );
  MUX U3921 ( .IN0(n6045), .IN1(n6043), .SEL(n6044), .F(n615) );
  IV U3922 ( .A(n615), .Z(n4566) );
  MUX U3923 ( .IN0(n6025), .IN1(n6023), .SEL(n6024), .F(n616) );
  IV U3924 ( .A(n616), .Z(n4555) );
  MUX U3925 ( .IN0(n6306), .IN1(n6304), .SEL(n6305), .F(n617) );
  IV U3926 ( .A(n617), .Z(n4713) );
  MUX U3927 ( .IN0(n6265), .IN1(n6263), .SEL(n6264), .F(n618) );
  IV U3928 ( .A(n618), .Z(n4690) );
  MUX U3929 ( .IN0(n6223), .IN1(n6221), .SEL(n6222), .F(n619) );
  IV U3930 ( .A(n619), .Z(n4664) );
  MUX U3931 ( .IN0(n6237), .IN1(n6235), .SEL(n6236), .F(n620) );
  IV U3932 ( .A(n620), .Z(n4672) );
  MUX U3933 ( .IN0(n6362), .IN1(n6360), .SEL(n6361), .F(n621) );
  IV U3934 ( .A(n621), .Z(n4745) );
  MUX U3935 ( .IN0(n6342), .IN1(n6340), .SEL(n6341), .F(n622) );
  IV U3936 ( .A(n622), .Z(n4734) );
  MUX U3937 ( .IN0(n6321), .IN1(n6319), .SEL(n6320), .F(n623) );
  IV U3938 ( .A(n623), .Z(n4722) );
  MUX U3939 ( .IN0(n6328), .IN1(n6326), .SEL(n6327), .F(n624) );
  IV U3940 ( .A(n624), .Z(n4726) );
  MUX U3941 ( .IN0(n6390), .IN1(n6388), .SEL(n6389), .F(n625) );
  IV U3942 ( .A(n625), .Z(n4761) );
  MUX U3943 ( .IN0(n6370), .IN1(n6368), .SEL(n6369), .F(n626) );
  IV U3944 ( .A(n626), .Z(n4750) );
  MUX U3945 ( .IN0(n6404), .IN1(n6402), .SEL(n6403), .F(n627) );
  IV U3946 ( .A(n627), .Z(n4771) );
  MUX U3947 ( .IN0(n6411), .IN1(n6409), .SEL(n6410), .F(n628) );
  IV U3948 ( .A(n628), .Z(n4775) );
  MUX U3949 ( .IN0(n5495), .IN1(n5493), .SEL(n5494), .F(n629) );
  IV U3950 ( .A(n629), .Z(n4257) );
  MUX U3951 ( .IN0(n5452), .IN1(n5450), .SEL(n5451), .F(n630) );
  IV U3952 ( .A(n630), .Z(n4235) );
  MUX U3953 ( .IN0(n5410), .IN1(n5408), .SEL(n5409), .F(n631) );
  IV U3954 ( .A(n631), .Z(n4207) );
  MUX U3955 ( .IN0(n5390), .IN1(n5388), .SEL(n5389), .F(n632) );
  IV U3956 ( .A(n632), .Z(n4196) );
  MUX U3957 ( .IN0(n5326), .IN1(n5324), .SEL(n5325), .F(n633) );
  IV U3958 ( .A(n633), .Z(n4159) );
  MUX U3959 ( .IN0(n5281), .IN1(n5279), .SEL(n5280), .F(n634) );
  IV U3960 ( .A(n634), .Z(n4138) );
  MUX U3961 ( .IN0(n5354), .IN1(n5352), .SEL(n5353), .F(n635) );
  IV U3962 ( .A(n635), .Z(n4175) );
  MUX U3963 ( .IN0(n5334), .IN1(n5332), .SEL(n5333), .F(n636) );
  IV U3964 ( .A(n636), .Z(n4164) );
  MUX U3965 ( .IN0(n5364), .IN1(n5362), .SEL(n5363), .F(n637) );
  IV U3966 ( .A(n637), .Z(n4178) );
  MUX U3967 ( .IN0(n5729), .IN1(n5727), .SEL(n5728), .F(n638) );
  IV U3968 ( .A(n638), .Z(n4389) );
  MUX U3969 ( .IN0(n5684), .IN1(n5682), .SEL(n5683), .F(n639) );
  IV U3970 ( .A(n639), .Z(n4368) );
  MUX U3971 ( .IN0(n5638), .IN1(n5636), .SEL(n5637), .F(n640) );
  IV U3972 ( .A(n640), .Z(n4341) );
  MUX U3973 ( .IN0(n5618), .IN1(n5616), .SEL(n5617), .F(n641) );
  IV U3974 ( .A(n641), .Z(n4330) );
  MUX U3975 ( .IN0(n5554), .IN1(n5552), .SEL(n5553), .F(n642) );
  IV U3976 ( .A(n642), .Z(n4289) );
  MUX U3977 ( .IN0(n5511), .IN1(n5509), .SEL(n5510), .F(n643) );
  IV U3978 ( .A(n643), .Z(n4267) );
  MUX U3979 ( .IN0(n5582), .IN1(n5580), .SEL(n5581), .F(n644) );
  IV U3980 ( .A(n644), .Z(n4305) );
  MUX U3981 ( .IN0(n5562), .IN1(n5560), .SEL(n5561), .F(n645) );
  IV U3982 ( .A(n645), .Z(n4294) );
  MUX U3983 ( .IN0(n5592), .IN1(n5590), .SEL(n5591), .F(n646) );
  IV U3984 ( .A(n646), .Z(n4308) );
  MUX U3985 ( .IN0(n5845), .IN1(n5843), .SEL(n5844), .F(n647) );
  IV U3986 ( .A(n647), .Z(n4453) );
  MUX U3987 ( .IN0(n5800), .IN1(n5798), .SEL(n5799), .F(n648) );
  IV U3988 ( .A(n648), .Z(n4432) );
  MUX U3989 ( .IN0(n5758), .IN1(n5756), .SEL(n5757), .F(n649) );
  IV U3990 ( .A(n649), .Z(n4406) );
  MUX U3991 ( .IN0(n5738), .IN1(n5736), .SEL(n5737), .F(n650) );
  IV U3992 ( .A(n650), .Z(n4395) );
  MUX U3993 ( .IN0(n5905), .IN1(n5903), .SEL(n5904), .F(n651) );
  IV U3994 ( .A(n651), .Z(n4485) );
  MUX U3995 ( .IN0(n5860), .IN1(n5858), .SEL(n5859), .F(n652) );
  IV U3996 ( .A(n652), .Z(n4464) );
  MUX U3997 ( .IN0(n5933), .IN1(n5931), .SEL(n5932), .F(n653) );
  IV U3998 ( .A(n653), .Z(n4501) );
  MUX U3999 ( .IN0(n5913), .IN1(n5911), .SEL(n5912), .F(n654) );
  IV U4000 ( .A(n654), .Z(n4490) );
  MUX U4001 ( .IN0(n2741), .IN1(n2743), .SEL(n2742), .F(n655) );
  IV U4002 ( .A(n655), .Z(n1832) );
  MUX U4003 ( .IN0(n2572), .IN1(n2574), .SEL(n2573), .F(n656) );
  IV U4004 ( .A(n656), .Z(n1736) );
  XOR U4005 ( .A(n4695), .B(n4693), .Z(n4687) );
  XOR U4006 ( .A(n4677), .B(n4675), .Z(n4669) );
  MUX U4007 ( .IN0(n6032), .IN1(n6034), .SEL(n6033), .F(n657) );
  IV U4008 ( .A(n657), .Z(n4557) );
  XOR U4009 ( .A(n4631), .B(n4630), .Z(n4624) );
  XOR U4010 ( .A(n4943), .B(n4941), .Z(n4951) );
  XOR U4011 ( .A(n5020), .B(n5019), .Z(n5013) );
  XOR U4012 ( .A(n4903), .B(n4902), .Z(n4896) );
  MUX U4013 ( .IN0(n6608), .IN1(n6610), .SEL(n6609), .F(n658) );
  IV U4014 ( .A(n658), .Z(n4880) );
  XOR U4015 ( .A(n4823), .B(n4822), .Z(n4816) );
  XOR U4016 ( .A(n4806), .B(n4805), .Z(n4799) );
  XOR U4017 ( .A(n4468), .B(n4467), .Z(n4461) );
  XOR U4018 ( .A(n4436), .B(n4435), .Z(n4429) );
  XOR U4019 ( .A(n4372), .B(n4371), .Z(n4365) );
  XOR U4020 ( .A(n4240), .B(n4238), .Z(n4232) );
  XOR U4021 ( .A(n4124), .B(n4122), .Z(n4116) );
  XOR U4022 ( .A(n4078), .B(n4076), .Z(n4070) );
  XOR U4023 ( .A(n4047), .B(n4046), .Z(n4040) );
  XOR U4024 ( .A(n4030), .B(n4028), .Z(n4022) );
  MUX U4025 ( .IN0(n4059), .IN1(n659), .SEL(n4060), .F(n3516) );
  IV U4026 ( .A(n4061), .Z(n659) );
  MUX U4027 ( .IN0(n4010), .IN1(n660), .SEL(n4011), .F(n3495) );
  IV U4028 ( .A(n4012), .Z(n660) );
  MUX U4029 ( .IN0(n4090), .IN1(n661), .SEL(n4091), .F(n3532) );
  IV U4030 ( .A(n4092), .Z(n661) );
  MUX U4031 ( .IN0(n4106), .IN1(n662), .SEL(n4107), .F(n3542) );
  IV U4032 ( .A(n4108), .Z(n662) );
  MUX U4033 ( .IN0(n3013), .IN1(n3011), .SEL(n3012), .F(n663) );
  IV U4034 ( .A(n663), .Z(n1990) );
  MUX U4035 ( .IN0(n2968), .IN1(n2966), .SEL(n2967), .F(n664) );
  IV U4036 ( .A(n664), .Z(n1970) );
  MUX U4037 ( .IN0(n2926), .IN1(n2924), .SEL(n2925), .F(n665) );
  IV U4038 ( .A(n665), .Z(n1944) );
  MUX U4039 ( .IN0(n2940), .IN1(n2938), .SEL(n2939), .F(n666) );
  IV U4040 ( .A(n666), .Z(n1954) );
  MUX U4041 ( .IN0(n2838), .IN1(n2836), .SEL(n2837), .F(n667) );
  IV U4042 ( .A(n667), .Z(n1894) );
  MUX U4043 ( .IN0(n2818), .IN1(n2816), .SEL(n2817), .F(n668) );
  IV U4044 ( .A(n668), .Z(n1883) );
  MUX U4045 ( .IN0(n2866), .IN1(n2864), .SEL(n2865), .F(n669) );
  IV U4046 ( .A(n669), .Z(n1910) );
  MUX U4047 ( .IN0(n2846), .IN1(n2844), .SEL(n2845), .F(n670) );
  IV U4048 ( .A(n670), .Z(n1899) );
  MUX U4049 ( .IN0(n2326), .IN1(n2324), .SEL(n2325), .F(n671) );
  MUX U4050 ( .IN0(n2289), .IN1(n2287), .SEL(n2288), .F(n672) );
  IV U4051 ( .A(n672), .Z(n1577) );
  MUX U4052 ( .IN0(n2296), .IN1(n2294), .SEL(n2295), .F(n673) );
  IV U4053 ( .A(n673), .Z(n1581) );
  MUX U4054 ( .IN0(n2234), .IN1(n2236), .SEL(n2235), .F(n674) );
  IV U4055 ( .A(n674), .Z(n1544) );
  MUX U4056 ( .IN0(n2247), .IN1(n2245), .SEL(n2246), .F(n675) );
  IV U4057 ( .A(n675), .Z(n1553) );
  MUX U4058 ( .IN0(n2227), .IN1(n2225), .SEL(n2226), .F(n676) );
  IV U4059 ( .A(n676), .Z(n1542) );
  MUX U4060 ( .IN0(n2261), .IN1(n2259), .SEL(n2260), .F(n677) );
  IV U4061 ( .A(n677), .Z(n1561) );
  MUX U4062 ( .IN0(n2268), .IN1(n2266), .SEL(n2267), .F(n678) );
  IV U4063 ( .A(n678), .Z(n1565) );
  MUX U4064 ( .IN0(n2163), .IN1(n2161), .SEL(n2162), .F(n679) );
  IV U4065 ( .A(n679), .Z(n1504) );
  MUX U4066 ( .IN0(n2122), .IN1(n2120), .SEL(n2121), .F(n680) );
  IV U4067 ( .A(n680), .Z(n1481) );
  MUX U4068 ( .IN0(n2187), .IN1(n2185), .SEL(n2186), .F(n681) );
  MUX U4069 ( .IN0(n2205), .IN1(n2203), .SEL(n2204), .F(n682) );
  IV U4070 ( .A(n682), .Z(n1529) );
  MUX U4071 ( .IN0(n2439), .IN1(n2437), .SEL(n2438), .F(n683) );
  MUX U4072 ( .IN0(n2402), .IN1(n2400), .SEL(n2401), .F(n684) );
  IV U4073 ( .A(n684), .Z(n1642) );
  MUX U4074 ( .IN0(n2409), .IN1(n2407), .SEL(n2408), .F(n685) );
  IV U4075 ( .A(n685), .Z(n1646) );
  MUX U4076 ( .IN0(n2359), .IN1(n2357), .SEL(n2358), .F(n686) );
  IV U4077 ( .A(n686), .Z(n1616) );
  XOR U4078 ( .A(n1606), .B(n1604), .Z(n1613) );
  MUX U4079 ( .IN0(n2373), .IN1(n2371), .SEL(n2372), .F(n687) );
  IV U4080 ( .A(n687), .Z(n1626) );
  MUX U4081 ( .IN0(n688), .IN1(n2385), .SEL(n2386), .F(n1631) );
  IV U4082 ( .A(n2387), .Z(n688) );
  MUX U4083 ( .IN0(n2497), .IN1(n2495), .SEL(n2496), .F(n689) );
  MUX U4084 ( .IN0(n2529), .IN1(n2527), .SEL(n2528), .F(n690) );
  IV U4085 ( .A(n690), .Z(n1712) );
  MUX U4086 ( .IN0(n2509), .IN1(n2507), .SEL(n2508), .F(n691) );
  IV U4087 ( .A(n691), .Z(n1701) );
  MUX U4088 ( .IN0(n2543), .IN1(n2541), .SEL(n2542), .F(n692) );
  IV U4089 ( .A(n692), .Z(n1721) );
  MUX U4090 ( .IN0(n2550), .IN1(n2548), .SEL(n2549), .F(n693) );
  IV U4091 ( .A(n693), .Z(n1725) );
  MUX U4092 ( .IN0(n1789), .IN1(n694), .SEL(n1790), .F(n1307) );
  IV U4093 ( .A(n1791), .Z(n694) );
  MUX U4094 ( .IN0(n1766), .IN1(n695), .SEL(n1767), .F(n1296) );
  IV U4095 ( .A(n1768), .Z(n695) );
  MUX U4096 ( .IN0(n1742), .IN1(n696), .SEL(n1743), .F(n1284) );
  IV U4097 ( .A(n1744), .Z(n696) );
  MUX U4098 ( .IN0(n1757), .IN1(n1760), .SEL(n1758), .F(n1289) );
  MUX U4099 ( .IN0(n1820), .IN1(n697), .SEL(n1821), .F(n1323) );
  IV U4100 ( .A(n1822), .Z(n697) );
  MUX U4101 ( .IN0(n1798), .IN1(n698), .SEL(n1799), .F(n1312) );
  IV U4102 ( .A(n1800), .Z(n698) );
  MUX U4103 ( .IN0(n1836), .IN1(n699), .SEL(n1837), .F(n1331) );
  IV U4104 ( .A(n1838), .Z(n699) );
  MUX U4105 ( .IN0(n1854), .IN1(n1857), .SEL(n1855), .F(n1335) );
  MUX U4106 ( .IN0(n5031), .IN1(n700), .SEL(n5032), .F(n3996) );
  IV U4107 ( .A(n5033), .Z(n700) );
  MUX U4108 ( .IN0(n4983), .IN1(n701), .SEL(n4984), .F(n3975) );
  IV U4109 ( .A(n4985), .Z(n701) );
  MUX U4110 ( .IN0(n4932), .IN1(n702), .SEL(n4933), .F(n3948) );
  IV U4111 ( .A(n4934), .Z(n702) );
  MUX U4112 ( .IN0(n4910), .IN1(n703), .SEL(n4911), .F(n3937) );
  IV U4113 ( .A(n4912), .Z(n703) );
  MUX U4114 ( .IN0(n4835), .IN1(n704), .SEL(n4836), .F(n3899) );
  IV U4115 ( .A(n4837), .Z(n704) );
  MUX U4116 ( .IN0(n4787), .IN1(n705), .SEL(n4788), .F(n3878) );
  IV U4117 ( .A(n4789), .Z(n705) );
  MUX U4118 ( .IN0(n4868), .IN1(n706), .SEL(n4869), .F(n3914) );
  IV U4119 ( .A(n4870), .Z(n706) );
  MUX U4120 ( .IN0(n4886), .IN1(n707), .SEL(n4887), .F(n3924) );
  IV U4121 ( .A(n4888), .Z(n707) );
  MUX U4122 ( .IN0(n4643), .IN1(n708), .SEL(n4644), .F(n3807) );
  IV U4123 ( .A(n4645), .Z(n708) );
  MUX U4124 ( .IN0(n4595), .IN1(n709), .SEL(n4596), .F(n3786) );
  IV U4125 ( .A(n4597), .Z(n709) );
  MUX U4126 ( .IN0(n4545), .IN1(n710), .SEL(n4546), .F(n3760) );
  IV U4127 ( .A(n4547), .Z(n710) );
  MUX U4128 ( .IN0(n4523), .IN1(n711), .SEL(n4524), .F(n3747) );
  IV U4129 ( .A(n4525), .Z(n711) );
  MUX U4130 ( .IN0(n4561), .IN1(n712), .SEL(n4562), .F(n3768) );
  IV U4131 ( .A(n4563), .Z(n712) );
  MUX U4132 ( .IN0(n4708), .IN1(n713), .SEL(n4709), .F(n3838) );
  IV U4133 ( .A(n4710), .Z(n713) );
  MUX U4134 ( .IN0(n4659), .IN1(n714), .SEL(n4660), .F(n3816) );
  IV U4135 ( .A(n4661), .Z(n714) );
  MUX U4136 ( .IN0(n4740), .IN1(n715), .SEL(n4741), .F(n3854) );
  IV U4137 ( .A(n4742), .Z(n715) );
  MUX U4138 ( .IN0(n4756), .IN1(n716), .SEL(n4757), .F(n3864) );
  IV U4139 ( .A(n4758), .Z(n716) );
  MUX U4140 ( .IN0(n4252), .IN1(n717), .SEL(n4253), .F(n3612) );
  IV U4141 ( .A(n4254), .Z(n717) );
  MUX U4142 ( .IN0(n4202), .IN1(n718), .SEL(n4203), .F(n3591) );
  IV U4143 ( .A(n4204), .Z(n718) );
  MUX U4144 ( .IN0(n4154), .IN1(n719), .SEL(n4155), .F(n3565) );
  IV U4145 ( .A(n4156), .Z(n719) );
  MUX U4146 ( .IN0(n4170), .IN1(n720), .SEL(n4171), .F(n3573) );
  IV U4147 ( .A(n4172), .Z(n720) );
  MUX U4148 ( .IN0(n4384), .IN1(n721), .SEL(n4385), .F(n3678) );
  IV U4149 ( .A(n4386), .Z(n721) );
  MUX U4150 ( .IN0(n4336), .IN1(n722), .SEL(n4337), .F(n3657) );
  IV U4151 ( .A(n4338), .Z(n722) );
  MUX U4152 ( .IN0(n4284), .IN1(n723), .SEL(n4285), .F(n3629) );
  IV U4153 ( .A(n4286), .Z(n723) );
  MUX U4154 ( .IN0(n4300), .IN1(n724), .SEL(n4301), .F(n3639) );
  IV U4155 ( .A(n4302), .Z(n724) );
  MUX U4156 ( .IN0(n4448), .IN1(n725), .SEL(n4449), .F(n3711) );
  IV U4157 ( .A(n4450), .Z(n725) );
  MUX U4158 ( .IN0(n4401), .IN1(n726), .SEL(n4402), .F(n3689) );
  IV U4159 ( .A(n4403), .Z(n726) );
  MUX U4160 ( .IN0(n4480), .IN1(n727), .SEL(n4481), .F(n3726) );
  IV U4161 ( .A(n4482), .Z(n727) );
  MUX U4162 ( .IN0(n4496), .IN1(n728), .SEL(n4497), .F(n3736) );
  IV U4163 ( .A(n4498), .Z(n728) );
  MUX U4164 ( .IN0(n2474), .IN1(n2476), .SEL(n2475), .F(n729) );
  IV U4165 ( .A(n729), .Z(n1680) );
  XOR U4166 ( .A(n4768), .B(n4767), .Z(n4754) );
  XOR U4167 ( .A(n4719), .B(n4718), .Z(n4738) );
  XOR U4168 ( .A(n4607), .B(n4606), .Z(n4593) );
  XOR U4169 ( .A(n4995), .B(n4994), .Z(n4981) );
  XOR U4170 ( .A(n4848), .B(n4847), .Z(n4866) );
  XOR U4171 ( .A(n4348), .B(n4347), .Z(n4334) );
  XOR U4172 ( .A(n4214), .B(n4213), .Z(n4200) );
  XOR U4173 ( .A(n3741), .B(n3739), .Z(n3733) );
  XOR U4174 ( .A(n3694), .B(n3692), .Z(n3686) );
  XOR U4175 ( .A(n3661), .B(n3660), .Z(n3654) );
  XOR U4176 ( .A(n3644), .B(n3642), .Z(n3636) );
  XOR U4177 ( .A(n3595), .B(n3594), .Z(n3588) );
  XOR U4178 ( .A(n3578), .B(n3576), .Z(n3570) );
  XOR U4179 ( .A(n3904), .B(n3903), .Z(n3911) );
  XOR U4180 ( .A(n3979), .B(n3978), .Z(n3972) );
  XOR U4181 ( .A(n3790), .B(n3789), .Z(n3783) );
  XOR U4182 ( .A(n3773), .B(n3771), .Z(n3765) );
  MUX U4183 ( .IN0(n4534), .IN1(n730), .SEL(n4535), .F(n3749) );
  IV U4184 ( .A(n4536), .Z(n730) );
  MUX U4185 ( .IN0(n3511), .IN1(n731), .SEL(n3512), .F(n3254) );
  IV U4186 ( .A(n3513), .Z(n731) );
  MUX U4187 ( .IN0(n3527), .IN1(n732), .SEL(n3528), .F(n3262) );
  IV U4188 ( .A(n3529), .Z(n732) );
  MUX U4189 ( .IN0(n1985), .IN1(n733), .SEL(n1986), .F(n1400) );
  IV U4190 ( .A(n1987), .Z(n733) );
  MUX U4191 ( .IN0(n1965), .IN1(n734), .SEL(n1966), .F(n1389) );
  IV U4192 ( .A(n1967), .Z(n734) );
  MUX U4193 ( .IN0(n1889), .IN1(n735), .SEL(n1890), .F(n1353) );
  IV U4194 ( .A(n1891), .Z(n735) );
  MUX U4195 ( .IN0(n1905), .IN1(n736), .SEL(n1906), .F(n1363) );
  IV U4196 ( .A(n1907), .Z(n736) );
  MUX U4197 ( .IN0(n1591), .IN1(n737), .SEL(n1592), .F(n1207) );
  IV U4198 ( .A(n1593), .Z(n737) );
  MUX U4199 ( .IN0(n1548), .IN1(n738), .SEL(n1549), .F(n1189) );
  IV U4200 ( .A(n1550), .Z(n738) );
  MUX U4201 ( .IN0(n1556), .IN1(n739), .SEL(n1557), .F(n1193) );
  IV U4202 ( .A(n1558), .Z(n739) );
  MUX U4203 ( .IN0(n1499), .IN1(n740), .SEL(n1500), .F(n1165) );
  IV U4204 ( .A(n1501), .Z(n740) );
  MUX U4205 ( .IN0(n1476), .IN1(n741), .SEL(n1477), .F(n1154) );
  IV U4206 ( .A(n1478), .Z(n741) );
  MUX U4207 ( .IN0(n1656), .IN1(n742), .SEL(n1657), .F(n1240) );
  IV U4208 ( .A(n1658), .Z(n742) );
  MUX U4209 ( .IN0(n1688), .IN1(n743), .SEL(n1689), .F(n1255) );
  IV U4210 ( .A(n1690), .Z(n743) );
  MUX U4211 ( .IN0(n1707), .IN1(n744), .SEL(n1708), .F(n1268) );
  IV U4212 ( .A(n1709), .Z(n744) );
  MUX U4213 ( .IN0(n1716), .IN1(n745), .SEL(n1717), .F(n1272) );
  IV U4214 ( .A(n1718), .Z(n745) );
  MUX U4215 ( .IN0(n1302), .IN1(n746), .SEL(n1303), .F(n1065) );
  IV U4216 ( .A(n1304), .Z(n746) );
  MUX U4217 ( .IN0(n1318), .IN1(n747), .SEL(n1319), .F(n1073) );
  IV U4218 ( .A(n1320), .Z(n747) );
  MUX U4219 ( .IN0(n3991), .IN1(n748), .SEL(n3992), .F(n3482) );
  IV U4220 ( .A(n3993), .Z(n748) );
  MUX U4221 ( .IN0(n3943), .IN1(n749), .SEL(n3944), .F(n3461) );
  IV U4222 ( .A(n3945), .Z(n749) );
  MUX U4223 ( .IN0(n3894), .IN1(n750), .SEL(n3895), .F(n3436) );
  IV U4224 ( .A(n3896), .Z(n750) );
  MUX U4225 ( .IN0(n3873), .IN1(n751), .SEL(n3874), .F(n3425) );
  IV U4226 ( .A(n3875), .Z(n751) );
  MUX U4227 ( .IN0(n3802), .IN1(n752), .SEL(n3803), .F(n3392) );
  IV U4228 ( .A(n3804), .Z(n752) );
  MUX U4229 ( .IN0(n3755), .IN1(n753), .SEL(n3756), .F(n3370) );
  IV U4230 ( .A(n3757), .Z(n753) );
  MUX U4231 ( .IN0(n3833), .IN1(n754), .SEL(n3834), .F(n3408) );
  IV U4232 ( .A(n3835), .Z(n754) );
  MUX U4233 ( .IN0(n3811), .IN1(n755), .SEL(n3812), .F(n3397) );
  IV U4234 ( .A(n3813), .Z(n755) );
  MUX U4235 ( .IN0(n3845), .IN1(n756), .SEL(n3846), .F(n3411) );
  IV U4236 ( .A(n3847), .Z(n756) );
  MUX U4237 ( .IN0(n3607), .IN1(n757), .SEL(n3608), .F(n3300) );
  IV U4238 ( .A(n3609), .Z(n757) );
  MUX U4239 ( .IN0(n3560), .IN1(n758), .SEL(n3561), .F(n3278) );
  IV U4240 ( .A(n3562), .Z(n758) );
  MUX U4241 ( .IN0(n3673), .IN1(n759), .SEL(n3674), .F(n3331) );
  IV U4242 ( .A(n3675), .Z(n759) );
  MUX U4243 ( .IN0(n3624), .IN1(n760), .SEL(n3625), .F(n3309) );
  IV U4244 ( .A(n3626), .Z(n760) );
  MUX U4245 ( .IN0(n3706), .IN1(n761), .SEL(n3707), .F(n3346) );
  IV U4246 ( .A(n3708), .Z(n761) );
  MUX U4247 ( .IN0(n3721), .IN1(n762), .SEL(n3722), .F(n3356) );
  IV U4248 ( .A(n3723), .Z(n762) );
  XOR U4249 ( .A(n2915), .B(n2914), .Z(n2986) );
  XOR U4250 ( .A(n5922), .B(n5921), .Z(n5878) );
  XOR U4251 ( .A(n5747), .B(n5746), .Z(n5818) );
  XOR U4252 ( .A(n5627), .B(n5626), .Z(n5702) );
  XOR U4253 ( .A(n5227), .B(n5226), .Z(n5183) );
  XOR U4254 ( .A(n5054), .B(n5053), .Z(n5125) );
  XOR U4255 ( .A(n5399), .B(n5398), .Z(n5468) );
  XOR U4256 ( .A(n6782), .B(n6781), .Z(n6853) );
  XOR U4257 ( .A(n6212), .B(n6211), .Z(n6281) );
  XOR U4258 ( .A(n6090), .B(n6089), .Z(n6165) );
  XOR U4259 ( .A(n1513), .B(n1512), .Z(n1489) );
  XOR U4260 ( .A(n1937), .B(n1936), .Z(n1976) );
  XOR U4261 ( .A(n1375), .B(n1374), .Z(n1393) );
  XOR U4262 ( .A(n3955), .B(n3954), .Z(n3941) );
  MUX U4263 ( .IN0(n2062), .IN1(n2060), .SEL(n2061), .F(n763) );
  IV U4264 ( .A(n763), .Z(n1446) );
  MUX U4265 ( .IN0(n2069), .IN1(n2067), .SEL(n2068), .F(n764) );
  IV U4266 ( .A(n764), .Z(n1450) );
  XOR U4267 ( .A(n3465), .B(n3464), .Z(n3458) );
  MUX U4268 ( .IN0(n2021), .IN1(n2019), .SEL(n2020), .F(n765) );
  IV U4269 ( .A(n765), .Z(n1421) );
  MUX U4270 ( .IN0(n2035), .IN1(n2033), .SEL(n2034), .F(n766) );
  IV U4271 ( .A(n766), .Z(n1431) );
  MUX U4272 ( .IN0(n2042), .IN1(n2040), .SEL(n2041), .F(n767) );
  IV U4273 ( .A(n767), .Z(n1435) );
  MUX U4274 ( .IN0(n3249), .IN1(n768), .SEL(n3250), .F(n3124) );
  IV U4275 ( .A(n3251), .Z(n768) );
  MUX U4276 ( .IN0(n3257), .IN1(n769), .SEL(n3258), .F(n3128) );
  IV U4277 ( .A(n3259), .Z(n769) );
  MUX U4278 ( .IN0(n1395), .IN1(n770), .SEL(n1396), .F(n1113) );
  IV U4279 ( .A(n1397), .Z(n770) );
  XOR U4280 ( .A(n1103), .B(n1101), .Z(n1110) );
  MUX U4281 ( .IN0(n1341), .IN1(n1343), .SEL(n1342), .F(n1092) );
  MUX U4282 ( .IN0(n1365), .IN1(n1367), .SEL(n1366), .F(n1095) );
  MUX U4283 ( .IN0(n1203), .IN1(n771), .SEL(n1204), .F(n1010) );
  IV U4284 ( .A(n1205), .Z(n771) );
  MUX U4285 ( .IN0(n1160), .IN1(n772), .SEL(n1161), .F(n992) );
  IV U4286 ( .A(n1162), .Z(n772) );
  MUX U4287 ( .IN0(n1168), .IN1(n773), .SEL(n1169), .F(n996) );
  IV U4288 ( .A(n1170), .Z(n773) );
  MUX U4289 ( .IN0(n1236), .IN1(n774), .SEL(n1237), .F(n1027) );
  IV U4290 ( .A(n1238), .Z(n774) );
  MUX U4291 ( .IN0(n1248), .IN1(n1250), .SEL(n1249), .F(n1041) );
  MUX U4292 ( .IN0(n3477), .IN1(n775), .SEL(n3478), .F(n3237) );
  IV U4293 ( .A(n3479), .Z(n775) );
  MUX U4294 ( .IN0(n3431), .IN1(n776), .SEL(n3432), .F(n3215) );
  IV U4295 ( .A(n3433), .Z(n776) );
  MUX U4296 ( .IN0(n3387), .IN1(n777), .SEL(n3388), .F(n3192) );
  IV U4297 ( .A(n3389), .Z(n777) );
  MUX U4298 ( .IN0(n3403), .IN1(n778), .SEL(n3404), .F(n3200) );
  IV U4299 ( .A(n3405), .Z(n778) );
  MUX U4300 ( .IN0(n3295), .IN1(n779), .SEL(n3296), .F(n3147) );
  IV U4301 ( .A(n3297), .Z(n779) );
  MUX U4302 ( .IN0(n3273), .IN1(n780), .SEL(n3274), .F(n3136) );
  IV U4303 ( .A(n3275), .Z(n780) );
  MUX U4304 ( .IN0(n3326), .IN1(n781), .SEL(n3327), .F(n3163) );
  IV U4305 ( .A(n3328), .Z(n781) );
  MUX U4306 ( .IN0(n3304), .IN1(n782), .SEL(n3305), .F(n3152) );
  IV U4307 ( .A(n3306), .Z(n782) );
  MUX U4308 ( .IN0(n3341), .IN1(n783), .SEL(n3342), .F(n3171) );
  IV U4309 ( .A(n3343), .Z(n783) );
  MUX U4310 ( .IN0(n3349), .IN1(n784), .SEL(n3350), .F(n3175) );
  IV U4311 ( .A(n3351), .Z(n784) );
  XOR U4312 ( .A(n2813), .B(n2812), .Z(n2956) );
  XOR U4313 ( .A(n5527), .B(n5526), .Z(n5672) );
  XOR U4314 ( .A(n5299), .B(n5298), .Z(n5440) );
  XOR U4315 ( .A(n6682), .B(n6681), .Z(n6823) );
  XOR U4316 ( .A(n1879), .B(n1878), .Z(n1962) );
  XOR U4317 ( .A(n4923), .B(n4922), .Z(n5006) );
  XOR U4318 ( .A(n4275), .B(n4274), .Z(n4358) );
  XOR U4319 ( .A(n4145), .B(n4144), .Z(n4225) );
  XOR U4320 ( .A(n1346), .B(n1345), .Z(n1385) );
  XOR U4321 ( .A(n1253), .B(n1252), .Z(n1230) );
  MUX U4322 ( .IN0(n1408), .IN1(n1411), .SEL(n1409), .F(n1128) );
  XOR U4323 ( .A(n3443), .B(n3442), .Z(n3429) );
  XOR U4324 ( .A(n3219), .B(n3218), .Z(n3212) );
  XOR U4325 ( .A(n3205), .B(n3203), .Z(n3197) );
  MUX U4326 ( .IN0(n3119), .IN1(n785), .SEL(n3120), .F(n3063) );
  IV U4327 ( .A(n3121), .Z(n785) );
  MUX U4328 ( .IN0(n1006), .IN1(n786), .SEL(n1007), .F(n911) );
  IV U4329 ( .A(n1008), .Z(n786) );
  MUX U4330 ( .IN0(n1018), .IN1(n1020), .SEL(n1019), .F(n925) );
  MUX U4331 ( .IN0(n3232), .IN1(n787), .SEL(n3233), .F(n3114) );
  IV U4332 ( .A(n3234), .Z(n787) );
  MUX U4333 ( .IN0(n3187), .IN1(n788), .SEL(n3188), .F(n3095) );
  IV U4334 ( .A(n3189), .Z(n788) );
  MUX U4335 ( .IN0(n3142), .IN1(n789), .SEL(n3143), .F(n3074) );
  IV U4336 ( .A(n3144), .Z(n789) );
  MUX U4337 ( .IN0(n3158), .IN1(n790), .SEL(n3159), .F(n3082) );
  IV U4338 ( .A(n3160), .Z(n790) );
  MUX U4339 ( .IN0(n3166), .IN1(n791), .SEL(n3167), .F(n3086) );
  IV U4340 ( .A(n3168), .Z(n791) );
  XOR U4341 ( .A(n2615), .B(n2614), .Z(n2900) );
  XOR U4342 ( .A(n6478), .B(n6477), .Z(n6767) );
  XOR U4343 ( .A(n1443), .B(n1442), .Z(n1461) );
  XOR U4344 ( .A(n1428), .B(n1427), .Z(n1414) );
  XOR U4345 ( .A(n1634), .B(n1633), .Z(n1537) );
  XOR U4346 ( .A(n1763), .B(n1762), .Z(n1928) );
  XOR U4347 ( .A(n4809), .B(n4808), .Z(n4972) );
  XOR U4348 ( .A(n4422), .B(n4421), .Z(n4325) );
  XOR U4349 ( .A(n4033), .B(n4032), .Z(n4191) );
  XOR U4350 ( .A(n1292), .B(n1291), .Z(n1370) );
  XOR U4351 ( .A(n3502), .B(n3501), .Z(n3581) );
  XOR U4352 ( .A(n3885), .B(n3884), .Z(n3965) );
  XOR U4353 ( .A(n1025), .B(n1024), .Z(n1000) );
  XOR U4354 ( .A(n1058), .B(n1057), .Z(n1098) );
  XOR U4355 ( .A(n936), .B(n935), .Z(n954) );
  MUX U4356 ( .IN0(n1146), .IN1(n1148), .SEL(n1147), .F(n1142) );
  MUX U4357 ( .IN0(n3109), .IN1(n792), .SEL(n3110), .F(n3057) );
  IV U4358 ( .A(n3111), .Z(n792) );
  MUX U4359 ( .IN0(n3090), .IN1(n793), .SEL(n3091), .F(n3049) );
  IV U4360 ( .A(n3092), .Z(n793) );
  MUX U4361 ( .IN0(n3065), .IN1(n794), .SEL(n3066), .F(n3035) );
  IV U4362 ( .A(n3067), .Z(n794) );
  XOR U4363 ( .A(n2221), .B(n2220), .Z(n2784) );
  XOR U4364 ( .A(n2010), .B(n2009), .Z(n2078) );
  XOR U4365 ( .A(n6075), .B(n6074), .Z(n6653) );
  XOR U4366 ( .A(n4584), .B(n4583), .Z(n4906) );
  XOR U4367 ( .A(n3647), .B(n3646), .Z(n3550) );
  XOR U4368 ( .A(n3776), .B(n3775), .Z(n3932) );
  XOR U4369 ( .A(n972), .B(n971), .Z(n979) );
  MUX U4370 ( .IN0(n1274), .IN1(n1132), .SEL(n1275), .F(n1046) );
  XOR U4371 ( .A(n3378), .B(n3377), .Z(n3453) );
  XOR U4372 ( .A(n909), .B(n908), .Z(n947) );
  MUX U4373 ( .IN0(n886), .IN1(n888), .SEL(n887), .F(n882) );
  XOR U4374 ( .A(n839), .B(n837), .Z(n847) );
  MUX U4375 ( .IN0(n3052), .IN1(n795), .SEL(n3053), .F(n3030) );
  IV U4376 ( .A(n3054), .Z(n795) );
  XOR U4377 ( .A(n5268), .B(n5267), .Z(n6886) );
  MUX U4378 ( .IN0(n796), .IN1(n1992), .SEL(n815), .F(n1402) );
  IV U4379 ( .A(n816), .Z(n796) );
  XOR U4380 ( .A(n3270), .B(n3269), .Z(n1117) );
  XOR U4381 ( .A(n3132), .B(n3131), .Z(n967) );
  MUX U4382 ( .IN0(n797), .IN1(n889), .SEL(n807), .F(n852) );
  IV U4383 ( .A(n808), .Z(n797) );
  XOR U4384 ( .A(n3026), .B(n3025), .Z(n833) );
  MUX U4385 ( .IN0(n817), .IN1(n798), .SEL(n800), .F(o[10]) );
  IV U4386 ( .A(n799), .Z(n798) );
  XNOR U4387 ( .A(n799), .B(n800), .Z(o[9]) );
  XOR U4388 ( .A(n801), .B(n802), .Z(o[8]) );
  XNOR U4389 ( .A(n803), .B(n804), .Z(o[7]) );
  XOR U4390 ( .A(n805), .B(n806), .Z(o[6]) );
  XOR U4391 ( .A(n807), .B(n808), .Z(o[5]) );
  XOR U4392 ( .A(n809), .B(n810), .Z(o[4]) );
  XOR U4393 ( .A(n811), .B(n812), .Z(o[3]) );
  XOR U4394 ( .A(n813), .B(n814), .Z(o[2]) );
  XOR U4395 ( .A(n815), .B(n816), .Z(o[1]) );
  NAND U4396 ( .A(n818), .B(n802), .Z(n799) );
  XOR U4397 ( .A(n821), .B(n822), .Z(n801) );
  XNOR U4398 ( .A(n823), .B(n820), .Z(n821) );
  XOR U4399 ( .A(n824), .B(n825), .Z(n802) );
  XNOR U4400 ( .A(n818), .B(n826), .Z(n824) );
  AND U4401 ( .A(n827), .B(n828), .Z(n826) );
  XNOR U4402 ( .A(n825), .B(n829), .Z(n828) );
  ANDN U4403 ( .B(n830), .A(n804), .Z(n818) );
  XNOR U4404 ( .A(n832), .B(n833), .Z(n803) );
  XNOR U4405 ( .A(n834), .B(n831), .Z(n832) );
  XOR U4406 ( .A(n835), .B(n829), .Z(n804) );
  XNOR U4407 ( .A(n827), .B(n830), .Z(n835) );
  XOR U4408 ( .A(n843), .B(n844), .Z(n827) );
  IV U4409 ( .A(n825), .Z(n844) );
  XNOR U4410 ( .A(n853), .B(n854), .Z(n805) );
  XNOR U4411 ( .A(n855), .B(n852), .Z(n853) );
  XOR U4412 ( .A(n841), .B(n842), .Z(n806) );
  NANDN U4413 ( .A(n856), .B(n857), .Z(n842) );
  XOR U4414 ( .A(n858), .B(n847), .Z(n841) );
  XOR U4415 ( .A(n859), .B(n836), .Z(n837) );
  IV U4416 ( .A(n838), .Z(n836) );
  XNOR U4417 ( .A(n846), .B(n840), .Z(n858) );
  IV U4418 ( .A(n857), .Z(n873) );
  XOR U4419 ( .A(n874), .B(n851), .Z(n846) );
  XNOR U4420 ( .A(n849), .B(n845), .Z(n874) );
  XOR U4421 ( .A(n882), .B(n848), .Z(n849) );
  IV U4422 ( .A(n850), .Z(n848) );
  XNOR U4423 ( .A(n890), .B(n891), .Z(n807) );
  XNOR U4424 ( .A(n892), .B(n889), .Z(n890) );
  XOR U4425 ( .A(n872), .B(n857), .Z(n808) );
  XOR U4426 ( .A(n893), .B(n894), .Z(n857) );
  XOR U4427 ( .A(n856), .B(n895), .Z(n893) );
  AND U4428 ( .A(n896), .B(n897), .Z(n895) );
  XOR U4429 ( .A(n894), .B(n898), .Z(n897) );
  OR U4430 ( .A(n899), .B(n900), .Z(n856) );
  XOR U4431 ( .A(n901), .B(n881), .Z(n872) );
  XOR U4432 ( .A(n902), .B(n866), .Z(n861) );
  XNOR U4433 ( .A(n864), .B(n860), .Z(n902) );
  XOR U4434 ( .A(n910), .B(n863), .Z(n864) );
  IV U4435 ( .A(n865), .Z(n863) );
  XOR U4436 ( .A(n918), .B(n867), .Z(n868) );
  IV U4437 ( .A(n869), .Z(n867) );
  XNOR U4438 ( .A(n880), .B(n871), .Z(n901) );
  XOR U4439 ( .A(n932), .B(n885), .Z(n880) );
  XOR U4440 ( .A(n933), .B(n875), .Z(n876) );
  IV U4441 ( .A(n877), .Z(n875) );
  XNOR U4442 ( .A(n884), .B(n879), .Z(n932) );
  XOR U4443 ( .A(n948), .B(n888), .Z(n884) );
  XNOR U4444 ( .A(n887), .B(n883), .Z(n948) );
  XOR U4445 ( .A(n955), .B(n886), .Z(n887) );
  AND U4446 ( .A(n958), .B(n959), .Z(n957) );
  XNOR U4447 ( .A(n956), .B(n960), .Z(n959) );
  XNOR U4448 ( .A(n966), .B(n967), .Z(n809) );
  XNOR U4449 ( .A(n968), .B(n965), .Z(n966) );
  XNOR U4450 ( .A(n931), .B(n900), .Z(n810) );
  XNOR U4451 ( .A(n969), .B(n898), .Z(n900) );
  XOR U4452 ( .A(n896), .B(n899), .Z(n969) );
  OR U4453 ( .A(n973), .B(n974), .Z(n899) );
  XOR U4454 ( .A(n975), .B(n976), .Z(n896) );
  IV U4455 ( .A(n894), .Z(n976) );
  XOR U4456 ( .A(n984), .B(n947), .Z(n931) );
  XOR U4457 ( .A(n985), .B(n913), .Z(n908) );
  XOR U4458 ( .A(n986), .B(n903), .Z(n904) );
  IV U4459 ( .A(n905), .Z(n903) );
  XNOR U4460 ( .A(n912), .B(n907), .Z(n985) );
  XOR U4461 ( .A(n1001), .B(n917), .Z(n912) );
  XNOR U4462 ( .A(n915), .B(n911), .Z(n1001) );
  XOR U4463 ( .A(n1009), .B(n914), .Z(n915) );
  IV U4464 ( .A(n916), .Z(n914) );
  XOR U4465 ( .A(n1017), .B(n925), .Z(n920) );
  XNOR U4466 ( .A(n923), .B(n919), .Z(n1017) );
  XOR U4467 ( .A(n1021), .B(n1022), .Z(n919) );
  AND U4468 ( .A(n1023), .B(n1024), .Z(n1022) );
  XNOR U4469 ( .A(n1021), .B(n1025), .Z(n1023) );
  XOR U4470 ( .A(n1026), .B(n922), .Z(n923) );
  IV U4471 ( .A(n924), .Z(n922) );
  XOR U4472 ( .A(n1034), .B(n926), .Z(n927) );
  IV U4473 ( .A(n928), .Z(n926) );
  XNOR U4474 ( .A(n946), .B(n930), .Z(n984) );
  XOR U4475 ( .A(n1048), .B(n954), .Z(n946) );
  XOR U4476 ( .A(n1049), .B(n940), .Z(n935) );
  XNOR U4477 ( .A(n938), .B(n934), .Z(n1049) );
  XOR U4478 ( .A(n1054), .B(n1055), .Z(n934) );
  AND U4479 ( .A(n1056), .B(n1057), .Z(n1055) );
  XNOR U4480 ( .A(n1054), .B(n1058), .Z(n1056) );
  XOR U4481 ( .A(n1059), .B(n937), .Z(n938) );
  IV U4482 ( .A(n939), .Z(n937) );
  XOR U4483 ( .A(n1067), .B(n941), .Z(n942) );
  IV U4484 ( .A(n943), .Z(n941) );
  XNOR U4485 ( .A(n953), .B(n945), .Z(n1048) );
  XOR U4486 ( .A(n1082), .B(n960), .Z(n953) );
  XOR U4487 ( .A(n1083), .B(n949), .Z(n950) );
  AND U4488 ( .A(n1086), .B(n1087), .Z(n1085) );
  XNOR U4489 ( .A(n1084), .B(n1088), .Z(n1086) );
  XNOR U4490 ( .A(n958), .B(n952), .Z(n1082) );
  XOR U4491 ( .A(n1099), .B(n964), .Z(n958) );
  XNOR U4492 ( .A(n962), .B(n956), .Z(n1099) );
  XOR U4493 ( .A(n1107), .B(n961), .Z(n962) );
  IV U4494 ( .A(n963), .Z(n961) );
  XNOR U4495 ( .A(n1116), .B(n1117), .Z(n811) );
  XNOR U4496 ( .A(n1118), .B(n1115), .Z(n1116) );
  XNOR U4497 ( .A(n1047), .B(n973), .Z(n812) );
  XOR U4498 ( .A(n1119), .B(n979), .Z(n973) );
  XOR U4499 ( .A(n1120), .B(n1121), .Z(n971) );
  IV U4500 ( .A(n970), .Z(n1121) );
  XOR U4501 ( .A(n978), .B(n974), .Z(n1119) );
  OR U4502 ( .A(n1132), .B(n1133), .Z(n974) );
  XOR U4503 ( .A(n1134), .B(n983), .Z(n978) );
  XNOR U4504 ( .A(n981), .B(n977), .Z(n1134) );
  XOR U4505 ( .A(n1142), .B(n980), .Z(n981) );
  IV U4506 ( .A(n982), .Z(n980) );
  XOR U4507 ( .A(n1149), .B(n1081), .Z(n1047) );
  XOR U4508 ( .A(n1150), .B(n1008), .Z(n999) );
  XOR U4509 ( .A(n1151), .B(n993), .Z(n988) );
  XNOR U4510 ( .A(n991), .B(n987), .Z(n1151) );
  XOR U4511 ( .A(n1159), .B(n990), .Z(n991) );
  IV U4512 ( .A(n992), .Z(n990) );
  XOR U4513 ( .A(n1167), .B(n994), .Z(n995) );
  IV U4514 ( .A(n996), .Z(n994) );
  XNOR U4515 ( .A(n1007), .B(n998), .Z(n1150) );
  XOR U4516 ( .A(n1182), .B(n1012), .Z(n1007) );
  XOR U4517 ( .A(n1183), .B(n1002), .Z(n1003) );
  IV U4518 ( .A(n1004), .Z(n1002) );
  XNOR U4519 ( .A(n1011), .B(n1006), .Z(n1182) );
  XOR U4520 ( .A(n1198), .B(n1016), .Z(n1011) );
  XNOR U4521 ( .A(n1014), .B(n1010), .Z(n1198) );
  XOR U4522 ( .A(n1206), .B(n1013), .Z(n1014) );
  IV U4523 ( .A(n1015), .Z(n1013) );
  XOR U4524 ( .A(n1214), .B(n1029), .Z(n1024) );
  XOR U4525 ( .A(n1215), .B(n1018), .Z(n1019) );
  AND U4526 ( .A(n1218), .B(n1219), .Z(n1217) );
  XNOR U4527 ( .A(n1216), .B(n1220), .Z(n1218) );
  XNOR U4528 ( .A(n1028), .B(n1021), .Z(n1214) );
  XOR U4529 ( .A(n1231), .B(n1033), .Z(n1028) );
  XNOR U4530 ( .A(n1031), .B(n1027), .Z(n1231) );
  XOR U4531 ( .A(n1239), .B(n1030), .Z(n1031) );
  IV U4532 ( .A(n1032), .Z(n1030) );
  XOR U4533 ( .A(n1247), .B(n1041), .Z(n1036) );
  XNOR U4534 ( .A(n1039), .B(n1035), .Z(n1247) );
  XOR U4535 ( .A(n1254), .B(n1038), .Z(n1039) );
  IV U4536 ( .A(n1040), .Z(n1038) );
  XOR U4537 ( .A(n1262), .B(n1042), .Z(n1043) );
  IV U4538 ( .A(n1044), .Z(n1042) );
  XNOR U4539 ( .A(n1080), .B(n1046), .Z(n1149) );
  XOR U4540 ( .A(n1276), .B(n1098), .Z(n1080) );
  XOR U4541 ( .A(n1277), .B(n1062), .Z(n1057) );
  XOR U4542 ( .A(n1278), .B(n1050), .Z(n1051) );
  IV U4543 ( .A(n1052), .Z(n1050) );
  XNOR U4544 ( .A(n1061), .B(n1054), .Z(n1277) );
  XOR U4545 ( .A(n1293), .B(n1066), .Z(n1061) );
  XNOR U4546 ( .A(n1064), .B(n1060), .Z(n1293) );
  XOR U4547 ( .A(n1301), .B(n1063), .Z(n1064) );
  IV U4548 ( .A(n1065), .Z(n1063) );
  XOR U4549 ( .A(n1309), .B(n1074), .Z(n1069) );
  XNOR U4550 ( .A(n1072), .B(n1068), .Z(n1309) );
  XOR U4551 ( .A(n1317), .B(n1071), .Z(n1072) );
  IV U4552 ( .A(n1073), .Z(n1071) );
  XOR U4553 ( .A(n1325), .B(n1075), .Z(n1076) );
  IV U4554 ( .A(n1077), .Z(n1075) );
  XNOR U4555 ( .A(n1097), .B(n1079), .Z(n1276) );
  XOR U4556 ( .A(n1339), .B(n1106), .Z(n1097) );
  XOR U4557 ( .A(n1340), .B(n1092), .Z(n1087) );
  XNOR U4558 ( .A(n1090), .B(n1084), .Z(n1340) );
  XOR U4559 ( .A(n1347), .B(n1089), .Z(n1090) );
  IV U4560 ( .A(n1091), .Z(n1089) );
  XOR U4561 ( .A(n1355), .B(n1093), .Z(n1094) );
  AND U4562 ( .A(n1358), .B(n1359), .Z(n1357) );
  XNOR U4563 ( .A(n1356), .B(n1360), .Z(n1358) );
  XNOR U4564 ( .A(n1105), .B(n1096), .Z(n1339) );
  XOR U4565 ( .A(n1371), .B(n1110), .Z(n1105) );
  XOR U4566 ( .A(n1372), .B(n1100), .Z(n1101) );
  IV U4567 ( .A(n1102), .Z(n1100) );
  XNOR U4568 ( .A(n1109), .B(n1104), .Z(n1371) );
  XOR U4569 ( .A(n1386), .B(n1114), .Z(n1109) );
  XNOR U4570 ( .A(n1112), .B(n1108), .Z(n1386) );
  XOR U4571 ( .A(n1394), .B(n1111), .Z(n1112) );
  IV U4572 ( .A(n1113), .Z(n1111) );
  XNOR U4573 ( .A(n1403), .B(n1404), .Z(n813) );
  XNOR U4574 ( .A(n1405), .B(n1402), .Z(n1403) );
  XNOR U4575 ( .A(n1275), .B(n1132), .Z(n814) );
  XOR U4576 ( .A(n1406), .B(n1141), .Z(n1132) );
  XOR U4577 ( .A(n1407), .B(n1128), .Z(n1123) );
  XNOR U4578 ( .A(n1126), .B(n1122), .Z(n1407) );
  XOR U4579 ( .A(n1415), .B(n1125), .Z(n1126) );
  IV U4580 ( .A(n1127), .Z(n1125) );
  XOR U4581 ( .A(n1423), .B(n1129), .Z(n1130) );
  AND U4582 ( .A(n1426), .B(n1427), .Z(n1425) );
  XNOR U4583 ( .A(n1424), .B(n1428), .Z(n1426) );
  XOR U4584 ( .A(n1140), .B(n1133), .Z(n1406) );
  OR U4585 ( .A(n1437), .B(n1438), .Z(n1133) );
  XOR U4586 ( .A(n1439), .B(n1145), .Z(n1140) );
  XOR U4587 ( .A(n1440), .B(n1135), .Z(n1136) );
  IV U4588 ( .A(n1137), .Z(n1135) );
  XNOR U4589 ( .A(n1144), .B(n1139), .Z(n1439) );
  XOR U4590 ( .A(n1455), .B(n1148), .Z(n1144) );
  XNOR U4591 ( .A(n1147), .B(n1143), .Z(n1455) );
  XOR U4592 ( .A(n1462), .B(n1146), .Z(n1147) );
  AND U4593 ( .A(n1465), .B(n1466), .Z(n1464) );
  XNOR U4594 ( .A(n1463), .B(n1467), .Z(n1466) );
  XOR U4595 ( .A(n1472), .B(n1338), .Z(n1275) );
  XOR U4596 ( .A(n1473), .B(n1197), .Z(n1180) );
  XOR U4597 ( .A(n1474), .B(n1162), .Z(n1157) );
  XOR U4598 ( .A(n1475), .B(n1152), .Z(n1153) );
  IV U4599 ( .A(n1154), .Z(n1152) );
  XNOR U4600 ( .A(n1161), .B(n1156), .Z(n1474) );
  XOR U4601 ( .A(n1490), .B(n1166), .Z(n1161) );
  XNOR U4602 ( .A(n1164), .B(n1160), .Z(n1490) );
  XOR U4603 ( .A(n1498), .B(n1163), .Z(n1164) );
  IV U4604 ( .A(n1165), .Z(n1163) );
  XOR U4605 ( .A(n1506), .B(n1174), .Z(n1169) );
  XNOR U4606 ( .A(n1172), .B(n1168), .Z(n1506) );
  XOR U4607 ( .A(n1514), .B(n1171), .Z(n1172) );
  IV U4608 ( .A(n1173), .Z(n1171) );
  XOR U4609 ( .A(n1521), .B(n1175), .Z(n1176) );
  IV U4610 ( .A(n1177), .Z(n1175) );
  XOR U4611 ( .A(n1525), .B(n1526), .Z(n1521) );
  AND U4612 ( .A(n1527), .B(n1528), .Z(n1526) );
  XNOR U4613 ( .A(n1529), .B(n1530), .Z(n1528) );
  XNOR U4614 ( .A(n1196), .B(n1179), .Z(n1473) );
  XOR U4615 ( .A(n1538), .B(n1205), .Z(n1196) );
  XOR U4616 ( .A(n1539), .B(n1190), .Z(n1185) );
  XNOR U4617 ( .A(n1188), .B(n1184), .Z(n1539) );
  XOR U4618 ( .A(n1547), .B(n1187), .Z(n1188) );
  IV U4619 ( .A(n1189), .Z(n1187) );
  XOR U4620 ( .A(n1555), .B(n1191), .Z(n1192) );
  IV U4621 ( .A(n1193), .Z(n1191) );
  XNOR U4622 ( .A(n1204), .B(n1195), .Z(n1538) );
  XOR U4623 ( .A(n1570), .B(n1209), .Z(n1204) );
  XOR U4624 ( .A(n1571), .B(n1199), .Z(n1200) );
  IV U4625 ( .A(n1201), .Z(n1199) );
  XNOR U4626 ( .A(n1208), .B(n1203), .Z(n1570) );
  XOR U4627 ( .A(n1586), .B(n1213), .Z(n1208) );
  XNOR U4628 ( .A(n1211), .B(n1207), .Z(n1586) );
  XOR U4629 ( .A(n1594), .B(n1210), .Z(n1211) );
  IV U4630 ( .A(n1212), .Z(n1210) );
  XOR U4631 ( .A(n1601), .B(n1238), .Z(n1229) );
  XOR U4632 ( .A(n1602), .B(n1224), .Z(n1219) );
  XNOR U4633 ( .A(n1222), .B(n1216), .Z(n1602) );
  XOR U4634 ( .A(n1610), .B(n1221), .Z(n1222) );
  IV U4635 ( .A(n1223), .Z(n1221) );
  XOR U4636 ( .A(n1618), .B(n1225), .Z(n1226) );
  AND U4637 ( .A(n1621), .B(n1622), .Z(n1620) );
  XNOR U4638 ( .A(n1619), .B(n1623), .Z(n1621) );
  XNOR U4639 ( .A(n1237), .B(n1228), .Z(n1601) );
  XOR U4640 ( .A(n1635), .B(n1242), .Z(n1237) );
  XOR U4641 ( .A(n1636), .B(n1232), .Z(n1233) );
  IV U4642 ( .A(n1234), .Z(n1232) );
  XNOR U4643 ( .A(n1241), .B(n1236), .Z(n1635) );
  XOR U4644 ( .A(n1651), .B(n1246), .Z(n1241) );
  XNOR U4645 ( .A(n1244), .B(n1240), .Z(n1651) );
  XOR U4646 ( .A(n1659), .B(n1243), .Z(n1244) );
  IV U4647 ( .A(n1245), .Z(n1243) );
  XOR U4648 ( .A(n1666), .B(n1257), .Z(n1252) );
  XOR U4649 ( .A(n1667), .B(n1248), .Z(n1249) );
  AND U4650 ( .A(n1670), .B(n1671), .Z(n1669) );
  XNOR U4651 ( .A(n1668), .B(n1672), .Z(n1670) );
  XNOR U4652 ( .A(n1256), .B(n1251), .Z(n1666) );
  XOR U4653 ( .A(n1683), .B(n1261), .Z(n1256) );
  XNOR U4654 ( .A(n1259), .B(n1255), .Z(n1683) );
  XOR U4655 ( .A(n1691), .B(n1258), .Z(n1259) );
  IV U4656 ( .A(n1260), .Z(n1258) );
  XOR U4657 ( .A(n1698), .B(n1269), .Z(n1264) );
  XNOR U4658 ( .A(n1267), .B(n1263), .Z(n1698) );
  XOR U4659 ( .A(n1706), .B(n1266), .Z(n1267) );
  IV U4660 ( .A(n1268), .Z(n1266) );
  XNOR U4661 ( .A(n1273), .B(n1714), .Z(n1265) );
  IV U4662 ( .A(n1271), .Z(n1714) );
  XOR U4663 ( .A(n1715), .B(n1270), .Z(n1271) );
  IV U4664 ( .A(n1272), .Z(n1270) );
  XNOR U4665 ( .A(n1337), .B(n1274), .Z(n1472) );
  XOR U4666 ( .A(n1729), .B(n1370), .Z(n1337) );
  XOR U4667 ( .A(n1730), .B(n1300), .Z(n1291) );
  XOR U4668 ( .A(n1731), .B(n1285), .Z(n1280) );
  XNOR U4669 ( .A(n1283), .B(n1279), .Z(n1731) );
  XOR U4670 ( .A(n1736), .B(n1737), .Z(n1279) );
  AND U4671 ( .A(n1738), .B(n1739), .Z(n1737) );
  XNOR U4672 ( .A(n1736), .B(n1740), .Z(n1738) );
  XOR U4673 ( .A(n1741), .B(n1282), .Z(n1283) );
  IV U4674 ( .A(n1284), .Z(n1282) );
  XOR U4675 ( .A(n1749), .B(n1286), .Z(n1287) );
  IV U4676 ( .A(n1288), .Z(n1286) );
  XNOR U4677 ( .A(n1299), .B(n1290), .Z(n1730) );
  XOR U4678 ( .A(n1764), .B(n1304), .Z(n1299) );
  XOR U4679 ( .A(n1765), .B(n1294), .Z(n1295) );
  IV U4680 ( .A(n1296), .Z(n1294) );
  XNOR U4681 ( .A(n1303), .B(n1298), .Z(n1764) );
  XOR U4682 ( .A(n1780), .B(n1308), .Z(n1303) );
  XNOR U4683 ( .A(n1306), .B(n1302), .Z(n1780) );
  XOR U4684 ( .A(n1788), .B(n1305), .Z(n1306) );
  IV U4685 ( .A(n1307), .Z(n1305) );
  XOR U4686 ( .A(n1796), .B(n1320), .Z(n1315) );
  XOR U4687 ( .A(n1797), .B(n1310), .Z(n1311) );
  IV U4688 ( .A(n1312), .Z(n1310) );
  XNOR U4689 ( .A(n1319), .B(n1314), .Z(n1796) );
  XOR U4690 ( .A(n1811), .B(n1324), .Z(n1319) );
  XNOR U4691 ( .A(n1322), .B(n1318), .Z(n1811) );
  XOR U4692 ( .A(n1819), .B(n1321), .Z(n1322) );
  IV U4693 ( .A(n1323), .Z(n1321) );
  XOR U4694 ( .A(n1827), .B(n1332), .Z(n1327) );
  XNOR U4695 ( .A(n1330), .B(n1326), .Z(n1827) );
  XOR U4696 ( .A(n1835), .B(n1329), .Z(n1330) );
  IV U4697 ( .A(n1331), .Z(n1329) );
  XNOR U4698 ( .A(n1335), .B(n1843), .Z(n1328) );
  IV U4699 ( .A(n1334), .Z(n1843) );
  XOR U4700 ( .A(n1844), .B(n1333), .Z(n1334) );
  AND U4701 ( .A(n1847), .B(n1848), .Z(n1846) );
  XNOR U4702 ( .A(n1845), .B(n1849), .Z(n1847) );
  XNOR U4703 ( .A(n1369), .B(n1336), .Z(n1729) );
  XOR U4704 ( .A(n1861), .B(n1385), .Z(n1369) );
  XOR U4705 ( .A(n1862), .B(n1350), .Z(n1345) );
  XOR U4706 ( .A(n1863), .B(n1341), .Z(n1342) );
  AND U4707 ( .A(n1866), .B(n1867), .Z(n1865) );
  XNOR U4708 ( .A(n1864), .B(n1868), .Z(n1866) );
  XNOR U4709 ( .A(n1349), .B(n1344), .Z(n1862) );
  XOR U4710 ( .A(n1880), .B(n1354), .Z(n1349) );
  XNOR U4711 ( .A(n1352), .B(n1348), .Z(n1880) );
  XOR U4712 ( .A(n1888), .B(n1351), .Z(n1352) );
  IV U4713 ( .A(n1353), .Z(n1351) );
  XOR U4714 ( .A(n1896), .B(n1364), .Z(n1359) );
  XNOR U4715 ( .A(n1362), .B(n1356), .Z(n1896) );
  XOR U4716 ( .A(n1904), .B(n1361), .Z(n1362) );
  IV U4717 ( .A(n1363), .Z(n1361) );
  XOR U4718 ( .A(n1912), .B(n1365), .Z(n1366) );
  AND U4719 ( .A(n1915), .B(n1916), .Z(n1914) );
  XNOR U4720 ( .A(n1913), .B(n1917), .Z(n1915) );
  XNOR U4721 ( .A(n1384), .B(n1368), .Z(n1861) );
  XOR U4722 ( .A(n1929), .B(n1393), .Z(n1384) );
  XOR U4723 ( .A(n1930), .B(n1379), .Z(n1374) );
  XNOR U4724 ( .A(n1377), .B(n1373), .Z(n1930) );
  XOR U4725 ( .A(n1938), .B(n1376), .Z(n1377) );
  IV U4726 ( .A(n1378), .Z(n1376) );
  XOR U4727 ( .A(n1946), .B(n1380), .Z(n1381) );
  AND U4728 ( .A(n1949), .B(n1950), .Z(n1948) );
  XNOR U4729 ( .A(n1947), .B(n1951), .Z(n1949) );
  XNOR U4730 ( .A(n1392), .B(n1383), .Z(n1929) );
  XOR U4731 ( .A(n1963), .B(n1397), .Z(n1392) );
  XOR U4732 ( .A(n1964), .B(n1387), .Z(n1388) );
  IV U4733 ( .A(n1389), .Z(n1387) );
  XNOR U4734 ( .A(n1396), .B(n1391), .Z(n1963) );
  XOR U4735 ( .A(n1977), .B(n1401), .Z(n1396) );
  XNOR U4736 ( .A(n1399), .B(n1395), .Z(n1977) );
  XOR U4737 ( .A(n1984), .B(n1398), .Z(n1399) );
  IV U4738 ( .A(n1400), .Z(n1398) );
  XNOR U4739 ( .A(n1993), .B(n1994), .Z(n815) );
  XNOR U4740 ( .A(n1995), .B(n1992), .Z(n1993) );
  XNOR U4741 ( .A(n1728), .B(n1437), .Z(n816) );
  XOR U4742 ( .A(n1996), .B(n1454), .Z(n1437) );
  XOR U4743 ( .A(n1997), .B(n1418), .Z(n1413) );
  XOR U4744 ( .A(n1998), .B(n1408), .Z(n1409) );
  IV U4745 ( .A(n1410), .Z(n1408) );
  XNOR U4746 ( .A(n1417), .B(n1412), .Z(n1997) );
  XOR U4747 ( .A(n2011), .B(n1422), .Z(n1417) );
  XNOR U4748 ( .A(n1420), .B(n1416), .Z(n2011) );
  XOR U4749 ( .A(n2018), .B(n1419), .Z(n1420) );
  IV U4750 ( .A(n1421), .Z(n1419) );
  XOR U4751 ( .A(n2025), .B(n1432), .Z(n1427) );
  XNOR U4752 ( .A(n1430), .B(n1424), .Z(n2025) );
  XOR U4753 ( .A(n2032), .B(n1429), .Z(n1430) );
  IV U4754 ( .A(n1431), .Z(n1429) );
  XOR U4755 ( .A(n2039), .B(n1433), .Z(n1434) );
  IV U4756 ( .A(n1435), .Z(n1433) );
  XOR U4757 ( .A(n1453), .B(n1438), .Z(n1996) );
  OR U4758 ( .A(n2049), .B(n2050), .Z(n1438) );
  XOR U4759 ( .A(n2051), .B(n1461), .Z(n1453) );
  XOR U4760 ( .A(n2052), .B(n1447), .Z(n1442) );
  XNOR U4761 ( .A(n1445), .B(n1441), .Z(n2052) );
  XOR U4762 ( .A(n2059), .B(n1444), .Z(n1445) );
  IV U4763 ( .A(n1446), .Z(n1444) );
  XOR U4764 ( .A(n2066), .B(n1448), .Z(n1449) );
  IV U4765 ( .A(n1450), .Z(n1448) );
  XNOR U4766 ( .A(n1460), .B(n1452), .Z(n2051) );
  XOR U4767 ( .A(n2079), .B(n1467), .Z(n1460) );
  XOR U4768 ( .A(n2080), .B(n1456), .Z(n1457) );
  ANDN U4769 ( .B(n2083), .A(n2084), .Z(n2082) );
  XOR U4770 ( .A(n2081), .B(n2085), .Z(n2083) );
  XNOR U4771 ( .A(n1465), .B(n1459), .Z(n2079) );
  XOR U4772 ( .A(n2095), .B(n1471), .Z(n1465) );
  XNOR U4773 ( .A(n1469), .B(n1463), .Z(n2095) );
  XOR U4774 ( .A(n2102), .B(n1468), .Z(n1469) );
  IV U4775 ( .A(n1470), .Z(n1468) );
  XOR U4776 ( .A(n2109), .B(n1860), .Z(n1728) );
  XOR U4777 ( .A(n2110), .B(n1569), .Z(n1536) );
  XOR U4778 ( .A(n2111), .B(n1497), .Z(n1488) );
  XOR U4779 ( .A(n2112), .B(n1482), .Z(n1477) );
  XNOR U4780 ( .A(n1480), .B(n1476), .Z(n2112) );
  XOR U4781 ( .A(n2119), .B(n1479), .Z(n1480) );
  IV U4782 ( .A(n1481), .Z(n1479) );
  XOR U4783 ( .A(n2126), .B(n1483), .Z(n1484) );
  IV U4784 ( .A(n1485), .Z(n1483) );
  XNOR U4785 ( .A(n1496), .B(n1487), .Z(n2111) );
  XOR U4786 ( .A(n2139), .B(n1501), .Z(n1496) );
  XOR U4787 ( .A(n2140), .B(n1491), .Z(n1492) );
  IV U4788 ( .A(n1493), .Z(n1491) );
  XNOR U4789 ( .A(n1500), .B(n1495), .Z(n2139) );
  XOR U4790 ( .A(n2153), .B(n1505), .Z(n1500) );
  XNOR U4791 ( .A(n1503), .B(n1499), .Z(n2153) );
  XOR U4792 ( .A(n2160), .B(n1502), .Z(n1503) );
  IV U4793 ( .A(n1504), .Z(n1502) );
  XOR U4794 ( .A(n2167), .B(n1516), .Z(n1512) );
  XOR U4795 ( .A(n2168), .B(n1507), .Z(n1508) );
  IV U4796 ( .A(n1509), .Z(n1507) );
  XNOR U4797 ( .A(n1515), .B(n1511), .Z(n2167) );
  XOR U4798 ( .A(n2181), .B(n1520), .Z(n1515) );
  XOR U4799 ( .A(n2188), .B(n1517), .Z(n1518) );
  IV U4800 ( .A(n1519), .Z(n1517) );
  XOR U4801 ( .A(n2195), .B(n1530), .Z(n1523) );
  XNOR U4802 ( .A(n1527), .B(n1522), .Z(n2195) );
  XOR U4803 ( .A(n2202), .B(n1525), .Z(n1527) );
  IV U4804 ( .A(n1529), .Z(n1525) );
  XOR U4805 ( .A(n2209), .B(n1531), .Z(n1532) );
  IV U4806 ( .A(n1533), .Z(n1531) );
  XNOR U4807 ( .A(n1568), .B(n1535), .Z(n2110) );
  XOR U4808 ( .A(n2222), .B(n1585), .Z(n1568) );
  XOR U4809 ( .A(n2223), .B(n1550), .Z(n1545) );
  XOR U4810 ( .A(n2224), .B(n1540), .Z(n1541) );
  IV U4811 ( .A(n1542), .Z(n1540) );
  XNOR U4812 ( .A(n1549), .B(n1544), .Z(n2223) );
  XOR U4813 ( .A(n2237), .B(n1554), .Z(n1549) );
  XNOR U4814 ( .A(n1552), .B(n1548), .Z(n2237) );
  XOR U4815 ( .A(n2244), .B(n1551), .Z(n1552) );
  IV U4816 ( .A(n1553), .Z(n1551) );
  XOR U4817 ( .A(n2251), .B(n1562), .Z(n1557) );
  XNOR U4818 ( .A(n1560), .B(n1556), .Z(n2251) );
  XOR U4819 ( .A(n2258), .B(n1559), .Z(n1560) );
  IV U4820 ( .A(n1561), .Z(n1559) );
  XOR U4821 ( .A(n2265), .B(n1563), .Z(n1564) );
  IV U4822 ( .A(n1565), .Z(n1563) );
  XNOR U4823 ( .A(n1584), .B(n1567), .Z(n2222) );
  XOR U4824 ( .A(n2278), .B(n1593), .Z(n1584) );
  XOR U4825 ( .A(n2279), .B(n1578), .Z(n1573) );
  XNOR U4826 ( .A(n1576), .B(n1572), .Z(n2279) );
  XOR U4827 ( .A(n2286), .B(n1575), .Z(n1576) );
  IV U4828 ( .A(n1577), .Z(n1575) );
  XOR U4829 ( .A(n2293), .B(n1579), .Z(n1580) );
  IV U4830 ( .A(n1581), .Z(n1579) );
  XNOR U4831 ( .A(n1592), .B(n1583), .Z(n2278) );
  XOR U4832 ( .A(n2306), .B(n1596), .Z(n1592) );
  XOR U4833 ( .A(n2307), .B(n1587), .Z(n1588) );
  IV U4834 ( .A(n1589), .Z(n1587) );
  XNOR U4835 ( .A(n1595), .B(n1591), .Z(n2306) );
  XOR U4836 ( .A(n2320), .B(n1600), .Z(n1595) );
  XOR U4837 ( .A(n2327), .B(n1597), .Z(n1598) );
  IV U4838 ( .A(n1599), .Z(n1597) );
  XOR U4839 ( .A(n2334), .B(n1650), .Z(n1633) );
  XOR U4840 ( .A(n2335), .B(n1613), .Z(n1608) );
  XOR U4841 ( .A(n2336), .B(n1603), .Z(n1604) );
  IV U4842 ( .A(n1605), .Z(n1603) );
  XNOR U4843 ( .A(n1612), .B(n1607), .Z(n2335) );
  XOR U4844 ( .A(n2349), .B(n1617), .Z(n1612) );
  XNOR U4845 ( .A(n1615), .B(n1611), .Z(n2349) );
  XOR U4846 ( .A(n2356), .B(n1614), .Z(n1615) );
  IV U4847 ( .A(n1616), .Z(n1614) );
  XOR U4848 ( .A(n2363), .B(n1627), .Z(n1622) );
  XNOR U4849 ( .A(n1625), .B(n1619), .Z(n2363) );
  XOR U4850 ( .A(n2370), .B(n1624), .Z(n1625) );
  IV U4851 ( .A(n1626), .Z(n1624) );
  XNOR U4852 ( .A(n1631), .B(n2377), .Z(n1623) );
  IV U4853 ( .A(n1629), .Z(n2377) );
  XOR U4854 ( .A(n2378), .B(n1628), .Z(n1629) );
  IV U4855 ( .A(n1630), .Z(n1628) );
  XNOR U4856 ( .A(n1649), .B(n1632), .Z(n2334) );
  XOR U4857 ( .A(n2391), .B(n1658), .Z(n1649) );
  XOR U4858 ( .A(n2392), .B(n1643), .Z(n1638) );
  XNOR U4859 ( .A(n1641), .B(n1637), .Z(n2392) );
  XOR U4860 ( .A(n2399), .B(n1640), .Z(n1641) );
  IV U4861 ( .A(n1642), .Z(n1640) );
  XOR U4862 ( .A(n2406), .B(n1644), .Z(n1645) );
  IV U4863 ( .A(n1646), .Z(n1644) );
  XNOR U4864 ( .A(n1657), .B(n1648), .Z(n2391) );
  XOR U4865 ( .A(n2419), .B(n1661), .Z(n1657) );
  XOR U4866 ( .A(n2420), .B(n1652), .Z(n1653) );
  IV U4867 ( .A(n1654), .Z(n1652) );
  XNOR U4868 ( .A(n1660), .B(n1656), .Z(n2419) );
  XOR U4869 ( .A(n2433), .B(n1665), .Z(n1660) );
  XOR U4870 ( .A(n2440), .B(n1662), .Z(n1663) );
  IV U4871 ( .A(n1664), .Z(n1662) );
  XOR U4872 ( .A(n2447), .B(n1690), .Z(n1681) );
  XOR U4873 ( .A(n2448), .B(n1676), .Z(n1671) );
  XNOR U4874 ( .A(n1674), .B(n1668), .Z(n2448) );
  XOR U4875 ( .A(n2455), .B(n1673), .Z(n1674) );
  IV U4876 ( .A(n1675), .Z(n1673) );
  XOR U4877 ( .A(n2462), .B(n1677), .Z(n1678) );
  ANDN U4878 ( .B(n2465), .A(n2466), .Z(n2464) );
  XOR U4879 ( .A(n2463), .B(n2467), .Z(n2465) );
  XNOR U4880 ( .A(n1689), .B(n1680), .Z(n2447) );
  XOR U4881 ( .A(n2477), .B(n1693), .Z(n1689) );
  XOR U4882 ( .A(n2478), .B(n1684), .Z(n1685) );
  IV U4883 ( .A(n1686), .Z(n1684) );
  XNOR U4884 ( .A(n1692), .B(n1688), .Z(n2477) );
  XOR U4885 ( .A(n2491), .B(n1697), .Z(n1692) );
  XOR U4886 ( .A(n2498), .B(n1694), .Z(n1695) );
  IV U4887 ( .A(n1696), .Z(n1694) );
  XOR U4888 ( .A(n2505), .B(n1709), .Z(n1704) );
  XOR U4889 ( .A(n2506), .B(n1699), .Z(n1700) );
  IV U4890 ( .A(n1701), .Z(n1699) );
  XNOR U4891 ( .A(n1708), .B(n1703), .Z(n2505) );
  XOR U4892 ( .A(n2519), .B(n1713), .Z(n1708) );
  XNOR U4893 ( .A(n1711), .B(n1707), .Z(n2519) );
  XOR U4894 ( .A(n2526), .B(n1710), .Z(n1711) );
  IV U4895 ( .A(n1712), .Z(n1710) );
  XOR U4896 ( .A(n2533), .B(n1722), .Z(n1717) );
  XNOR U4897 ( .A(n1720), .B(n1716), .Z(n2533) );
  XOR U4898 ( .A(n2540), .B(n1719), .Z(n1720) );
  IV U4899 ( .A(n1721), .Z(n1719) );
  XOR U4900 ( .A(n2547), .B(n1723), .Z(n1724) );
  IV U4901 ( .A(n1725), .Z(n1723) );
  XNOR U4902 ( .A(n1859), .B(n1727), .Z(n2109) );
  XOR U4903 ( .A(n2559), .B(n1928), .Z(n1859) );
  XOR U4904 ( .A(n2560), .B(n1779), .Z(n1762) );
  XOR U4905 ( .A(n2561), .B(n1744), .Z(n1739) );
  XOR U4906 ( .A(n2562), .B(n1732), .Z(n1733) );
  IV U4907 ( .A(n1734), .Z(n1732) );
  XNOR U4908 ( .A(n1743), .B(n1736), .Z(n2561) );
  XOR U4909 ( .A(n2575), .B(n1748), .Z(n1743) );
  XNOR U4910 ( .A(n1746), .B(n1742), .Z(n2575) );
  XOR U4911 ( .A(n2582), .B(n1745), .Z(n1746) );
  IV U4912 ( .A(n1747), .Z(n1745) );
  XOR U4913 ( .A(n2589), .B(n1756), .Z(n1751) );
  XNOR U4914 ( .A(n1754), .B(n1750), .Z(n2589) );
  XOR U4915 ( .A(n2596), .B(n1753), .Z(n1754) );
  IV U4916 ( .A(n1755), .Z(n1753) );
  XOR U4917 ( .A(n2603), .B(n1757), .Z(n1758) );
  IV U4918 ( .A(n1759), .Z(n1757) );
  XNOR U4919 ( .A(n1778), .B(n1761), .Z(n2560) );
  XOR U4920 ( .A(n2616), .B(n1787), .Z(n1778) );
  XOR U4921 ( .A(n2617), .B(n1772), .Z(n1767) );
  XNOR U4922 ( .A(n1770), .B(n1766), .Z(n2617) );
  XOR U4923 ( .A(n2624), .B(n1769), .Z(n1770) );
  IV U4924 ( .A(n1771), .Z(n1769) );
  XOR U4925 ( .A(n2631), .B(n1773), .Z(n1774) );
  IV U4926 ( .A(n1775), .Z(n1773) );
  XNOR U4927 ( .A(n1786), .B(n1777), .Z(n2616) );
  XOR U4928 ( .A(n2644), .B(n1791), .Z(n1786) );
  XOR U4929 ( .A(n2645), .B(n1781), .Z(n1782) );
  IV U4930 ( .A(n1783), .Z(n1781) );
  XNOR U4931 ( .A(n1790), .B(n1785), .Z(n2644) );
  XOR U4932 ( .A(n2658), .B(n1795), .Z(n1790) );
  XNOR U4933 ( .A(n1793), .B(n1789), .Z(n2658) );
  XOR U4934 ( .A(n2665), .B(n1792), .Z(n1793) );
  IV U4935 ( .A(n1794), .Z(n1792) );
  XOR U4936 ( .A(n2672), .B(n1818), .Z(n1809) );
  XOR U4937 ( .A(n2673), .B(n1804), .Z(n1799) );
  XNOR U4938 ( .A(n1802), .B(n1798), .Z(n2673) );
  XOR U4939 ( .A(n2680), .B(n1801), .Z(n1802) );
  IV U4940 ( .A(n1803), .Z(n1801) );
  XOR U4941 ( .A(n2687), .B(n1805), .Z(n1806) );
  ANDN U4942 ( .B(n2690), .A(n2691), .Z(n2689) );
  XOR U4943 ( .A(n2688), .B(n2692), .Z(n2690) );
  XNOR U4944 ( .A(n1817), .B(n1808), .Z(n2672) );
  XOR U4945 ( .A(n2702), .B(n1822), .Z(n1817) );
  XOR U4946 ( .A(n2703), .B(n1812), .Z(n1813) );
  IV U4947 ( .A(n1814), .Z(n1812) );
  XNOR U4948 ( .A(n1821), .B(n1816), .Z(n2702) );
  XOR U4949 ( .A(n2716), .B(n1826), .Z(n1821) );
  XNOR U4950 ( .A(n1824), .B(n1820), .Z(n2716) );
  XOR U4951 ( .A(n2723), .B(n1823), .Z(n1824) );
  IV U4952 ( .A(n1825), .Z(n1823) );
  XOR U4953 ( .A(n2730), .B(n1838), .Z(n1833) );
  XOR U4954 ( .A(n2731), .B(n1828), .Z(n1829) );
  IV U4955 ( .A(n1830), .Z(n1828) );
  XNOR U4956 ( .A(n1837), .B(n1832), .Z(n2730) );
  XOR U4957 ( .A(n2744), .B(n1842), .Z(n1837) );
  XNOR U4958 ( .A(n1840), .B(n1836), .Z(n2744) );
  XOR U4959 ( .A(n2751), .B(n1839), .Z(n1840) );
  IV U4960 ( .A(n1841), .Z(n1839) );
  XOR U4961 ( .A(n2758), .B(n1853), .Z(n1848) );
  XNOR U4962 ( .A(n1851), .B(n1845), .Z(n2758) );
  XOR U4963 ( .A(n2765), .B(n1850), .Z(n1851) );
  IV U4964 ( .A(n1852), .Z(n1850) );
  XOR U4965 ( .A(n2772), .B(n1854), .Z(n1855) );
  IV U4966 ( .A(n1856), .Z(n1854) );
  XNOR U4967 ( .A(n1927), .B(n1858), .Z(n2559) );
  XOR U4968 ( .A(n2785), .B(n1962), .Z(n1927) );
  XOR U4969 ( .A(n2786), .B(n1887), .Z(n1878) );
  XOR U4970 ( .A(n2787), .B(n1872), .Z(n1867) );
  XNOR U4971 ( .A(n1870), .B(n1864), .Z(n2787) );
  XOR U4972 ( .A(n2794), .B(n1869), .Z(n1870) );
  IV U4973 ( .A(n1871), .Z(n1869) );
  XOR U4974 ( .A(n2801), .B(n1873), .Z(n1874) );
  IV U4975 ( .A(n1875), .Z(n1873) );
  XNOR U4976 ( .A(n1886), .B(n1877), .Z(n2786) );
  XOR U4977 ( .A(n2814), .B(n1891), .Z(n1886) );
  XOR U4978 ( .A(n2815), .B(n1881), .Z(n1882) );
  IV U4979 ( .A(n1883), .Z(n1881) );
  XNOR U4980 ( .A(n1890), .B(n1885), .Z(n2814) );
  XOR U4981 ( .A(n2828), .B(n1895), .Z(n1890) );
  XNOR U4982 ( .A(n1893), .B(n1889), .Z(n2828) );
  XOR U4983 ( .A(n2835), .B(n1892), .Z(n1893) );
  IV U4984 ( .A(n1894), .Z(n1892) );
  XOR U4985 ( .A(n2842), .B(n1907), .Z(n1902) );
  XOR U4986 ( .A(n2843), .B(n1897), .Z(n1898) );
  IV U4987 ( .A(n1899), .Z(n1897) );
  XNOR U4988 ( .A(n1906), .B(n1901), .Z(n2842) );
  XOR U4989 ( .A(n2856), .B(n1911), .Z(n1906) );
  XNOR U4990 ( .A(n1909), .B(n1905), .Z(n2856) );
  XOR U4991 ( .A(n2863), .B(n1908), .Z(n1909) );
  IV U4992 ( .A(n1910), .Z(n1908) );
  XOR U4993 ( .A(n2870), .B(n1921), .Z(n1916) );
  XNOR U4994 ( .A(n1919), .B(n1913), .Z(n2870) );
  XNOR U4995 ( .A(n2874), .B(n2875), .Z(n1913) );
  ANDN U4996 ( .B(n2876), .A(n2877), .Z(n2875) );
  XOR U4997 ( .A(n2874), .B(n2878), .Z(n2876) );
  XOR U4998 ( .A(n2879), .B(n1918), .Z(n1919) );
  IV U4999 ( .A(n1920), .Z(n1918) );
  XOR U5000 ( .A(n2883), .B(n2884), .Z(n2879) );
  ANDN U5001 ( .B(n2885), .A(n2886), .Z(n2884) );
  XOR U5002 ( .A(n2883), .B(n2887), .Z(n2885) );
  XOR U5003 ( .A(n2888), .B(n1922), .Z(n1923) );
  IV U5004 ( .A(n1924), .Z(n1922) );
  XNOR U5005 ( .A(n1961), .B(n1926), .Z(n2785) );
  XOR U5006 ( .A(n2901), .B(n1976), .Z(n1961) );
  XOR U5007 ( .A(n2902), .B(n1941), .Z(n1936) );
  XOR U5008 ( .A(n2903), .B(n1931), .Z(n1932) );
  IV U5009 ( .A(n1933), .Z(n1931) );
  XNOR U5010 ( .A(n1940), .B(n1935), .Z(n2902) );
  XOR U5011 ( .A(n2916), .B(n1945), .Z(n1940) );
  XNOR U5012 ( .A(n1943), .B(n1939), .Z(n2916) );
  XOR U5013 ( .A(n2923), .B(n1942), .Z(n1943) );
  IV U5014 ( .A(n1944), .Z(n1942) );
  XOR U5015 ( .A(n2930), .B(n1955), .Z(n1950) );
  XNOR U5016 ( .A(n1953), .B(n1947), .Z(n2930) );
  XOR U5017 ( .A(n2937), .B(n1952), .Z(n1953) );
  IV U5018 ( .A(n1954), .Z(n1952) );
  XOR U5019 ( .A(n2944), .B(n1956), .Z(n1957) );
  IV U5020 ( .A(n1958), .Z(n1956) );
  XNOR U5021 ( .A(n1975), .B(n1960), .Z(n2901) );
  XOR U5022 ( .A(n2957), .B(n1983), .Z(n1975) );
  XOR U5023 ( .A(n2958), .B(n1971), .Z(n1966) );
  XNOR U5024 ( .A(n1969), .B(n1965), .Z(n2958) );
  XOR U5025 ( .A(n2965), .B(n1968), .Z(n1969) );
  IV U5026 ( .A(n1970), .Z(n1968) );
  XOR U5027 ( .A(n2972), .B(n1972), .Z(n1973) );
  ANDN U5028 ( .B(n2975), .A(n2976), .Z(n2974) );
  XOR U5029 ( .A(n2973), .B(n2977), .Z(n2975) );
  XOR U5030 ( .A(n2987), .B(n1987), .Z(n1982) );
  XOR U5031 ( .A(n2988), .B(n1978), .Z(n1979) );
  ANDN U5032 ( .B(n2991), .A(n2992), .Z(n2990) );
  XOR U5033 ( .A(n2989), .B(n2993), .Z(n2991) );
  XNOR U5034 ( .A(n1986), .B(n1981), .Z(n2987) );
  XOR U5035 ( .A(n3003), .B(n1991), .Z(n1986) );
  XNOR U5036 ( .A(n1989), .B(n1985), .Z(n3003) );
  XOR U5037 ( .A(n3010), .B(n1988), .Z(n1989) );
  IV U5038 ( .A(n1990), .Z(n1988) );
  XOR U5039 ( .A(n3020), .B(n3021), .Z(n819) );
  AND U5040 ( .A(n823), .B(n3022), .Z(n3021) );
  XOR U5041 ( .A(n3023), .B(n822), .Z(n3022) );
  XOR U5042 ( .A(n3027), .B(n3020), .Z(n823) );
  IV U5043 ( .A(n3023), .Z(n3020) );
  XOR U5044 ( .A(n3033), .B(n3034), .Z(n3025) );
  IV U5045 ( .A(n3024), .Z(n3034) );
  XOR U5046 ( .A(n3046), .B(n3031), .Z(n834) );
  XNOR U5047 ( .A(n3029), .B(n3032), .Z(n3046) );
  XOR U5048 ( .A(n3051), .B(n3028), .Z(n3029) );
  IV U5049 ( .A(n3030), .Z(n3028) );
  XOR U5050 ( .A(n3060), .B(n3041), .Z(n3036) );
  XNOR U5051 ( .A(n3039), .B(n3035), .Z(n3060) );
  XOR U5052 ( .A(n3068), .B(n3038), .Z(n3039) );
  IV U5053 ( .A(n3040), .Z(n3038) );
  XOR U5054 ( .A(n3076), .B(n3042), .Z(n3043) );
  IV U5055 ( .A(n3044), .Z(n3042) );
  XOR U5056 ( .A(n3088), .B(n3054), .Z(n855) );
  XOR U5057 ( .A(n3089), .B(n3047), .Z(n3048) );
  IV U5058 ( .A(n3049), .Z(n3047) );
  XNOR U5059 ( .A(n3053), .B(n3059), .Z(n3088) );
  XOR U5060 ( .A(n3101), .B(n3058), .Z(n3053) );
  XNOR U5061 ( .A(n3056), .B(n3052), .Z(n3101) );
  XOR U5062 ( .A(n3108), .B(n3055), .Z(n3056) );
  IV U5063 ( .A(n3057), .Z(n3055) );
  XOR U5064 ( .A(n3117), .B(n3071), .Z(n3066) );
  XOR U5065 ( .A(n3118), .B(n3061), .Z(n3062) );
  IV U5066 ( .A(n3063), .Z(n3061) );
  XNOR U5067 ( .A(n3070), .B(n3065), .Z(n3117) );
  XOR U5068 ( .A(n3133), .B(n3075), .Z(n3070) );
  XNOR U5069 ( .A(n3073), .B(n3069), .Z(n3133) );
  XOR U5070 ( .A(n3141), .B(n3072), .Z(n3073) );
  IV U5071 ( .A(n3074), .Z(n3072) );
  XOR U5072 ( .A(n3149), .B(n3083), .Z(n3078) );
  XNOR U5073 ( .A(n3081), .B(n3077), .Z(n3149) );
  XOR U5074 ( .A(n3157), .B(n3080), .Z(n3081) );
  IV U5075 ( .A(n3082), .Z(n3080) );
  XOR U5076 ( .A(n3165), .B(n3084), .Z(n3085) );
  IV U5077 ( .A(n3086), .Z(n3084) );
  XOR U5078 ( .A(n3177), .B(n3107), .Z(n892) );
  XOR U5079 ( .A(n3178), .B(n3096), .Z(n3091) );
  XNOR U5080 ( .A(n3094), .B(n3090), .Z(n3178) );
  XOR U5081 ( .A(n3186), .B(n3093), .Z(n3094) );
  IV U5082 ( .A(n3095), .Z(n3093) );
  XOR U5083 ( .A(n3194), .B(n3097), .Z(n3098) );
  IV U5084 ( .A(n3099), .Z(n3097) );
  XNOR U5085 ( .A(n3106), .B(n3116), .Z(n3177) );
  XOR U5086 ( .A(n3206), .B(n3111), .Z(n3106) );
  XOR U5087 ( .A(n3207), .B(n3102), .Z(n3103) );
  AND U5088 ( .A(n3210), .B(n3211), .Z(n3209) );
  XNOR U5089 ( .A(n3208), .B(n3212), .Z(n3210) );
  XNOR U5090 ( .A(n3110), .B(n3105), .Z(n3206) );
  XOR U5091 ( .A(n3223), .B(n3115), .Z(n3110) );
  XNOR U5092 ( .A(n3113), .B(n3109), .Z(n3223) );
  XOR U5093 ( .A(n3231), .B(n3112), .Z(n3113) );
  IV U5094 ( .A(n3114), .Z(n3112) );
  XOR U5095 ( .A(n3240), .B(n3140), .Z(n3131) );
  XOR U5096 ( .A(n3241), .B(n3125), .Z(n3120) );
  XNOR U5097 ( .A(n3123), .B(n3119), .Z(n3241) );
  XOR U5098 ( .A(n3248), .B(n3122), .Z(n3123) );
  IV U5099 ( .A(n3124), .Z(n3122) );
  XOR U5100 ( .A(n3256), .B(n3126), .Z(n3127) );
  IV U5101 ( .A(n3128), .Z(n3126) );
  XNOR U5102 ( .A(n3139), .B(n3130), .Z(n3240) );
  XOR U5103 ( .A(n3271), .B(n3144), .Z(n3139) );
  XOR U5104 ( .A(n3272), .B(n3134), .Z(n3135) );
  IV U5105 ( .A(n3136), .Z(n3134) );
  XNOR U5106 ( .A(n3143), .B(n3138), .Z(n3271) );
  XOR U5107 ( .A(n3287), .B(n3148), .Z(n3143) );
  XNOR U5108 ( .A(n3146), .B(n3142), .Z(n3287) );
  XOR U5109 ( .A(n3294), .B(n3145), .Z(n3146) );
  IV U5110 ( .A(n3147), .Z(n3145) );
  XOR U5111 ( .A(n3302), .B(n3160), .Z(n3155) );
  XOR U5112 ( .A(n3303), .B(n3150), .Z(n3151) );
  IV U5113 ( .A(n3152), .Z(n3150) );
  XNOR U5114 ( .A(n3159), .B(n3154), .Z(n3302) );
  XOR U5115 ( .A(n3318), .B(n3164), .Z(n3159) );
  XNOR U5116 ( .A(n3162), .B(n3158), .Z(n3318) );
  XOR U5117 ( .A(n3325), .B(n3161), .Z(n3162) );
  IV U5118 ( .A(n3163), .Z(n3161) );
  XOR U5119 ( .A(n3333), .B(n3172), .Z(n3167) );
  XNOR U5120 ( .A(n3170), .B(n3166), .Z(n3333) );
  XOR U5121 ( .A(n3340), .B(n3169), .Z(n3170) );
  IV U5122 ( .A(n3171), .Z(n3169) );
  XOR U5123 ( .A(n3348), .B(n3173), .Z(n3174) );
  IV U5124 ( .A(n3175), .Z(n3173) );
  XOR U5125 ( .A(n3352), .B(n3353), .Z(n3348) );
  AND U5126 ( .A(n3354), .B(n3355), .Z(n3353) );
  XNOR U5127 ( .A(n3356), .B(n3357), .Z(n3355) );
  XOR U5128 ( .A(n3362), .B(n3222), .Z(n968) );
  XOR U5129 ( .A(n3363), .B(n3189), .Z(n3184) );
  XOR U5130 ( .A(n3364), .B(n3179), .Z(n3180) );
  IV U5131 ( .A(n3181), .Z(n3179) );
  XNOR U5132 ( .A(n3188), .B(n3183), .Z(n3363) );
  XOR U5133 ( .A(n3379), .B(n3193), .Z(n3188) );
  XNOR U5134 ( .A(n3191), .B(n3187), .Z(n3379) );
  XOR U5135 ( .A(n3386), .B(n3190), .Z(n3191) );
  IV U5136 ( .A(n3192), .Z(n3190) );
  XOR U5137 ( .A(n3394), .B(n3201), .Z(n3196) );
  XNOR U5138 ( .A(n3199), .B(n3195), .Z(n3394) );
  XOR U5139 ( .A(n3402), .B(n3198), .Z(n3199) );
  IV U5140 ( .A(n3200), .Z(n3198) );
  XOR U5141 ( .A(n3410), .B(n3202), .Z(n3203) );
  IV U5142 ( .A(n3204), .Z(n3202) );
  XNOR U5143 ( .A(n3221), .B(n3239), .Z(n3362) );
  XOR U5144 ( .A(n3421), .B(n3230), .Z(n3221) );
  XOR U5145 ( .A(n3422), .B(n3216), .Z(n3211) );
  XNOR U5146 ( .A(n3214), .B(n3208), .Z(n3422) );
  XOR U5147 ( .A(n3430), .B(n3213), .Z(n3214) );
  IV U5148 ( .A(n3215), .Z(n3213) );
  XOR U5149 ( .A(n3438), .B(n3217), .Z(n3218) );
  AND U5150 ( .A(n3441), .B(n3442), .Z(n3440) );
  XNOR U5151 ( .A(n3439), .B(n3443), .Z(n3441) );
  XNOR U5152 ( .A(n3229), .B(n3220), .Z(n3421) );
  XOR U5153 ( .A(n3454), .B(n3234), .Z(n3229) );
  XOR U5154 ( .A(n3455), .B(n3224), .Z(n3225) );
  IV U5155 ( .A(n3226), .Z(n3224) );
  XNOR U5156 ( .A(n3233), .B(n3228), .Z(n3454) );
  XOR U5157 ( .A(n3469), .B(n3238), .Z(n3233) );
  XNOR U5158 ( .A(n3236), .B(n3232), .Z(n3469) );
  XOR U5159 ( .A(n3476), .B(n3235), .Z(n3236) );
  IV U5160 ( .A(n3237), .Z(n3235) );
  XOR U5161 ( .A(n3485), .B(n3286), .Z(n3269) );
  XOR U5162 ( .A(n3486), .B(n3251), .Z(n3246) );
  XOR U5163 ( .A(n3487), .B(n3242), .Z(n3243) );
  AND U5164 ( .A(n3490), .B(n3491), .Z(n3489) );
  XNOR U5165 ( .A(n3488), .B(n3492), .Z(n3490) );
  XNOR U5166 ( .A(n3250), .B(n3245), .Z(n3486) );
  XOR U5167 ( .A(n3503), .B(n3255), .Z(n3250) );
  XNOR U5168 ( .A(n3253), .B(n3249), .Z(n3503) );
  XOR U5169 ( .A(n3510), .B(n3252), .Z(n3253) );
  IV U5170 ( .A(n3254), .Z(n3252) );
  XOR U5171 ( .A(n3518), .B(n3263), .Z(n3258) );
  XNOR U5172 ( .A(n3261), .B(n3257), .Z(n3518) );
  XOR U5173 ( .A(n3526), .B(n3260), .Z(n3261) );
  IV U5174 ( .A(n3262), .Z(n3260) );
  XOR U5175 ( .A(n3534), .B(n3264), .Z(n3265) );
  IV U5176 ( .A(n3266), .Z(n3264) );
  XOR U5177 ( .A(n3535), .B(n3536), .Z(n3266) );
  AND U5178 ( .A(n3537), .B(n3538), .Z(n3536) );
  XNOR U5179 ( .A(n3535), .B(n3539), .Z(n3537) );
  XNOR U5180 ( .A(n3285), .B(n3268), .Z(n3485) );
  XOR U5181 ( .A(n3551), .B(n3293), .Z(n3285) );
  XOR U5182 ( .A(n3552), .B(n3279), .Z(n3274) );
  XNOR U5183 ( .A(n3277), .B(n3273), .Z(n3552) );
  XOR U5184 ( .A(n3559), .B(n3276), .Z(n3277) );
  IV U5185 ( .A(n3278), .Z(n3276) );
  XOR U5186 ( .A(n3567), .B(n3280), .Z(n3281) );
  IV U5187 ( .A(n3282), .Z(n3280) );
  XNOR U5188 ( .A(n3292), .B(n3284), .Z(n3551) );
  XOR U5189 ( .A(n3582), .B(n3297), .Z(n3292) );
  XOR U5190 ( .A(n3583), .B(n3288), .Z(n3289) );
  AND U5191 ( .A(n3586), .B(n3587), .Z(n3585) );
  XNOR U5192 ( .A(n3584), .B(n3588), .Z(n3586) );
  XNOR U5193 ( .A(n3296), .B(n3291), .Z(n3582) );
  XOR U5194 ( .A(n3599), .B(n3301), .Z(n3296) );
  XNOR U5195 ( .A(n3299), .B(n3295), .Z(n3599) );
  XOR U5196 ( .A(n3606), .B(n3298), .Z(n3299) );
  IV U5197 ( .A(n3300), .Z(n3298) );
  XOR U5198 ( .A(n3614), .B(n3324), .Z(n3316) );
  XOR U5199 ( .A(n3615), .B(n3310), .Z(n3305) );
  XNOR U5200 ( .A(n3308), .B(n3304), .Z(n3615) );
  XOR U5201 ( .A(n3623), .B(n3307), .Z(n3308) );
  IV U5202 ( .A(n3309), .Z(n3307) );
  XOR U5203 ( .A(n3631), .B(n3311), .Z(n3312) );
  IV U5204 ( .A(n3313), .Z(n3311) );
  XOR U5205 ( .A(n3632), .B(n3633), .Z(n3313) );
  AND U5206 ( .A(n3634), .B(n3635), .Z(n3633) );
  XNOR U5207 ( .A(n3632), .B(n3636), .Z(n3634) );
  XNOR U5208 ( .A(n3323), .B(n3315), .Z(n3614) );
  XOR U5209 ( .A(n3648), .B(n3328), .Z(n3323) );
  XOR U5210 ( .A(n3649), .B(n3319), .Z(n3320) );
  AND U5211 ( .A(n3652), .B(n3653), .Z(n3651) );
  XNOR U5212 ( .A(n3650), .B(n3654), .Z(n3652) );
  XNOR U5213 ( .A(n3327), .B(n3322), .Z(n3648) );
  XOR U5214 ( .A(n3665), .B(n3332), .Z(n3327) );
  XNOR U5215 ( .A(n3330), .B(n3326), .Z(n3665) );
  XOR U5216 ( .A(n3672), .B(n3329), .Z(n3330) );
  IV U5217 ( .A(n3331), .Z(n3329) );
  XOR U5218 ( .A(n3680), .B(n3343), .Z(n3338) );
  XOR U5219 ( .A(n3681), .B(n3334), .Z(n3335) );
  AND U5220 ( .A(n3684), .B(n3685), .Z(n3683) );
  XNOR U5221 ( .A(n3682), .B(n3686), .Z(n3684) );
  XNOR U5222 ( .A(n3342), .B(n3337), .Z(n3680) );
  XOR U5223 ( .A(n3698), .B(n3347), .Z(n3342) );
  XNOR U5224 ( .A(n3345), .B(n3341), .Z(n3698) );
  XOR U5225 ( .A(n3705), .B(n3344), .Z(n3345) );
  IV U5226 ( .A(n3346), .Z(n3344) );
  XOR U5227 ( .A(n3713), .B(n3357), .Z(n3350) );
  XNOR U5228 ( .A(n3354), .B(n3349), .Z(n3713) );
  XOR U5229 ( .A(n3720), .B(n3352), .Z(n3354) );
  IV U5230 ( .A(n3356), .Z(n3352) );
  XOR U5231 ( .A(n3728), .B(n3358), .Z(n3359) );
  IV U5232 ( .A(n3360), .Z(n3358) );
  XOR U5233 ( .A(n3729), .B(n3730), .Z(n3360) );
  AND U5234 ( .A(n3731), .B(n3732), .Z(n3730) );
  XNOR U5235 ( .A(n3729), .B(n3733), .Z(n3731) );
  XOR U5236 ( .A(n3742), .B(n3453), .Z(n1118) );
  XOR U5237 ( .A(n3743), .B(n3385), .Z(n3377) );
  XOR U5238 ( .A(n3744), .B(n3371), .Z(n3366) );
  XNOR U5239 ( .A(n3369), .B(n3365), .Z(n3744) );
  XOR U5240 ( .A(n3749), .B(n3750), .Z(n3365) );
  AND U5241 ( .A(n3751), .B(n3752), .Z(n3750) );
  XNOR U5242 ( .A(n3749), .B(n3753), .Z(n3751) );
  XOR U5243 ( .A(n3754), .B(n3368), .Z(n3369) );
  IV U5244 ( .A(n3370), .Z(n3368) );
  XOR U5245 ( .A(n3762), .B(n3372), .Z(n3373) );
  IV U5246 ( .A(n3374), .Z(n3372) );
  XNOR U5247 ( .A(n3384), .B(n3376), .Z(n3743) );
  XOR U5248 ( .A(n3777), .B(n3389), .Z(n3384) );
  XOR U5249 ( .A(n3778), .B(n3380), .Z(n3381) );
  AND U5250 ( .A(n3781), .B(n3782), .Z(n3780) );
  XNOR U5251 ( .A(n3779), .B(n3783), .Z(n3781) );
  XNOR U5252 ( .A(n3388), .B(n3383), .Z(n3777) );
  XOR U5253 ( .A(n3794), .B(n3393), .Z(n3388) );
  XNOR U5254 ( .A(n3391), .B(n3387), .Z(n3794) );
  XOR U5255 ( .A(n3801), .B(n3390), .Z(n3391) );
  IV U5256 ( .A(n3392), .Z(n3390) );
  XOR U5257 ( .A(n3809), .B(n3405), .Z(n3400) );
  XOR U5258 ( .A(n3810), .B(n3395), .Z(n3396) );
  IV U5259 ( .A(n3397), .Z(n3395) );
  XNOR U5260 ( .A(n3404), .B(n3399), .Z(n3809) );
  XOR U5261 ( .A(n3825), .B(n3409), .Z(n3404) );
  XNOR U5262 ( .A(n3407), .B(n3403), .Z(n3825) );
  XOR U5263 ( .A(n3832), .B(n3406), .Z(n3407) );
  IV U5264 ( .A(n3408), .Z(n3406) );
  XOR U5265 ( .A(n3840), .B(n3417), .Z(n3412) );
  XNOR U5266 ( .A(n3415), .B(n3411), .Z(n3840) );
  XOR U5267 ( .A(n3848), .B(n3414), .Z(n3415) );
  IV U5268 ( .A(n3416), .Z(n3414) );
  XOR U5269 ( .A(n3856), .B(n3418), .Z(n3419) );
  AND U5270 ( .A(n3859), .B(n3860), .Z(n3858) );
  XNOR U5271 ( .A(n3857), .B(n3861), .Z(n3859) );
  XNOR U5272 ( .A(n3452), .B(n3484), .Z(n3742) );
  XOR U5273 ( .A(n3870), .B(n3468), .Z(n3452) );
  XOR U5274 ( .A(n3871), .B(n3433), .Z(n3428) );
  XOR U5275 ( .A(n3872), .B(n3423), .Z(n3424) );
  IV U5276 ( .A(n3425), .Z(n3423) );
  XNOR U5277 ( .A(n3432), .B(n3427), .Z(n3871) );
  XOR U5278 ( .A(n3886), .B(n3437), .Z(n3432) );
  XNOR U5279 ( .A(n3435), .B(n3431), .Z(n3886) );
  XOR U5280 ( .A(n3893), .B(n3434), .Z(n3435) );
  IV U5281 ( .A(n3436), .Z(n3434) );
  XOR U5282 ( .A(n3901), .B(n3447), .Z(n3442) );
  XNOR U5283 ( .A(n3445), .B(n3439), .Z(n3901) );
  XOR U5284 ( .A(n3908), .B(n3444), .Z(n3445) );
  IV U5285 ( .A(n3446), .Z(n3444) );
  XOR U5286 ( .A(n3916), .B(n3448), .Z(n3449) );
  AND U5287 ( .A(n3919), .B(n3920), .Z(n3918) );
  XNOR U5288 ( .A(n3917), .B(n3921), .Z(n3919) );
  XNOR U5289 ( .A(n3467), .B(n3451), .Z(n3870) );
  XOR U5290 ( .A(n3933), .B(n3475), .Z(n3467) );
  XOR U5291 ( .A(n3934), .B(n3462), .Z(n3457) );
  XNOR U5292 ( .A(n3460), .B(n3456), .Z(n3934) );
  XOR U5293 ( .A(n3942), .B(n3459), .Z(n3460) );
  IV U5294 ( .A(n3461), .Z(n3459) );
  XOR U5295 ( .A(n3950), .B(n3463), .Z(n3464) );
  AND U5296 ( .A(n3953), .B(n3954), .Z(n3952) );
  XNOR U5297 ( .A(n3951), .B(n3955), .Z(n3953) );
  XNOR U5298 ( .A(n3474), .B(n3466), .Z(n3933) );
  XOR U5299 ( .A(n3966), .B(n3479), .Z(n3474) );
  XOR U5300 ( .A(n3967), .B(n3470), .Z(n3471) );
  AND U5301 ( .A(n3970), .B(n3971), .Z(n3969) );
  XNOR U5302 ( .A(n3968), .B(n3972), .Z(n3970) );
  XNOR U5303 ( .A(n3478), .B(n3473), .Z(n3966) );
  XOR U5304 ( .A(n3983), .B(n3483), .Z(n3478) );
  XNOR U5305 ( .A(n3481), .B(n3477), .Z(n3983) );
  XOR U5306 ( .A(n3990), .B(n3480), .Z(n3481) );
  IV U5307 ( .A(n3482), .Z(n3480) );
  XOR U5308 ( .A(n3999), .B(n3581), .Z(n3549) );
  XOR U5309 ( .A(n4000), .B(n3509), .Z(n3501) );
  XOR U5310 ( .A(n4001), .B(n3496), .Z(n3491) );
  XNOR U5311 ( .A(n3494), .B(n3488), .Z(n4001) );
  XOR U5312 ( .A(n4009), .B(n3493), .Z(n3494) );
  IV U5313 ( .A(n3495), .Z(n3493) );
  XOR U5314 ( .A(n4017), .B(n3497), .Z(n3498) );
  AND U5315 ( .A(n4020), .B(n4021), .Z(n4019) );
  XNOR U5316 ( .A(n4018), .B(n4022), .Z(n4020) );
  XNOR U5317 ( .A(n3508), .B(n3500), .Z(n4000) );
  XOR U5318 ( .A(n4034), .B(n3513), .Z(n3508) );
  XOR U5319 ( .A(n4035), .B(n3504), .Z(n3505) );
  AND U5320 ( .A(n4038), .B(n4039), .Z(n4037) );
  XNOR U5321 ( .A(n4036), .B(n4040), .Z(n4038) );
  XNOR U5322 ( .A(n3512), .B(n3507), .Z(n4034) );
  XOR U5323 ( .A(n4051), .B(n3517), .Z(n3512) );
  XNOR U5324 ( .A(n3515), .B(n3511), .Z(n4051) );
  XOR U5325 ( .A(n4058), .B(n3514), .Z(n3515) );
  IV U5326 ( .A(n3516), .Z(n3514) );
  XOR U5327 ( .A(n4066), .B(n3529), .Z(n3524) );
  XOR U5328 ( .A(n4067), .B(n3519), .Z(n3520) );
  IV U5329 ( .A(n3521), .Z(n3519) );
  XNOR U5330 ( .A(n3528), .B(n3523), .Z(n4066) );
  XOR U5331 ( .A(n4082), .B(n3533), .Z(n3528) );
  XNOR U5332 ( .A(n3531), .B(n3527), .Z(n4082) );
  XOR U5333 ( .A(n4089), .B(n3530), .Z(n3531) );
  IV U5334 ( .A(n3532), .Z(n3530) );
  XOR U5335 ( .A(n4097), .B(n3543), .Z(n3538) );
  XNOR U5336 ( .A(n3541), .B(n3535), .Z(n4097) );
  XOR U5337 ( .A(n4105), .B(n3540), .Z(n3541) );
  IV U5338 ( .A(n3542), .Z(n3540) );
  XOR U5339 ( .A(n4113), .B(n3544), .Z(n3545) );
  IV U5340 ( .A(n3546), .Z(n3544) );
  XNOR U5341 ( .A(n3580), .B(n3548), .Z(n3999) );
  XOR U5342 ( .A(n4128), .B(n3598), .Z(n3580) );
  XOR U5343 ( .A(n4129), .B(n3562), .Z(n3557) );
  XOR U5344 ( .A(n4130), .B(n3553), .Z(n3554) );
  AND U5345 ( .A(n4133), .B(n4134), .Z(n4132) );
  XNOR U5346 ( .A(n4131), .B(n4135), .Z(n4133) );
  XNOR U5347 ( .A(n3561), .B(n3556), .Z(n4129) );
  XOR U5348 ( .A(n4146), .B(n3566), .Z(n3561) );
  XNOR U5349 ( .A(n3564), .B(n3560), .Z(n4146) );
  XOR U5350 ( .A(n4153), .B(n3563), .Z(n3564) );
  IV U5351 ( .A(n3565), .Z(n3563) );
  XOR U5352 ( .A(n4161), .B(n3574), .Z(n3569) );
  XNOR U5353 ( .A(n3572), .B(n3568), .Z(n4161) );
  XOR U5354 ( .A(n4169), .B(n3571), .Z(n3572) );
  IV U5355 ( .A(n3573), .Z(n3571) );
  XOR U5356 ( .A(n4177), .B(n3575), .Z(n3576) );
  IV U5357 ( .A(n3577), .Z(n3575) );
  XNOR U5358 ( .A(n3597), .B(n3579), .Z(n4128) );
  XOR U5359 ( .A(n4192), .B(n3605), .Z(n3597) );
  XOR U5360 ( .A(n4193), .B(n3592), .Z(n3587) );
  XNOR U5361 ( .A(n3590), .B(n3584), .Z(n4193) );
  XOR U5362 ( .A(n4201), .B(n3589), .Z(n3590) );
  IV U5363 ( .A(n3591), .Z(n3589) );
  XOR U5364 ( .A(n4209), .B(n3593), .Z(n3594) );
  AND U5365 ( .A(n4212), .B(n4213), .Z(n4211) );
  XNOR U5366 ( .A(n4210), .B(n4214), .Z(n4212) );
  XNOR U5367 ( .A(n3604), .B(n3596), .Z(n4192) );
  XOR U5368 ( .A(n4226), .B(n3609), .Z(n3604) );
  XOR U5369 ( .A(n4227), .B(n3600), .Z(n3601) );
  AND U5370 ( .A(n4230), .B(n4231), .Z(n4229) );
  XNOR U5371 ( .A(n4228), .B(n4232), .Z(n4230) );
  XNOR U5372 ( .A(n3608), .B(n3603), .Z(n4226) );
  XOR U5373 ( .A(n4244), .B(n3613), .Z(n3608) );
  XNOR U5374 ( .A(n3611), .B(n3607), .Z(n4244) );
  XOR U5375 ( .A(n4251), .B(n3610), .Z(n3611) );
  IV U5376 ( .A(n3612), .Z(n3610) );
  XOR U5377 ( .A(n4259), .B(n3664), .Z(n3646) );
  XOR U5378 ( .A(n4260), .B(n3626), .Z(n3621) );
  XOR U5379 ( .A(n4261), .B(n3616), .Z(n3617) );
  IV U5380 ( .A(n3618), .Z(n3616) );
  XNOR U5381 ( .A(n3625), .B(n3620), .Z(n4260) );
  XOR U5382 ( .A(n4276), .B(n3630), .Z(n3625) );
  XNOR U5383 ( .A(n3628), .B(n3624), .Z(n4276) );
  XOR U5384 ( .A(n4283), .B(n3627), .Z(n3628) );
  IV U5385 ( .A(n3629), .Z(n3627) );
  XOR U5386 ( .A(n4291), .B(n3640), .Z(n3635) );
  XNOR U5387 ( .A(n3638), .B(n3632), .Z(n4291) );
  XOR U5388 ( .A(n4299), .B(n3637), .Z(n3638) );
  IV U5389 ( .A(n3639), .Z(n3637) );
  XOR U5390 ( .A(n4307), .B(n3641), .Z(n3642) );
  IV U5391 ( .A(n3643), .Z(n3641) );
  XOR U5392 ( .A(n4308), .B(n4309), .Z(n3643) );
  AND U5393 ( .A(n4310), .B(n4311), .Z(n4309) );
  XNOR U5394 ( .A(n4308), .B(n4312), .Z(n4310) );
  XNOR U5395 ( .A(n3663), .B(n3645), .Z(n4259) );
  XOR U5396 ( .A(n4321), .B(n4322), .Z(n3645) );
  AND U5397 ( .A(n4323), .B(n4324), .Z(n4322) );
  XNOR U5398 ( .A(n4321), .B(n4325), .Z(n4323) );
  XOR U5399 ( .A(n4326), .B(n3671), .Z(n3663) );
  XOR U5400 ( .A(n4327), .B(n3658), .Z(n3653) );
  XNOR U5401 ( .A(n3656), .B(n3650), .Z(n4327) );
  XOR U5402 ( .A(n4335), .B(n3655), .Z(n3656) );
  IV U5403 ( .A(n3657), .Z(n3655) );
  XOR U5404 ( .A(n4343), .B(n3659), .Z(n3660) );
  AND U5405 ( .A(n4346), .B(n4347), .Z(n4345) );
  XNOR U5406 ( .A(n4344), .B(n4348), .Z(n4346) );
  XNOR U5407 ( .A(n3670), .B(n3662), .Z(n4326) );
  XOR U5408 ( .A(n4359), .B(n3675), .Z(n3670) );
  XOR U5409 ( .A(n4360), .B(n3666), .Z(n3667) );
  AND U5410 ( .A(n4363), .B(n4364), .Z(n4362) );
  XNOR U5411 ( .A(n4361), .B(n4365), .Z(n4363) );
  XNOR U5412 ( .A(n3674), .B(n3669), .Z(n4359) );
  XOR U5413 ( .A(n4376), .B(n3679), .Z(n3674) );
  XNOR U5414 ( .A(n3677), .B(n3673), .Z(n4376) );
  XOR U5415 ( .A(n4383), .B(n3676), .Z(n3677) );
  IV U5416 ( .A(n3678), .Z(n3676) );
  XOR U5417 ( .A(n4391), .B(n3704), .Z(n3696) );
  XOR U5418 ( .A(n4392), .B(n3690), .Z(n3685) );
  XNOR U5419 ( .A(n3688), .B(n3682), .Z(n4392) );
  XOR U5420 ( .A(n4400), .B(n3687), .Z(n3688) );
  IV U5421 ( .A(n3689), .Z(n3687) );
  XOR U5422 ( .A(n4408), .B(n3691), .Z(n3692) );
  IV U5423 ( .A(n3693), .Z(n3691) );
  XNOR U5424 ( .A(n3703), .B(n3695), .Z(n4391) );
  XOR U5425 ( .A(n4423), .B(n3708), .Z(n3703) );
  XOR U5426 ( .A(n4424), .B(n3699), .Z(n3700) );
  AND U5427 ( .A(n4427), .B(n4428), .Z(n4426) );
  XNOR U5428 ( .A(n4425), .B(n4429), .Z(n4427) );
  XNOR U5429 ( .A(n3707), .B(n3702), .Z(n4423) );
  XOR U5430 ( .A(n4440), .B(n3712), .Z(n3707) );
  XNOR U5431 ( .A(n3710), .B(n3706), .Z(n4440) );
  XOR U5432 ( .A(n4447), .B(n3709), .Z(n3710) );
  IV U5433 ( .A(n3711), .Z(n3709) );
  XOR U5434 ( .A(n4455), .B(n3723), .Z(n3718) );
  XOR U5435 ( .A(n4456), .B(n3714), .Z(n3715) );
  AND U5436 ( .A(n4459), .B(n4460), .Z(n4458) );
  XNOR U5437 ( .A(n4457), .B(n4461), .Z(n4459) );
  XNOR U5438 ( .A(n3722), .B(n3717), .Z(n4455) );
  XOR U5439 ( .A(n4472), .B(n3727), .Z(n3722) );
  XNOR U5440 ( .A(n3725), .B(n3721), .Z(n4472) );
  XOR U5441 ( .A(n4479), .B(n3724), .Z(n3725) );
  IV U5442 ( .A(n3726), .Z(n3724) );
  XOR U5443 ( .A(n4487), .B(n3737), .Z(n3732) );
  XNOR U5444 ( .A(n3735), .B(n3729), .Z(n4487) );
  XOR U5445 ( .A(n4495), .B(n3734), .Z(n3735) );
  IV U5446 ( .A(n3736), .Z(n3734) );
  XOR U5447 ( .A(n4503), .B(n3738), .Z(n3739) );
  IV U5448 ( .A(n3740), .Z(n3738) );
  XOR U5449 ( .A(n4504), .B(n4505), .Z(n3740) );
  AND U5450 ( .A(n4506), .B(n4507), .Z(n4505) );
  XNOR U5451 ( .A(n4504), .B(n4508), .Z(n4506) );
  XOR U5452 ( .A(n4509), .B(n4510), .Z(n4503) );
  AND U5453 ( .A(n4511), .B(n4512), .Z(n4510) );
  XNOR U5454 ( .A(n4513), .B(n4514), .Z(n4512) );
  XOR U5455 ( .A(n4519), .B(n3932), .Z(n1405) );
  XOR U5456 ( .A(n4520), .B(n3793), .Z(n3775) );
  XOR U5457 ( .A(n4521), .B(n3757), .Z(n3752) );
  XOR U5458 ( .A(n4522), .B(n3745), .Z(n3746) );
  IV U5459 ( .A(n3747), .Z(n3745) );
  XNOR U5460 ( .A(n3756), .B(n3749), .Z(n4521) );
  XOR U5461 ( .A(n4537), .B(n3761), .Z(n3756) );
  XNOR U5462 ( .A(n3759), .B(n3755), .Z(n4537) );
  XOR U5463 ( .A(n4544), .B(n3758), .Z(n3759) );
  IV U5464 ( .A(n3760), .Z(n3758) );
  XOR U5465 ( .A(n4552), .B(n3769), .Z(n3764) );
  XNOR U5466 ( .A(n3767), .B(n3763), .Z(n4552) );
  XOR U5467 ( .A(n4560), .B(n3766), .Z(n3767) );
  IV U5468 ( .A(n3768), .Z(n3766) );
  XOR U5469 ( .A(n4568), .B(n3770), .Z(n3771) );
  IV U5470 ( .A(n3772), .Z(n3770) );
  XOR U5471 ( .A(n4572), .B(n4573), .Z(n4568) );
  AND U5472 ( .A(n4574), .B(n4575), .Z(n4573) );
  XNOR U5473 ( .A(n4576), .B(n4577), .Z(n4575) );
  XNOR U5474 ( .A(n3792), .B(n3774), .Z(n4520) );
  XOR U5475 ( .A(n4585), .B(n3800), .Z(n3792) );
  XOR U5476 ( .A(n4586), .B(n3787), .Z(n3782) );
  XNOR U5477 ( .A(n3785), .B(n3779), .Z(n4586) );
  XOR U5478 ( .A(n4594), .B(n3784), .Z(n3785) );
  IV U5479 ( .A(n3786), .Z(n3784) );
  XOR U5480 ( .A(n4602), .B(n3788), .Z(n3789) );
  AND U5481 ( .A(n4605), .B(n4606), .Z(n4604) );
  XNOR U5482 ( .A(n4603), .B(n4607), .Z(n4605) );
  XNOR U5483 ( .A(n3799), .B(n3791), .Z(n4585) );
  XOR U5484 ( .A(n4618), .B(n3804), .Z(n3799) );
  XOR U5485 ( .A(n4619), .B(n3795), .Z(n3796) );
  AND U5486 ( .A(n4622), .B(n4623), .Z(n4621) );
  XNOR U5487 ( .A(n4620), .B(n4624), .Z(n4622) );
  XNOR U5488 ( .A(n3803), .B(n3798), .Z(n4618) );
  XOR U5489 ( .A(n4635), .B(n3808), .Z(n3803) );
  XNOR U5490 ( .A(n3806), .B(n3802), .Z(n4635) );
  XOR U5491 ( .A(n4642), .B(n3805), .Z(n3806) );
  IV U5492 ( .A(n3807), .Z(n3805) );
  XOR U5493 ( .A(n4650), .B(n3831), .Z(n3823) );
  XOR U5494 ( .A(n4651), .B(n3817), .Z(n3812) );
  XNOR U5495 ( .A(n3815), .B(n3811), .Z(n4651) );
  XOR U5496 ( .A(n4658), .B(n3814), .Z(n3815) );
  IV U5497 ( .A(n3816), .Z(n3814) );
  XOR U5498 ( .A(n4666), .B(n3818), .Z(n3819) );
  IV U5499 ( .A(n3820), .Z(n3818) );
  XNOR U5500 ( .A(n3830), .B(n3822), .Z(n4650) );
  XOR U5501 ( .A(n4681), .B(n3835), .Z(n3830) );
  XOR U5502 ( .A(n4682), .B(n3826), .Z(n3827) );
  AND U5503 ( .A(n4685), .B(n4686), .Z(n4684) );
  XNOR U5504 ( .A(n4683), .B(n4687), .Z(n4685) );
  XNOR U5505 ( .A(n3834), .B(n3829), .Z(n4681) );
  XOR U5506 ( .A(n4699), .B(n3839), .Z(n3834) );
  XNOR U5507 ( .A(n3837), .B(n3833), .Z(n4699) );
  XOR U5508 ( .A(n4707), .B(n3836), .Z(n3837) );
  IV U5509 ( .A(n3838), .Z(n3836) );
  XOR U5510 ( .A(n4715), .B(n3851), .Z(n3846) );
  XOR U5511 ( .A(n4716), .B(n3841), .Z(n3842) );
  IV U5512 ( .A(n3843), .Z(n3841) );
  XNOR U5513 ( .A(n3850), .B(n3845), .Z(n4715) );
  XOR U5514 ( .A(n4731), .B(n3855), .Z(n3850) );
  XNOR U5515 ( .A(n3853), .B(n3849), .Z(n4731) );
  XOR U5516 ( .A(n4739), .B(n3852), .Z(n3853) );
  IV U5517 ( .A(n3854), .Z(n3852) );
  XOR U5518 ( .A(n4747), .B(n3865), .Z(n3860) );
  XNOR U5519 ( .A(n3863), .B(n3857), .Z(n4747) );
  XOR U5520 ( .A(n4755), .B(n3862), .Z(n3863) );
  IV U5521 ( .A(n3864), .Z(n3862) );
  XOR U5522 ( .A(n4763), .B(n3866), .Z(n3867) );
  IV U5523 ( .A(n3868), .Z(n3866) );
  XOR U5524 ( .A(n4764), .B(n4765), .Z(n3868) );
  AND U5525 ( .A(n4766), .B(n4767), .Z(n4765) );
  XNOR U5526 ( .A(n4764), .B(n4768), .Z(n4766) );
  XNOR U5527 ( .A(n3931), .B(n3998), .Z(n4519) );
  XOR U5528 ( .A(n4777), .B(n3965), .Z(n3931) );
  XOR U5529 ( .A(n4778), .B(n3892), .Z(n3884) );
  XOR U5530 ( .A(n4779), .B(n3879), .Z(n3874) );
  XNOR U5531 ( .A(n3877), .B(n3873), .Z(n4779) );
  XOR U5532 ( .A(n4786), .B(n3876), .Z(n3877) );
  IV U5533 ( .A(n3878), .Z(n3876) );
  XOR U5534 ( .A(n4794), .B(n3880), .Z(n3881) );
  AND U5535 ( .A(n4797), .B(n4798), .Z(n4796) );
  XNOR U5536 ( .A(n4795), .B(n4799), .Z(n4797) );
  XNOR U5537 ( .A(n3891), .B(n3883), .Z(n4778) );
  XOR U5538 ( .A(n4810), .B(n3896), .Z(n3891) );
  XOR U5539 ( .A(n4811), .B(n3887), .Z(n3888) );
  AND U5540 ( .A(n4814), .B(n4815), .Z(n4813) );
  XNOR U5541 ( .A(n4812), .B(n4816), .Z(n4814) );
  XNOR U5542 ( .A(n3895), .B(n3890), .Z(n4810) );
  XOR U5543 ( .A(n4827), .B(n3900), .Z(n3895) );
  XNOR U5544 ( .A(n3898), .B(n3894), .Z(n4827) );
  XOR U5545 ( .A(n4834), .B(n3897), .Z(n3898) );
  IV U5546 ( .A(n3899), .Z(n3897) );
  XOR U5547 ( .A(n4842), .B(n3911), .Z(n3906) );
  XOR U5548 ( .A(n4843), .B(n3902), .Z(n3903) );
  AND U5549 ( .A(n4846), .B(n4847), .Z(n4845) );
  XNOR U5550 ( .A(n4844), .B(n4848), .Z(n4846) );
  XNOR U5551 ( .A(n3910), .B(n3905), .Z(n4842) );
  XOR U5552 ( .A(n4859), .B(n3915), .Z(n3910) );
  XNOR U5553 ( .A(n3913), .B(n3909), .Z(n4859) );
  XOR U5554 ( .A(n4867), .B(n3912), .Z(n3913) );
  IV U5555 ( .A(n3914), .Z(n3912) );
  XOR U5556 ( .A(n4875), .B(n3925), .Z(n3920) );
  XNOR U5557 ( .A(n3923), .B(n3917), .Z(n4875) );
  XOR U5558 ( .A(n4880), .B(n4881), .Z(n3917) );
  AND U5559 ( .A(n4882), .B(n4883), .Z(n4881) );
  XNOR U5560 ( .A(n4880), .B(n4884), .Z(n4882) );
  XOR U5561 ( .A(n4885), .B(n3922), .Z(n3923) );
  IV U5562 ( .A(n3924), .Z(n3922) );
  XOR U5563 ( .A(n4893), .B(n3926), .Z(n3927) );
  IV U5564 ( .A(n3928), .Z(n3926) );
  XNOR U5565 ( .A(n3964), .B(n3930), .Z(n4777) );
  XOR U5566 ( .A(n4907), .B(n3982), .Z(n3964) );
  XOR U5567 ( .A(n4908), .B(n3945), .Z(n3940) );
  XOR U5568 ( .A(n4909), .B(n3935), .Z(n3936) );
  IV U5569 ( .A(n3937), .Z(n3935) );
  XNOR U5570 ( .A(n3944), .B(n3939), .Z(n4908) );
  XOR U5571 ( .A(n4924), .B(n3949), .Z(n3944) );
  XNOR U5572 ( .A(n3947), .B(n3943), .Z(n4924) );
  XOR U5573 ( .A(n4931), .B(n3946), .Z(n3947) );
  IV U5574 ( .A(n3948), .Z(n3946) );
  XOR U5575 ( .A(n4939), .B(n3959), .Z(n3954) );
  XNOR U5576 ( .A(n3957), .B(n3951), .Z(n4939) );
  XOR U5577 ( .A(n4944), .B(n4945), .Z(n3951) );
  AND U5578 ( .A(n4946), .B(n4947), .Z(n4945) );
  XNOR U5579 ( .A(n4944), .B(n4948), .Z(n4946) );
  XOR U5580 ( .A(n4949), .B(n3956), .Z(n3957) );
  IV U5581 ( .A(n3958), .Z(n3956) );
  XOR U5582 ( .A(n4956), .B(n3960), .Z(n3961) );
  AND U5583 ( .A(n4959), .B(n4960), .Z(n4958) );
  XNOR U5584 ( .A(n4957), .B(n4961), .Z(n4959) );
  XNOR U5585 ( .A(n3981), .B(n3963), .Z(n4907) );
  XOR U5586 ( .A(n4973), .B(n3989), .Z(n3981) );
  XOR U5587 ( .A(n4974), .B(n3976), .Z(n3971) );
  XNOR U5588 ( .A(n3974), .B(n3968), .Z(n4974) );
  XOR U5589 ( .A(n4982), .B(n3973), .Z(n3974) );
  IV U5590 ( .A(n3975), .Z(n3973) );
  XOR U5591 ( .A(n4990), .B(n3977), .Z(n3978) );
  AND U5592 ( .A(n4993), .B(n4994), .Z(n4992) );
  XNOR U5593 ( .A(n4991), .B(n4995), .Z(n4993) );
  XNOR U5594 ( .A(n3988), .B(n3980), .Z(n4973) );
  XOR U5595 ( .A(n5007), .B(n3993), .Z(n3988) );
  XOR U5596 ( .A(n5008), .B(n3984), .Z(n3985) );
  AND U5597 ( .A(n5011), .B(n5012), .Z(n5010) );
  XNOR U5598 ( .A(n5009), .B(n5013), .Z(n5011) );
  XNOR U5599 ( .A(n3992), .B(n3987), .Z(n5007) );
  XOR U5600 ( .A(n5023), .B(n3997), .Z(n3992) );
  XNOR U5601 ( .A(n3995), .B(n3991), .Z(n5023) );
  XOR U5602 ( .A(n5030), .B(n3994), .Z(n3995) );
  IV U5603 ( .A(n3996), .Z(n3994) );
  XOR U5604 ( .A(n5039), .B(n4191), .Z(n4126) );
  XOR U5605 ( .A(n5040), .B(n4050), .Z(n4032) );
  XOR U5606 ( .A(n5041), .B(n4012), .Z(n4007) );
  XOR U5607 ( .A(n5042), .B(n4002), .Z(n4003) );
  IV U5608 ( .A(n4004), .Z(n4002) );
  XNOR U5609 ( .A(n4011), .B(n4006), .Z(n5041) );
  XOR U5610 ( .A(n5055), .B(n4016), .Z(n4011) );
  XNOR U5611 ( .A(n4014), .B(n4010), .Z(n5055) );
  XOR U5612 ( .A(n5062), .B(n4013), .Z(n4014) );
  IV U5613 ( .A(n4015), .Z(n4013) );
  XOR U5614 ( .A(n5069), .B(n4026), .Z(n4021) );
  XNOR U5615 ( .A(n4024), .B(n4018), .Z(n5069) );
  XOR U5616 ( .A(n5076), .B(n4023), .Z(n4024) );
  IV U5617 ( .A(n4025), .Z(n4023) );
  XOR U5618 ( .A(n5083), .B(n4027), .Z(n4028) );
  IV U5619 ( .A(n4029), .Z(n4027) );
  XNOR U5620 ( .A(n4049), .B(n4031), .Z(n5040) );
  XOR U5621 ( .A(n5096), .B(n4057), .Z(n4049) );
  XOR U5622 ( .A(n5097), .B(n4044), .Z(n4039) );
  XNOR U5623 ( .A(n4042), .B(n4036), .Z(n5097) );
  XOR U5624 ( .A(n5104), .B(n4041), .Z(n4042) );
  IV U5625 ( .A(n4043), .Z(n4041) );
  XOR U5626 ( .A(n5111), .B(n4045), .Z(n4046) );
  ANDN U5627 ( .B(n5114), .A(n5115), .Z(n5113) );
  XOR U5628 ( .A(n5112), .B(n5116), .Z(n5114) );
  XNOR U5629 ( .A(n4056), .B(n4048), .Z(n5096) );
  XOR U5630 ( .A(n5126), .B(n4061), .Z(n4056) );
  XOR U5631 ( .A(n5127), .B(n4052), .Z(n4053) );
  ANDN U5632 ( .B(n5130), .A(n5131), .Z(n5129) );
  XOR U5633 ( .A(n5128), .B(n5132), .Z(n5130) );
  XNOR U5634 ( .A(n4060), .B(n4055), .Z(n5126) );
  XOR U5635 ( .A(n5142), .B(n4065), .Z(n4060) );
  XNOR U5636 ( .A(n4063), .B(n4059), .Z(n5142) );
  XOR U5637 ( .A(n5149), .B(n4062), .Z(n4063) );
  IV U5638 ( .A(n4064), .Z(n4062) );
  XOR U5639 ( .A(n5156), .B(n4088), .Z(n4080) );
  XOR U5640 ( .A(n5157), .B(n4074), .Z(n4069) );
  XNOR U5641 ( .A(n4072), .B(n4068), .Z(n5157) );
  XOR U5642 ( .A(n5164), .B(n4071), .Z(n4072) );
  IV U5643 ( .A(n4073), .Z(n4071) );
  XOR U5644 ( .A(n5171), .B(n4075), .Z(n4076) );
  IV U5645 ( .A(n4077), .Z(n4075) );
  XNOR U5646 ( .A(n4087), .B(n4079), .Z(n5156) );
  XOR U5647 ( .A(n5184), .B(n4092), .Z(n4087) );
  XOR U5648 ( .A(n5185), .B(n4083), .Z(n4084) );
  ANDN U5649 ( .B(n5188), .A(n5189), .Z(n5187) );
  XOR U5650 ( .A(n5186), .B(n5190), .Z(n5188) );
  XNOR U5651 ( .A(n4091), .B(n4086), .Z(n5184) );
  XOR U5652 ( .A(n5200), .B(n4096), .Z(n4091) );
  XNOR U5653 ( .A(n4094), .B(n4090), .Z(n5200) );
  XOR U5654 ( .A(n5207), .B(n4093), .Z(n4094) );
  IV U5655 ( .A(n4095), .Z(n4093) );
  XOR U5656 ( .A(n5214), .B(n4108), .Z(n4103) );
  XOR U5657 ( .A(n5215), .B(n4098), .Z(n4099) );
  IV U5658 ( .A(n4100), .Z(n4098) );
  XNOR U5659 ( .A(n4107), .B(n4102), .Z(n5214) );
  XOR U5660 ( .A(n5228), .B(n4112), .Z(n4107) );
  XNOR U5661 ( .A(n4110), .B(n4106), .Z(n5228) );
  XOR U5662 ( .A(n5235), .B(n4109), .Z(n4110) );
  IV U5663 ( .A(n4111), .Z(n4109) );
  XOR U5664 ( .A(n5242), .B(n4120), .Z(n4115) );
  XNOR U5665 ( .A(n4118), .B(n4114), .Z(n5242) );
  XOR U5666 ( .A(n5249), .B(n4117), .Z(n4118) );
  IV U5667 ( .A(n4119), .Z(n4117) );
  XOR U5668 ( .A(n5256), .B(n4121), .Z(n4122) );
  IV U5669 ( .A(n4123), .Z(n4121) );
  XNOR U5670 ( .A(n4190), .B(n4125), .Z(n5039) );
  XOR U5671 ( .A(n5269), .B(n4225), .Z(n4190) );
  XOR U5672 ( .A(n5270), .B(n4152), .Z(n4144) );
  XOR U5673 ( .A(n5271), .B(n4139), .Z(n4134) );
  XNOR U5674 ( .A(n4137), .B(n4131), .Z(n5271) );
  XOR U5675 ( .A(n5278), .B(n4136), .Z(n4137) );
  IV U5676 ( .A(n4138), .Z(n4136) );
  XOR U5677 ( .A(n5285), .B(n4140), .Z(n4141) );
  ANDN U5678 ( .B(n5288), .A(n5289), .Z(n5287) );
  XOR U5679 ( .A(n5286), .B(n5290), .Z(n5288) );
  XNOR U5680 ( .A(n4151), .B(n4143), .Z(n5270) );
  XOR U5681 ( .A(n5300), .B(n4156), .Z(n4151) );
  XOR U5682 ( .A(n5301), .B(n4147), .Z(n4148) );
  ANDN U5683 ( .B(n5304), .A(n5305), .Z(n5303) );
  XOR U5684 ( .A(n5302), .B(n5306), .Z(n5304) );
  XNOR U5685 ( .A(n4155), .B(n4150), .Z(n5300) );
  XOR U5686 ( .A(n5316), .B(n4160), .Z(n4155) );
  XNOR U5687 ( .A(n4158), .B(n4154), .Z(n5316) );
  XOR U5688 ( .A(n5323), .B(n4157), .Z(n4158) );
  IV U5689 ( .A(n4159), .Z(n4157) );
  XOR U5690 ( .A(n5330), .B(n4172), .Z(n4167) );
  XOR U5691 ( .A(n5331), .B(n4162), .Z(n4163) );
  IV U5692 ( .A(n4164), .Z(n4162) );
  XNOR U5693 ( .A(n4171), .B(n4166), .Z(n5330) );
  XOR U5694 ( .A(n5344), .B(n4176), .Z(n4171) );
  XNOR U5695 ( .A(n4174), .B(n4170), .Z(n5344) );
  XOR U5696 ( .A(n5351), .B(n4173), .Z(n4174) );
  IV U5697 ( .A(n4175), .Z(n4173) );
  XOR U5698 ( .A(n5358), .B(n4184), .Z(n4179) );
  XNOR U5699 ( .A(n4182), .B(n4178), .Z(n5358) );
  XOR U5700 ( .A(n5365), .B(n4181), .Z(n4182) );
  IV U5701 ( .A(n4183), .Z(n4181) );
  XOR U5702 ( .A(n5372), .B(n4185), .Z(n4186) );
  IV U5703 ( .A(n4187), .Z(n4185) );
  XNOR U5704 ( .A(n4224), .B(n4189), .Z(n5269) );
  XOR U5705 ( .A(n5385), .B(n4243), .Z(n4224) );
  XOR U5706 ( .A(n5386), .B(n4204), .Z(n4199) );
  XOR U5707 ( .A(n5387), .B(n4194), .Z(n4195) );
  IV U5708 ( .A(n4196), .Z(n4194) );
  XNOR U5709 ( .A(n4203), .B(n4198), .Z(n5386) );
  XOR U5710 ( .A(n5400), .B(n4208), .Z(n4203) );
  XNOR U5711 ( .A(n4206), .B(n4202), .Z(n5400) );
  XOR U5712 ( .A(n5407), .B(n4205), .Z(n4206) );
  IV U5713 ( .A(n4207), .Z(n4205) );
  XOR U5714 ( .A(n5414), .B(n4218), .Z(n4213) );
  XNOR U5715 ( .A(n4216), .B(n4210), .Z(n5414) );
  XOR U5716 ( .A(n5421), .B(n4215), .Z(n4216) );
  IV U5717 ( .A(n4217), .Z(n4215) );
  XOR U5718 ( .A(n5428), .B(n4219), .Z(n4220) );
  IV U5719 ( .A(n4221), .Z(n4219) );
  XNOR U5720 ( .A(n4242), .B(n4223), .Z(n5385) );
  XOR U5721 ( .A(n5441), .B(n4250), .Z(n4242) );
  XOR U5722 ( .A(n5442), .B(n4236), .Z(n4231) );
  XNOR U5723 ( .A(n4234), .B(n4228), .Z(n5442) );
  XOR U5724 ( .A(n5449), .B(n4233), .Z(n4234) );
  IV U5725 ( .A(n4235), .Z(n4233) );
  XOR U5726 ( .A(n5456), .B(n4237), .Z(n4238) );
  IV U5727 ( .A(n4239), .Z(n4237) );
  XNOR U5728 ( .A(n4249), .B(n4241), .Z(n5441) );
  XOR U5729 ( .A(n5469), .B(n4254), .Z(n4249) );
  XOR U5730 ( .A(n5470), .B(n4245), .Z(n4246) );
  ANDN U5731 ( .B(n5473), .A(n5474), .Z(n5472) );
  XOR U5732 ( .A(n5471), .B(n5475), .Z(n5473) );
  XNOR U5733 ( .A(n4253), .B(n4248), .Z(n5469) );
  XOR U5734 ( .A(n5485), .B(n4258), .Z(n4253) );
  XNOR U5735 ( .A(n4256), .B(n4252), .Z(n5485) );
  XOR U5736 ( .A(n5492), .B(n4255), .Z(n4256) );
  IV U5737 ( .A(n4257), .Z(n4255) );
  XOR U5738 ( .A(n5499), .B(n4358), .Z(n4324) );
  XOR U5739 ( .A(n5500), .B(n4282), .Z(n4274) );
  XOR U5740 ( .A(n5501), .B(n4268), .Z(n4263) );
  XNOR U5741 ( .A(n4266), .B(n4262), .Z(n5501) );
  XOR U5742 ( .A(n5508), .B(n4265), .Z(n4266) );
  IV U5743 ( .A(n4267), .Z(n4265) );
  XOR U5744 ( .A(n5515), .B(n4269), .Z(n4270) );
  IV U5745 ( .A(n4271), .Z(n4269) );
  XNOR U5746 ( .A(n4281), .B(n4273), .Z(n5500) );
  XOR U5747 ( .A(n5528), .B(n4286), .Z(n4281) );
  XOR U5748 ( .A(n5529), .B(n4277), .Z(n4278) );
  ANDN U5749 ( .B(n5532), .A(n5533), .Z(n5531) );
  XOR U5750 ( .A(n5530), .B(n5534), .Z(n5532) );
  XNOR U5751 ( .A(n4285), .B(n4280), .Z(n5528) );
  XOR U5752 ( .A(n5544), .B(n4290), .Z(n4285) );
  XNOR U5753 ( .A(n4288), .B(n4284), .Z(n5544) );
  XOR U5754 ( .A(n5551), .B(n4287), .Z(n4288) );
  IV U5755 ( .A(n4289), .Z(n4287) );
  XOR U5756 ( .A(n5558), .B(n4302), .Z(n4297) );
  XOR U5757 ( .A(n5559), .B(n4292), .Z(n4293) );
  IV U5758 ( .A(n4294), .Z(n4292) );
  XNOR U5759 ( .A(n4301), .B(n4296), .Z(n5558) );
  XOR U5760 ( .A(n5572), .B(n4306), .Z(n4301) );
  XNOR U5761 ( .A(n4304), .B(n4300), .Z(n5572) );
  XOR U5762 ( .A(n5579), .B(n4303), .Z(n4304) );
  IV U5763 ( .A(n4305), .Z(n4303) );
  XOR U5764 ( .A(n5586), .B(n4316), .Z(n4311) );
  XNOR U5765 ( .A(n4314), .B(n4308), .Z(n5586) );
  XOR U5766 ( .A(n5593), .B(n4313), .Z(n4314) );
  IV U5767 ( .A(n4315), .Z(n4313) );
  XOR U5768 ( .A(n5600), .B(n4317), .Z(n4318) );
  IV U5769 ( .A(n4319), .Z(n4317) );
  XNOR U5770 ( .A(n4357), .B(n4321), .Z(n5499) );
  XOR U5771 ( .A(n5613), .B(n4375), .Z(n4357) );
  XOR U5772 ( .A(n5614), .B(n4338), .Z(n4333) );
  XOR U5773 ( .A(n5615), .B(n4328), .Z(n4329) );
  IV U5774 ( .A(n4330), .Z(n4328) );
  XNOR U5775 ( .A(n4337), .B(n4332), .Z(n5614) );
  XOR U5776 ( .A(n5628), .B(n4342), .Z(n4337) );
  XNOR U5777 ( .A(n4340), .B(n4336), .Z(n5628) );
  XOR U5778 ( .A(n5635), .B(n4339), .Z(n4340) );
  IV U5779 ( .A(n4341), .Z(n4339) );
  XOR U5780 ( .A(n5642), .B(n4352), .Z(n4347) );
  XNOR U5781 ( .A(n4350), .B(n4344), .Z(n5642) );
  XNOR U5782 ( .A(n5646), .B(n5647), .Z(n4344) );
  ANDN U5783 ( .B(n5648), .A(n5649), .Z(n5647) );
  XOR U5784 ( .A(n5646), .B(n5650), .Z(n5648) );
  XOR U5785 ( .A(n5651), .B(n4349), .Z(n4350) );
  IV U5786 ( .A(n4351), .Z(n4349) );
  XOR U5787 ( .A(n5658), .B(n4353), .Z(n4354) );
  ANDN U5788 ( .B(n5661), .A(n5662), .Z(n5660) );
  XOR U5789 ( .A(n5659), .B(n5663), .Z(n5661) );
  XNOR U5790 ( .A(n4374), .B(n4356), .Z(n5613) );
  XOR U5791 ( .A(n5673), .B(n4382), .Z(n4374) );
  XOR U5792 ( .A(n5674), .B(n4369), .Z(n4364) );
  XNOR U5793 ( .A(n4367), .B(n4361), .Z(n5674) );
  XOR U5794 ( .A(n5681), .B(n4366), .Z(n4367) );
  IV U5795 ( .A(n4368), .Z(n4366) );
  XOR U5796 ( .A(n5688), .B(n4370), .Z(n4371) );
  ANDN U5797 ( .B(n5691), .A(n5692), .Z(n5690) );
  XOR U5798 ( .A(n5689), .B(n5693), .Z(n5691) );
  XNOR U5799 ( .A(n4381), .B(n4373), .Z(n5673) );
  XOR U5800 ( .A(n5703), .B(n4386), .Z(n4381) );
  XOR U5801 ( .A(n5704), .B(n4377), .Z(n4378) );
  ANDN U5802 ( .B(n5707), .A(n5708), .Z(n5706) );
  XOR U5803 ( .A(n5705), .B(n5709), .Z(n5707) );
  XNOR U5804 ( .A(n4385), .B(n4380), .Z(n5703) );
  XOR U5805 ( .A(n5719), .B(n4390), .Z(n4385) );
  XNOR U5806 ( .A(n4388), .B(n4384), .Z(n5719) );
  XOR U5807 ( .A(n5726), .B(n4387), .Z(n4388) );
  IV U5808 ( .A(n4389), .Z(n4387) );
  XOR U5809 ( .A(n5733), .B(n4439), .Z(n4421) );
  XOR U5810 ( .A(n5734), .B(n4403), .Z(n4398) );
  XOR U5811 ( .A(n5735), .B(n4393), .Z(n4394) );
  IV U5812 ( .A(n4395), .Z(n4393) );
  XNOR U5813 ( .A(n4402), .B(n4397), .Z(n5734) );
  XOR U5814 ( .A(n5748), .B(n4407), .Z(n4402) );
  XNOR U5815 ( .A(n4405), .B(n4401), .Z(n5748) );
  XOR U5816 ( .A(n5755), .B(n4404), .Z(n4405) );
  IV U5817 ( .A(n4406), .Z(n4404) );
  XOR U5818 ( .A(n5762), .B(n4415), .Z(n4410) );
  XNOR U5819 ( .A(n4413), .B(n4409), .Z(n5762) );
  XOR U5820 ( .A(n5769), .B(n4412), .Z(n4413) );
  IV U5821 ( .A(n4414), .Z(n4412) );
  XOR U5822 ( .A(n5776), .B(n4416), .Z(n4417) );
  IV U5823 ( .A(n4418), .Z(n4416) );
  XNOR U5824 ( .A(n4438), .B(n4420), .Z(n5733) );
  XOR U5825 ( .A(n5789), .B(n4446), .Z(n4438) );
  XOR U5826 ( .A(n5790), .B(n4433), .Z(n4428) );
  XNOR U5827 ( .A(n4431), .B(n4425), .Z(n5790) );
  XOR U5828 ( .A(n5797), .B(n4430), .Z(n4431) );
  IV U5829 ( .A(n4432), .Z(n4430) );
  XOR U5830 ( .A(n5804), .B(n4434), .Z(n4435) );
  ANDN U5831 ( .B(n5807), .A(n5808), .Z(n5806) );
  XOR U5832 ( .A(n5805), .B(n5809), .Z(n5807) );
  XNOR U5833 ( .A(n4445), .B(n4437), .Z(n5789) );
  XOR U5834 ( .A(n5819), .B(n4450), .Z(n4445) );
  XOR U5835 ( .A(n5820), .B(n4441), .Z(n4442) );
  ANDN U5836 ( .B(n5823), .A(n5824), .Z(n5822) );
  XOR U5837 ( .A(n5821), .B(n5825), .Z(n5823) );
  XNOR U5838 ( .A(n4449), .B(n4444), .Z(n5819) );
  XOR U5839 ( .A(n5835), .B(n4454), .Z(n4449) );
  XNOR U5840 ( .A(n4452), .B(n4448), .Z(n5835) );
  XOR U5841 ( .A(n5842), .B(n4451), .Z(n4452) );
  IV U5842 ( .A(n4453), .Z(n4451) );
  XOR U5843 ( .A(n5849), .B(n4478), .Z(n4470) );
  XOR U5844 ( .A(n5850), .B(n4465), .Z(n4460) );
  XNOR U5845 ( .A(n4463), .B(n4457), .Z(n5850) );
  XOR U5846 ( .A(n5857), .B(n4462), .Z(n4463) );
  IV U5847 ( .A(n4464), .Z(n4462) );
  XOR U5848 ( .A(n5864), .B(n4466), .Z(n4467) );
  ANDN U5849 ( .B(n5867), .A(n5868), .Z(n5866) );
  XOR U5850 ( .A(n5865), .B(n5869), .Z(n5867) );
  XNOR U5851 ( .A(n4477), .B(n4469), .Z(n5849) );
  XOR U5852 ( .A(n5879), .B(n4482), .Z(n4477) );
  XOR U5853 ( .A(n5880), .B(n4473), .Z(n4474) );
  ANDN U5854 ( .B(n5883), .A(n5884), .Z(n5882) );
  XOR U5855 ( .A(n5881), .B(n5885), .Z(n5883) );
  XNOR U5856 ( .A(n4481), .B(n4476), .Z(n5879) );
  XOR U5857 ( .A(n5895), .B(n4486), .Z(n4481) );
  XNOR U5858 ( .A(n4484), .B(n4480), .Z(n5895) );
  XOR U5859 ( .A(n5902), .B(n4483), .Z(n4484) );
  IV U5860 ( .A(n4485), .Z(n4483) );
  XOR U5861 ( .A(n5909), .B(n4498), .Z(n4493) );
  XOR U5862 ( .A(n5910), .B(n4488), .Z(n4489) );
  IV U5863 ( .A(n4490), .Z(n4488) );
  XNOR U5864 ( .A(n4497), .B(n4492), .Z(n5909) );
  XOR U5865 ( .A(n5923), .B(n4502), .Z(n4497) );
  XNOR U5866 ( .A(n4500), .B(n4496), .Z(n5923) );
  XOR U5867 ( .A(n5930), .B(n4499), .Z(n4500) );
  IV U5868 ( .A(n4501), .Z(n4499) );
  XOR U5869 ( .A(n5937), .B(n4514), .Z(n4507) );
  XNOR U5870 ( .A(n4511), .B(n4504), .Z(n5937) );
  XOR U5871 ( .A(n5944), .B(n4509), .Z(n4511) );
  IV U5872 ( .A(n4513), .Z(n4509) );
  XOR U5873 ( .A(n5951), .B(n4515), .Z(n4516) );
  IV U5874 ( .A(n4517), .Z(n4515) );
  XOR U5875 ( .A(n5961), .B(n4906), .Z(n1995) );
  XOR U5876 ( .A(n5962), .B(n4617), .Z(n4583) );
  XOR U5877 ( .A(n5963), .B(n4543), .Z(n4535) );
  XOR U5878 ( .A(n5964), .B(n4529), .Z(n4524) );
  XNOR U5879 ( .A(n4527), .B(n4523), .Z(n5964) );
  XOR U5880 ( .A(n5971), .B(n4526), .Z(n4527) );
  IV U5881 ( .A(n4528), .Z(n4526) );
  XOR U5882 ( .A(n5978), .B(n4530), .Z(n4531) );
  IV U5883 ( .A(n4532), .Z(n4530) );
  XNOR U5884 ( .A(n4542), .B(n4534), .Z(n5963) );
  XOR U5885 ( .A(n5991), .B(n4547), .Z(n4542) );
  XOR U5886 ( .A(n5992), .B(n4538), .Z(n4539) );
  ANDN U5887 ( .B(n5995), .A(n5996), .Z(n5994) );
  XOR U5888 ( .A(n5993), .B(n5997), .Z(n5995) );
  XNOR U5889 ( .A(n4546), .B(n4541), .Z(n5991) );
  XOR U5890 ( .A(n6007), .B(n4551), .Z(n4546) );
  XNOR U5891 ( .A(n4549), .B(n4545), .Z(n6007) );
  XOR U5892 ( .A(n6014), .B(n4548), .Z(n4549) );
  IV U5893 ( .A(n4550), .Z(n4548) );
  XOR U5894 ( .A(n6021), .B(n4563), .Z(n4558) );
  XOR U5895 ( .A(n6022), .B(n4553), .Z(n4554) );
  IV U5896 ( .A(n4555), .Z(n4553) );
  XNOR U5897 ( .A(n4562), .B(n4557), .Z(n6021) );
  XOR U5898 ( .A(n6035), .B(n4567), .Z(n4562) );
  XNOR U5899 ( .A(n4565), .B(n4561), .Z(n6035) );
  XOR U5900 ( .A(n6042), .B(n4564), .Z(n4565) );
  IV U5901 ( .A(n4566), .Z(n4564) );
  XOR U5902 ( .A(n6049), .B(n4577), .Z(n4570) );
  XNOR U5903 ( .A(n4574), .B(n4569), .Z(n6049) );
  XOR U5904 ( .A(n6056), .B(n4572), .Z(n4574) );
  IV U5905 ( .A(n4576), .Z(n4572) );
  XOR U5906 ( .A(n6063), .B(n4578), .Z(n4579) );
  IV U5907 ( .A(n4580), .Z(n4578) );
  XNOR U5908 ( .A(n4616), .B(n4582), .Z(n5962) );
  XOR U5909 ( .A(n6076), .B(n4634), .Z(n4616) );
  XOR U5910 ( .A(n6077), .B(n4597), .Z(n4592) );
  XOR U5911 ( .A(n6078), .B(n4587), .Z(n4588) );
  IV U5912 ( .A(n4589), .Z(n4587) );
  XNOR U5913 ( .A(n4596), .B(n4591), .Z(n6077) );
  XOR U5914 ( .A(n6091), .B(n4601), .Z(n4596) );
  XNOR U5915 ( .A(n4599), .B(n4595), .Z(n6091) );
  XOR U5916 ( .A(n6098), .B(n4598), .Z(n4599) );
  IV U5917 ( .A(n4600), .Z(n4598) );
  XOR U5918 ( .A(n6105), .B(n4611), .Z(n4606) );
  XNOR U5919 ( .A(n4609), .B(n4603), .Z(n6105) );
  XNOR U5920 ( .A(n6109), .B(n6110), .Z(n4603) );
  ANDN U5921 ( .B(n6111), .A(n6112), .Z(n6110) );
  XOR U5922 ( .A(n6109), .B(n6113), .Z(n6111) );
  XOR U5923 ( .A(n6114), .B(n4608), .Z(n4609) );
  IV U5924 ( .A(n4610), .Z(n4608) );
  XOR U5925 ( .A(n6121), .B(n4612), .Z(n4613) );
  ANDN U5926 ( .B(n6124), .A(n6125), .Z(n6123) );
  XOR U5927 ( .A(n6122), .B(n6126), .Z(n6124) );
  XNOR U5928 ( .A(n4633), .B(n4615), .Z(n6076) );
  XOR U5929 ( .A(n6136), .B(n4641), .Z(n4633) );
  XOR U5930 ( .A(n6137), .B(n4628), .Z(n4623) );
  XNOR U5931 ( .A(n4626), .B(n4620), .Z(n6137) );
  XOR U5932 ( .A(n6144), .B(n4625), .Z(n4626) );
  IV U5933 ( .A(n4627), .Z(n4625) );
  XOR U5934 ( .A(n6151), .B(n4629), .Z(n4630) );
  ANDN U5935 ( .B(n6154), .A(n6155), .Z(n6153) );
  XOR U5936 ( .A(n6152), .B(n6156), .Z(n6154) );
  XNOR U5937 ( .A(n4640), .B(n4632), .Z(n6136) );
  XOR U5938 ( .A(n6166), .B(n4645), .Z(n4640) );
  XOR U5939 ( .A(n6167), .B(n4636), .Z(n4637) );
  ANDN U5940 ( .B(n6170), .A(n6171), .Z(n6169) );
  XOR U5941 ( .A(n6168), .B(n6172), .Z(n6170) );
  XNOR U5942 ( .A(n4644), .B(n4639), .Z(n6166) );
  XOR U5943 ( .A(n6182), .B(n4649), .Z(n4644) );
  XNOR U5944 ( .A(n4647), .B(n4643), .Z(n6182) );
  XOR U5945 ( .A(n6189), .B(n4646), .Z(n4647) );
  IV U5946 ( .A(n4648), .Z(n4646) );
  XOR U5947 ( .A(n6196), .B(n4698), .Z(n4679) );
  XOR U5948 ( .A(n6197), .B(n4661), .Z(n4656) );
  XOR U5949 ( .A(n6198), .B(n4652), .Z(n4653) );
  ANDN U5950 ( .B(n6201), .A(n6202), .Z(n6200) );
  XOR U5951 ( .A(n6199), .B(n6203), .Z(n6201) );
  XNOR U5952 ( .A(n4660), .B(n4655), .Z(n6197) );
  XOR U5953 ( .A(n6213), .B(n4665), .Z(n4660) );
  XNOR U5954 ( .A(n4663), .B(n4659), .Z(n6213) );
  XOR U5955 ( .A(n6220), .B(n4662), .Z(n4663) );
  IV U5956 ( .A(n4664), .Z(n4662) );
  XOR U5957 ( .A(n6227), .B(n4673), .Z(n4668) );
  XNOR U5958 ( .A(n4671), .B(n4667), .Z(n6227) );
  XOR U5959 ( .A(n6234), .B(n4670), .Z(n4671) );
  IV U5960 ( .A(n4672), .Z(n4670) );
  XOR U5961 ( .A(n6241), .B(n4674), .Z(n4675) );
  IV U5962 ( .A(n4676), .Z(n4674) );
  XNOR U5963 ( .A(n4697), .B(n4678), .Z(n6196) );
  XOR U5964 ( .A(n6254), .B(n4706), .Z(n4697) );
  XOR U5965 ( .A(n6255), .B(n4691), .Z(n4686) );
  XNOR U5966 ( .A(n4689), .B(n4683), .Z(n6255) );
  XOR U5967 ( .A(n6262), .B(n4688), .Z(n4689) );
  IV U5968 ( .A(n4690), .Z(n4688) );
  XOR U5969 ( .A(n6269), .B(n4692), .Z(n4693) );
  IV U5970 ( .A(n4694), .Z(n4692) );
  XNOR U5971 ( .A(n4705), .B(n4696), .Z(n6254) );
  XOR U5972 ( .A(n6282), .B(n4710), .Z(n4705) );
  XOR U5973 ( .A(n6283), .B(n4700), .Z(n4701) );
  IV U5974 ( .A(n4702), .Z(n4700) );
  XNOR U5975 ( .A(n4709), .B(n4704), .Z(n6282) );
  XOR U5976 ( .A(n6296), .B(n4714), .Z(n4709) );
  XNOR U5977 ( .A(n4712), .B(n4708), .Z(n6296) );
  XOR U5978 ( .A(n6303), .B(n4711), .Z(n4712) );
  IV U5979 ( .A(n4713), .Z(n4711) );
  XOR U5980 ( .A(n6310), .B(n4738), .Z(n4729) );
  XOR U5981 ( .A(n6311), .B(n4723), .Z(n4718) );
  XNOR U5982 ( .A(n4721), .B(n4717), .Z(n6311) );
  XOR U5983 ( .A(n6318), .B(n4720), .Z(n4721) );
  IV U5984 ( .A(n4722), .Z(n4720) );
  XOR U5985 ( .A(n6325), .B(n4724), .Z(n4725) );
  IV U5986 ( .A(n4726), .Z(n4724) );
  XNOR U5987 ( .A(n4737), .B(n4728), .Z(n6310) );
  XOR U5988 ( .A(n6338), .B(n4742), .Z(n4737) );
  XOR U5989 ( .A(n6339), .B(n4732), .Z(n4733) );
  IV U5990 ( .A(n4734), .Z(n4732) );
  XNOR U5991 ( .A(n4741), .B(n4736), .Z(n6338) );
  XOR U5992 ( .A(n6352), .B(n4746), .Z(n4741) );
  XNOR U5993 ( .A(n4744), .B(n4740), .Z(n6352) );
  XOR U5994 ( .A(n6359), .B(n4743), .Z(n4744) );
  IV U5995 ( .A(n4745), .Z(n4743) );
  XOR U5996 ( .A(n6366), .B(n4758), .Z(n4753) );
  XOR U5997 ( .A(n6367), .B(n4748), .Z(n4749) );
  IV U5998 ( .A(n4750), .Z(n4748) );
  XNOR U5999 ( .A(n4757), .B(n4752), .Z(n6366) );
  XOR U6000 ( .A(n6380), .B(n4762), .Z(n4757) );
  XNOR U6001 ( .A(n4760), .B(n4756), .Z(n6380) );
  XOR U6002 ( .A(n6387), .B(n4759), .Z(n4760) );
  IV U6003 ( .A(n4761), .Z(n4759) );
  XOR U6004 ( .A(n6394), .B(n4772), .Z(n4767) );
  XNOR U6005 ( .A(n4770), .B(n4764), .Z(n6394) );
  XOR U6006 ( .A(n6401), .B(n4769), .Z(n4770) );
  IV U6007 ( .A(n4771), .Z(n4769) );
  XOR U6008 ( .A(n6408), .B(n4773), .Z(n4774) );
  IV U6009 ( .A(n4775), .Z(n4773) );
  XNOR U6010 ( .A(n4905), .B(n5038), .Z(n5961) );
  XOR U6011 ( .A(n6418), .B(n4972), .Z(n4905) );
  XOR U6012 ( .A(n6419), .B(n4826), .Z(n4808) );
  XOR U6013 ( .A(n6420), .B(n4789), .Z(n4784) );
  XOR U6014 ( .A(n6421), .B(n4780), .Z(n4781) );
  ANDN U6015 ( .B(n6424), .A(n6425), .Z(n6423) );
  XOR U6016 ( .A(n6422), .B(n6426), .Z(n6424) );
  XNOR U6017 ( .A(n4788), .B(n4783), .Z(n6420) );
  XOR U6018 ( .A(n6436), .B(n4793), .Z(n4788) );
  XNOR U6019 ( .A(n4791), .B(n4787), .Z(n6436) );
  XOR U6020 ( .A(n6443), .B(n4790), .Z(n4791) );
  IV U6021 ( .A(n4792), .Z(n4790) );
  XOR U6022 ( .A(n6450), .B(n4803), .Z(n4798) );
  XNOR U6023 ( .A(n4801), .B(n4795), .Z(n6450) );
  XOR U6024 ( .A(n6457), .B(n4800), .Z(n4801) );
  IV U6025 ( .A(n4802), .Z(n4800) );
  XOR U6026 ( .A(n6464), .B(n4804), .Z(n4805) );
  ANDN U6027 ( .B(n6467), .A(n6468), .Z(n6466) );
  XOR U6028 ( .A(n6465), .B(n6469), .Z(n6467) );
  XNOR U6029 ( .A(n4825), .B(n4807), .Z(n6419) );
  XOR U6030 ( .A(n6479), .B(n4833), .Z(n4825) );
  XOR U6031 ( .A(n6480), .B(n4820), .Z(n4815) );
  XNOR U6032 ( .A(n4818), .B(n4812), .Z(n6480) );
  XOR U6033 ( .A(n6487), .B(n4817), .Z(n4818) );
  IV U6034 ( .A(n4819), .Z(n4817) );
  XOR U6035 ( .A(n6494), .B(n4821), .Z(n4822) );
  ANDN U6036 ( .B(n6497), .A(n6498), .Z(n6496) );
  XOR U6037 ( .A(n6495), .B(n6499), .Z(n6497) );
  XNOR U6038 ( .A(n4832), .B(n4824), .Z(n6479) );
  XOR U6039 ( .A(n6509), .B(n4837), .Z(n4832) );
  XOR U6040 ( .A(n6510), .B(n4828), .Z(n4829) );
  ANDN U6041 ( .B(n6513), .A(n6514), .Z(n6512) );
  XOR U6042 ( .A(n6511), .B(n6515), .Z(n6513) );
  XNOR U6043 ( .A(n4836), .B(n4831), .Z(n6509) );
  XOR U6044 ( .A(n6525), .B(n4841), .Z(n4836) );
  XNOR U6045 ( .A(n4839), .B(n4835), .Z(n6525) );
  XOR U6046 ( .A(n6532), .B(n4838), .Z(n4839) );
  IV U6047 ( .A(n4840), .Z(n4838) );
  XOR U6048 ( .A(n6539), .B(n4866), .Z(n4857) );
  XOR U6049 ( .A(n6540), .B(n4852), .Z(n4847) );
  XNOR U6050 ( .A(n4850), .B(n4844), .Z(n6540) );
  XOR U6051 ( .A(n6547), .B(n4849), .Z(n4850) );
  IV U6052 ( .A(n4851), .Z(n4849) );
  XOR U6053 ( .A(n6554), .B(n4853), .Z(n4854) );
  ANDN U6054 ( .B(n6557), .A(n6558), .Z(n6556) );
  XOR U6055 ( .A(n6555), .B(n6559), .Z(n6557) );
  XNOR U6056 ( .A(n4865), .B(n4856), .Z(n6539) );
  XOR U6057 ( .A(n6569), .B(n4870), .Z(n4865) );
  XOR U6058 ( .A(n6570), .B(n4860), .Z(n4861) );
  IV U6059 ( .A(n4862), .Z(n4860) );
  XNOR U6060 ( .A(n4869), .B(n4864), .Z(n6569) );
  XOR U6061 ( .A(n6583), .B(n4874), .Z(n4869) );
  XNOR U6062 ( .A(n4872), .B(n4868), .Z(n6583) );
  XOR U6063 ( .A(n6590), .B(n4871), .Z(n4872) );
  IV U6064 ( .A(n4873), .Z(n4871) );
  XOR U6065 ( .A(n6597), .B(n4888), .Z(n4883) );
  XOR U6066 ( .A(n6598), .B(n4876), .Z(n4877) );
  IV U6067 ( .A(n4878), .Z(n4876) );
  XNOR U6068 ( .A(n4887), .B(n4880), .Z(n6597) );
  XOR U6069 ( .A(n6611), .B(n4892), .Z(n4887) );
  XNOR U6070 ( .A(n4890), .B(n4886), .Z(n6611) );
  XOR U6071 ( .A(n6618), .B(n4889), .Z(n4890) );
  IV U6072 ( .A(n4891), .Z(n4889) );
  XOR U6073 ( .A(n6625), .B(n4900), .Z(n4895) );
  XNOR U6074 ( .A(n4898), .B(n4894), .Z(n6625) );
  XOR U6075 ( .A(n6632), .B(n4897), .Z(n4898) );
  IV U6076 ( .A(n4899), .Z(n4897) );
  XOR U6077 ( .A(n6639), .B(n4901), .Z(n4902) );
  ANDN U6078 ( .B(n6642), .A(n6643), .Z(n6641) );
  XOR U6079 ( .A(n6640), .B(n6644), .Z(n6642) );
  XNOR U6080 ( .A(n4971), .B(n4904), .Z(n6418) );
  XOR U6081 ( .A(n6654), .B(n5006), .Z(n4971) );
  XOR U6082 ( .A(n6655), .B(n4930), .Z(n4922) );
  XOR U6083 ( .A(n6656), .B(n4916), .Z(n4911) );
  XNOR U6084 ( .A(n4914), .B(n4910), .Z(n6656) );
  XOR U6085 ( .A(n6663), .B(n4913), .Z(n4914) );
  IV U6086 ( .A(n4915), .Z(n4913) );
  XOR U6087 ( .A(n6670), .B(n4917), .Z(n4918) );
  IV U6088 ( .A(n4919), .Z(n4917) );
  XNOR U6089 ( .A(n4929), .B(n4921), .Z(n6655) );
  XOR U6090 ( .A(n6683), .B(n4934), .Z(n4929) );
  XOR U6091 ( .A(n6684), .B(n4925), .Z(n4926) );
  ANDN U6092 ( .B(n6687), .A(n6688), .Z(n6686) );
  XOR U6093 ( .A(n6685), .B(n6689), .Z(n6687) );
  XNOR U6094 ( .A(n4933), .B(n4928), .Z(n6683) );
  XOR U6095 ( .A(n6699), .B(n4938), .Z(n4933) );
  XNOR U6096 ( .A(n4936), .B(n4932), .Z(n6699) );
  XOR U6097 ( .A(n6706), .B(n4935), .Z(n4936) );
  IV U6098 ( .A(n4937), .Z(n4935) );
  XOR U6099 ( .A(n6713), .B(n4951), .Z(n4947) );
  XOR U6100 ( .A(n6714), .B(n4940), .Z(n4941) );
  IV U6101 ( .A(n4942), .Z(n4940) );
  XNOR U6102 ( .A(n4950), .B(n4944), .Z(n6713) );
  XOR U6103 ( .A(n6727), .B(n4955), .Z(n4950) );
  XOR U6104 ( .A(n6734), .B(n4952), .Z(n4953) );
  IV U6105 ( .A(n4954), .Z(n4952) );
  XOR U6106 ( .A(n6741), .B(n4965), .Z(n4960) );
  XNOR U6107 ( .A(n4963), .B(n4957), .Z(n6741) );
  XOR U6108 ( .A(n6748), .B(n4962), .Z(n4963) );
  IV U6109 ( .A(n4964), .Z(n4962) );
  XOR U6110 ( .A(n6755), .B(n4966), .Z(n4967) );
  IV U6111 ( .A(n4968), .Z(n4966) );
  XNOR U6112 ( .A(n5005), .B(n4970), .Z(n6654) );
  XOR U6113 ( .A(n6768), .B(n5022), .Z(n5005) );
  XOR U6114 ( .A(n6769), .B(n4985), .Z(n4980) );
  XOR U6115 ( .A(n6770), .B(n4975), .Z(n4976) );
  IV U6116 ( .A(n4977), .Z(n4975) );
  XNOR U6117 ( .A(n4984), .B(n4979), .Z(n6769) );
  XOR U6118 ( .A(n6783), .B(n4989), .Z(n4984) );
  XNOR U6119 ( .A(n4987), .B(n4983), .Z(n6783) );
  XOR U6120 ( .A(n6790), .B(n4986), .Z(n4987) );
  IV U6121 ( .A(n4988), .Z(n4986) );
  XOR U6122 ( .A(n6797), .B(n4999), .Z(n4994) );
  XNOR U6123 ( .A(n4997), .B(n4991), .Z(n6797) );
  XOR U6124 ( .A(n6804), .B(n4996), .Z(n4997) );
  IV U6125 ( .A(n4998), .Z(n4996) );
  XOR U6126 ( .A(n6811), .B(n5000), .Z(n5001) );
  IV U6127 ( .A(n5002), .Z(n5000) );
  XNOR U6128 ( .A(n5021), .B(n5004), .Z(n6768) );
  XOR U6129 ( .A(n6824), .B(n5029), .Z(n5021) );
  XOR U6130 ( .A(n6825), .B(n5017), .Z(n5012) );
  XNOR U6131 ( .A(n5015), .B(n5009), .Z(n6825) );
  XOR U6132 ( .A(n6832), .B(n5014), .Z(n5015) );
  IV U6133 ( .A(n5016), .Z(n5014) );
  XOR U6134 ( .A(n6839), .B(n5018), .Z(n5019) );
  ANDN U6135 ( .B(n6842), .A(n6843), .Z(n6841) );
  XOR U6136 ( .A(n6840), .B(n6844), .Z(n6842) );
  XOR U6137 ( .A(n6854), .B(n5033), .Z(n5028) );
  XOR U6138 ( .A(n6855), .B(n5024), .Z(n5025) );
  ANDN U6139 ( .B(n6858), .A(n6859), .Z(n6857) );
  XOR U6140 ( .A(n6856), .B(n6860), .Z(n6858) );
  XNOR U6141 ( .A(n5032), .B(n5027), .Z(n6854) );
  XOR U6142 ( .A(n6870), .B(n5037), .Z(n5032) );
  XNOR U6143 ( .A(n5035), .B(n5031), .Z(n6870) );
  XOR U6144 ( .A(n6877), .B(n5034), .Z(n5035) );
  IV U6145 ( .A(n5036), .Z(n5034) );
  XOR U6146 ( .A(n3018), .B(n3019), .Z(o[0]) );
  XNOR U6147 ( .A(n2558), .B(n2049), .Z(n3019) );
  XOR U6148 ( .A(n6887), .B(n2078), .Z(n2049) );
  XOR U6149 ( .A(n6888), .B(n2017), .Z(n2009) );
  XNOR U6150 ( .A(n2001), .B(n2000), .Z(n2017) );
  XNOR U6151 ( .A(n6889), .B(n2004), .Z(n2000) );
  XNOR U6152 ( .A(y[27]), .B(x[27]), .Z(n2004) );
  XNOR U6153 ( .A(n2003), .B(n1999), .Z(n6889) );
  XNOR U6154 ( .A(y[21]), .B(x[21]), .Z(n1999) );
  XNOR U6155 ( .A(n6890), .B(n2002), .Z(n2003) );
  XNOR U6156 ( .A(y[25]), .B(x[25]), .Z(n2002) );
  XNOR U6157 ( .A(y[26]), .B(x[26]), .Z(n6890) );
  XOR U6158 ( .A(n2007), .B(n2006), .Z(n2001) );
  XNOR U6159 ( .A(n6891), .B(n2005), .Z(n2006) );
  XNOR U6160 ( .A(y[22]), .B(x[22]), .Z(n2005) );
  XNOR U6161 ( .A(y[23]), .B(x[23]), .Z(n6891) );
  XOR U6162 ( .A(y[24]), .B(x[24]), .Z(n2007) );
  XNOR U6163 ( .A(n2016), .B(n2008), .Z(n6888) );
  XNOR U6164 ( .A(y[4]), .B(x[4]), .Z(n2008) );
  XNOR U6165 ( .A(n6892), .B(n2021), .Z(n2016) );
  XNOR U6166 ( .A(n2014), .B(n2013), .Z(n2021) );
  XNOR U6167 ( .A(n6893), .B(n2012), .Z(n2013) );
  XNOR U6168 ( .A(y[29]), .B(x[29]), .Z(n2012) );
  XNOR U6169 ( .A(y[30]), .B(x[30]), .Z(n6893) );
  XNOR U6170 ( .A(y[31]), .B(x[31]), .Z(n2014) );
  XNOR U6171 ( .A(n2020), .B(n2015), .Z(n6892) );
  XNOR U6172 ( .A(y[20]), .B(x[20]), .Z(n2015) );
  XNOR U6173 ( .A(n6894), .B(n2024), .Z(n2020) );
  XNOR U6174 ( .A(y[34]), .B(x[34]), .Z(n2024) );
  XNOR U6175 ( .A(n2023), .B(n2019), .Z(n6894) );
  XNOR U6176 ( .A(y[28]), .B(x[28]), .Z(n2019) );
  XNOR U6177 ( .A(n6895), .B(n2022), .Z(n2023) );
  XNOR U6178 ( .A(y[32]), .B(x[32]), .Z(n2022) );
  XNOR U6179 ( .A(y[33]), .B(x[33]), .Z(n6895) );
  XNOR U6180 ( .A(n2031), .B(n2030), .Z(n2010) );
  XNOR U6181 ( .A(n6896), .B(n2035), .Z(n2030) );
  XNOR U6182 ( .A(n2028), .B(n2027), .Z(n2035) );
  XNOR U6183 ( .A(n6897), .B(n2026), .Z(n2027) );
  XNOR U6184 ( .A(y[14]), .B(x[14]), .Z(n2026) );
  XNOR U6185 ( .A(y[15]), .B(x[15]), .Z(n6897) );
  XNOR U6186 ( .A(y[16]), .B(x[16]), .Z(n2028) );
  XNOR U6187 ( .A(n2034), .B(n2029), .Z(n6896) );
  XNOR U6188 ( .A(y[5]), .B(x[5]), .Z(n2029) );
  XNOR U6189 ( .A(n6898), .B(n2038), .Z(n2034) );
  XNOR U6190 ( .A(y[19]), .B(x[19]), .Z(n2038) );
  XNOR U6191 ( .A(n2037), .B(n2033), .Z(n6898) );
  XNOR U6192 ( .A(y[13]), .B(x[13]), .Z(n2033) );
  XNOR U6193 ( .A(n6899), .B(n2036), .Z(n2037) );
  XNOR U6194 ( .A(y[17]), .B(x[17]), .Z(n2036) );
  XNOR U6195 ( .A(y[18]), .B(x[18]), .Z(n6899) );
  XNOR U6196 ( .A(n2042), .B(n2041), .Z(n2031) );
  XNOR U6197 ( .A(n6900), .B(n2045), .Z(n2041) );
  XNOR U6198 ( .A(y[12]), .B(x[12]), .Z(n2045) );
  XNOR U6199 ( .A(n2044), .B(n2040), .Z(n6900) );
  XNOR U6200 ( .A(y[6]), .B(x[6]), .Z(n2040) );
  XNOR U6201 ( .A(n6901), .B(n2043), .Z(n2044) );
  XNOR U6202 ( .A(y[10]), .B(x[10]), .Z(n2043) );
  XNOR U6203 ( .A(y[11]), .B(x[11]), .Z(n6901) );
  XOR U6204 ( .A(n2048), .B(n2047), .Z(n2042) );
  XNOR U6205 ( .A(n6902), .B(n2046), .Z(n2047) );
  XNOR U6206 ( .A(y[7]), .B(x[7]), .Z(n2046) );
  XNOR U6207 ( .A(y[8]), .B(x[8]), .Z(n6902) );
  XOR U6208 ( .A(y[9]), .B(x[9]), .Z(n2048) );
  XOR U6209 ( .A(n2077), .B(n2050), .Z(n6887) );
  XNOR U6210 ( .A(y[2]), .B(x[2]), .Z(n2050) );
  XOR U6211 ( .A(n6903), .B(n2094), .Z(n2077) );
  XNOR U6212 ( .A(n2058), .B(n2057), .Z(n2094) );
  XNOR U6213 ( .A(n6904), .B(n2062), .Z(n2057) );
  XNOR U6214 ( .A(n2055), .B(n2054), .Z(n2062) );
  XNOR U6215 ( .A(n6905), .B(n2053), .Z(n2054) );
  XNOR U6216 ( .A(y[45]), .B(x[45]), .Z(n2053) );
  XNOR U6217 ( .A(y[46]), .B(x[46]), .Z(n6905) );
  XNOR U6218 ( .A(y[47]), .B(x[47]), .Z(n2055) );
  XNOR U6219 ( .A(n2061), .B(n2056), .Z(n6904) );
  XNOR U6220 ( .A(y[36]), .B(x[36]), .Z(n2056) );
  XNOR U6221 ( .A(n6906), .B(n2065), .Z(n2061) );
  XNOR U6222 ( .A(y[50]), .B(x[50]), .Z(n2065) );
  XNOR U6223 ( .A(n2064), .B(n2060), .Z(n6906) );
  XNOR U6224 ( .A(y[44]), .B(x[44]), .Z(n2060) );
  XNOR U6225 ( .A(n6907), .B(n2063), .Z(n2064) );
  XNOR U6226 ( .A(y[48]), .B(x[48]), .Z(n2063) );
  XNOR U6227 ( .A(y[49]), .B(x[49]), .Z(n6907) );
  XNOR U6228 ( .A(n2069), .B(n2068), .Z(n2058) );
  XNOR U6229 ( .A(n6908), .B(n2072), .Z(n2068) );
  XNOR U6230 ( .A(y[43]), .B(x[43]), .Z(n2072) );
  XNOR U6231 ( .A(n2071), .B(n2067), .Z(n6908) );
  XNOR U6232 ( .A(y[37]), .B(x[37]), .Z(n2067) );
  XNOR U6233 ( .A(n6909), .B(n2070), .Z(n2071) );
  XNOR U6234 ( .A(y[41]), .B(x[41]), .Z(n2070) );
  XNOR U6235 ( .A(y[42]), .B(x[42]), .Z(n6909) );
  XOR U6236 ( .A(n2075), .B(n2074), .Z(n2069) );
  XNOR U6237 ( .A(n6910), .B(n2073), .Z(n2074) );
  XNOR U6238 ( .A(y[38]), .B(x[38]), .Z(n2073) );
  XNOR U6239 ( .A(y[39]), .B(x[39]), .Z(n6910) );
  XOR U6240 ( .A(y[40]), .B(x[40]), .Z(n2075) );
  XOR U6241 ( .A(n2093), .B(n2076), .Z(n6903) );
  XNOR U6242 ( .A(y[3]), .B(x[3]), .Z(n2076) );
  XOR U6243 ( .A(n6911), .B(n2101), .Z(n2093) );
  XNOR U6244 ( .A(n2085), .B(n2084), .Z(n2101) );
  XNOR U6245 ( .A(n6912), .B(n2088), .Z(n2084) );
  XNOR U6246 ( .A(y[58]), .B(x[58]), .Z(n2088) );
  XNOR U6247 ( .A(n2087), .B(n2081), .Z(n6912) );
  XNOR U6248 ( .A(y[52]), .B(x[52]), .Z(n2081) );
  XNOR U6249 ( .A(n6913), .B(n2086), .Z(n2087) );
  XNOR U6250 ( .A(y[56]), .B(x[56]), .Z(n2086) );
  XNOR U6251 ( .A(y[57]), .B(x[57]), .Z(n6913) );
  XOR U6252 ( .A(n2091), .B(n2090), .Z(n2085) );
  XNOR U6253 ( .A(n6914), .B(n2089), .Z(n2090) );
  XNOR U6254 ( .A(y[53]), .B(x[53]), .Z(n2089) );
  XNOR U6255 ( .A(y[54]), .B(x[54]), .Z(n6914) );
  XOR U6256 ( .A(y[55]), .B(x[55]), .Z(n2091) );
  XNOR U6257 ( .A(n2100), .B(n2092), .Z(n6911) );
  XNOR U6258 ( .A(y[35]), .B(x[35]), .Z(n2092) );
  XNOR U6259 ( .A(n6915), .B(n2105), .Z(n2100) );
  XNOR U6260 ( .A(n2098), .B(n2097), .Z(n2105) );
  XNOR U6261 ( .A(n6916), .B(n2096), .Z(n2097) );
  XNOR U6262 ( .A(y[60]), .B(x[60]), .Z(n2096) );
  XNOR U6263 ( .A(y[61]), .B(x[61]), .Z(n6916) );
  XNOR U6264 ( .A(y[62]), .B(x[62]), .Z(n2098) );
  XNOR U6265 ( .A(n2104), .B(n2099), .Z(n6915) );
  XNOR U6266 ( .A(y[51]), .B(x[51]), .Z(n2099) );
  XNOR U6267 ( .A(n6917), .B(n2108), .Z(n2104) );
  XNOR U6268 ( .A(y[65]), .B(x[65]), .Z(n2108) );
  XNOR U6269 ( .A(n2107), .B(n2103), .Z(n6917) );
  XNOR U6270 ( .A(y[59]), .B(x[59]), .Z(n2103) );
  XNOR U6271 ( .A(n6918), .B(n2106), .Z(n2107) );
  XNOR U6272 ( .A(y[63]), .B(x[63]), .Z(n2106) );
  XNOR U6273 ( .A(y[64]), .B(x[64]), .Z(n6918) );
  XOR U6274 ( .A(n6919), .B(n2784), .Z(n2558) );
  XOR U6275 ( .A(n6920), .B(n2277), .Z(n2220) );
  XOR U6276 ( .A(n6921), .B(n2152), .Z(n2137) );
  XNOR U6277 ( .A(n2118), .B(n2117), .Z(n2152) );
  XNOR U6278 ( .A(n6922), .B(n2122), .Z(n2117) );
  XNOR U6279 ( .A(n2115), .B(n2114), .Z(n2122) );
  XNOR U6280 ( .A(n6923), .B(n2113), .Z(n2114) );
  XNOR U6281 ( .A(y[238]), .B(x[238]), .Z(n2113) );
  XNOR U6282 ( .A(y[239]), .B(x[239]), .Z(n6923) );
  XNOR U6283 ( .A(y[240]), .B(x[240]), .Z(n2115) );
  XNOR U6284 ( .A(n2121), .B(n2116), .Z(n6922) );
  XNOR U6285 ( .A(y[229]), .B(x[229]), .Z(n2116) );
  XNOR U6286 ( .A(n6924), .B(n2125), .Z(n2121) );
  XNOR U6287 ( .A(y[243]), .B(x[243]), .Z(n2125) );
  XNOR U6288 ( .A(n2124), .B(n2120), .Z(n6924) );
  XNOR U6289 ( .A(y[237]), .B(x[237]), .Z(n2120) );
  XNOR U6290 ( .A(n6925), .B(n2123), .Z(n2124) );
  XNOR U6291 ( .A(y[241]), .B(x[241]), .Z(n2123) );
  XNOR U6292 ( .A(y[242]), .B(x[242]), .Z(n6925) );
  XNOR U6293 ( .A(n2129), .B(n2128), .Z(n2118) );
  XNOR U6294 ( .A(n6926), .B(n2132), .Z(n2128) );
  XNOR U6295 ( .A(y[236]), .B(x[236]), .Z(n2132) );
  XNOR U6296 ( .A(n2131), .B(n2127), .Z(n6926) );
  XNOR U6297 ( .A(y[230]), .B(x[230]), .Z(n2127) );
  XNOR U6298 ( .A(n6927), .B(n2130), .Z(n2131) );
  XNOR U6299 ( .A(y[234]), .B(x[234]), .Z(n2130) );
  XNOR U6300 ( .A(y[235]), .B(x[235]), .Z(n6927) );
  XOR U6301 ( .A(n2135), .B(n2134), .Z(n2129) );
  XNOR U6302 ( .A(n6928), .B(n2133), .Z(n2134) );
  XNOR U6303 ( .A(y[231]), .B(x[231]), .Z(n2133) );
  XNOR U6304 ( .A(y[232]), .B(x[232]), .Z(n6928) );
  XOR U6305 ( .A(y[233]), .B(x[233]), .Z(n2135) );
  XOR U6306 ( .A(n2151), .B(n2136), .Z(n6921) );
  XNOR U6307 ( .A(y[196]), .B(x[196]), .Z(n2136) );
  XOR U6308 ( .A(n6929), .B(n2159), .Z(n2151) );
  XNOR U6309 ( .A(n2143), .B(n2142), .Z(n2159) );
  XNOR U6310 ( .A(n6930), .B(n2146), .Z(n2142) );
  XNOR U6311 ( .A(y[251]), .B(x[251]), .Z(n2146) );
  XNOR U6312 ( .A(n2145), .B(n2141), .Z(n6930) );
  XNOR U6313 ( .A(y[245]), .B(x[245]), .Z(n2141) );
  XNOR U6314 ( .A(n6931), .B(n2144), .Z(n2145) );
  XNOR U6315 ( .A(y[249]), .B(x[249]), .Z(n2144) );
  XNOR U6316 ( .A(y[250]), .B(x[250]), .Z(n6931) );
  XOR U6317 ( .A(n2149), .B(n2148), .Z(n2143) );
  XNOR U6318 ( .A(n6932), .B(n2147), .Z(n2148) );
  XNOR U6319 ( .A(y[246]), .B(x[246]), .Z(n2147) );
  XNOR U6320 ( .A(y[247]), .B(x[247]), .Z(n6932) );
  XOR U6321 ( .A(y[248]), .B(x[248]), .Z(n2149) );
  XNOR U6322 ( .A(n2158), .B(n2150), .Z(n6929) );
  XNOR U6323 ( .A(y[228]), .B(x[228]), .Z(n2150) );
  XNOR U6324 ( .A(n6933), .B(n2163), .Z(n2158) );
  XNOR U6325 ( .A(n2156), .B(n2155), .Z(n2163) );
  XNOR U6326 ( .A(n6934), .B(n2154), .Z(n2155) );
  XNOR U6327 ( .A(y[253]), .B(x[253]), .Z(n2154) );
  XNOR U6328 ( .A(y[254]), .B(x[254]), .Z(n6934) );
  XNOR U6329 ( .A(y[255]), .B(x[255]), .Z(n2156) );
  XNOR U6330 ( .A(n2162), .B(n2157), .Z(n6933) );
  XNOR U6331 ( .A(y[244]), .B(x[244]), .Z(n2157) );
  XNOR U6332 ( .A(n6935), .B(n2166), .Z(n2162) );
  XNOR U6333 ( .A(y[258]), .B(x[258]), .Z(n2166) );
  XNOR U6334 ( .A(n2165), .B(n2161), .Z(n6935) );
  XNOR U6335 ( .A(y[252]), .B(x[252]), .Z(n2161) );
  XNOR U6336 ( .A(n6936), .B(n2164), .Z(n2165) );
  XNOR U6337 ( .A(y[256]), .B(x[256]), .Z(n2164) );
  XNOR U6338 ( .A(y[257]), .B(x[257]), .Z(n6936) );
  XOR U6339 ( .A(n6937), .B(n2187), .Z(n2179) );
  XNOR U6340 ( .A(n2171), .B(n2170), .Z(n2187) );
  XNOR U6341 ( .A(n6938), .B(n2174), .Z(n2170) );
  XNOR U6342 ( .A(y[220]), .B(x[220]), .Z(n2174) );
  XNOR U6343 ( .A(n2173), .B(n2169), .Z(n6938) );
  XNOR U6344 ( .A(y[214]), .B(x[214]), .Z(n2169) );
  XNOR U6345 ( .A(n6939), .B(n2172), .Z(n2173) );
  XNOR U6346 ( .A(y[218]), .B(x[218]), .Z(n2172) );
  XNOR U6347 ( .A(y[219]), .B(x[219]), .Z(n6939) );
  XOR U6348 ( .A(n2177), .B(n2176), .Z(n2171) );
  XNOR U6349 ( .A(n6940), .B(n2175), .Z(n2176) );
  XNOR U6350 ( .A(y[215]), .B(x[215]), .Z(n2175) );
  XNOR U6351 ( .A(y[216]), .B(x[216]), .Z(n6940) );
  XOR U6352 ( .A(y[217]), .B(x[217]), .Z(n2177) );
  XNOR U6353 ( .A(n2186), .B(n2178), .Z(n6937) );
  XNOR U6354 ( .A(y[197]), .B(x[197]), .Z(n2178) );
  XNOR U6355 ( .A(n6941), .B(n2191), .Z(n2186) );
  XNOR U6356 ( .A(n2184), .B(n2183), .Z(n2191) );
  XNOR U6357 ( .A(n6942), .B(n2182), .Z(n2183) );
  XNOR U6358 ( .A(y[222]), .B(x[222]), .Z(n2182) );
  XNOR U6359 ( .A(y[223]), .B(x[223]), .Z(n6942) );
  XNOR U6360 ( .A(y[224]), .B(x[224]), .Z(n2184) );
  XNOR U6361 ( .A(n2190), .B(n2185), .Z(n6941) );
  XNOR U6362 ( .A(y[213]), .B(x[213]), .Z(n2185) );
  XNOR U6363 ( .A(n6943), .B(n2194), .Z(n2190) );
  XNOR U6364 ( .A(y[227]), .B(x[227]), .Z(n2194) );
  XNOR U6365 ( .A(n2193), .B(n2189), .Z(n6943) );
  XNOR U6366 ( .A(y[221]), .B(x[221]), .Z(n2189) );
  XNOR U6367 ( .A(n6944), .B(n2192), .Z(n2193) );
  XNOR U6368 ( .A(y[225]), .B(x[225]), .Z(n2192) );
  XNOR U6369 ( .A(y[226]), .B(x[226]), .Z(n6944) );
  XNOR U6370 ( .A(n2201), .B(n2200), .Z(n2180) );
  XNOR U6371 ( .A(n6945), .B(n2205), .Z(n2200) );
  XNOR U6372 ( .A(n2198), .B(n2197), .Z(n2205) );
  XNOR U6373 ( .A(n6946), .B(n2196), .Z(n2197) );
  XNOR U6374 ( .A(y[207]), .B(x[207]), .Z(n2196) );
  XNOR U6375 ( .A(y[208]), .B(x[208]), .Z(n6946) );
  XNOR U6376 ( .A(y[209]), .B(x[209]), .Z(n2198) );
  XNOR U6377 ( .A(n2204), .B(n2199), .Z(n6945) );
  XNOR U6378 ( .A(y[198]), .B(x[198]), .Z(n2199) );
  XNOR U6379 ( .A(n6947), .B(n2208), .Z(n2204) );
  XNOR U6380 ( .A(y[212]), .B(x[212]), .Z(n2208) );
  XNOR U6381 ( .A(n2207), .B(n2203), .Z(n6947) );
  XNOR U6382 ( .A(y[206]), .B(x[206]), .Z(n2203) );
  XNOR U6383 ( .A(n6948), .B(n2206), .Z(n2207) );
  XNOR U6384 ( .A(y[210]), .B(x[210]), .Z(n2206) );
  XNOR U6385 ( .A(y[211]), .B(x[211]), .Z(n6948) );
  XNOR U6386 ( .A(n2212), .B(n2211), .Z(n2201) );
  XNOR U6387 ( .A(n6949), .B(n2215), .Z(n2211) );
  XNOR U6388 ( .A(y[205]), .B(x[205]), .Z(n2215) );
  XNOR U6389 ( .A(n2214), .B(n2210), .Z(n6949) );
  XNOR U6390 ( .A(y[199]), .B(x[199]), .Z(n2210) );
  XNOR U6391 ( .A(n6950), .B(n2213), .Z(n2214) );
  XNOR U6392 ( .A(y[203]), .B(x[203]), .Z(n2213) );
  XNOR U6393 ( .A(y[204]), .B(x[204]), .Z(n6950) );
  XOR U6394 ( .A(n2218), .B(n2217), .Z(n2212) );
  XNOR U6395 ( .A(n6951), .B(n2216), .Z(n2217) );
  XNOR U6396 ( .A(y[200]), .B(x[200]), .Z(n2216) );
  XNOR U6397 ( .A(y[201]), .B(x[201]), .Z(n6951) );
  XOR U6398 ( .A(y[202]), .B(x[202]), .Z(n2218) );
  XOR U6399 ( .A(n2276), .B(n2219), .Z(n6920) );
  XNOR U6400 ( .A(y[67]), .B(x[67]), .Z(n2219) );
  XOR U6401 ( .A(n6952), .B(n2305), .Z(n2276) );
  XOR U6402 ( .A(n6953), .B(n2243), .Z(n2235) );
  XNOR U6403 ( .A(n2227), .B(n2226), .Z(n2243) );
  XNOR U6404 ( .A(n6954), .B(n2230), .Z(n2226) );
  XNOR U6405 ( .A(y[283]), .B(x[283]), .Z(n2230) );
  XNOR U6406 ( .A(n2229), .B(n2225), .Z(n6954) );
  XNOR U6407 ( .A(y[277]), .B(x[277]), .Z(n2225) );
  XNOR U6408 ( .A(n6955), .B(n2228), .Z(n2229) );
  XNOR U6409 ( .A(y[281]), .B(x[281]), .Z(n2228) );
  XNOR U6410 ( .A(y[282]), .B(x[282]), .Z(n6955) );
  XOR U6411 ( .A(n2233), .B(n2232), .Z(n2227) );
  XNOR U6412 ( .A(n6956), .B(n2231), .Z(n2232) );
  XNOR U6413 ( .A(y[278]), .B(x[278]), .Z(n2231) );
  XNOR U6414 ( .A(y[279]), .B(x[279]), .Z(n6956) );
  XOR U6415 ( .A(y[280]), .B(x[280]), .Z(n2233) );
  XNOR U6416 ( .A(n2242), .B(n2234), .Z(n6953) );
  XNOR U6417 ( .A(y[260]), .B(x[260]), .Z(n2234) );
  XNOR U6418 ( .A(n6957), .B(n2247), .Z(n2242) );
  XNOR U6419 ( .A(n2240), .B(n2239), .Z(n2247) );
  XNOR U6420 ( .A(n6958), .B(n2238), .Z(n2239) );
  XNOR U6421 ( .A(y[285]), .B(x[285]), .Z(n2238) );
  XNOR U6422 ( .A(y[286]), .B(x[286]), .Z(n6958) );
  XNOR U6423 ( .A(y[287]), .B(x[287]), .Z(n2240) );
  XNOR U6424 ( .A(n2246), .B(n2241), .Z(n6957) );
  XNOR U6425 ( .A(y[276]), .B(x[276]), .Z(n2241) );
  XNOR U6426 ( .A(n6959), .B(n2250), .Z(n2246) );
  XNOR U6427 ( .A(y[290]), .B(x[290]), .Z(n2250) );
  XNOR U6428 ( .A(n2249), .B(n2245), .Z(n6959) );
  XNOR U6429 ( .A(y[284]), .B(x[284]), .Z(n2245) );
  XNOR U6430 ( .A(n6960), .B(n2248), .Z(n2249) );
  XNOR U6431 ( .A(y[288]), .B(x[288]), .Z(n2248) );
  XNOR U6432 ( .A(y[289]), .B(x[289]), .Z(n6960) );
  XNOR U6433 ( .A(n2257), .B(n2256), .Z(n2236) );
  XNOR U6434 ( .A(n6961), .B(n2261), .Z(n2256) );
  XNOR U6435 ( .A(n2254), .B(n2253), .Z(n2261) );
  XNOR U6436 ( .A(n6962), .B(n2252), .Z(n2253) );
  XNOR U6437 ( .A(y[270]), .B(x[270]), .Z(n2252) );
  XNOR U6438 ( .A(y[271]), .B(x[271]), .Z(n6962) );
  XNOR U6439 ( .A(y[272]), .B(x[272]), .Z(n2254) );
  XNOR U6440 ( .A(n2260), .B(n2255), .Z(n6961) );
  XNOR U6441 ( .A(y[261]), .B(x[261]), .Z(n2255) );
  XNOR U6442 ( .A(n6963), .B(n2264), .Z(n2260) );
  XNOR U6443 ( .A(y[275]), .B(x[275]), .Z(n2264) );
  XNOR U6444 ( .A(n2263), .B(n2259), .Z(n6963) );
  XNOR U6445 ( .A(y[269]), .B(x[269]), .Z(n2259) );
  XNOR U6446 ( .A(n6964), .B(n2262), .Z(n2263) );
  XNOR U6447 ( .A(y[273]), .B(x[273]), .Z(n2262) );
  XNOR U6448 ( .A(y[274]), .B(x[274]), .Z(n6964) );
  XNOR U6449 ( .A(n2268), .B(n2267), .Z(n2257) );
  XNOR U6450 ( .A(n6965), .B(n2271), .Z(n2267) );
  XNOR U6451 ( .A(y[268]), .B(x[268]), .Z(n2271) );
  XNOR U6452 ( .A(n2270), .B(n2266), .Z(n6965) );
  XNOR U6453 ( .A(y[262]), .B(x[262]), .Z(n2266) );
  XNOR U6454 ( .A(n6966), .B(n2269), .Z(n2270) );
  XNOR U6455 ( .A(y[266]), .B(x[266]), .Z(n2269) );
  XNOR U6456 ( .A(y[267]), .B(x[267]), .Z(n6966) );
  XOR U6457 ( .A(n2274), .B(n2273), .Z(n2268) );
  XNOR U6458 ( .A(n6967), .B(n2272), .Z(n2273) );
  XNOR U6459 ( .A(y[263]), .B(x[263]), .Z(n2272) );
  XNOR U6460 ( .A(y[264]), .B(x[264]), .Z(n6967) );
  XOR U6461 ( .A(y[265]), .B(x[265]), .Z(n2274) );
  XOR U6462 ( .A(n2304), .B(n2275), .Z(n6952) );
  XNOR U6463 ( .A(y[195]), .B(x[195]), .Z(n2275) );
  XOR U6464 ( .A(n6968), .B(n2319), .Z(n2304) );
  XNOR U6465 ( .A(n2285), .B(n2284), .Z(n2319) );
  XNOR U6466 ( .A(n6969), .B(n2289), .Z(n2284) );
  XNOR U6467 ( .A(n2282), .B(n2281), .Z(n2289) );
  XNOR U6468 ( .A(n6970), .B(n2280), .Z(n2281) );
  XNOR U6469 ( .A(y[301]), .B(x[301]), .Z(n2280) );
  XNOR U6470 ( .A(y[302]), .B(x[302]), .Z(n6970) );
  XNOR U6471 ( .A(y[303]), .B(x[303]), .Z(n2282) );
  XNOR U6472 ( .A(n2288), .B(n2283), .Z(n6969) );
  XNOR U6473 ( .A(y[292]), .B(x[292]), .Z(n2283) );
  XNOR U6474 ( .A(n6971), .B(n2292), .Z(n2288) );
  XNOR U6475 ( .A(y[306]), .B(x[306]), .Z(n2292) );
  XNOR U6476 ( .A(n2291), .B(n2287), .Z(n6971) );
  XNOR U6477 ( .A(y[300]), .B(x[300]), .Z(n2287) );
  XNOR U6478 ( .A(n6972), .B(n2290), .Z(n2291) );
  XNOR U6479 ( .A(y[304]), .B(x[304]), .Z(n2290) );
  XNOR U6480 ( .A(y[305]), .B(x[305]), .Z(n6972) );
  XNOR U6481 ( .A(n2296), .B(n2295), .Z(n2285) );
  XNOR U6482 ( .A(n6973), .B(n2299), .Z(n2295) );
  XNOR U6483 ( .A(y[299]), .B(x[299]), .Z(n2299) );
  XNOR U6484 ( .A(n2298), .B(n2294), .Z(n6973) );
  XNOR U6485 ( .A(y[293]), .B(x[293]), .Z(n2294) );
  XNOR U6486 ( .A(n6974), .B(n2297), .Z(n2298) );
  XNOR U6487 ( .A(y[297]), .B(x[297]), .Z(n2297) );
  XNOR U6488 ( .A(y[298]), .B(x[298]), .Z(n6974) );
  XOR U6489 ( .A(n2302), .B(n2301), .Z(n2296) );
  XNOR U6490 ( .A(n6975), .B(n2300), .Z(n2301) );
  XNOR U6491 ( .A(y[294]), .B(x[294]), .Z(n2300) );
  XNOR U6492 ( .A(y[295]), .B(x[295]), .Z(n6975) );
  XOR U6493 ( .A(y[296]), .B(x[296]), .Z(n2302) );
  XOR U6494 ( .A(n2318), .B(n2303), .Z(n6968) );
  XNOR U6495 ( .A(y[259]), .B(x[259]), .Z(n2303) );
  XOR U6496 ( .A(n6976), .B(n2326), .Z(n2318) );
  XNOR U6497 ( .A(n2310), .B(n2309), .Z(n2326) );
  XNOR U6498 ( .A(n6977), .B(n2313), .Z(n2309) );
  XNOR U6499 ( .A(y[314]), .B(x[314]), .Z(n2313) );
  XNOR U6500 ( .A(n2312), .B(n2308), .Z(n6977) );
  XNOR U6501 ( .A(y[308]), .B(x[308]), .Z(n2308) );
  XNOR U6502 ( .A(n6978), .B(n2311), .Z(n2312) );
  XNOR U6503 ( .A(y[312]), .B(x[312]), .Z(n2311) );
  XNOR U6504 ( .A(y[313]), .B(x[313]), .Z(n6978) );
  XOR U6505 ( .A(n2316), .B(n2315), .Z(n2310) );
  XNOR U6506 ( .A(n6979), .B(n2314), .Z(n2315) );
  XNOR U6507 ( .A(y[309]), .B(x[309]), .Z(n2314) );
  XNOR U6508 ( .A(y[310]), .B(x[310]), .Z(n6979) );
  XOR U6509 ( .A(y[311]), .B(x[311]), .Z(n2316) );
  XNOR U6510 ( .A(n2325), .B(n2317), .Z(n6976) );
  XNOR U6511 ( .A(y[291]), .B(x[291]), .Z(n2317) );
  XNOR U6512 ( .A(n6980), .B(n2330), .Z(n2325) );
  XNOR U6513 ( .A(n2323), .B(n2322), .Z(n2330) );
  XNOR U6514 ( .A(n6981), .B(n2321), .Z(n2322) );
  XNOR U6515 ( .A(y[316]), .B(x[316]), .Z(n2321) );
  XNOR U6516 ( .A(y[317]), .B(x[317]), .Z(n6981) );
  XNOR U6517 ( .A(y[318]), .B(x[318]), .Z(n2323) );
  XNOR U6518 ( .A(n2329), .B(n2324), .Z(n6980) );
  XNOR U6519 ( .A(y[307]), .B(x[307]), .Z(n2324) );
  XNOR U6520 ( .A(n6982), .B(n2333), .Z(n2329) );
  XNOR U6521 ( .A(y[321]), .B(x[321]), .Z(n2333) );
  XNOR U6522 ( .A(n2332), .B(n2328), .Z(n6982) );
  XNOR U6523 ( .A(y[315]), .B(x[315]), .Z(n2328) );
  XNOR U6524 ( .A(n6983), .B(n2331), .Z(n2332) );
  XNOR U6525 ( .A(y[319]), .B(x[319]), .Z(n2331) );
  XNOR U6526 ( .A(y[320]), .B(x[320]), .Z(n6983) );
  XOR U6527 ( .A(n6984), .B(n2418), .Z(n2389) );
  XOR U6528 ( .A(n6985), .B(n2355), .Z(n2347) );
  XNOR U6529 ( .A(n2339), .B(n2338), .Z(n2355) );
  XNOR U6530 ( .A(n6986), .B(n2342), .Z(n2338) );
  XNOR U6531 ( .A(y[156]), .B(x[156]), .Z(n2342) );
  XNOR U6532 ( .A(n2341), .B(n2337), .Z(n6986) );
  XNOR U6533 ( .A(y[150]), .B(x[150]), .Z(n2337) );
  XNOR U6534 ( .A(n6987), .B(n2340), .Z(n2341) );
  XNOR U6535 ( .A(y[154]), .B(x[154]), .Z(n2340) );
  XNOR U6536 ( .A(y[155]), .B(x[155]), .Z(n6987) );
  XOR U6537 ( .A(n2345), .B(n2344), .Z(n2339) );
  XNOR U6538 ( .A(n6988), .B(n2343), .Z(n2344) );
  XNOR U6539 ( .A(y[151]), .B(x[151]), .Z(n2343) );
  XNOR U6540 ( .A(y[152]), .B(x[152]), .Z(n6988) );
  XOR U6541 ( .A(y[153]), .B(x[153]), .Z(n2345) );
  XNOR U6542 ( .A(n2354), .B(n2346), .Z(n6985) );
  XNOR U6543 ( .A(y[133]), .B(x[133]), .Z(n2346) );
  XNOR U6544 ( .A(n6989), .B(n2359), .Z(n2354) );
  XNOR U6545 ( .A(n2352), .B(n2351), .Z(n2359) );
  XNOR U6546 ( .A(n6990), .B(n2350), .Z(n2351) );
  XNOR U6547 ( .A(y[158]), .B(x[158]), .Z(n2350) );
  XNOR U6548 ( .A(y[159]), .B(x[159]), .Z(n6990) );
  XNOR U6549 ( .A(y[160]), .B(x[160]), .Z(n2352) );
  XNOR U6550 ( .A(n2358), .B(n2353), .Z(n6989) );
  XNOR U6551 ( .A(y[149]), .B(x[149]), .Z(n2353) );
  XNOR U6552 ( .A(n6991), .B(n2362), .Z(n2358) );
  XNOR U6553 ( .A(y[163]), .B(x[163]), .Z(n2362) );
  XNOR U6554 ( .A(n2361), .B(n2357), .Z(n6991) );
  XNOR U6555 ( .A(y[157]), .B(x[157]), .Z(n2357) );
  XNOR U6556 ( .A(n6992), .B(n2360), .Z(n2361) );
  XNOR U6557 ( .A(y[161]), .B(x[161]), .Z(n2360) );
  XNOR U6558 ( .A(y[162]), .B(x[162]), .Z(n6992) );
  XNOR U6559 ( .A(n2369), .B(n2368), .Z(n2348) );
  XNOR U6560 ( .A(n6993), .B(n2373), .Z(n2368) );
  XNOR U6561 ( .A(n2366), .B(n2365), .Z(n2373) );
  XNOR U6562 ( .A(n6994), .B(n2364), .Z(n2365) );
  XNOR U6563 ( .A(y[143]), .B(x[143]), .Z(n2364) );
  XNOR U6564 ( .A(y[144]), .B(x[144]), .Z(n6994) );
  XNOR U6565 ( .A(y[145]), .B(x[145]), .Z(n2366) );
  XNOR U6566 ( .A(n2372), .B(n2367), .Z(n6993) );
  XNOR U6567 ( .A(y[134]), .B(x[134]), .Z(n2367) );
  XNOR U6568 ( .A(n6995), .B(n2376), .Z(n2372) );
  XNOR U6569 ( .A(y[148]), .B(x[148]), .Z(n2376) );
  XNOR U6570 ( .A(n2375), .B(n2371), .Z(n6995) );
  XNOR U6571 ( .A(y[142]), .B(x[142]), .Z(n2371) );
  XNOR U6572 ( .A(n6996), .B(n2374), .Z(n2375) );
  XNOR U6573 ( .A(y[146]), .B(x[146]), .Z(n2374) );
  XNOR U6574 ( .A(y[147]), .B(x[147]), .Z(n6996) );
  XNOR U6575 ( .A(n2381), .B(n2380), .Z(n2369) );
  XNOR U6576 ( .A(n6997), .B(n2384), .Z(n2380) );
  XNOR U6577 ( .A(y[141]), .B(x[141]), .Z(n2384) );
  XNOR U6578 ( .A(n2383), .B(n2379), .Z(n6997) );
  XNOR U6579 ( .A(y[135]), .B(x[135]), .Z(n2379) );
  XNOR U6580 ( .A(n6998), .B(n2382), .Z(n2383) );
  XNOR U6581 ( .A(y[139]), .B(x[139]), .Z(n2382) );
  XNOR U6582 ( .A(y[140]), .B(x[140]), .Z(n6998) );
  XOR U6583 ( .A(n2387), .B(n2386), .Z(n2381) );
  XNOR U6584 ( .A(n6999), .B(n2385), .Z(n2386) );
  XNOR U6585 ( .A(y[136]), .B(x[136]), .Z(n2385) );
  XNOR U6586 ( .A(y[137]), .B(x[137]), .Z(n6999) );
  XOR U6587 ( .A(y[138]), .B(x[138]), .Z(n2387) );
  XOR U6588 ( .A(n2417), .B(n2388), .Z(n6984) );
  XNOR U6589 ( .A(y[68]), .B(x[68]), .Z(n2388) );
  XOR U6590 ( .A(n7000), .B(n2432), .Z(n2417) );
  XNOR U6591 ( .A(n2398), .B(n2397), .Z(n2432) );
  XNOR U6592 ( .A(n7001), .B(n2402), .Z(n2397) );
  XNOR U6593 ( .A(n2395), .B(n2394), .Z(n2402) );
  XNOR U6594 ( .A(n7002), .B(n2393), .Z(n2394) );
  XNOR U6595 ( .A(y[174]), .B(x[174]), .Z(n2393) );
  XNOR U6596 ( .A(y[175]), .B(x[175]), .Z(n7002) );
  XNOR U6597 ( .A(y[176]), .B(x[176]), .Z(n2395) );
  XNOR U6598 ( .A(n2401), .B(n2396), .Z(n7001) );
  XNOR U6599 ( .A(y[165]), .B(x[165]), .Z(n2396) );
  XNOR U6600 ( .A(n7003), .B(n2405), .Z(n2401) );
  XNOR U6601 ( .A(y[179]), .B(x[179]), .Z(n2405) );
  XNOR U6602 ( .A(n2404), .B(n2400), .Z(n7003) );
  XNOR U6603 ( .A(y[173]), .B(x[173]), .Z(n2400) );
  XNOR U6604 ( .A(n7004), .B(n2403), .Z(n2404) );
  XNOR U6605 ( .A(y[177]), .B(x[177]), .Z(n2403) );
  XNOR U6606 ( .A(y[178]), .B(x[178]), .Z(n7004) );
  XNOR U6607 ( .A(n2409), .B(n2408), .Z(n2398) );
  XNOR U6608 ( .A(n7005), .B(n2412), .Z(n2408) );
  XNOR U6609 ( .A(y[172]), .B(x[172]), .Z(n2412) );
  XNOR U6610 ( .A(n2411), .B(n2407), .Z(n7005) );
  XNOR U6611 ( .A(y[166]), .B(x[166]), .Z(n2407) );
  XNOR U6612 ( .A(n7006), .B(n2410), .Z(n2411) );
  XNOR U6613 ( .A(y[170]), .B(x[170]), .Z(n2410) );
  XNOR U6614 ( .A(y[171]), .B(x[171]), .Z(n7006) );
  XOR U6615 ( .A(n2415), .B(n2414), .Z(n2409) );
  XNOR U6616 ( .A(n7007), .B(n2413), .Z(n2414) );
  XNOR U6617 ( .A(y[167]), .B(x[167]), .Z(n2413) );
  XNOR U6618 ( .A(y[168]), .B(x[168]), .Z(n7007) );
  XOR U6619 ( .A(y[169]), .B(x[169]), .Z(n2415) );
  XOR U6620 ( .A(n2431), .B(n2416), .Z(n7000) );
  XNOR U6621 ( .A(y[132]), .B(x[132]), .Z(n2416) );
  XOR U6622 ( .A(n7008), .B(n2439), .Z(n2431) );
  XNOR U6623 ( .A(n2423), .B(n2422), .Z(n2439) );
  XNOR U6624 ( .A(n7009), .B(n2426), .Z(n2422) );
  XNOR U6625 ( .A(y[187]), .B(x[187]), .Z(n2426) );
  XNOR U6626 ( .A(n2425), .B(n2421), .Z(n7009) );
  XNOR U6627 ( .A(y[181]), .B(x[181]), .Z(n2421) );
  XNOR U6628 ( .A(n7010), .B(n2424), .Z(n2425) );
  XNOR U6629 ( .A(y[185]), .B(x[185]), .Z(n2424) );
  XNOR U6630 ( .A(y[186]), .B(x[186]), .Z(n7010) );
  XOR U6631 ( .A(n2429), .B(n2428), .Z(n2423) );
  XNOR U6632 ( .A(n7011), .B(n2427), .Z(n2428) );
  XNOR U6633 ( .A(y[182]), .B(x[182]), .Z(n2427) );
  XNOR U6634 ( .A(y[183]), .B(x[183]), .Z(n7011) );
  XOR U6635 ( .A(y[184]), .B(x[184]), .Z(n2429) );
  XNOR U6636 ( .A(n2438), .B(n2430), .Z(n7008) );
  XNOR U6637 ( .A(y[164]), .B(x[164]), .Z(n2430) );
  XNOR U6638 ( .A(n7012), .B(n2443), .Z(n2438) );
  XNOR U6639 ( .A(n2436), .B(n2435), .Z(n2443) );
  XNOR U6640 ( .A(n7013), .B(n2434), .Z(n2435) );
  XNOR U6641 ( .A(y[189]), .B(x[189]), .Z(n2434) );
  XNOR U6642 ( .A(y[190]), .B(x[190]), .Z(n7013) );
  XNOR U6643 ( .A(y[191]), .B(x[191]), .Z(n2436) );
  XNOR U6644 ( .A(n2442), .B(n2437), .Z(n7012) );
  XNOR U6645 ( .A(y[180]), .B(x[180]), .Z(n2437) );
  XNOR U6646 ( .A(n7014), .B(n2446), .Z(n2442) );
  XNOR U6647 ( .A(y[194]), .B(x[194]), .Z(n2446) );
  XNOR U6648 ( .A(n2445), .B(n2441), .Z(n7014) );
  XNOR U6649 ( .A(y[188]), .B(x[188]), .Z(n2441) );
  XNOR U6650 ( .A(n7015), .B(n2444), .Z(n2445) );
  XNOR U6651 ( .A(y[192]), .B(x[192]), .Z(n2444) );
  XNOR U6652 ( .A(y[193]), .B(x[193]), .Z(n7015) );
  XOR U6653 ( .A(n7016), .B(n2490), .Z(n2475) );
  XNOR U6654 ( .A(n2454), .B(n2453), .Z(n2490) );
  XNOR U6655 ( .A(n7017), .B(n2458), .Z(n2453) );
  XNOR U6656 ( .A(n2451), .B(n2450), .Z(n2458) );
  XNOR U6657 ( .A(n7018), .B(n2449), .Z(n2450) );
  XNOR U6658 ( .A(y[111]), .B(x[111]), .Z(n2449) );
  XNOR U6659 ( .A(y[112]), .B(x[112]), .Z(n7018) );
  XNOR U6660 ( .A(y[113]), .B(x[113]), .Z(n2451) );
  XNOR U6661 ( .A(n2457), .B(n2452), .Z(n7017) );
  XNOR U6662 ( .A(y[102]), .B(x[102]), .Z(n2452) );
  XNOR U6663 ( .A(n7019), .B(n2461), .Z(n2457) );
  XNOR U6664 ( .A(y[116]), .B(x[116]), .Z(n2461) );
  XNOR U6665 ( .A(n2460), .B(n2456), .Z(n7019) );
  XNOR U6666 ( .A(y[110]), .B(x[110]), .Z(n2456) );
  XNOR U6667 ( .A(n7020), .B(n2459), .Z(n2460) );
  XNOR U6668 ( .A(y[114]), .B(x[114]), .Z(n2459) );
  XNOR U6669 ( .A(y[115]), .B(x[115]), .Z(n7020) );
  XNOR U6670 ( .A(n2467), .B(n2466), .Z(n2454) );
  XNOR U6671 ( .A(n7021), .B(n2470), .Z(n2466) );
  XNOR U6672 ( .A(y[109]), .B(x[109]), .Z(n2470) );
  XNOR U6673 ( .A(n2469), .B(n2463), .Z(n7021) );
  XNOR U6674 ( .A(y[103]), .B(x[103]), .Z(n2463) );
  XNOR U6675 ( .A(n7022), .B(n2468), .Z(n2469) );
  XNOR U6676 ( .A(y[107]), .B(x[107]), .Z(n2468) );
  XNOR U6677 ( .A(y[108]), .B(x[108]), .Z(n7022) );
  XOR U6678 ( .A(n2473), .B(n2472), .Z(n2467) );
  XNOR U6679 ( .A(n7023), .B(n2471), .Z(n2472) );
  XNOR U6680 ( .A(y[104]), .B(x[104]), .Z(n2471) );
  XNOR U6681 ( .A(y[105]), .B(x[105]), .Z(n7023) );
  XOR U6682 ( .A(y[106]), .B(x[106]), .Z(n2473) );
  XOR U6683 ( .A(n2489), .B(n2474), .Z(n7016) );
  XNOR U6684 ( .A(y[69]), .B(x[69]), .Z(n2474) );
  XOR U6685 ( .A(n7024), .B(n2497), .Z(n2489) );
  XNOR U6686 ( .A(n2481), .B(n2480), .Z(n2497) );
  XNOR U6687 ( .A(n7025), .B(n2484), .Z(n2480) );
  XNOR U6688 ( .A(y[124]), .B(x[124]), .Z(n2484) );
  XNOR U6689 ( .A(n2483), .B(n2479), .Z(n7025) );
  XNOR U6690 ( .A(y[118]), .B(x[118]), .Z(n2479) );
  XNOR U6691 ( .A(n7026), .B(n2482), .Z(n2483) );
  XNOR U6692 ( .A(y[122]), .B(x[122]), .Z(n2482) );
  XNOR U6693 ( .A(y[123]), .B(x[123]), .Z(n7026) );
  XOR U6694 ( .A(n2487), .B(n2486), .Z(n2481) );
  XNOR U6695 ( .A(n7027), .B(n2485), .Z(n2486) );
  XNOR U6696 ( .A(y[119]), .B(x[119]), .Z(n2485) );
  XNOR U6697 ( .A(y[120]), .B(x[120]), .Z(n7027) );
  XOR U6698 ( .A(y[121]), .B(x[121]), .Z(n2487) );
  XNOR U6699 ( .A(n2496), .B(n2488), .Z(n7024) );
  XNOR U6700 ( .A(y[101]), .B(x[101]), .Z(n2488) );
  XNOR U6701 ( .A(n7028), .B(n2501), .Z(n2496) );
  XNOR U6702 ( .A(n2494), .B(n2493), .Z(n2501) );
  XNOR U6703 ( .A(n7029), .B(n2492), .Z(n2493) );
  XNOR U6704 ( .A(y[126]), .B(x[126]), .Z(n2492) );
  XNOR U6705 ( .A(y[127]), .B(x[127]), .Z(n7029) );
  XNOR U6706 ( .A(y[128]), .B(x[128]), .Z(n2494) );
  XNOR U6707 ( .A(n2500), .B(n2495), .Z(n7028) );
  XNOR U6708 ( .A(y[117]), .B(x[117]), .Z(n2495) );
  XNOR U6709 ( .A(n7030), .B(n2504), .Z(n2500) );
  XNOR U6710 ( .A(y[131]), .B(x[131]), .Z(n2504) );
  XNOR U6711 ( .A(n2503), .B(n2499), .Z(n7030) );
  XNOR U6712 ( .A(y[125]), .B(x[125]), .Z(n2499) );
  XNOR U6713 ( .A(n7031), .B(n2502), .Z(n2503) );
  XNOR U6714 ( .A(y[129]), .B(x[129]), .Z(n2502) );
  XNOR U6715 ( .A(y[130]), .B(x[130]), .Z(n7031) );
  XOR U6716 ( .A(n7032), .B(n2525), .Z(n2517) );
  XNOR U6717 ( .A(n2509), .B(n2508), .Z(n2525) );
  XNOR U6718 ( .A(n7033), .B(n2512), .Z(n2508) );
  XNOR U6719 ( .A(y[93]), .B(x[93]), .Z(n2512) );
  XNOR U6720 ( .A(n2511), .B(n2507), .Z(n7033) );
  XNOR U6721 ( .A(y[87]), .B(x[87]), .Z(n2507) );
  XNOR U6722 ( .A(n7034), .B(n2510), .Z(n2511) );
  XNOR U6723 ( .A(y[91]), .B(x[91]), .Z(n2510) );
  XNOR U6724 ( .A(y[92]), .B(x[92]), .Z(n7034) );
  XOR U6725 ( .A(n2515), .B(n2514), .Z(n2509) );
  XNOR U6726 ( .A(n7035), .B(n2513), .Z(n2514) );
  XNOR U6727 ( .A(y[88]), .B(x[88]), .Z(n2513) );
  XNOR U6728 ( .A(y[89]), .B(x[89]), .Z(n7035) );
  XOR U6729 ( .A(y[90]), .B(x[90]), .Z(n2515) );
  XNOR U6730 ( .A(n2524), .B(n2516), .Z(n7032) );
  XNOR U6731 ( .A(y[70]), .B(x[70]), .Z(n2516) );
  XNOR U6732 ( .A(n7036), .B(n2529), .Z(n2524) );
  XNOR U6733 ( .A(n2522), .B(n2521), .Z(n2529) );
  XNOR U6734 ( .A(n7037), .B(n2520), .Z(n2521) );
  XNOR U6735 ( .A(y[95]), .B(x[95]), .Z(n2520) );
  XNOR U6736 ( .A(y[96]), .B(x[96]), .Z(n7037) );
  XNOR U6737 ( .A(y[97]), .B(x[97]), .Z(n2522) );
  XNOR U6738 ( .A(n2528), .B(n2523), .Z(n7036) );
  XNOR U6739 ( .A(y[86]), .B(x[86]), .Z(n2523) );
  XNOR U6740 ( .A(n7038), .B(n2532), .Z(n2528) );
  XNOR U6741 ( .A(y[100]), .B(x[100]), .Z(n2532) );
  XNOR U6742 ( .A(n2531), .B(n2527), .Z(n7038) );
  XNOR U6743 ( .A(y[94]), .B(x[94]), .Z(n2527) );
  XNOR U6744 ( .A(n7039), .B(n2530), .Z(n2531) );
  XNOR U6745 ( .A(y[98]), .B(x[98]), .Z(n2530) );
  XNOR U6746 ( .A(y[99]), .B(x[99]), .Z(n7039) );
  XNOR U6747 ( .A(n2539), .B(n2538), .Z(n2518) );
  XNOR U6748 ( .A(n7040), .B(n2543), .Z(n2538) );
  XNOR U6749 ( .A(n2536), .B(n2535), .Z(n2543) );
  XNOR U6750 ( .A(n7041), .B(n2534), .Z(n2535) );
  XNOR U6751 ( .A(y[80]), .B(x[80]), .Z(n2534) );
  XNOR U6752 ( .A(y[81]), .B(x[81]), .Z(n7041) );
  XNOR U6753 ( .A(y[82]), .B(x[82]), .Z(n2536) );
  XNOR U6754 ( .A(n2542), .B(n2537), .Z(n7040) );
  XNOR U6755 ( .A(y[71]), .B(x[71]), .Z(n2537) );
  XNOR U6756 ( .A(n7042), .B(n2546), .Z(n2542) );
  XNOR U6757 ( .A(y[85]), .B(x[85]), .Z(n2546) );
  XNOR U6758 ( .A(n2545), .B(n2541), .Z(n7042) );
  XNOR U6759 ( .A(y[79]), .B(x[79]), .Z(n2541) );
  XNOR U6760 ( .A(n7043), .B(n2544), .Z(n2545) );
  XNOR U6761 ( .A(y[83]), .B(x[83]), .Z(n2544) );
  XNOR U6762 ( .A(y[84]), .B(x[84]), .Z(n7043) );
  XNOR U6763 ( .A(n2550), .B(n2549), .Z(n2539) );
  XNOR U6764 ( .A(n7044), .B(n2553), .Z(n2549) );
  XNOR U6765 ( .A(y[78]), .B(x[78]), .Z(n2553) );
  XNOR U6766 ( .A(n2552), .B(n2548), .Z(n7044) );
  XNOR U6767 ( .A(y[72]), .B(x[72]), .Z(n2548) );
  XNOR U6768 ( .A(n7045), .B(n2551), .Z(n2552) );
  XNOR U6769 ( .A(y[76]), .B(x[76]), .Z(n2551) );
  XNOR U6770 ( .A(y[77]), .B(x[77]), .Z(n7045) );
  XOR U6771 ( .A(n2556), .B(n2555), .Z(n2550) );
  XNOR U6772 ( .A(n7046), .B(n2554), .Z(n2555) );
  XNOR U6773 ( .A(y[73]), .B(x[73]), .Z(n2554) );
  XNOR U6774 ( .A(y[74]), .B(x[74]), .Z(n7046) );
  XOR U6775 ( .A(y[75]), .B(x[75]), .Z(n2556) );
  XOR U6776 ( .A(n2783), .B(n2557), .Z(n6919) );
  XNOR U6777 ( .A(y[1]), .B(x[1]), .Z(n2557) );
  XOR U6778 ( .A(n7047), .B(n2900), .Z(n2783) );
  XOR U6779 ( .A(n7048), .B(n2643), .Z(n2614) );
  XOR U6780 ( .A(n7049), .B(n2581), .Z(n2573) );
  XNOR U6781 ( .A(n2565), .B(n2564), .Z(n2581) );
  XNOR U6782 ( .A(n7050), .B(n2568), .Z(n2564) );
  XNOR U6783 ( .A(y[411]), .B(x[411]), .Z(n2568) );
  XNOR U6784 ( .A(n2567), .B(n2563), .Z(n7050) );
  XNOR U6785 ( .A(y[405]), .B(x[405]), .Z(n2563) );
  XNOR U6786 ( .A(n7051), .B(n2566), .Z(n2567) );
  XNOR U6787 ( .A(y[409]), .B(x[409]), .Z(n2566) );
  XNOR U6788 ( .A(y[410]), .B(x[410]), .Z(n7051) );
  XOR U6789 ( .A(n2571), .B(n2570), .Z(n2565) );
  XNOR U6790 ( .A(n7052), .B(n2569), .Z(n2570) );
  XNOR U6791 ( .A(y[406]), .B(x[406]), .Z(n2569) );
  XNOR U6792 ( .A(y[407]), .B(x[407]), .Z(n7052) );
  XOR U6793 ( .A(y[408]), .B(x[408]), .Z(n2571) );
  XNOR U6794 ( .A(n2580), .B(n2572), .Z(n7049) );
  XNOR U6795 ( .A(y[388]), .B(x[388]), .Z(n2572) );
  XNOR U6796 ( .A(n7053), .B(n2585), .Z(n2580) );
  XNOR U6797 ( .A(n2578), .B(n2577), .Z(n2585) );
  XNOR U6798 ( .A(n7054), .B(n2576), .Z(n2577) );
  XNOR U6799 ( .A(y[413]), .B(x[413]), .Z(n2576) );
  XNOR U6800 ( .A(y[414]), .B(x[414]), .Z(n7054) );
  XNOR U6801 ( .A(y[415]), .B(x[415]), .Z(n2578) );
  XNOR U6802 ( .A(n2584), .B(n2579), .Z(n7053) );
  XNOR U6803 ( .A(y[404]), .B(x[404]), .Z(n2579) );
  XNOR U6804 ( .A(n7055), .B(n2588), .Z(n2584) );
  XNOR U6805 ( .A(y[418]), .B(x[418]), .Z(n2588) );
  XNOR U6806 ( .A(n2587), .B(n2583), .Z(n7055) );
  XNOR U6807 ( .A(y[412]), .B(x[412]), .Z(n2583) );
  XNOR U6808 ( .A(n7056), .B(n2586), .Z(n2587) );
  XNOR U6809 ( .A(y[416]), .B(x[416]), .Z(n2586) );
  XNOR U6810 ( .A(y[417]), .B(x[417]), .Z(n7056) );
  XNOR U6811 ( .A(n2595), .B(n2594), .Z(n2574) );
  XNOR U6812 ( .A(n7057), .B(n2599), .Z(n2594) );
  XNOR U6813 ( .A(n2592), .B(n2591), .Z(n2599) );
  XNOR U6814 ( .A(n7058), .B(n2590), .Z(n2591) );
  XNOR U6815 ( .A(y[398]), .B(x[398]), .Z(n2590) );
  XNOR U6816 ( .A(y[399]), .B(x[399]), .Z(n7058) );
  XNOR U6817 ( .A(y[400]), .B(x[400]), .Z(n2592) );
  XNOR U6818 ( .A(n2598), .B(n2593), .Z(n7057) );
  XNOR U6819 ( .A(y[389]), .B(x[389]), .Z(n2593) );
  XNOR U6820 ( .A(n7059), .B(n2602), .Z(n2598) );
  XNOR U6821 ( .A(y[403]), .B(x[403]), .Z(n2602) );
  XNOR U6822 ( .A(n2601), .B(n2597), .Z(n7059) );
  XNOR U6823 ( .A(y[397]), .B(x[397]), .Z(n2597) );
  XNOR U6824 ( .A(n7060), .B(n2600), .Z(n2601) );
  XNOR U6825 ( .A(y[401]), .B(x[401]), .Z(n2600) );
  XNOR U6826 ( .A(y[402]), .B(x[402]), .Z(n7060) );
  XNOR U6827 ( .A(n2606), .B(n2605), .Z(n2595) );
  XNOR U6828 ( .A(n7061), .B(n2609), .Z(n2605) );
  XNOR U6829 ( .A(y[396]), .B(x[396]), .Z(n2609) );
  XNOR U6830 ( .A(n2608), .B(n2604), .Z(n7061) );
  XNOR U6831 ( .A(y[390]), .B(x[390]), .Z(n2604) );
  XNOR U6832 ( .A(n7062), .B(n2607), .Z(n2608) );
  XNOR U6833 ( .A(y[394]), .B(x[394]), .Z(n2607) );
  XNOR U6834 ( .A(y[395]), .B(x[395]), .Z(n7062) );
  XOR U6835 ( .A(n2612), .B(n2611), .Z(n2606) );
  XNOR U6836 ( .A(n7063), .B(n2610), .Z(n2611) );
  XNOR U6837 ( .A(y[391]), .B(x[391]), .Z(n2610) );
  XNOR U6838 ( .A(y[392]), .B(x[392]), .Z(n7063) );
  XOR U6839 ( .A(y[393]), .B(x[393]), .Z(n2612) );
  XOR U6840 ( .A(n2642), .B(n2613), .Z(n7048) );
  XNOR U6841 ( .A(y[323]), .B(x[323]), .Z(n2613) );
  XOR U6842 ( .A(n7064), .B(n2657), .Z(n2642) );
  XNOR U6843 ( .A(n2623), .B(n2622), .Z(n2657) );
  XNOR U6844 ( .A(n7065), .B(n2627), .Z(n2622) );
  XNOR U6845 ( .A(n2620), .B(n2619), .Z(n2627) );
  XNOR U6846 ( .A(n7066), .B(n2618), .Z(n2619) );
  XNOR U6847 ( .A(y[429]), .B(x[429]), .Z(n2618) );
  XNOR U6848 ( .A(y[430]), .B(x[430]), .Z(n7066) );
  XNOR U6849 ( .A(y[431]), .B(x[431]), .Z(n2620) );
  XNOR U6850 ( .A(n2626), .B(n2621), .Z(n7065) );
  XNOR U6851 ( .A(y[420]), .B(x[420]), .Z(n2621) );
  XNOR U6852 ( .A(n7067), .B(n2630), .Z(n2626) );
  XNOR U6853 ( .A(y[434]), .B(x[434]), .Z(n2630) );
  XNOR U6854 ( .A(n2629), .B(n2625), .Z(n7067) );
  XNOR U6855 ( .A(y[428]), .B(x[428]), .Z(n2625) );
  XNOR U6856 ( .A(n7068), .B(n2628), .Z(n2629) );
  XNOR U6857 ( .A(y[432]), .B(x[432]), .Z(n2628) );
  XNOR U6858 ( .A(y[433]), .B(x[433]), .Z(n7068) );
  XNOR U6859 ( .A(n2634), .B(n2633), .Z(n2623) );
  XNOR U6860 ( .A(n7069), .B(n2637), .Z(n2633) );
  XNOR U6861 ( .A(y[427]), .B(x[427]), .Z(n2637) );
  XNOR U6862 ( .A(n2636), .B(n2632), .Z(n7069) );
  XNOR U6863 ( .A(y[421]), .B(x[421]), .Z(n2632) );
  XNOR U6864 ( .A(n7070), .B(n2635), .Z(n2636) );
  XNOR U6865 ( .A(y[425]), .B(x[425]), .Z(n2635) );
  XNOR U6866 ( .A(y[426]), .B(x[426]), .Z(n7070) );
  XOR U6867 ( .A(n2640), .B(n2639), .Z(n2634) );
  XNOR U6868 ( .A(n7071), .B(n2638), .Z(n2639) );
  XNOR U6869 ( .A(y[422]), .B(x[422]), .Z(n2638) );
  XNOR U6870 ( .A(y[423]), .B(x[423]), .Z(n7071) );
  XOR U6871 ( .A(y[424]), .B(x[424]), .Z(n2640) );
  XOR U6872 ( .A(n2656), .B(n2641), .Z(n7064) );
  XNOR U6873 ( .A(y[387]), .B(x[387]), .Z(n2641) );
  XOR U6874 ( .A(n7072), .B(n2664), .Z(n2656) );
  XNOR U6875 ( .A(n2648), .B(n2647), .Z(n2664) );
  XNOR U6876 ( .A(n7073), .B(n2651), .Z(n2647) );
  XNOR U6877 ( .A(y[442]), .B(x[442]), .Z(n2651) );
  XNOR U6878 ( .A(n2650), .B(n2646), .Z(n7073) );
  XNOR U6879 ( .A(y[436]), .B(x[436]), .Z(n2646) );
  XNOR U6880 ( .A(n7074), .B(n2649), .Z(n2650) );
  XNOR U6881 ( .A(y[440]), .B(x[440]), .Z(n2649) );
  XNOR U6882 ( .A(y[441]), .B(x[441]), .Z(n7074) );
  XOR U6883 ( .A(n2654), .B(n2653), .Z(n2648) );
  XNOR U6884 ( .A(n7075), .B(n2652), .Z(n2653) );
  XNOR U6885 ( .A(y[437]), .B(x[437]), .Z(n2652) );
  XNOR U6886 ( .A(y[438]), .B(x[438]), .Z(n7075) );
  XOR U6887 ( .A(y[439]), .B(x[439]), .Z(n2654) );
  XNOR U6888 ( .A(n2663), .B(n2655), .Z(n7072) );
  XNOR U6889 ( .A(y[419]), .B(x[419]), .Z(n2655) );
  XNOR U6890 ( .A(n7076), .B(n2668), .Z(n2663) );
  XNOR U6891 ( .A(n2661), .B(n2660), .Z(n2668) );
  XNOR U6892 ( .A(n7077), .B(n2659), .Z(n2660) );
  XNOR U6893 ( .A(y[444]), .B(x[444]), .Z(n2659) );
  XNOR U6894 ( .A(y[445]), .B(x[445]), .Z(n7077) );
  XNOR U6895 ( .A(y[446]), .B(x[446]), .Z(n2661) );
  XNOR U6896 ( .A(n2667), .B(n2662), .Z(n7076) );
  XNOR U6897 ( .A(y[435]), .B(x[435]), .Z(n2662) );
  XNOR U6898 ( .A(n7078), .B(n2671), .Z(n2667) );
  XNOR U6899 ( .A(y[449]), .B(x[449]), .Z(n2671) );
  XNOR U6900 ( .A(n2670), .B(n2666), .Z(n7078) );
  XNOR U6901 ( .A(y[443]), .B(x[443]), .Z(n2666) );
  XNOR U6902 ( .A(n7079), .B(n2669), .Z(n2670) );
  XNOR U6903 ( .A(y[447]), .B(x[447]), .Z(n2669) );
  XNOR U6904 ( .A(y[448]), .B(x[448]), .Z(n7079) );
  XOR U6905 ( .A(n7080), .B(n2715), .Z(n2700) );
  XNOR U6906 ( .A(n2679), .B(n2678), .Z(n2715) );
  XNOR U6907 ( .A(n7081), .B(n2683), .Z(n2678) );
  XNOR U6908 ( .A(n2676), .B(n2675), .Z(n2683) );
  XNOR U6909 ( .A(n7082), .B(n2674), .Z(n2675) );
  XNOR U6910 ( .A(y[366]), .B(x[366]), .Z(n2674) );
  XNOR U6911 ( .A(y[367]), .B(x[367]), .Z(n7082) );
  XNOR U6912 ( .A(y[368]), .B(x[368]), .Z(n2676) );
  XNOR U6913 ( .A(n2682), .B(n2677), .Z(n7081) );
  XNOR U6914 ( .A(y[357]), .B(x[357]), .Z(n2677) );
  XNOR U6915 ( .A(n7083), .B(n2686), .Z(n2682) );
  XNOR U6916 ( .A(y[371]), .B(x[371]), .Z(n2686) );
  XNOR U6917 ( .A(n2685), .B(n2681), .Z(n7083) );
  XNOR U6918 ( .A(y[365]), .B(x[365]), .Z(n2681) );
  XNOR U6919 ( .A(n7084), .B(n2684), .Z(n2685) );
  XNOR U6920 ( .A(y[369]), .B(x[369]), .Z(n2684) );
  XNOR U6921 ( .A(y[370]), .B(x[370]), .Z(n7084) );
  XNOR U6922 ( .A(n2692), .B(n2691), .Z(n2679) );
  XNOR U6923 ( .A(n7085), .B(n2695), .Z(n2691) );
  XNOR U6924 ( .A(y[364]), .B(x[364]), .Z(n2695) );
  XNOR U6925 ( .A(n2694), .B(n2688), .Z(n7085) );
  XNOR U6926 ( .A(y[358]), .B(x[358]), .Z(n2688) );
  XNOR U6927 ( .A(n7086), .B(n2693), .Z(n2694) );
  XNOR U6928 ( .A(y[362]), .B(x[362]), .Z(n2693) );
  XNOR U6929 ( .A(y[363]), .B(x[363]), .Z(n7086) );
  XOR U6930 ( .A(n2698), .B(n2697), .Z(n2692) );
  XNOR U6931 ( .A(n7087), .B(n2696), .Z(n2697) );
  XNOR U6932 ( .A(y[359]), .B(x[359]), .Z(n2696) );
  XNOR U6933 ( .A(y[360]), .B(x[360]), .Z(n7087) );
  XOR U6934 ( .A(y[361]), .B(x[361]), .Z(n2698) );
  XOR U6935 ( .A(n2714), .B(n2699), .Z(n7080) );
  XNOR U6936 ( .A(y[324]), .B(x[324]), .Z(n2699) );
  XOR U6937 ( .A(n7088), .B(n2722), .Z(n2714) );
  XNOR U6938 ( .A(n2706), .B(n2705), .Z(n2722) );
  XNOR U6939 ( .A(n7089), .B(n2709), .Z(n2705) );
  XNOR U6940 ( .A(y[379]), .B(x[379]), .Z(n2709) );
  XNOR U6941 ( .A(n2708), .B(n2704), .Z(n7089) );
  XNOR U6942 ( .A(y[373]), .B(x[373]), .Z(n2704) );
  XNOR U6943 ( .A(n7090), .B(n2707), .Z(n2708) );
  XNOR U6944 ( .A(y[377]), .B(x[377]), .Z(n2707) );
  XNOR U6945 ( .A(y[378]), .B(x[378]), .Z(n7090) );
  XOR U6946 ( .A(n2712), .B(n2711), .Z(n2706) );
  XNOR U6947 ( .A(n7091), .B(n2710), .Z(n2711) );
  XNOR U6948 ( .A(y[374]), .B(x[374]), .Z(n2710) );
  XNOR U6949 ( .A(y[375]), .B(x[375]), .Z(n7091) );
  XOR U6950 ( .A(y[376]), .B(x[376]), .Z(n2712) );
  XNOR U6951 ( .A(n2721), .B(n2713), .Z(n7088) );
  XNOR U6952 ( .A(y[356]), .B(x[356]), .Z(n2713) );
  XNOR U6953 ( .A(n7092), .B(n2726), .Z(n2721) );
  XNOR U6954 ( .A(n2719), .B(n2718), .Z(n2726) );
  XNOR U6955 ( .A(n7093), .B(n2717), .Z(n2718) );
  XNOR U6956 ( .A(y[381]), .B(x[381]), .Z(n2717) );
  XNOR U6957 ( .A(y[382]), .B(x[382]), .Z(n7093) );
  XNOR U6958 ( .A(y[383]), .B(x[383]), .Z(n2719) );
  XNOR U6959 ( .A(n2725), .B(n2720), .Z(n7092) );
  XNOR U6960 ( .A(y[372]), .B(x[372]), .Z(n2720) );
  XNOR U6961 ( .A(n7094), .B(n2729), .Z(n2725) );
  XNOR U6962 ( .A(y[386]), .B(x[386]), .Z(n2729) );
  XNOR U6963 ( .A(n2728), .B(n2724), .Z(n7094) );
  XNOR U6964 ( .A(y[380]), .B(x[380]), .Z(n2724) );
  XNOR U6965 ( .A(n7095), .B(n2727), .Z(n2728) );
  XNOR U6966 ( .A(y[384]), .B(x[384]), .Z(n2727) );
  XNOR U6967 ( .A(y[385]), .B(x[385]), .Z(n7095) );
  XOR U6968 ( .A(n7096), .B(n2750), .Z(n2742) );
  XNOR U6969 ( .A(n2734), .B(n2733), .Z(n2750) );
  XNOR U6970 ( .A(n7097), .B(n2737), .Z(n2733) );
  XNOR U6971 ( .A(y[348]), .B(x[348]), .Z(n2737) );
  XNOR U6972 ( .A(n2736), .B(n2732), .Z(n7097) );
  XNOR U6973 ( .A(y[342]), .B(x[342]), .Z(n2732) );
  XNOR U6974 ( .A(n7098), .B(n2735), .Z(n2736) );
  XNOR U6975 ( .A(y[346]), .B(x[346]), .Z(n2735) );
  XNOR U6976 ( .A(y[347]), .B(x[347]), .Z(n7098) );
  XOR U6977 ( .A(n2740), .B(n2739), .Z(n2734) );
  XNOR U6978 ( .A(n7099), .B(n2738), .Z(n2739) );
  XNOR U6979 ( .A(y[343]), .B(x[343]), .Z(n2738) );
  XNOR U6980 ( .A(y[344]), .B(x[344]), .Z(n7099) );
  XOR U6981 ( .A(y[345]), .B(x[345]), .Z(n2740) );
  XNOR U6982 ( .A(n2749), .B(n2741), .Z(n7096) );
  XNOR U6983 ( .A(y[325]), .B(x[325]), .Z(n2741) );
  XNOR U6984 ( .A(n7100), .B(n2754), .Z(n2749) );
  XNOR U6985 ( .A(n2747), .B(n2746), .Z(n2754) );
  XNOR U6986 ( .A(n7101), .B(n2745), .Z(n2746) );
  XNOR U6987 ( .A(y[350]), .B(x[350]), .Z(n2745) );
  XNOR U6988 ( .A(y[351]), .B(x[351]), .Z(n7101) );
  XNOR U6989 ( .A(y[352]), .B(x[352]), .Z(n2747) );
  XNOR U6990 ( .A(n2753), .B(n2748), .Z(n7100) );
  XNOR U6991 ( .A(y[341]), .B(x[341]), .Z(n2748) );
  XNOR U6992 ( .A(n7102), .B(n2757), .Z(n2753) );
  XNOR U6993 ( .A(y[355]), .B(x[355]), .Z(n2757) );
  XNOR U6994 ( .A(n2756), .B(n2752), .Z(n7102) );
  XNOR U6995 ( .A(y[349]), .B(x[349]), .Z(n2752) );
  XNOR U6996 ( .A(n7103), .B(n2755), .Z(n2756) );
  XNOR U6997 ( .A(y[353]), .B(x[353]), .Z(n2755) );
  XNOR U6998 ( .A(y[354]), .B(x[354]), .Z(n7103) );
  XNOR U6999 ( .A(n2764), .B(n2763), .Z(n2743) );
  XNOR U7000 ( .A(n7104), .B(n2768), .Z(n2763) );
  XNOR U7001 ( .A(n2761), .B(n2760), .Z(n2768) );
  XNOR U7002 ( .A(n7105), .B(n2759), .Z(n2760) );
  XNOR U7003 ( .A(y[335]), .B(x[335]), .Z(n2759) );
  XNOR U7004 ( .A(y[336]), .B(x[336]), .Z(n7105) );
  XNOR U7005 ( .A(y[337]), .B(x[337]), .Z(n2761) );
  XNOR U7006 ( .A(n2767), .B(n2762), .Z(n7104) );
  XNOR U7007 ( .A(y[326]), .B(x[326]), .Z(n2762) );
  XNOR U7008 ( .A(n7106), .B(n2771), .Z(n2767) );
  XNOR U7009 ( .A(y[340]), .B(x[340]), .Z(n2771) );
  XNOR U7010 ( .A(n2770), .B(n2766), .Z(n7106) );
  XNOR U7011 ( .A(y[334]), .B(x[334]), .Z(n2766) );
  XNOR U7012 ( .A(n7107), .B(n2769), .Z(n2770) );
  XNOR U7013 ( .A(y[338]), .B(x[338]), .Z(n2769) );
  XNOR U7014 ( .A(y[339]), .B(x[339]), .Z(n7107) );
  XNOR U7015 ( .A(n2775), .B(n2774), .Z(n2764) );
  XNOR U7016 ( .A(n7108), .B(n2778), .Z(n2774) );
  XNOR U7017 ( .A(y[333]), .B(x[333]), .Z(n2778) );
  XNOR U7018 ( .A(n2777), .B(n2773), .Z(n7108) );
  XNOR U7019 ( .A(y[327]), .B(x[327]), .Z(n2773) );
  XNOR U7020 ( .A(n7109), .B(n2776), .Z(n2777) );
  XNOR U7021 ( .A(y[331]), .B(x[331]), .Z(n2776) );
  XNOR U7022 ( .A(y[332]), .B(x[332]), .Z(n7109) );
  XOR U7023 ( .A(n2781), .B(n2780), .Z(n2775) );
  XNOR U7024 ( .A(n7110), .B(n2779), .Z(n2780) );
  XNOR U7025 ( .A(y[328]), .B(x[328]), .Z(n2779) );
  XNOR U7026 ( .A(y[329]), .B(x[329]), .Z(n7110) );
  XOR U7027 ( .A(y[330]), .B(x[330]), .Z(n2781) );
  XOR U7028 ( .A(n2899), .B(n2782), .Z(n7047) );
  XNOR U7029 ( .A(y[66]), .B(x[66]), .Z(n2782) );
  XOR U7030 ( .A(n7111), .B(n2956), .Z(n2899) );
  XOR U7031 ( .A(n7112), .B(n2827), .Z(n2812) );
  XNOR U7032 ( .A(n2793), .B(n2792), .Z(n2827) );
  XNOR U7033 ( .A(n7113), .B(n2797), .Z(n2792) );
  XNOR U7034 ( .A(n2790), .B(n2789), .Z(n2797) );
  XNOR U7035 ( .A(n7114), .B(n2788), .Z(n2789) );
  XNOR U7036 ( .A(y[493]), .B(x[493]), .Z(n2788) );
  XNOR U7037 ( .A(y[494]), .B(x[494]), .Z(n7114) );
  XNOR U7038 ( .A(y[495]), .B(x[495]), .Z(n2790) );
  XNOR U7039 ( .A(n2796), .B(n2791), .Z(n7113) );
  XNOR U7040 ( .A(y[484]), .B(x[484]), .Z(n2791) );
  XNOR U7041 ( .A(n7115), .B(n2800), .Z(n2796) );
  XNOR U7042 ( .A(y[498]), .B(x[498]), .Z(n2800) );
  XNOR U7043 ( .A(n2799), .B(n2795), .Z(n7115) );
  XNOR U7044 ( .A(y[492]), .B(x[492]), .Z(n2795) );
  XNOR U7045 ( .A(n7116), .B(n2798), .Z(n2799) );
  XNOR U7046 ( .A(y[496]), .B(x[496]), .Z(n2798) );
  XNOR U7047 ( .A(y[497]), .B(x[497]), .Z(n7116) );
  XNOR U7048 ( .A(n2804), .B(n2803), .Z(n2793) );
  XNOR U7049 ( .A(n7117), .B(n2807), .Z(n2803) );
  XNOR U7050 ( .A(y[491]), .B(x[491]), .Z(n2807) );
  XNOR U7051 ( .A(n2806), .B(n2802), .Z(n7117) );
  XNOR U7052 ( .A(y[485]), .B(x[485]), .Z(n2802) );
  XNOR U7053 ( .A(n7118), .B(n2805), .Z(n2806) );
  XNOR U7054 ( .A(y[489]), .B(x[489]), .Z(n2805) );
  XNOR U7055 ( .A(y[490]), .B(x[490]), .Z(n7118) );
  XOR U7056 ( .A(n2810), .B(n2809), .Z(n2804) );
  XNOR U7057 ( .A(n7119), .B(n2808), .Z(n2809) );
  XNOR U7058 ( .A(y[486]), .B(x[486]), .Z(n2808) );
  XNOR U7059 ( .A(y[487]), .B(x[487]), .Z(n7119) );
  XOR U7060 ( .A(y[488]), .B(x[488]), .Z(n2810) );
  XOR U7061 ( .A(n2826), .B(n2811), .Z(n7112) );
  XNOR U7062 ( .A(y[451]), .B(x[451]), .Z(n2811) );
  XOR U7063 ( .A(n7120), .B(n2834), .Z(n2826) );
  XNOR U7064 ( .A(n2818), .B(n2817), .Z(n2834) );
  XNOR U7065 ( .A(n7121), .B(n2821), .Z(n2817) );
  XNOR U7066 ( .A(y[506]), .B(x[506]), .Z(n2821) );
  XNOR U7067 ( .A(n2820), .B(n2816), .Z(n7121) );
  XNOR U7068 ( .A(y[500]), .B(x[500]), .Z(n2816) );
  XNOR U7069 ( .A(n7122), .B(n2819), .Z(n2820) );
  XNOR U7070 ( .A(y[504]), .B(x[504]), .Z(n2819) );
  XNOR U7071 ( .A(y[505]), .B(x[505]), .Z(n7122) );
  XOR U7072 ( .A(n2824), .B(n2823), .Z(n2818) );
  XNOR U7073 ( .A(n7123), .B(n2822), .Z(n2823) );
  XNOR U7074 ( .A(y[501]), .B(x[501]), .Z(n2822) );
  XNOR U7075 ( .A(y[502]), .B(x[502]), .Z(n7123) );
  XOR U7076 ( .A(y[503]), .B(x[503]), .Z(n2824) );
  XNOR U7077 ( .A(n2833), .B(n2825), .Z(n7120) );
  XNOR U7078 ( .A(y[483]), .B(x[483]), .Z(n2825) );
  XNOR U7079 ( .A(n7124), .B(n2838), .Z(n2833) );
  XNOR U7080 ( .A(n2831), .B(n2830), .Z(n2838) );
  XNOR U7081 ( .A(n7125), .B(n2829), .Z(n2830) );
  XNOR U7082 ( .A(y[508]), .B(x[508]), .Z(n2829) );
  XNOR U7083 ( .A(y[509]), .B(x[509]), .Z(n7125) );
  XNOR U7084 ( .A(y[510]), .B(x[510]), .Z(n2831) );
  XNOR U7085 ( .A(n2837), .B(n2832), .Z(n7124) );
  XNOR U7086 ( .A(y[499]), .B(x[499]), .Z(n2832) );
  XNOR U7087 ( .A(n7126), .B(n2841), .Z(n2837) );
  XNOR U7088 ( .A(y[513]), .B(x[513]), .Z(n2841) );
  XNOR U7089 ( .A(n2840), .B(n2836), .Z(n7126) );
  XNOR U7090 ( .A(y[507]), .B(x[507]), .Z(n2836) );
  XNOR U7091 ( .A(n7127), .B(n2839), .Z(n2840) );
  XNOR U7092 ( .A(y[511]), .B(x[511]), .Z(n2839) );
  XNOR U7093 ( .A(y[512]), .B(x[512]), .Z(n7127) );
  XOR U7094 ( .A(n7128), .B(n2862), .Z(n2854) );
  XNOR U7095 ( .A(n2846), .B(n2845), .Z(n2862) );
  XNOR U7096 ( .A(n7129), .B(n2849), .Z(n2845) );
  XNOR U7097 ( .A(y[475]), .B(x[475]), .Z(n2849) );
  XNOR U7098 ( .A(n2848), .B(n2844), .Z(n7129) );
  XNOR U7099 ( .A(y[469]), .B(x[469]), .Z(n2844) );
  XNOR U7100 ( .A(n7130), .B(n2847), .Z(n2848) );
  XNOR U7101 ( .A(y[473]), .B(x[473]), .Z(n2847) );
  XNOR U7102 ( .A(y[474]), .B(x[474]), .Z(n7130) );
  XOR U7103 ( .A(n2852), .B(n2851), .Z(n2846) );
  XNOR U7104 ( .A(n7131), .B(n2850), .Z(n2851) );
  XNOR U7105 ( .A(y[470]), .B(x[470]), .Z(n2850) );
  XNOR U7106 ( .A(y[471]), .B(x[471]), .Z(n7131) );
  XOR U7107 ( .A(y[472]), .B(x[472]), .Z(n2852) );
  XNOR U7108 ( .A(n2861), .B(n2853), .Z(n7128) );
  XNOR U7109 ( .A(y[452]), .B(x[452]), .Z(n2853) );
  XNOR U7110 ( .A(n7132), .B(n2866), .Z(n2861) );
  XNOR U7111 ( .A(n2859), .B(n2858), .Z(n2866) );
  XNOR U7112 ( .A(n7133), .B(n2857), .Z(n2858) );
  XNOR U7113 ( .A(y[477]), .B(x[477]), .Z(n2857) );
  XNOR U7114 ( .A(y[478]), .B(x[478]), .Z(n7133) );
  XNOR U7115 ( .A(y[479]), .B(x[479]), .Z(n2859) );
  XNOR U7116 ( .A(n2865), .B(n2860), .Z(n7132) );
  XNOR U7117 ( .A(y[468]), .B(x[468]), .Z(n2860) );
  XNOR U7118 ( .A(n7134), .B(n2869), .Z(n2865) );
  XNOR U7119 ( .A(y[482]), .B(x[482]), .Z(n2869) );
  XNOR U7120 ( .A(n2868), .B(n2864), .Z(n7134) );
  XNOR U7121 ( .A(y[476]), .B(x[476]), .Z(n2864) );
  XNOR U7122 ( .A(n7135), .B(n2867), .Z(n2868) );
  XNOR U7123 ( .A(y[480]), .B(x[480]), .Z(n2867) );
  XNOR U7124 ( .A(y[481]), .B(x[481]), .Z(n7135) );
  XNOR U7125 ( .A(n2878), .B(n2877), .Z(n2855) );
  XNOR U7126 ( .A(n7136), .B(n2882), .Z(n2877) );
  XNOR U7127 ( .A(n2873), .B(n2872), .Z(n2882) );
  XNOR U7128 ( .A(n7137), .B(n2871), .Z(n2872) );
  XNOR U7129 ( .A(y[462]), .B(x[462]), .Z(n2871) );
  XNOR U7130 ( .A(y[463]), .B(x[463]), .Z(n7137) );
  XNOR U7131 ( .A(y[464]), .B(x[464]), .Z(n2873) );
  XNOR U7132 ( .A(n2881), .B(n2874), .Z(n7136) );
  XNOR U7133 ( .A(y[453]), .B(x[453]), .Z(n2874) );
  XNOR U7134 ( .A(n7138), .B(n2887), .Z(n2881) );
  XNOR U7135 ( .A(y[467]), .B(x[467]), .Z(n2887) );
  XNOR U7136 ( .A(n2886), .B(n2880), .Z(n7138) );
  XNOR U7137 ( .A(y[461]), .B(x[461]), .Z(n2880) );
  XNOR U7138 ( .A(n7139), .B(n2883), .Z(n2886) );
  XNOR U7139 ( .A(y[465]), .B(x[465]), .Z(n2883) );
  XNOR U7140 ( .A(y[466]), .B(x[466]), .Z(n7139) );
  XNOR U7141 ( .A(n2891), .B(n2890), .Z(n2878) );
  XNOR U7142 ( .A(n7140), .B(n2894), .Z(n2890) );
  XNOR U7143 ( .A(y[460]), .B(x[460]), .Z(n2894) );
  XNOR U7144 ( .A(n2893), .B(n2889), .Z(n7140) );
  XNOR U7145 ( .A(y[454]), .B(x[454]), .Z(n2889) );
  XNOR U7146 ( .A(n7141), .B(n2892), .Z(n2893) );
  XNOR U7147 ( .A(y[458]), .B(x[458]), .Z(n2892) );
  XNOR U7148 ( .A(y[459]), .B(x[459]), .Z(n7141) );
  XOR U7149 ( .A(n2897), .B(n2896), .Z(n2891) );
  XNOR U7150 ( .A(n7142), .B(n2895), .Z(n2896) );
  XNOR U7151 ( .A(y[455]), .B(x[455]), .Z(n2895) );
  XNOR U7152 ( .A(y[456]), .B(x[456]), .Z(n7142) );
  XOR U7153 ( .A(y[457]), .B(x[457]), .Z(n2897) );
  XOR U7154 ( .A(n2955), .B(n2898), .Z(n7111) );
  XNOR U7155 ( .A(y[322]), .B(x[322]), .Z(n2898) );
  XOR U7156 ( .A(n7143), .B(n2986), .Z(n2955) );
  XOR U7157 ( .A(n7144), .B(n2922), .Z(n2914) );
  XNOR U7158 ( .A(n2906), .B(n2905), .Z(n2922) );
  XNOR U7159 ( .A(n7145), .B(n2909), .Z(n2905) );
  XNOR U7160 ( .A(y[538]), .B(x[538]), .Z(n2909) );
  XNOR U7161 ( .A(n2908), .B(n2904), .Z(n7145) );
  XNOR U7162 ( .A(y[532]), .B(x[532]), .Z(n2904) );
  XNOR U7163 ( .A(n7146), .B(n2907), .Z(n2908) );
  XNOR U7164 ( .A(y[536]), .B(x[536]), .Z(n2907) );
  XNOR U7165 ( .A(y[537]), .B(x[537]), .Z(n7146) );
  XOR U7166 ( .A(n2912), .B(n2911), .Z(n2906) );
  XNOR U7167 ( .A(n7147), .B(n2910), .Z(n2911) );
  XNOR U7168 ( .A(y[533]), .B(x[533]), .Z(n2910) );
  XNOR U7169 ( .A(y[534]), .B(x[534]), .Z(n7147) );
  XOR U7170 ( .A(y[535]), .B(x[535]), .Z(n2912) );
  XNOR U7171 ( .A(n2921), .B(n2913), .Z(n7144) );
  XNOR U7172 ( .A(y[515]), .B(x[515]), .Z(n2913) );
  XNOR U7173 ( .A(n7148), .B(n2926), .Z(n2921) );
  XNOR U7174 ( .A(n2919), .B(n2918), .Z(n2926) );
  XNOR U7175 ( .A(n7149), .B(n2917), .Z(n2918) );
  XNOR U7176 ( .A(y[540]), .B(x[540]), .Z(n2917) );
  XNOR U7177 ( .A(y[541]), .B(x[541]), .Z(n7149) );
  XNOR U7178 ( .A(y[542]), .B(x[542]), .Z(n2919) );
  XNOR U7179 ( .A(n2925), .B(n2920), .Z(n7148) );
  XNOR U7180 ( .A(y[531]), .B(x[531]), .Z(n2920) );
  XNOR U7181 ( .A(n7150), .B(n2929), .Z(n2925) );
  XNOR U7182 ( .A(y[545]), .B(x[545]), .Z(n2929) );
  XNOR U7183 ( .A(n2928), .B(n2924), .Z(n7150) );
  XNOR U7184 ( .A(y[539]), .B(x[539]), .Z(n2924) );
  XNOR U7185 ( .A(n7151), .B(n2927), .Z(n2928) );
  XNOR U7186 ( .A(y[543]), .B(x[543]), .Z(n2927) );
  XNOR U7187 ( .A(y[544]), .B(x[544]), .Z(n7151) );
  XNOR U7188 ( .A(n2936), .B(n2935), .Z(n2915) );
  XNOR U7189 ( .A(n7152), .B(n2940), .Z(n2935) );
  XNOR U7190 ( .A(n2933), .B(n2932), .Z(n2940) );
  XNOR U7191 ( .A(n7153), .B(n2931), .Z(n2932) );
  XNOR U7192 ( .A(y[525]), .B(x[525]), .Z(n2931) );
  XNOR U7193 ( .A(y[526]), .B(x[526]), .Z(n7153) );
  XNOR U7194 ( .A(y[527]), .B(x[527]), .Z(n2933) );
  XNOR U7195 ( .A(n2939), .B(n2934), .Z(n7152) );
  XNOR U7196 ( .A(y[516]), .B(x[516]), .Z(n2934) );
  XNOR U7197 ( .A(n7154), .B(n2943), .Z(n2939) );
  XNOR U7198 ( .A(y[530]), .B(x[530]), .Z(n2943) );
  XNOR U7199 ( .A(n2942), .B(n2938), .Z(n7154) );
  XNOR U7200 ( .A(y[524]), .B(x[524]), .Z(n2938) );
  XNOR U7201 ( .A(n7155), .B(n2941), .Z(n2942) );
  XNOR U7202 ( .A(y[528]), .B(x[528]), .Z(n2941) );
  XNOR U7203 ( .A(y[529]), .B(x[529]), .Z(n7155) );
  XNOR U7204 ( .A(n2947), .B(n2946), .Z(n2936) );
  XNOR U7205 ( .A(n7156), .B(n2950), .Z(n2946) );
  XNOR U7206 ( .A(y[523]), .B(x[523]), .Z(n2950) );
  XNOR U7207 ( .A(n2949), .B(n2945), .Z(n7156) );
  XNOR U7208 ( .A(y[517]), .B(x[517]), .Z(n2945) );
  XNOR U7209 ( .A(n7157), .B(n2948), .Z(n2949) );
  XNOR U7210 ( .A(y[521]), .B(x[521]), .Z(n2948) );
  XNOR U7211 ( .A(y[522]), .B(x[522]), .Z(n7157) );
  XOR U7212 ( .A(n2953), .B(n2952), .Z(n2947) );
  XNOR U7213 ( .A(n7158), .B(n2951), .Z(n2952) );
  XNOR U7214 ( .A(y[518]), .B(x[518]), .Z(n2951) );
  XNOR U7215 ( .A(y[519]), .B(x[519]), .Z(n7158) );
  XOR U7216 ( .A(y[520]), .B(x[520]), .Z(n2953) );
  XOR U7217 ( .A(n2985), .B(n2954), .Z(n7143) );
  XNOR U7218 ( .A(y[450]), .B(x[450]), .Z(n2954) );
  XOR U7219 ( .A(n7159), .B(n3002), .Z(n2985) );
  XNOR U7220 ( .A(n2964), .B(n2963), .Z(n3002) );
  XNOR U7221 ( .A(n7160), .B(n2968), .Z(n2963) );
  XNOR U7222 ( .A(n2961), .B(n2960), .Z(n2968) );
  XNOR U7223 ( .A(n7161), .B(n2959), .Z(n2960) );
  XNOR U7224 ( .A(y[556]), .B(x[556]), .Z(n2959) );
  XNOR U7225 ( .A(y[557]), .B(x[557]), .Z(n7161) );
  XNOR U7226 ( .A(y[558]), .B(x[558]), .Z(n2961) );
  XNOR U7227 ( .A(n2967), .B(n2962), .Z(n7160) );
  XNOR U7228 ( .A(y[547]), .B(x[547]), .Z(n2962) );
  XNOR U7229 ( .A(n7162), .B(n2971), .Z(n2967) );
  XNOR U7230 ( .A(y[561]), .B(x[561]), .Z(n2971) );
  XNOR U7231 ( .A(n2970), .B(n2966), .Z(n7162) );
  XNOR U7232 ( .A(y[555]), .B(x[555]), .Z(n2966) );
  XNOR U7233 ( .A(n7163), .B(n2969), .Z(n2970) );
  XNOR U7234 ( .A(y[559]), .B(x[559]), .Z(n2969) );
  XNOR U7235 ( .A(y[560]), .B(x[560]), .Z(n7163) );
  XNOR U7236 ( .A(n2977), .B(n2976), .Z(n2964) );
  XNOR U7237 ( .A(n7164), .B(n2980), .Z(n2976) );
  XNOR U7238 ( .A(y[554]), .B(x[554]), .Z(n2980) );
  XNOR U7239 ( .A(n2979), .B(n2973), .Z(n7164) );
  XNOR U7240 ( .A(y[548]), .B(x[548]), .Z(n2973) );
  XNOR U7241 ( .A(n7165), .B(n2978), .Z(n2979) );
  XNOR U7242 ( .A(y[552]), .B(x[552]), .Z(n2978) );
  XNOR U7243 ( .A(y[553]), .B(x[553]), .Z(n7165) );
  XOR U7244 ( .A(n2983), .B(n2982), .Z(n2977) );
  XNOR U7245 ( .A(n7166), .B(n2981), .Z(n2982) );
  XNOR U7246 ( .A(y[549]), .B(x[549]), .Z(n2981) );
  XNOR U7247 ( .A(y[550]), .B(x[550]), .Z(n7166) );
  XOR U7248 ( .A(y[551]), .B(x[551]), .Z(n2983) );
  XOR U7249 ( .A(n3001), .B(n2984), .Z(n7159) );
  XNOR U7250 ( .A(y[514]), .B(x[514]), .Z(n2984) );
  XOR U7251 ( .A(n7167), .B(n3009), .Z(n3001) );
  XNOR U7252 ( .A(n2993), .B(n2992), .Z(n3009) );
  XNOR U7253 ( .A(n7168), .B(n2996), .Z(n2992) );
  XNOR U7254 ( .A(y[569]), .B(x[569]), .Z(n2996) );
  XNOR U7255 ( .A(n2995), .B(n2989), .Z(n7168) );
  XNOR U7256 ( .A(y[563]), .B(x[563]), .Z(n2989) );
  XNOR U7257 ( .A(n7169), .B(n2994), .Z(n2995) );
  XNOR U7258 ( .A(y[567]), .B(x[567]), .Z(n2994) );
  XNOR U7259 ( .A(y[568]), .B(x[568]), .Z(n7169) );
  XOR U7260 ( .A(n2999), .B(n2998), .Z(n2993) );
  XNOR U7261 ( .A(n7170), .B(n2997), .Z(n2998) );
  XNOR U7262 ( .A(y[564]), .B(x[564]), .Z(n2997) );
  XNOR U7263 ( .A(y[565]), .B(x[565]), .Z(n7170) );
  XOR U7264 ( .A(y[566]), .B(x[566]), .Z(n2999) );
  XNOR U7265 ( .A(n3008), .B(n3000), .Z(n7167) );
  XNOR U7266 ( .A(y[546]), .B(x[546]), .Z(n3000) );
  XNOR U7267 ( .A(n7171), .B(n3013), .Z(n3008) );
  XNOR U7268 ( .A(n3006), .B(n3005), .Z(n3013) );
  XNOR U7269 ( .A(n7172), .B(n3004), .Z(n3005) );
  XNOR U7270 ( .A(y[571]), .B(x[571]), .Z(n3004) );
  XNOR U7271 ( .A(y[572]), .B(x[572]), .Z(n7172) );
  XNOR U7272 ( .A(y[573]), .B(x[573]), .Z(n3006) );
  XNOR U7273 ( .A(n3012), .B(n3007), .Z(n7171) );
  XNOR U7274 ( .A(y[562]), .B(x[562]), .Z(n3007) );
  XNOR U7275 ( .A(n7173), .B(n3016), .Z(n3012) );
  XNOR U7276 ( .A(y[576]), .B(x[576]), .Z(n3016) );
  XNOR U7277 ( .A(n3015), .B(n3011), .Z(n7173) );
  XNOR U7278 ( .A(y[570]), .B(x[570]), .Z(n3011) );
  XNOR U7279 ( .A(n7174), .B(n3014), .Z(n3015) );
  XNOR U7280 ( .A(y[574]), .B(x[574]), .Z(n3014) );
  XNOR U7281 ( .A(y[575]), .B(x[575]), .Z(n7174) );
  XNOR U7282 ( .A(n7175), .B(n6886), .Z(n3018) );
  XOR U7283 ( .A(n7176), .B(n5384), .Z(n5267) );
  XOR U7284 ( .A(n7177), .B(n5125), .Z(n5094) );
  XOR U7285 ( .A(n7178), .B(n5061), .Z(n5053) );
  XNOR U7286 ( .A(n5045), .B(n5044), .Z(n5061) );
  XNOR U7287 ( .A(n7179), .B(n5048), .Z(n5044) );
  XNOR U7288 ( .A(y[923]), .B(x[923]), .Z(n5048) );
  XNOR U7289 ( .A(n5047), .B(n5043), .Z(n7179) );
  XNOR U7290 ( .A(y[917]), .B(x[917]), .Z(n5043) );
  XNOR U7291 ( .A(n7180), .B(n5046), .Z(n5047) );
  XNOR U7292 ( .A(y[921]), .B(x[921]), .Z(n5046) );
  XNOR U7293 ( .A(y[922]), .B(x[922]), .Z(n7180) );
  XOR U7294 ( .A(n5051), .B(n5050), .Z(n5045) );
  XNOR U7295 ( .A(n7181), .B(n5049), .Z(n5050) );
  XNOR U7296 ( .A(y[918]), .B(x[918]), .Z(n5049) );
  XNOR U7297 ( .A(y[919]), .B(x[919]), .Z(n7181) );
  XOR U7298 ( .A(y[920]), .B(x[920]), .Z(n5051) );
  XNOR U7299 ( .A(n5060), .B(n5052), .Z(n7178) );
  XNOR U7300 ( .A(y[900]), .B(x[900]), .Z(n5052) );
  XNOR U7301 ( .A(n7182), .B(n5065), .Z(n5060) );
  XNOR U7302 ( .A(n5058), .B(n5057), .Z(n5065) );
  XNOR U7303 ( .A(n7183), .B(n5056), .Z(n5057) );
  XNOR U7304 ( .A(y[925]), .B(x[925]), .Z(n5056) );
  XNOR U7305 ( .A(y[926]), .B(x[926]), .Z(n7183) );
  XNOR U7306 ( .A(y[927]), .B(x[927]), .Z(n5058) );
  XNOR U7307 ( .A(n5064), .B(n5059), .Z(n7182) );
  XNOR U7308 ( .A(y[916]), .B(x[916]), .Z(n5059) );
  XNOR U7309 ( .A(n7184), .B(n5068), .Z(n5064) );
  XNOR U7310 ( .A(y[930]), .B(x[930]), .Z(n5068) );
  XNOR U7311 ( .A(n5067), .B(n5063), .Z(n7184) );
  XNOR U7312 ( .A(y[924]), .B(x[924]), .Z(n5063) );
  XNOR U7313 ( .A(n7185), .B(n5066), .Z(n5067) );
  XNOR U7314 ( .A(y[928]), .B(x[928]), .Z(n5066) );
  XNOR U7315 ( .A(y[929]), .B(x[929]), .Z(n7185) );
  XNOR U7316 ( .A(n5075), .B(n5074), .Z(n5054) );
  XNOR U7317 ( .A(n7186), .B(n5079), .Z(n5074) );
  XNOR U7318 ( .A(n5072), .B(n5071), .Z(n5079) );
  XNOR U7319 ( .A(n7187), .B(n5070), .Z(n5071) );
  XNOR U7320 ( .A(y[910]), .B(x[910]), .Z(n5070) );
  XNOR U7321 ( .A(y[911]), .B(x[911]), .Z(n7187) );
  XNOR U7322 ( .A(y[912]), .B(x[912]), .Z(n5072) );
  XNOR U7323 ( .A(n5078), .B(n5073), .Z(n7186) );
  XNOR U7324 ( .A(y[901]), .B(x[901]), .Z(n5073) );
  XNOR U7325 ( .A(n7188), .B(n5082), .Z(n5078) );
  XNOR U7326 ( .A(y[915]), .B(x[915]), .Z(n5082) );
  XNOR U7327 ( .A(n5081), .B(n5077), .Z(n7188) );
  XNOR U7328 ( .A(y[909]), .B(x[909]), .Z(n5077) );
  XNOR U7329 ( .A(n7189), .B(n5080), .Z(n5081) );
  XNOR U7330 ( .A(y[913]), .B(x[913]), .Z(n5080) );
  XNOR U7331 ( .A(y[914]), .B(x[914]), .Z(n7189) );
  XNOR U7332 ( .A(n5086), .B(n5085), .Z(n5075) );
  XNOR U7333 ( .A(n7190), .B(n5089), .Z(n5085) );
  XNOR U7334 ( .A(y[908]), .B(x[908]), .Z(n5089) );
  XNOR U7335 ( .A(n5088), .B(n5084), .Z(n7190) );
  XNOR U7336 ( .A(y[902]), .B(x[902]), .Z(n5084) );
  XNOR U7337 ( .A(n7191), .B(n5087), .Z(n5088) );
  XNOR U7338 ( .A(y[906]), .B(x[906]), .Z(n5087) );
  XNOR U7339 ( .A(y[907]), .B(x[907]), .Z(n7191) );
  XOR U7340 ( .A(n5092), .B(n5091), .Z(n5086) );
  XNOR U7341 ( .A(n7192), .B(n5090), .Z(n5091) );
  XNOR U7342 ( .A(y[903]), .B(x[903]), .Z(n5090) );
  XNOR U7343 ( .A(y[904]), .B(x[904]), .Z(n7192) );
  XOR U7344 ( .A(y[905]), .B(x[905]), .Z(n5092) );
  XOR U7345 ( .A(n5124), .B(n5093), .Z(n7177) );
  XNOR U7346 ( .A(y[835]), .B(x[835]), .Z(n5093) );
  XOR U7347 ( .A(n7193), .B(n5141), .Z(n5124) );
  XNOR U7348 ( .A(n5103), .B(n5102), .Z(n5141) );
  XNOR U7349 ( .A(n7194), .B(n5107), .Z(n5102) );
  XNOR U7350 ( .A(n5100), .B(n5099), .Z(n5107) );
  XNOR U7351 ( .A(n7195), .B(n5098), .Z(n5099) );
  XNOR U7352 ( .A(y[941]), .B(x[941]), .Z(n5098) );
  XNOR U7353 ( .A(y[942]), .B(x[942]), .Z(n7195) );
  XNOR U7354 ( .A(y[943]), .B(x[943]), .Z(n5100) );
  XNOR U7355 ( .A(n5106), .B(n5101), .Z(n7194) );
  XNOR U7356 ( .A(y[932]), .B(x[932]), .Z(n5101) );
  XNOR U7357 ( .A(n7196), .B(n5110), .Z(n5106) );
  XNOR U7358 ( .A(y[946]), .B(x[946]), .Z(n5110) );
  XNOR U7359 ( .A(n5109), .B(n5105), .Z(n7196) );
  XNOR U7360 ( .A(y[940]), .B(x[940]), .Z(n5105) );
  XNOR U7361 ( .A(n7197), .B(n5108), .Z(n5109) );
  XNOR U7362 ( .A(y[944]), .B(x[944]), .Z(n5108) );
  XNOR U7363 ( .A(y[945]), .B(x[945]), .Z(n7197) );
  XNOR U7364 ( .A(n5116), .B(n5115), .Z(n5103) );
  XNOR U7365 ( .A(n7198), .B(n5119), .Z(n5115) );
  XNOR U7366 ( .A(y[939]), .B(x[939]), .Z(n5119) );
  XNOR U7367 ( .A(n5118), .B(n5112), .Z(n7198) );
  XNOR U7368 ( .A(y[933]), .B(x[933]), .Z(n5112) );
  XNOR U7369 ( .A(n7199), .B(n5117), .Z(n5118) );
  XNOR U7370 ( .A(y[937]), .B(x[937]), .Z(n5117) );
  XNOR U7371 ( .A(y[938]), .B(x[938]), .Z(n7199) );
  XOR U7372 ( .A(n5122), .B(n5121), .Z(n5116) );
  XNOR U7373 ( .A(n7200), .B(n5120), .Z(n5121) );
  XNOR U7374 ( .A(y[934]), .B(x[934]), .Z(n5120) );
  XNOR U7375 ( .A(y[935]), .B(x[935]), .Z(n7200) );
  XOR U7376 ( .A(y[936]), .B(x[936]), .Z(n5122) );
  XOR U7377 ( .A(n5140), .B(n5123), .Z(n7193) );
  XNOR U7378 ( .A(y[899]), .B(x[899]), .Z(n5123) );
  XOR U7379 ( .A(n7201), .B(n5148), .Z(n5140) );
  XNOR U7380 ( .A(n5132), .B(n5131), .Z(n5148) );
  XNOR U7381 ( .A(n7202), .B(n5135), .Z(n5131) );
  XNOR U7382 ( .A(y[954]), .B(x[954]), .Z(n5135) );
  XNOR U7383 ( .A(n5134), .B(n5128), .Z(n7202) );
  XNOR U7384 ( .A(y[948]), .B(x[948]), .Z(n5128) );
  XNOR U7385 ( .A(n7203), .B(n5133), .Z(n5134) );
  XNOR U7386 ( .A(y[952]), .B(x[952]), .Z(n5133) );
  XNOR U7387 ( .A(y[953]), .B(x[953]), .Z(n7203) );
  XOR U7388 ( .A(n5138), .B(n5137), .Z(n5132) );
  XNOR U7389 ( .A(n7204), .B(n5136), .Z(n5137) );
  XNOR U7390 ( .A(y[949]), .B(x[949]), .Z(n5136) );
  XNOR U7391 ( .A(y[950]), .B(x[950]), .Z(n7204) );
  XOR U7392 ( .A(y[951]), .B(x[951]), .Z(n5138) );
  XNOR U7393 ( .A(n5147), .B(n5139), .Z(n7201) );
  XNOR U7394 ( .A(y[931]), .B(x[931]), .Z(n5139) );
  XNOR U7395 ( .A(n7205), .B(n5152), .Z(n5147) );
  XNOR U7396 ( .A(n5145), .B(n5144), .Z(n5152) );
  XNOR U7397 ( .A(n7206), .B(n5143), .Z(n5144) );
  XNOR U7398 ( .A(y[956]), .B(x[956]), .Z(n5143) );
  XNOR U7399 ( .A(y[957]), .B(x[957]), .Z(n7206) );
  XNOR U7400 ( .A(y[958]), .B(x[958]), .Z(n5145) );
  XNOR U7401 ( .A(n5151), .B(n5146), .Z(n7205) );
  XNOR U7402 ( .A(y[947]), .B(x[947]), .Z(n5146) );
  XNOR U7403 ( .A(n7207), .B(n5155), .Z(n5151) );
  XNOR U7404 ( .A(y[961]), .B(x[961]), .Z(n5155) );
  XNOR U7405 ( .A(n5154), .B(n5150), .Z(n7207) );
  XNOR U7406 ( .A(y[955]), .B(x[955]), .Z(n5150) );
  XNOR U7407 ( .A(n7208), .B(n5153), .Z(n5154) );
  XNOR U7408 ( .A(y[959]), .B(x[959]), .Z(n5153) );
  XNOR U7409 ( .A(y[960]), .B(x[960]), .Z(n7208) );
  XOR U7410 ( .A(n7209), .B(n5199), .Z(n5182) );
  XNOR U7411 ( .A(n5163), .B(n5162), .Z(n5199) );
  XNOR U7412 ( .A(n7210), .B(n5167), .Z(n5162) );
  XNOR U7413 ( .A(n5160), .B(n5159), .Z(n5167) );
  XNOR U7414 ( .A(n7211), .B(n5158), .Z(n5159) );
  XNOR U7415 ( .A(y[878]), .B(x[878]), .Z(n5158) );
  XNOR U7416 ( .A(y[879]), .B(x[879]), .Z(n7211) );
  XNOR U7417 ( .A(y[880]), .B(x[880]), .Z(n5160) );
  XNOR U7418 ( .A(n5166), .B(n5161), .Z(n7210) );
  XNOR U7419 ( .A(y[869]), .B(x[869]), .Z(n5161) );
  XNOR U7420 ( .A(n7212), .B(n5170), .Z(n5166) );
  XNOR U7421 ( .A(y[883]), .B(x[883]), .Z(n5170) );
  XNOR U7422 ( .A(n5169), .B(n5165), .Z(n7212) );
  XNOR U7423 ( .A(y[877]), .B(x[877]), .Z(n5165) );
  XNOR U7424 ( .A(n7213), .B(n5168), .Z(n5169) );
  XNOR U7425 ( .A(y[881]), .B(x[881]), .Z(n5168) );
  XNOR U7426 ( .A(y[882]), .B(x[882]), .Z(n7213) );
  XNOR U7427 ( .A(n5174), .B(n5173), .Z(n5163) );
  XNOR U7428 ( .A(n7214), .B(n5177), .Z(n5173) );
  XNOR U7429 ( .A(y[876]), .B(x[876]), .Z(n5177) );
  XNOR U7430 ( .A(n5176), .B(n5172), .Z(n7214) );
  XNOR U7431 ( .A(y[870]), .B(x[870]), .Z(n5172) );
  XNOR U7432 ( .A(n7215), .B(n5175), .Z(n5176) );
  XNOR U7433 ( .A(y[874]), .B(x[874]), .Z(n5175) );
  XNOR U7434 ( .A(y[875]), .B(x[875]), .Z(n7215) );
  XOR U7435 ( .A(n5180), .B(n5179), .Z(n5174) );
  XNOR U7436 ( .A(n7216), .B(n5178), .Z(n5179) );
  XNOR U7437 ( .A(y[871]), .B(x[871]), .Z(n5178) );
  XNOR U7438 ( .A(y[872]), .B(x[872]), .Z(n7216) );
  XOR U7439 ( .A(y[873]), .B(x[873]), .Z(n5180) );
  XOR U7440 ( .A(n5198), .B(n5181), .Z(n7209) );
  XNOR U7441 ( .A(y[836]), .B(x[836]), .Z(n5181) );
  XOR U7442 ( .A(n7217), .B(n5206), .Z(n5198) );
  XNOR U7443 ( .A(n5190), .B(n5189), .Z(n5206) );
  XNOR U7444 ( .A(n7218), .B(n5193), .Z(n5189) );
  XNOR U7445 ( .A(y[891]), .B(x[891]), .Z(n5193) );
  XNOR U7446 ( .A(n5192), .B(n5186), .Z(n7218) );
  XNOR U7447 ( .A(y[885]), .B(x[885]), .Z(n5186) );
  XNOR U7448 ( .A(n7219), .B(n5191), .Z(n5192) );
  XNOR U7449 ( .A(y[889]), .B(x[889]), .Z(n5191) );
  XNOR U7450 ( .A(y[890]), .B(x[890]), .Z(n7219) );
  XOR U7451 ( .A(n5196), .B(n5195), .Z(n5190) );
  XNOR U7452 ( .A(n7220), .B(n5194), .Z(n5195) );
  XNOR U7453 ( .A(y[886]), .B(x[886]), .Z(n5194) );
  XNOR U7454 ( .A(y[887]), .B(x[887]), .Z(n7220) );
  XOR U7455 ( .A(y[888]), .B(x[888]), .Z(n5196) );
  XNOR U7456 ( .A(n5205), .B(n5197), .Z(n7217) );
  XNOR U7457 ( .A(y[868]), .B(x[868]), .Z(n5197) );
  XNOR U7458 ( .A(n7221), .B(n5210), .Z(n5205) );
  XNOR U7459 ( .A(n5203), .B(n5202), .Z(n5210) );
  XNOR U7460 ( .A(n7222), .B(n5201), .Z(n5202) );
  XNOR U7461 ( .A(y[893]), .B(x[893]), .Z(n5201) );
  XNOR U7462 ( .A(y[894]), .B(x[894]), .Z(n7222) );
  XNOR U7463 ( .A(y[895]), .B(x[895]), .Z(n5203) );
  XNOR U7464 ( .A(n5209), .B(n5204), .Z(n7221) );
  XNOR U7465 ( .A(y[884]), .B(x[884]), .Z(n5204) );
  XNOR U7466 ( .A(n7223), .B(n5213), .Z(n5209) );
  XNOR U7467 ( .A(y[898]), .B(x[898]), .Z(n5213) );
  XNOR U7468 ( .A(n5212), .B(n5208), .Z(n7223) );
  XNOR U7469 ( .A(y[892]), .B(x[892]), .Z(n5208) );
  XNOR U7470 ( .A(n7224), .B(n5211), .Z(n5212) );
  XNOR U7471 ( .A(y[896]), .B(x[896]), .Z(n5211) );
  XNOR U7472 ( .A(y[897]), .B(x[897]), .Z(n7224) );
  XOR U7473 ( .A(n7225), .B(n5234), .Z(n5226) );
  XNOR U7474 ( .A(n5218), .B(n5217), .Z(n5234) );
  XNOR U7475 ( .A(n7226), .B(n5221), .Z(n5217) );
  XNOR U7476 ( .A(y[860]), .B(x[860]), .Z(n5221) );
  XNOR U7477 ( .A(n5220), .B(n5216), .Z(n7226) );
  XNOR U7478 ( .A(y[854]), .B(x[854]), .Z(n5216) );
  XNOR U7479 ( .A(n7227), .B(n5219), .Z(n5220) );
  XNOR U7480 ( .A(y[858]), .B(x[858]), .Z(n5219) );
  XNOR U7481 ( .A(y[859]), .B(x[859]), .Z(n7227) );
  XOR U7482 ( .A(n5224), .B(n5223), .Z(n5218) );
  XNOR U7483 ( .A(n7228), .B(n5222), .Z(n5223) );
  XNOR U7484 ( .A(y[855]), .B(x[855]), .Z(n5222) );
  XNOR U7485 ( .A(y[856]), .B(x[856]), .Z(n7228) );
  XOR U7486 ( .A(y[857]), .B(x[857]), .Z(n5224) );
  XNOR U7487 ( .A(n5233), .B(n5225), .Z(n7225) );
  XNOR U7488 ( .A(y[837]), .B(x[837]), .Z(n5225) );
  XNOR U7489 ( .A(n7229), .B(n5238), .Z(n5233) );
  XNOR U7490 ( .A(n5231), .B(n5230), .Z(n5238) );
  XNOR U7491 ( .A(n7230), .B(n5229), .Z(n5230) );
  XNOR U7492 ( .A(y[862]), .B(x[862]), .Z(n5229) );
  XNOR U7493 ( .A(y[863]), .B(x[863]), .Z(n7230) );
  XNOR U7494 ( .A(y[864]), .B(x[864]), .Z(n5231) );
  XNOR U7495 ( .A(n5237), .B(n5232), .Z(n7229) );
  XNOR U7496 ( .A(y[853]), .B(x[853]), .Z(n5232) );
  XNOR U7497 ( .A(n7231), .B(n5241), .Z(n5237) );
  XNOR U7498 ( .A(y[867]), .B(x[867]), .Z(n5241) );
  XNOR U7499 ( .A(n5240), .B(n5236), .Z(n7231) );
  XNOR U7500 ( .A(y[861]), .B(x[861]), .Z(n5236) );
  XNOR U7501 ( .A(n7232), .B(n5239), .Z(n5240) );
  XNOR U7502 ( .A(y[865]), .B(x[865]), .Z(n5239) );
  XNOR U7503 ( .A(y[866]), .B(x[866]), .Z(n7232) );
  XNOR U7504 ( .A(n5248), .B(n5247), .Z(n5227) );
  XNOR U7505 ( .A(n7233), .B(n5252), .Z(n5247) );
  XNOR U7506 ( .A(n5245), .B(n5244), .Z(n5252) );
  XNOR U7507 ( .A(n7234), .B(n5243), .Z(n5244) );
  XNOR U7508 ( .A(y[847]), .B(x[847]), .Z(n5243) );
  XNOR U7509 ( .A(y[848]), .B(x[848]), .Z(n7234) );
  XNOR U7510 ( .A(y[849]), .B(x[849]), .Z(n5245) );
  XNOR U7511 ( .A(n5251), .B(n5246), .Z(n7233) );
  XNOR U7512 ( .A(y[838]), .B(x[838]), .Z(n5246) );
  XNOR U7513 ( .A(n7235), .B(n5255), .Z(n5251) );
  XNOR U7514 ( .A(y[852]), .B(x[852]), .Z(n5255) );
  XNOR U7515 ( .A(n5254), .B(n5250), .Z(n7235) );
  XNOR U7516 ( .A(y[846]), .B(x[846]), .Z(n5250) );
  XNOR U7517 ( .A(n7236), .B(n5253), .Z(n5254) );
  XNOR U7518 ( .A(y[850]), .B(x[850]), .Z(n5253) );
  XNOR U7519 ( .A(y[851]), .B(x[851]), .Z(n7236) );
  XNOR U7520 ( .A(n5259), .B(n5258), .Z(n5248) );
  XNOR U7521 ( .A(n7237), .B(n5262), .Z(n5258) );
  XNOR U7522 ( .A(y[845]), .B(x[845]), .Z(n5262) );
  XNOR U7523 ( .A(n5261), .B(n5257), .Z(n7237) );
  XNOR U7524 ( .A(y[839]), .B(x[839]), .Z(n5257) );
  XNOR U7525 ( .A(n7238), .B(n5260), .Z(n5261) );
  XNOR U7526 ( .A(y[843]), .B(x[843]), .Z(n5260) );
  XNOR U7527 ( .A(y[844]), .B(x[844]), .Z(n7238) );
  XOR U7528 ( .A(n5265), .B(n5264), .Z(n5259) );
  XNOR U7529 ( .A(n7239), .B(n5263), .Z(n5264) );
  XNOR U7530 ( .A(y[840]), .B(x[840]), .Z(n5263) );
  XNOR U7531 ( .A(y[841]), .B(x[841]), .Z(n7239) );
  XOR U7532 ( .A(y[842]), .B(x[842]), .Z(n5265) );
  XOR U7533 ( .A(n5383), .B(n5266), .Z(n7176) );
  XNOR U7534 ( .A(y[578]), .B(x[578]), .Z(n5266) );
  XOR U7535 ( .A(n7240), .B(n5440), .Z(n5383) );
  XOR U7536 ( .A(n7241), .B(n5315), .Z(n5298) );
  XNOR U7537 ( .A(n5277), .B(n5276), .Z(n5315) );
  XNOR U7538 ( .A(n7242), .B(n5281), .Z(n5276) );
  XNOR U7539 ( .A(n5274), .B(n5273), .Z(n5281) );
  XNOR U7540 ( .A(n7243), .B(n5272), .Z(n5273) );
  XNOR U7541 ( .A(y[1005]), .B(x[1005]), .Z(n5272) );
  XNOR U7542 ( .A(y[1006]), .B(x[1006]), .Z(n7243) );
  XNOR U7543 ( .A(y[1007]), .B(x[1007]), .Z(n5274) );
  XNOR U7544 ( .A(n5280), .B(n5275), .Z(n7242) );
  XNOR U7545 ( .A(y[996]), .B(x[996]), .Z(n5275) );
  XNOR U7546 ( .A(n7244), .B(n5284), .Z(n5280) );
  XNOR U7547 ( .A(y[1010]), .B(x[1010]), .Z(n5284) );
  XNOR U7548 ( .A(n5283), .B(n5279), .Z(n7244) );
  XNOR U7549 ( .A(y[1004]), .B(x[1004]), .Z(n5279) );
  XNOR U7550 ( .A(n7245), .B(n5282), .Z(n5283) );
  XNOR U7551 ( .A(y[1008]), .B(x[1008]), .Z(n5282) );
  XNOR U7552 ( .A(y[1009]), .B(x[1009]), .Z(n7245) );
  XNOR U7553 ( .A(n5290), .B(n5289), .Z(n5277) );
  XNOR U7554 ( .A(n7246), .B(n5293), .Z(n5289) );
  XNOR U7555 ( .A(y[1003]), .B(x[1003]), .Z(n5293) );
  XNOR U7556 ( .A(n5292), .B(n5286), .Z(n7246) );
  XNOR U7557 ( .A(y[997]), .B(x[997]), .Z(n5286) );
  XNOR U7558 ( .A(n7247), .B(n5291), .Z(n5292) );
  XNOR U7559 ( .A(y[1001]), .B(x[1001]), .Z(n5291) );
  XNOR U7560 ( .A(y[1002]), .B(x[1002]), .Z(n7247) );
  XOR U7561 ( .A(n5296), .B(n5295), .Z(n5290) );
  XNOR U7562 ( .A(n7248), .B(n5294), .Z(n5295) );
  XNOR U7563 ( .A(y[998]), .B(x[998]), .Z(n5294) );
  XNOR U7564 ( .A(y[999]), .B(x[999]), .Z(n7248) );
  XOR U7565 ( .A(y[1000]), .B(x[1000]), .Z(n5296) );
  XOR U7566 ( .A(n5314), .B(n5297), .Z(n7241) );
  XNOR U7567 ( .A(y[963]), .B(x[963]), .Z(n5297) );
  XOR U7568 ( .A(n7249), .B(n5322), .Z(n5314) );
  XNOR U7569 ( .A(n5306), .B(n5305), .Z(n5322) );
  XNOR U7570 ( .A(n7250), .B(n5309), .Z(n5305) );
  XNOR U7571 ( .A(y[1018]), .B(x[1018]), .Z(n5309) );
  XNOR U7572 ( .A(n5308), .B(n5302), .Z(n7250) );
  XNOR U7573 ( .A(y[1012]), .B(x[1012]), .Z(n5302) );
  XNOR U7574 ( .A(n7251), .B(n5307), .Z(n5308) );
  XNOR U7575 ( .A(y[1016]), .B(x[1016]), .Z(n5307) );
  XNOR U7576 ( .A(y[1017]), .B(x[1017]), .Z(n7251) );
  XOR U7577 ( .A(n5312), .B(n5311), .Z(n5306) );
  XNOR U7578 ( .A(n7252), .B(n5310), .Z(n5311) );
  XNOR U7579 ( .A(y[1013]), .B(x[1013]), .Z(n5310) );
  XNOR U7580 ( .A(y[1014]), .B(x[1014]), .Z(n7252) );
  XOR U7581 ( .A(y[1015]), .B(x[1015]), .Z(n5312) );
  XNOR U7582 ( .A(n5321), .B(n5313), .Z(n7249) );
  XNOR U7583 ( .A(y[995]), .B(x[995]), .Z(n5313) );
  XNOR U7584 ( .A(n7253), .B(n5326), .Z(n5321) );
  XNOR U7585 ( .A(n5319), .B(n5318), .Z(n5326) );
  XNOR U7586 ( .A(n7254), .B(n5317), .Z(n5318) );
  XNOR U7587 ( .A(y[1020]), .B(x[1020]), .Z(n5317) );
  XNOR U7588 ( .A(y[1021]), .B(x[1021]), .Z(n7254) );
  XNOR U7589 ( .A(y[1022]), .B(x[1022]), .Z(n5319) );
  XNOR U7590 ( .A(n5325), .B(n5320), .Z(n7253) );
  XNOR U7591 ( .A(y[1011]), .B(x[1011]), .Z(n5320) );
  XNOR U7592 ( .A(n7255), .B(n5329), .Z(n5325) );
  XNOR U7593 ( .A(y[1025]), .B(x[1025]), .Z(n5329) );
  XNOR U7594 ( .A(n5328), .B(n5324), .Z(n7255) );
  XNOR U7595 ( .A(y[1019]), .B(x[1019]), .Z(n5324) );
  XNOR U7596 ( .A(n7256), .B(n5327), .Z(n5328) );
  XNOR U7597 ( .A(y[1023]), .B(x[1023]), .Z(n5327) );
  XNOR U7598 ( .A(y[1024]), .B(x[1024]), .Z(n7256) );
  XOR U7599 ( .A(n7257), .B(n5350), .Z(n5342) );
  XNOR U7600 ( .A(n5334), .B(n5333), .Z(n5350) );
  XNOR U7601 ( .A(n7258), .B(n5337), .Z(n5333) );
  XNOR U7602 ( .A(y[987]), .B(x[987]), .Z(n5337) );
  XNOR U7603 ( .A(n5336), .B(n5332), .Z(n7258) );
  XNOR U7604 ( .A(y[981]), .B(x[981]), .Z(n5332) );
  XNOR U7605 ( .A(n7259), .B(n5335), .Z(n5336) );
  XNOR U7606 ( .A(y[985]), .B(x[985]), .Z(n5335) );
  XNOR U7607 ( .A(y[986]), .B(x[986]), .Z(n7259) );
  XOR U7608 ( .A(n5340), .B(n5339), .Z(n5334) );
  XNOR U7609 ( .A(n7260), .B(n5338), .Z(n5339) );
  XNOR U7610 ( .A(y[982]), .B(x[982]), .Z(n5338) );
  XNOR U7611 ( .A(y[983]), .B(x[983]), .Z(n7260) );
  XOR U7612 ( .A(y[984]), .B(x[984]), .Z(n5340) );
  XNOR U7613 ( .A(n5349), .B(n5341), .Z(n7257) );
  XNOR U7614 ( .A(y[964]), .B(x[964]), .Z(n5341) );
  XNOR U7615 ( .A(n7261), .B(n5354), .Z(n5349) );
  XNOR U7616 ( .A(n5347), .B(n5346), .Z(n5354) );
  XNOR U7617 ( .A(n7262), .B(n5345), .Z(n5346) );
  XNOR U7618 ( .A(y[989]), .B(x[989]), .Z(n5345) );
  XNOR U7619 ( .A(y[990]), .B(x[990]), .Z(n7262) );
  XNOR U7620 ( .A(y[991]), .B(x[991]), .Z(n5347) );
  XNOR U7621 ( .A(n5353), .B(n5348), .Z(n7261) );
  XNOR U7622 ( .A(y[980]), .B(x[980]), .Z(n5348) );
  XNOR U7623 ( .A(n7263), .B(n5357), .Z(n5353) );
  XNOR U7624 ( .A(y[994]), .B(x[994]), .Z(n5357) );
  XNOR U7625 ( .A(n5356), .B(n5352), .Z(n7263) );
  XNOR U7626 ( .A(y[988]), .B(x[988]), .Z(n5352) );
  XNOR U7627 ( .A(n7264), .B(n5355), .Z(n5356) );
  XNOR U7628 ( .A(y[992]), .B(x[992]), .Z(n5355) );
  XNOR U7629 ( .A(y[993]), .B(x[993]), .Z(n7264) );
  XNOR U7630 ( .A(n5364), .B(n5363), .Z(n5343) );
  XNOR U7631 ( .A(n7265), .B(n5368), .Z(n5363) );
  XNOR U7632 ( .A(n5361), .B(n5360), .Z(n5368) );
  XNOR U7633 ( .A(n7266), .B(n5359), .Z(n5360) );
  XNOR U7634 ( .A(y[974]), .B(x[974]), .Z(n5359) );
  XNOR U7635 ( .A(y[975]), .B(x[975]), .Z(n7266) );
  XNOR U7636 ( .A(y[976]), .B(x[976]), .Z(n5361) );
  XNOR U7637 ( .A(n5367), .B(n5362), .Z(n7265) );
  XNOR U7638 ( .A(y[965]), .B(x[965]), .Z(n5362) );
  XNOR U7639 ( .A(n7267), .B(n5371), .Z(n5367) );
  XNOR U7640 ( .A(y[979]), .B(x[979]), .Z(n5371) );
  XNOR U7641 ( .A(n5370), .B(n5366), .Z(n7267) );
  XNOR U7642 ( .A(y[973]), .B(x[973]), .Z(n5366) );
  XNOR U7643 ( .A(n7268), .B(n5369), .Z(n5370) );
  XNOR U7644 ( .A(y[977]), .B(x[977]), .Z(n5369) );
  XNOR U7645 ( .A(y[978]), .B(x[978]), .Z(n7268) );
  XNOR U7646 ( .A(n5375), .B(n5374), .Z(n5364) );
  XNOR U7647 ( .A(n7269), .B(n5378), .Z(n5374) );
  XNOR U7648 ( .A(y[972]), .B(x[972]), .Z(n5378) );
  XNOR U7649 ( .A(n5377), .B(n5373), .Z(n7269) );
  XNOR U7650 ( .A(y[966]), .B(x[966]), .Z(n5373) );
  XNOR U7651 ( .A(n7270), .B(n5376), .Z(n5377) );
  XNOR U7652 ( .A(y[970]), .B(x[970]), .Z(n5376) );
  XNOR U7653 ( .A(y[971]), .B(x[971]), .Z(n7270) );
  XOR U7654 ( .A(n5381), .B(n5380), .Z(n5375) );
  XNOR U7655 ( .A(n7271), .B(n5379), .Z(n5380) );
  XNOR U7656 ( .A(y[967]), .B(x[967]), .Z(n5379) );
  XNOR U7657 ( .A(y[968]), .B(x[968]), .Z(n7271) );
  XOR U7658 ( .A(y[969]), .B(x[969]), .Z(n5381) );
  XOR U7659 ( .A(n5439), .B(n5382), .Z(n7240) );
  XNOR U7660 ( .A(y[834]), .B(x[834]), .Z(n5382) );
  XOR U7661 ( .A(n7272), .B(n5468), .Z(n5439) );
  XOR U7662 ( .A(n7273), .B(n5406), .Z(n5398) );
  XNOR U7663 ( .A(n5390), .B(n5389), .Z(n5406) );
  XNOR U7664 ( .A(n7274), .B(n5393), .Z(n5389) );
  XNOR U7665 ( .A(y[1050]), .B(x[1050]), .Z(n5393) );
  XNOR U7666 ( .A(n5392), .B(n5388), .Z(n7274) );
  XNOR U7667 ( .A(y[1044]), .B(x[1044]), .Z(n5388) );
  XNOR U7668 ( .A(n7275), .B(n5391), .Z(n5392) );
  XNOR U7669 ( .A(y[1048]), .B(x[1048]), .Z(n5391) );
  XNOR U7670 ( .A(y[1049]), .B(x[1049]), .Z(n7275) );
  XOR U7671 ( .A(n5396), .B(n5395), .Z(n5390) );
  XNOR U7672 ( .A(n7276), .B(n5394), .Z(n5395) );
  XNOR U7673 ( .A(y[1045]), .B(x[1045]), .Z(n5394) );
  XNOR U7674 ( .A(y[1046]), .B(x[1046]), .Z(n7276) );
  XOR U7675 ( .A(y[1047]), .B(x[1047]), .Z(n5396) );
  XNOR U7676 ( .A(n5405), .B(n5397), .Z(n7273) );
  XNOR U7677 ( .A(y[1027]), .B(x[1027]), .Z(n5397) );
  XNOR U7678 ( .A(n7277), .B(n5410), .Z(n5405) );
  XNOR U7679 ( .A(n5403), .B(n5402), .Z(n5410) );
  XNOR U7680 ( .A(n7278), .B(n5401), .Z(n5402) );
  XNOR U7681 ( .A(y[1052]), .B(x[1052]), .Z(n5401) );
  XNOR U7682 ( .A(y[1053]), .B(x[1053]), .Z(n7278) );
  XNOR U7683 ( .A(y[1054]), .B(x[1054]), .Z(n5403) );
  XNOR U7684 ( .A(n5409), .B(n5404), .Z(n7277) );
  XNOR U7685 ( .A(y[1043]), .B(x[1043]), .Z(n5404) );
  XNOR U7686 ( .A(n7279), .B(n5413), .Z(n5409) );
  XNOR U7687 ( .A(y[1057]), .B(x[1057]), .Z(n5413) );
  XNOR U7688 ( .A(n5412), .B(n5408), .Z(n7279) );
  XNOR U7689 ( .A(y[1051]), .B(x[1051]), .Z(n5408) );
  XNOR U7690 ( .A(n7280), .B(n5411), .Z(n5412) );
  XNOR U7691 ( .A(y[1055]), .B(x[1055]), .Z(n5411) );
  XNOR U7692 ( .A(y[1056]), .B(x[1056]), .Z(n7280) );
  XNOR U7693 ( .A(n5420), .B(n5419), .Z(n5399) );
  XNOR U7694 ( .A(n7281), .B(n5424), .Z(n5419) );
  XNOR U7695 ( .A(n5417), .B(n5416), .Z(n5424) );
  XNOR U7696 ( .A(n7282), .B(n5415), .Z(n5416) );
  XNOR U7697 ( .A(y[1037]), .B(x[1037]), .Z(n5415) );
  XNOR U7698 ( .A(y[1038]), .B(x[1038]), .Z(n7282) );
  XNOR U7699 ( .A(y[1039]), .B(x[1039]), .Z(n5417) );
  XNOR U7700 ( .A(n5423), .B(n5418), .Z(n7281) );
  XNOR U7701 ( .A(y[1028]), .B(x[1028]), .Z(n5418) );
  XNOR U7702 ( .A(n7283), .B(n5427), .Z(n5423) );
  XNOR U7703 ( .A(y[1042]), .B(x[1042]), .Z(n5427) );
  XNOR U7704 ( .A(n5426), .B(n5422), .Z(n7283) );
  XNOR U7705 ( .A(y[1036]), .B(x[1036]), .Z(n5422) );
  XNOR U7706 ( .A(n7284), .B(n5425), .Z(n5426) );
  XNOR U7707 ( .A(y[1040]), .B(x[1040]), .Z(n5425) );
  XNOR U7708 ( .A(y[1041]), .B(x[1041]), .Z(n7284) );
  XNOR U7709 ( .A(n5431), .B(n5430), .Z(n5420) );
  XNOR U7710 ( .A(n7285), .B(n5434), .Z(n5430) );
  XNOR U7711 ( .A(y[1035]), .B(x[1035]), .Z(n5434) );
  XNOR U7712 ( .A(n5433), .B(n5429), .Z(n7285) );
  XNOR U7713 ( .A(y[1029]), .B(x[1029]), .Z(n5429) );
  XNOR U7714 ( .A(n7286), .B(n5432), .Z(n5433) );
  XNOR U7715 ( .A(y[1033]), .B(x[1033]), .Z(n5432) );
  XNOR U7716 ( .A(y[1034]), .B(x[1034]), .Z(n7286) );
  XOR U7717 ( .A(n5437), .B(n5436), .Z(n5431) );
  XNOR U7718 ( .A(n7287), .B(n5435), .Z(n5436) );
  XNOR U7719 ( .A(y[1030]), .B(x[1030]), .Z(n5435) );
  XNOR U7720 ( .A(y[1031]), .B(x[1031]), .Z(n7287) );
  XOR U7721 ( .A(y[1032]), .B(x[1032]), .Z(n5437) );
  XOR U7722 ( .A(n5467), .B(n5438), .Z(n7272) );
  XNOR U7723 ( .A(y[962]), .B(x[962]), .Z(n5438) );
  XOR U7724 ( .A(n7288), .B(n5484), .Z(n5467) );
  XNOR U7725 ( .A(n5448), .B(n5447), .Z(n5484) );
  XNOR U7726 ( .A(n7289), .B(n5452), .Z(n5447) );
  XNOR U7727 ( .A(n5445), .B(n5444), .Z(n5452) );
  XNOR U7728 ( .A(n7290), .B(n5443), .Z(n5444) );
  XNOR U7729 ( .A(y[1068]), .B(x[1068]), .Z(n5443) );
  XNOR U7730 ( .A(y[1069]), .B(x[1069]), .Z(n7290) );
  XNOR U7731 ( .A(y[1070]), .B(x[1070]), .Z(n5445) );
  XNOR U7732 ( .A(n5451), .B(n5446), .Z(n7289) );
  XNOR U7733 ( .A(y[1059]), .B(x[1059]), .Z(n5446) );
  XNOR U7734 ( .A(n7291), .B(n5455), .Z(n5451) );
  XNOR U7735 ( .A(y[1073]), .B(x[1073]), .Z(n5455) );
  XNOR U7736 ( .A(n5454), .B(n5450), .Z(n7291) );
  XNOR U7737 ( .A(y[1067]), .B(x[1067]), .Z(n5450) );
  XNOR U7738 ( .A(n7292), .B(n5453), .Z(n5454) );
  XNOR U7739 ( .A(y[1071]), .B(x[1071]), .Z(n5453) );
  XNOR U7740 ( .A(y[1072]), .B(x[1072]), .Z(n7292) );
  XNOR U7741 ( .A(n5459), .B(n5458), .Z(n5448) );
  XNOR U7742 ( .A(n7293), .B(n5462), .Z(n5458) );
  XNOR U7743 ( .A(y[1066]), .B(x[1066]), .Z(n5462) );
  XNOR U7744 ( .A(n5461), .B(n5457), .Z(n7293) );
  XNOR U7745 ( .A(y[1060]), .B(x[1060]), .Z(n5457) );
  XNOR U7746 ( .A(n7294), .B(n5460), .Z(n5461) );
  XNOR U7747 ( .A(y[1064]), .B(x[1064]), .Z(n5460) );
  XNOR U7748 ( .A(y[1065]), .B(x[1065]), .Z(n7294) );
  XOR U7749 ( .A(n5465), .B(n5464), .Z(n5459) );
  XNOR U7750 ( .A(n7295), .B(n5463), .Z(n5464) );
  XNOR U7751 ( .A(y[1061]), .B(x[1061]), .Z(n5463) );
  XNOR U7752 ( .A(y[1062]), .B(x[1062]), .Z(n7295) );
  XOR U7753 ( .A(y[1063]), .B(x[1063]), .Z(n5465) );
  XOR U7754 ( .A(n5483), .B(n5466), .Z(n7288) );
  XNOR U7755 ( .A(y[1026]), .B(x[1026]), .Z(n5466) );
  XOR U7756 ( .A(n7296), .B(n5491), .Z(n5483) );
  XNOR U7757 ( .A(n5475), .B(n5474), .Z(n5491) );
  XNOR U7758 ( .A(n7297), .B(n5478), .Z(n5474) );
  XNOR U7759 ( .A(y[1081]), .B(x[1081]), .Z(n5478) );
  XNOR U7760 ( .A(n5477), .B(n5471), .Z(n7297) );
  XNOR U7761 ( .A(y[1075]), .B(x[1075]), .Z(n5471) );
  XNOR U7762 ( .A(n7298), .B(n5476), .Z(n5477) );
  XNOR U7763 ( .A(y[1079]), .B(x[1079]), .Z(n5476) );
  XNOR U7764 ( .A(y[1080]), .B(x[1080]), .Z(n7298) );
  XOR U7765 ( .A(n5481), .B(n5480), .Z(n5475) );
  XNOR U7766 ( .A(n7299), .B(n5479), .Z(n5480) );
  XNOR U7767 ( .A(y[1076]), .B(x[1076]), .Z(n5479) );
  XNOR U7768 ( .A(y[1077]), .B(x[1077]), .Z(n7299) );
  XOR U7769 ( .A(y[1078]), .B(x[1078]), .Z(n5481) );
  XNOR U7770 ( .A(n5490), .B(n5482), .Z(n7296) );
  XNOR U7771 ( .A(y[1058]), .B(x[1058]), .Z(n5482) );
  XNOR U7772 ( .A(n7300), .B(n5495), .Z(n5490) );
  XNOR U7773 ( .A(n5488), .B(n5487), .Z(n5495) );
  XNOR U7774 ( .A(n7301), .B(n5486), .Z(n5487) );
  XNOR U7775 ( .A(y[1083]), .B(x[1083]), .Z(n5486) );
  XNOR U7776 ( .A(y[1084]), .B(x[1084]), .Z(n7301) );
  XNOR U7777 ( .A(y[1085]), .B(x[1085]), .Z(n5488) );
  XNOR U7778 ( .A(n5494), .B(n5489), .Z(n7300) );
  XNOR U7779 ( .A(y[1074]), .B(x[1074]), .Z(n5489) );
  XNOR U7780 ( .A(n7302), .B(n5498), .Z(n5494) );
  XNOR U7781 ( .A(y[1088]), .B(x[1088]), .Z(n5498) );
  XNOR U7782 ( .A(n5497), .B(n5493), .Z(n7302) );
  XNOR U7783 ( .A(y[1082]), .B(x[1082]), .Z(n5493) );
  XNOR U7784 ( .A(n7303), .B(n5496), .Z(n5497) );
  XNOR U7785 ( .A(y[1086]), .B(x[1086]), .Z(n5496) );
  XNOR U7786 ( .A(y[1087]), .B(x[1087]), .Z(n7303) );
  XOR U7787 ( .A(n7304), .B(n5672), .Z(n5611) );
  XOR U7788 ( .A(n7305), .B(n5543), .Z(n5526) );
  XNOR U7789 ( .A(n5507), .B(n5506), .Z(n5543) );
  XNOR U7790 ( .A(n7306), .B(n5511), .Z(n5506) );
  XNOR U7791 ( .A(n5504), .B(n5503), .Z(n5511) );
  XNOR U7792 ( .A(n7307), .B(n5502), .Z(n5503) );
  XNOR U7793 ( .A(y[750]), .B(x[750]), .Z(n5502) );
  XNOR U7794 ( .A(y[751]), .B(x[751]), .Z(n7307) );
  XNOR U7795 ( .A(y[752]), .B(x[752]), .Z(n5504) );
  XNOR U7796 ( .A(n5510), .B(n5505), .Z(n7306) );
  XNOR U7797 ( .A(y[741]), .B(x[741]), .Z(n5505) );
  XNOR U7798 ( .A(n7308), .B(n5514), .Z(n5510) );
  XNOR U7799 ( .A(y[755]), .B(x[755]), .Z(n5514) );
  XNOR U7800 ( .A(n5513), .B(n5509), .Z(n7308) );
  XNOR U7801 ( .A(y[749]), .B(x[749]), .Z(n5509) );
  XNOR U7802 ( .A(n7309), .B(n5512), .Z(n5513) );
  XNOR U7803 ( .A(y[753]), .B(x[753]), .Z(n5512) );
  XNOR U7804 ( .A(y[754]), .B(x[754]), .Z(n7309) );
  XNOR U7805 ( .A(n5518), .B(n5517), .Z(n5507) );
  XNOR U7806 ( .A(n7310), .B(n5521), .Z(n5517) );
  XNOR U7807 ( .A(y[748]), .B(x[748]), .Z(n5521) );
  XNOR U7808 ( .A(n5520), .B(n5516), .Z(n7310) );
  XNOR U7809 ( .A(y[742]), .B(x[742]), .Z(n5516) );
  XNOR U7810 ( .A(n7311), .B(n5519), .Z(n5520) );
  XNOR U7811 ( .A(y[746]), .B(x[746]), .Z(n5519) );
  XNOR U7812 ( .A(y[747]), .B(x[747]), .Z(n7311) );
  XOR U7813 ( .A(n5524), .B(n5523), .Z(n5518) );
  XNOR U7814 ( .A(n7312), .B(n5522), .Z(n5523) );
  XNOR U7815 ( .A(y[743]), .B(x[743]), .Z(n5522) );
  XNOR U7816 ( .A(y[744]), .B(x[744]), .Z(n7312) );
  XOR U7817 ( .A(y[745]), .B(x[745]), .Z(n5524) );
  XOR U7818 ( .A(n5542), .B(n5525), .Z(n7305) );
  XNOR U7819 ( .A(y[708]), .B(x[708]), .Z(n5525) );
  XOR U7820 ( .A(n7313), .B(n5550), .Z(n5542) );
  XNOR U7821 ( .A(n5534), .B(n5533), .Z(n5550) );
  XNOR U7822 ( .A(n7314), .B(n5537), .Z(n5533) );
  XNOR U7823 ( .A(y[763]), .B(x[763]), .Z(n5537) );
  XNOR U7824 ( .A(n5536), .B(n5530), .Z(n7314) );
  XNOR U7825 ( .A(y[757]), .B(x[757]), .Z(n5530) );
  XNOR U7826 ( .A(n7315), .B(n5535), .Z(n5536) );
  XNOR U7827 ( .A(y[761]), .B(x[761]), .Z(n5535) );
  XNOR U7828 ( .A(y[762]), .B(x[762]), .Z(n7315) );
  XOR U7829 ( .A(n5540), .B(n5539), .Z(n5534) );
  XNOR U7830 ( .A(n7316), .B(n5538), .Z(n5539) );
  XNOR U7831 ( .A(y[758]), .B(x[758]), .Z(n5538) );
  XNOR U7832 ( .A(y[759]), .B(x[759]), .Z(n7316) );
  XOR U7833 ( .A(y[760]), .B(x[760]), .Z(n5540) );
  XNOR U7834 ( .A(n5549), .B(n5541), .Z(n7313) );
  XNOR U7835 ( .A(y[740]), .B(x[740]), .Z(n5541) );
  XNOR U7836 ( .A(n7317), .B(n5554), .Z(n5549) );
  XNOR U7837 ( .A(n5547), .B(n5546), .Z(n5554) );
  XNOR U7838 ( .A(n7318), .B(n5545), .Z(n5546) );
  XNOR U7839 ( .A(y[765]), .B(x[765]), .Z(n5545) );
  XNOR U7840 ( .A(y[766]), .B(x[766]), .Z(n7318) );
  XNOR U7841 ( .A(y[767]), .B(x[767]), .Z(n5547) );
  XNOR U7842 ( .A(n5553), .B(n5548), .Z(n7317) );
  XNOR U7843 ( .A(y[756]), .B(x[756]), .Z(n5548) );
  XNOR U7844 ( .A(n7319), .B(n5557), .Z(n5553) );
  XNOR U7845 ( .A(y[770]), .B(x[770]), .Z(n5557) );
  XNOR U7846 ( .A(n5556), .B(n5552), .Z(n7319) );
  XNOR U7847 ( .A(y[764]), .B(x[764]), .Z(n5552) );
  XNOR U7848 ( .A(n7320), .B(n5555), .Z(n5556) );
  XNOR U7849 ( .A(y[768]), .B(x[768]), .Z(n5555) );
  XNOR U7850 ( .A(y[769]), .B(x[769]), .Z(n7320) );
  XOR U7851 ( .A(n7321), .B(n5578), .Z(n5570) );
  XNOR U7852 ( .A(n5562), .B(n5561), .Z(n5578) );
  XNOR U7853 ( .A(n7322), .B(n5565), .Z(n5561) );
  XNOR U7854 ( .A(y[732]), .B(x[732]), .Z(n5565) );
  XNOR U7855 ( .A(n5564), .B(n5560), .Z(n7322) );
  XNOR U7856 ( .A(y[726]), .B(x[726]), .Z(n5560) );
  XNOR U7857 ( .A(n7323), .B(n5563), .Z(n5564) );
  XNOR U7858 ( .A(y[730]), .B(x[730]), .Z(n5563) );
  XNOR U7859 ( .A(y[731]), .B(x[731]), .Z(n7323) );
  XOR U7860 ( .A(n5568), .B(n5567), .Z(n5562) );
  XNOR U7861 ( .A(n7324), .B(n5566), .Z(n5567) );
  XNOR U7862 ( .A(y[727]), .B(x[727]), .Z(n5566) );
  XNOR U7863 ( .A(y[728]), .B(x[728]), .Z(n7324) );
  XOR U7864 ( .A(y[729]), .B(x[729]), .Z(n5568) );
  XNOR U7865 ( .A(n5577), .B(n5569), .Z(n7321) );
  XNOR U7866 ( .A(y[709]), .B(x[709]), .Z(n5569) );
  XNOR U7867 ( .A(n7325), .B(n5582), .Z(n5577) );
  XNOR U7868 ( .A(n5575), .B(n5574), .Z(n5582) );
  XNOR U7869 ( .A(n7326), .B(n5573), .Z(n5574) );
  XNOR U7870 ( .A(y[734]), .B(x[734]), .Z(n5573) );
  XNOR U7871 ( .A(y[735]), .B(x[735]), .Z(n7326) );
  XNOR U7872 ( .A(y[736]), .B(x[736]), .Z(n5575) );
  XNOR U7873 ( .A(n5581), .B(n5576), .Z(n7325) );
  XNOR U7874 ( .A(y[725]), .B(x[725]), .Z(n5576) );
  XNOR U7875 ( .A(n7327), .B(n5585), .Z(n5581) );
  XNOR U7876 ( .A(y[739]), .B(x[739]), .Z(n5585) );
  XNOR U7877 ( .A(n5584), .B(n5580), .Z(n7327) );
  XNOR U7878 ( .A(y[733]), .B(x[733]), .Z(n5580) );
  XNOR U7879 ( .A(n7328), .B(n5583), .Z(n5584) );
  XNOR U7880 ( .A(y[737]), .B(x[737]), .Z(n5583) );
  XNOR U7881 ( .A(y[738]), .B(x[738]), .Z(n7328) );
  XNOR U7882 ( .A(n5592), .B(n5591), .Z(n5571) );
  XNOR U7883 ( .A(n7329), .B(n5596), .Z(n5591) );
  XNOR U7884 ( .A(n5589), .B(n5588), .Z(n5596) );
  XNOR U7885 ( .A(n7330), .B(n5587), .Z(n5588) );
  XNOR U7886 ( .A(y[719]), .B(x[719]), .Z(n5587) );
  XNOR U7887 ( .A(y[720]), .B(x[720]), .Z(n7330) );
  XNOR U7888 ( .A(y[721]), .B(x[721]), .Z(n5589) );
  XNOR U7889 ( .A(n5595), .B(n5590), .Z(n7329) );
  XNOR U7890 ( .A(y[710]), .B(x[710]), .Z(n5590) );
  XNOR U7891 ( .A(n7331), .B(n5599), .Z(n5595) );
  XNOR U7892 ( .A(y[724]), .B(x[724]), .Z(n5599) );
  XNOR U7893 ( .A(n5598), .B(n5594), .Z(n7331) );
  XNOR U7894 ( .A(y[718]), .B(x[718]), .Z(n5594) );
  XNOR U7895 ( .A(n7332), .B(n5597), .Z(n5598) );
  XNOR U7896 ( .A(y[722]), .B(x[722]), .Z(n5597) );
  XNOR U7897 ( .A(y[723]), .B(x[723]), .Z(n7332) );
  XNOR U7898 ( .A(n5603), .B(n5602), .Z(n5592) );
  XNOR U7899 ( .A(n7333), .B(n5606), .Z(n5602) );
  XNOR U7900 ( .A(y[717]), .B(x[717]), .Z(n5606) );
  XNOR U7901 ( .A(n5605), .B(n5601), .Z(n7333) );
  XNOR U7902 ( .A(y[711]), .B(x[711]), .Z(n5601) );
  XNOR U7903 ( .A(n7334), .B(n5604), .Z(n5605) );
  XNOR U7904 ( .A(y[715]), .B(x[715]), .Z(n5604) );
  XNOR U7905 ( .A(y[716]), .B(x[716]), .Z(n7334) );
  XOR U7906 ( .A(n5609), .B(n5608), .Z(n5603) );
  XNOR U7907 ( .A(n7335), .B(n5607), .Z(n5608) );
  XNOR U7908 ( .A(y[712]), .B(x[712]), .Z(n5607) );
  XNOR U7909 ( .A(y[713]), .B(x[713]), .Z(n7335) );
  XOR U7910 ( .A(y[714]), .B(x[714]), .Z(n5609) );
  XOR U7911 ( .A(n5671), .B(n5610), .Z(n7304) );
  XNOR U7912 ( .A(y[579]), .B(x[579]), .Z(n5610) );
  XOR U7913 ( .A(n7336), .B(n5702), .Z(n5671) );
  XOR U7914 ( .A(n7337), .B(n5634), .Z(n5626) );
  XNOR U7915 ( .A(n5618), .B(n5617), .Z(n5634) );
  XNOR U7916 ( .A(n7338), .B(n5621), .Z(n5617) );
  XNOR U7917 ( .A(y[795]), .B(x[795]), .Z(n5621) );
  XNOR U7918 ( .A(n5620), .B(n5616), .Z(n7338) );
  XNOR U7919 ( .A(y[789]), .B(x[789]), .Z(n5616) );
  XNOR U7920 ( .A(n7339), .B(n5619), .Z(n5620) );
  XNOR U7921 ( .A(y[793]), .B(x[793]), .Z(n5619) );
  XNOR U7922 ( .A(y[794]), .B(x[794]), .Z(n7339) );
  XOR U7923 ( .A(n5624), .B(n5623), .Z(n5618) );
  XNOR U7924 ( .A(n7340), .B(n5622), .Z(n5623) );
  XNOR U7925 ( .A(y[790]), .B(x[790]), .Z(n5622) );
  XNOR U7926 ( .A(y[791]), .B(x[791]), .Z(n7340) );
  XOR U7927 ( .A(y[792]), .B(x[792]), .Z(n5624) );
  XNOR U7928 ( .A(n5633), .B(n5625), .Z(n7337) );
  XNOR U7929 ( .A(y[772]), .B(x[772]), .Z(n5625) );
  XNOR U7930 ( .A(n7341), .B(n5638), .Z(n5633) );
  XNOR U7931 ( .A(n5631), .B(n5630), .Z(n5638) );
  XNOR U7932 ( .A(n7342), .B(n5629), .Z(n5630) );
  XNOR U7933 ( .A(y[797]), .B(x[797]), .Z(n5629) );
  XNOR U7934 ( .A(y[798]), .B(x[798]), .Z(n7342) );
  XNOR U7935 ( .A(y[799]), .B(x[799]), .Z(n5631) );
  XNOR U7936 ( .A(n5637), .B(n5632), .Z(n7341) );
  XNOR U7937 ( .A(y[788]), .B(x[788]), .Z(n5632) );
  XNOR U7938 ( .A(n7343), .B(n5641), .Z(n5637) );
  XNOR U7939 ( .A(y[802]), .B(x[802]), .Z(n5641) );
  XNOR U7940 ( .A(n5640), .B(n5636), .Z(n7343) );
  XNOR U7941 ( .A(y[796]), .B(x[796]), .Z(n5636) );
  XNOR U7942 ( .A(n7344), .B(n5639), .Z(n5640) );
  XNOR U7943 ( .A(y[800]), .B(x[800]), .Z(n5639) );
  XNOR U7944 ( .A(y[801]), .B(x[801]), .Z(n7344) );
  XNOR U7945 ( .A(n5650), .B(n5649), .Z(n5627) );
  XNOR U7946 ( .A(n7345), .B(n5654), .Z(n5649) );
  XNOR U7947 ( .A(n5645), .B(n5644), .Z(n5654) );
  XNOR U7948 ( .A(n7346), .B(n5643), .Z(n5644) );
  XNOR U7949 ( .A(y[782]), .B(x[782]), .Z(n5643) );
  XNOR U7950 ( .A(y[783]), .B(x[783]), .Z(n7346) );
  XNOR U7951 ( .A(y[784]), .B(x[784]), .Z(n5645) );
  XNOR U7952 ( .A(n5653), .B(n5646), .Z(n7345) );
  XNOR U7953 ( .A(y[773]), .B(x[773]), .Z(n5646) );
  XNOR U7954 ( .A(n7347), .B(n5657), .Z(n5653) );
  XNOR U7955 ( .A(y[787]), .B(x[787]), .Z(n5657) );
  XNOR U7956 ( .A(n5656), .B(n5652), .Z(n7347) );
  XNOR U7957 ( .A(y[781]), .B(x[781]), .Z(n5652) );
  XNOR U7958 ( .A(n7348), .B(n5655), .Z(n5656) );
  XNOR U7959 ( .A(y[785]), .B(x[785]), .Z(n5655) );
  XNOR U7960 ( .A(y[786]), .B(x[786]), .Z(n7348) );
  XNOR U7961 ( .A(n5663), .B(n5662), .Z(n5650) );
  XNOR U7962 ( .A(n7349), .B(n5666), .Z(n5662) );
  XNOR U7963 ( .A(y[780]), .B(x[780]), .Z(n5666) );
  XNOR U7964 ( .A(n5665), .B(n5659), .Z(n7349) );
  XNOR U7965 ( .A(y[774]), .B(x[774]), .Z(n5659) );
  XNOR U7966 ( .A(n7350), .B(n5664), .Z(n5665) );
  XNOR U7967 ( .A(y[778]), .B(x[778]), .Z(n5664) );
  XNOR U7968 ( .A(y[779]), .B(x[779]), .Z(n7350) );
  XOR U7969 ( .A(n5669), .B(n5668), .Z(n5663) );
  XNOR U7970 ( .A(n7351), .B(n5667), .Z(n5668) );
  XNOR U7971 ( .A(y[775]), .B(x[775]), .Z(n5667) );
  XNOR U7972 ( .A(y[776]), .B(x[776]), .Z(n7351) );
  XOR U7973 ( .A(y[777]), .B(x[777]), .Z(n5669) );
  XOR U7974 ( .A(n5701), .B(n5670), .Z(n7336) );
  XNOR U7975 ( .A(y[707]), .B(x[707]), .Z(n5670) );
  XOR U7976 ( .A(n7352), .B(n5718), .Z(n5701) );
  XNOR U7977 ( .A(n5680), .B(n5679), .Z(n5718) );
  XNOR U7978 ( .A(n7353), .B(n5684), .Z(n5679) );
  XNOR U7979 ( .A(n5677), .B(n5676), .Z(n5684) );
  XNOR U7980 ( .A(n7354), .B(n5675), .Z(n5676) );
  XNOR U7981 ( .A(y[813]), .B(x[813]), .Z(n5675) );
  XNOR U7982 ( .A(y[814]), .B(x[814]), .Z(n7354) );
  XNOR U7983 ( .A(y[815]), .B(x[815]), .Z(n5677) );
  XNOR U7984 ( .A(n5683), .B(n5678), .Z(n7353) );
  XNOR U7985 ( .A(y[804]), .B(x[804]), .Z(n5678) );
  XNOR U7986 ( .A(n7355), .B(n5687), .Z(n5683) );
  XNOR U7987 ( .A(y[818]), .B(x[818]), .Z(n5687) );
  XNOR U7988 ( .A(n5686), .B(n5682), .Z(n7355) );
  XNOR U7989 ( .A(y[812]), .B(x[812]), .Z(n5682) );
  XNOR U7990 ( .A(n7356), .B(n5685), .Z(n5686) );
  XNOR U7991 ( .A(y[816]), .B(x[816]), .Z(n5685) );
  XNOR U7992 ( .A(y[817]), .B(x[817]), .Z(n7356) );
  XNOR U7993 ( .A(n5693), .B(n5692), .Z(n5680) );
  XNOR U7994 ( .A(n7357), .B(n5696), .Z(n5692) );
  XNOR U7995 ( .A(y[811]), .B(x[811]), .Z(n5696) );
  XNOR U7996 ( .A(n5695), .B(n5689), .Z(n7357) );
  XNOR U7997 ( .A(y[805]), .B(x[805]), .Z(n5689) );
  XNOR U7998 ( .A(n7358), .B(n5694), .Z(n5695) );
  XNOR U7999 ( .A(y[809]), .B(x[809]), .Z(n5694) );
  XNOR U8000 ( .A(y[810]), .B(x[810]), .Z(n7358) );
  XOR U8001 ( .A(n5699), .B(n5698), .Z(n5693) );
  XNOR U8002 ( .A(n7359), .B(n5697), .Z(n5698) );
  XNOR U8003 ( .A(y[806]), .B(x[806]), .Z(n5697) );
  XNOR U8004 ( .A(y[807]), .B(x[807]), .Z(n7359) );
  XOR U8005 ( .A(y[808]), .B(x[808]), .Z(n5699) );
  XOR U8006 ( .A(n5717), .B(n5700), .Z(n7352) );
  XNOR U8007 ( .A(y[771]), .B(x[771]), .Z(n5700) );
  XOR U8008 ( .A(n7360), .B(n5725), .Z(n5717) );
  XNOR U8009 ( .A(n5709), .B(n5708), .Z(n5725) );
  XNOR U8010 ( .A(n7361), .B(n5712), .Z(n5708) );
  XNOR U8011 ( .A(y[826]), .B(x[826]), .Z(n5712) );
  XNOR U8012 ( .A(n5711), .B(n5705), .Z(n7361) );
  XNOR U8013 ( .A(y[820]), .B(x[820]), .Z(n5705) );
  XNOR U8014 ( .A(n7362), .B(n5710), .Z(n5711) );
  XNOR U8015 ( .A(y[824]), .B(x[824]), .Z(n5710) );
  XNOR U8016 ( .A(y[825]), .B(x[825]), .Z(n7362) );
  XOR U8017 ( .A(n5715), .B(n5714), .Z(n5709) );
  XNOR U8018 ( .A(n7363), .B(n5713), .Z(n5714) );
  XNOR U8019 ( .A(y[821]), .B(x[821]), .Z(n5713) );
  XNOR U8020 ( .A(y[822]), .B(x[822]), .Z(n7363) );
  XOR U8021 ( .A(y[823]), .B(x[823]), .Z(n5715) );
  XNOR U8022 ( .A(n5724), .B(n5716), .Z(n7360) );
  XNOR U8023 ( .A(y[803]), .B(x[803]), .Z(n5716) );
  XNOR U8024 ( .A(n7364), .B(n5729), .Z(n5724) );
  XNOR U8025 ( .A(n5722), .B(n5721), .Z(n5729) );
  XNOR U8026 ( .A(n7365), .B(n5720), .Z(n5721) );
  XNOR U8027 ( .A(y[828]), .B(x[828]), .Z(n5720) );
  XNOR U8028 ( .A(y[829]), .B(x[829]), .Z(n7365) );
  XNOR U8029 ( .A(y[830]), .B(x[830]), .Z(n5722) );
  XNOR U8030 ( .A(n5728), .B(n5723), .Z(n7364) );
  XNOR U8031 ( .A(y[819]), .B(x[819]), .Z(n5723) );
  XNOR U8032 ( .A(n7366), .B(n5732), .Z(n5728) );
  XNOR U8033 ( .A(y[833]), .B(x[833]), .Z(n5732) );
  XNOR U8034 ( .A(n5731), .B(n5727), .Z(n7366) );
  XNOR U8035 ( .A(y[827]), .B(x[827]), .Z(n5727) );
  XNOR U8036 ( .A(n7367), .B(n5730), .Z(n5731) );
  XNOR U8037 ( .A(y[831]), .B(x[831]), .Z(n5730) );
  XNOR U8038 ( .A(y[832]), .B(x[832]), .Z(n7367) );
  XOR U8039 ( .A(n7368), .B(n5818), .Z(n5787) );
  XOR U8040 ( .A(n7369), .B(n5754), .Z(n5746) );
  XNOR U8041 ( .A(n5738), .B(n5737), .Z(n5754) );
  XNOR U8042 ( .A(n7370), .B(n5741), .Z(n5737) );
  XNOR U8043 ( .A(y[668]), .B(x[668]), .Z(n5741) );
  XNOR U8044 ( .A(n5740), .B(n5736), .Z(n7370) );
  XNOR U8045 ( .A(y[662]), .B(x[662]), .Z(n5736) );
  XNOR U8046 ( .A(n7371), .B(n5739), .Z(n5740) );
  XNOR U8047 ( .A(y[666]), .B(x[666]), .Z(n5739) );
  XNOR U8048 ( .A(y[667]), .B(x[667]), .Z(n7371) );
  XOR U8049 ( .A(n5744), .B(n5743), .Z(n5738) );
  XNOR U8050 ( .A(n7372), .B(n5742), .Z(n5743) );
  XNOR U8051 ( .A(y[663]), .B(x[663]), .Z(n5742) );
  XNOR U8052 ( .A(y[664]), .B(x[664]), .Z(n7372) );
  XOR U8053 ( .A(y[665]), .B(x[665]), .Z(n5744) );
  XNOR U8054 ( .A(n5753), .B(n5745), .Z(n7369) );
  XNOR U8055 ( .A(y[645]), .B(x[645]), .Z(n5745) );
  XNOR U8056 ( .A(n7373), .B(n5758), .Z(n5753) );
  XNOR U8057 ( .A(n5751), .B(n5750), .Z(n5758) );
  XNOR U8058 ( .A(n7374), .B(n5749), .Z(n5750) );
  XNOR U8059 ( .A(y[670]), .B(x[670]), .Z(n5749) );
  XNOR U8060 ( .A(y[671]), .B(x[671]), .Z(n7374) );
  XNOR U8061 ( .A(y[672]), .B(x[672]), .Z(n5751) );
  XNOR U8062 ( .A(n5757), .B(n5752), .Z(n7373) );
  XNOR U8063 ( .A(y[661]), .B(x[661]), .Z(n5752) );
  XNOR U8064 ( .A(n7375), .B(n5761), .Z(n5757) );
  XNOR U8065 ( .A(y[675]), .B(x[675]), .Z(n5761) );
  XNOR U8066 ( .A(n5760), .B(n5756), .Z(n7375) );
  XNOR U8067 ( .A(y[669]), .B(x[669]), .Z(n5756) );
  XNOR U8068 ( .A(n7376), .B(n5759), .Z(n5760) );
  XNOR U8069 ( .A(y[673]), .B(x[673]), .Z(n5759) );
  XNOR U8070 ( .A(y[674]), .B(x[674]), .Z(n7376) );
  XNOR U8071 ( .A(n5768), .B(n5767), .Z(n5747) );
  XNOR U8072 ( .A(n7377), .B(n5772), .Z(n5767) );
  XNOR U8073 ( .A(n5765), .B(n5764), .Z(n5772) );
  XNOR U8074 ( .A(n7378), .B(n5763), .Z(n5764) );
  XNOR U8075 ( .A(y[655]), .B(x[655]), .Z(n5763) );
  XNOR U8076 ( .A(y[656]), .B(x[656]), .Z(n7378) );
  XNOR U8077 ( .A(y[657]), .B(x[657]), .Z(n5765) );
  XNOR U8078 ( .A(n5771), .B(n5766), .Z(n7377) );
  XNOR U8079 ( .A(y[646]), .B(x[646]), .Z(n5766) );
  XNOR U8080 ( .A(n7379), .B(n5775), .Z(n5771) );
  XNOR U8081 ( .A(y[660]), .B(x[660]), .Z(n5775) );
  XNOR U8082 ( .A(n5774), .B(n5770), .Z(n7379) );
  XNOR U8083 ( .A(y[654]), .B(x[654]), .Z(n5770) );
  XNOR U8084 ( .A(n7380), .B(n5773), .Z(n5774) );
  XNOR U8085 ( .A(y[658]), .B(x[658]), .Z(n5773) );
  XNOR U8086 ( .A(y[659]), .B(x[659]), .Z(n7380) );
  XNOR U8087 ( .A(n5779), .B(n5778), .Z(n5768) );
  XNOR U8088 ( .A(n7381), .B(n5782), .Z(n5778) );
  XNOR U8089 ( .A(y[653]), .B(x[653]), .Z(n5782) );
  XNOR U8090 ( .A(n5781), .B(n5777), .Z(n7381) );
  XNOR U8091 ( .A(y[647]), .B(x[647]), .Z(n5777) );
  XNOR U8092 ( .A(n7382), .B(n5780), .Z(n5781) );
  XNOR U8093 ( .A(y[651]), .B(x[651]), .Z(n5780) );
  XNOR U8094 ( .A(y[652]), .B(x[652]), .Z(n7382) );
  XOR U8095 ( .A(n5785), .B(n5784), .Z(n5779) );
  XNOR U8096 ( .A(n7383), .B(n5783), .Z(n5784) );
  XNOR U8097 ( .A(y[648]), .B(x[648]), .Z(n5783) );
  XNOR U8098 ( .A(y[649]), .B(x[649]), .Z(n7383) );
  XOR U8099 ( .A(y[650]), .B(x[650]), .Z(n5785) );
  XOR U8100 ( .A(n5817), .B(n5786), .Z(n7368) );
  XNOR U8101 ( .A(y[580]), .B(x[580]), .Z(n5786) );
  XOR U8102 ( .A(n7384), .B(n5834), .Z(n5817) );
  XNOR U8103 ( .A(n5796), .B(n5795), .Z(n5834) );
  XNOR U8104 ( .A(n7385), .B(n5800), .Z(n5795) );
  XNOR U8105 ( .A(n5793), .B(n5792), .Z(n5800) );
  XNOR U8106 ( .A(n7386), .B(n5791), .Z(n5792) );
  XNOR U8107 ( .A(y[686]), .B(x[686]), .Z(n5791) );
  XNOR U8108 ( .A(y[687]), .B(x[687]), .Z(n7386) );
  XNOR U8109 ( .A(y[688]), .B(x[688]), .Z(n5793) );
  XNOR U8110 ( .A(n5799), .B(n5794), .Z(n7385) );
  XNOR U8111 ( .A(y[677]), .B(x[677]), .Z(n5794) );
  XNOR U8112 ( .A(n7387), .B(n5803), .Z(n5799) );
  XNOR U8113 ( .A(y[691]), .B(x[691]), .Z(n5803) );
  XNOR U8114 ( .A(n5802), .B(n5798), .Z(n7387) );
  XNOR U8115 ( .A(y[685]), .B(x[685]), .Z(n5798) );
  XNOR U8116 ( .A(n7388), .B(n5801), .Z(n5802) );
  XNOR U8117 ( .A(y[689]), .B(x[689]), .Z(n5801) );
  XNOR U8118 ( .A(y[690]), .B(x[690]), .Z(n7388) );
  XNOR U8119 ( .A(n5809), .B(n5808), .Z(n5796) );
  XNOR U8120 ( .A(n7389), .B(n5812), .Z(n5808) );
  XNOR U8121 ( .A(y[684]), .B(x[684]), .Z(n5812) );
  XNOR U8122 ( .A(n5811), .B(n5805), .Z(n7389) );
  XNOR U8123 ( .A(y[678]), .B(x[678]), .Z(n5805) );
  XNOR U8124 ( .A(n7390), .B(n5810), .Z(n5811) );
  XNOR U8125 ( .A(y[682]), .B(x[682]), .Z(n5810) );
  XNOR U8126 ( .A(y[683]), .B(x[683]), .Z(n7390) );
  XOR U8127 ( .A(n5815), .B(n5814), .Z(n5809) );
  XNOR U8128 ( .A(n7391), .B(n5813), .Z(n5814) );
  XNOR U8129 ( .A(y[679]), .B(x[679]), .Z(n5813) );
  XNOR U8130 ( .A(y[680]), .B(x[680]), .Z(n7391) );
  XOR U8131 ( .A(y[681]), .B(x[681]), .Z(n5815) );
  XOR U8132 ( .A(n5833), .B(n5816), .Z(n7384) );
  XNOR U8133 ( .A(y[644]), .B(x[644]), .Z(n5816) );
  XOR U8134 ( .A(n7392), .B(n5841), .Z(n5833) );
  XNOR U8135 ( .A(n5825), .B(n5824), .Z(n5841) );
  XNOR U8136 ( .A(n7393), .B(n5828), .Z(n5824) );
  XNOR U8137 ( .A(y[699]), .B(x[699]), .Z(n5828) );
  XNOR U8138 ( .A(n5827), .B(n5821), .Z(n7393) );
  XNOR U8139 ( .A(y[693]), .B(x[693]), .Z(n5821) );
  XNOR U8140 ( .A(n7394), .B(n5826), .Z(n5827) );
  XNOR U8141 ( .A(y[697]), .B(x[697]), .Z(n5826) );
  XNOR U8142 ( .A(y[698]), .B(x[698]), .Z(n7394) );
  XOR U8143 ( .A(n5831), .B(n5830), .Z(n5825) );
  XNOR U8144 ( .A(n7395), .B(n5829), .Z(n5830) );
  XNOR U8145 ( .A(y[694]), .B(x[694]), .Z(n5829) );
  XNOR U8146 ( .A(y[695]), .B(x[695]), .Z(n7395) );
  XOR U8147 ( .A(y[696]), .B(x[696]), .Z(n5831) );
  XNOR U8148 ( .A(n5840), .B(n5832), .Z(n7392) );
  XNOR U8149 ( .A(y[676]), .B(x[676]), .Z(n5832) );
  XNOR U8150 ( .A(n7396), .B(n5845), .Z(n5840) );
  XNOR U8151 ( .A(n5838), .B(n5837), .Z(n5845) );
  XNOR U8152 ( .A(n7397), .B(n5836), .Z(n5837) );
  XNOR U8153 ( .A(y[701]), .B(x[701]), .Z(n5836) );
  XNOR U8154 ( .A(y[702]), .B(x[702]), .Z(n7397) );
  XNOR U8155 ( .A(y[703]), .B(x[703]), .Z(n5838) );
  XNOR U8156 ( .A(n5844), .B(n5839), .Z(n7396) );
  XNOR U8157 ( .A(y[692]), .B(x[692]), .Z(n5839) );
  XNOR U8158 ( .A(n7398), .B(n5848), .Z(n5844) );
  XNOR U8159 ( .A(y[706]), .B(x[706]), .Z(n5848) );
  XNOR U8160 ( .A(n5847), .B(n5843), .Z(n7398) );
  XNOR U8161 ( .A(y[700]), .B(x[700]), .Z(n5843) );
  XNOR U8162 ( .A(n7399), .B(n5846), .Z(n5847) );
  XNOR U8163 ( .A(y[704]), .B(x[704]), .Z(n5846) );
  XNOR U8164 ( .A(y[705]), .B(x[705]), .Z(n7399) );
  XOR U8165 ( .A(n7400), .B(n5894), .Z(n5877) );
  XNOR U8166 ( .A(n5856), .B(n5855), .Z(n5894) );
  XNOR U8167 ( .A(n7401), .B(n5860), .Z(n5855) );
  XNOR U8168 ( .A(n5853), .B(n5852), .Z(n5860) );
  XNOR U8169 ( .A(n7402), .B(n5851), .Z(n5852) );
  XNOR U8170 ( .A(y[623]), .B(x[623]), .Z(n5851) );
  XNOR U8171 ( .A(y[624]), .B(x[624]), .Z(n7402) );
  XNOR U8172 ( .A(y[625]), .B(x[625]), .Z(n5853) );
  XNOR U8173 ( .A(n5859), .B(n5854), .Z(n7401) );
  XNOR U8174 ( .A(y[614]), .B(x[614]), .Z(n5854) );
  XNOR U8175 ( .A(n7403), .B(n5863), .Z(n5859) );
  XNOR U8176 ( .A(y[628]), .B(x[628]), .Z(n5863) );
  XNOR U8177 ( .A(n5862), .B(n5858), .Z(n7403) );
  XNOR U8178 ( .A(y[622]), .B(x[622]), .Z(n5858) );
  XNOR U8179 ( .A(n7404), .B(n5861), .Z(n5862) );
  XNOR U8180 ( .A(y[626]), .B(x[626]), .Z(n5861) );
  XNOR U8181 ( .A(y[627]), .B(x[627]), .Z(n7404) );
  XNOR U8182 ( .A(n5869), .B(n5868), .Z(n5856) );
  XNOR U8183 ( .A(n7405), .B(n5872), .Z(n5868) );
  XNOR U8184 ( .A(y[621]), .B(x[621]), .Z(n5872) );
  XNOR U8185 ( .A(n5871), .B(n5865), .Z(n7405) );
  XNOR U8186 ( .A(y[615]), .B(x[615]), .Z(n5865) );
  XNOR U8187 ( .A(n7406), .B(n5870), .Z(n5871) );
  XNOR U8188 ( .A(y[619]), .B(x[619]), .Z(n5870) );
  XNOR U8189 ( .A(y[620]), .B(x[620]), .Z(n7406) );
  XOR U8190 ( .A(n5875), .B(n5874), .Z(n5869) );
  XNOR U8191 ( .A(n7407), .B(n5873), .Z(n5874) );
  XNOR U8192 ( .A(y[616]), .B(x[616]), .Z(n5873) );
  XNOR U8193 ( .A(y[617]), .B(x[617]), .Z(n7407) );
  XOR U8194 ( .A(y[618]), .B(x[618]), .Z(n5875) );
  XOR U8195 ( .A(n5893), .B(n5876), .Z(n7400) );
  XNOR U8196 ( .A(y[581]), .B(x[581]), .Z(n5876) );
  XOR U8197 ( .A(n7408), .B(n5901), .Z(n5893) );
  XNOR U8198 ( .A(n5885), .B(n5884), .Z(n5901) );
  XNOR U8199 ( .A(n7409), .B(n5888), .Z(n5884) );
  XNOR U8200 ( .A(y[636]), .B(x[636]), .Z(n5888) );
  XNOR U8201 ( .A(n5887), .B(n5881), .Z(n7409) );
  XNOR U8202 ( .A(y[630]), .B(x[630]), .Z(n5881) );
  XNOR U8203 ( .A(n7410), .B(n5886), .Z(n5887) );
  XNOR U8204 ( .A(y[634]), .B(x[634]), .Z(n5886) );
  XNOR U8205 ( .A(y[635]), .B(x[635]), .Z(n7410) );
  XOR U8206 ( .A(n5891), .B(n5890), .Z(n5885) );
  XNOR U8207 ( .A(n7411), .B(n5889), .Z(n5890) );
  XNOR U8208 ( .A(y[631]), .B(x[631]), .Z(n5889) );
  XNOR U8209 ( .A(y[632]), .B(x[632]), .Z(n7411) );
  XOR U8210 ( .A(y[633]), .B(x[633]), .Z(n5891) );
  XNOR U8211 ( .A(n5900), .B(n5892), .Z(n7408) );
  XNOR U8212 ( .A(y[613]), .B(x[613]), .Z(n5892) );
  XNOR U8213 ( .A(n7412), .B(n5905), .Z(n5900) );
  XNOR U8214 ( .A(n5898), .B(n5897), .Z(n5905) );
  XNOR U8215 ( .A(n7413), .B(n5896), .Z(n5897) );
  XNOR U8216 ( .A(y[638]), .B(x[638]), .Z(n5896) );
  XNOR U8217 ( .A(y[639]), .B(x[639]), .Z(n7413) );
  XNOR U8218 ( .A(y[640]), .B(x[640]), .Z(n5898) );
  XNOR U8219 ( .A(n5904), .B(n5899), .Z(n7412) );
  XNOR U8220 ( .A(y[629]), .B(x[629]), .Z(n5899) );
  XNOR U8221 ( .A(n7414), .B(n5908), .Z(n5904) );
  XNOR U8222 ( .A(y[643]), .B(x[643]), .Z(n5908) );
  XNOR U8223 ( .A(n5907), .B(n5903), .Z(n7414) );
  XNOR U8224 ( .A(y[637]), .B(x[637]), .Z(n5903) );
  XNOR U8225 ( .A(n7415), .B(n5906), .Z(n5907) );
  XNOR U8226 ( .A(y[641]), .B(x[641]), .Z(n5906) );
  XNOR U8227 ( .A(y[642]), .B(x[642]), .Z(n7415) );
  XOR U8228 ( .A(n7416), .B(n5929), .Z(n5921) );
  XNOR U8229 ( .A(n5913), .B(n5912), .Z(n5929) );
  XNOR U8230 ( .A(n7417), .B(n5916), .Z(n5912) );
  XNOR U8231 ( .A(y[605]), .B(x[605]), .Z(n5916) );
  XNOR U8232 ( .A(n5915), .B(n5911), .Z(n7417) );
  XNOR U8233 ( .A(y[599]), .B(x[599]), .Z(n5911) );
  XNOR U8234 ( .A(n7418), .B(n5914), .Z(n5915) );
  XNOR U8235 ( .A(y[603]), .B(x[603]), .Z(n5914) );
  XNOR U8236 ( .A(y[604]), .B(x[604]), .Z(n7418) );
  XOR U8237 ( .A(n5919), .B(n5918), .Z(n5913) );
  XNOR U8238 ( .A(n7419), .B(n5917), .Z(n5918) );
  XNOR U8239 ( .A(y[600]), .B(x[600]), .Z(n5917) );
  XNOR U8240 ( .A(y[601]), .B(x[601]), .Z(n7419) );
  XOR U8241 ( .A(y[602]), .B(x[602]), .Z(n5919) );
  XNOR U8242 ( .A(n5928), .B(n5920), .Z(n7416) );
  XNOR U8243 ( .A(y[582]), .B(x[582]), .Z(n5920) );
  XNOR U8244 ( .A(n7420), .B(n5933), .Z(n5928) );
  XNOR U8245 ( .A(n5926), .B(n5925), .Z(n5933) );
  XNOR U8246 ( .A(n7421), .B(n5924), .Z(n5925) );
  XNOR U8247 ( .A(y[607]), .B(x[607]), .Z(n5924) );
  XNOR U8248 ( .A(y[608]), .B(x[608]), .Z(n7421) );
  XNOR U8249 ( .A(y[609]), .B(x[609]), .Z(n5926) );
  XNOR U8250 ( .A(n5932), .B(n5927), .Z(n7420) );
  XNOR U8251 ( .A(y[598]), .B(x[598]), .Z(n5927) );
  XNOR U8252 ( .A(n7422), .B(n5936), .Z(n5932) );
  XNOR U8253 ( .A(y[612]), .B(x[612]), .Z(n5936) );
  XNOR U8254 ( .A(n5935), .B(n5931), .Z(n7422) );
  XNOR U8255 ( .A(y[606]), .B(x[606]), .Z(n5931) );
  XNOR U8256 ( .A(n7423), .B(n5934), .Z(n5935) );
  XNOR U8257 ( .A(y[610]), .B(x[610]), .Z(n5934) );
  XNOR U8258 ( .A(y[611]), .B(x[611]), .Z(n7423) );
  XNOR U8259 ( .A(n5943), .B(n5942), .Z(n5922) );
  XNOR U8260 ( .A(n7424), .B(n5947), .Z(n5942) );
  XNOR U8261 ( .A(n5940), .B(n5939), .Z(n5947) );
  XNOR U8262 ( .A(n7425), .B(n5938), .Z(n5939) );
  XNOR U8263 ( .A(y[592]), .B(x[592]), .Z(n5938) );
  XNOR U8264 ( .A(y[593]), .B(x[593]), .Z(n7425) );
  XNOR U8265 ( .A(y[594]), .B(x[594]), .Z(n5940) );
  XNOR U8266 ( .A(n5946), .B(n5941), .Z(n7424) );
  XNOR U8267 ( .A(y[583]), .B(x[583]), .Z(n5941) );
  XNOR U8268 ( .A(n7426), .B(n5950), .Z(n5946) );
  XNOR U8269 ( .A(y[597]), .B(x[597]), .Z(n5950) );
  XNOR U8270 ( .A(n5949), .B(n5945), .Z(n7426) );
  XNOR U8271 ( .A(y[591]), .B(x[591]), .Z(n5945) );
  XNOR U8272 ( .A(n7427), .B(n5948), .Z(n5949) );
  XNOR U8273 ( .A(y[595]), .B(x[595]), .Z(n5948) );
  XNOR U8274 ( .A(y[596]), .B(x[596]), .Z(n7427) );
  XNOR U8275 ( .A(n5954), .B(n5953), .Z(n5943) );
  XNOR U8276 ( .A(n7428), .B(n5957), .Z(n5953) );
  XNOR U8277 ( .A(y[590]), .B(x[590]), .Z(n5957) );
  XNOR U8278 ( .A(n5956), .B(n5952), .Z(n7428) );
  XNOR U8279 ( .A(y[584]), .B(x[584]), .Z(n5952) );
  XNOR U8280 ( .A(n7429), .B(n5955), .Z(n5956) );
  XNOR U8281 ( .A(y[588]), .B(x[588]), .Z(n5955) );
  XNOR U8282 ( .A(y[589]), .B(x[589]), .Z(n7429) );
  XOR U8283 ( .A(n5960), .B(n5959), .Z(n5954) );
  XNOR U8284 ( .A(n7430), .B(n5958), .Z(n5959) );
  XNOR U8285 ( .A(y[585]), .B(x[585]), .Z(n5958) );
  XNOR U8286 ( .A(y[586]), .B(x[586]), .Z(n7430) );
  XOR U8287 ( .A(y[587]), .B(x[587]), .Z(n5960) );
  XOR U8288 ( .A(n6885), .B(n3017), .Z(n7175) );
  XNOR U8289 ( .A(y[0]), .B(x[0]), .Z(n3017) );
  XOR U8290 ( .A(n7431), .B(n6653), .Z(n6885) );
  XOR U8291 ( .A(n7432), .B(n6135), .Z(n6074) );
  XOR U8292 ( .A(n7433), .B(n6006), .Z(n5989) );
  XNOR U8293 ( .A(n5970), .B(n5969), .Z(n6006) );
  XNOR U8294 ( .A(n7434), .B(n5974), .Z(n5969) );
  XNOR U8295 ( .A(n5967), .B(n5966), .Z(n5974) );
  XNOR U8296 ( .A(n7435), .B(n5965), .Z(n5966) );
  XNOR U8297 ( .A(y[1261]), .B(x[1261]), .Z(n5965) );
  XNOR U8298 ( .A(y[1262]), .B(x[1262]), .Z(n7435) );
  XNOR U8299 ( .A(y[1263]), .B(x[1263]), .Z(n5967) );
  XNOR U8300 ( .A(n5973), .B(n5968), .Z(n7434) );
  XNOR U8301 ( .A(y[1252]), .B(x[1252]), .Z(n5968) );
  XNOR U8302 ( .A(n7436), .B(n5977), .Z(n5973) );
  XNOR U8303 ( .A(y[1266]), .B(x[1266]), .Z(n5977) );
  XNOR U8304 ( .A(n5976), .B(n5972), .Z(n7436) );
  XNOR U8305 ( .A(y[1260]), .B(x[1260]), .Z(n5972) );
  XNOR U8306 ( .A(n7437), .B(n5975), .Z(n5976) );
  XNOR U8307 ( .A(y[1264]), .B(x[1264]), .Z(n5975) );
  XNOR U8308 ( .A(y[1265]), .B(x[1265]), .Z(n7437) );
  XNOR U8309 ( .A(n5981), .B(n5980), .Z(n5970) );
  XNOR U8310 ( .A(n7438), .B(n5984), .Z(n5980) );
  XNOR U8311 ( .A(y[1259]), .B(x[1259]), .Z(n5984) );
  XNOR U8312 ( .A(n5983), .B(n5979), .Z(n7438) );
  XNOR U8313 ( .A(y[1253]), .B(x[1253]), .Z(n5979) );
  XNOR U8314 ( .A(n7439), .B(n5982), .Z(n5983) );
  XNOR U8315 ( .A(y[1257]), .B(x[1257]), .Z(n5982) );
  XNOR U8316 ( .A(y[1258]), .B(x[1258]), .Z(n7439) );
  XOR U8317 ( .A(n5987), .B(n5986), .Z(n5981) );
  XNOR U8318 ( .A(n7440), .B(n5985), .Z(n5986) );
  XNOR U8319 ( .A(y[1254]), .B(x[1254]), .Z(n5985) );
  XNOR U8320 ( .A(y[1255]), .B(x[1255]), .Z(n7440) );
  XOR U8321 ( .A(y[1256]), .B(x[1256]), .Z(n5987) );
  XOR U8322 ( .A(n6005), .B(n5988), .Z(n7433) );
  XNOR U8323 ( .A(y[1219]), .B(x[1219]), .Z(n5988) );
  XOR U8324 ( .A(n7441), .B(n6013), .Z(n6005) );
  XNOR U8325 ( .A(n5997), .B(n5996), .Z(n6013) );
  XNOR U8326 ( .A(n7442), .B(n6000), .Z(n5996) );
  XNOR U8327 ( .A(y[1274]), .B(x[1274]), .Z(n6000) );
  XNOR U8328 ( .A(n5999), .B(n5993), .Z(n7442) );
  XNOR U8329 ( .A(y[1268]), .B(x[1268]), .Z(n5993) );
  XNOR U8330 ( .A(n7443), .B(n5998), .Z(n5999) );
  XNOR U8331 ( .A(y[1272]), .B(x[1272]), .Z(n5998) );
  XNOR U8332 ( .A(y[1273]), .B(x[1273]), .Z(n7443) );
  XOR U8333 ( .A(n6003), .B(n6002), .Z(n5997) );
  XNOR U8334 ( .A(n7444), .B(n6001), .Z(n6002) );
  XNOR U8335 ( .A(y[1269]), .B(x[1269]), .Z(n6001) );
  XNOR U8336 ( .A(y[1270]), .B(x[1270]), .Z(n7444) );
  XOR U8337 ( .A(y[1271]), .B(x[1271]), .Z(n6003) );
  XNOR U8338 ( .A(n6012), .B(n6004), .Z(n7441) );
  XNOR U8339 ( .A(y[1251]), .B(x[1251]), .Z(n6004) );
  XNOR U8340 ( .A(n7445), .B(n6017), .Z(n6012) );
  XNOR U8341 ( .A(n6010), .B(n6009), .Z(n6017) );
  XNOR U8342 ( .A(n7446), .B(n6008), .Z(n6009) );
  XNOR U8343 ( .A(y[1276]), .B(x[1276]), .Z(n6008) );
  XNOR U8344 ( .A(y[1277]), .B(x[1277]), .Z(n7446) );
  XNOR U8345 ( .A(y[1278]), .B(x[1278]), .Z(n6010) );
  XNOR U8346 ( .A(n6016), .B(n6011), .Z(n7445) );
  XNOR U8347 ( .A(y[1267]), .B(x[1267]), .Z(n6011) );
  XNOR U8348 ( .A(n7447), .B(n6020), .Z(n6016) );
  XNOR U8349 ( .A(y[1281]), .B(x[1281]), .Z(n6020) );
  XNOR U8350 ( .A(n6019), .B(n6015), .Z(n7447) );
  XNOR U8351 ( .A(y[1275]), .B(x[1275]), .Z(n6015) );
  XNOR U8352 ( .A(n7448), .B(n6018), .Z(n6019) );
  XNOR U8353 ( .A(y[1279]), .B(x[1279]), .Z(n6018) );
  XNOR U8354 ( .A(y[1280]), .B(x[1280]), .Z(n7448) );
  XOR U8355 ( .A(n7449), .B(n6041), .Z(n6033) );
  XNOR U8356 ( .A(n6025), .B(n6024), .Z(n6041) );
  XNOR U8357 ( .A(n7450), .B(n6028), .Z(n6024) );
  XNOR U8358 ( .A(y[1243]), .B(x[1243]), .Z(n6028) );
  XNOR U8359 ( .A(n6027), .B(n6023), .Z(n7450) );
  XNOR U8360 ( .A(y[1237]), .B(x[1237]), .Z(n6023) );
  XNOR U8361 ( .A(n7451), .B(n6026), .Z(n6027) );
  XNOR U8362 ( .A(y[1241]), .B(x[1241]), .Z(n6026) );
  XNOR U8363 ( .A(y[1242]), .B(x[1242]), .Z(n7451) );
  XOR U8364 ( .A(n6031), .B(n6030), .Z(n6025) );
  XNOR U8365 ( .A(n7452), .B(n6029), .Z(n6030) );
  XNOR U8366 ( .A(y[1238]), .B(x[1238]), .Z(n6029) );
  XNOR U8367 ( .A(y[1239]), .B(x[1239]), .Z(n7452) );
  XOR U8368 ( .A(y[1240]), .B(x[1240]), .Z(n6031) );
  XNOR U8369 ( .A(n6040), .B(n6032), .Z(n7449) );
  XNOR U8370 ( .A(y[1220]), .B(x[1220]), .Z(n6032) );
  XNOR U8371 ( .A(n7453), .B(n6045), .Z(n6040) );
  XNOR U8372 ( .A(n6038), .B(n6037), .Z(n6045) );
  XNOR U8373 ( .A(n7454), .B(n6036), .Z(n6037) );
  XNOR U8374 ( .A(y[1245]), .B(x[1245]), .Z(n6036) );
  XNOR U8375 ( .A(y[1246]), .B(x[1246]), .Z(n7454) );
  XNOR U8376 ( .A(y[1247]), .B(x[1247]), .Z(n6038) );
  XNOR U8377 ( .A(n6044), .B(n6039), .Z(n7453) );
  XNOR U8378 ( .A(y[1236]), .B(x[1236]), .Z(n6039) );
  XNOR U8379 ( .A(n7455), .B(n6048), .Z(n6044) );
  XNOR U8380 ( .A(y[1250]), .B(x[1250]), .Z(n6048) );
  XNOR U8381 ( .A(n6047), .B(n6043), .Z(n7455) );
  XNOR U8382 ( .A(y[1244]), .B(x[1244]), .Z(n6043) );
  XNOR U8383 ( .A(n7456), .B(n6046), .Z(n6047) );
  XNOR U8384 ( .A(y[1248]), .B(x[1248]), .Z(n6046) );
  XNOR U8385 ( .A(y[1249]), .B(x[1249]), .Z(n7456) );
  XNOR U8386 ( .A(n6055), .B(n6054), .Z(n6034) );
  XNOR U8387 ( .A(n7457), .B(n6059), .Z(n6054) );
  XNOR U8388 ( .A(n6052), .B(n6051), .Z(n6059) );
  XNOR U8389 ( .A(n7458), .B(n6050), .Z(n6051) );
  XNOR U8390 ( .A(y[1230]), .B(x[1230]), .Z(n6050) );
  XNOR U8391 ( .A(y[1231]), .B(x[1231]), .Z(n7458) );
  XNOR U8392 ( .A(y[1232]), .B(x[1232]), .Z(n6052) );
  XNOR U8393 ( .A(n6058), .B(n6053), .Z(n7457) );
  XNOR U8394 ( .A(y[1221]), .B(x[1221]), .Z(n6053) );
  XNOR U8395 ( .A(n7459), .B(n6062), .Z(n6058) );
  XNOR U8396 ( .A(y[1235]), .B(x[1235]), .Z(n6062) );
  XNOR U8397 ( .A(n6061), .B(n6057), .Z(n7459) );
  XNOR U8398 ( .A(y[1229]), .B(x[1229]), .Z(n6057) );
  XNOR U8399 ( .A(n7460), .B(n6060), .Z(n6061) );
  XNOR U8400 ( .A(y[1233]), .B(x[1233]), .Z(n6060) );
  XNOR U8401 ( .A(y[1234]), .B(x[1234]), .Z(n7460) );
  XNOR U8402 ( .A(n6066), .B(n6065), .Z(n6055) );
  XNOR U8403 ( .A(n7461), .B(n6069), .Z(n6065) );
  XNOR U8404 ( .A(y[1228]), .B(x[1228]), .Z(n6069) );
  XNOR U8405 ( .A(n6068), .B(n6064), .Z(n7461) );
  XNOR U8406 ( .A(y[1222]), .B(x[1222]), .Z(n6064) );
  XNOR U8407 ( .A(n7462), .B(n6067), .Z(n6068) );
  XNOR U8408 ( .A(y[1226]), .B(x[1226]), .Z(n6067) );
  XNOR U8409 ( .A(y[1227]), .B(x[1227]), .Z(n7462) );
  XOR U8410 ( .A(n6072), .B(n6071), .Z(n6066) );
  XNOR U8411 ( .A(n7463), .B(n6070), .Z(n6071) );
  XNOR U8412 ( .A(y[1223]), .B(x[1223]), .Z(n6070) );
  XNOR U8413 ( .A(y[1224]), .B(x[1224]), .Z(n7463) );
  XOR U8414 ( .A(y[1225]), .B(x[1225]), .Z(n6072) );
  XOR U8415 ( .A(n6134), .B(n6073), .Z(n7432) );
  XNOR U8416 ( .A(y[1090]), .B(x[1090]), .Z(n6073) );
  XOR U8417 ( .A(n7464), .B(n6165), .Z(n6134) );
  XOR U8418 ( .A(n7465), .B(n6097), .Z(n6089) );
  XNOR U8419 ( .A(n6081), .B(n6080), .Z(n6097) );
  XNOR U8420 ( .A(n7466), .B(n6084), .Z(n6080) );
  XNOR U8421 ( .A(y[1306]), .B(x[1306]), .Z(n6084) );
  XNOR U8422 ( .A(n6083), .B(n6079), .Z(n7466) );
  XNOR U8423 ( .A(y[1300]), .B(x[1300]), .Z(n6079) );
  XNOR U8424 ( .A(n7467), .B(n6082), .Z(n6083) );
  XNOR U8425 ( .A(y[1304]), .B(x[1304]), .Z(n6082) );
  XNOR U8426 ( .A(y[1305]), .B(x[1305]), .Z(n7467) );
  XOR U8427 ( .A(n6087), .B(n6086), .Z(n6081) );
  XNOR U8428 ( .A(n7468), .B(n6085), .Z(n6086) );
  XNOR U8429 ( .A(y[1301]), .B(x[1301]), .Z(n6085) );
  XNOR U8430 ( .A(y[1302]), .B(x[1302]), .Z(n7468) );
  XOR U8431 ( .A(y[1303]), .B(x[1303]), .Z(n6087) );
  XNOR U8432 ( .A(n6096), .B(n6088), .Z(n7465) );
  XNOR U8433 ( .A(y[1283]), .B(x[1283]), .Z(n6088) );
  XNOR U8434 ( .A(n7469), .B(n6101), .Z(n6096) );
  XNOR U8435 ( .A(n6094), .B(n6093), .Z(n6101) );
  XNOR U8436 ( .A(n7470), .B(n6092), .Z(n6093) );
  XNOR U8437 ( .A(y[1308]), .B(x[1308]), .Z(n6092) );
  XNOR U8438 ( .A(y[1309]), .B(x[1309]), .Z(n7470) );
  XNOR U8439 ( .A(y[1310]), .B(x[1310]), .Z(n6094) );
  XNOR U8440 ( .A(n6100), .B(n6095), .Z(n7469) );
  XNOR U8441 ( .A(y[1299]), .B(x[1299]), .Z(n6095) );
  XNOR U8442 ( .A(n7471), .B(n6104), .Z(n6100) );
  XNOR U8443 ( .A(y[1313]), .B(x[1313]), .Z(n6104) );
  XNOR U8444 ( .A(n6103), .B(n6099), .Z(n7471) );
  XNOR U8445 ( .A(y[1307]), .B(x[1307]), .Z(n6099) );
  XNOR U8446 ( .A(n7472), .B(n6102), .Z(n6103) );
  XNOR U8447 ( .A(y[1311]), .B(x[1311]), .Z(n6102) );
  XNOR U8448 ( .A(y[1312]), .B(x[1312]), .Z(n7472) );
  XNOR U8449 ( .A(n6113), .B(n6112), .Z(n6090) );
  XNOR U8450 ( .A(n7473), .B(n6117), .Z(n6112) );
  XNOR U8451 ( .A(n6108), .B(n6107), .Z(n6117) );
  XNOR U8452 ( .A(n7474), .B(n6106), .Z(n6107) );
  XNOR U8453 ( .A(y[1293]), .B(x[1293]), .Z(n6106) );
  XNOR U8454 ( .A(y[1294]), .B(x[1294]), .Z(n7474) );
  XNOR U8455 ( .A(y[1295]), .B(x[1295]), .Z(n6108) );
  XNOR U8456 ( .A(n6116), .B(n6109), .Z(n7473) );
  XNOR U8457 ( .A(y[1284]), .B(x[1284]), .Z(n6109) );
  XNOR U8458 ( .A(n7475), .B(n6120), .Z(n6116) );
  XNOR U8459 ( .A(y[1298]), .B(x[1298]), .Z(n6120) );
  XNOR U8460 ( .A(n6119), .B(n6115), .Z(n7475) );
  XNOR U8461 ( .A(y[1292]), .B(x[1292]), .Z(n6115) );
  XNOR U8462 ( .A(n7476), .B(n6118), .Z(n6119) );
  XNOR U8463 ( .A(y[1296]), .B(x[1296]), .Z(n6118) );
  XNOR U8464 ( .A(y[1297]), .B(x[1297]), .Z(n7476) );
  XNOR U8465 ( .A(n6126), .B(n6125), .Z(n6113) );
  XNOR U8466 ( .A(n7477), .B(n6129), .Z(n6125) );
  XNOR U8467 ( .A(y[1291]), .B(x[1291]), .Z(n6129) );
  XNOR U8468 ( .A(n6128), .B(n6122), .Z(n7477) );
  XNOR U8469 ( .A(y[1285]), .B(x[1285]), .Z(n6122) );
  XNOR U8470 ( .A(n7478), .B(n6127), .Z(n6128) );
  XNOR U8471 ( .A(y[1289]), .B(x[1289]), .Z(n6127) );
  XNOR U8472 ( .A(y[1290]), .B(x[1290]), .Z(n7478) );
  XOR U8473 ( .A(n6132), .B(n6131), .Z(n6126) );
  XNOR U8474 ( .A(n7479), .B(n6130), .Z(n6131) );
  XNOR U8475 ( .A(y[1286]), .B(x[1286]), .Z(n6130) );
  XNOR U8476 ( .A(y[1287]), .B(x[1287]), .Z(n7479) );
  XOR U8477 ( .A(y[1288]), .B(x[1288]), .Z(n6132) );
  XOR U8478 ( .A(n6164), .B(n6133), .Z(n7464) );
  XNOR U8479 ( .A(y[1218]), .B(x[1218]), .Z(n6133) );
  XOR U8480 ( .A(n7480), .B(n6181), .Z(n6164) );
  XNOR U8481 ( .A(n6143), .B(n6142), .Z(n6181) );
  XNOR U8482 ( .A(n7481), .B(n6147), .Z(n6142) );
  XNOR U8483 ( .A(n6140), .B(n6139), .Z(n6147) );
  XNOR U8484 ( .A(n7482), .B(n6138), .Z(n6139) );
  XNOR U8485 ( .A(y[1324]), .B(x[1324]), .Z(n6138) );
  XNOR U8486 ( .A(y[1325]), .B(x[1325]), .Z(n7482) );
  XNOR U8487 ( .A(y[1326]), .B(x[1326]), .Z(n6140) );
  XNOR U8488 ( .A(n6146), .B(n6141), .Z(n7481) );
  XNOR U8489 ( .A(y[1315]), .B(x[1315]), .Z(n6141) );
  XNOR U8490 ( .A(n7483), .B(n6150), .Z(n6146) );
  XNOR U8491 ( .A(y[1329]), .B(x[1329]), .Z(n6150) );
  XNOR U8492 ( .A(n6149), .B(n6145), .Z(n7483) );
  XNOR U8493 ( .A(y[1323]), .B(x[1323]), .Z(n6145) );
  XNOR U8494 ( .A(n7484), .B(n6148), .Z(n6149) );
  XNOR U8495 ( .A(y[1327]), .B(x[1327]), .Z(n6148) );
  XNOR U8496 ( .A(y[1328]), .B(x[1328]), .Z(n7484) );
  XNOR U8497 ( .A(n6156), .B(n6155), .Z(n6143) );
  XNOR U8498 ( .A(n7485), .B(n6159), .Z(n6155) );
  XNOR U8499 ( .A(y[1322]), .B(x[1322]), .Z(n6159) );
  XNOR U8500 ( .A(n6158), .B(n6152), .Z(n7485) );
  XNOR U8501 ( .A(y[1316]), .B(x[1316]), .Z(n6152) );
  XNOR U8502 ( .A(n7486), .B(n6157), .Z(n6158) );
  XNOR U8503 ( .A(y[1320]), .B(x[1320]), .Z(n6157) );
  XNOR U8504 ( .A(y[1321]), .B(x[1321]), .Z(n7486) );
  XOR U8505 ( .A(n6162), .B(n6161), .Z(n6156) );
  XNOR U8506 ( .A(n7487), .B(n6160), .Z(n6161) );
  XNOR U8507 ( .A(y[1317]), .B(x[1317]), .Z(n6160) );
  XNOR U8508 ( .A(y[1318]), .B(x[1318]), .Z(n7487) );
  XOR U8509 ( .A(y[1319]), .B(x[1319]), .Z(n6162) );
  XOR U8510 ( .A(n6180), .B(n6163), .Z(n7480) );
  XNOR U8511 ( .A(y[1282]), .B(x[1282]), .Z(n6163) );
  XOR U8512 ( .A(n7488), .B(n6188), .Z(n6180) );
  XNOR U8513 ( .A(n6172), .B(n6171), .Z(n6188) );
  XNOR U8514 ( .A(n7489), .B(n6175), .Z(n6171) );
  XNOR U8515 ( .A(y[1337]), .B(x[1337]), .Z(n6175) );
  XNOR U8516 ( .A(n6174), .B(n6168), .Z(n7489) );
  XNOR U8517 ( .A(y[1331]), .B(x[1331]), .Z(n6168) );
  XNOR U8518 ( .A(n7490), .B(n6173), .Z(n6174) );
  XNOR U8519 ( .A(y[1335]), .B(x[1335]), .Z(n6173) );
  XNOR U8520 ( .A(y[1336]), .B(x[1336]), .Z(n7490) );
  XOR U8521 ( .A(n6178), .B(n6177), .Z(n6172) );
  XNOR U8522 ( .A(n7491), .B(n6176), .Z(n6177) );
  XNOR U8523 ( .A(y[1332]), .B(x[1332]), .Z(n6176) );
  XNOR U8524 ( .A(y[1333]), .B(x[1333]), .Z(n7491) );
  XOR U8525 ( .A(y[1334]), .B(x[1334]), .Z(n6178) );
  XNOR U8526 ( .A(n6187), .B(n6179), .Z(n7488) );
  XNOR U8527 ( .A(y[1314]), .B(x[1314]), .Z(n6179) );
  XNOR U8528 ( .A(n7492), .B(n6192), .Z(n6187) );
  XNOR U8529 ( .A(n6185), .B(n6184), .Z(n6192) );
  XNOR U8530 ( .A(n7493), .B(n6183), .Z(n6184) );
  XNOR U8531 ( .A(y[1339]), .B(x[1339]), .Z(n6183) );
  XNOR U8532 ( .A(y[1340]), .B(x[1340]), .Z(n7493) );
  XNOR U8533 ( .A(y[1341]), .B(x[1341]), .Z(n6185) );
  XNOR U8534 ( .A(n6191), .B(n6186), .Z(n7492) );
  XNOR U8535 ( .A(y[1330]), .B(x[1330]), .Z(n6186) );
  XNOR U8536 ( .A(n7494), .B(n6195), .Z(n6191) );
  XNOR U8537 ( .A(y[1344]), .B(x[1344]), .Z(n6195) );
  XNOR U8538 ( .A(n6194), .B(n6190), .Z(n7494) );
  XNOR U8539 ( .A(y[1338]), .B(x[1338]), .Z(n6190) );
  XNOR U8540 ( .A(n7495), .B(n6193), .Z(n6194) );
  XNOR U8541 ( .A(y[1342]), .B(x[1342]), .Z(n6193) );
  XNOR U8542 ( .A(y[1343]), .B(x[1343]), .Z(n7495) );
  XOR U8543 ( .A(n7496), .B(n6281), .Z(n6252) );
  XOR U8544 ( .A(n7497), .B(n6219), .Z(n6211) );
  XNOR U8545 ( .A(n6203), .B(n6202), .Z(n6219) );
  XNOR U8546 ( .A(n7498), .B(n6206), .Z(n6202) );
  XNOR U8547 ( .A(y[1179]), .B(x[1179]), .Z(n6206) );
  XNOR U8548 ( .A(n6205), .B(n6199), .Z(n7498) );
  XNOR U8549 ( .A(y[1173]), .B(x[1173]), .Z(n6199) );
  XNOR U8550 ( .A(n7499), .B(n6204), .Z(n6205) );
  XNOR U8551 ( .A(y[1177]), .B(x[1177]), .Z(n6204) );
  XNOR U8552 ( .A(y[1178]), .B(x[1178]), .Z(n7499) );
  XOR U8553 ( .A(n6209), .B(n6208), .Z(n6203) );
  XNOR U8554 ( .A(n7500), .B(n6207), .Z(n6208) );
  XNOR U8555 ( .A(y[1174]), .B(x[1174]), .Z(n6207) );
  XNOR U8556 ( .A(y[1175]), .B(x[1175]), .Z(n7500) );
  XOR U8557 ( .A(y[1176]), .B(x[1176]), .Z(n6209) );
  XNOR U8558 ( .A(n6218), .B(n6210), .Z(n7497) );
  XNOR U8559 ( .A(y[1156]), .B(x[1156]), .Z(n6210) );
  XNOR U8560 ( .A(n7501), .B(n6223), .Z(n6218) );
  XNOR U8561 ( .A(n6216), .B(n6215), .Z(n6223) );
  XNOR U8562 ( .A(n7502), .B(n6214), .Z(n6215) );
  XNOR U8563 ( .A(y[1181]), .B(x[1181]), .Z(n6214) );
  XNOR U8564 ( .A(y[1182]), .B(x[1182]), .Z(n7502) );
  XNOR U8565 ( .A(y[1183]), .B(x[1183]), .Z(n6216) );
  XNOR U8566 ( .A(n6222), .B(n6217), .Z(n7501) );
  XNOR U8567 ( .A(y[1172]), .B(x[1172]), .Z(n6217) );
  XNOR U8568 ( .A(n7503), .B(n6226), .Z(n6222) );
  XNOR U8569 ( .A(y[1186]), .B(x[1186]), .Z(n6226) );
  XNOR U8570 ( .A(n6225), .B(n6221), .Z(n7503) );
  XNOR U8571 ( .A(y[1180]), .B(x[1180]), .Z(n6221) );
  XNOR U8572 ( .A(n7504), .B(n6224), .Z(n6225) );
  XNOR U8573 ( .A(y[1184]), .B(x[1184]), .Z(n6224) );
  XNOR U8574 ( .A(y[1185]), .B(x[1185]), .Z(n7504) );
  XNOR U8575 ( .A(n6233), .B(n6232), .Z(n6212) );
  XNOR U8576 ( .A(n7505), .B(n6237), .Z(n6232) );
  XNOR U8577 ( .A(n6230), .B(n6229), .Z(n6237) );
  XNOR U8578 ( .A(n7506), .B(n6228), .Z(n6229) );
  XNOR U8579 ( .A(y[1166]), .B(x[1166]), .Z(n6228) );
  XNOR U8580 ( .A(y[1167]), .B(x[1167]), .Z(n7506) );
  XNOR U8581 ( .A(y[1168]), .B(x[1168]), .Z(n6230) );
  XNOR U8582 ( .A(n6236), .B(n6231), .Z(n7505) );
  XNOR U8583 ( .A(y[1157]), .B(x[1157]), .Z(n6231) );
  XNOR U8584 ( .A(n7507), .B(n6240), .Z(n6236) );
  XNOR U8585 ( .A(y[1171]), .B(x[1171]), .Z(n6240) );
  XNOR U8586 ( .A(n6239), .B(n6235), .Z(n7507) );
  XNOR U8587 ( .A(y[1165]), .B(x[1165]), .Z(n6235) );
  XNOR U8588 ( .A(n7508), .B(n6238), .Z(n6239) );
  XNOR U8589 ( .A(y[1169]), .B(x[1169]), .Z(n6238) );
  XNOR U8590 ( .A(y[1170]), .B(x[1170]), .Z(n7508) );
  XNOR U8591 ( .A(n6244), .B(n6243), .Z(n6233) );
  XNOR U8592 ( .A(n7509), .B(n6247), .Z(n6243) );
  XNOR U8593 ( .A(y[1164]), .B(x[1164]), .Z(n6247) );
  XNOR U8594 ( .A(n6246), .B(n6242), .Z(n7509) );
  XNOR U8595 ( .A(y[1158]), .B(x[1158]), .Z(n6242) );
  XNOR U8596 ( .A(n7510), .B(n6245), .Z(n6246) );
  XNOR U8597 ( .A(y[1162]), .B(x[1162]), .Z(n6245) );
  XNOR U8598 ( .A(y[1163]), .B(x[1163]), .Z(n7510) );
  XOR U8599 ( .A(n6250), .B(n6249), .Z(n6244) );
  XNOR U8600 ( .A(n7511), .B(n6248), .Z(n6249) );
  XNOR U8601 ( .A(y[1159]), .B(x[1159]), .Z(n6248) );
  XNOR U8602 ( .A(y[1160]), .B(x[1160]), .Z(n7511) );
  XOR U8603 ( .A(y[1161]), .B(x[1161]), .Z(n6250) );
  XOR U8604 ( .A(n6280), .B(n6251), .Z(n7496) );
  XNOR U8605 ( .A(y[1091]), .B(x[1091]), .Z(n6251) );
  XOR U8606 ( .A(n7512), .B(n6295), .Z(n6280) );
  XNOR U8607 ( .A(n6261), .B(n6260), .Z(n6295) );
  XNOR U8608 ( .A(n7513), .B(n6265), .Z(n6260) );
  XNOR U8609 ( .A(n6258), .B(n6257), .Z(n6265) );
  XNOR U8610 ( .A(n7514), .B(n6256), .Z(n6257) );
  XNOR U8611 ( .A(y[1197]), .B(x[1197]), .Z(n6256) );
  XNOR U8612 ( .A(y[1198]), .B(x[1198]), .Z(n7514) );
  XNOR U8613 ( .A(y[1199]), .B(x[1199]), .Z(n6258) );
  XNOR U8614 ( .A(n6264), .B(n6259), .Z(n7513) );
  XNOR U8615 ( .A(y[1188]), .B(x[1188]), .Z(n6259) );
  XNOR U8616 ( .A(n7515), .B(n6268), .Z(n6264) );
  XNOR U8617 ( .A(y[1202]), .B(x[1202]), .Z(n6268) );
  XNOR U8618 ( .A(n6267), .B(n6263), .Z(n7515) );
  XNOR U8619 ( .A(y[1196]), .B(x[1196]), .Z(n6263) );
  XNOR U8620 ( .A(n7516), .B(n6266), .Z(n6267) );
  XNOR U8621 ( .A(y[1200]), .B(x[1200]), .Z(n6266) );
  XNOR U8622 ( .A(y[1201]), .B(x[1201]), .Z(n7516) );
  XNOR U8623 ( .A(n6272), .B(n6271), .Z(n6261) );
  XNOR U8624 ( .A(n7517), .B(n6275), .Z(n6271) );
  XNOR U8625 ( .A(y[1195]), .B(x[1195]), .Z(n6275) );
  XNOR U8626 ( .A(n6274), .B(n6270), .Z(n7517) );
  XNOR U8627 ( .A(y[1189]), .B(x[1189]), .Z(n6270) );
  XNOR U8628 ( .A(n7518), .B(n6273), .Z(n6274) );
  XNOR U8629 ( .A(y[1193]), .B(x[1193]), .Z(n6273) );
  XNOR U8630 ( .A(y[1194]), .B(x[1194]), .Z(n7518) );
  XOR U8631 ( .A(n6278), .B(n6277), .Z(n6272) );
  XNOR U8632 ( .A(n7519), .B(n6276), .Z(n6277) );
  XNOR U8633 ( .A(y[1190]), .B(x[1190]), .Z(n6276) );
  XNOR U8634 ( .A(y[1191]), .B(x[1191]), .Z(n7519) );
  XOR U8635 ( .A(y[1192]), .B(x[1192]), .Z(n6278) );
  XOR U8636 ( .A(n6294), .B(n6279), .Z(n7512) );
  XNOR U8637 ( .A(y[1155]), .B(x[1155]), .Z(n6279) );
  XOR U8638 ( .A(n7520), .B(n6302), .Z(n6294) );
  XNOR U8639 ( .A(n6286), .B(n6285), .Z(n6302) );
  XNOR U8640 ( .A(n7521), .B(n6289), .Z(n6285) );
  XNOR U8641 ( .A(y[1210]), .B(x[1210]), .Z(n6289) );
  XNOR U8642 ( .A(n6288), .B(n6284), .Z(n7521) );
  XNOR U8643 ( .A(y[1204]), .B(x[1204]), .Z(n6284) );
  XNOR U8644 ( .A(n7522), .B(n6287), .Z(n6288) );
  XNOR U8645 ( .A(y[1208]), .B(x[1208]), .Z(n6287) );
  XNOR U8646 ( .A(y[1209]), .B(x[1209]), .Z(n7522) );
  XOR U8647 ( .A(n6292), .B(n6291), .Z(n6286) );
  XNOR U8648 ( .A(n7523), .B(n6290), .Z(n6291) );
  XNOR U8649 ( .A(y[1205]), .B(x[1205]), .Z(n6290) );
  XNOR U8650 ( .A(y[1206]), .B(x[1206]), .Z(n7523) );
  XOR U8651 ( .A(y[1207]), .B(x[1207]), .Z(n6292) );
  XNOR U8652 ( .A(n6301), .B(n6293), .Z(n7520) );
  XNOR U8653 ( .A(y[1187]), .B(x[1187]), .Z(n6293) );
  XNOR U8654 ( .A(n7524), .B(n6306), .Z(n6301) );
  XNOR U8655 ( .A(n6299), .B(n6298), .Z(n6306) );
  XNOR U8656 ( .A(n7525), .B(n6297), .Z(n6298) );
  XNOR U8657 ( .A(y[1212]), .B(x[1212]), .Z(n6297) );
  XNOR U8658 ( .A(y[1213]), .B(x[1213]), .Z(n7525) );
  XNOR U8659 ( .A(y[1214]), .B(x[1214]), .Z(n6299) );
  XNOR U8660 ( .A(n6305), .B(n6300), .Z(n7524) );
  XNOR U8661 ( .A(y[1203]), .B(x[1203]), .Z(n6300) );
  XNOR U8662 ( .A(n7526), .B(n6309), .Z(n6305) );
  XNOR U8663 ( .A(y[1217]), .B(x[1217]), .Z(n6309) );
  XNOR U8664 ( .A(n6308), .B(n6304), .Z(n7526) );
  XNOR U8665 ( .A(y[1211]), .B(x[1211]), .Z(n6304) );
  XNOR U8666 ( .A(n7527), .B(n6307), .Z(n6308) );
  XNOR U8667 ( .A(y[1215]), .B(x[1215]), .Z(n6307) );
  XNOR U8668 ( .A(y[1216]), .B(x[1216]), .Z(n7527) );
  XOR U8669 ( .A(n7528), .B(n6351), .Z(n6336) );
  XNOR U8670 ( .A(n6317), .B(n6316), .Z(n6351) );
  XNOR U8671 ( .A(n7529), .B(n6321), .Z(n6316) );
  XNOR U8672 ( .A(n6314), .B(n6313), .Z(n6321) );
  XNOR U8673 ( .A(n7530), .B(n6312), .Z(n6313) );
  XNOR U8674 ( .A(y[1134]), .B(x[1134]), .Z(n6312) );
  XNOR U8675 ( .A(y[1135]), .B(x[1135]), .Z(n7530) );
  XNOR U8676 ( .A(y[1136]), .B(x[1136]), .Z(n6314) );
  XNOR U8677 ( .A(n6320), .B(n6315), .Z(n7529) );
  XNOR U8678 ( .A(y[1125]), .B(x[1125]), .Z(n6315) );
  XNOR U8679 ( .A(n7531), .B(n6324), .Z(n6320) );
  XNOR U8680 ( .A(y[1139]), .B(x[1139]), .Z(n6324) );
  XNOR U8681 ( .A(n6323), .B(n6319), .Z(n7531) );
  XNOR U8682 ( .A(y[1133]), .B(x[1133]), .Z(n6319) );
  XNOR U8683 ( .A(n7532), .B(n6322), .Z(n6323) );
  XNOR U8684 ( .A(y[1137]), .B(x[1137]), .Z(n6322) );
  XNOR U8685 ( .A(y[1138]), .B(x[1138]), .Z(n7532) );
  XNOR U8686 ( .A(n6328), .B(n6327), .Z(n6317) );
  XNOR U8687 ( .A(n7533), .B(n6331), .Z(n6327) );
  XNOR U8688 ( .A(y[1132]), .B(x[1132]), .Z(n6331) );
  XNOR U8689 ( .A(n6330), .B(n6326), .Z(n7533) );
  XNOR U8690 ( .A(y[1126]), .B(x[1126]), .Z(n6326) );
  XNOR U8691 ( .A(n7534), .B(n6329), .Z(n6330) );
  XNOR U8692 ( .A(y[1130]), .B(x[1130]), .Z(n6329) );
  XNOR U8693 ( .A(y[1131]), .B(x[1131]), .Z(n7534) );
  XOR U8694 ( .A(n6334), .B(n6333), .Z(n6328) );
  XNOR U8695 ( .A(n7535), .B(n6332), .Z(n6333) );
  XNOR U8696 ( .A(y[1127]), .B(x[1127]), .Z(n6332) );
  XNOR U8697 ( .A(y[1128]), .B(x[1128]), .Z(n7535) );
  XOR U8698 ( .A(y[1129]), .B(x[1129]), .Z(n6334) );
  XOR U8699 ( .A(n6350), .B(n6335), .Z(n7528) );
  XNOR U8700 ( .A(y[1092]), .B(x[1092]), .Z(n6335) );
  XOR U8701 ( .A(n7536), .B(n6358), .Z(n6350) );
  XNOR U8702 ( .A(n6342), .B(n6341), .Z(n6358) );
  XNOR U8703 ( .A(n7537), .B(n6345), .Z(n6341) );
  XNOR U8704 ( .A(y[1147]), .B(x[1147]), .Z(n6345) );
  XNOR U8705 ( .A(n6344), .B(n6340), .Z(n7537) );
  XNOR U8706 ( .A(y[1141]), .B(x[1141]), .Z(n6340) );
  XNOR U8707 ( .A(n7538), .B(n6343), .Z(n6344) );
  XNOR U8708 ( .A(y[1145]), .B(x[1145]), .Z(n6343) );
  XNOR U8709 ( .A(y[1146]), .B(x[1146]), .Z(n7538) );
  XOR U8710 ( .A(n6348), .B(n6347), .Z(n6342) );
  XNOR U8711 ( .A(n7539), .B(n6346), .Z(n6347) );
  XNOR U8712 ( .A(y[1142]), .B(x[1142]), .Z(n6346) );
  XNOR U8713 ( .A(y[1143]), .B(x[1143]), .Z(n7539) );
  XOR U8714 ( .A(y[1144]), .B(x[1144]), .Z(n6348) );
  XNOR U8715 ( .A(n6357), .B(n6349), .Z(n7536) );
  XNOR U8716 ( .A(y[1124]), .B(x[1124]), .Z(n6349) );
  XNOR U8717 ( .A(n7540), .B(n6362), .Z(n6357) );
  XNOR U8718 ( .A(n6355), .B(n6354), .Z(n6362) );
  XNOR U8719 ( .A(n7541), .B(n6353), .Z(n6354) );
  XNOR U8720 ( .A(y[1149]), .B(x[1149]), .Z(n6353) );
  XNOR U8721 ( .A(y[1150]), .B(x[1150]), .Z(n7541) );
  XNOR U8722 ( .A(y[1151]), .B(x[1151]), .Z(n6355) );
  XNOR U8723 ( .A(n6361), .B(n6356), .Z(n7540) );
  XNOR U8724 ( .A(y[1140]), .B(x[1140]), .Z(n6356) );
  XNOR U8725 ( .A(n7542), .B(n6365), .Z(n6361) );
  XNOR U8726 ( .A(y[1154]), .B(x[1154]), .Z(n6365) );
  XNOR U8727 ( .A(n6364), .B(n6360), .Z(n7542) );
  XNOR U8728 ( .A(y[1148]), .B(x[1148]), .Z(n6360) );
  XNOR U8729 ( .A(n7543), .B(n6363), .Z(n6364) );
  XNOR U8730 ( .A(y[1152]), .B(x[1152]), .Z(n6363) );
  XNOR U8731 ( .A(y[1153]), .B(x[1153]), .Z(n7543) );
  XOR U8732 ( .A(n7544), .B(n6386), .Z(n6378) );
  XNOR U8733 ( .A(n6370), .B(n6369), .Z(n6386) );
  XNOR U8734 ( .A(n7545), .B(n6373), .Z(n6369) );
  XNOR U8735 ( .A(y[1116]), .B(x[1116]), .Z(n6373) );
  XNOR U8736 ( .A(n6372), .B(n6368), .Z(n7545) );
  XNOR U8737 ( .A(y[1110]), .B(x[1110]), .Z(n6368) );
  XNOR U8738 ( .A(n7546), .B(n6371), .Z(n6372) );
  XNOR U8739 ( .A(y[1114]), .B(x[1114]), .Z(n6371) );
  XNOR U8740 ( .A(y[1115]), .B(x[1115]), .Z(n7546) );
  XOR U8741 ( .A(n6376), .B(n6375), .Z(n6370) );
  XNOR U8742 ( .A(n7547), .B(n6374), .Z(n6375) );
  XNOR U8743 ( .A(y[1111]), .B(x[1111]), .Z(n6374) );
  XNOR U8744 ( .A(y[1112]), .B(x[1112]), .Z(n7547) );
  XOR U8745 ( .A(y[1113]), .B(x[1113]), .Z(n6376) );
  XNOR U8746 ( .A(n6385), .B(n6377), .Z(n7544) );
  XNOR U8747 ( .A(y[1093]), .B(x[1093]), .Z(n6377) );
  XNOR U8748 ( .A(n7548), .B(n6390), .Z(n6385) );
  XNOR U8749 ( .A(n6383), .B(n6382), .Z(n6390) );
  XNOR U8750 ( .A(n7549), .B(n6381), .Z(n6382) );
  XNOR U8751 ( .A(y[1118]), .B(x[1118]), .Z(n6381) );
  XNOR U8752 ( .A(y[1119]), .B(x[1119]), .Z(n7549) );
  XNOR U8753 ( .A(y[1120]), .B(x[1120]), .Z(n6383) );
  XNOR U8754 ( .A(n6389), .B(n6384), .Z(n7548) );
  XNOR U8755 ( .A(y[1109]), .B(x[1109]), .Z(n6384) );
  XNOR U8756 ( .A(n7550), .B(n6393), .Z(n6389) );
  XNOR U8757 ( .A(y[1123]), .B(x[1123]), .Z(n6393) );
  XNOR U8758 ( .A(n6392), .B(n6388), .Z(n7550) );
  XNOR U8759 ( .A(y[1117]), .B(x[1117]), .Z(n6388) );
  XNOR U8760 ( .A(n7551), .B(n6391), .Z(n6392) );
  XNOR U8761 ( .A(y[1121]), .B(x[1121]), .Z(n6391) );
  XNOR U8762 ( .A(y[1122]), .B(x[1122]), .Z(n7551) );
  XNOR U8763 ( .A(n6400), .B(n6399), .Z(n6379) );
  XNOR U8764 ( .A(n7552), .B(n6404), .Z(n6399) );
  XNOR U8765 ( .A(n6397), .B(n6396), .Z(n6404) );
  XNOR U8766 ( .A(n7553), .B(n6395), .Z(n6396) );
  XNOR U8767 ( .A(y[1103]), .B(x[1103]), .Z(n6395) );
  XNOR U8768 ( .A(y[1104]), .B(x[1104]), .Z(n7553) );
  XNOR U8769 ( .A(y[1105]), .B(x[1105]), .Z(n6397) );
  XNOR U8770 ( .A(n6403), .B(n6398), .Z(n7552) );
  XNOR U8771 ( .A(y[1094]), .B(x[1094]), .Z(n6398) );
  XNOR U8772 ( .A(n7554), .B(n6407), .Z(n6403) );
  XNOR U8773 ( .A(y[1108]), .B(x[1108]), .Z(n6407) );
  XNOR U8774 ( .A(n6406), .B(n6402), .Z(n7554) );
  XNOR U8775 ( .A(y[1102]), .B(x[1102]), .Z(n6402) );
  XNOR U8776 ( .A(n7555), .B(n6405), .Z(n6406) );
  XNOR U8777 ( .A(y[1106]), .B(x[1106]), .Z(n6405) );
  XNOR U8778 ( .A(y[1107]), .B(x[1107]), .Z(n7555) );
  XNOR U8779 ( .A(n6411), .B(n6410), .Z(n6400) );
  XNOR U8780 ( .A(n7556), .B(n6414), .Z(n6410) );
  XNOR U8781 ( .A(y[1101]), .B(x[1101]), .Z(n6414) );
  XNOR U8782 ( .A(n6413), .B(n6409), .Z(n7556) );
  XNOR U8783 ( .A(y[1095]), .B(x[1095]), .Z(n6409) );
  XNOR U8784 ( .A(n7557), .B(n6412), .Z(n6413) );
  XNOR U8785 ( .A(y[1099]), .B(x[1099]), .Z(n6412) );
  XNOR U8786 ( .A(y[1100]), .B(x[1100]), .Z(n7557) );
  XOR U8787 ( .A(n6417), .B(n6416), .Z(n6411) );
  XNOR U8788 ( .A(n7558), .B(n6415), .Z(n6416) );
  XNOR U8789 ( .A(y[1096]), .B(x[1096]), .Z(n6415) );
  XNOR U8790 ( .A(y[1097]), .B(x[1097]), .Z(n7558) );
  XOR U8791 ( .A(y[1098]), .B(x[1098]), .Z(n6417) );
  XOR U8792 ( .A(n6652), .B(n6884), .Z(n7431) );
  XNOR U8793 ( .A(y[577]), .B(x[577]), .Z(n6884) );
  XOR U8794 ( .A(n7559), .B(n6767), .Z(n6652) );
  XOR U8795 ( .A(n7560), .B(n6508), .Z(n6477) );
  XOR U8796 ( .A(n7561), .B(n6442), .Z(n6434) );
  XNOR U8797 ( .A(n6426), .B(n6425), .Z(n6442) );
  XNOR U8798 ( .A(n7562), .B(n6429), .Z(n6425) );
  XNOR U8799 ( .A(y[1434]), .B(x[1434]), .Z(n6429) );
  XNOR U8800 ( .A(n6428), .B(n6422), .Z(n7562) );
  XNOR U8801 ( .A(y[1428]), .B(x[1428]), .Z(n6422) );
  XNOR U8802 ( .A(n7563), .B(n6427), .Z(n6428) );
  XNOR U8803 ( .A(y[1432]), .B(x[1432]), .Z(n6427) );
  XNOR U8804 ( .A(y[1433]), .B(x[1433]), .Z(n7563) );
  XOR U8805 ( .A(n6432), .B(n6431), .Z(n6426) );
  XNOR U8806 ( .A(n7564), .B(n6430), .Z(n6431) );
  XNOR U8807 ( .A(y[1429]), .B(x[1429]), .Z(n6430) );
  XNOR U8808 ( .A(y[1430]), .B(x[1430]), .Z(n7564) );
  XOR U8809 ( .A(y[1431]), .B(x[1431]), .Z(n6432) );
  XNOR U8810 ( .A(n6441), .B(n6433), .Z(n7561) );
  XNOR U8811 ( .A(y[1411]), .B(x[1411]), .Z(n6433) );
  XNOR U8812 ( .A(n7565), .B(n6446), .Z(n6441) );
  XNOR U8813 ( .A(n6439), .B(n6438), .Z(n6446) );
  XNOR U8814 ( .A(n7566), .B(n6437), .Z(n6438) );
  XNOR U8815 ( .A(y[1436]), .B(x[1436]), .Z(n6437) );
  XNOR U8816 ( .A(y[1437]), .B(x[1437]), .Z(n7566) );
  XNOR U8817 ( .A(y[1438]), .B(x[1438]), .Z(n6439) );
  XNOR U8818 ( .A(n6445), .B(n6440), .Z(n7565) );
  XNOR U8819 ( .A(y[1427]), .B(x[1427]), .Z(n6440) );
  XNOR U8820 ( .A(n7567), .B(n6449), .Z(n6445) );
  XNOR U8821 ( .A(y[1441]), .B(x[1441]), .Z(n6449) );
  XNOR U8822 ( .A(n6448), .B(n6444), .Z(n7567) );
  XNOR U8823 ( .A(y[1435]), .B(x[1435]), .Z(n6444) );
  XNOR U8824 ( .A(n7568), .B(n6447), .Z(n6448) );
  XNOR U8825 ( .A(y[1439]), .B(x[1439]), .Z(n6447) );
  XNOR U8826 ( .A(y[1440]), .B(x[1440]), .Z(n7568) );
  XNOR U8827 ( .A(n6456), .B(n6455), .Z(n6435) );
  XNOR U8828 ( .A(n7569), .B(n6460), .Z(n6455) );
  XNOR U8829 ( .A(n6453), .B(n6452), .Z(n6460) );
  XNOR U8830 ( .A(n7570), .B(n6451), .Z(n6452) );
  XNOR U8831 ( .A(y[1421]), .B(x[1421]), .Z(n6451) );
  XNOR U8832 ( .A(y[1422]), .B(x[1422]), .Z(n7570) );
  XNOR U8833 ( .A(y[1423]), .B(x[1423]), .Z(n6453) );
  XNOR U8834 ( .A(n6459), .B(n6454), .Z(n7569) );
  XNOR U8835 ( .A(y[1412]), .B(x[1412]), .Z(n6454) );
  XNOR U8836 ( .A(n7571), .B(n6463), .Z(n6459) );
  XNOR U8837 ( .A(y[1426]), .B(x[1426]), .Z(n6463) );
  XNOR U8838 ( .A(n6462), .B(n6458), .Z(n7571) );
  XNOR U8839 ( .A(y[1420]), .B(x[1420]), .Z(n6458) );
  XNOR U8840 ( .A(n7572), .B(n6461), .Z(n6462) );
  XNOR U8841 ( .A(y[1424]), .B(x[1424]), .Z(n6461) );
  XNOR U8842 ( .A(y[1425]), .B(x[1425]), .Z(n7572) );
  XNOR U8843 ( .A(n6469), .B(n6468), .Z(n6456) );
  XNOR U8844 ( .A(n7573), .B(n6472), .Z(n6468) );
  XNOR U8845 ( .A(y[1419]), .B(x[1419]), .Z(n6472) );
  XNOR U8846 ( .A(n6471), .B(n6465), .Z(n7573) );
  XNOR U8847 ( .A(y[1413]), .B(x[1413]), .Z(n6465) );
  XNOR U8848 ( .A(n7574), .B(n6470), .Z(n6471) );
  XNOR U8849 ( .A(y[1417]), .B(x[1417]), .Z(n6470) );
  XNOR U8850 ( .A(y[1418]), .B(x[1418]), .Z(n7574) );
  XOR U8851 ( .A(n6475), .B(n6474), .Z(n6469) );
  XNOR U8852 ( .A(n7575), .B(n6473), .Z(n6474) );
  XNOR U8853 ( .A(y[1414]), .B(x[1414]), .Z(n6473) );
  XNOR U8854 ( .A(y[1415]), .B(x[1415]), .Z(n7575) );
  XOR U8855 ( .A(y[1416]), .B(x[1416]), .Z(n6475) );
  XOR U8856 ( .A(n6507), .B(n6476), .Z(n7560) );
  XNOR U8857 ( .A(y[1346]), .B(x[1346]), .Z(n6476) );
  XOR U8858 ( .A(n7576), .B(n6524), .Z(n6507) );
  XNOR U8859 ( .A(n6486), .B(n6485), .Z(n6524) );
  XNOR U8860 ( .A(n7577), .B(n6490), .Z(n6485) );
  XNOR U8861 ( .A(n6483), .B(n6482), .Z(n6490) );
  XNOR U8862 ( .A(n7578), .B(n6481), .Z(n6482) );
  XNOR U8863 ( .A(y[1452]), .B(x[1452]), .Z(n6481) );
  XNOR U8864 ( .A(y[1453]), .B(x[1453]), .Z(n7578) );
  XNOR U8865 ( .A(y[1454]), .B(x[1454]), .Z(n6483) );
  XNOR U8866 ( .A(n6489), .B(n6484), .Z(n7577) );
  XNOR U8867 ( .A(y[1443]), .B(x[1443]), .Z(n6484) );
  XNOR U8868 ( .A(n7579), .B(n6493), .Z(n6489) );
  XNOR U8869 ( .A(y[1457]), .B(x[1457]), .Z(n6493) );
  XNOR U8870 ( .A(n6492), .B(n6488), .Z(n7579) );
  XNOR U8871 ( .A(y[1451]), .B(x[1451]), .Z(n6488) );
  XNOR U8872 ( .A(n7580), .B(n6491), .Z(n6492) );
  XNOR U8873 ( .A(y[1455]), .B(x[1455]), .Z(n6491) );
  XNOR U8874 ( .A(y[1456]), .B(x[1456]), .Z(n7580) );
  XNOR U8875 ( .A(n6499), .B(n6498), .Z(n6486) );
  XNOR U8876 ( .A(n7581), .B(n6502), .Z(n6498) );
  XNOR U8877 ( .A(y[1450]), .B(x[1450]), .Z(n6502) );
  XNOR U8878 ( .A(n6501), .B(n6495), .Z(n7581) );
  XNOR U8879 ( .A(y[1444]), .B(x[1444]), .Z(n6495) );
  XNOR U8880 ( .A(n7582), .B(n6500), .Z(n6501) );
  XNOR U8881 ( .A(y[1448]), .B(x[1448]), .Z(n6500) );
  XNOR U8882 ( .A(y[1449]), .B(x[1449]), .Z(n7582) );
  XOR U8883 ( .A(n6505), .B(n6504), .Z(n6499) );
  XNOR U8884 ( .A(n7583), .B(n6503), .Z(n6504) );
  XNOR U8885 ( .A(y[1445]), .B(x[1445]), .Z(n6503) );
  XNOR U8886 ( .A(y[1446]), .B(x[1446]), .Z(n7583) );
  XOR U8887 ( .A(y[1447]), .B(x[1447]), .Z(n6505) );
  XOR U8888 ( .A(n6523), .B(n6506), .Z(n7576) );
  XNOR U8889 ( .A(y[1410]), .B(x[1410]), .Z(n6506) );
  XOR U8890 ( .A(n7584), .B(n6531), .Z(n6523) );
  XNOR U8891 ( .A(n6515), .B(n6514), .Z(n6531) );
  XNOR U8892 ( .A(n7585), .B(n6518), .Z(n6514) );
  XNOR U8893 ( .A(y[1465]), .B(x[1465]), .Z(n6518) );
  XNOR U8894 ( .A(n6517), .B(n6511), .Z(n7585) );
  XNOR U8895 ( .A(y[1459]), .B(x[1459]), .Z(n6511) );
  XNOR U8896 ( .A(n7586), .B(n6516), .Z(n6517) );
  XNOR U8897 ( .A(y[1463]), .B(x[1463]), .Z(n6516) );
  XNOR U8898 ( .A(y[1464]), .B(x[1464]), .Z(n7586) );
  XOR U8899 ( .A(n6521), .B(n6520), .Z(n6515) );
  XNOR U8900 ( .A(n7587), .B(n6519), .Z(n6520) );
  XNOR U8901 ( .A(y[1460]), .B(x[1460]), .Z(n6519) );
  XNOR U8902 ( .A(y[1461]), .B(x[1461]), .Z(n7587) );
  XOR U8903 ( .A(y[1462]), .B(x[1462]), .Z(n6521) );
  XNOR U8904 ( .A(n6530), .B(n6522), .Z(n7584) );
  XNOR U8905 ( .A(y[1442]), .B(x[1442]), .Z(n6522) );
  XNOR U8906 ( .A(n7588), .B(n6535), .Z(n6530) );
  XNOR U8907 ( .A(n6528), .B(n6527), .Z(n6535) );
  XNOR U8908 ( .A(n7589), .B(n6526), .Z(n6527) );
  XNOR U8909 ( .A(y[1467]), .B(x[1467]), .Z(n6526) );
  XNOR U8910 ( .A(y[1468]), .B(x[1468]), .Z(n7589) );
  XNOR U8911 ( .A(y[1469]), .B(x[1469]), .Z(n6528) );
  XNOR U8912 ( .A(n6534), .B(n6529), .Z(n7588) );
  XNOR U8913 ( .A(y[1458]), .B(x[1458]), .Z(n6529) );
  XNOR U8914 ( .A(n7590), .B(n6538), .Z(n6534) );
  XNOR U8915 ( .A(y[1472]), .B(x[1472]), .Z(n6538) );
  XNOR U8916 ( .A(n6537), .B(n6533), .Z(n7590) );
  XNOR U8917 ( .A(y[1466]), .B(x[1466]), .Z(n6533) );
  XNOR U8918 ( .A(n7591), .B(n6536), .Z(n6537) );
  XNOR U8919 ( .A(y[1470]), .B(x[1470]), .Z(n6536) );
  XNOR U8920 ( .A(y[1471]), .B(x[1471]), .Z(n7591) );
  XOR U8921 ( .A(n7592), .B(n6582), .Z(n6567) );
  XNOR U8922 ( .A(n6546), .B(n6545), .Z(n6582) );
  XNOR U8923 ( .A(n7593), .B(n6550), .Z(n6545) );
  XNOR U8924 ( .A(n6543), .B(n6542), .Z(n6550) );
  XNOR U8925 ( .A(n7594), .B(n6541), .Z(n6542) );
  XNOR U8926 ( .A(y[1389]), .B(x[1389]), .Z(n6541) );
  XNOR U8927 ( .A(y[1390]), .B(x[1390]), .Z(n7594) );
  XNOR U8928 ( .A(y[1391]), .B(x[1391]), .Z(n6543) );
  XNOR U8929 ( .A(n6549), .B(n6544), .Z(n7593) );
  XNOR U8930 ( .A(y[1380]), .B(x[1380]), .Z(n6544) );
  XNOR U8931 ( .A(n7595), .B(n6553), .Z(n6549) );
  XNOR U8932 ( .A(y[1394]), .B(x[1394]), .Z(n6553) );
  XNOR U8933 ( .A(n6552), .B(n6548), .Z(n7595) );
  XNOR U8934 ( .A(y[1388]), .B(x[1388]), .Z(n6548) );
  XNOR U8935 ( .A(n7596), .B(n6551), .Z(n6552) );
  XNOR U8936 ( .A(y[1392]), .B(x[1392]), .Z(n6551) );
  XNOR U8937 ( .A(y[1393]), .B(x[1393]), .Z(n7596) );
  XNOR U8938 ( .A(n6559), .B(n6558), .Z(n6546) );
  XNOR U8939 ( .A(n7597), .B(n6562), .Z(n6558) );
  XNOR U8940 ( .A(y[1387]), .B(x[1387]), .Z(n6562) );
  XNOR U8941 ( .A(n6561), .B(n6555), .Z(n7597) );
  XNOR U8942 ( .A(y[1381]), .B(x[1381]), .Z(n6555) );
  XNOR U8943 ( .A(n7598), .B(n6560), .Z(n6561) );
  XNOR U8944 ( .A(y[1385]), .B(x[1385]), .Z(n6560) );
  XNOR U8945 ( .A(y[1386]), .B(x[1386]), .Z(n7598) );
  XOR U8946 ( .A(n6565), .B(n6564), .Z(n6559) );
  XNOR U8947 ( .A(n7599), .B(n6563), .Z(n6564) );
  XNOR U8948 ( .A(y[1382]), .B(x[1382]), .Z(n6563) );
  XNOR U8949 ( .A(y[1383]), .B(x[1383]), .Z(n7599) );
  XOR U8950 ( .A(y[1384]), .B(x[1384]), .Z(n6565) );
  XOR U8951 ( .A(n6581), .B(n6566), .Z(n7592) );
  XNOR U8952 ( .A(y[1347]), .B(x[1347]), .Z(n6566) );
  XOR U8953 ( .A(n7600), .B(n6589), .Z(n6581) );
  XNOR U8954 ( .A(n6573), .B(n6572), .Z(n6589) );
  XNOR U8955 ( .A(n7601), .B(n6576), .Z(n6572) );
  XNOR U8956 ( .A(y[1402]), .B(x[1402]), .Z(n6576) );
  XNOR U8957 ( .A(n6575), .B(n6571), .Z(n7601) );
  XNOR U8958 ( .A(y[1396]), .B(x[1396]), .Z(n6571) );
  XNOR U8959 ( .A(n7602), .B(n6574), .Z(n6575) );
  XNOR U8960 ( .A(y[1400]), .B(x[1400]), .Z(n6574) );
  XNOR U8961 ( .A(y[1401]), .B(x[1401]), .Z(n7602) );
  XOR U8962 ( .A(n6579), .B(n6578), .Z(n6573) );
  XNOR U8963 ( .A(n7603), .B(n6577), .Z(n6578) );
  XNOR U8964 ( .A(y[1397]), .B(x[1397]), .Z(n6577) );
  XNOR U8965 ( .A(y[1398]), .B(x[1398]), .Z(n7603) );
  XOR U8966 ( .A(y[1399]), .B(x[1399]), .Z(n6579) );
  XNOR U8967 ( .A(n6588), .B(n6580), .Z(n7600) );
  XNOR U8968 ( .A(y[1379]), .B(x[1379]), .Z(n6580) );
  XNOR U8969 ( .A(n7604), .B(n6593), .Z(n6588) );
  XNOR U8970 ( .A(n6586), .B(n6585), .Z(n6593) );
  XNOR U8971 ( .A(n7605), .B(n6584), .Z(n6585) );
  XNOR U8972 ( .A(y[1404]), .B(x[1404]), .Z(n6584) );
  XNOR U8973 ( .A(y[1405]), .B(x[1405]), .Z(n7605) );
  XNOR U8974 ( .A(y[1406]), .B(x[1406]), .Z(n6586) );
  XNOR U8975 ( .A(n6592), .B(n6587), .Z(n7604) );
  XNOR U8976 ( .A(y[1395]), .B(x[1395]), .Z(n6587) );
  XNOR U8977 ( .A(n7606), .B(n6596), .Z(n6592) );
  XNOR U8978 ( .A(y[1409]), .B(x[1409]), .Z(n6596) );
  XNOR U8979 ( .A(n6595), .B(n6591), .Z(n7606) );
  XNOR U8980 ( .A(y[1403]), .B(x[1403]), .Z(n6591) );
  XNOR U8981 ( .A(n7607), .B(n6594), .Z(n6595) );
  XNOR U8982 ( .A(y[1407]), .B(x[1407]), .Z(n6594) );
  XNOR U8983 ( .A(y[1408]), .B(x[1408]), .Z(n7607) );
  XOR U8984 ( .A(n7608), .B(n6617), .Z(n6609) );
  XNOR U8985 ( .A(n6601), .B(n6600), .Z(n6617) );
  XNOR U8986 ( .A(n7609), .B(n6604), .Z(n6600) );
  XNOR U8987 ( .A(y[1371]), .B(x[1371]), .Z(n6604) );
  XNOR U8988 ( .A(n6603), .B(n6599), .Z(n7609) );
  XNOR U8989 ( .A(y[1365]), .B(x[1365]), .Z(n6599) );
  XNOR U8990 ( .A(n7610), .B(n6602), .Z(n6603) );
  XNOR U8991 ( .A(y[1369]), .B(x[1369]), .Z(n6602) );
  XNOR U8992 ( .A(y[1370]), .B(x[1370]), .Z(n7610) );
  XOR U8993 ( .A(n6607), .B(n6606), .Z(n6601) );
  XNOR U8994 ( .A(n7611), .B(n6605), .Z(n6606) );
  XNOR U8995 ( .A(y[1366]), .B(x[1366]), .Z(n6605) );
  XNOR U8996 ( .A(y[1367]), .B(x[1367]), .Z(n7611) );
  XOR U8997 ( .A(y[1368]), .B(x[1368]), .Z(n6607) );
  XNOR U8998 ( .A(n6616), .B(n6608), .Z(n7608) );
  XNOR U8999 ( .A(y[1348]), .B(x[1348]), .Z(n6608) );
  XNOR U9000 ( .A(n7612), .B(n6621), .Z(n6616) );
  XNOR U9001 ( .A(n6614), .B(n6613), .Z(n6621) );
  XNOR U9002 ( .A(n7613), .B(n6612), .Z(n6613) );
  XNOR U9003 ( .A(y[1373]), .B(x[1373]), .Z(n6612) );
  XNOR U9004 ( .A(y[1374]), .B(x[1374]), .Z(n7613) );
  XNOR U9005 ( .A(y[1375]), .B(x[1375]), .Z(n6614) );
  XNOR U9006 ( .A(n6620), .B(n6615), .Z(n7612) );
  XNOR U9007 ( .A(y[1364]), .B(x[1364]), .Z(n6615) );
  XNOR U9008 ( .A(n7614), .B(n6624), .Z(n6620) );
  XNOR U9009 ( .A(y[1378]), .B(x[1378]), .Z(n6624) );
  XNOR U9010 ( .A(n6623), .B(n6619), .Z(n7614) );
  XNOR U9011 ( .A(y[1372]), .B(x[1372]), .Z(n6619) );
  XNOR U9012 ( .A(n7615), .B(n6622), .Z(n6623) );
  XNOR U9013 ( .A(y[1376]), .B(x[1376]), .Z(n6622) );
  XNOR U9014 ( .A(y[1377]), .B(x[1377]), .Z(n7615) );
  XNOR U9015 ( .A(n6631), .B(n6630), .Z(n6610) );
  XNOR U9016 ( .A(n7616), .B(n6635), .Z(n6630) );
  XNOR U9017 ( .A(n6628), .B(n6627), .Z(n6635) );
  XNOR U9018 ( .A(n7617), .B(n6626), .Z(n6627) );
  XNOR U9019 ( .A(y[1358]), .B(x[1358]), .Z(n6626) );
  XNOR U9020 ( .A(y[1359]), .B(x[1359]), .Z(n7617) );
  XNOR U9021 ( .A(y[1360]), .B(x[1360]), .Z(n6628) );
  XNOR U9022 ( .A(n6634), .B(n6629), .Z(n7616) );
  XNOR U9023 ( .A(y[1349]), .B(x[1349]), .Z(n6629) );
  XNOR U9024 ( .A(n7618), .B(n6638), .Z(n6634) );
  XNOR U9025 ( .A(y[1363]), .B(x[1363]), .Z(n6638) );
  XNOR U9026 ( .A(n6637), .B(n6633), .Z(n7618) );
  XNOR U9027 ( .A(y[1357]), .B(x[1357]), .Z(n6633) );
  XNOR U9028 ( .A(n7619), .B(n6636), .Z(n6637) );
  XNOR U9029 ( .A(y[1361]), .B(x[1361]), .Z(n6636) );
  XNOR U9030 ( .A(y[1362]), .B(x[1362]), .Z(n7619) );
  XNOR U9031 ( .A(n6644), .B(n6643), .Z(n6631) );
  XNOR U9032 ( .A(n7620), .B(n6647), .Z(n6643) );
  XNOR U9033 ( .A(y[1356]), .B(x[1356]), .Z(n6647) );
  XNOR U9034 ( .A(n6646), .B(n6640), .Z(n7620) );
  XNOR U9035 ( .A(y[1350]), .B(x[1350]), .Z(n6640) );
  XNOR U9036 ( .A(n7621), .B(n6645), .Z(n6646) );
  XNOR U9037 ( .A(y[1354]), .B(x[1354]), .Z(n6645) );
  XNOR U9038 ( .A(y[1355]), .B(x[1355]), .Z(n7621) );
  XOR U9039 ( .A(n6650), .B(n6649), .Z(n6644) );
  XNOR U9040 ( .A(n7622), .B(n6648), .Z(n6649) );
  XNOR U9041 ( .A(y[1351]), .B(x[1351]), .Z(n6648) );
  XNOR U9042 ( .A(y[1352]), .B(x[1352]), .Z(n7622) );
  XOR U9043 ( .A(y[1353]), .B(x[1353]), .Z(n6650) );
  XOR U9044 ( .A(n6766), .B(n6651), .Z(n7559) );
  XNOR U9045 ( .A(y[1089]), .B(x[1089]), .Z(n6651) );
  XOR U9046 ( .A(n7623), .B(n6823), .Z(n6766) );
  XOR U9047 ( .A(n7624), .B(n6698), .Z(n6681) );
  XNOR U9048 ( .A(n6662), .B(n6661), .Z(n6698) );
  XNOR U9049 ( .A(n7625), .B(n6666), .Z(n6661) );
  XNOR U9050 ( .A(n6659), .B(n6658), .Z(n6666) );
  XNOR U9051 ( .A(n7626), .B(n6657), .Z(n6658) );
  XNOR U9052 ( .A(y[1516]), .B(x[1516]), .Z(n6657) );
  XNOR U9053 ( .A(y[1517]), .B(x[1517]), .Z(n7626) );
  XNOR U9054 ( .A(y[1518]), .B(x[1518]), .Z(n6659) );
  XNOR U9055 ( .A(n6665), .B(n6660), .Z(n7625) );
  XNOR U9056 ( .A(y[1507]), .B(x[1507]), .Z(n6660) );
  XNOR U9057 ( .A(n7627), .B(n6669), .Z(n6665) );
  XNOR U9058 ( .A(y[1521]), .B(x[1521]), .Z(n6669) );
  XNOR U9059 ( .A(n6668), .B(n6664), .Z(n7627) );
  XNOR U9060 ( .A(y[1515]), .B(x[1515]), .Z(n6664) );
  XNOR U9061 ( .A(n7628), .B(n6667), .Z(n6668) );
  XNOR U9062 ( .A(y[1519]), .B(x[1519]), .Z(n6667) );
  XNOR U9063 ( .A(y[1520]), .B(x[1520]), .Z(n7628) );
  XNOR U9064 ( .A(n6673), .B(n6672), .Z(n6662) );
  XNOR U9065 ( .A(n7629), .B(n6676), .Z(n6672) );
  XNOR U9066 ( .A(y[1514]), .B(x[1514]), .Z(n6676) );
  XNOR U9067 ( .A(n6675), .B(n6671), .Z(n7629) );
  XNOR U9068 ( .A(y[1508]), .B(x[1508]), .Z(n6671) );
  XNOR U9069 ( .A(n7630), .B(n6674), .Z(n6675) );
  XNOR U9070 ( .A(y[1512]), .B(x[1512]), .Z(n6674) );
  XNOR U9071 ( .A(y[1513]), .B(x[1513]), .Z(n7630) );
  XOR U9072 ( .A(n6679), .B(n6678), .Z(n6673) );
  XNOR U9073 ( .A(n7631), .B(n6677), .Z(n6678) );
  XNOR U9074 ( .A(y[1509]), .B(x[1509]), .Z(n6677) );
  XNOR U9075 ( .A(y[1510]), .B(x[1510]), .Z(n7631) );
  XOR U9076 ( .A(y[1511]), .B(x[1511]), .Z(n6679) );
  XOR U9077 ( .A(n6697), .B(n6680), .Z(n7624) );
  XNOR U9078 ( .A(y[1474]), .B(x[1474]), .Z(n6680) );
  XOR U9079 ( .A(n7632), .B(n6705), .Z(n6697) );
  XNOR U9080 ( .A(n6689), .B(n6688), .Z(n6705) );
  XNOR U9081 ( .A(n7633), .B(n6692), .Z(n6688) );
  XNOR U9082 ( .A(y[1529]), .B(x[1529]), .Z(n6692) );
  XNOR U9083 ( .A(n6691), .B(n6685), .Z(n7633) );
  XNOR U9084 ( .A(y[1523]), .B(x[1523]), .Z(n6685) );
  XNOR U9085 ( .A(n7634), .B(n6690), .Z(n6691) );
  XNOR U9086 ( .A(y[1527]), .B(x[1527]), .Z(n6690) );
  XNOR U9087 ( .A(y[1528]), .B(x[1528]), .Z(n7634) );
  XOR U9088 ( .A(n6695), .B(n6694), .Z(n6689) );
  XNOR U9089 ( .A(n7635), .B(n6693), .Z(n6694) );
  XNOR U9090 ( .A(y[1524]), .B(x[1524]), .Z(n6693) );
  XNOR U9091 ( .A(y[1525]), .B(x[1525]), .Z(n7635) );
  XOR U9092 ( .A(y[1526]), .B(x[1526]), .Z(n6695) );
  XNOR U9093 ( .A(n6704), .B(n6696), .Z(n7632) );
  XNOR U9094 ( .A(y[1506]), .B(x[1506]), .Z(n6696) );
  XNOR U9095 ( .A(n7636), .B(n6709), .Z(n6704) );
  XNOR U9096 ( .A(n6702), .B(n6701), .Z(n6709) );
  XNOR U9097 ( .A(n7637), .B(n6700), .Z(n6701) );
  XNOR U9098 ( .A(y[1531]), .B(x[1531]), .Z(n6700) );
  XNOR U9099 ( .A(y[1532]), .B(x[1532]), .Z(n7637) );
  XNOR U9100 ( .A(y[1533]), .B(x[1533]), .Z(n6702) );
  XNOR U9101 ( .A(n6708), .B(n6703), .Z(n7636) );
  XNOR U9102 ( .A(y[1522]), .B(x[1522]), .Z(n6703) );
  XNOR U9103 ( .A(n7638), .B(n6712), .Z(n6708) );
  XNOR U9104 ( .A(y[1536]), .B(x[1536]), .Z(n6712) );
  XNOR U9105 ( .A(n6711), .B(n6707), .Z(n7638) );
  XNOR U9106 ( .A(y[1530]), .B(x[1530]), .Z(n6707) );
  XNOR U9107 ( .A(n7639), .B(n6710), .Z(n6711) );
  XNOR U9108 ( .A(y[1534]), .B(x[1534]), .Z(n6710) );
  XNOR U9109 ( .A(y[1535]), .B(x[1535]), .Z(n7639) );
  XOR U9110 ( .A(n7640), .B(n6733), .Z(n6725) );
  XNOR U9111 ( .A(n6717), .B(n6716), .Z(n6733) );
  XNOR U9112 ( .A(n7641), .B(n6720), .Z(n6716) );
  XNOR U9113 ( .A(y[1498]), .B(x[1498]), .Z(n6720) );
  XNOR U9114 ( .A(n6719), .B(n6715), .Z(n7641) );
  XNOR U9115 ( .A(y[1492]), .B(x[1492]), .Z(n6715) );
  XNOR U9116 ( .A(n7642), .B(n6718), .Z(n6719) );
  XNOR U9117 ( .A(y[1496]), .B(x[1496]), .Z(n6718) );
  XNOR U9118 ( .A(y[1497]), .B(x[1497]), .Z(n7642) );
  XOR U9119 ( .A(n6723), .B(n6722), .Z(n6717) );
  XNOR U9120 ( .A(n7643), .B(n6721), .Z(n6722) );
  XNOR U9121 ( .A(y[1493]), .B(x[1493]), .Z(n6721) );
  XNOR U9122 ( .A(y[1494]), .B(x[1494]), .Z(n7643) );
  XOR U9123 ( .A(y[1495]), .B(x[1495]), .Z(n6723) );
  XNOR U9124 ( .A(n6732), .B(n6724), .Z(n7640) );
  XNOR U9125 ( .A(y[1475]), .B(x[1475]), .Z(n6724) );
  XNOR U9126 ( .A(n7644), .B(n6737), .Z(n6732) );
  XNOR U9127 ( .A(n6730), .B(n6729), .Z(n6737) );
  XNOR U9128 ( .A(n7645), .B(n6728), .Z(n6729) );
  XNOR U9129 ( .A(y[1500]), .B(x[1500]), .Z(n6728) );
  XNOR U9130 ( .A(y[1501]), .B(x[1501]), .Z(n7645) );
  XNOR U9131 ( .A(y[1502]), .B(x[1502]), .Z(n6730) );
  XNOR U9132 ( .A(n6736), .B(n6731), .Z(n7644) );
  XNOR U9133 ( .A(y[1491]), .B(x[1491]), .Z(n6731) );
  XNOR U9134 ( .A(n7646), .B(n6740), .Z(n6736) );
  XNOR U9135 ( .A(y[1505]), .B(x[1505]), .Z(n6740) );
  XNOR U9136 ( .A(n6739), .B(n6735), .Z(n7646) );
  XNOR U9137 ( .A(y[1499]), .B(x[1499]), .Z(n6735) );
  XNOR U9138 ( .A(n7647), .B(n6738), .Z(n6739) );
  XNOR U9139 ( .A(y[1503]), .B(x[1503]), .Z(n6738) );
  XNOR U9140 ( .A(y[1504]), .B(x[1504]), .Z(n7647) );
  XNOR U9141 ( .A(n6747), .B(n6746), .Z(n6726) );
  XNOR U9142 ( .A(n7648), .B(n6751), .Z(n6746) );
  XNOR U9143 ( .A(n6744), .B(n6743), .Z(n6751) );
  XNOR U9144 ( .A(n7649), .B(n6742), .Z(n6743) );
  XNOR U9145 ( .A(y[1485]), .B(x[1485]), .Z(n6742) );
  XNOR U9146 ( .A(y[1486]), .B(x[1486]), .Z(n7649) );
  XNOR U9147 ( .A(y[1487]), .B(x[1487]), .Z(n6744) );
  XNOR U9148 ( .A(n6750), .B(n6745), .Z(n7648) );
  XNOR U9149 ( .A(y[1476]), .B(x[1476]), .Z(n6745) );
  XNOR U9150 ( .A(n7650), .B(n6754), .Z(n6750) );
  XNOR U9151 ( .A(y[1490]), .B(x[1490]), .Z(n6754) );
  XNOR U9152 ( .A(n6753), .B(n6749), .Z(n7650) );
  XNOR U9153 ( .A(y[1484]), .B(x[1484]), .Z(n6749) );
  XNOR U9154 ( .A(n7651), .B(n6752), .Z(n6753) );
  XNOR U9155 ( .A(y[1488]), .B(x[1488]), .Z(n6752) );
  XNOR U9156 ( .A(y[1489]), .B(x[1489]), .Z(n7651) );
  XNOR U9157 ( .A(n6758), .B(n6757), .Z(n6747) );
  XNOR U9158 ( .A(n7652), .B(n6761), .Z(n6757) );
  XNOR U9159 ( .A(y[1483]), .B(x[1483]), .Z(n6761) );
  XNOR U9160 ( .A(n6760), .B(n6756), .Z(n7652) );
  XNOR U9161 ( .A(y[1477]), .B(x[1477]), .Z(n6756) );
  XNOR U9162 ( .A(n7653), .B(n6759), .Z(n6760) );
  XNOR U9163 ( .A(y[1481]), .B(x[1481]), .Z(n6759) );
  XNOR U9164 ( .A(y[1482]), .B(x[1482]), .Z(n7653) );
  XOR U9165 ( .A(n6764), .B(n6763), .Z(n6758) );
  XNOR U9166 ( .A(n7654), .B(n6762), .Z(n6763) );
  XNOR U9167 ( .A(y[1478]), .B(x[1478]), .Z(n6762) );
  XNOR U9168 ( .A(y[1479]), .B(x[1479]), .Z(n7654) );
  XOR U9169 ( .A(y[1480]), .B(x[1480]), .Z(n6764) );
  XOR U9170 ( .A(n6822), .B(n6765), .Z(n7623) );
  XNOR U9171 ( .A(y[1345]), .B(x[1345]), .Z(n6765) );
  XOR U9172 ( .A(n7655), .B(n6853), .Z(n6822) );
  XOR U9173 ( .A(n7656), .B(n6789), .Z(n6781) );
  XNOR U9174 ( .A(n6773), .B(n6772), .Z(n6789) );
  XNOR U9175 ( .A(n7657), .B(n6776), .Z(n6772) );
  XNOR U9176 ( .A(y[1561]), .B(x[1561]), .Z(n6776) );
  XNOR U9177 ( .A(n6775), .B(n6771), .Z(n7657) );
  XNOR U9178 ( .A(y[1555]), .B(x[1555]), .Z(n6771) );
  XNOR U9179 ( .A(n7658), .B(n6774), .Z(n6775) );
  XNOR U9180 ( .A(y[1559]), .B(x[1559]), .Z(n6774) );
  XNOR U9181 ( .A(y[1560]), .B(x[1560]), .Z(n7658) );
  XOR U9182 ( .A(n6779), .B(n6778), .Z(n6773) );
  XNOR U9183 ( .A(n7659), .B(n6777), .Z(n6778) );
  XNOR U9184 ( .A(y[1556]), .B(x[1556]), .Z(n6777) );
  XNOR U9185 ( .A(y[1557]), .B(x[1557]), .Z(n7659) );
  XOR U9186 ( .A(y[1558]), .B(x[1558]), .Z(n6779) );
  XNOR U9187 ( .A(n6788), .B(n6780), .Z(n7656) );
  XNOR U9188 ( .A(y[1538]), .B(x[1538]), .Z(n6780) );
  XNOR U9189 ( .A(n7660), .B(n6793), .Z(n6788) );
  XNOR U9190 ( .A(n6786), .B(n6785), .Z(n6793) );
  XNOR U9191 ( .A(n7661), .B(n6784), .Z(n6785) );
  XNOR U9192 ( .A(y[1563]), .B(x[1563]), .Z(n6784) );
  XNOR U9193 ( .A(y[1564]), .B(x[1564]), .Z(n7661) );
  XNOR U9194 ( .A(y[1565]), .B(x[1565]), .Z(n6786) );
  XNOR U9195 ( .A(n6792), .B(n6787), .Z(n7660) );
  XNOR U9196 ( .A(y[1554]), .B(x[1554]), .Z(n6787) );
  XNOR U9197 ( .A(n7662), .B(n6796), .Z(n6792) );
  XNOR U9198 ( .A(y[1568]), .B(x[1568]), .Z(n6796) );
  XNOR U9199 ( .A(n6795), .B(n6791), .Z(n7662) );
  XNOR U9200 ( .A(y[1562]), .B(x[1562]), .Z(n6791) );
  XNOR U9201 ( .A(n7663), .B(n6794), .Z(n6795) );
  XNOR U9202 ( .A(y[1566]), .B(x[1566]), .Z(n6794) );
  XNOR U9203 ( .A(y[1567]), .B(x[1567]), .Z(n7663) );
  XNOR U9204 ( .A(n6803), .B(n6802), .Z(n6782) );
  XNOR U9205 ( .A(n7664), .B(n6807), .Z(n6802) );
  XNOR U9206 ( .A(n6800), .B(n6799), .Z(n6807) );
  XNOR U9207 ( .A(n7665), .B(n6798), .Z(n6799) );
  XNOR U9208 ( .A(y[1548]), .B(x[1548]), .Z(n6798) );
  XNOR U9209 ( .A(y[1549]), .B(x[1549]), .Z(n7665) );
  XNOR U9210 ( .A(y[1550]), .B(x[1550]), .Z(n6800) );
  XNOR U9211 ( .A(n6806), .B(n6801), .Z(n7664) );
  XNOR U9212 ( .A(y[1539]), .B(x[1539]), .Z(n6801) );
  XNOR U9213 ( .A(n7666), .B(n6810), .Z(n6806) );
  XNOR U9214 ( .A(y[1553]), .B(x[1553]), .Z(n6810) );
  XNOR U9215 ( .A(n6809), .B(n6805), .Z(n7666) );
  XNOR U9216 ( .A(y[1547]), .B(x[1547]), .Z(n6805) );
  XNOR U9217 ( .A(n7667), .B(n6808), .Z(n6809) );
  XNOR U9218 ( .A(y[1551]), .B(x[1551]), .Z(n6808) );
  XNOR U9219 ( .A(y[1552]), .B(x[1552]), .Z(n7667) );
  XNOR U9220 ( .A(n6814), .B(n6813), .Z(n6803) );
  XNOR U9221 ( .A(n7668), .B(n6817), .Z(n6813) );
  XNOR U9222 ( .A(y[1546]), .B(x[1546]), .Z(n6817) );
  XNOR U9223 ( .A(n6816), .B(n6812), .Z(n7668) );
  XNOR U9224 ( .A(y[1540]), .B(x[1540]), .Z(n6812) );
  XNOR U9225 ( .A(n7669), .B(n6815), .Z(n6816) );
  XNOR U9226 ( .A(y[1544]), .B(x[1544]), .Z(n6815) );
  XNOR U9227 ( .A(y[1545]), .B(x[1545]), .Z(n7669) );
  XOR U9228 ( .A(n6820), .B(n6819), .Z(n6814) );
  XNOR U9229 ( .A(n7670), .B(n6818), .Z(n6819) );
  XNOR U9230 ( .A(y[1541]), .B(x[1541]), .Z(n6818) );
  XNOR U9231 ( .A(y[1542]), .B(x[1542]), .Z(n7670) );
  XOR U9232 ( .A(y[1543]), .B(x[1543]), .Z(n6820) );
  XOR U9233 ( .A(n6852), .B(n6821), .Z(n7655) );
  XNOR U9234 ( .A(y[1473]), .B(x[1473]), .Z(n6821) );
  XOR U9235 ( .A(n7671), .B(n6869), .Z(n6852) );
  XNOR U9236 ( .A(n6831), .B(n6830), .Z(n6869) );
  XNOR U9237 ( .A(n7672), .B(n6835), .Z(n6830) );
  XNOR U9238 ( .A(n6828), .B(n6827), .Z(n6835) );
  XNOR U9239 ( .A(n7673), .B(n6826), .Z(n6827) );
  XNOR U9240 ( .A(y[1579]), .B(x[1579]), .Z(n6826) );
  XNOR U9241 ( .A(y[1580]), .B(x[1580]), .Z(n7673) );
  XNOR U9242 ( .A(y[1581]), .B(x[1581]), .Z(n6828) );
  XNOR U9243 ( .A(n6834), .B(n6829), .Z(n7672) );
  XNOR U9244 ( .A(y[1570]), .B(x[1570]), .Z(n6829) );
  XNOR U9245 ( .A(n7674), .B(n6838), .Z(n6834) );
  XNOR U9246 ( .A(y[1584]), .B(x[1584]), .Z(n6838) );
  XNOR U9247 ( .A(n6837), .B(n6833), .Z(n7674) );
  XNOR U9248 ( .A(y[1578]), .B(x[1578]), .Z(n6833) );
  XNOR U9249 ( .A(n7675), .B(n6836), .Z(n6837) );
  XNOR U9250 ( .A(y[1582]), .B(x[1582]), .Z(n6836) );
  XNOR U9251 ( .A(y[1583]), .B(x[1583]), .Z(n7675) );
  XNOR U9252 ( .A(n6844), .B(n6843), .Z(n6831) );
  XNOR U9253 ( .A(n7676), .B(n6847), .Z(n6843) );
  XNOR U9254 ( .A(y[1577]), .B(x[1577]), .Z(n6847) );
  XNOR U9255 ( .A(n6846), .B(n6840), .Z(n7676) );
  XNOR U9256 ( .A(y[1571]), .B(x[1571]), .Z(n6840) );
  XNOR U9257 ( .A(n7677), .B(n6845), .Z(n6846) );
  XNOR U9258 ( .A(y[1575]), .B(x[1575]), .Z(n6845) );
  XNOR U9259 ( .A(y[1576]), .B(x[1576]), .Z(n7677) );
  XOR U9260 ( .A(n6850), .B(n6849), .Z(n6844) );
  XNOR U9261 ( .A(n7678), .B(n6848), .Z(n6849) );
  XNOR U9262 ( .A(y[1572]), .B(x[1572]), .Z(n6848) );
  XNOR U9263 ( .A(y[1573]), .B(x[1573]), .Z(n7678) );
  XOR U9264 ( .A(y[1574]), .B(x[1574]), .Z(n6850) );
  XOR U9265 ( .A(n6868), .B(n6851), .Z(n7671) );
  XNOR U9266 ( .A(y[1537]), .B(x[1537]), .Z(n6851) );
  XOR U9267 ( .A(n7679), .B(n6876), .Z(n6868) );
  XNOR U9268 ( .A(n6860), .B(n6859), .Z(n6876) );
  XNOR U9269 ( .A(n7680), .B(n6863), .Z(n6859) );
  XNOR U9270 ( .A(y[1592]), .B(x[1592]), .Z(n6863) );
  XNOR U9271 ( .A(n6862), .B(n6856), .Z(n7680) );
  XNOR U9272 ( .A(y[1586]), .B(x[1586]), .Z(n6856) );
  XNOR U9273 ( .A(n7681), .B(n6861), .Z(n6862) );
  XNOR U9274 ( .A(y[1590]), .B(x[1590]), .Z(n6861) );
  XNOR U9275 ( .A(y[1591]), .B(x[1591]), .Z(n7681) );
  XOR U9276 ( .A(n6866), .B(n6865), .Z(n6860) );
  XNOR U9277 ( .A(n7682), .B(n6864), .Z(n6865) );
  XNOR U9278 ( .A(y[1587]), .B(x[1587]), .Z(n6864) );
  XNOR U9279 ( .A(y[1588]), .B(x[1588]), .Z(n7682) );
  XOR U9280 ( .A(y[1589]), .B(x[1589]), .Z(n6866) );
  XNOR U9281 ( .A(n6875), .B(n6867), .Z(n7679) );
  XNOR U9282 ( .A(y[1569]), .B(x[1569]), .Z(n6867) );
  XNOR U9283 ( .A(n7683), .B(n6880), .Z(n6875) );
  XNOR U9284 ( .A(n6873), .B(n6872), .Z(n6880) );
  XNOR U9285 ( .A(n7684), .B(n6871), .Z(n6872) );
  XNOR U9286 ( .A(y[1594]), .B(x[1594]), .Z(n6871) );
  XNOR U9287 ( .A(y[1595]), .B(x[1595]), .Z(n7684) );
  XNOR U9288 ( .A(y[1596]), .B(x[1596]), .Z(n6873) );
  XNOR U9289 ( .A(n6879), .B(n6874), .Z(n7683) );
  XNOR U9290 ( .A(y[1585]), .B(x[1585]), .Z(n6874) );
  XNOR U9291 ( .A(n7685), .B(n6883), .Z(n6879) );
  XNOR U9292 ( .A(y[1599]), .B(x[1599]), .Z(n6883) );
  XNOR U9293 ( .A(n6882), .B(n6878), .Z(n7685) );
  XNOR U9294 ( .A(y[1593]), .B(x[1593]), .Z(n6878) );
  XNOR U9295 ( .A(n7686), .B(n6881), .Z(n6882) );
  XNOR U9296 ( .A(y[1597]), .B(x[1597]), .Z(n6881) );
  XNOR U9297 ( .A(y[1598]), .B(x[1598]), .Z(n7686) );
endmodule

