
module hamming_N16000_CC32 ( clk, rst, x, y, o );
  input [499:0] x;
  input [499:0] y;
  output [13:0] o;
  input clk, rst;
  wire   n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056;
  wire   [13:0] oglobal;

  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[0]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[1]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[2]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[3]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[4]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[5]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[6]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[7]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[8]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[9]) );
  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[10]) );
  DFF \oglobal_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[11]) );
  DFF \oglobal_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[12]) );
  DFF \oglobal_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[13]) );
  XNOR U517 ( .A(n410), .B(n795), .Z(n416) );
  XNOR U518 ( .A(n476), .B(n477), .Z(n489) );
  XNOR U519 ( .A(n554), .B(n1023), .Z(n560) );
  XNOR U520 ( .A(n190), .B(n362), .Z(n192) );
  XNOR U521 ( .A(n268), .B(n514), .Z(n274) );
  XNOR U522 ( .A(n292), .B(n562), .Z(n298) );
  XNOR U523 ( .A(n341), .B(n658), .Z(n347) );
  XNOR U524 ( .A(n124), .B(n227), .Z(n130) );
  XNOR U525 ( .A(n174), .B(n325), .Z(n180) );
  XNOR U526 ( .A(n154), .B(n251), .Z(n137) );
  XNOR U527 ( .A(n379), .B(n682), .Z(n354) );
  XNOR U528 ( .A(n530), .B(n985), .Z(n536) );
  XNOR U529 ( .A(n500), .B(n501), .Z(n513) );
  XNOR U530 ( .A(n620), .B(n621), .Z(n633) );
  XNOR U531 ( .A(n668), .B(n669), .Z(n681) );
  XNOR U532 ( .A(n723), .B(n1289), .Z(n729) );
  XNOR U533 ( .A(n692), .B(n693), .Z(n705) );
  XNOR U534 ( .A(n243), .B(n466), .Z(n249) );
  XNOR U535 ( .A(n608), .B(n609), .Z(n616) );
  XNOR U536 ( .A(n656), .B(n657), .Z(n664) );
  XNOR U537 ( .A(n753), .B(n754), .Z(n761) );
  XNOR U538 ( .A(n1026), .B(n1028), .Z(n1047) );
  XNOR U539 ( .A(n1102), .B(n1104), .Z(n1123) );
  XNOR U540 ( .A(n198), .B(n374), .Z(n204) );
  XNOR U541 ( .A(n225), .B(n226), .Z(n233) );
  XNOR U542 ( .A(n423), .B(n424), .Z(n448) );
  XNOR U543 ( .A(n567), .B(n1004), .Z(n543) );
  XNOR U544 ( .A(n817), .B(n819), .Z(n857) );
  XNOR U545 ( .A(n103), .B(n182), .Z(n109) );
  XNOR U546 ( .A(n281), .B(n490), .Z(n256) );
  XNOR U547 ( .A(n58), .B(n87), .Z(n64) );
  XNOR U548 ( .A(n354), .B(n586), .Z(n305) );
  XNOR U549 ( .A(n458), .B(n871), .Z(n464) );
  XNOR U550 ( .A(n506), .B(n947), .Z(n512) );
  XNOR U551 ( .A(n602), .B(n1099), .Z(n608) );
  XNOR U552 ( .A(n626), .B(n1137), .Z(n632) );
  XNOR U553 ( .A(n650), .B(n1175), .Z(n656) );
  XNOR U554 ( .A(n674), .B(n1213), .Z(n680) );
  XNOR U555 ( .A(n698), .B(n1251), .Z(n704) );
  XNOR U556 ( .A(n747), .B(n1327), .Z(n753) );
  XNOR U557 ( .A(n765), .B(n766), .Z(n778) );
  XNOR U558 ( .A(n219), .B(n418), .Z(n225) );
  XNOR U559 ( .A(n317), .B(n610), .Z(n323) );
  XNOR U560 ( .A(n536), .B(n966), .Z(n519) );
  XNOR U561 ( .A(n729), .B(n1270), .Z(n712) );
  XNOR U562 ( .A(n1064), .B(n1678), .Z(n1045) );
  XNOR U563 ( .A(n1330), .B(n1332), .Z(n1351) );
  XNOR U564 ( .A(n117), .B(n119), .Z(n131) );
  XNOR U565 ( .A(n148), .B(n276), .Z(n154) );
  XNOR U566 ( .A(n249), .B(n442), .Z(n232) );
  XNOR U567 ( .A(n347), .B(n634), .Z(n330) );
  XNOR U568 ( .A(n969), .B(n971), .Z(n1009) );
  XNOR U569 ( .A(n1273), .B(n1275), .Z(n1313) );
  XNOR U570 ( .A(n79), .B(n132), .Z(n85) );
  XNOR U571 ( .A(n204), .B(n349), .Z(n187) );
  XNOR U572 ( .A(n447), .B(n448), .Z(n496) );
  XNOR U573 ( .A(n855), .B(n857), .Z(n933) );
  XNOR U574 ( .A(n1159), .B(n1161), .Z(n1237) );
  XNOR U575 ( .A(n109), .B(n156), .Z(n92) );
  XNOR U576 ( .A(n687), .B(n1080), .Z(n591) );
  XOR U577 ( .A(oglobal[7]), .B(n46), .Z(n17) );
  XOR U578 ( .A(oglobal[4]), .B(n207), .Z(n23) );
  ANDN U579 ( .B(n1822), .A(n1181), .Z(n1183) );
  ANDN U580 ( .B(n2036), .A(n1371), .Z(n1373) );
  XNOR U581 ( .A(n235), .B(n454), .Z(n237) );
  XNOR U582 ( .A(n382), .B(n743), .Z(n384) );
  XNOR U583 ( .A(n548), .B(n549), .Z(n561) );
  XNOR U584 ( .A(n578), .B(n1061), .Z(n584) );
  XNOR U585 ( .A(n644), .B(n645), .Z(n657) );
  XNOR U586 ( .A(n717), .B(n718), .Z(n730) );
  XNOR U587 ( .A(n2024), .B(n2023), .Z(n2043) );
  XNOR U588 ( .A(n2003), .B(n2002), .Z(n2000) );
  XNOR U589 ( .A(n1961), .B(n1960), .Z(n1958) );
  XNOR U590 ( .A(n1919), .B(n1918), .Z(n1916) );
  XNOR U591 ( .A(n1877), .B(n1876), .Z(n1874) );
  XNOR U592 ( .A(n1812), .B(n1811), .Z(n1829) );
  XNOR U593 ( .A(n1770), .B(n1769), .Z(n1789) );
  XNOR U594 ( .A(n1751), .B(n1750), .Z(n1748) );
  XNOR U595 ( .A(n1625), .B(n1624), .Z(n1622) );
  XNOR U596 ( .A(n1583), .B(n1582), .Z(n1580) );
  XNOR U597 ( .A(n1543), .B(n1542), .Z(n1540) );
  XNOR U598 ( .A(n1499), .B(n1498), .Z(n1496) );
  XNOR U599 ( .A(n1459), .B(n1458), .Z(n1456) );
  XNOR U600 ( .A(n1417), .B(n1416), .Z(n1414) );
  XNOR U601 ( .A(n140), .B(n264), .Z(n142) );
  XNOR U602 ( .A(n310), .B(n312), .Z(n324) );
  XNOR U603 ( .A(n390), .B(n755), .Z(n396) );
  XNOR U604 ( .A(n440), .B(n814), .Z(n423) );
  XNOR U605 ( .A(n704), .B(n705), .Z(n713) );
  XNOR U606 ( .A(n874), .B(n876), .Z(n895) );
  XNOR U607 ( .A(n950), .B(n952), .Z(n971) );
  XNOR U608 ( .A(n1178), .B(n1180), .Z(n1199) );
  XNOR U609 ( .A(n298), .B(n538), .Z(n281) );
  XNOR U610 ( .A(n471), .B(n852), .Z(n447) );
  XNOR U611 ( .A(n760), .B(n1308), .Z(n736) );
  XNOR U612 ( .A(n1121), .B(n1123), .Z(n1161) );
  XNOR U613 ( .A(n72), .B(n74), .Z(n86) );
  XNOR U614 ( .A(n130), .B(n131), .Z(n138) );
  XNOR U615 ( .A(n232), .B(n233), .Z(n257) );
  XNOR U616 ( .A(n543), .B(n928), .Z(n495) );
  XNOR U617 ( .A(n639), .B(n640), .Z(n688) );
  XNOR U618 ( .A(n1311), .B(n1888), .Z(n1235) );
  XNOR U619 ( .A(n41), .B(n54), .Z(n43) );
  XNOR U620 ( .A(n187), .B(n300), .Z(n161) );
  XNOR U621 ( .A(n931), .B(n933), .Z(n1085) );
  XOR U622 ( .A(oglobal[6]), .B(n67), .Z(n19) );
  XOR U623 ( .A(oglobal[3]), .B(n399), .Z(n25) );
  ANDN U624 ( .B(n1448), .A(n839), .Z(n841) );
  ANDN U625 ( .B(n1532), .A(n915), .Z(n917) );
  XNOR U626 ( .A(n284), .B(n550), .Z(n286) );
  XNOR U627 ( .A(n333), .B(n646), .Z(n335) );
  XNOR U628 ( .A(n404), .B(n405), .Z(n417) );
  XNOR U629 ( .A(n428), .B(n429), .Z(n441) );
  XNOR U630 ( .A(n452), .B(n453), .Z(n465) );
  XNOR U631 ( .A(n524), .B(n525), .Z(n537) );
  XNOR U632 ( .A(n572), .B(n573), .Z(n585) );
  XNOR U633 ( .A(n596), .B(n597), .Z(n609) );
  XNOR U634 ( .A(n741), .B(n742), .Z(n754) );
  XNOR U635 ( .A(n771), .B(n1365), .Z(n777) );
  XNOR U636 ( .A(n1938), .B(n1937), .Z(n1957) );
  XNOR U637 ( .A(n1898), .B(n1897), .Z(n1915) );
  XNOR U638 ( .A(n1793), .B(n1792), .Z(n1790) );
  XNOR U639 ( .A(n1730), .B(n1729), .Z(n1747) );
  XNOR U640 ( .A(n1711), .B(n1710), .Z(n1708) );
  XNOR U641 ( .A(n1667), .B(n1666), .Z(n1664) );
  XNOR U642 ( .A(n1602), .B(n1601), .Z(n1621) );
  XNOR U643 ( .A(n1562), .B(n1561), .Z(n1579) );
  XNOR U644 ( .A(n1520), .B(n1519), .Z(n1539) );
  XNOR U645 ( .A(n1478), .B(n1477), .Z(n1495) );
  XNOR U646 ( .A(n1436), .B(n1435), .Z(n1455) );
  XNOR U647 ( .A(n1396), .B(n1395), .Z(n1413) );
  XNOR U648 ( .A(n261), .B(n263), .Z(n275) );
  XNOR U649 ( .A(n359), .B(n361), .Z(n373) );
  XNOR U650 ( .A(n488), .B(n890), .Z(n471) );
  XNOR U651 ( .A(n512), .B(n513), .Z(n520) );
  XNOR U652 ( .A(n560), .B(n561), .Z(n568) );
  XNOR U653 ( .A(n632), .B(n1118), .Z(n615) );
  XNOR U654 ( .A(n798), .B(n800), .Z(n819) );
  XNOR U655 ( .A(n1216), .B(n1844), .Z(n1197) );
  XNOR U656 ( .A(n1254), .B(n1256), .Z(n1275) );
  XNOR U657 ( .A(n1368), .B(n2014), .Z(n1349) );
  XNOR U658 ( .A(n396), .B(n731), .Z(n379) );
  XNOR U659 ( .A(n663), .B(n1156), .Z(n639) );
  XNOR U660 ( .A(n893), .B(n1468), .Z(n855) );
  XNOR U661 ( .A(n97), .B(n98), .Z(n110) );
  XNOR U662 ( .A(n180), .B(n181), .Z(n188) );
  XNOR U663 ( .A(n330), .B(n331), .Z(n355) );
  XNOR U664 ( .A(n736), .B(n1232), .Z(n687) );
  XNOR U665 ( .A(n1007), .B(n1552), .Z(n931) );
  XNOR U666 ( .A(n51), .B(n53), .Z(n65) );
  XNOR U667 ( .A(n85), .B(n86), .Z(n93) );
  XNOR U668 ( .A(n137), .B(n138), .Z(n162) );
  XNOR U669 ( .A(n256), .B(n257), .Z(n306) );
  XNOR U670 ( .A(n495), .B(n496), .Z(n592) );
  XNOR U671 ( .A(n1235), .B(n1720), .Z(n1083) );
  XOR U672 ( .A(oglobal[8]), .B(n38), .Z(n15) );
  XOR U673 ( .A(oglobal[5]), .B(n112), .Z(n21) );
  XOR U674 ( .A(oglobal[2]), .B(n780), .Z(n27) );
  ANDN U675 ( .B(n1406), .A(n801), .Z(n803) );
  ANDN U676 ( .B(n1488), .A(n877), .Z(n879) );
  ANDN U677 ( .B(n1572), .A(n953), .Z(n955) );
  ANDN U678 ( .B(n1614), .A(n991), .Z(n993) );
  ANDN U679 ( .B(n1656), .A(n1029), .Z(n1031) );
  ANDN U680 ( .B(n1700), .A(n1067), .Z(n1069) );
  ANDN U681 ( .B(n1740), .A(n1105), .Z(n1107) );
  ANDN U682 ( .B(n1782), .A(n1143), .Z(n1145) );
  ANDN U683 ( .B(n1866), .A(n1219), .Z(n1221) );
  ANDN U684 ( .B(n1908), .A(n1257), .Z(n1259) );
  ANDN U685 ( .B(n1950), .A(n1295), .Z(n1297) );
  ANDN U686 ( .B(n1992), .A(n1333), .Z(n1335) );
  XNOR U687 ( .A(n434), .B(n833), .Z(n440) );
  XNOR U688 ( .A(n482), .B(n909), .Z(n488) );
  XNOR U689 ( .A(n2047), .B(n2046), .Z(n2044) );
  XNOR U690 ( .A(n1982), .B(n1981), .Z(n1999) );
  XNOR U691 ( .A(n1854), .B(n1853), .Z(n1873) );
  XNOR U692 ( .A(n1833), .B(n1832), .Z(n1830) );
  XNOR U693 ( .A(n1688), .B(n1687), .Z(n1707) );
  XNOR U694 ( .A(n1646), .B(n1645), .Z(n1663) );
  XNOR U695 ( .A(n212), .B(n214), .Z(n226) );
  XNOR U696 ( .A(n237), .B(n238), .Z(n250) );
  XNOR U697 ( .A(n286), .B(n287), .Z(n299) );
  XNOR U698 ( .A(n335), .B(n336), .Z(n348) );
  XNOR U699 ( .A(n384), .B(n385), .Z(n397) );
  XNOR U700 ( .A(n416), .B(n417), .Z(n424) );
  XNOR U701 ( .A(n464), .B(n465), .Z(n472) );
  XNOR U702 ( .A(n584), .B(n1042), .Z(n567) );
  XNOR U703 ( .A(n680), .B(n1194), .Z(n663) );
  XNOR U704 ( .A(n777), .B(n1346), .Z(n760) );
  XNOR U705 ( .A(n836), .B(n1426), .Z(n817) );
  XNOR U706 ( .A(n912), .B(n1510), .Z(n893) );
  XNOR U707 ( .A(n988), .B(n1592), .Z(n969) );
  XNOR U708 ( .A(n1140), .B(n1760), .Z(n1121) );
  XNOR U709 ( .A(n1292), .B(n1928), .Z(n1273) );
  XNOR U710 ( .A(n142), .B(n143), .Z(n155) );
  XNOR U711 ( .A(n166), .B(n168), .Z(n181) );
  XNOR U712 ( .A(n192), .B(n193), .Z(n205) );
  XNOR U713 ( .A(n274), .B(n275), .Z(n282) );
  XNOR U714 ( .A(n323), .B(n324), .Z(n331) );
  XNOR U715 ( .A(n372), .B(n373), .Z(n380) );
  XNOR U716 ( .A(n519), .B(n520), .Z(n544) );
  XNOR U717 ( .A(n615), .B(n616), .Z(n640) );
  XNOR U718 ( .A(n712), .B(n713), .Z(n737) );
  XNOR U719 ( .A(n1045), .B(n1636), .Z(n1007) );
  XNOR U720 ( .A(n1197), .B(n1802), .Z(n1159) );
  XNOR U721 ( .A(n1349), .B(n1972), .Z(n1311) );
  XNOR U722 ( .A(n43), .B(n44), .Z(n18) );
  XNOR U723 ( .A(n64), .B(n65), .Z(n20) );
  XNOR U724 ( .A(n92), .B(n93), .Z(n22) );
  XNOR U725 ( .A(n161), .B(n162), .Z(n24) );
  XNOR U726 ( .A(n305), .B(n306), .Z(n26) );
  XNOR U727 ( .A(n591), .B(n592), .Z(n28) );
  XNOR U728 ( .A(n1083), .B(n1085), .Z(n30) );
  XNOR U729 ( .A(n15), .B(n16), .Z(o[8]) );
  XOR U730 ( .A(n17), .B(n18), .Z(o[7]) );
  XOR U731 ( .A(n19), .B(n20), .Z(o[6]) );
  XOR U732 ( .A(n21), .B(n22), .Z(o[5]) );
  XOR U733 ( .A(n23), .B(n24), .Z(o[4]) );
  XOR U734 ( .A(n25), .B(n26), .Z(o[3]) );
  XOR U735 ( .A(n27), .B(n28), .Z(o[2]) );
  XOR U736 ( .A(n29), .B(n30), .Z(o[1]) );
  XOR U737 ( .A(n31), .B(n32), .Z(o[13]) );
  XOR U738 ( .A(oglobal[13]), .B(n33), .Z(n32) );
  AND U739 ( .A(n31), .B(o[12]), .Z(n33) );
  XOR U740 ( .A(oglobal[12]), .B(n31), .Z(o[12]) );
  ANDN U741 ( .B(n34), .A(o[11]), .Z(n31) );
  XOR U742 ( .A(oglobal[11]), .B(n34), .Z(o[11]) );
  ANDN U743 ( .B(n35), .A(o[10]), .Z(n34) );
  XOR U744 ( .A(oglobal[10]), .B(n35), .Z(o[10]) );
  ANDN U745 ( .B(n36), .A(o[9]), .Z(n35) );
  XOR U746 ( .A(oglobal[9]), .B(n36), .Z(o[9]) );
  XNOR U747 ( .A(n37), .B(n38), .Z(n36) );
  ANDN U748 ( .B(n39), .A(n15), .Z(n37) );
  XNOR U749 ( .A(n38), .B(n16), .Z(n39) );
  XNOR U750 ( .A(n40), .B(n41), .Z(n16) );
  ANDN U751 ( .B(n42), .A(n43), .Z(n40) );
  XOR U752 ( .A(n41), .B(n44), .Z(n42) );
  XOR U753 ( .A(n45), .B(n46), .Z(n38) );
  ANDN U754 ( .B(n47), .A(n17), .Z(n45) );
  XOR U755 ( .A(n46), .B(n18), .Z(n47) );
  XNOR U756 ( .A(n48), .B(n49), .Z(n44) );
  ANDN U757 ( .B(n50), .A(n51), .Z(n48) );
  XOR U758 ( .A(n52), .B(n53), .Z(n50) );
  XNOR U759 ( .A(n55), .B(n56), .Z(n54) );
  ANDN U760 ( .B(n57), .A(n58), .Z(n55) );
  XNOR U761 ( .A(n59), .B(n60), .Z(n57) );
  XOR U762 ( .A(n61), .B(n62), .Z(n41) );
  ANDN U763 ( .B(n63), .A(n64), .Z(n61) );
  XOR U764 ( .A(n62), .B(n65), .Z(n63) );
  XOR U765 ( .A(n66), .B(n67), .Z(n46) );
  ANDN U766 ( .B(n68), .A(n19), .Z(n66) );
  XOR U767 ( .A(n67), .B(n20), .Z(n68) );
  XNOR U768 ( .A(n69), .B(n70), .Z(n53) );
  ANDN U769 ( .B(n71), .A(n72), .Z(n69) );
  XOR U770 ( .A(n73), .B(n74), .Z(n71) );
  XOR U771 ( .A(n49), .B(n75), .Z(n51) );
  XNOR U772 ( .A(n76), .B(n77), .Z(n75) );
  ANDN U773 ( .B(n78), .A(n79), .Z(n76) );
  XNOR U774 ( .A(n80), .B(n81), .Z(n78) );
  IV U775 ( .A(n52), .Z(n49) );
  XOR U776 ( .A(n82), .B(n83), .Z(n52) );
  ANDN U777 ( .B(n84), .A(n85), .Z(n82) );
  XOR U778 ( .A(n83), .B(n86), .Z(n84) );
  XNOR U779 ( .A(n59), .B(n88), .Z(n87) );
  IV U780 ( .A(n62), .Z(n88) );
  XOR U781 ( .A(n89), .B(n90), .Z(n62) );
  ANDN U782 ( .B(n91), .A(n92), .Z(n89) );
  XOR U783 ( .A(n90), .B(n93), .Z(n91) );
  XNOR U784 ( .A(n94), .B(n95), .Z(n59) );
  ANDN U785 ( .B(n96), .A(n97), .Z(n94) );
  XOR U786 ( .A(n95), .B(n98), .Z(n96) );
  XOR U787 ( .A(n56), .B(n99), .Z(n58) );
  XNOR U788 ( .A(n100), .B(n101), .Z(n99) );
  ANDN U789 ( .B(n102), .A(n103), .Z(n100) );
  XNOR U790 ( .A(n104), .B(n105), .Z(n102) );
  IV U791 ( .A(n60), .Z(n56) );
  XOR U792 ( .A(n106), .B(n107), .Z(n60) );
  ANDN U793 ( .B(n108), .A(n109), .Z(n106) );
  XOR U794 ( .A(n110), .B(n107), .Z(n108) );
  XOR U795 ( .A(n111), .B(n112), .Z(n67) );
  ANDN U796 ( .B(n113), .A(n21), .Z(n111) );
  XOR U797 ( .A(n112), .B(n22), .Z(n113) );
  XNOR U798 ( .A(n114), .B(n115), .Z(n74) );
  ANDN U799 ( .B(n116), .A(n117), .Z(n114) );
  XOR U800 ( .A(n118), .B(n119), .Z(n116) );
  XOR U801 ( .A(n70), .B(n120), .Z(n72) );
  XNOR U802 ( .A(n121), .B(n122), .Z(n120) );
  ANDN U803 ( .B(n123), .A(n124), .Z(n121) );
  XNOR U804 ( .A(n125), .B(n126), .Z(n123) );
  IV U805 ( .A(n73), .Z(n70) );
  XOR U806 ( .A(n127), .B(n128), .Z(n73) );
  ANDN U807 ( .B(n129), .A(n130), .Z(n127) );
  XOR U808 ( .A(n128), .B(n131), .Z(n129) );
  XNOR U809 ( .A(n80), .B(n133), .Z(n132) );
  IV U810 ( .A(n83), .Z(n133) );
  XOR U811 ( .A(n134), .B(n135), .Z(n83) );
  ANDN U812 ( .B(n136), .A(n137), .Z(n134) );
  XOR U813 ( .A(n135), .B(n138), .Z(n136) );
  XNOR U814 ( .A(n139), .B(n140), .Z(n80) );
  ANDN U815 ( .B(n141), .A(n142), .Z(n139) );
  XOR U816 ( .A(n140), .B(n143), .Z(n141) );
  XOR U817 ( .A(n77), .B(n144), .Z(n79) );
  XNOR U818 ( .A(n145), .B(n146), .Z(n144) );
  ANDN U819 ( .B(n147), .A(n148), .Z(n145) );
  XNOR U820 ( .A(n149), .B(n150), .Z(n147) );
  IV U821 ( .A(n81), .Z(n77) );
  XOR U822 ( .A(n151), .B(n152), .Z(n81) );
  ANDN U823 ( .B(n153), .A(n154), .Z(n151) );
  XOR U824 ( .A(n155), .B(n152), .Z(n153) );
  XOR U825 ( .A(n110), .B(n157), .Z(n156) );
  IV U826 ( .A(n90), .Z(n157) );
  XOR U827 ( .A(n158), .B(n159), .Z(n90) );
  ANDN U828 ( .B(n160), .A(n161), .Z(n158) );
  XOR U829 ( .A(n159), .B(n162), .Z(n160) );
  XNOR U830 ( .A(n163), .B(n164), .Z(n98) );
  ANDN U831 ( .B(n165), .A(n166), .Z(n163) );
  XOR U832 ( .A(n167), .B(n168), .Z(n165) );
  XOR U833 ( .A(n169), .B(n170), .Z(n97) );
  XNOR U834 ( .A(n171), .B(n172), .Z(n170) );
  ANDN U835 ( .B(n173), .A(n174), .Z(n171) );
  XNOR U836 ( .A(n175), .B(n176), .Z(n173) );
  IV U837 ( .A(n95), .Z(n169) );
  XOR U838 ( .A(n177), .B(n178), .Z(n95) );
  ANDN U839 ( .B(n179), .A(n180), .Z(n177) );
  XOR U840 ( .A(n178), .B(n181), .Z(n179) );
  XNOR U841 ( .A(n104), .B(n183), .Z(n182) );
  IV U842 ( .A(n107), .Z(n183) );
  XOR U843 ( .A(n184), .B(n185), .Z(n107) );
  ANDN U844 ( .B(n186), .A(n187), .Z(n184) );
  XOR U845 ( .A(n188), .B(n185), .Z(n186) );
  XNOR U846 ( .A(n189), .B(n190), .Z(n104) );
  ANDN U847 ( .B(n191), .A(n192), .Z(n189) );
  XOR U848 ( .A(n190), .B(n193), .Z(n191) );
  XOR U849 ( .A(n101), .B(n194), .Z(n103) );
  XNOR U850 ( .A(n195), .B(n196), .Z(n194) );
  ANDN U851 ( .B(n197), .A(n198), .Z(n195) );
  XNOR U852 ( .A(n199), .B(n200), .Z(n197) );
  IV U853 ( .A(n105), .Z(n101) );
  XOR U854 ( .A(n201), .B(n202), .Z(n105) );
  ANDN U855 ( .B(n203), .A(n204), .Z(n201) );
  XOR U856 ( .A(n205), .B(n202), .Z(n203) );
  XOR U857 ( .A(n206), .B(n207), .Z(n112) );
  ANDN U858 ( .B(n208), .A(n23), .Z(n206) );
  XOR U859 ( .A(n207), .B(n24), .Z(n208) );
  XNOR U860 ( .A(n209), .B(n210), .Z(n119) );
  ANDN U861 ( .B(n211), .A(n212), .Z(n209) );
  XOR U862 ( .A(n213), .B(n214), .Z(n211) );
  XOR U863 ( .A(n115), .B(n215), .Z(n117) );
  XNOR U864 ( .A(n216), .B(n217), .Z(n215) );
  ANDN U865 ( .B(n218), .A(n219), .Z(n216) );
  XNOR U866 ( .A(n220), .B(n221), .Z(n218) );
  IV U867 ( .A(n118), .Z(n115) );
  XOR U868 ( .A(n222), .B(n223), .Z(n118) );
  ANDN U869 ( .B(n224), .A(n225), .Z(n222) );
  XOR U870 ( .A(n223), .B(n226), .Z(n224) );
  XNOR U871 ( .A(n125), .B(n228), .Z(n227) );
  IV U872 ( .A(n128), .Z(n228) );
  XOR U873 ( .A(n229), .B(n230), .Z(n128) );
  ANDN U874 ( .B(n231), .A(n232), .Z(n229) );
  XOR U875 ( .A(n230), .B(n233), .Z(n231) );
  XNOR U876 ( .A(n234), .B(n235), .Z(n125) );
  ANDN U877 ( .B(n236), .A(n237), .Z(n234) );
  XOR U878 ( .A(n235), .B(n238), .Z(n236) );
  XOR U879 ( .A(n122), .B(n239), .Z(n124) );
  XNOR U880 ( .A(n240), .B(n241), .Z(n239) );
  ANDN U881 ( .B(n242), .A(n243), .Z(n240) );
  XNOR U882 ( .A(n244), .B(n245), .Z(n242) );
  IV U883 ( .A(n126), .Z(n122) );
  XOR U884 ( .A(n246), .B(n247), .Z(n126) );
  ANDN U885 ( .B(n248), .A(n249), .Z(n246) );
  XOR U886 ( .A(n250), .B(n247), .Z(n248) );
  XOR U887 ( .A(n155), .B(n252), .Z(n251) );
  IV U888 ( .A(n135), .Z(n252) );
  XOR U889 ( .A(n253), .B(n254), .Z(n135) );
  ANDN U890 ( .B(n255), .A(n256), .Z(n253) );
  XOR U891 ( .A(n254), .B(n257), .Z(n255) );
  XNOR U892 ( .A(n258), .B(n259), .Z(n143) );
  ANDN U893 ( .B(n260), .A(n261), .Z(n258) );
  XOR U894 ( .A(n262), .B(n263), .Z(n260) );
  XNOR U895 ( .A(n265), .B(n266), .Z(n264) );
  ANDN U896 ( .B(n267), .A(n268), .Z(n265) );
  XNOR U897 ( .A(n269), .B(n270), .Z(n267) );
  XOR U898 ( .A(n271), .B(n272), .Z(n140) );
  ANDN U899 ( .B(n273), .A(n274), .Z(n271) );
  XOR U900 ( .A(n272), .B(n275), .Z(n273) );
  XNOR U901 ( .A(n149), .B(n277), .Z(n276) );
  IV U902 ( .A(n152), .Z(n277) );
  XOR U903 ( .A(n278), .B(n279), .Z(n152) );
  ANDN U904 ( .B(n280), .A(n281), .Z(n278) );
  XOR U905 ( .A(n282), .B(n279), .Z(n280) );
  XNOR U906 ( .A(n283), .B(n284), .Z(n149) );
  ANDN U907 ( .B(n285), .A(n286), .Z(n283) );
  XOR U908 ( .A(n284), .B(n287), .Z(n285) );
  XOR U909 ( .A(n146), .B(n288), .Z(n148) );
  XNOR U910 ( .A(n289), .B(n290), .Z(n288) );
  ANDN U911 ( .B(n291), .A(n292), .Z(n289) );
  XNOR U912 ( .A(n293), .B(n294), .Z(n291) );
  IV U913 ( .A(n150), .Z(n146) );
  XOR U914 ( .A(n295), .B(n296), .Z(n150) );
  ANDN U915 ( .B(n297), .A(n298), .Z(n295) );
  XOR U916 ( .A(n299), .B(n296), .Z(n297) );
  XOR U917 ( .A(n188), .B(n301), .Z(n300) );
  IV U918 ( .A(n159), .Z(n301) );
  XOR U919 ( .A(n302), .B(n303), .Z(n159) );
  ANDN U920 ( .B(n304), .A(n305), .Z(n302) );
  XOR U921 ( .A(n303), .B(n306), .Z(n304) );
  XNOR U922 ( .A(n307), .B(n308), .Z(n168) );
  ANDN U923 ( .B(n309), .A(n310), .Z(n307) );
  XOR U924 ( .A(n311), .B(n312), .Z(n309) );
  XOR U925 ( .A(n164), .B(n313), .Z(n166) );
  XNOR U926 ( .A(n314), .B(n315), .Z(n313) );
  ANDN U927 ( .B(n316), .A(n317), .Z(n314) );
  XNOR U928 ( .A(n318), .B(n319), .Z(n316) );
  IV U929 ( .A(n167), .Z(n164) );
  XOR U930 ( .A(n320), .B(n321), .Z(n167) );
  ANDN U931 ( .B(n322), .A(n323), .Z(n320) );
  XOR U932 ( .A(n321), .B(n324), .Z(n322) );
  XNOR U933 ( .A(n175), .B(n326), .Z(n325) );
  IV U934 ( .A(n178), .Z(n326) );
  XOR U935 ( .A(n327), .B(n328), .Z(n178) );
  ANDN U936 ( .B(n329), .A(n330), .Z(n327) );
  XOR U937 ( .A(n328), .B(n331), .Z(n329) );
  XNOR U938 ( .A(n332), .B(n333), .Z(n175) );
  ANDN U939 ( .B(n334), .A(n335), .Z(n332) );
  XOR U940 ( .A(n333), .B(n336), .Z(n334) );
  XOR U941 ( .A(n172), .B(n337), .Z(n174) );
  XNOR U942 ( .A(n338), .B(n339), .Z(n337) );
  ANDN U943 ( .B(n340), .A(n341), .Z(n338) );
  XNOR U944 ( .A(n342), .B(n343), .Z(n340) );
  IV U945 ( .A(n176), .Z(n172) );
  XOR U946 ( .A(n344), .B(n345), .Z(n176) );
  ANDN U947 ( .B(n346), .A(n347), .Z(n344) );
  XOR U948 ( .A(n348), .B(n345), .Z(n346) );
  XOR U949 ( .A(n205), .B(n350), .Z(n349) );
  IV U950 ( .A(n185), .Z(n350) );
  XOR U951 ( .A(n351), .B(n352), .Z(n185) );
  ANDN U952 ( .B(n353), .A(n354), .Z(n351) );
  XOR U953 ( .A(n355), .B(n352), .Z(n353) );
  XNOR U954 ( .A(n356), .B(n357), .Z(n193) );
  ANDN U955 ( .B(n358), .A(n359), .Z(n356) );
  XOR U956 ( .A(n360), .B(n361), .Z(n358) );
  XNOR U957 ( .A(n363), .B(n364), .Z(n362) );
  ANDN U958 ( .B(n365), .A(n366), .Z(n363) );
  XNOR U959 ( .A(n367), .B(n368), .Z(n365) );
  XOR U960 ( .A(n369), .B(n370), .Z(n190) );
  ANDN U961 ( .B(n371), .A(n372), .Z(n369) );
  XOR U962 ( .A(n370), .B(n373), .Z(n371) );
  XNOR U963 ( .A(n199), .B(n375), .Z(n374) );
  IV U964 ( .A(n202), .Z(n375) );
  XOR U965 ( .A(n376), .B(n377), .Z(n202) );
  ANDN U966 ( .B(n378), .A(n379), .Z(n376) );
  XOR U967 ( .A(n380), .B(n377), .Z(n378) );
  XNOR U968 ( .A(n381), .B(n382), .Z(n199) );
  ANDN U969 ( .B(n383), .A(n384), .Z(n381) );
  XOR U970 ( .A(n382), .B(n385), .Z(n383) );
  XOR U971 ( .A(n196), .B(n386), .Z(n198) );
  XNOR U972 ( .A(n387), .B(n388), .Z(n386) );
  ANDN U973 ( .B(n389), .A(n390), .Z(n387) );
  XNOR U974 ( .A(n391), .B(n392), .Z(n389) );
  IV U975 ( .A(n200), .Z(n196) );
  XOR U976 ( .A(n393), .B(n394), .Z(n200) );
  ANDN U977 ( .B(n395), .A(n396), .Z(n393) );
  XOR U978 ( .A(n397), .B(n394), .Z(n395) );
  XOR U979 ( .A(n398), .B(n399), .Z(n207) );
  ANDN U980 ( .B(n400), .A(n25), .Z(n398) );
  XOR U981 ( .A(n399), .B(n26), .Z(n400) );
  XNOR U982 ( .A(n401), .B(n402), .Z(n214) );
  ANDN U983 ( .B(n403), .A(n404), .Z(n401) );
  XNOR U984 ( .A(n402), .B(n405), .Z(n403) );
  XOR U985 ( .A(n210), .B(n406), .Z(n212) );
  XNOR U986 ( .A(n407), .B(n408), .Z(n406) );
  ANDN U987 ( .B(n409), .A(n410), .Z(n407) );
  XNOR U988 ( .A(n411), .B(n412), .Z(n409) );
  IV U989 ( .A(n213), .Z(n210) );
  XOR U990 ( .A(n413), .B(n414), .Z(n213) );
  ANDN U991 ( .B(n415), .A(n416), .Z(n413) );
  XOR U992 ( .A(n414), .B(n417), .Z(n415) );
  XNOR U993 ( .A(n220), .B(n419), .Z(n418) );
  IV U994 ( .A(n223), .Z(n419) );
  XOR U995 ( .A(n420), .B(n421), .Z(n223) );
  ANDN U996 ( .B(n422), .A(n423), .Z(n420) );
  XOR U997 ( .A(n421), .B(n424), .Z(n422) );
  XOR U998 ( .A(n425), .B(n426), .Z(n220) );
  ANDN U999 ( .B(n427), .A(n428), .Z(n425) );
  XNOR U1000 ( .A(n426), .B(n429), .Z(n427) );
  XOR U1001 ( .A(n217), .B(n430), .Z(n219) );
  XNOR U1002 ( .A(n431), .B(n432), .Z(n430) );
  ANDN U1003 ( .B(n433), .A(n434), .Z(n431) );
  XNOR U1004 ( .A(n435), .B(n436), .Z(n433) );
  IV U1005 ( .A(n221), .Z(n217) );
  XOR U1006 ( .A(n437), .B(n438), .Z(n221) );
  ANDN U1007 ( .B(n439), .A(n440), .Z(n437) );
  XOR U1008 ( .A(n441), .B(n438), .Z(n439) );
  XOR U1009 ( .A(n250), .B(n443), .Z(n442) );
  IV U1010 ( .A(n230), .Z(n443) );
  XOR U1011 ( .A(n444), .B(n445), .Z(n230) );
  ANDN U1012 ( .B(n446), .A(n447), .Z(n444) );
  XOR U1013 ( .A(n445), .B(n448), .Z(n446) );
  XNOR U1014 ( .A(n449), .B(n450), .Z(n238) );
  ANDN U1015 ( .B(n451), .A(n452), .Z(n449) );
  XNOR U1016 ( .A(n450), .B(n453), .Z(n451) );
  XNOR U1017 ( .A(n455), .B(n456), .Z(n454) );
  ANDN U1018 ( .B(n457), .A(n458), .Z(n455) );
  XNOR U1019 ( .A(n459), .B(n460), .Z(n457) );
  XOR U1020 ( .A(n461), .B(n462), .Z(n235) );
  ANDN U1021 ( .B(n463), .A(n464), .Z(n461) );
  XOR U1022 ( .A(n462), .B(n465), .Z(n463) );
  XNOR U1023 ( .A(n244), .B(n467), .Z(n466) );
  IV U1024 ( .A(n247), .Z(n467) );
  XOR U1025 ( .A(n468), .B(n469), .Z(n247) );
  ANDN U1026 ( .B(n470), .A(n471), .Z(n468) );
  XOR U1027 ( .A(n472), .B(n469), .Z(n470) );
  XOR U1028 ( .A(n473), .B(n474), .Z(n244) );
  ANDN U1029 ( .B(n475), .A(n476), .Z(n473) );
  XNOR U1030 ( .A(n474), .B(n477), .Z(n475) );
  XOR U1031 ( .A(n241), .B(n478), .Z(n243) );
  XNOR U1032 ( .A(n479), .B(n480), .Z(n478) );
  ANDN U1033 ( .B(n481), .A(n482), .Z(n479) );
  XNOR U1034 ( .A(n483), .B(n484), .Z(n481) );
  IV U1035 ( .A(n245), .Z(n241) );
  XOR U1036 ( .A(n485), .B(n486), .Z(n245) );
  ANDN U1037 ( .B(n487), .A(n488), .Z(n485) );
  XOR U1038 ( .A(n489), .B(n486), .Z(n487) );
  XOR U1039 ( .A(n282), .B(n491), .Z(n490) );
  IV U1040 ( .A(n254), .Z(n491) );
  XOR U1041 ( .A(n492), .B(n493), .Z(n254) );
  ANDN U1042 ( .B(n494), .A(n495), .Z(n492) );
  XOR U1043 ( .A(n493), .B(n496), .Z(n494) );
  XNOR U1044 ( .A(n497), .B(n498), .Z(n263) );
  ANDN U1045 ( .B(n499), .A(n500), .Z(n497) );
  XNOR U1046 ( .A(n498), .B(n501), .Z(n499) );
  XOR U1047 ( .A(n259), .B(n502), .Z(n261) );
  XNOR U1048 ( .A(n503), .B(n504), .Z(n502) );
  ANDN U1049 ( .B(n505), .A(n506), .Z(n503) );
  XNOR U1050 ( .A(n507), .B(n508), .Z(n505) );
  IV U1051 ( .A(n262), .Z(n259) );
  XOR U1052 ( .A(n509), .B(n510), .Z(n262) );
  ANDN U1053 ( .B(n511), .A(n512), .Z(n509) );
  XOR U1054 ( .A(n510), .B(n513), .Z(n511) );
  XNOR U1055 ( .A(n269), .B(n515), .Z(n514) );
  IV U1056 ( .A(n272), .Z(n515) );
  XOR U1057 ( .A(n516), .B(n517), .Z(n272) );
  ANDN U1058 ( .B(n518), .A(n519), .Z(n516) );
  XOR U1059 ( .A(n517), .B(n520), .Z(n518) );
  XOR U1060 ( .A(n521), .B(n522), .Z(n269) );
  ANDN U1061 ( .B(n523), .A(n524), .Z(n521) );
  XNOR U1062 ( .A(n522), .B(n525), .Z(n523) );
  XOR U1063 ( .A(n266), .B(n526), .Z(n268) );
  XNOR U1064 ( .A(n527), .B(n528), .Z(n526) );
  ANDN U1065 ( .B(n529), .A(n530), .Z(n527) );
  XNOR U1066 ( .A(n531), .B(n532), .Z(n529) );
  IV U1067 ( .A(n270), .Z(n266) );
  XOR U1068 ( .A(n533), .B(n534), .Z(n270) );
  ANDN U1069 ( .B(n535), .A(n536), .Z(n533) );
  XOR U1070 ( .A(n537), .B(n534), .Z(n535) );
  XOR U1071 ( .A(n299), .B(n539), .Z(n538) );
  IV U1072 ( .A(n279), .Z(n539) );
  XOR U1073 ( .A(n540), .B(n541), .Z(n279) );
  ANDN U1074 ( .B(n542), .A(n543), .Z(n540) );
  XOR U1075 ( .A(n544), .B(n541), .Z(n542) );
  XNOR U1076 ( .A(n545), .B(n546), .Z(n287) );
  ANDN U1077 ( .B(n547), .A(n548), .Z(n545) );
  XNOR U1078 ( .A(n546), .B(n549), .Z(n547) );
  XNOR U1079 ( .A(n551), .B(n552), .Z(n550) );
  ANDN U1080 ( .B(n553), .A(n554), .Z(n551) );
  XNOR U1081 ( .A(n555), .B(n556), .Z(n553) );
  XOR U1082 ( .A(n557), .B(n558), .Z(n284) );
  ANDN U1083 ( .B(n559), .A(n560), .Z(n557) );
  XOR U1084 ( .A(n558), .B(n561), .Z(n559) );
  XNOR U1085 ( .A(n293), .B(n563), .Z(n562) );
  IV U1086 ( .A(n296), .Z(n563) );
  XOR U1087 ( .A(n564), .B(n565), .Z(n296) );
  ANDN U1088 ( .B(n566), .A(n567), .Z(n564) );
  XOR U1089 ( .A(n568), .B(n565), .Z(n566) );
  XOR U1090 ( .A(n569), .B(n570), .Z(n293) );
  ANDN U1091 ( .B(n571), .A(n572), .Z(n569) );
  XNOR U1092 ( .A(n570), .B(n573), .Z(n571) );
  XOR U1093 ( .A(n290), .B(n574), .Z(n292) );
  XNOR U1094 ( .A(n575), .B(n576), .Z(n574) );
  ANDN U1095 ( .B(n577), .A(n578), .Z(n575) );
  XNOR U1096 ( .A(n579), .B(n580), .Z(n577) );
  IV U1097 ( .A(n294), .Z(n290) );
  XOR U1098 ( .A(n581), .B(n582), .Z(n294) );
  ANDN U1099 ( .B(n583), .A(n584), .Z(n581) );
  XOR U1100 ( .A(n585), .B(n582), .Z(n583) );
  XOR U1101 ( .A(n355), .B(n587), .Z(n586) );
  IV U1102 ( .A(n303), .Z(n587) );
  XOR U1103 ( .A(n588), .B(n589), .Z(n303) );
  ANDN U1104 ( .B(n590), .A(n591), .Z(n588) );
  XOR U1105 ( .A(n589), .B(n592), .Z(n590) );
  XNOR U1106 ( .A(n593), .B(n594), .Z(n312) );
  ANDN U1107 ( .B(n595), .A(n596), .Z(n593) );
  XNOR U1108 ( .A(n594), .B(n597), .Z(n595) );
  XOR U1109 ( .A(n308), .B(n598), .Z(n310) );
  XNOR U1110 ( .A(n599), .B(n600), .Z(n598) );
  ANDN U1111 ( .B(n601), .A(n602), .Z(n599) );
  XNOR U1112 ( .A(n603), .B(n604), .Z(n601) );
  IV U1113 ( .A(n311), .Z(n308) );
  XOR U1114 ( .A(n605), .B(n606), .Z(n311) );
  ANDN U1115 ( .B(n607), .A(n608), .Z(n605) );
  XOR U1116 ( .A(n606), .B(n609), .Z(n607) );
  XNOR U1117 ( .A(n318), .B(n611), .Z(n610) );
  IV U1118 ( .A(n321), .Z(n611) );
  XOR U1119 ( .A(n612), .B(n613), .Z(n321) );
  ANDN U1120 ( .B(n614), .A(n615), .Z(n612) );
  XOR U1121 ( .A(n613), .B(n616), .Z(n614) );
  XOR U1122 ( .A(n617), .B(n618), .Z(n318) );
  ANDN U1123 ( .B(n619), .A(n620), .Z(n617) );
  XNOR U1124 ( .A(n618), .B(n621), .Z(n619) );
  XOR U1125 ( .A(n315), .B(n622), .Z(n317) );
  XNOR U1126 ( .A(n623), .B(n624), .Z(n622) );
  ANDN U1127 ( .B(n625), .A(n626), .Z(n623) );
  XNOR U1128 ( .A(n627), .B(n628), .Z(n625) );
  IV U1129 ( .A(n319), .Z(n315) );
  XOR U1130 ( .A(n629), .B(n630), .Z(n319) );
  ANDN U1131 ( .B(n631), .A(n632), .Z(n629) );
  XOR U1132 ( .A(n633), .B(n630), .Z(n631) );
  XOR U1133 ( .A(n348), .B(n635), .Z(n634) );
  IV U1134 ( .A(n328), .Z(n635) );
  XOR U1135 ( .A(n636), .B(n637), .Z(n328) );
  ANDN U1136 ( .B(n638), .A(n639), .Z(n636) );
  XOR U1137 ( .A(n637), .B(n640), .Z(n638) );
  XNOR U1138 ( .A(n641), .B(n642), .Z(n336) );
  ANDN U1139 ( .B(n643), .A(n644), .Z(n641) );
  XNOR U1140 ( .A(n642), .B(n645), .Z(n643) );
  XNOR U1141 ( .A(n647), .B(n648), .Z(n646) );
  ANDN U1142 ( .B(n649), .A(n650), .Z(n647) );
  XNOR U1143 ( .A(n651), .B(n652), .Z(n649) );
  XOR U1144 ( .A(n653), .B(n654), .Z(n333) );
  ANDN U1145 ( .B(n655), .A(n656), .Z(n653) );
  XOR U1146 ( .A(n654), .B(n657), .Z(n655) );
  XNOR U1147 ( .A(n342), .B(n659), .Z(n658) );
  IV U1148 ( .A(n345), .Z(n659) );
  XOR U1149 ( .A(n660), .B(n661), .Z(n345) );
  ANDN U1150 ( .B(n662), .A(n663), .Z(n660) );
  XOR U1151 ( .A(n664), .B(n661), .Z(n662) );
  XOR U1152 ( .A(n665), .B(n666), .Z(n342) );
  ANDN U1153 ( .B(n667), .A(n668), .Z(n665) );
  XNOR U1154 ( .A(n666), .B(n669), .Z(n667) );
  XOR U1155 ( .A(n339), .B(n670), .Z(n341) );
  XNOR U1156 ( .A(n671), .B(n672), .Z(n670) );
  ANDN U1157 ( .B(n673), .A(n674), .Z(n671) );
  XNOR U1158 ( .A(n675), .B(n676), .Z(n673) );
  IV U1159 ( .A(n343), .Z(n339) );
  XOR U1160 ( .A(n677), .B(n678), .Z(n343) );
  ANDN U1161 ( .B(n679), .A(n680), .Z(n677) );
  XOR U1162 ( .A(n681), .B(n678), .Z(n679) );
  XOR U1163 ( .A(n380), .B(n683), .Z(n682) );
  IV U1164 ( .A(n352), .Z(n683) );
  XOR U1165 ( .A(n684), .B(n685), .Z(n352) );
  ANDN U1166 ( .B(n686), .A(n687), .Z(n684) );
  XOR U1167 ( .A(n688), .B(n685), .Z(n686) );
  XNOR U1168 ( .A(n689), .B(n690), .Z(n361) );
  ANDN U1169 ( .B(n691), .A(n692), .Z(n689) );
  XNOR U1170 ( .A(n690), .B(n693), .Z(n691) );
  XOR U1171 ( .A(n357), .B(n694), .Z(n359) );
  XNOR U1172 ( .A(n695), .B(n696), .Z(n694) );
  ANDN U1173 ( .B(n697), .A(n698), .Z(n695) );
  XNOR U1174 ( .A(n699), .B(n700), .Z(n697) );
  IV U1175 ( .A(n360), .Z(n357) );
  XOR U1176 ( .A(n701), .B(n702), .Z(n360) );
  ANDN U1177 ( .B(n703), .A(n704), .Z(n701) );
  XOR U1178 ( .A(n702), .B(n705), .Z(n703) );
  XOR U1179 ( .A(n706), .B(n707), .Z(n372) );
  XNOR U1180 ( .A(n367), .B(n708), .Z(n707) );
  IV U1181 ( .A(n370), .Z(n708) );
  XOR U1182 ( .A(n709), .B(n710), .Z(n370) );
  ANDN U1183 ( .B(n711), .A(n712), .Z(n709) );
  XOR U1184 ( .A(n710), .B(n713), .Z(n711) );
  XOR U1185 ( .A(n714), .B(n715), .Z(n367) );
  ANDN U1186 ( .B(n716), .A(n717), .Z(n714) );
  XNOR U1187 ( .A(n715), .B(n718), .Z(n716) );
  IV U1188 ( .A(n366), .Z(n706) );
  XOR U1189 ( .A(n364), .B(n719), .Z(n366) );
  XNOR U1190 ( .A(n720), .B(n721), .Z(n719) );
  ANDN U1191 ( .B(n722), .A(n723), .Z(n720) );
  XNOR U1192 ( .A(n724), .B(n725), .Z(n722) );
  IV U1193 ( .A(n368), .Z(n364) );
  XOR U1194 ( .A(n726), .B(n727), .Z(n368) );
  ANDN U1195 ( .B(n728), .A(n729), .Z(n726) );
  XOR U1196 ( .A(n730), .B(n727), .Z(n728) );
  XOR U1197 ( .A(n397), .B(n732), .Z(n731) );
  IV U1198 ( .A(n377), .Z(n732) );
  XOR U1199 ( .A(n733), .B(n734), .Z(n377) );
  ANDN U1200 ( .B(n735), .A(n736), .Z(n733) );
  XOR U1201 ( .A(n737), .B(n734), .Z(n735) );
  XNOR U1202 ( .A(n738), .B(n739), .Z(n385) );
  ANDN U1203 ( .B(n740), .A(n741), .Z(n738) );
  XNOR U1204 ( .A(n739), .B(n742), .Z(n740) );
  XNOR U1205 ( .A(n744), .B(n745), .Z(n743) );
  ANDN U1206 ( .B(n746), .A(n747), .Z(n744) );
  XNOR U1207 ( .A(n748), .B(n749), .Z(n746) );
  XOR U1208 ( .A(n750), .B(n751), .Z(n382) );
  ANDN U1209 ( .B(n752), .A(n753), .Z(n750) );
  XOR U1210 ( .A(n751), .B(n754), .Z(n752) );
  XNOR U1211 ( .A(n391), .B(n756), .Z(n755) );
  IV U1212 ( .A(n394), .Z(n756) );
  XOR U1213 ( .A(n757), .B(n758), .Z(n394) );
  ANDN U1214 ( .B(n759), .A(n760), .Z(n757) );
  XOR U1215 ( .A(n761), .B(n758), .Z(n759) );
  XOR U1216 ( .A(n762), .B(n763), .Z(n391) );
  ANDN U1217 ( .B(n764), .A(n765), .Z(n762) );
  XNOR U1218 ( .A(n763), .B(n766), .Z(n764) );
  XOR U1219 ( .A(n388), .B(n767), .Z(n390) );
  XNOR U1220 ( .A(n768), .B(n769), .Z(n767) );
  ANDN U1221 ( .B(n770), .A(n771), .Z(n768) );
  XNOR U1222 ( .A(n772), .B(n773), .Z(n770) );
  IV U1223 ( .A(n392), .Z(n388) );
  XOR U1224 ( .A(n774), .B(n775), .Z(n392) );
  ANDN U1225 ( .B(n776), .A(n777), .Z(n774) );
  XOR U1226 ( .A(n778), .B(n775), .Z(n776) );
  XOR U1227 ( .A(n779), .B(n780), .Z(n399) );
  ANDN U1228 ( .B(n781), .A(n27), .Z(n779) );
  XOR U1229 ( .A(n780), .B(n28), .Z(n781) );
  XNOR U1230 ( .A(n782), .B(n783), .Z(n405) );
  NANDN U1231 ( .A(n784), .B(n785), .Z(n783) );
  NANDN U1232 ( .A(n786), .B(n782), .Z(n785) );
  XNOR U1233 ( .A(n787), .B(n402), .Z(n404) );
  XNOR U1234 ( .A(n788), .B(n789), .Z(n402) );
  NAND U1235 ( .A(n790), .B(n791), .Z(n789) );
  XNOR U1236 ( .A(n788), .B(n792), .Z(n790) );
  NOR U1237 ( .A(n793), .B(n794), .Z(n787) );
  XOR U1238 ( .A(n411), .B(n414), .Z(n795) );
  XNOR U1239 ( .A(n796), .B(n797), .Z(n414) );
  NANDN U1240 ( .A(n798), .B(n799), .Z(n797) );
  XOR U1241 ( .A(n796), .B(n800), .Z(n799) );
  XNOR U1242 ( .A(n801), .B(n802), .Z(n411) );
  NANDN U1243 ( .A(n803), .B(n804), .Z(n802) );
  NANDN U1244 ( .A(n801), .B(n805), .Z(n804) );
  XOR U1245 ( .A(n806), .B(n412), .Z(n410) );
  IV U1246 ( .A(n408), .Z(n412) );
  XNOR U1247 ( .A(n807), .B(n808), .Z(n408) );
  NAND U1248 ( .A(n809), .B(n810), .Z(n808) );
  XOR U1249 ( .A(n807), .B(n811), .Z(n809) );
  NOR U1250 ( .A(n812), .B(n813), .Z(n806) );
  XNOR U1251 ( .A(n441), .B(n421), .Z(n814) );
  XNOR U1252 ( .A(n815), .B(n816), .Z(n421) );
  NANDN U1253 ( .A(n817), .B(n818), .Z(n816) );
  XOR U1254 ( .A(n815), .B(n819), .Z(n818) );
  XNOR U1255 ( .A(n820), .B(n821), .Z(n429) );
  NANDN U1256 ( .A(n822), .B(n823), .Z(n821) );
  NANDN U1257 ( .A(n824), .B(n820), .Z(n823) );
  XNOR U1258 ( .A(n825), .B(n426), .Z(n428) );
  XNOR U1259 ( .A(n826), .B(n827), .Z(n426) );
  NAND U1260 ( .A(n828), .B(n829), .Z(n827) );
  XNOR U1261 ( .A(n826), .B(n830), .Z(n828) );
  NOR U1262 ( .A(n831), .B(n832), .Z(n825) );
  XOR U1263 ( .A(n435), .B(n438), .Z(n833) );
  XNOR U1264 ( .A(n834), .B(n835), .Z(n438) );
  NANDN U1265 ( .A(n836), .B(n837), .Z(n835) );
  XNOR U1266 ( .A(n834), .B(n838), .Z(n837) );
  XNOR U1267 ( .A(n839), .B(n840), .Z(n435) );
  NANDN U1268 ( .A(n841), .B(n842), .Z(n840) );
  NANDN U1269 ( .A(n839), .B(n843), .Z(n842) );
  XOR U1270 ( .A(n844), .B(n436), .Z(n434) );
  IV U1271 ( .A(n432), .Z(n436) );
  XNOR U1272 ( .A(n845), .B(n846), .Z(n432) );
  NAND U1273 ( .A(n847), .B(n848), .Z(n846) );
  XOR U1274 ( .A(n845), .B(n849), .Z(n847) );
  NOR U1275 ( .A(n850), .B(n851), .Z(n844) );
  XNOR U1276 ( .A(n472), .B(n445), .Z(n852) );
  XNOR U1277 ( .A(n853), .B(n854), .Z(n445) );
  NANDN U1278 ( .A(n855), .B(n856), .Z(n854) );
  XOR U1279 ( .A(n853), .B(n857), .Z(n856) );
  XNOR U1280 ( .A(n858), .B(n859), .Z(n453) );
  NANDN U1281 ( .A(n860), .B(n861), .Z(n859) );
  NANDN U1282 ( .A(n862), .B(n858), .Z(n861) );
  XNOR U1283 ( .A(n863), .B(n450), .Z(n452) );
  XNOR U1284 ( .A(n864), .B(n865), .Z(n450) );
  NAND U1285 ( .A(n866), .B(n867), .Z(n865) );
  XNOR U1286 ( .A(n864), .B(n868), .Z(n866) );
  NOR U1287 ( .A(n869), .B(n870), .Z(n863) );
  XOR U1288 ( .A(n459), .B(n462), .Z(n871) );
  XNOR U1289 ( .A(n872), .B(n873), .Z(n462) );
  NANDN U1290 ( .A(n874), .B(n875), .Z(n873) );
  XOR U1291 ( .A(n872), .B(n876), .Z(n875) );
  XNOR U1292 ( .A(n877), .B(n878), .Z(n459) );
  NANDN U1293 ( .A(n879), .B(n880), .Z(n878) );
  NANDN U1294 ( .A(n877), .B(n881), .Z(n880) );
  XOR U1295 ( .A(n882), .B(n460), .Z(n458) );
  IV U1296 ( .A(n456), .Z(n460) );
  XNOR U1297 ( .A(n883), .B(n884), .Z(n456) );
  NAND U1298 ( .A(n885), .B(n886), .Z(n884) );
  XOR U1299 ( .A(n883), .B(n887), .Z(n885) );
  NOR U1300 ( .A(n888), .B(n889), .Z(n882) );
  XNOR U1301 ( .A(n489), .B(n469), .Z(n890) );
  XNOR U1302 ( .A(n891), .B(n892), .Z(n469) );
  NANDN U1303 ( .A(n893), .B(n894), .Z(n892) );
  XOR U1304 ( .A(n891), .B(n895), .Z(n894) );
  XNOR U1305 ( .A(n896), .B(n897), .Z(n477) );
  NANDN U1306 ( .A(n898), .B(n899), .Z(n897) );
  NANDN U1307 ( .A(n900), .B(n896), .Z(n899) );
  XNOR U1308 ( .A(n901), .B(n474), .Z(n476) );
  XNOR U1309 ( .A(n902), .B(n903), .Z(n474) );
  NAND U1310 ( .A(n904), .B(n905), .Z(n903) );
  XNOR U1311 ( .A(n902), .B(n906), .Z(n904) );
  NOR U1312 ( .A(n907), .B(n908), .Z(n901) );
  XOR U1313 ( .A(n483), .B(n486), .Z(n909) );
  XNOR U1314 ( .A(n910), .B(n911), .Z(n486) );
  NANDN U1315 ( .A(n912), .B(n913), .Z(n911) );
  XNOR U1316 ( .A(n910), .B(n914), .Z(n913) );
  XNOR U1317 ( .A(n915), .B(n916), .Z(n483) );
  NANDN U1318 ( .A(n917), .B(n918), .Z(n916) );
  NANDN U1319 ( .A(n915), .B(n919), .Z(n918) );
  XOR U1320 ( .A(n920), .B(n484), .Z(n482) );
  IV U1321 ( .A(n480), .Z(n484) );
  XNOR U1322 ( .A(n921), .B(n922), .Z(n480) );
  NAND U1323 ( .A(n923), .B(n924), .Z(n922) );
  XOR U1324 ( .A(n921), .B(n925), .Z(n923) );
  NOR U1325 ( .A(n926), .B(n927), .Z(n920) );
  XNOR U1326 ( .A(n544), .B(n493), .Z(n928) );
  XNOR U1327 ( .A(n929), .B(n930), .Z(n493) );
  NANDN U1328 ( .A(n931), .B(n932), .Z(n930) );
  XOR U1329 ( .A(n929), .B(n933), .Z(n932) );
  XNOR U1330 ( .A(n934), .B(n935), .Z(n501) );
  NANDN U1331 ( .A(n936), .B(n937), .Z(n935) );
  NANDN U1332 ( .A(n938), .B(n934), .Z(n937) );
  XNOR U1333 ( .A(n939), .B(n498), .Z(n500) );
  XNOR U1334 ( .A(n940), .B(n941), .Z(n498) );
  NAND U1335 ( .A(n942), .B(n943), .Z(n941) );
  XNOR U1336 ( .A(n940), .B(n944), .Z(n942) );
  NOR U1337 ( .A(n945), .B(n946), .Z(n939) );
  XOR U1338 ( .A(n507), .B(n510), .Z(n947) );
  XNOR U1339 ( .A(n948), .B(n949), .Z(n510) );
  NANDN U1340 ( .A(n950), .B(n951), .Z(n949) );
  XOR U1341 ( .A(n948), .B(n952), .Z(n951) );
  XNOR U1342 ( .A(n953), .B(n954), .Z(n507) );
  NANDN U1343 ( .A(n955), .B(n956), .Z(n954) );
  NANDN U1344 ( .A(n953), .B(n957), .Z(n956) );
  XOR U1345 ( .A(n958), .B(n508), .Z(n506) );
  IV U1346 ( .A(n504), .Z(n508) );
  XNOR U1347 ( .A(n959), .B(n960), .Z(n504) );
  NAND U1348 ( .A(n961), .B(n962), .Z(n960) );
  XOR U1349 ( .A(n959), .B(n963), .Z(n961) );
  NOR U1350 ( .A(n964), .B(n965), .Z(n958) );
  XNOR U1351 ( .A(n537), .B(n517), .Z(n966) );
  XNOR U1352 ( .A(n967), .B(n968), .Z(n517) );
  NANDN U1353 ( .A(n969), .B(n970), .Z(n968) );
  XOR U1354 ( .A(n967), .B(n971), .Z(n970) );
  XNOR U1355 ( .A(n972), .B(n973), .Z(n525) );
  NANDN U1356 ( .A(n974), .B(n975), .Z(n973) );
  NANDN U1357 ( .A(n976), .B(n972), .Z(n975) );
  XNOR U1358 ( .A(n977), .B(n522), .Z(n524) );
  XNOR U1359 ( .A(n978), .B(n979), .Z(n522) );
  NAND U1360 ( .A(n980), .B(n981), .Z(n979) );
  XNOR U1361 ( .A(n978), .B(n982), .Z(n980) );
  NOR U1362 ( .A(n983), .B(n984), .Z(n977) );
  XOR U1363 ( .A(n531), .B(n534), .Z(n985) );
  XNOR U1364 ( .A(n986), .B(n987), .Z(n534) );
  NANDN U1365 ( .A(n988), .B(n989), .Z(n987) );
  XNOR U1366 ( .A(n986), .B(n990), .Z(n989) );
  XNOR U1367 ( .A(n991), .B(n992), .Z(n531) );
  NANDN U1368 ( .A(n993), .B(n994), .Z(n992) );
  NANDN U1369 ( .A(n991), .B(n995), .Z(n994) );
  XOR U1370 ( .A(n996), .B(n532), .Z(n530) );
  IV U1371 ( .A(n528), .Z(n532) );
  XNOR U1372 ( .A(n997), .B(n998), .Z(n528) );
  NAND U1373 ( .A(n999), .B(n1000), .Z(n998) );
  XOR U1374 ( .A(n997), .B(n1001), .Z(n999) );
  NOR U1375 ( .A(n1002), .B(n1003), .Z(n996) );
  XNOR U1376 ( .A(n568), .B(n541), .Z(n1004) );
  XNOR U1377 ( .A(n1005), .B(n1006), .Z(n541) );
  NANDN U1378 ( .A(n1007), .B(n1008), .Z(n1006) );
  XOR U1379 ( .A(n1005), .B(n1009), .Z(n1008) );
  XNOR U1380 ( .A(n1010), .B(n1011), .Z(n549) );
  NANDN U1381 ( .A(n1012), .B(n1013), .Z(n1011) );
  NANDN U1382 ( .A(n1014), .B(n1010), .Z(n1013) );
  XNOR U1383 ( .A(n1015), .B(n546), .Z(n548) );
  XNOR U1384 ( .A(n1016), .B(n1017), .Z(n546) );
  NAND U1385 ( .A(n1018), .B(n1019), .Z(n1017) );
  XNOR U1386 ( .A(n1016), .B(n1020), .Z(n1018) );
  NOR U1387 ( .A(n1021), .B(n1022), .Z(n1015) );
  XOR U1388 ( .A(n555), .B(n558), .Z(n1023) );
  XNOR U1389 ( .A(n1024), .B(n1025), .Z(n558) );
  NANDN U1390 ( .A(n1026), .B(n1027), .Z(n1025) );
  XOR U1391 ( .A(n1024), .B(n1028), .Z(n1027) );
  XNOR U1392 ( .A(n1029), .B(n1030), .Z(n555) );
  NANDN U1393 ( .A(n1031), .B(n1032), .Z(n1030) );
  NANDN U1394 ( .A(n1029), .B(n1033), .Z(n1032) );
  XOR U1395 ( .A(n1034), .B(n556), .Z(n554) );
  IV U1396 ( .A(n552), .Z(n556) );
  XNOR U1397 ( .A(n1035), .B(n1036), .Z(n552) );
  NAND U1398 ( .A(n1037), .B(n1038), .Z(n1036) );
  XOR U1399 ( .A(n1035), .B(n1039), .Z(n1037) );
  NOR U1400 ( .A(n1040), .B(n1041), .Z(n1034) );
  XNOR U1401 ( .A(n585), .B(n565), .Z(n1042) );
  XNOR U1402 ( .A(n1043), .B(n1044), .Z(n565) );
  NANDN U1403 ( .A(n1045), .B(n1046), .Z(n1044) );
  XOR U1404 ( .A(n1043), .B(n1047), .Z(n1046) );
  XNOR U1405 ( .A(n1048), .B(n1049), .Z(n573) );
  NANDN U1406 ( .A(n1050), .B(n1051), .Z(n1049) );
  NANDN U1407 ( .A(n1052), .B(n1048), .Z(n1051) );
  XNOR U1408 ( .A(n1053), .B(n570), .Z(n572) );
  XNOR U1409 ( .A(n1054), .B(n1055), .Z(n570) );
  NAND U1410 ( .A(n1056), .B(n1057), .Z(n1055) );
  XNOR U1411 ( .A(n1054), .B(n1058), .Z(n1056) );
  NOR U1412 ( .A(n1059), .B(n1060), .Z(n1053) );
  XOR U1413 ( .A(n579), .B(n582), .Z(n1061) );
  XNOR U1414 ( .A(n1062), .B(n1063), .Z(n582) );
  NANDN U1415 ( .A(n1064), .B(n1065), .Z(n1063) );
  XNOR U1416 ( .A(n1062), .B(n1066), .Z(n1065) );
  XNOR U1417 ( .A(n1067), .B(n1068), .Z(n579) );
  NANDN U1418 ( .A(n1069), .B(n1070), .Z(n1068) );
  NANDN U1419 ( .A(n1067), .B(n1071), .Z(n1070) );
  XOR U1420 ( .A(n1072), .B(n580), .Z(n578) );
  IV U1421 ( .A(n576), .Z(n580) );
  XNOR U1422 ( .A(n1073), .B(n1074), .Z(n576) );
  NAND U1423 ( .A(n1075), .B(n1076), .Z(n1074) );
  XOR U1424 ( .A(n1073), .B(n1077), .Z(n1075) );
  NOR U1425 ( .A(n1078), .B(n1079), .Z(n1072) );
  XNOR U1426 ( .A(n688), .B(n589), .Z(n1080) );
  XNOR U1427 ( .A(n1081), .B(n1082), .Z(n589) );
  NANDN U1428 ( .A(n1083), .B(n1084), .Z(n1082) );
  XOR U1429 ( .A(n1081), .B(n1085), .Z(n1084) );
  XNOR U1430 ( .A(n1086), .B(n1087), .Z(n597) );
  NANDN U1431 ( .A(n1088), .B(n1089), .Z(n1087) );
  NANDN U1432 ( .A(n1090), .B(n1086), .Z(n1089) );
  XNOR U1433 ( .A(n1091), .B(n594), .Z(n596) );
  XNOR U1434 ( .A(n1092), .B(n1093), .Z(n594) );
  NAND U1435 ( .A(n1094), .B(n1095), .Z(n1093) );
  XNOR U1436 ( .A(n1092), .B(n1096), .Z(n1094) );
  NOR U1437 ( .A(n1097), .B(n1098), .Z(n1091) );
  XOR U1438 ( .A(n603), .B(n606), .Z(n1099) );
  XNOR U1439 ( .A(n1100), .B(n1101), .Z(n606) );
  NANDN U1440 ( .A(n1102), .B(n1103), .Z(n1101) );
  XOR U1441 ( .A(n1100), .B(n1104), .Z(n1103) );
  XNOR U1442 ( .A(n1105), .B(n1106), .Z(n603) );
  NANDN U1443 ( .A(n1107), .B(n1108), .Z(n1106) );
  NANDN U1444 ( .A(n1105), .B(n1109), .Z(n1108) );
  XOR U1445 ( .A(n1110), .B(n604), .Z(n602) );
  IV U1446 ( .A(n600), .Z(n604) );
  XNOR U1447 ( .A(n1111), .B(n1112), .Z(n600) );
  NAND U1448 ( .A(n1113), .B(n1114), .Z(n1112) );
  XOR U1449 ( .A(n1111), .B(n1115), .Z(n1113) );
  NOR U1450 ( .A(n1116), .B(n1117), .Z(n1110) );
  XNOR U1451 ( .A(n633), .B(n613), .Z(n1118) );
  XNOR U1452 ( .A(n1119), .B(n1120), .Z(n613) );
  NANDN U1453 ( .A(n1121), .B(n1122), .Z(n1120) );
  XOR U1454 ( .A(n1119), .B(n1123), .Z(n1122) );
  XNOR U1455 ( .A(n1124), .B(n1125), .Z(n621) );
  NANDN U1456 ( .A(n1126), .B(n1127), .Z(n1125) );
  NANDN U1457 ( .A(n1128), .B(n1124), .Z(n1127) );
  XNOR U1458 ( .A(n1129), .B(n618), .Z(n620) );
  XNOR U1459 ( .A(n1130), .B(n1131), .Z(n618) );
  NAND U1460 ( .A(n1132), .B(n1133), .Z(n1131) );
  XNOR U1461 ( .A(n1130), .B(n1134), .Z(n1132) );
  NOR U1462 ( .A(n1135), .B(n1136), .Z(n1129) );
  XOR U1463 ( .A(n627), .B(n630), .Z(n1137) );
  XNOR U1464 ( .A(n1138), .B(n1139), .Z(n630) );
  NANDN U1465 ( .A(n1140), .B(n1141), .Z(n1139) );
  XNOR U1466 ( .A(n1138), .B(n1142), .Z(n1141) );
  XNOR U1467 ( .A(n1143), .B(n1144), .Z(n627) );
  NANDN U1468 ( .A(n1145), .B(n1146), .Z(n1144) );
  NANDN U1469 ( .A(n1143), .B(n1147), .Z(n1146) );
  XOR U1470 ( .A(n1148), .B(n628), .Z(n626) );
  IV U1471 ( .A(n624), .Z(n628) );
  XNOR U1472 ( .A(n1149), .B(n1150), .Z(n624) );
  NAND U1473 ( .A(n1151), .B(n1152), .Z(n1150) );
  XOR U1474 ( .A(n1149), .B(n1153), .Z(n1151) );
  NOR U1475 ( .A(n1154), .B(n1155), .Z(n1148) );
  XNOR U1476 ( .A(n664), .B(n637), .Z(n1156) );
  XNOR U1477 ( .A(n1157), .B(n1158), .Z(n637) );
  NANDN U1478 ( .A(n1159), .B(n1160), .Z(n1158) );
  XOR U1479 ( .A(n1157), .B(n1161), .Z(n1160) );
  XNOR U1480 ( .A(n1162), .B(n1163), .Z(n645) );
  NANDN U1481 ( .A(n1164), .B(n1165), .Z(n1163) );
  NANDN U1482 ( .A(n1166), .B(n1162), .Z(n1165) );
  XNOR U1483 ( .A(n1167), .B(n642), .Z(n644) );
  XNOR U1484 ( .A(n1168), .B(n1169), .Z(n642) );
  NAND U1485 ( .A(n1170), .B(n1171), .Z(n1169) );
  XNOR U1486 ( .A(n1168), .B(n1172), .Z(n1170) );
  NOR U1487 ( .A(n1173), .B(n1174), .Z(n1167) );
  XOR U1488 ( .A(n651), .B(n654), .Z(n1175) );
  XNOR U1489 ( .A(n1176), .B(n1177), .Z(n654) );
  NANDN U1490 ( .A(n1178), .B(n1179), .Z(n1177) );
  XOR U1491 ( .A(n1176), .B(n1180), .Z(n1179) );
  XNOR U1492 ( .A(n1181), .B(n1182), .Z(n651) );
  NANDN U1493 ( .A(n1183), .B(n1184), .Z(n1182) );
  NANDN U1494 ( .A(n1181), .B(n1185), .Z(n1184) );
  XOR U1495 ( .A(n1186), .B(n652), .Z(n650) );
  IV U1496 ( .A(n648), .Z(n652) );
  XNOR U1497 ( .A(n1187), .B(n1188), .Z(n648) );
  NAND U1498 ( .A(n1189), .B(n1190), .Z(n1188) );
  XOR U1499 ( .A(n1187), .B(n1191), .Z(n1189) );
  NOR U1500 ( .A(n1192), .B(n1193), .Z(n1186) );
  XNOR U1501 ( .A(n681), .B(n661), .Z(n1194) );
  XNOR U1502 ( .A(n1195), .B(n1196), .Z(n661) );
  NANDN U1503 ( .A(n1197), .B(n1198), .Z(n1196) );
  XOR U1504 ( .A(n1195), .B(n1199), .Z(n1198) );
  XNOR U1505 ( .A(n1200), .B(n1201), .Z(n669) );
  NANDN U1506 ( .A(n1202), .B(n1203), .Z(n1201) );
  NANDN U1507 ( .A(n1204), .B(n1200), .Z(n1203) );
  XNOR U1508 ( .A(n1205), .B(n666), .Z(n668) );
  XNOR U1509 ( .A(n1206), .B(n1207), .Z(n666) );
  NAND U1510 ( .A(n1208), .B(n1209), .Z(n1207) );
  XNOR U1511 ( .A(n1206), .B(n1210), .Z(n1208) );
  NOR U1512 ( .A(n1211), .B(n1212), .Z(n1205) );
  XOR U1513 ( .A(n675), .B(n678), .Z(n1213) );
  XNOR U1514 ( .A(n1214), .B(n1215), .Z(n678) );
  NANDN U1515 ( .A(n1216), .B(n1217), .Z(n1215) );
  XNOR U1516 ( .A(n1214), .B(n1218), .Z(n1217) );
  XNOR U1517 ( .A(n1219), .B(n1220), .Z(n675) );
  NANDN U1518 ( .A(n1221), .B(n1222), .Z(n1220) );
  NANDN U1519 ( .A(n1219), .B(n1223), .Z(n1222) );
  XOR U1520 ( .A(n1224), .B(n676), .Z(n674) );
  IV U1521 ( .A(n672), .Z(n676) );
  XNOR U1522 ( .A(n1225), .B(n1226), .Z(n672) );
  NAND U1523 ( .A(n1227), .B(n1228), .Z(n1226) );
  XOR U1524 ( .A(n1225), .B(n1229), .Z(n1227) );
  NOR U1525 ( .A(n1230), .B(n1231), .Z(n1224) );
  XNOR U1526 ( .A(n737), .B(n685), .Z(n1232) );
  XNOR U1527 ( .A(n1233), .B(n1234), .Z(n685) );
  NANDN U1528 ( .A(n1235), .B(n1236), .Z(n1234) );
  XOR U1529 ( .A(n1233), .B(n1237), .Z(n1236) );
  XNOR U1530 ( .A(n1238), .B(n1239), .Z(n693) );
  NANDN U1531 ( .A(n1240), .B(n1241), .Z(n1239) );
  NANDN U1532 ( .A(n1242), .B(n1238), .Z(n1241) );
  XNOR U1533 ( .A(n1243), .B(n690), .Z(n692) );
  XNOR U1534 ( .A(n1244), .B(n1245), .Z(n690) );
  NAND U1535 ( .A(n1246), .B(n1247), .Z(n1245) );
  XNOR U1536 ( .A(n1244), .B(n1248), .Z(n1246) );
  NOR U1537 ( .A(n1249), .B(n1250), .Z(n1243) );
  XOR U1538 ( .A(n699), .B(n702), .Z(n1251) );
  XNOR U1539 ( .A(n1252), .B(n1253), .Z(n702) );
  NANDN U1540 ( .A(n1254), .B(n1255), .Z(n1253) );
  XOR U1541 ( .A(n1252), .B(n1256), .Z(n1255) );
  XNOR U1542 ( .A(n1257), .B(n1258), .Z(n699) );
  NANDN U1543 ( .A(n1259), .B(n1260), .Z(n1258) );
  NANDN U1544 ( .A(n1257), .B(n1261), .Z(n1260) );
  XOR U1545 ( .A(n1262), .B(n700), .Z(n698) );
  IV U1546 ( .A(n696), .Z(n700) );
  XNOR U1547 ( .A(n1263), .B(n1264), .Z(n696) );
  NAND U1548 ( .A(n1265), .B(n1266), .Z(n1264) );
  XOR U1549 ( .A(n1263), .B(n1267), .Z(n1265) );
  NOR U1550 ( .A(n1268), .B(n1269), .Z(n1262) );
  XNOR U1551 ( .A(n730), .B(n710), .Z(n1270) );
  XNOR U1552 ( .A(n1271), .B(n1272), .Z(n710) );
  NANDN U1553 ( .A(n1273), .B(n1274), .Z(n1272) );
  XOR U1554 ( .A(n1271), .B(n1275), .Z(n1274) );
  XNOR U1555 ( .A(n1276), .B(n1277), .Z(n718) );
  NANDN U1556 ( .A(n1278), .B(n1279), .Z(n1277) );
  NANDN U1557 ( .A(n1280), .B(n1276), .Z(n1279) );
  XNOR U1558 ( .A(n1281), .B(n715), .Z(n717) );
  XNOR U1559 ( .A(n1282), .B(n1283), .Z(n715) );
  NAND U1560 ( .A(n1284), .B(n1285), .Z(n1283) );
  XNOR U1561 ( .A(n1282), .B(n1286), .Z(n1284) );
  NOR U1562 ( .A(n1287), .B(n1288), .Z(n1281) );
  XOR U1563 ( .A(n724), .B(n727), .Z(n1289) );
  XNOR U1564 ( .A(n1290), .B(n1291), .Z(n727) );
  NANDN U1565 ( .A(n1292), .B(n1293), .Z(n1291) );
  XNOR U1566 ( .A(n1290), .B(n1294), .Z(n1293) );
  XNOR U1567 ( .A(n1295), .B(n1296), .Z(n724) );
  NANDN U1568 ( .A(n1297), .B(n1298), .Z(n1296) );
  NANDN U1569 ( .A(n1295), .B(n1299), .Z(n1298) );
  XOR U1570 ( .A(n1300), .B(n725), .Z(n723) );
  IV U1571 ( .A(n721), .Z(n725) );
  XNOR U1572 ( .A(n1301), .B(n1302), .Z(n721) );
  NAND U1573 ( .A(n1303), .B(n1304), .Z(n1302) );
  XOR U1574 ( .A(n1301), .B(n1305), .Z(n1303) );
  NOR U1575 ( .A(n1306), .B(n1307), .Z(n1300) );
  XNOR U1576 ( .A(n761), .B(n734), .Z(n1308) );
  XNOR U1577 ( .A(n1309), .B(n1310), .Z(n734) );
  NANDN U1578 ( .A(n1311), .B(n1312), .Z(n1310) );
  XOR U1579 ( .A(n1309), .B(n1313), .Z(n1312) );
  XNOR U1580 ( .A(n1314), .B(n1315), .Z(n742) );
  NANDN U1581 ( .A(n1316), .B(n1317), .Z(n1315) );
  NANDN U1582 ( .A(n1318), .B(n1314), .Z(n1317) );
  XNOR U1583 ( .A(n1319), .B(n739), .Z(n741) );
  XNOR U1584 ( .A(n1320), .B(n1321), .Z(n739) );
  NAND U1585 ( .A(n1322), .B(n1323), .Z(n1321) );
  XNOR U1586 ( .A(n1320), .B(n1324), .Z(n1322) );
  NOR U1587 ( .A(n1325), .B(n1326), .Z(n1319) );
  XOR U1588 ( .A(n748), .B(n751), .Z(n1327) );
  XNOR U1589 ( .A(n1328), .B(n1329), .Z(n751) );
  NANDN U1590 ( .A(n1330), .B(n1331), .Z(n1329) );
  XOR U1591 ( .A(n1328), .B(n1332), .Z(n1331) );
  XNOR U1592 ( .A(n1333), .B(n1334), .Z(n748) );
  NANDN U1593 ( .A(n1335), .B(n1336), .Z(n1334) );
  NANDN U1594 ( .A(n1333), .B(n1337), .Z(n1336) );
  XOR U1595 ( .A(n1338), .B(n749), .Z(n747) );
  IV U1596 ( .A(n745), .Z(n749) );
  XNOR U1597 ( .A(n1339), .B(n1340), .Z(n745) );
  NAND U1598 ( .A(n1341), .B(n1342), .Z(n1340) );
  XOR U1599 ( .A(n1339), .B(n1343), .Z(n1341) );
  NOR U1600 ( .A(n1344), .B(n1345), .Z(n1338) );
  XNOR U1601 ( .A(n778), .B(n758), .Z(n1346) );
  XNOR U1602 ( .A(n1347), .B(n1348), .Z(n758) );
  NANDN U1603 ( .A(n1349), .B(n1350), .Z(n1348) );
  XOR U1604 ( .A(n1347), .B(n1351), .Z(n1350) );
  XNOR U1605 ( .A(n1352), .B(n1353), .Z(n766) );
  NANDN U1606 ( .A(n1354), .B(n1355), .Z(n1353) );
  NANDN U1607 ( .A(n1356), .B(n1352), .Z(n1355) );
  XNOR U1608 ( .A(n1357), .B(n763), .Z(n765) );
  XNOR U1609 ( .A(n1358), .B(n1359), .Z(n763) );
  NAND U1610 ( .A(n1360), .B(n1361), .Z(n1359) );
  XNOR U1611 ( .A(n1358), .B(n1362), .Z(n1360) );
  NOR U1612 ( .A(n1363), .B(n1364), .Z(n1357) );
  XOR U1613 ( .A(n772), .B(n775), .Z(n1365) );
  XNOR U1614 ( .A(n1366), .B(n1367), .Z(n775) );
  NANDN U1615 ( .A(n1368), .B(n1369), .Z(n1367) );
  XNOR U1616 ( .A(n1366), .B(n1370), .Z(n1369) );
  XNOR U1617 ( .A(n1371), .B(n1372), .Z(n772) );
  NANDN U1618 ( .A(n1373), .B(n1374), .Z(n1372) );
  NANDN U1619 ( .A(n1371), .B(n1375), .Z(n1374) );
  XOR U1620 ( .A(n1376), .B(n773), .Z(n771) );
  IV U1621 ( .A(n769), .Z(n773) );
  XNOR U1622 ( .A(n1377), .B(n1378), .Z(n769) );
  NAND U1623 ( .A(n1379), .B(n1380), .Z(n1378) );
  XOR U1624 ( .A(n1377), .B(n1381), .Z(n1379) );
  NOR U1625 ( .A(n1382), .B(n1383), .Z(n1376) );
  XOR U1626 ( .A(n1384), .B(n1385), .Z(n780) );
  NANDN U1627 ( .A(n29), .B(n1386), .Z(n1385) );
  XNOR U1628 ( .A(n1384), .B(n30), .Z(n1386) );
  XOR U1629 ( .A(n791), .B(n792), .Z(n800) );
  XOR U1630 ( .A(n786), .B(n784), .Z(n792) );
  AND U1631 ( .A(n1387), .B(n782), .Z(n784) );
  OR U1632 ( .A(n1388), .B(n1389), .Z(n782) );
  OR U1633 ( .A(n1390), .B(n1391), .Z(n1387) );
  NOR U1634 ( .A(n1392), .B(n1393), .Z(n786) );
  XOR U1635 ( .A(n793), .B(n1394), .Z(n791) );
  XOR U1636 ( .A(n794), .B(n788), .Z(n1394) );
  NOR U1637 ( .A(n1395), .B(n1396), .Z(n788) );
  OR U1638 ( .A(n1397), .B(n1398), .Z(n794) );
  AND U1639 ( .A(n1399), .B(n1400), .Z(n793) );
  OR U1640 ( .A(n1401), .B(n1402), .Z(n1400) );
  OR U1641 ( .A(n1403), .B(n1404), .Z(n1399) );
  XNOR U1642 ( .A(n810), .B(n1405), .Z(n798) );
  XNOR U1643 ( .A(n796), .B(n811), .Z(n1405) );
  XOR U1644 ( .A(n805), .B(n803), .Z(n811) );
  NOR U1645 ( .A(n1407), .B(n1408), .Z(n801) );
  OR U1646 ( .A(n1409), .B(n1410), .Z(n1406) );
  OR U1647 ( .A(n1411), .B(n1412), .Z(n805) );
  OR U1648 ( .A(n1413), .B(n1414), .Z(n796) );
  XOR U1649 ( .A(n812), .B(n1415), .Z(n810) );
  XOR U1650 ( .A(n813), .B(n807), .Z(n1415) );
  NOR U1651 ( .A(n1416), .B(n1417), .Z(n807) );
  OR U1652 ( .A(n1418), .B(n1419), .Z(n813) );
  AND U1653 ( .A(n1420), .B(n1421), .Z(n812) );
  OR U1654 ( .A(n1422), .B(n1423), .Z(n1421) );
  OR U1655 ( .A(n1424), .B(n1425), .Z(n1420) );
  XOR U1656 ( .A(n815), .B(n838), .Z(n1426) );
  XNOR U1657 ( .A(n829), .B(n830), .Z(n838) );
  XOR U1658 ( .A(n824), .B(n822), .Z(n830) );
  AND U1659 ( .A(n1427), .B(n820), .Z(n822) );
  OR U1660 ( .A(n1428), .B(n1429), .Z(n820) );
  OR U1661 ( .A(n1430), .B(n1431), .Z(n1427) );
  NOR U1662 ( .A(n1432), .B(n1433), .Z(n824) );
  XOR U1663 ( .A(n831), .B(n1434), .Z(n829) );
  XOR U1664 ( .A(n832), .B(n826), .Z(n1434) );
  NOR U1665 ( .A(n1435), .B(n1436), .Z(n826) );
  OR U1666 ( .A(n1437), .B(n1438), .Z(n832) );
  AND U1667 ( .A(n1439), .B(n1440), .Z(n831) );
  OR U1668 ( .A(n1441), .B(n1442), .Z(n1440) );
  OR U1669 ( .A(n1443), .B(n1444), .Z(n1439) );
  OR U1670 ( .A(n1445), .B(n1446), .Z(n815) );
  XNOR U1671 ( .A(n848), .B(n1447), .Z(n836) );
  XNOR U1672 ( .A(n834), .B(n849), .Z(n1447) );
  XOR U1673 ( .A(n843), .B(n841), .Z(n849) );
  NOR U1674 ( .A(n1449), .B(n1450), .Z(n839) );
  OR U1675 ( .A(n1451), .B(n1452), .Z(n1448) );
  OR U1676 ( .A(n1453), .B(n1454), .Z(n843) );
  OR U1677 ( .A(n1455), .B(n1456), .Z(n834) );
  XOR U1678 ( .A(n850), .B(n1457), .Z(n848) );
  XOR U1679 ( .A(n851), .B(n845), .Z(n1457) );
  NOR U1680 ( .A(n1458), .B(n1459), .Z(n845) );
  OR U1681 ( .A(n1460), .B(n1461), .Z(n851) );
  AND U1682 ( .A(n1462), .B(n1463), .Z(n850) );
  OR U1683 ( .A(n1464), .B(n1465), .Z(n1463) );
  OR U1684 ( .A(n1466), .B(n1467), .Z(n1462) );
  XNOR U1685 ( .A(n853), .B(n895), .Z(n1468) );
  XOR U1686 ( .A(n867), .B(n868), .Z(n876) );
  XOR U1687 ( .A(n862), .B(n860), .Z(n868) );
  AND U1688 ( .A(n1469), .B(n858), .Z(n860) );
  OR U1689 ( .A(n1470), .B(n1471), .Z(n858) );
  OR U1690 ( .A(n1472), .B(n1473), .Z(n1469) );
  NOR U1691 ( .A(n1474), .B(n1475), .Z(n862) );
  XOR U1692 ( .A(n869), .B(n1476), .Z(n867) );
  XOR U1693 ( .A(n870), .B(n864), .Z(n1476) );
  NOR U1694 ( .A(n1477), .B(n1478), .Z(n864) );
  OR U1695 ( .A(n1479), .B(n1480), .Z(n870) );
  AND U1696 ( .A(n1481), .B(n1482), .Z(n869) );
  OR U1697 ( .A(n1483), .B(n1484), .Z(n1482) );
  OR U1698 ( .A(n1485), .B(n1486), .Z(n1481) );
  XNOR U1699 ( .A(n886), .B(n1487), .Z(n874) );
  XNOR U1700 ( .A(n872), .B(n887), .Z(n1487) );
  XOR U1701 ( .A(n881), .B(n879), .Z(n887) );
  NOR U1702 ( .A(n1489), .B(n1490), .Z(n877) );
  OR U1703 ( .A(n1491), .B(n1492), .Z(n1488) );
  OR U1704 ( .A(n1493), .B(n1494), .Z(n881) );
  OR U1705 ( .A(n1495), .B(n1496), .Z(n872) );
  XOR U1706 ( .A(n888), .B(n1497), .Z(n886) );
  XOR U1707 ( .A(n889), .B(n883), .Z(n1497) );
  NOR U1708 ( .A(n1498), .B(n1499), .Z(n883) );
  OR U1709 ( .A(n1500), .B(n1501), .Z(n889) );
  AND U1710 ( .A(n1502), .B(n1503), .Z(n888) );
  OR U1711 ( .A(n1504), .B(n1505), .Z(n1503) );
  OR U1712 ( .A(n1506), .B(n1507), .Z(n1502) );
  OR U1713 ( .A(n1508), .B(n1509), .Z(n853) );
  XOR U1714 ( .A(n891), .B(n914), .Z(n1510) );
  XNOR U1715 ( .A(n905), .B(n906), .Z(n914) );
  XOR U1716 ( .A(n900), .B(n898), .Z(n906) );
  AND U1717 ( .A(n1511), .B(n896), .Z(n898) );
  OR U1718 ( .A(n1512), .B(n1513), .Z(n896) );
  OR U1719 ( .A(n1514), .B(n1515), .Z(n1511) );
  NOR U1720 ( .A(n1516), .B(n1517), .Z(n900) );
  XOR U1721 ( .A(n907), .B(n1518), .Z(n905) );
  XOR U1722 ( .A(n908), .B(n902), .Z(n1518) );
  NOR U1723 ( .A(n1519), .B(n1520), .Z(n902) );
  OR U1724 ( .A(n1521), .B(n1522), .Z(n908) );
  AND U1725 ( .A(n1523), .B(n1524), .Z(n907) );
  OR U1726 ( .A(n1525), .B(n1526), .Z(n1524) );
  OR U1727 ( .A(n1527), .B(n1528), .Z(n1523) );
  OR U1728 ( .A(n1529), .B(n1530), .Z(n891) );
  XNOR U1729 ( .A(n924), .B(n1531), .Z(n912) );
  XNOR U1730 ( .A(n910), .B(n925), .Z(n1531) );
  XOR U1731 ( .A(n919), .B(n917), .Z(n925) );
  NOR U1732 ( .A(n1533), .B(n1534), .Z(n915) );
  OR U1733 ( .A(n1535), .B(n1536), .Z(n1532) );
  OR U1734 ( .A(n1537), .B(n1538), .Z(n919) );
  OR U1735 ( .A(n1539), .B(n1540), .Z(n910) );
  XOR U1736 ( .A(n926), .B(n1541), .Z(n924) );
  XOR U1737 ( .A(n927), .B(n921), .Z(n1541) );
  NOR U1738 ( .A(n1542), .B(n1543), .Z(n921) );
  OR U1739 ( .A(n1544), .B(n1545), .Z(n927) );
  AND U1740 ( .A(n1546), .B(n1547), .Z(n926) );
  OR U1741 ( .A(n1548), .B(n1549), .Z(n1547) );
  OR U1742 ( .A(n1550), .B(n1551), .Z(n1546) );
  XNOR U1743 ( .A(n929), .B(n1009), .Z(n1552) );
  XOR U1744 ( .A(n943), .B(n944), .Z(n952) );
  XOR U1745 ( .A(n938), .B(n936), .Z(n944) );
  AND U1746 ( .A(n1553), .B(n934), .Z(n936) );
  OR U1747 ( .A(n1554), .B(n1555), .Z(n934) );
  OR U1748 ( .A(n1556), .B(n1557), .Z(n1553) );
  NOR U1749 ( .A(n1558), .B(n1559), .Z(n938) );
  XOR U1750 ( .A(n945), .B(n1560), .Z(n943) );
  XOR U1751 ( .A(n946), .B(n940), .Z(n1560) );
  NOR U1752 ( .A(n1561), .B(n1562), .Z(n940) );
  OR U1753 ( .A(n1563), .B(n1564), .Z(n946) );
  AND U1754 ( .A(n1565), .B(n1566), .Z(n945) );
  OR U1755 ( .A(n1567), .B(n1568), .Z(n1566) );
  OR U1756 ( .A(n1569), .B(n1570), .Z(n1565) );
  XNOR U1757 ( .A(n962), .B(n1571), .Z(n950) );
  XNOR U1758 ( .A(n948), .B(n963), .Z(n1571) );
  XOR U1759 ( .A(n957), .B(n955), .Z(n963) );
  NOR U1760 ( .A(n1573), .B(n1574), .Z(n953) );
  OR U1761 ( .A(n1575), .B(n1576), .Z(n1572) );
  OR U1762 ( .A(n1577), .B(n1578), .Z(n957) );
  OR U1763 ( .A(n1579), .B(n1580), .Z(n948) );
  XOR U1764 ( .A(n964), .B(n1581), .Z(n962) );
  XOR U1765 ( .A(n965), .B(n959), .Z(n1581) );
  NOR U1766 ( .A(n1582), .B(n1583), .Z(n959) );
  OR U1767 ( .A(n1584), .B(n1585), .Z(n965) );
  AND U1768 ( .A(n1586), .B(n1587), .Z(n964) );
  OR U1769 ( .A(n1588), .B(n1589), .Z(n1587) );
  OR U1770 ( .A(n1590), .B(n1591), .Z(n1586) );
  XOR U1771 ( .A(n967), .B(n990), .Z(n1592) );
  XNOR U1772 ( .A(n981), .B(n982), .Z(n990) );
  XOR U1773 ( .A(n976), .B(n974), .Z(n982) );
  AND U1774 ( .A(n1593), .B(n972), .Z(n974) );
  OR U1775 ( .A(n1594), .B(n1595), .Z(n972) );
  OR U1776 ( .A(n1596), .B(n1597), .Z(n1593) );
  NOR U1777 ( .A(n1598), .B(n1599), .Z(n976) );
  XOR U1778 ( .A(n983), .B(n1600), .Z(n981) );
  XOR U1779 ( .A(n984), .B(n978), .Z(n1600) );
  NOR U1780 ( .A(n1601), .B(n1602), .Z(n978) );
  OR U1781 ( .A(n1603), .B(n1604), .Z(n984) );
  AND U1782 ( .A(n1605), .B(n1606), .Z(n983) );
  OR U1783 ( .A(n1607), .B(n1608), .Z(n1606) );
  OR U1784 ( .A(n1609), .B(n1610), .Z(n1605) );
  OR U1785 ( .A(n1611), .B(n1612), .Z(n967) );
  XNOR U1786 ( .A(n1000), .B(n1613), .Z(n988) );
  XNOR U1787 ( .A(n986), .B(n1001), .Z(n1613) );
  XOR U1788 ( .A(n995), .B(n993), .Z(n1001) );
  NOR U1789 ( .A(n1615), .B(n1616), .Z(n991) );
  OR U1790 ( .A(n1617), .B(n1618), .Z(n1614) );
  OR U1791 ( .A(n1619), .B(n1620), .Z(n995) );
  OR U1792 ( .A(n1621), .B(n1622), .Z(n986) );
  XOR U1793 ( .A(n1002), .B(n1623), .Z(n1000) );
  XOR U1794 ( .A(n1003), .B(n997), .Z(n1623) );
  NOR U1795 ( .A(n1624), .B(n1625), .Z(n997) );
  OR U1796 ( .A(n1626), .B(n1627), .Z(n1003) );
  AND U1797 ( .A(n1628), .B(n1629), .Z(n1002) );
  OR U1798 ( .A(n1630), .B(n1631), .Z(n1629) );
  OR U1799 ( .A(n1632), .B(n1633), .Z(n1628) );
  OR U1800 ( .A(n1634), .B(n1635), .Z(n929) );
  XNOR U1801 ( .A(n1005), .B(n1047), .Z(n1636) );
  XOR U1802 ( .A(n1019), .B(n1020), .Z(n1028) );
  XOR U1803 ( .A(n1014), .B(n1012), .Z(n1020) );
  AND U1804 ( .A(n1637), .B(n1010), .Z(n1012) );
  OR U1805 ( .A(n1638), .B(n1639), .Z(n1010) );
  OR U1806 ( .A(n1640), .B(n1641), .Z(n1637) );
  NOR U1807 ( .A(n1642), .B(n1643), .Z(n1014) );
  XOR U1808 ( .A(n1021), .B(n1644), .Z(n1019) );
  XOR U1809 ( .A(n1022), .B(n1016), .Z(n1644) );
  NOR U1810 ( .A(n1645), .B(n1646), .Z(n1016) );
  OR U1811 ( .A(n1647), .B(n1648), .Z(n1022) );
  AND U1812 ( .A(n1649), .B(n1650), .Z(n1021) );
  OR U1813 ( .A(n1651), .B(n1652), .Z(n1650) );
  OR U1814 ( .A(n1653), .B(n1654), .Z(n1649) );
  XNOR U1815 ( .A(n1038), .B(n1655), .Z(n1026) );
  XNOR U1816 ( .A(n1024), .B(n1039), .Z(n1655) );
  XOR U1817 ( .A(n1033), .B(n1031), .Z(n1039) );
  NOR U1818 ( .A(n1657), .B(n1658), .Z(n1029) );
  OR U1819 ( .A(n1659), .B(n1660), .Z(n1656) );
  OR U1820 ( .A(n1661), .B(n1662), .Z(n1033) );
  OR U1821 ( .A(n1663), .B(n1664), .Z(n1024) );
  XOR U1822 ( .A(n1040), .B(n1665), .Z(n1038) );
  XOR U1823 ( .A(n1041), .B(n1035), .Z(n1665) );
  NOR U1824 ( .A(n1666), .B(n1667), .Z(n1035) );
  OR U1825 ( .A(n1668), .B(n1669), .Z(n1041) );
  AND U1826 ( .A(n1670), .B(n1671), .Z(n1040) );
  OR U1827 ( .A(n1672), .B(n1673), .Z(n1671) );
  OR U1828 ( .A(n1674), .B(n1675), .Z(n1670) );
  OR U1829 ( .A(n1676), .B(n1677), .Z(n1005) );
  XOR U1830 ( .A(n1043), .B(n1066), .Z(n1678) );
  XNOR U1831 ( .A(n1057), .B(n1058), .Z(n1066) );
  XOR U1832 ( .A(n1052), .B(n1050), .Z(n1058) );
  AND U1833 ( .A(n1679), .B(n1048), .Z(n1050) );
  OR U1834 ( .A(n1680), .B(n1681), .Z(n1048) );
  OR U1835 ( .A(n1682), .B(n1683), .Z(n1679) );
  NOR U1836 ( .A(n1684), .B(n1685), .Z(n1052) );
  XOR U1837 ( .A(n1059), .B(n1686), .Z(n1057) );
  XOR U1838 ( .A(n1060), .B(n1054), .Z(n1686) );
  NOR U1839 ( .A(n1687), .B(n1688), .Z(n1054) );
  OR U1840 ( .A(n1689), .B(n1690), .Z(n1060) );
  AND U1841 ( .A(n1691), .B(n1692), .Z(n1059) );
  OR U1842 ( .A(n1693), .B(n1694), .Z(n1692) );
  OR U1843 ( .A(n1695), .B(n1696), .Z(n1691) );
  OR U1844 ( .A(n1697), .B(n1698), .Z(n1043) );
  XNOR U1845 ( .A(n1076), .B(n1699), .Z(n1064) );
  XNOR U1846 ( .A(n1062), .B(n1077), .Z(n1699) );
  XOR U1847 ( .A(n1071), .B(n1069), .Z(n1077) );
  NOR U1848 ( .A(n1701), .B(n1702), .Z(n1067) );
  OR U1849 ( .A(n1703), .B(n1704), .Z(n1700) );
  OR U1850 ( .A(n1705), .B(n1706), .Z(n1071) );
  OR U1851 ( .A(n1707), .B(n1708), .Z(n1062) );
  XOR U1852 ( .A(n1078), .B(n1709), .Z(n1076) );
  XOR U1853 ( .A(n1079), .B(n1073), .Z(n1709) );
  NOR U1854 ( .A(n1710), .B(n1711), .Z(n1073) );
  OR U1855 ( .A(n1712), .B(n1713), .Z(n1079) );
  AND U1856 ( .A(n1714), .B(n1715), .Z(n1078) );
  OR U1857 ( .A(n1716), .B(n1717), .Z(n1715) );
  OR U1858 ( .A(n1718), .B(n1719), .Z(n1714) );
  XNOR U1859 ( .A(n1081), .B(n1237), .Z(n1720) );
  XOR U1860 ( .A(n1095), .B(n1096), .Z(n1104) );
  XOR U1861 ( .A(n1090), .B(n1088), .Z(n1096) );
  AND U1862 ( .A(n1721), .B(n1086), .Z(n1088) );
  OR U1863 ( .A(n1722), .B(n1723), .Z(n1086) );
  OR U1864 ( .A(n1724), .B(n1725), .Z(n1721) );
  NOR U1865 ( .A(n1726), .B(n1727), .Z(n1090) );
  XOR U1866 ( .A(n1097), .B(n1728), .Z(n1095) );
  XOR U1867 ( .A(n1098), .B(n1092), .Z(n1728) );
  NOR U1868 ( .A(n1729), .B(n1730), .Z(n1092) );
  OR U1869 ( .A(n1731), .B(n1732), .Z(n1098) );
  AND U1870 ( .A(n1733), .B(n1734), .Z(n1097) );
  OR U1871 ( .A(n1735), .B(n1736), .Z(n1734) );
  OR U1872 ( .A(n1737), .B(n1738), .Z(n1733) );
  XNOR U1873 ( .A(n1114), .B(n1739), .Z(n1102) );
  XNOR U1874 ( .A(n1100), .B(n1115), .Z(n1739) );
  XOR U1875 ( .A(n1109), .B(n1107), .Z(n1115) );
  NOR U1876 ( .A(n1741), .B(n1742), .Z(n1105) );
  OR U1877 ( .A(n1743), .B(n1744), .Z(n1740) );
  OR U1878 ( .A(n1745), .B(n1746), .Z(n1109) );
  OR U1879 ( .A(n1747), .B(n1748), .Z(n1100) );
  XOR U1880 ( .A(n1116), .B(n1749), .Z(n1114) );
  XOR U1881 ( .A(n1117), .B(n1111), .Z(n1749) );
  NOR U1882 ( .A(n1750), .B(n1751), .Z(n1111) );
  OR U1883 ( .A(n1752), .B(n1753), .Z(n1117) );
  AND U1884 ( .A(n1754), .B(n1755), .Z(n1116) );
  OR U1885 ( .A(n1756), .B(n1757), .Z(n1755) );
  OR U1886 ( .A(n1758), .B(n1759), .Z(n1754) );
  XOR U1887 ( .A(n1119), .B(n1142), .Z(n1760) );
  XNOR U1888 ( .A(n1133), .B(n1134), .Z(n1142) );
  XOR U1889 ( .A(n1128), .B(n1126), .Z(n1134) );
  AND U1890 ( .A(n1761), .B(n1124), .Z(n1126) );
  OR U1891 ( .A(n1762), .B(n1763), .Z(n1124) );
  OR U1892 ( .A(n1764), .B(n1765), .Z(n1761) );
  NOR U1893 ( .A(n1766), .B(n1767), .Z(n1128) );
  XOR U1894 ( .A(n1135), .B(n1768), .Z(n1133) );
  XOR U1895 ( .A(n1136), .B(n1130), .Z(n1768) );
  NOR U1896 ( .A(n1769), .B(n1770), .Z(n1130) );
  OR U1897 ( .A(n1771), .B(n1772), .Z(n1136) );
  AND U1898 ( .A(n1773), .B(n1774), .Z(n1135) );
  OR U1899 ( .A(n1775), .B(n1776), .Z(n1774) );
  OR U1900 ( .A(n1777), .B(n1778), .Z(n1773) );
  OR U1901 ( .A(n1779), .B(n1780), .Z(n1119) );
  XNOR U1902 ( .A(n1152), .B(n1781), .Z(n1140) );
  XNOR U1903 ( .A(n1138), .B(n1153), .Z(n1781) );
  XOR U1904 ( .A(n1147), .B(n1145), .Z(n1153) );
  NOR U1905 ( .A(n1783), .B(n1784), .Z(n1143) );
  OR U1906 ( .A(n1785), .B(n1786), .Z(n1782) );
  OR U1907 ( .A(n1787), .B(n1788), .Z(n1147) );
  OR U1908 ( .A(n1789), .B(n1790), .Z(n1138) );
  XOR U1909 ( .A(n1154), .B(n1791), .Z(n1152) );
  XOR U1910 ( .A(n1155), .B(n1149), .Z(n1791) );
  NOR U1911 ( .A(n1792), .B(n1793), .Z(n1149) );
  OR U1912 ( .A(n1794), .B(n1795), .Z(n1155) );
  AND U1913 ( .A(n1796), .B(n1797), .Z(n1154) );
  OR U1914 ( .A(n1798), .B(n1799), .Z(n1797) );
  OR U1915 ( .A(n1800), .B(n1801), .Z(n1796) );
  XNOR U1916 ( .A(n1157), .B(n1199), .Z(n1802) );
  XOR U1917 ( .A(n1171), .B(n1172), .Z(n1180) );
  XOR U1918 ( .A(n1166), .B(n1164), .Z(n1172) );
  AND U1919 ( .A(n1803), .B(n1162), .Z(n1164) );
  OR U1920 ( .A(n1804), .B(n1805), .Z(n1162) );
  OR U1921 ( .A(n1806), .B(n1807), .Z(n1803) );
  NOR U1922 ( .A(n1808), .B(n1809), .Z(n1166) );
  XOR U1923 ( .A(n1173), .B(n1810), .Z(n1171) );
  XOR U1924 ( .A(n1174), .B(n1168), .Z(n1810) );
  NOR U1925 ( .A(n1811), .B(n1812), .Z(n1168) );
  OR U1926 ( .A(n1813), .B(n1814), .Z(n1174) );
  AND U1927 ( .A(n1815), .B(n1816), .Z(n1173) );
  OR U1928 ( .A(n1817), .B(n1818), .Z(n1816) );
  OR U1929 ( .A(n1819), .B(n1820), .Z(n1815) );
  XNOR U1930 ( .A(n1190), .B(n1821), .Z(n1178) );
  XNOR U1931 ( .A(n1176), .B(n1191), .Z(n1821) );
  XOR U1932 ( .A(n1185), .B(n1183), .Z(n1191) );
  NOR U1933 ( .A(n1823), .B(n1824), .Z(n1181) );
  OR U1934 ( .A(n1825), .B(n1826), .Z(n1822) );
  OR U1935 ( .A(n1827), .B(n1828), .Z(n1185) );
  OR U1936 ( .A(n1829), .B(n1830), .Z(n1176) );
  XOR U1937 ( .A(n1192), .B(n1831), .Z(n1190) );
  XOR U1938 ( .A(n1193), .B(n1187), .Z(n1831) );
  NOR U1939 ( .A(n1832), .B(n1833), .Z(n1187) );
  OR U1940 ( .A(n1834), .B(n1835), .Z(n1193) );
  AND U1941 ( .A(n1836), .B(n1837), .Z(n1192) );
  OR U1942 ( .A(n1838), .B(n1839), .Z(n1837) );
  OR U1943 ( .A(n1840), .B(n1841), .Z(n1836) );
  OR U1944 ( .A(n1842), .B(n1843), .Z(n1157) );
  XOR U1945 ( .A(n1195), .B(n1218), .Z(n1844) );
  XNOR U1946 ( .A(n1209), .B(n1210), .Z(n1218) );
  XOR U1947 ( .A(n1204), .B(n1202), .Z(n1210) );
  AND U1948 ( .A(n1845), .B(n1200), .Z(n1202) );
  OR U1949 ( .A(n1846), .B(n1847), .Z(n1200) );
  OR U1950 ( .A(n1848), .B(n1849), .Z(n1845) );
  NOR U1951 ( .A(n1850), .B(n1851), .Z(n1204) );
  XOR U1952 ( .A(n1211), .B(n1852), .Z(n1209) );
  XOR U1953 ( .A(n1212), .B(n1206), .Z(n1852) );
  NOR U1954 ( .A(n1853), .B(n1854), .Z(n1206) );
  OR U1955 ( .A(n1855), .B(n1856), .Z(n1212) );
  AND U1956 ( .A(n1857), .B(n1858), .Z(n1211) );
  OR U1957 ( .A(n1859), .B(n1860), .Z(n1858) );
  OR U1958 ( .A(n1861), .B(n1862), .Z(n1857) );
  OR U1959 ( .A(n1863), .B(n1864), .Z(n1195) );
  XNOR U1960 ( .A(n1228), .B(n1865), .Z(n1216) );
  XNOR U1961 ( .A(n1214), .B(n1229), .Z(n1865) );
  XOR U1962 ( .A(n1223), .B(n1221), .Z(n1229) );
  NOR U1963 ( .A(n1867), .B(n1868), .Z(n1219) );
  OR U1964 ( .A(n1869), .B(n1870), .Z(n1866) );
  OR U1965 ( .A(n1871), .B(n1872), .Z(n1223) );
  OR U1966 ( .A(n1873), .B(n1874), .Z(n1214) );
  XOR U1967 ( .A(n1230), .B(n1875), .Z(n1228) );
  XOR U1968 ( .A(n1231), .B(n1225), .Z(n1875) );
  NOR U1969 ( .A(n1876), .B(n1877), .Z(n1225) );
  OR U1970 ( .A(n1878), .B(n1879), .Z(n1231) );
  AND U1971 ( .A(n1880), .B(n1881), .Z(n1230) );
  OR U1972 ( .A(n1882), .B(n1883), .Z(n1881) );
  OR U1973 ( .A(n1884), .B(n1885), .Z(n1880) );
  OR U1974 ( .A(n1886), .B(n1887), .Z(n1081) );
  XNOR U1975 ( .A(n1233), .B(n1313), .Z(n1888) );
  XOR U1976 ( .A(n1247), .B(n1248), .Z(n1256) );
  XOR U1977 ( .A(n1242), .B(n1240), .Z(n1248) );
  AND U1978 ( .A(n1889), .B(n1238), .Z(n1240) );
  OR U1979 ( .A(n1890), .B(n1891), .Z(n1238) );
  OR U1980 ( .A(n1892), .B(n1893), .Z(n1889) );
  NOR U1981 ( .A(n1894), .B(n1895), .Z(n1242) );
  XOR U1982 ( .A(n1249), .B(n1896), .Z(n1247) );
  XOR U1983 ( .A(n1250), .B(n1244), .Z(n1896) );
  NOR U1984 ( .A(n1897), .B(n1898), .Z(n1244) );
  OR U1985 ( .A(n1899), .B(n1900), .Z(n1250) );
  AND U1986 ( .A(n1901), .B(n1902), .Z(n1249) );
  OR U1987 ( .A(n1903), .B(n1904), .Z(n1902) );
  OR U1988 ( .A(n1905), .B(n1906), .Z(n1901) );
  XNOR U1989 ( .A(n1266), .B(n1907), .Z(n1254) );
  XNOR U1990 ( .A(n1252), .B(n1267), .Z(n1907) );
  XOR U1991 ( .A(n1261), .B(n1259), .Z(n1267) );
  NOR U1992 ( .A(n1909), .B(n1910), .Z(n1257) );
  OR U1993 ( .A(n1911), .B(n1912), .Z(n1908) );
  OR U1994 ( .A(n1913), .B(n1914), .Z(n1261) );
  OR U1995 ( .A(n1915), .B(n1916), .Z(n1252) );
  XOR U1996 ( .A(n1268), .B(n1917), .Z(n1266) );
  XOR U1997 ( .A(n1269), .B(n1263), .Z(n1917) );
  NOR U1998 ( .A(n1918), .B(n1919), .Z(n1263) );
  OR U1999 ( .A(n1920), .B(n1921), .Z(n1269) );
  AND U2000 ( .A(n1922), .B(n1923), .Z(n1268) );
  OR U2001 ( .A(n1924), .B(n1925), .Z(n1923) );
  OR U2002 ( .A(n1926), .B(n1927), .Z(n1922) );
  XOR U2003 ( .A(n1271), .B(n1294), .Z(n1928) );
  XNOR U2004 ( .A(n1285), .B(n1286), .Z(n1294) );
  XOR U2005 ( .A(n1280), .B(n1278), .Z(n1286) );
  AND U2006 ( .A(n1929), .B(n1276), .Z(n1278) );
  OR U2007 ( .A(n1930), .B(n1931), .Z(n1276) );
  OR U2008 ( .A(n1932), .B(n1933), .Z(n1929) );
  NOR U2009 ( .A(n1934), .B(n1935), .Z(n1280) );
  XOR U2010 ( .A(n1287), .B(n1936), .Z(n1285) );
  XOR U2011 ( .A(n1288), .B(n1282), .Z(n1936) );
  NOR U2012 ( .A(n1937), .B(n1938), .Z(n1282) );
  OR U2013 ( .A(n1939), .B(n1940), .Z(n1288) );
  AND U2014 ( .A(n1941), .B(n1942), .Z(n1287) );
  OR U2015 ( .A(n1943), .B(n1944), .Z(n1942) );
  OR U2016 ( .A(n1945), .B(n1946), .Z(n1941) );
  OR U2017 ( .A(n1947), .B(n1948), .Z(n1271) );
  XNOR U2018 ( .A(n1304), .B(n1949), .Z(n1292) );
  XNOR U2019 ( .A(n1290), .B(n1305), .Z(n1949) );
  XOR U2020 ( .A(n1299), .B(n1297), .Z(n1305) );
  NOR U2021 ( .A(n1951), .B(n1952), .Z(n1295) );
  OR U2022 ( .A(n1953), .B(n1954), .Z(n1950) );
  OR U2023 ( .A(n1955), .B(n1956), .Z(n1299) );
  OR U2024 ( .A(n1957), .B(n1958), .Z(n1290) );
  XOR U2025 ( .A(n1306), .B(n1959), .Z(n1304) );
  XOR U2026 ( .A(n1307), .B(n1301), .Z(n1959) );
  NOR U2027 ( .A(n1960), .B(n1961), .Z(n1301) );
  OR U2028 ( .A(n1962), .B(n1963), .Z(n1307) );
  AND U2029 ( .A(n1964), .B(n1965), .Z(n1306) );
  OR U2030 ( .A(n1966), .B(n1967), .Z(n1965) );
  OR U2031 ( .A(n1968), .B(n1969), .Z(n1964) );
  OR U2032 ( .A(n1970), .B(n1971), .Z(n1233) );
  XNOR U2033 ( .A(n1309), .B(n1351), .Z(n1972) );
  XOR U2034 ( .A(n1323), .B(n1324), .Z(n1332) );
  XOR U2035 ( .A(n1318), .B(n1316), .Z(n1324) );
  AND U2036 ( .A(n1973), .B(n1314), .Z(n1316) );
  OR U2037 ( .A(n1974), .B(n1975), .Z(n1314) );
  OR U2038 ( .A(n1976), .B(n1977), .Z(n1973) );
  NOR U2039 ( .A(n1978), .B(n1979), .Z(n1318) );
  XOR U2040 ( .A(n1325), .B(n1980), .Z(n1323) );
  XOR U2041 ( .A(n1326), .B(n1320), .Z(n1980) );
  NOR U2042 ( .A(n1981), .B(n1982), .Z(n1320) );
  OR U2043 ( .A(n1983), .B(n1984), .Z(n1326) );
  AND U2044 ( .A(n1985), .B(n1986), .Z(n1325) );
  OR U2045 ( .A(n1987), .B(n1988), .Z(n1986) );
  OR U2046 ( .A(n1989), .B(n1990), .Z(n1985) );
  XNOR U2047 ( .A(n1342), .B(n1991), .Z(n1330) );
  XNOR U2048 ( .A(n1328), .B(n1343), .Z(n1991) );
  XOR U2049 ( .A(n1337), .B(n1335), .Z(n1343) );
  NOR U2050 ( .A(n1993), .B(n1994), .Z(n1333) );
  OR U2051 ( .A(n1995), .B(n1996), .Z(n1992) );
  OR U2052 ( .A(n1997), .B(n1998), .Z(n1337) );
  OR U2053 ( .A(n1999), .B(n2000), .Z(n1328) );
  XOR U2054 ( .A(n1344), .B(n2001), .Z(n1342) );
  XOR U2055 ( .A(n1345), .B(n1339), .Z(n2001) );
  NOR U2056 ( .A(n2002), .B(n2003), .Z(n1339) );
  OR U2057 ( .A(n2004), .B(n2005), .Z(n1345) );
  AND U2058 ( .A(n2006), .B(n2007), .Z(n1344) );
  OR U2059 ( .A(n2008), .B(n2009), .Z(n2007) );
  OR U2060 ( .A(n2010), .B(n2011), .Z(n2006) );
  OR U2061 ( .A(n2012), .B(n2013), .Z(n1309) );
  XOR U2062 ( .A(n1347), .B(n1370), .Z(n2014) );
  XNOR U2063 ( .A(n1361), .B(n1362), .Z(n1370) );
  XOR U2064 ( .A(n1356), .B(n1354), .Z(n1362) );
  AND U2065 ( .A(n2015), .B(n1352), .Z(n1354) );
  OR U2066 ( .A(n2016), .B(n2017), .Z(n1352) );
  OR U2067 ( .A(n2018), .B(n2019), .Z(n2015) );
  NOR U2068 ( .A(n2020), .B(n2021), .Z(n1356) );
  XOR U2069 ( .A(n1363), .B(n2022), .Z(n1361) );
  XOR U2070 ( .A(n1364), .B(n1358), .Z(n2022) );
  NOR U2071 ( .A(n2023), .B(n2024), .Z(n1358) );
  OR U2072 ( .A(n2025), .B(n2026), .Z(n1364) );
  AND U2073 ( .A(n2027), .B(n2028), .Z(n1363) );
  OR U2074 ( .A(n2029), .B(n2030), .Z(n2028) );
  OR U2075 ( .A(n2031), .B(n2032), .Z(n2027) );
  OR U2076 ( .A(n2033), .B(n2034), .Z(n1347) );
  XNOR U2077 ( .A(n1380), .B(n2035), .Z(n1368) );
  XNOR U2078 ( .A(n1366), .B(n1381), .Z(n2035) );
  XOR U2079 ( .A(n1375), .B(n1373), .Z(n1381) );
  NOR U2080 ( .A(n2037), .B(n2038), .Z(n1371) );
  OR U2081 ( .A(n2039), .B(n2040), .Z(n2036) );
  OR U2082 ( .A(n2041), .B(n2042), .Z(n1375) );
  OR U2083 ( .A(n2043), .B(n2044), .Z(n1366) );
  XOR U2084 ( .A(n1382), .B(n2045), .Z(n1380) );
  XOR U2085 ( .A(n1383), .B(n1377), .Z(n2045) );
  NOR U2086 ( .A(n2046), .B(n2047), .Z(n1377) );
  OR U2087 ( .A(n2048), .B(n2049), .Z(n1383) );
  AND U2088 ( .A(n2050), .B(n2051), .Z(n1382) );
  OR U2089 ( .A(n2052), .B(n2053), .Z(n2051) );
  OR U2090 ( .A(n2054), .B(n2055), .Z(n2050) );
  XNOR U2091 ( .A(oglobal[1]), .B(n1384), .Z(n29) );
  ANDN U2092 ( .B(oglobal[0]), .A(n2056), .Z(n1384) );
  XNOR U2093 ( .A(oglobal[0]), .B(n2056), .Z(o[0]) );
  XNOR U2094 ( .A(n1887), .B(n1886), .Z(n2056) );
  XNOR U2095 ( .A(n1635), .B(n1634), .Z(n1886) );
  XNOR U2096 ( .A(n1509), .B(n1508), .Z(n1634) );
  XNOR U2097 ( .A(n1446), .B(n1445), .Z(n1508) );
  XNOR U2098 ( .A(n1414), .B(n1413), .Z(n1445) );
  XNOR U2099 ( .A(n1388), .B(n1389), .Z(n1395) );
  XNOR U2100 ( .A(n1392), .B(n1393), .Z(n1389) );
  XNOR U2101 ( .A(y[255]), .B(x[255]), .Z(n1393) );
  XNOR U2102 ( .A(y[254]), .B(x[254]), .Z(n1392) );
  XNOR U2103 ( .A(n1390), .B(n1391), .Z(n1388) );
  XNOR U2104 ( .A(y[253]), .B(x[253]), .Z(n1391) );
  XNOR U2105 ( .A(y[252]), .B(x[252]), .Z(n1390) );
  XNOR U2106 ( .A(n1403), .B(n1404), .Z(n1396) );
  XNOR U2107 ( .A(n1398), .B(n1397), .Z(n1404) );
  XNOR U2108 ( .A(y[251]), .B(x[251]), .Z(n1397) );
  XNOR U2109 ( .A(y[250]), .B(x[250]), .Z(n1398) );
  XNOR U2110 ( .A(n1401), .B(n1402), .Z(n1403) );
  XNOR U2111 ( .A(y[249]), .B(x[249]), .Z(n1402) );
  XNOR U2112 ( .A(y[248]), .B(x[248]), .Z(n1401) );
  XNOR U2113 ( .A(n1407), .B(n1408), .Z(n1416) );
  XNOR U2114 ( .A(n1411), .B(n1412), .Z(n1408) );
  XNOR U2115 ( .A(y[247]), .B(x[247]), .Z(n1412) );
  XNOR U2116 ( .A(y[246]), .B(x[246]), .Z(n1411) );
  XNOR U2117 ( .A(n1409), .B(n1410), .Z(n1407) );
  XNOR U2118 ( .A(y[245]), .B(x[245]), .Z(n1410) );
  XNOR U2119 ( .A(y[244]), .B(x[244]), .Z(n1409) );
  XNOR U2120 ( .A(n1424), .B(n1425), .Z(n1417) );
  XNOR U2121 ( .A(n1419), .B(n1418), .Z(n1425) );
  XNOR U2122 ( .A(y[243]), .B(x[243]), .Z(n1418) );
  XNOR U2123 ( .A(y[242]), .B(x[242]), .Z(n1419) );
  XNOR U2124 ( .A(n1422), .B(n1423), .Z(n1424) );
  XNOR U2125 ( .A(y[241]), .B(x[241]), .Z(n1423) );
  XNOR U2126 ( .A(y[240]), .B(x[240]), .Z(n1422) );
  XNOR U2127 ( .A(n1456), .B(n1455), .Z(n1446) );
  XNOR U2128 ( .A(n1428), .B(n1429), .Z(n1435) );
  XNOR U2129 ( .A(n1432), .B(n1433), .Z(n1429) );
  XNOR U2130 ( .A(y[239]), .B(x[239]), .Z(n1433) );
  XNOR U2131 ( .A(y[238]), .B(x[238]), .Z(n1432) );
  XNOR U2132 ( .A(n1430), .B(n1431), .Z(n1428) );
  XNOR U2133 ( .A(y[237]), .B(x[237]), .Z(n1431) );
  XNOR U2134 ( .A(y[236]), .B(x[236]), .Z(n1430) );
  XNOR U2135 ( .A(n1443), .B(n1444), .Z(n1436) );
  XNOR U2136 ( .A(n1438), .B(n1437), .Z(n1444) );
  XNOR U2137 ( .A(y[235]), .B(x[235]), .Z(n1437) );
  XNOR U2138 ( .A(y[234]), .B(x[234]), .Z(n1438) );
  XNOR U2139 ( .A(n1441), .B(n1442), .Z(n1443) );
  XNOR U2140 ( .A(y[233]), .B(x[233]), .Z(n1442) );
  XNOR U2141 ( .A(y[232]), .B(x[232]), .Z(n1441) );
  XNOR U2142 ( .A(n1449), .B(n1450), .Z(n1458) );
  XNOR U2143 ( .A(n1453), .B(n1454), .Z(n1450) );
  XNOR U2144 ( .A(y[231]), .B(x[231]), .Z(n1454) );
  XNOR U2145 ( .A(y[230]), .B(x[230]), .Z(n1453) );
  XNOR U2146 ( .A(n1451), .B(n1452), .Z(n1449) );
  XNOR U2147 ( .A(y[229]), .B(x[229]), .Z(n1452) );
  XNOR U2148 ( .A(y[228]), .B(x[228]), .Z(n1451) );
  XNOR U2149 ( .A(n1466), .B(n1467), .Z(n1459) );
  XNOR U2150 ( .A(n1461), .B(n1460), .Z(n1467) );
  XNOR U2151 ( .A(y[227]), .B(x[227]), .Z(n1460) );
  XNOR U2152 ( .A(y[226]), .B(x[226]), .Z(n1461) );
  XNOR U2153 ( .A(n1464), .B(n1465), .Z(n1466) );
  XNOR U2154 ( .A(y[225]), .B(x[225]), .Z(n1465) );
  XNOR U2155 ( .A(y[224]), .B(x[224]), .Z(n1464) );
  XNOR U2156 ( .A(n1530), .B(n1529), .Z(n1509) );
  XNOR U2157 ( .A(n1496), .B(n1495), .Z(n1529) );
  XNOR U2158 ( .A(n1470), .B(n1471), .Z(n1477) );
  XNOR U2159 ( .A(n1474), .B(n1475), .Z(n1471) );
  XNOR U2160 ( .A(y[223]), .B(x[223]), .Z(n1475) );
  XNOR U2161 ( .A(y[222]), .B(x[222]), .Z(n1474) );
  XNOR U2162 ( .A(n1472), .B(n1473), .Z(n1470) );
  XNOR U2163 ( .A(y[221]), .B(x[221]), .Z(n1473) );
  XNOR U2164 ( .A(y[220]), .B(x[220]), .Z(n1472) );
  XNOR U2165 ( .A(n1485), .B(n1486), .Z(n1478) );
  XNOR U2166 ( .A(n1480), .B(n1479), .Z(n1486) );
  XNOR U2167 ( .A(y[219]), .B(x[219]), .Z(n1479) );
  XNOR U2168 ( .A(y[218]), .B(x[218]), .Z(n1480) );
  XNOR U2169 ( .A(n1483), .B(n1484), .Z(n1485) );
  XNOR U2170 ( .A(y[217]), .B(x[217]), .Z(n1484) );
  XNOR U2171 ( .A(y[216]), .B(x[216]), .Z(n1483) );
  XNOR U2172 ( .A(n1489), .B(n1490), .Z(n1498) );
  XNOR U2173 ( .A(n1493), .B(n1494), .Z(n1490) );
  XNOR U2174 ( .A(y[215]), .B(x[215]), .Z(n1494) );
  XNOR U2175 ( .A(y[214]), .B(x[214]), .Z(n1493) );
  XNOR U2176 ( .A(n1491), .B(n1492), .Z(n1489) );
  XNOR U2177 ( .A(y[213]), .B(x[213]), .Z(n1492) );
  XNOR U2178 ( .A(y[212]), .B(x[212]), .Z(n1491) );
  XNOR U2179 ( .A(n1506), .B(n1507), .Z(n1499) );
  XNOR U2180 ( .A(n1501), .B(n1500), .Z(n1507) );
  XNOR U2181 ( .A(y[211]), .B(x[211]), .Z(n1500) );
  XNOR U2182 ( .A(y[210]), .B(x[210]), .Z(n1501) );
  XNOR U2183 ( .A(n1504), .B(n1505), .Z(n1506) );
  XNOR U2184 ( .A(y[209]), .B(x[209]), .Z(n1505) );
  XNOR U2185 ( .A(y[208]), .B(x[208]), .Z(n1504) );
  XNOR U2186 ( .A(n1540), .B(n1539), .Z(n1530) );
  XNOR U2187 ( .A(n1512), .B(n1513), .Z(n1519) );
  XNOR U2188 ( .A(n1516), .B(n1517), .Z(n1513) );
  XNOR U2189 ( .A(y[207]), .B(x[207]), .Z(n1517) );
  XNOR U2190 ( .A(y[206]), .B(x[206]), .Z(n1516) );
  XNOR U2191 ( .A(n1514), .B(n1515), .Z(n1512) );
  XNOR U2192 ( .A(y[205]), .B(x[205]), .Z(n1515) );
  XNOR U2193 ( .A(y[204]), .B(x[204]), .Z(n1514) );
  XNOR U2194 ( .A(n1527), .B(n1528), .Z(n1520) );
  XNOR U2195 ( .A(n1522), .B(n1521), .Z(n1528) );
  XNOR U2196 ( .A(y[203]), .B(x[203]), .Z(n1521) );
  XNOR U2197 ( .A(y[202]), .B(x[202]), .Z(n1522) );
  XNOR U2198 ( .A(n1525), .B(n1526), .Z(n1527) );
  XNOR U2199 ( .A(y[201]), .B(x[201]), .Z(n1526) );
  XNOR U2200 ( .A(y[200]), .B(x[200]), .Z(n1525) );
  XNOR U2201 ( .A(n1533), .B(n1534), .Z(n1542) );
  XNOR U2202 ( .A(n1537), .B(n1538), .Z(n1534) );
  XNOR U2203 ( .A(y[199]), .B(x[199]), .Z(n1538) );
  XNOR U2204 ( .A(y[198]), .B(x[198]), .Z(n1537) );
  XNOR U2205 ( .A(n1535), .B(n1536), .Z(n1533) );
  XNOR U2206 ( .A(y[197]), .B(x[197]), .Z(n1536) );
  XNOR U2207 ( .A(y[196]), .B(x[196]), .Z(n1535) );
  XNOR U2208 ( .A(n1550), .B(n1551), .Z(n1543) );
  XNOR U2209 ( .A(n1545), .B(n1544), .Z(n1551) );
  XNOR U2210 ( .A(y[195]), .B(x[195]), .Z(n1544) );
  XNOR U2211 ( .A(y[194]), .B(x[194]), .Z(n1545) );
  XNOR U2212 ( .A(n1548), .B(n1549), .Z(n1550) );
  XNOR U2213 ( .A(y[193]), .B(x[193]), .Z(n1549) );
  XNOR U2214 ( .A(y[192]), .B(x[192]), .Z(n1548) );
  XNOR U2215 ( .A(n1677), .B(n1676), .Z(n1635) );
  XNOR U2216 ( .A(n1612), .B(n1611), .Z(n1676) );
  XNOR U2217 ( .A(n1580), .B(n1579), .Z(n1611) );
  XNOR U2218 ( .A(n1554), .B(n1555), .Z(n1561) );
  XNOR U2219 ( .A(n1558), .B(n1559), .Z(n1555) );
  XNOR U2220 ( .A(y[191]), .B(x[191]), .Z(n1559) );
  XNOR U2221 ( .A(y[190]), .B(x[190]), .Z(n1558) );
  XNOR U2222 ( .A(n1556), .B(n1557), .Z(n1554) );
  XNOR U2223 ( .A(y[189]), .B(x[189]), .Z(n1557) );
  XNOR U2224 ( .A(y[188]), .B(x[188]), .Z(n1556) );
  XNOR U2225 ( .A(n1569), .B(n1570), .Z(n1562) );
  XNOR U2226 ( .A(n1564), .B(n1563), .Z(n1570) );
  XNOR U2227 ( .A(y[187]), .B(x[187]), .Z(n1563) );
  XNOR U2228 ( .A(y[186]), .B(x[186]), .Z(n1564) );
  XNOR U2229 ( .A(n1567), .B(n1568), .Z(n1569) );
  XNOR U2230 ( .A(y[185]), .B(x[185]), .Z(n1568) );
  XNOR U2231 ( .A(y[184]), .B(x[184]), .Z(n1567) );
  XNOR U2232 ( .A(n1573), .B(n1574), .Z(n1582) );
  XNOR U2233 ( .A(n1577), .B(n1578), .Z(n1574) );
  XNOR U2234 ( .A(y[183]), .B(x[183]), .Z(n1578) );
  XNOR U2235 ( .A(y[182]), .B(x[182]), .Z(n1577) );
  XNOR U2236 ( .A(n1575), .B(n1576), .Z(n1573) );
  XNOR U2237 ( .A(y[181]), .B(x[181]), .Z(n1576) );
  XNOR U2238 ( .A(y[180]), .B(x[180]), .Z(n1575) );
  XNOR U2239 ( .A(n1590), .B(n1591), .Z(n1583) );
  XNOR U2240 ( .A(n1585), .B(n1584), .Z(n1591) );
  XNOR U2241 ( .A(y[179]), .B(x[179]), .Z(n1584) );
  XNOR U2242 ( .A(y[178]), .B(x[178]), .Z(n1585) );
  XNOR U2243 ( .A(n1588), .B(n1589), .Z(n1590) );
  XNOR U2244 ( .A(y[177]), .B(x[177]), .Z(n1589) );
  XNOR U2245 ( .A(y[176]), .B(x[176]), .Z(n1588) );
  XNOR U2246 ( .A(n1622), .B(n1621), .Z(n1612) );
  XNOR U2247 ( .A(n1594), .B(n1595), .Z(n1601) );
  XNOR U2248 ( .A(n1598), .B(n1599), .Z(n1595) );
  XNOR U2249 ( .A(y[175]), .B(x[175]), .Z(n1599) );
  XNOR U2250 ( .A(y[174]), .B(x[174]), .Z(n1598) );
  XNOR U2251 ( .A(n1596), .B(n1597), .Z(n1594) );
  XNOR U2252 ( .A(y[173]), .B(x[173]), .Z(n1597) );
  XNOR U2253 ( .A(y[172]), .B(x[172]), .Z(n1596) );
  XNOR U2254 ( .A(n1609), .B(n1610), .Z(n1602) );
  XNOR U2255 ( .A(n1604), .B(n1603), .Z(n1610) );
  XNOR U2256 ( .A(y[171]), .B(x[171]), .Z(n1603) );
  XNOR U2257 ( .A(y[170]), .B(x[170]), .Z(n1604) );
  XNOR U2258 ( .A(n1607), .B(n1608), .Z(n1609) );
  XNOR U2259 ( .A(y[169]), .B(x[169]), .Z(n1608) );
  XNOR U2260 ( .A(y[168]), .B(x[168]), .Z(n1607) );
  XNOR U2261 ( .A(n1615), .B(n1616), .Z(n1624) );
  XNOR U2262 ( .A(n1619), .B(n1620), .Z(n1616) );
  XNOR U2263 ( .A(y[167]), .B(x[167]), .Z(n1620) );
  XNOR U2264 ( .A(y[166]), .B(x[166]), .Z(n1619) );
  XNOR U2265 ( .A(n1617), .B(n1618), .Z(n1615) );
  XNOR U2266 ( .A(y[165]), .B(x[165]), .Z(n1618) );
  XNOR U2267 ( .A(y[164]), .B(x[164]), .Z(n1617) );
  XNOR U2268 ( .A(n1632), .B(n1633), .Z(n1625) );
  XNOR U2269 ( .A(n1627), .B(n1626), .Z(n1633) );
  XNOR U2270 ( .A(y[163]), .B(x[163]), .Z(n1626) );
  XNOR U2271 ( .A(y[162]), .B(x[162]), .Z(n1627) );
  XNOR U2272 ( .A(n1630), .B(n1631), .Z(n1632) );
  XNOR U2273 ( .A(y[161]), .B(x[161]), .Z(n1631) );
  XNOR U2274 ( .A(y[160]), .B(x[160]), .Z(n1630) );
  XNOR U2275 ( .A(n1698), .B(n1697), .Z(n1677) );
  XNOR U2276 ( .A(n1664), .B(n1663), .Z(n1697) );
  XNOR U2277 ( .A(n1638), .B(n1639), .Z(n1645) );
  XNOR U2278 ( .A(n1642), .B(n1643), .Z(n1639) );
  XNOR U2279 ( .A(y[159]), .B(x[159]), .Z(n1643) );
  XNOR U2280 ( .A(y[158]), .B(x[158]), .Z(n1642) );
  XNOR U2281 ( .A(n1640), .B(n1641), .Z(n1638) );
  XNOR U2282 ( .A(y[157]), .B(x[157]), .Z(n1641) );
  XNOR U2283 ( .A(y[156]), .B(x[156]), .Z(n1640) );
  XNOR U2284 ( .A(n1653), .B(n1654), .Z(n1646) );
  XNOR U2285 ( .A(n1648), .B(n1647), .Z(n1654) );
  XNOR U2286 ( .A(y[155]), .B(x[155]), .Z(n1647) );
  XNOR U2287 ( .A(y[154]), .B(x[154]), .Z(n1648) );
  XNOR U2288 ( .A(n1651), .B(n1652), .Z(n1653) );
  XNOR U2289 ( .A(y[153]), .B(x[153]), .Z(n1652) );
  XNOR U2290 ( .A(y[152]), .B(x[152]), .Z(n1651) );
  XNOR U2291 ( .A(n1657), .B(n1658), .Z(n1666) );
  XNOR U2292 ( .A(n1661), .B(n1662), .Z(n1658) );
  XNOR U2293 ( .A(y[151]), .B(x[151]), .Z(n1662) );
  XNOR U2294 ( .A(y[150]), .B(x[150]), .Z(n1661) );
  XNOR U2295 ( .A(n1659), .B(n1660), .Z(n1657) );
  XNOR U2296 ( .A(y[149]), .B(x[149]), .Z(n1660) );
  XNOR U2297 ( .A(y[148]), .B(x[148]), .Z(n1659) );
  XNOR U2298 ( .A(n1674), .B(n1675), .Z(n1667) );
  XNOR U2299 ( .A(n1669), .B(n1668), .Z(n1675) );
  XNOR U2300 ( .A(y[147]), .B(x[147]), .Z(n1668) );
  XNOR U2301 ( .A(y[146]), .B(x[146]), .Z(n1669) );
  XNOR U2302 ( .A(n1672), .B(n1673), .Z(n1674) );
  XNOR U2303 ( .A(y[145]), .B(x[145]), .Z(n1673) );
  XNOR U2304 ( .A(y[144]), .B(x[144]), .Z(n1672) );
  XNOR U2305 ( .A(n1708), .B(n1707), .Z(n1698) );
  XNOR U2306 ( .A(n1680), .B(n1681), .Z(n1687) );
  XNOR U2307 ( .A(n1684), .B(n1685), .Z(n1681) );
  XNOR U2308 ( .A(y[143]), .B(x[143]), .Z(n1685) );
  XNOR U2309 ( .A(y[142]), .B(x[142]), .Z(n1684) );
  XNOR U2310 ( .A(n1682), .B(n1683), .Z(n1680) );
  XNOR U2311 ( .A(y[141]), .B(x[141]), .Z(n1683) );
  XNOR U2312 ( .A(y[140]), .B(x[140]), .Z(n1682) );
  XNOR U2313 ( .A(n1695), .B(n1696), .Z(n1688) );
  XNOR U2314 ( .A(n1690), .B(n1689), .Z(n1696) );
  XNOR U2315 ( .A(y[139]), .B(x[139]), .Z(n1689) );
  XNOR U2316 ( .A(y[138]), .B(x[138]), .Z(n1690) );
  XNOR U2317 ( .A(n1693), .B(n1694), .Z(n1695) );
  XNOR U2318 ( .A(y[137]), .B(x[137]), .Z(n1694) );
  XNOR U2319 ( .A(y[136]), .B(x[136]), .Z(n1693) );
  XNOR U2320 ( .A(n1701), .B(n1702), .Z(n1710) );
  XNOR U2321 ( .A(n1705), .B(n1706), .Z(n1702) );
  XNOR U2322 ( .A(y[135]), .B(x[135]), .Z(n1706) );
  XNOR U2323 ( .A(y[134]), .B(x[134]), .Z(n1705) );
  XNOR U2324 ( .A(n1703), .B(n1704), .Z(n1701) );
  XNOR U2325 ( .A(y[133]), .B(x[133]), .Z(n1704) );
  XNOR U2326 ( .A(y[132]), .B(x[132]), .Z(n1703) );
  XNOR U2327 ( .A(n1718), .B(n1719), .Z(n1711) );
  XNOR U2328 ( .A(n1713), .B(n1712), .Z(n1719) );
  XNOR U2329 ( .A(y[131]), .B(x[131]), .Z(n1712) );
  XNOR U2330 ( .A(y[130]), .B(x[130]), .Z(n1713) );
  XNOR U2331 ( .A(n1716), .B(n1717), .Z(n1718) );
  XNOR U2332 ( .A(y[129]), .B(x[129]), .Z(n1717) );
  XNOR U2333 ( .A(y[128]), .B(x[128]), .Z(n1716) );
  XNOR U2334 ( .A(n1971), .B(n1970), .Z(n1887) );
  XNOR U2335 ( .A(n1843), .B(n1842), .Z(n1970) );
  XNOR U2336 ( .A(n1780), .B(n1779), .Z(n1842) );
  XNOR U2337 ( .A(n1748), .B(n1747), .Z(n1779) );
  XNOR U2338 ( .A(n1722), .B(n1723), .Z(n1729) );
  XNOR U2339 ( .A(n1726), .B(n1727), .Z(n1723) );
  XNOR U2340 ( .A(y[127]), .B(x[127]), .Z(n1727) );
  XNOR U2341 ( .A(y[126]), .B(x[126]), .Z(n1726) );
  XNOR U2342 ( .A(n1724), .B(n1725), .Z(n1722) );
  XNOR U2343 ( .A(y[125]), .B(x[125]), .Z(n1725) );
  XNOR U2344 ( .A(y[124]), .B(x[124]), .Z(n1724) );
  XNOR U2345 ( .A(n1737), .B(n1738), .Z(n1730) );
  XNOR U2346 ( .A(n1732), .B(n1731), .Z(n1738) );
  XNOR U2347 ( .A(y[123]), .B(x[123]), .Z(n1731) );
  XNOR U2348 ( .A(y[122]), .B(x[122]), .Z(n1732) );
  XNOR U2349 ( .A(n1735), .B(n1736), .Z(n1737) );
  XNOR U2350 ( .A(y[121]), .B(x[121]), .Z(n1736) );
  XNOR U2351 ( .A(y[120]), .B(x[120]), .Z(n1735) );
  XNOR U2352 ( .A(n1741), .B(n1742), .Z(n1750) );
  XNOR U2353 ( .A(n1745), .B(n1746), .Z(n1742) );
  XNOR U2354 ( .A(y[119]), .B(x[119]), .Z(n1746) );
  XNOR U2355 ( .A(y[118]), .B(x[118]), .Z(n1745) );
  XNOR U2356 ( .A(n1743), .B(n1744), .Z(n1741) );
  XNOR U2357 ( .A(y[117]), .B(x[117]), .Z(n1744) );
  XNOR U2358 ( .A(y[116]), .B(x[116]), .Z(n1743) );
  XNOR U2359 ( .A(n1758), .B(n1759), .Z(n1751) );
  XNOR U2360 ( .A(n1753), .B(n1752), .Z(n1759) );
  XNOR U2361 ( .A(y[115]), .B(x[115]), .Z(n1752) );
  XNOR U2362 ( .A(y[114]), .B(x[114]), .Z(n1753) );
  XNOR U2363 ( .A(n1756), .B(n1757), .Z(n1758) );
  XNOR U2364 ( .A(y[113]), .B(x[113]), .Z(n1757) );
  XNOR U2365 ( .A(y[112]), .B(x[112]), .Z(n1756) );
  XNOR U2366 ( .A(n1790), .B(n1789), .Z(n1780) );
  XNOR U2367 ( .A(n1762), .B(n1763), .Z(n1769) );
  XNOR U2368 ( .A(n1766), .B(n1767), .Z(n1763) );
  XNOR U2369 ( .A(y[111]), .B(x[111]), .Z(n1767) );
  XNOR U2370 ( .A(y[110]), .B(x[110]), .Z(n1766) );
  XNOR U2371 ( .A(n1764), .B(n1765), .Z(n1762) );
  XNOR U2372 ( .A(y[109]), .B(x[109]), .Z(n1765) );
  XNOR U2373 ( .A(y[108]), .B(x[108]), .Z(n1764) );
  XNOR U2374 ( .A(n1777), .B(n1778), .Z(n1770) );
  XNOR U2375 ( .A(n1772), .B(n1771), .Z(n1778) );
  XNOR U2376 ( .A(y[107]), .B(x[107]), .Z(n1771) );
  XNOR U2377 ( .A(y[106]), .B(x[106]), .Z(n1772) );
  XNOR U2378 ( .A(n1775), .B(n1776), .Z(n1777) );
  XNOR U2379 ( .A(y[105]), .B(x[105]), .Z(n1776) );
  XNOR U2380 ( .A(y[104]), .B(x[104]), .Z(n1775) );
  XNOR U2381 ( .A(n1783), .B(n1784), .Z(n1792) );
  XNOR U2382 ( .A(n1787), .B(n1788), .Z(n1784) );
  XNOR U2383 ( .A(y[103]), .B(x[103]), .Z(n1788) );
  XNOR U2384 ( .A(y[102]), .B(x[102]), .Z(n1787) );
  XNOR U2385 ( .A(n1785), .B(n1786), .Z(n1783) );
  XNOR U2386 ( .A(y[101]), .B(x[101]), .Z(n1786) );
  XNOR U2387 ( .A(y[100]), .B(x[100]), .Z(n1785) );
  XNOR U2388 ( .A(n1800), .B(n1801), .Z(n1793) );
  XNOR U2389 ( .A(n1795), .B(n1794), .Z(n1801) );
  XNOR U2390 ( .A(y[99]), .B(x[99]), .Z(n1794) );
  XNOR U2391 ( .A(y[98]), .B(x[98]), .Z(n1795) );
  XNOR U2392 ( .A(n1798), .B(n1799), .Z(n1800) );
  XNOR U2393 ( .A(y[97]), .B(x[97]), .Z(n1799) );
  XNOR U2394 ( .A(y[96]), .B(x[96]), .Z(n1798) );
  XNOR U2395 ( .A(n1864), .B(n1863), .Z(n1843) );
  XNOR U2396 ( .A(n1830), .B(n1829), .Z(n1863) );
  XNOR U2397 ( .A(n1804), .B(n1805), .Z(n1811) );
  XNOR U2398 ( .A(n1808), .B(n1809), .Z(n1805) );
  XNOR U2399 ( .A(y[95]), .B(x[95]), .Z(n1809) );
  XNOR U2400 ( .A(y[94]), .B(x[94]), .Z(n1808) );
  XNOR U2401 ( .A(n1806), .B(n1807), .Z(n1804) );
  XNOR U2402 ( .A(y[93]), .B(x[93]), .Z(n1807) );
  XNOR U2403 ( .A(y[92]), .B(x[92]), .Z(n1806) );
  XNOR U2404 ( .A(n1819), .B(n1820), .Z(n1812) );
  XNOR U2405 ( .A(n1814), .B(n1813), .Z(n1820) );
  XNOR U2406 ( .A(y[91]), .B(x[91]), .Z(n1813) );
  XNOR U2407 ( .A(y[90]), .B(x[90]), .Z(n1814) );
  XNOR U2408 ( .A(n1817), .B(n1818), .Z(n1819) );
  XNOR U2409 ( .A(y[89]), .B(x[89]), .Z(n1818) );
  XNOR U2410 ( .A(y[88]), .B(x[88]), .Z(n1817) );
  XNOR U2411 ( .A(n1823), .B(n1824), .Z(n1832) );
  XNOR U2412 ( .A(n1827), .B(n1828), .Z(n1824) );
  XNOR U2413 ( .A(y[87]), .B(x[87]), .Z(n1828) );
  XNOR U2414 ( .A(y[86]), .B(x[86]), .Z(n1827) );
  XNOR U2415 ( .A(n1825), .B(n1826), .Z(n1823) );
  XNOR U2416 ( .A(y[85]), .B(x[85]), .Z(n1826) );
  XNOR U2417 ( .A(y[84]), .B(x[84]), .Z(n1825) );
  XNOR U2418 ( .A(n1840), .B(n1841), .Z(n1833) );
  XNOR U2419 ( .A(n1835), .B(n1834), .Z(n1841) );
  XNOR U2420 ( .A(y[83]), .B(x[83]), .Z(n1834) );
  XNOR U2421 ( .A(y[82]), .B(x[82]), .Z(n1835) );
  XNOR U2422 ( .A(n1838), .B(n1839), .Z(n1840) );
  XNOR U2423 ( .A(y[81]), .B(x[81]), .Z(n1839) );
  XNOR U2424 ( .A(y[80]), .B(x[80]), .Z(n1838) );
  XNOR U2425 ( .A(n1874), .B(n1873), .Z(n1864) );
  XNOR U2426 ( .A(n1846), .B(n1847), .Z(n1853) );
  XNOR U2427 ( .A(n1850), .B(n1851), .Z(n1847) );
  XNOR U2428 ( .A(y[79]), .B(x[79]), .Z(n1851) );
  XNOR U2429 ( .A(y[78]), .B(x[78]), .Z(n1850) );
  XNOR U2430 ( .A(n1848), .B(n1849), .Z(n1846) );
  XNOR U2431 ( .A(y[77]), .B(x[77]), .Z(n1849) );
  XNOR U2432 ( .A(y[76]), .B(x[76]), .Z(n1848) );
  XNOR U2433 ( .A(n1861), .B(n1862), .Z(n1854) );
  XNOR U2434 ( .A(n1856), .B(n1855), .Z(n1862) );
  XNOR U2435 ( .A(y[75]), .B(x[75]), .Z(n1855) );
  XNOR U2436 ( .A(y[74]), .B(x[74]), .Z(n1856) );
  XNOR U2437 ( .A(n1859), .B(n1860), .Z(n1861) );
  XNOR U2438 ( .A(y[73]), .B(x[73]), .Z(n1860) );
  XNOR U2439 ( .A(y[72]), .B(x[72]), .Z(n1859) );
  XNOR U2440 ( .A(n1867), .B(n1868), .Z(n1876) );
  XNOR U2441 ( .A(n1871), .B(n1872), .Z(n1868) );
  XNOR U2442 ( .A(y[71]), .B(x[71]), .Z(n1872) );
  XNOR U2443 ( .A(y[70]), .B(x[70]), .Z(n1871) );
  XNOR U2444 ( .A(n1869), .B(n1870), .Z(n1867) );
  XNOR U2445 ( .A(y[69]), .B(x[69]), .Z(n1870) );
  XNOR U2446 ( .A(y[68]), .B(x[68]), .Z(n1869) );
  XNOR U2447 ( .A(n1884), .B(n1885), .Z(n1877) );
  XNOR U2448 ( .A(n1879), .B(n1878), .Z(n1885) );
  XNOR U2449 ( .A(y[67]), .B(x[67]), .Z(n1878) );
  XNOR U2450 ( .A(y[66]), .B(x[66]), .Z(n1879) );
  XNOR U2451 ( .A(n1882), .B(n1883), .Z(n1884) );
  XNOR U2452 ( .A(y[65]), .B(x[65]), .Z(n1883) );
  XNOR U2453 ( .A(y[64]), .B(x[64]), .Z(n1882) );
  XNOR U2454 ( .A(n2013), .B(n2012), .Z(n1971) );
  XNOR U2455 ( .A(n1948), .B(n1947), .Z(n2012) );
  XNOR U2456 ( .A(n1916), .B(n1915), .Z(n1947) );
  XNOR U2457 ( .A(n1890), .B(n1891), .Z(n1897) );
  XNOR U2458 ( .A(n1894), .B(n1895), .Z(n1891) );
  XNOR U2459 ( .A(y[63]), .B(x[63]), .Z(n1895) );
  XNOR U2460 ( .A(y[62]), .B(x[62]), .Z(n1894) );
  XNOR U2461 ( .A(n1892), .B(n1893), .Z(n1890) );
  XNOR U2462 ( .A(y[61]), .B(x[61]), .Z(n1893) );
  XNOR U2463 ( .A(y[60]), .B(x[60]), .Z(n1892) );
  XNOR U2464 ( .A(n1905), .B(n1906), .Z(n1898) );
  XNOR U2465 ( .A(n1900), .B(n1899), .Z(n1906) );
  XNOR U2466 ( .A(y[59]), .B(x[59]), .Z(n1899) );
  XNOR U2467 ( .A(y[58]), .B(x[58]), .Z(n1900) );
  XNOR U2468 ( .A(n1903), .B(n1904), .Z(n1905) );
  XNOR U2469 ( .A(y[57]), .B(x[57]), .Z(n1904) );
  XNOR U2470 ( .A(y[56]), .B(x[56]), .Z(n1903) );
  XNOR U2471 ( .A(n1909), .B(n1910), .Z(n1918) );
  XNOR U2472 ( .A(n1913), .B(n1914), .Z(n1910) );
  XNOR U2473 ( .A(y[55]), .B(x[55]), .Z(n1914) );
  XNOR U2474 ( .A(y[54]), .B(x[54]), .Z(n1913) );
  XNOR U2475 ( .A(n1911), .B(n1912), .Z(n1909) );
  XNOR U2476 ( .A(y[53]), .B(x[53]), .Z(n1912) );
  XNOR U2477 ( .A(y[52]), .B(x[52]), .Z(n1911) );
  XNOR U2478 ( .A(n1926), .B(n1927), .Z(n1919) );
  XNOR U2479 ( .A(n1921), .B(n1920), .Z(n1927) );
  XNOR U2480 ( .A(y[51]), .B(x[51]), .Z(n1920) );
  XNOR U2481 ( .A(y[50]), .B(x[50]), .Z(n1921) );
  XNOR U2482 ( .A(n1924), .B(n1925), .Z(n1926) );
  XNOR U2483 ( .A(y[49]), .B(x[49]), .Z(n1925) );
  XNOR U2484 ( .A(y[48]), .B(x[48]), .Z(n1924) );
  XNOR U2485 ( .A(n1958), .B(n1957), .Z(n1948) );
  XNOR U2486 ( .A(n1930), .B(n1931), .Z(n1937) );
  XNOR U2487 ( .A(n1934), .B(n1935), .Z(n1931) );
  XNOR U2488 ( .A(y[47]), .B(x[47]), .Z(n1935) );
  XNOR U2489 ( .A(y[46]), .B(x[46]), .Z(n1934) );
  XNOR U2490 ( .A(n1932), .B(n1933), .Z(n1930) );
  XNOR U2491 ( .A(y[45]), .B(x[45]), .Z(n1933) );
  XNOR U2492 ( .A(y[44]), .B(x[44]), .Z(n1932) );
  XNOR U2493 ( .A(n1945), .B(n1946), .Z(n1938) );
  XNOR U2494 ( .A(n1940), .B(n1939), .Z(n1946) );
  XNOR U2495 ( .A(y[43]), .B(x[43]), .Z(n1939) );
  XNOR U2496 ( .A(y[42]), .B(x[42]), .Z(n1940) );
  XNOR U2497 ( .A(n1943), .B(n1944), .Z(n1945) );
  XNOR U2498 ( .A(y[41]), .B(x[41]), .Z(n1944) );
  XNOR U2499 ( .A(y[40]), .B(x[40]), .Z(n1943) );
  XNOR U2500 ( .A(n1951), .B(n1952), .Z(n1960) );
  XNOR U2501 ( .A(n1955), .B(n1956), .Z(n1952) );
  XNOR U2502 ( .A(y[39]), .B(x[39]), .Z(n1956) );
  XNOR U2503 ( .A(y[38]), .B(x[38]), .Z(n1955) );
  XNOR U2504 ( .A(n1953), .B(n1954), .Z(n1951) );
  XNOR U2505 ( .A(y[37]), .B(x[37]), .Z(n1954) );
  XNOR U2506 ( .A(y[36]), .B(x[36]), .Z(n1953) );
  XNOR U2507 ( .A(n1968), .B(n1969), .Z(n1961) );
  XNOR U2508 ( .A(n1963), .B(n1962), .Z(n1969) );
  XNOR U2509 ( .A(y[35]), .B(x[35]), .Z(n1962) );
  XNOR U2510 ( .A(y[34]), .B(x[34]), .Z(n1963) );
  XNOR U2511 ( .A(n1966), .B(n1967), .Z(n1968) );
  XNOR U2512 ( .A(y[33]), .B(x[33]), .Z(n1967) );
  XNOR U2513 ( .A(y[32]), .B(x[32]), .Z(n1966) );
  XNOR U2514 ( .A(n2034), .B(n2033), .Z(n2013) );
  XNOR U2515 ( .A(n2000), .B(n1999), .Z(n2033) );
  XNOR U2516 ( .A(n1974), .B(n1975), .Z(n1981) );
  XNOR U2517 ( .A(n1978), .B(n1979), .Z(n1975) );
  XNOR U2518 ( .A(y[31]), .B(x[31]), .Z(n1979) );
  XNOR U2519 ( .A(y[30]), .B(x[30]), .Z(n1978) );
  XNOR U2520 ( .A(n1976), .B(n1977), .Z(n1974) );
  XNOR U2521 ( .A(y[29]), .B(x[29]), .Z(n1977) );
  XNOR U2522 ( .A(y[28]), .B(x[28]), .Z(n1976) );
  XNOR U2523 ( .A(n1989), .B(n1990), .Z(n1982) );
  XNOR U2524 ( .A(n1984), .B(n1983), .Z(n1990) );
  XNOR U2525 ( .A(y[27]), .B(x[27]), .Z(n1983) );
  XNOR U2526 ( .A(y[26]), .B(x[26]), .Z(n1984) );
  XNOR U2527 ( .A(n1987), .B(n1988), .Z(n1989) );
  XNOR U2528 ( .A(y[25]), .B(x[25]), .Z(n1988) );
  XNOR U2529 ( .A(y[24]), .B(x[24]), .Z(n1987) );
  XNOR U2530 ( .A(n1993), .B(n1994), .Z(n2002) );
  XNOR U2531 ( .A(n1997), .B(n1998), .Z(n1994) );
  XNOR U2532 ( .A(y[23]), .B(x[23]), .Z(n1998) );
  XNOR U2533 ( .A(y[22]), .B(x[22]), .Z(n1997) );
  XNOR U2534 ( .A(n1995), .B(n1996), .Z(n1993) );
  XNOR U2535 ( .A(y[21]), .B(x[21]), .Z(n1996) );
  XNOR U2536 ( .A(y[20]), .B(x[20]), .Z(n1995) );
  XNOR U2537 ( .A(n2010), .B(n2011), .Z(n2003) );
  XNOR U2538 ( .A(n2005), .B(n2004), .Z(n2011) );
  XNOR U2539 ( .A(y[19]), .B(x[19]), .Z(n2004) );
  XNOR U2540 ( .A(y[18]), .B(x[18]), .Z(n2005) );
  XNOR U2541 ( .A(n2008), .B(n2009), .Z(n2010) );
  XNOR U2542 ( .A(y[17]), .B(x[17]), .Z(n2009) );
  XNOR U2543 ( .A(y[16]), .B(x[16]), .Z(n2008) );
  XNOR U2544 ( .A(n2044), .B(n2043), .Z(n2034) );
  XNOR U2545 ( .A(n2016), .B(n2017), .Z(n2023) );
  XNOR U2546 ( .A(n2020), .B(n2021), .Z(n2017) );
  XNOR U2547 ( .A(y[15]), .B(x[15]), .Z(n2021) );
  XNOR U2548 ( .A(y[14]), .B(x[14]), .Z(n2020) );
  XNOR U2549 ( .A(n2018), .B(n2019), .Z(n2016) );
  XNOR U2550 ( .A(y[13]), .B(x[13]), .Z(n2019) );
  XNOR U2551 ( .A(y[12]), .B(x[12]), .Z(n2018) );
  XNOR U2552 ( .A(n2031), .B(n2032), .Z(n2024) );
  XNOR U2553 ( .A(n2026), .B(n2025), .Z(n2032) );
  XNOR U2554 ( .A(y[11]), .B(x[11]), .Z(n2025) );
  XNOR U2555 ( .A(y[10]), .B(x[10]), .Z(n2026) );
  XNOR U2556 ( .A(n2029), .B(n2030), .Z(n2031) );
  XNOR U2557 ( .A(y[9]), .B(x[9]), .Z(n2030) );
  XNOR U2558 ( .A(y[8]), .B(x[8]), .Z(n2029) );
  XNOR U2559 ( .A(n2037), .B(n2038), .Z(n2046) );
  XNOR U2560 ( .A(n2041), .B(n2042), .Z(n2038) );
  XNOR U2561 ( .A(y[7]), .B(x[7]), .Z(n2042) );
  XNOR U2562 ( .A(y[6]), .B(x[6]), .Z(n2041) );
  XNOR U2563 ( .A(n2039), .B(n2040), .Z(n2037) );
  XNOR U2564 ( .A(y[5]), .B(x[5]), .Z(n2040) );
  XNOR U2565 ( .A(y[4]), .B(x[4]), .Z(n2039) );
  XNOR U2566 ( .A(n2054), .B(n2055), .Z(n2047) );
  XNOR U2567 ( .A(n2049), .B(n2048), .Z(n2055) );
  XNOR U2568 ( .A(y[3]), .B(x[3]), .Z(n2048) );
  XNOR U2569 ( .A(y[2]), .B(x[2]), .Z(n2049) );
  XNOR U2570 ( .A(n2052), .B(n2053), .Z(n2054) );
  XNOR U2571 ( .A(y[1]), .B(x[1]), .Z(n2053) );
  XNOR U2572 ( .A(y[0]), .B(x[0]), .Z(n2052) );
endmodule

