
module mult_N1024_CC1024 ( clk, rst, a, b, c );
  input [1023:0] a;
  input [0:0] b;
  output [2047:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183;
  wire   [2047:0] sreg;

  DFF \sreg_reg[2046]  ( .D(c[2047]), .CLK(clk), .RST(rst), .Q(sreg[2046]) );
  DFF \sreg_reg[2045]  ( .D(c[2046]), .CLK(clk), .RST(rst), .Q(sreg[2045]) );
  DFF \sreg_reg[2044]  ( .D(c[2045]), .CLK(clk), .RST(rst), .Q(sreg[2044]) );
  DFF \sreg_reg[2043]  ( .D(c[2044]), .CLK(clk), .RST(rst), .Q(sreg[2043]) );
  DFF \sreg_reg[2042]  ( .D(c[2043]), .CLK(clk), .RST(rst), .Q(sreg[2042]) );
  DFF \sreg_reg[2041]  ( .D(c[2042]), .CLK(clk), .RST(rst), .Q(sreg[2041]) );
  DFF \sreg_reg[2040]  ( .D(c[2041]), .CLK(clk), .RST(rst), .Q(sreg[2040]) );
  DFF \sreg_reg[2039]  ( .D(c[2040]), .CLK(clk), .RST(rst), .Q(sreg[2039]) );
  DFF \sreg_reg[2038]  ( .D(c[2039]), .CLK(clk), .RST(rst), .Q(sreg[2038]) );
  DFF \sreg_reg[2037]  ( .D(c[2038]), .CLK(clk), .RST(rst), .Q(sreg[2037]) );
  DFF \sreg_reg[2036]  ( .D(c[2037]), .CLK(clk), .RST(rst), .Q(sreg[2036]) );
  DFF \sreg_reg[2035]  ( .D(c[2036]), .CLK(clk), .RST(rst), .Q(sreg[2035]) );
  DFF \sreg_reg[2034]  ( .D(c[2035]), .CLK(clk), .RST(rst), .Q(sreg[2034]) );
  DFF \sreg_reg[2033]  ( .D(c[2034]), .CLK(clk), .RST(rst), .Q(sreg[2033]) );
  DFF \sreg_reg[2032]  ( .D(c[2033]), .CLK(clk), .RST(rst), .Q(sreg[2032]) );
  DFF \sreg_reg[2031]  ( .D(c[2032]), .CLK(clk), .RST(rst), .Q(sreg[2031]) );
  DFF \sreg_reg[2030]  ( .D(c[2031]), .CLK(clk), .RST(rst), .Q(sreg[2030]) );
  DFF \sreg_reg[2029]  ( .D(c[2030]), .CLK(clk), .RST(rst), .Q(sreg[2029]) );
  DFF \sreg_reg[2028]  ( .D(c[2029]), .CLK(clk), .RST(rst), .Q(sreg[2028]) );
  DFF \sreg_reg[2027]  ( .D(c[2028]), .CLK(clk), .RST(rst), .Q(sreg[2027]) );
  DFF \sreg_reg[2026]  ( .D(c[2027]), .CLK(clk), .RST(rst), .Q(sreg[2026]) );
  DFF \sreg_reg[2025]  ( .D(c[2026]), .CLK(clk), .RST(rst), .Q(sreg[2025]) );
  DFF \sreg_reg[2024]  ( .D(c[2025]), .CLK(clk), .RST(rst), .Q(sreg[2024]) );
  DFF \sreg_reg[2023]  ( .D(c[2024]), .CLK(clk), .RST(rst), .Q(sreg[2023]) );
  DFF \sreg_reg[2022]  ( .D(c[2023]), .CLK(clk), .RST(rst), .Q(sreg[2022]) );
  DFF \sreg_reg[2021]  ( .D(c[2022]), .CLK(clk), .RST(rst), .Q(sreg[2021]) );
  DFF \sreg_reg[2020]  ( .D(c[2021]), .CLK(clk), .RST(rst), .Q(sreg[2020]) );
  DFF \sreg_reg[2019]  ( .D(c[2020]), .CLK(clk), .RST(rst), .Q(sreg[2019]) );
  DFF \sreg_reg[2018]  ( .D(c[2019]), .CLK(clk), .RST(rst), .Q(sreg[2018]) );
  DFF \sreg_reg[2017]  ( .D(c[2018]), .CLK(clk), .RST(rst), .Q(sreg[2017]) );
  DFF \sreg_reg[2016]  ( .D(c[2017]), .CLK(clk), .RST(rst), .Q(sreg[2016]) );
  DFF \sreg_reg[2015]  ( .D(c[2016]), .CLK(clk), .RST(rst), .Q(sreg[2015]) );
  DFF \sreg_reg[2014]  ( .D(c[2015]), .CLK(clk), .RST(rst), .Q(sreg[2014]) );
  DFF \sreg_reg[2013]  ( .D(c[2014]), .CLK(clk), .RST(rst), .Q(sreg[2013]) );
  DFF \sreg_reg[2012]  ( .D(c[2013]), .CLK(clk), .RST(rst), .Q(sreg[2012]) );
  DFF \sreg_reg[2011]  ( .D(c[2012]), .CLK(clk), .RST(rst), .Q(sreg[2011]) );
  DFF \sreg_reg[2010]  ( .D(c[2011]), .CLK(clk), .RST(rst), .Q(sreg[2010]) );
  DFF \sreg_reg[2009]  ( .D(c[2010]), .CLK(clk), .RST(rst), .Q(sreg[2009]) );
  DFF \sreg_reg[2008]  ( .D(c[2009]), .CLK(clk), .RST(rst), .Q(sreg[2008]) );
  DFF \sreg_reg[2007]  ( .D(c[2008]), .CLK(clk), .RST(rst), .Q(sreg[2007]) );
  DFF \sreg_reg[2006]  ( .D(c[2007]), .CLK(clk), .RST(rst), .Q(sreg[2006]) );
  DFF \sreg_reg[2005]  ( .D(c[2006]), .CLK(clk), .RST(rst), .Q(sreg[2005]) );
  DFF \sreg_reg[2004]  ( .D(c[2005]), .CLK(clk), .RST(rst), .Q(sreg[2004]) );
  DFF \sreg_reg[2003]  ( .D(c[2004]), .CLK(clk), .RST(rst), .Q(sreg[2003]) );
  DFF \sreg_reg[2002]  ( .D(c[2003]), .CLK(clk), .RST(rst), .Q(sreg[2002]) );
  DFF \sreg_reg[2001]  ( .D(c[2002]), .CLK(clk), .RST(rst), .Q(sreg[2001]) );
  DFF \sreg_reg[2000]  ( .D(c[2001]), .CLK(clk), .RST(rst), .Q(sreg[2000]) );
  DFF \sreg_reg[1999]  ( .D(c[2000]), .CLK(clk), .RST(rst), .Q(sreg[1999]) );
  DFF \sreg_reg[1998]  ( .D(c[1999]), .CLK(clk), .RST(rst), .Q(sreg[1998]) );
  DFF \sreg_reg[1997]  ( .D(c[1998]), .CLK(clk), .RST(rst), .Q(sreg[1997]) );
  DFF \sreg_reg[1996]  ( .D(c[1997]), .CLK(clk), .RST(rst), .Q(sreg[1996]) );
  DFF \sreg_reg[1995]  ( .D(c[1996]), .CLK(clk), .RST(rst), .Q(sreg[1995]) );
  DFF \sreg_reg[1994]  ( .D(c[1995]), .CLK(clk), .RST(rst), .Q(sreg[1994]) );
  DFF \sreg_reg[1993]  ( .D(c[1994]), .CLK(clk), .RST(rst), .Q(sreg[1993]) );
  DFF \sreg_reg[1992]  ( .D(c[1993]), .CLK(clk), .RST(rst), .Q(sreg[1992]) );
  DFF \sreg_reg[1991]  ( .D(c[1992]), .CLK(clk), .RST(rst), .Q(sreg[1991]) );
  DFF \sreg_reg[1990]  ( .D(c[1991]), .CLK(clk), .RST(rst), .Q(sreg[1990]) );
  DFF \sreg_reg[1989]  ( .D(c[1990]), .CLK(clk), .RST(rst), .Q(sreg[1989]) );
  DFF \sreg_reg[1988]  ( .D(c[1989]), .CLK(clk), .RST(rst), .Q(sreg[1988]) );
  DFF \sreg_reg[1987]  ( .D(c[1988]), .CLK(clk), .RST(rst), .Q(sreg[1987]) );
  DFF \sreg_reg[1986]  ( .D(c[1987]), .CLK(clk), .RST(rst), .Q(sreg[1986]) );
  DFF \sreg_reg[1985]  ( .D(c[1986]), .CLK(clk), .RST(rst), .Q(sreg[1985]) );
  DFF \sreg_reg[1984]  ( .D(c[1985]), .CLK(clk), .RST(rst), .Q(sreg[1984]) );
  DFF \sreg_reg[1983]  ( .D(c[1984]), .CLK(clk), .RST(rst), .Q(sreg[1983]) );
  DFF \sreg_reg[1982]  ( .D(c[1983]), .CLK(clk), .RST(rst), .Q(sreg[1982]) );
  DFF \sreg_reg[1981]  ( .D(c[1982]), .CLK(clk), .RST(rst), .Q(sreg[1981]) );
  DFF \sreg_reg[1980]  ( .D(c[1981]), .CLK(clk), .RST(rst), .Q(sreg[1980]) );
  DFF \sreg_reg[1979]  ( .D(c[1980]), .CLK(clk), .RST(rst), .Q(sreg[1979]) );
  DFF \sreg_reg[1978]  ( .D(c[1979]), .CLK(clk), .RST(rst), .Q(sreg[1978]) );
  DFF \sreg_reg[1977]  ( .D(c[1978]), .CLK(clk), .RST(rst), .Q(sreg[1977]) );
  DFF \sreg_reg[1976]  ( .D(c[1977]), .CLK(clk), .RST(rst), .Q(sreg[1976]) );
  DFF \sreg_reg[1975]  ( .D(c[1976]), .CLK(clk), .RST(rst), .Q(sreg[1975]) );
  DFF \sreg_reg[1974]  ( .D(c[1975]), .CLK(clk), .RST(rst), .Q(sreg[1974]) );
  DFF \sreg_reg[1973]  ( .D(c[1974]), .CLK(clk), .RST(rst), .Q(sreg[1973]) );
  DFF \sreg_reg[1972]  ( .D(c[1973]), .CLK(clk), .RST(rst), .Q(sreg[1972]) );
  DFF \sreg_reg[1971]  ( .D(c[1972]), .CLK(clk), .RST(rst), .Q(sreg[1971]) );
  DFF \sreg_reg[1970]  ( .D(c[1971]), .CLK(clk), .RST(rst), .Q(sreg[1970]) );
  DFF \sreg_reg[1969]  ( .D(c[1970]), .CLK(clk), .RST(rst), .Q(sreg[1969]) );
  DFF \sreg_reg[1968]  ( .D(c[1969]), .CLK(clk), .RST(rst), .Q(sreg[1968]) );
  DFF \sreg_reg[1967]  ( .D(c[1968]), .CLK(clk), .RST(rst), .Q(sreg[1967]) );
  DFF \sreg_reg[1966]  ( .D(c[1967]), .CLK(clk), .RST(rst), .Q(sreg[1966]) );
  DFF \sreg_reg[1965]  ( .D(c[1966]), .CLK(clk), .RST(rst), .Q(sreg[1965]) );
  DFF \sreg_reg[1964]  ( .D(c[1965]), .CLK(clk), .RST(rst), .Q(sreg[1964]) );
  DFF \sreg_reg[1963]  ( .D(c[1964]), .CLK(clk), .RST(rst), .Q(sreg[1963]) );
  DFF \sreg_reg[1962]  ( .D(c[1963]), .CLK(clk), .RST(rst), .Q(sreg[1962]) );
  DFF \sreg_reg[1961]  ( .D(c[1962]), .CLK(clk), .RST(rst), .Q(sreg[1961]) );
  DFF \sreg_reg[1960]  ( .D(c[1961]), .CLK(clk), .RST(rst), .Q(sreg[1960]) );
  DFF \sreg_reg[1959]  ( .D(c[1960]), .CLK(clk), .RST(rst), .Q(sreg[1959]) );
  DFF \sreg_reg[1958]  ( .D(c[1959]), .CLK(clk), .RST(rst), .Q(sreg[1958]) );
  DFF \sreg_reg[1957]  ( .D(c[1958]), .CLK(clk), .RST(rst), .Q(sreg[1957]) );
  DFF \sreg_reg[1956]  ( .D(c[1957]), .CLK(clk), .RST(rst), .Q(sreg[1956]) );
  DFF \sreg_reg[1955]  ( .D(c[1956]), .CLK(clk), .RST(rst), .Q(sreg[1955]) );
  DFF \sreg_reg[1954]  ( .D(c[1955]), .CLK(clk), .RST(rst), .Q(sreg[1954]) );
  DFF \sreg_reg[1953]  ( .D(c[1954]), .CLK(clk), .RST(rst), .Q(sreg[1953]) );
  DFF \sreg_reg[1952]  ( .D(c[1953]), .CLK(clk), .RST(rst), .Q(sreg[1952]) );
  DFF \sreg_reg[1951]  ( .D(c[1952]), .CLK(clk), .RST(rst), .Q(sreg[1951]) );
  DFF \sreg_reg[1950]  ( .D(c[1951]), .CLK(clk), .RST(rst), .Q(sreg[1950]) );
  DFF \sreg_reg[1949]  ( .D(c[1950]), .CLK(clk), .RST(rst), .Q(sreg[1949]) );
  DFF \sreg_reg[1948]  ( .D(c[1949]), .CLK(clk), .RST(rst), .Q(sreg[1948]) );
  DFF \sreg_reg[1947]  ( .D(c[1948]), .CLK(clk), .RST(rst), .Q(sreg[1947]) );
  DFF \sreg_reg[1946]  ( .D(c[1947]), .CLK(clk), .RST(rst), .Q(sreg[1946]) );
  DFF \sreg_reg[1945]  ( .D(c[1946]), .CLK(clk), .RST(rst), .Q(sreg[1945]) );
  DFF \sreg_reg[1944]  ( .D(c[1945]), .CLK(clk), .RST(rst), .Q(sreg[1944]) );
  DFF \sreg_reg[1943]  ( .D(c[1944]), .CLK(clk), .RST(rst), .Q(sreg[1943]) );
  DFF \sreg_reg[1942]  ( .D(c[1943]), .CLK(clk), .RST(rst), .Q(sreg[1942]) );
  DFF \sreg_reg[1941]  ( .D(c[1942]), .CLK(clk), .RST(rst), .Q(sreg[1941]) );
  DFF \sreg_reg[1940]  ( .D(c[1941]), .CLK(clk), .RST(rst), .Q(sreg[1940]) );
  DFF \sreg_reg[1939]  ( .D(c[1940]), .CLK(clk), .RST(rst), .Q(sreg[1939]) );
  DFF \sreg_reg[1938]  ( .D(c[1939]), .CLK(clk), .RST(rst), .Q(sreg[1938]) );
  DFF \sreg_reg[1937]  ( .D(c[1938]), .CLK(clk), .RST(rst), .Q(sreg[1937]) );
  DFF \sreg_reg[1936]  ( .D(c[1937]), .CLK(clk), .RST(rst), .Q(sreg[1936]) );
  DFF \sreg_reg[1935]  ( .D(c[1936]), .CLK(clk), .RST(rst), .Q(sreg[1935]) );
  DFF \sreg_reg[1934]  ( .D(c[1935]), .CLK(clk), .RST(rst), .Q(sreg[1934]) );
  DFF \sreg_reg[1933]  ( .D(c[1934]), .CLK(clk), .RST(rst), .Q(sreg[1933]) );
  DFF \sreg_reg[1932]  ( .D(c[1933]), .CLK(clk), .RST(rst), .Q(sreg[1932]) );
  DFF \sreg_reg[1931]  ( .D(c[1932]), .CLK(clk), .RST(rst), .Q(sreg[1931]) );
  DFF \sreg_reg[1930]  ( .D(c[1931]), .CLK(clk), .RST(rst), .Q(sreg[1930]) );
  DFF \sreg_reg[1929]  ( .D(c[1930]), .CLK(clk), .RST(rst), .Q(sreg[1929]) );
  DFF \sreg_reg[1928]  ( .D(c[1929]), .CLK(clk), .RST(rst), .Q(sreg[1928]) );
  DFF \sreg_reg[1927]  ( .D(c[1928]), .CLK(clk), .RST(rst), .Q(sreg[1927]) );
  DFF \sreg_reg[1926]  ( .D(c[1927]), .CLK(clk), .RST(rst), .Q(sreg[1926]) );
  DFF \sreg_reg[1925]  ( .D(c[1926]), .CLK(clk), .RST(rst), .Q(sreg[1925]) );
  DFF \sreg_reg[1924]  ( .D(c[1925]), .CLK(clk), .RST(rst), .Q(sreg[1924]) );
  DFF \sreg_reg[1923]  ( .D(c[1924]), .CLK(clk), .RST(rst), .Q(sreg[1923]) );
  DFF \sreg_reg[1922]  ( .D(c[1923]), .CLK(clk), .RST(rst), .Q(sreg[1922]) );
  DFF \sreg_reg[1921]  ( .D(c[1922]), .CLK(clk), .RST(rst), .Q(sreg[1921]) );
  DFF \sreg_reg[1920]  ( .D(c[1921]), .CLK(clk), .RST(rst), .Q(sreg[1920]) );
  DFF \sreg_reg[1919]  ( .D(c[1920]), .CLK(clk), .RST(rst), .Q(sreg[1919]) );
  DFF \sreg_reg[1918]  ( .D(c[1919]), .CLK(clk), .RST(rst), .Q(sreg[1918]) );
  DFF \sreg_reg[1917]  ( .D(c[1918]), .CLK(clk), .RST(rst), .Q(sreg[1917]) );
  DFF \sreg_reg[1916]  ( .D(c[1917]), .CLK(clk), .RST(rst), .Q(sreg[1916]) );
  DFF \sreg_reg[1915]  ( .D(c[1916]), .CLK(clk), .RST(rst), .Q(sreg[1915]) );
  DFF \sreg_reg[1914]  ( .D(c[1915]), .CLK(clk), .RST(rst), .Q(sreg[1914]) );
  DFF \sreg_reg[1913]  ( .D(c[1914]), .CLK(clk), .RST(rst), .Q(sreg[1913]) );
  DFF \sreg_reg[1912]  ( .D(c[1913]), .CLK(clk), .RST(rst), .Q(sreg[1912]) );
  DFF \sreg_reg[1911]  ( .D(c[1912]), .CLK(clk), .RST(rst), .Q(sreg[1911]) );
  DFF \sreg_reg[1910]  ( .D(c[1911]), .CLK(clk), .RST(rst), .Q(sreg[1910]) );
  DFF \sreg_reg[1909]  ( .D(c[1910]), .CLK(clk), .RST(rst), .Q(sreg[1909]) );
  DFF \sreg_reg[1908]  ( .D(c[1909]), .CLK(clk), .RST(rst), .Q(sreg[1908]) );
  DFF \sreg_reg[1907]  ( .D(c[1908]), .CLK(clk), .RST(rst), .Q(sreg[1907]) );
  DFF \sreg_reg[1906]  ( .D(c[1907]), .CLK(clk), .RST(rst), .Q(sreg[1906]) );
  DFF \sreg_reg[1905]  ( .D(c[1906]), .CLK(clk), .RST(rst), .Q(sreg[1905]) );
  DFF \sreg_reg[1904]  ( .D(c[1905]), .CLK(clk), .RST(rst), .Q(sreg[1904]) );
  DFF \sreg_reg[1903]  ( .D(c[1904]), .CLK(clk), .RST(rst), .Q(sreg[1903]) );
  DFF \sreg_reg[1902]  ( .D(c[1903]), .CLK(clk), .RST(rst), .Q(sreg[1902]) );
  DFF \sreg_reg[1901]  ( .D(c[1902]), .CLK(clk), .RST(rst), .Q(sreg[1901]) );
  DFF \sreg_reg[1900]  ( .D(c[1901]), .CLK(clk), .RST(rst), .Q(sreg[1900]) );
  DFF \sreg_reg[1899]  ( .D(c[1900]), .CLK(clk), .RST(rst), .Q(sreg[1899]) );
  DFF \sreg_reg[1898]  ( .D(c[1899]), .CLK(clk), .RST(rst), .Q(sreg[1898]) );
  DFF \sreg_reg[1897]  ( .D(c[1898]), .CLK(clk), .RST(rst), .Q(sreg[1897]) );
  DFF \sreg_reg[1896]  ( .D(c[1897]), .CLK(clk), .RST(rst), .Q(sreg[1896]) );
  DFF \sreg_reg[1895]  ( .D(c[1896]), .CLK(clk), .RST(rst), .Q(sreg[1895]) );
  DFF \sreg_reg[1894]  ( .D(c[1895]), .CLK(clk), .RST(rst), .Q(sreg[1894]) );
  DFF \sreg_reg[1893]  ( .D(c[1894]), .CLK(clk), .RST(rst), .Q(sreg[1893]) );
  DFF \sreg_reg[1892]  ( .D(c[1893]), .CLK(clk), .RST(rst), .Q(sreg[1892]) );
  DFF \sreg_reg[1891]  ( .D(c[1892]), .CLK(clk), .RST(rst), .Q(sreg[1891]) );
  DFF \sreg_reg[1890]  ( .D(c[1891]), .CLK(clk), .RST(rst), .Q(sreg[1890]) );
  DFF \sreg_reg[1889]  ( .D(c[1890]), .CLK(clk), .RST(rst), .Q(sreg[1889]) );
  DFF \sreg_reg[1888]  ( .D(c[1889]), .CLK(clk), .RST(rst), .Q(sreg[1888]) );
  DFF \sreg_reg[1887]  ( .D(c[1888]), .CLK(clk), .RST(rst), .Q(sreg[1887]) );
  DFF \sreg_reg[1886]  ( .D(c[1887]), .CLK(clk), .RST(rst), .Q(sreg[1886]) );
  DFF \sreg_reg[1885]  ( .D(c[1886]), .CLK(clk), .RST(rst), .Q(sreg[1885]) );
  DFF \sreg_reg[1884]  ( .D(c[1885]), .CLK(clk), .RST(rst), .Q(sreg[1884]) );
  DFF \sreg_reg[1883]  ( .D(c[1884]), .CLK(clk), .RST(rst), .Q(sreg[1883]) );
  DFF \sreg_reg[1882]  ( .D(c[1883]), .CLK(clk), .RST(rst), .Q(sreg[1882]) );
  DFF \sreg_reg[1881]  ( .D(c[1882]), .CLK(clk), .RST(rst), .Q(sreg[1881]) );
  DFF \sreg_reg[1880]  ( .D(c[1881]), .CLK(clk), .RST(rst), .Q(sreg[1880]) );
  DFF \sreg_reg[1879]  ( .D(c[1880]), .CLK(clk), .RST(rst), .Q(sreg[1879]) );
  DFF \sreg_reg[1878]  ( .D(c[1879]), .CLK(clk), .RST(rst), .Q(sreg[1878]) );
  DFF \sreg_reg[1877]  ( .D(c[1878]), .CLK(clk), .RST(rst), .Q(sreg[1877]) );
  DFF \sreg_reg[1876]  ( .D(c[1877]), .CLK(clk), .RST(rst), .Q(sreg[1876]) );
  DFF \sreg_reg[1875]  ( .D(c[1876]), .CLK(clk), .RST(rst), .Q(sreg[1875]) );
  DFF \sreg_reg[1874]  ( .D(c[1875]), .CLK(clk), .RST(rst), .Q(sreg[1874]) );
  DFF \sreg_reg[1873]  ( .D(c[1874]), .CLK(clk), .RST(rst), .Q(sreg[1873]) );
  DFF \sreg_reg[1872]  ( .D(c[1873]), .CLK(clk), .RST(rst), .Q(sreg[1872]) );
  DFF \sreg_reg[1871]  ( .D(c[1872]), .CLK(clk), .RST(rst), .Q(sreg[1871]) );
  DFF \sreg_reg[1870]  ( .D(c[1871]), .CLK(clk), .RST(rst), .Q(sreg[1870]) );
  DFF \sreg_reg[1869]  ( .D(c[1870]), .CLK(clk), .RST(rst), .Q(sreg[1869]) );
  DFF \sreg_reg[1868]  ( .D(c[1869]), .CLK(clk), .RST(rst), .Q(sreg[1868]) );
  DFF \sreg_reg[1867]  ( .D(c[1868]), .CLK(clk), .RST(rst), .Q(sreg[1867]) );
  DFF \sreg_reg[1866]  ( .D(c[1867]), .CLK(clk), .RST(rst), .Q(sreg[1866]) );
  DFF \sreg_reg[1865]  ( .D(c[1866]), .CLK(clk), .RST(rst), .Q(sreg[1865]) );
  DFF \sreg_reg[1864]  ( .D(c[1865]), .CLK(clk), .RST(rst), .Q(sreg[1864]) );
  DFF \sreg_reg[1863]  ( .D(c[1864]), .CLK(clk), .RST(rst), .Q(sreg[1863]) );
  DFF \sreg_reg[1862]  ( .D(c[1863]), .CLK(clk), .RST(rst), .Q(sreg[1862]) );
  DFF \sreg_reg[1861]  ( .D(c[1862]), .CLK(clk), .RST(rst), .Q(sreg[1861]) );
  DFF \sreg_reg[1860]  ( .D(c[1861]), .CLK(clk), .RST(rst), .Q(sreg[1860]) );
  DFF \sreg_reg[1859]  ( .D(c[1860]), .CLK(clk), .RST(rst), .Q(sreg[1859]) );
  DFF \sreg_reg[1858]  ( .D(c[1859]), .CLK(clk), .RST(rst), .Q(sreg[1858]) );
  DFF \sreg_reg[1857]  ( .D(c[1858]), .CLK(clk), .RST(rst), .Q(sreg[1857]) );
  DFF \sreg_reg[1856]  ( .D(c[1857]), .CLK(clk), .RST(rst), .Q(sreg[1856]) );
  DFF \sreg_reg[1855]  ( .D(c[1856]), .CLK(clk), .RST(rst), .Q(sreg[1855]) );
  DFF \sreg_reg[1854]  ( .D(c[1855]), .CLK(clk), .RST(rst), .Q(sreg[1854]) );
  DFF \sreg_reg[1853]  ( .D(c[1854]), .CLK(clk), .RST(rst), .Q(sreg[1853]) );
  DFF \sreg_reg[1852]  ( .D(c[1853]), .CLK(clk), .RST(rst), .Q(sreg[1852]) );
  DFF \sreg_reg[1851]  ( .D(c[1852]), .CLK(clk), .RST(rst), .Q(sreg[1851]) );
  DFF \sreg_reg[1850]  ( .D(c[1851]), .CLK(clk), .RST(rst), .Q(sreg[1850]) );
  DFF \sreg_reg[1849]  ( .D(c[1850]), .CLK(clk), .RST(rst), .Q(sreg[1849]) );
  DFF \sreg_reg[1848]  ( .D(c[1849]), .CLK(clk), .RST(rst), .Q(sreg[1848]) );
  DFF \sreg_reg[1847]  ( .D(c[1848]), .CLK(clk), .RST(rst), .Q(sreg[1847]) );
  DFF \sreg_reg[1846]  ( .D(c[1847]), .CLK(clk), .RST(rst), .Q(sreg[1846]) );
  DFF \sreg_reg[1845]  ( .D(c[1846]), .CLK(clk), .RST(rst), .Q(sreg[1845]) );
  DFF \sreg_reg[1844]  ( .D(c[1845]), .CLK(clk), .RST(rst), .Q(sreg[1844]) );
  DFF \sreg_reg[1843]  ( .D(c[1844]), .CLK(clk), .RST(rst), .Q(sreg[1843]) );
  DFF \sreg_reg[1842]  ( .D(c[1843]), .CLK(clk), .RST(rst), .Q(sreg[1842]) );
  DFF \sreg_reg[1841]  ( .D(c[1842]), .CLK(clk), .RST(rst), .Q(sreg[1841]) );
  DFF \sreg_reg[1840]  ( .D(c[1841]), .CLK(clk), .RST(rst), .Q(sreg[1840]) );
  DFF \sreg_reg[1839]  ( .D(c[1840]), .CLK(clk), .RST(rst), .Q(sreg[1839]) );
  DFF \sreg_reg[1838]  ( .D(c[1839]), .CLK(clk), .RST(rst), .Q(sreg[1838]) );
  DFF \sreg_reg[1837]  ( .D(c[1838]), .CLK(clk), .RST(rst), .Q(sreg[1837]) );
  DFF \sreg_reg[1836]  ( .D(c[1837]), .CLK(clk), .RST(rst), .Q(sreg[1836]) );
  DFF \sreg_reg[1835]  ( .D(c[1836]), .CLK(clk), .RST(rst), .Q(sreg[1835]) );
  DFF \sreg_reg[1834]  ( .D(c[1835]), .CLK(clk), .RST(rst), .Q(sreg[1834]) );
  DFF \sreg_reg[1833]  ( .D(c[1834]), .CLK(clk), .RST(rst), .Q(sreg[1833]) );
  DFF \sreg_reg[1832]  ( .D(c[1833]), .CLK(clk), .RST(rst), .Q(sreg[1832]) );
  DFF \sreg_reg[1831]  ( .D(c[1832]), .CLK(clk), .RST(rst), .Q(sreg[1831]) );
  DFF \sreg_reg[1830]  ( .D(c[1831]), .CLK(clk), .RST(rst), .Q(sreg[1830]) );
  DFF \sreg_reg[1829]  ( .D(c[1830]), .CLK(clk), .RST(rst), .Q(sreg[1829]) );
  DFF \sreg_reg[1828]  ( .D(c[1829]), .CLK(clk), .RST(rst), .Q(sreg[1828]) );
  DFF \sreg_reg[1827]  ( .D(c[1828]), .CLK(clk), .RST(rst), .Q(sreg[1827]) );
  DFF \sreg_reg[1826]  ( .D(c[1827]), .CLK(clk), .RST(rst), .Q(sreg[1826]) );
  DFF \sreg_reg[1825]  ( .D(c[1826]), .CLK(clk), .RST(rst), .Q(sreg[1825]) );
  DFF \sreg_reg[1824]  ( .D(c[1825]), .CLK(clk), .RST(rst), .Q(sreg[1824]) );
  DFF \sreg_reg[1823]  ( .D(c[1824]), .CLK(clk), .RST(rst), .Q(sreg[1823]) );
  DFF \sreg_reg[1822]  ( .D(c[1823]), .CLK(clk), .RST(rst), .Q(sreg[1822]) );
  DFF \sreg_reg[1821]  ( .D(c[1822]), .CLK(clk), .RST(rst), .Q(sreg[1821]) );
  DFF \sreg_reg[1820]  ( .D(c[1821]), .CLK(clk), .RST(rst), .Q(sreg[1820]) );
  DFF \sreg_reg[1819]  ( .D(c[1820]), .CLK(clk), .RST(rst), .Q(sreg[1819]) );
  DFF \sreg_reg[1818]  ( .D(c[1819]), .CLK(clk), .RST(rst), .Q(sreg[1818]) );
  DFF \sreg_reg[1817]  ( .D(c[1818]), .CLK(clk), .RST(rst), .Q(sreg[1817]) );
  DFF \sreg_reg[1816]  ( .D(c[1817]), .CLK(clk), .RST(rst), .Q(sreg[1816]) );
  DFF \sreg_reg[1815]  ( .D(c[1816]), .CLK(clk), .RST(rst), .Q(sreg[1815]) );
  DFF \sreg_reg[1814]  ( .D(c[1815]), .CLK(clk), .RST(rst), .Q(sreg[1814]) );
  DFF \sreg_reg[1813]  ( .D(c[1814]), .CLK(clk), .RST(rst), .Q(sreg[1813]) );
  DFF \sreg_reg[1812]  ( .D(c[1813]), .CLK(clk), .RST(rst), .Q(sreg[1812]) );
  DFF \sreg_reg[1811]  ( .D(c[1812]), .CLK(clk), .RST(rst), .Q(sreg[1811]) );
  DFF \sreg_reg[1810]  ( .D(c[1811]), .CLK(clk), .RST(rst), .Q(sreg[1810]) );
  DFF \sreg_reg[1809]  ( .D(c[1810]), .CLK(clk), .RST(rst), .Q(sreg[1809]) );
  DFF \sreg_reg[1808]  ( .D(c[1809]), .CLK(clk), .RST(rst), .Q(sreg[1808]) );
  DFF \sreg_reg[1807]  ( .D(c[1808]), .CLK(clk), .RST(rst), .Q(sreg[1807]) );
  DFF \sreg_reg[1806]  ( .D(c[1807]), .CLK(clk), .RST(rst), .Q(sreg[1806]) );
  DFF \sreg_reg[1805]  ( .D(c[1806]), .CLK(clk), .RST(rst), .Q(sreg[1805]) );
  DFF \sreg_reg[1804]  ( .D(c[1805]), .CLK(clk), .RST(rst), .Q(sreg[1804]) );
  DFF \sreg_reg[1803]  ( .D(c[1804]), .CLK(clk), .RST(rst), .Q(sreg[1803]) );
  DFF \sreg_reg[1802]  ( .D(c[1803]), .CLK(clk), .RST(rst), .Q(sreg[1802]) );
  DFF \sreg_reg[1801]  ( .D(c[1802]), .CLK(clk), .RST(rst), .Q(sreg[1801]) );
  DFF \sreg_reg[1800]  ( .D(c[1801]), .CLK(clk), .RST(rst), .Q(sreg[1800]) );
  DFF \sreg_reg[1799]  ( .D(c[1800]), .CLK(clk), .RST(rst), .Q(sreg[1799]) );
  DFF \sreg_reg[1798]  ( .D(c[1799]), .CLK(clk), .RST(rst), .Q(sreg[1798]) );
  DFF \sreg_reg[1797]  ( .D(c[1798]), .CLK(clk), .RST(rst), .Q(sreg[1797]) );
  DFF \sreg_reg[1796]  ( .D(c[1797]), .CLK(clk), .RST(rst), .Q(sreg[1796]) );
  DFF \sreg_reg[1795]  ( .D(c[1796]), .CLK(clk), .RST(rst), .Q(sreg[1795]) );
  DFF \sreg_reg[1794]  ( .D(c[1795]), .CLK(clk), .RST(rst), .Q(sreg[1794]) );
  DFF \sreg_reg[1793]  ( .D(c[1794]), .CLK(clk), .RST(rst), .Q(sreg[1793]) );
  DFF \sreg_reg[1792]  ( .D(c[1793]), .CLK(clk), .RST(rst), .Q(sreg[1792]) );
  DFF \sreg_reg[1791]  ( .D(c[1792]), .CLK(clk), .RST(rst), .Q(sreg[1791]) );
  DFF \sreg_reg[1790]  ( .D(c[1791]), .CLK(clk), .RST(rst), .Q(sreg[1790]) );
  DFF \sreg_reg[1789]  ( .D(c[1790]), .CLK(clk), .RST(rst), .Q(sreg[1789]) );
  DFF \sreg_reg[1788]  ( .D(c[1789]), .CLK(clk), .RST(rst), .Q(sreg[1788]) );
  DFF \sreg_reg[1787]  ( .D(c[1788]), .CLK(clk), .RST(rst), .Q(sreg[1787]) );
  DFF \sreg_reg[1786]  ( .D(c[1787]), .CLK(clk), .RST(rst), .Q(sreg[1786]) );
  DFF \sreg_reg[1785]  ( .D(c[1786]), .CLK(clk), .RST(rst), .Q(sreg[1785]) );
  DFF \sreg_reg[1784]  ( .D(c[1785]), .CLK(clk), .RST(rst), .Q(sreg[1784]) );
  DFF \sreg_reg[1783]  ( .D(c[1784]), .CLK(clk), .RST(rst), .Q(sreg[1783]) );
  DFF \sreg_reg[1782]  ( .D(c[1783]), .CLK(clk), .RST(rst), .Q(sreg[1782]) );
  DFF \sreg_reg[1781]  ( .D(c[1782]), .CLK(clk), .RST(rst), .Q(sreg[1781]) );
  DFF \sreg_reg[1780]  ( .D(c[1781]), .CLK(clk), .RST(rst), .Q(sreg[1780]) );
  DFF \sreg_reg[1779]  ( .D(c[1780]), .CLK(clk), .RST(rst), .Q(sreg[1779]) );
  DFF \sreg_reg[1778]  ( .D(c[1779]), .CLK(clk), .RST(rst), .Q(sreg[1778]) );
  DFF \sreg_reg[1777]  ( .D(c[1778]), .CLK(clk), .RST(rst), .Q(sreg[1777]) );
  DFF \sreg_reg[1776]  ( .D(c[1777]), .CLK(clk), .RST(rst), .Q(sreg[1776]) );
  DFF \sreg_reg[1775]  ( .D(c[1776]), .CLK(clk), .RST(rst), .Q(sreg[1775]) );
  DFF \sreg_reg[1774]  ( .D(c[1775]), .CLK(clk), .RST(rst), .Q(sreg[1774]) );
  DFF \sreg_reg[1773]  ( .D(c[1774]), .CLK(clk), .RST(rst), .Q(sreg[1773]) );
  DFF \sreg_reg[1772]  ( .D(c[1773]), .CLK(clk), .RST(rst), .Q(sreg[1772]) );
  DFF \sreg_reg[1771]  ( .D(c[1772]), .CLK(clk), .RST(rst), .Q(sreg[1771]) );
  DFF \sreg_reg[1770]  ( .D(c[1771]), .CLK(clk), .RST(rst), .Q(sreg[1770]) );
  DFF \sreg_reg[1769]  ( .D(c[1770]), .CLK(clk), .RST(rst), .Q(sreg[1769]) );
  DFF \sreg_reg[1768]  ( .D(c[1769]), .CLK(clk), .RST(rst), .Q(sreg[1768]) );
  DFF \sreg_reg[1767]  ( .D(c[1768]), .CLK(clk), .RST(rst), .Q(sreg[1767]) );
  DFF \sreg_reg[1766]  ( .D(c[1767]), .CLK(clk), .RST(rst), .Q(sreg[1766]) );
  DFF \sreg_reg[1765]  ( .D(c[1766]), .CLK(clk), .RST(rst), .Q(sreg[1765]) );
  DFF \sreg_reg[1764]  ( .D(c[1765]), .CLK(clk), .RST(rst), .Q(sreg[1764]) );
  DFF \sreg_reg[1763]  ( .D(c[1764]), .CLK(clk), .RST(rst), .Q(sreg[1763]) );
  DFF \sreg_reg[1762]  ( .D(c[1763]), .CLK(clk), .RST(rst), .Q(sreg[1762]) );
  DFF \sreg_reg[1761]  ( .D(c[1762]), .CLK(clk), .RST(rst), .Q(sreg[1761]) );
  DFF \sreg_reg[1760]  ( .D(c[1761]), .CLK(clk), .RST(rst), .Q(sreg[1760]) );
  DFF \sreg_reg[1759]  ( .D(c[1760]), .CLK(clk), .RST(rst), .Q(sreg[1759]) );
  DFF \sreg_reg[1758]  ( .D(c[1759]), .CLK(clk), .RST(rst), .Q(sreg[1758]) );
  DFF \sreg_reg[1757]  ( .D(c[1758]), .CLK(clk), .RST(rst), .Q(sreg[1757]) );
  DFF \sreg_reg[1756]  ( .D(c[1757]), .CLK(clk), .RST(rst), .Q(sreg[1756]) );
  DFF \sreg_reg[1755]  ( .D(c[1756]), .CLK(clk), .RST(rst), .Q(sreg[1755]) );
  DFF \sreg_reg[1754]  ( .D(c[1755]), .CLK(clk), .RST(rst), .Q(sreg[1754]) );
  DFF \sreg_reg[1753]  ( .D(c[1754]), .CLK(clk), .RST(rst), .Q(sreg[1753]) );
  DFF \sreg_reg[1752]  ( .D(c[1753]), .CLK(clk), .RST(rst), .Q(sreg[1752]) );
  DFF \sreg_reg[1751]  ( .D(c[1752]), .CLK(clk), .RST(rst), .Q(sreg[1751]) );
  DFF \sreg_reg[1750]  ( .D(c[1751]), .CLK(clk), .RST(rst), .Q(sreg[1750]) );
  DFF \sreg_reg[1749]  ( .D(c[1750]), .CLK(clk), .RST(rst), .Q(sreg[1749]) );
  DFF \sreg_reg[1748]  ( .D(c[1749]), .CLK(clk), .RST(rst), .Q(sreg[1748]) );
  DFF \sreg_reg[1747]  ( .D(c[1748]), .CLK(clk), .RST(rst), .Q(sreg[1747]) );
  DFF \sreg_reg[1746]  ( .D(c[1747]), .CLK(clk), .RST(rst), .Q(sreg[1746]) );
  DFF \sreg_reg[1745]  ( .D(c[1746]), .CLK(clk), .RST(rst), .Q(sreg[1745]) );
  DFF \sreg_reg[1744]  ( .D(c[1745]), .CLK(clk), .RST(rst), .Q(sreg[1744]) );
  DFF \sreg_reg[1743]  ( .D(c[1744]), .CLK(clk), .RST(rst), .Q(sreg[1743]) );
  DFF \sreg_reg[1742]  ( .D(c[1743]), .CLK(clk), .RST(rst), .Q(sreg[1742]) );
  DFF \sreg_reg[1741]  ( .D(c[1742]), .CLK(clk), .RST(rst), .Q(sreg[1741]) );
  DFF \sreg_reg[1740]  ( .D(c[1741]), .CLK(clk), .RST(rst), .Q(sreg[1740]) );
  DFF \sreg_reg[1739]  ( .D(c[1740]), .CLK(clk), .RST(rst), .Q(sreg[1739]) );
  DFF \sreg_reg[1738]  ( .D(c[1739]), .CLK(clk), .RST(rst), .Q(sreg[1738]) );
  DFF \sreg_reg[1737]  ( .D(c[1738]), .CLK(clk), .RST(rst), .Q(sreg[1737]) );
  DFF \sreg_reg[1736]  ( .D(c[1737]), .CLK(clk), .RST(rst), .Q(sreg[1736]) );
  DFF \sreg_reg[1735]  ( .D(c[1736]), .CLK(clk), .RST(rst), .Q(sreg[1735]) );
  DFF \sreg_reg[1734]  ( .D(c[1735]), .CLK(clk), .RST(rst), .Q(sreg[1734]) );
  DFF \sreg_reg[1733]  ( .D(c[1734]), .CLK(clk), .RST(rst), .Q(sreg[1733]) );
  DFF \sreg_reg[1732]  ( .D(c[1733]), .CLK(clk), .RST(rst), .Q(sreg[1732]) );
  DFF \sreg_reg[1731]  ( .D(c[1732]), .CLK(clk), .RST(rst), .Q(sreg[1731]) );
  DFF \sreg_reg[1730]  ( .D(c[1731]), .CLK(clk), .RST(rst), .Q(sreg[1730]) );
  DFF \sreg_reg[1729]  ( .D(c[1730]), .CLK(clk), .RST(rst), .Q(sreg[1729]) );
  DFF \sreg_reg[1728]  ( .D(c[1729]), .CLK(clk), .RST(rst), .Q(sreg[1728]) );
  DFF \sreg_reg[1727]  ( .D(c[1728]), .CLK(clk), .RST(rst), .Q(sreg[1727]) );
  DFF \sreg_reg[1726]  ( .D(c[1727]), .CLK(clk), .RST(rst), .Q(sreg[1726]) );
  DFF \sreg_reg[1725]  ( .D(c[1726]), .CLK(clk), .RST(rst), .Q(sreg[1725]) );
  DFF \sreg_reg[1724]  ( .D(c[1725]), .CLK(clk), .RST(rst), .Q(sreg[1724]) );
  DFF \sreg_reg[1723]  ( .D(c[1724]), .CLK(clk), .RST(rst), .Q(sreg[1723]) );
  DFF \sreg_reg[1722]  ( .D(c[1723]), .CLK(clk), .RST(rst), .Q(sreg[1722]) );
  DFF \sreg_reg[1721]  ( .D(c[1722]), .CLK(clk), .RST(rst), .Q(sreg[1721]) );
  DFF \sreg_reg[1720]  ( .D(c[1721]), .CLK(clk), .RST(rst), .Q(sreg[1720]) );
  DFF \sreg_reg[1719]  ( .D(c[1720]), .CLK(clk), .RST(rst), .Q(sreg[1719]) );
  DFF \sreg_reg[1718]  ( .D(c[1719]), .CLK(clk), .RST(rst), .Q(sreg[1718]) );
  DFF \sreg_reg[1717]  ( .D(c[1718]), .CLK(clk), .RST(rst), .Q(sreg[1717]) );
  DFF \sreg_reg[1716]  ( .D(c[1717]), .CLK(clk), .RST(rst), .Q(sreg[1716]) );
  DFF \sreg_reg[1715]  ( .D(c[1716]), .CLK(clk), .RST(rst), .Q(sreg[1715]) );
  DFF \sreg_reg[1714]  ( .D(c[1715]), .CLK(clk), .RST(rst), .Q(sreg[1714]) );
  DFF \sreg_reg[1713]  ( .D(c[1714]), .CLK(clk), .RST(rst), .Q(sreg[1713]) );
  DFF \sreg_reg[1712]  ( .D(c[1713]), .CLK(clk), .RST(rst), .Q(sreg[1712]) );
  DFF \sreg_reg[1711]  ( .D(c[1712]), .CLK(clk), .RST(rst), .Q(sreg[1711]) );
  DFF \sreg_reg[1710]  ( .D(c[1711]), .CLK(clk), .RST(rst), .Q(sreg[1710]) );
  DFF \sreg_reg[1709]  ( .D(c[1710]), .CLK(clk), .RST(rst), .Q(sreg[1709]) );
  DFF \sreg_reg[1708]  ( .D(c[1709]), .CLK(clk), .RST(rst), .Q(sreg[1708]) );
  DFF \sreg_reg[1707]  ( .D(c[1708]), .CLK(clk), .RST(rst), .Q(sreg[1707]) );
  DFF \sreg_reg[1706]  ( .D(c[1707]), .CLK(clk), .RST(rst), .Q(sreg[1706]) );
  DFF \sreg_reg[1705]  ( .D(c[1706]), .CLK(clk), .RST(rst), .Q(sreg[1705]) );
  DFF \sreg_reg[1704]  ( .D(c[1705]), .CLK(clk), .RST(rst), .Q(sreg[1704]) );
  DFF \sreg_reg[1703]  ( .D(c[1704]), .CLK(clk), .RST(rst), .Q(sreg[1703]) );
  DFF \sreg_reg[1702]  ( .D(c[1703]), .CLK(clk), .RST(rst), .Q(sreg[1702]) );
  DFF \sreg_reg[1701]  ( .D(c[1702]), .CLK(clk), .RST(rst), .Q(sreg[1701]) );
  DFF \sreg_reg[1700]  ( .D(c[1701]), .CLK(clk), .RST(rst), .Q(sreg[1700]) );
  DFF \sreg_reg[1699]  ( .D(c[1700]), .CLK(clk), .RST(rst), .Q(sreg[1699]) );
  DFF \sreg_reg[1698]  ( .D(c[1699]), .CLK(clk), .RST(rst), .Q(sreg[1698]) );
  DFF \sreg_reg[1697]  ( .D(c[1698]), .CLK(clk), .RST(rst), .Q(sreg[1697]) );
  DFF \sreg_reg[1696]  ( .D(c[1697]), .CLK(clk), .RST(rst), .Q(sreg[1696]) );
  DFF \sreg_reg[1695]  ( .D(c[1696]), .CLK(clk), .RST(rst), .Q(sreg[1695]) );
  DFF \sreg_reg[1694]  ( .D(c[1695]), .CLK(clk), .RST(rst), .Q(sreg[1694]) );
  DFF \sreg_reg[1693]  ( .D(c[1694]), .CLK(clk), .RST(rst), .Q(sreg[1693]) );
  DFF \sreg_reg[1692]  ( .D(c[1693]), .CLK(clk), .RST(rst), .Q(sreg[1692]) );
  DFF \sreg_reg[1691]  ( .D(c[1692]), .CLK(clk), .RST(rst), .Q(sreg[1691]) );
  DFF \sreg_reg[1690]  ( .D(c[1691]), .CLK(clk), .RST(rst), .Q(sreg[1690]) );
  DFF \sreg_reg[1689]  ( .D(c[1690]), .CLK(clk), .RST(rst), .Q(sreg[1689]) );
  DFF \sreg_reg[1688]  ( .D(c[1689]), .CLK(clk), .RST(rst), .Q(sreg[1688]) );
  DFF \sreg_reg[1687]  ( .D(c[1688]), .CLK(clk), .RST(rst), .Q(sreg[1687]) );
  DFF \sreg_reg[1686]  ( .D(c[1687]), .CLK(clk), .RST(rst), .Q(sreg[1686]) );
  DFF \sreg_reg[1685]  ( .D(c[1686]), .CLK(clk), .RST(rst), .Q(sreg[1685]) );
  DFF \sreg_reg[1684]  ( .D(c[1685]), .CLK(clk), .RST(rst), .Q(sreg[1684]) );
  DFF \sreg_reg[1683]  ( .D(c[1684]), .CLK(clk), .RST(rst), .Q(sreg[1683]) );
  DFF \sreg_reg[1682]  ( .D(c[1683]), .CLK(clk), .RST(rst), .Q(sreg[1682]) );
  DFF \sreg_reg[1681]  ( .D(c[1682]), .CLK(clk), .RST(rst), .Q(sreg[1681]) );
  DFF \sreg_reg[1680]  ( .D(c[1681]), .CLK(clk), .RST(rst), .Q(sreg[1680]) );
  DFF \sreg_reg[1679]  ( .D(c[1680]), .CLK(clk), .RST(rst), .Q(sreg[1679]) );
  DFF \sreg_reg[1678]  ( .D(c[1679]), .CLK(clk), .RST(rst), .Q(sreg[1678]) );
  DFF \sreg_reg[1677]  ( .D(c[1678]), .CLK(clk), .RST(rst), .Q(sreg[1677]) );
  DFF \sreg_reg[1676]  ( .D(c[1677]), .CLK(clk), .RST(rst), .Q(sreg[1676]) );
  DFF \sreg_reg[1675]  ( .D(c[1676]), .CLK(clk), .RST(rst), .Q(sreg[1675]) );
  DFF \sreg_reg[1674]  ( .D(c[1675]), .CLK(clk), .RST(rst), .Q(sreg[1674]) );
  DFF \sreg_reg[1673]  ( .D(c[1674]), .CLK(clk), .RST(rst), .Q(sreg[1673]) );
  DFF \sreg_reg[1672]  ( .D(c[1673]), .CLK(clk), .RST(rst), .Q(sreg[1672]) );
  DFF \sreg_reg[1671]  ( .D(c[1672]), .CLK(clk), .RST(rst), .Q(sreg[1671]) );
  DFF \sreg_reg[1670]  ( .D(c[1671]), .CLK(clk), .RST(rst), .Q(sreg[1670]) );
  DFF \sreg_reg[1669]  ( .D(c[1670]), .CLK(clk), .RST(rst), .Q(sreg[1669]) );
  DFF \sreg_reg[1668]  ( .D(c[1669]), .CLK(clk), .RST(rst), .Q(sreg[1668]) );
  DFF \sreg_reg[1667]  ( .D(c[1668]), .CLK(clk), .RST(rst), .Q(sreg[1667]) );
  DFF \sreg_reg[1666]  ( .D(c[1667]), .CLK(clk), .RST(rst), .Q(sreg[1666]) );
  DFF \sreg_reg[1665]  ( .D(c[1666]), .CLK(clk), .RST(rst), .Q(sreg[1665]) );
  DFF \sreg_reg[1664]  ( .D(c[1665]), .CLK(clk), .RST(rst), .Q(sreg[1664]) );
  DFF \sreg_reg[1663]  ( .D(c[1664]), .CLK(clk), .RST(rst), .Q(sreg[1663]) );
  DFF \sreg_reg[1662]  ( .D(c[1663]), .CLK(clk), .RST(rst), .Q(sreg[1662]) );
  DFF \sreg_reg[1661]  ( .D(c[1662]), .CLK(clk), .RST(rst), .Q(sreg[1661]) );
  DFF \sreg_reg[1660]  ( .D(c[1661]), .CLK(clk), .RST(rst), .Q(sreg[1660]) );
  DFF \sreg_reg[1659]  ( .D(c[1660]), .CLK(clk), .RST(rst), .Q(sreg[1659]) );
  DFF \sreg_reg[1658]  ( .D(c[1659]), .CLK(clk), .RST(rst), .Q(sreg[1658]) );
  DFF \sreg_reg[1657]  ( .D(c[1658]), .CLK(clk), .RST(rst), .Q(sreg[1657]) );
  DFF \sreg_reg[1656]  ( .D(c[1657]), .CLK(clk), .RST(rst), .Q(sreg[1656]) );
  DFF \sreg_reg[1655]  ( .D(c[1656]), .CLK(clk), .RST(rst), .Q(sreg[1655]) );
  DFF \sreg_reg[1654]  ( .D(c[1655]), .CLK(clk), .RST(rst), .Q(sreg[1654]) );
  DFF \sreg_reg[1653]  ( .D(c[1654]), .CLK(clk), .RST(rst), .Q(sreg[1653]) );
  DFF \sreg_reg[1652]  ( .D(c[1653]), .CLK(clk), .RST(rst), .Q(sreg[1652]) );
  DFF \sreg_reg[1651]  ( .D(c[1652]), .CLK(clk), .RST(rst), .Q(sreg[1651]) );
  DFF \sreg_reg[1650]  ( .D(c[1651]), .CLK(clk), .RST(rst), .Q(sreg[1650]) );
  DFF \sreg_reg[1649]  ( .D(c[1650]), .CLK(clk), .RST(rst), .Q(sreg[1649]) );
  DFF \sreg_reg[1648]  ( .D(c[1649]), .CLK(clk), .RST(rst), .Q(sreg[1648]) );
  DFF \sreg_reg[1647]  ( .D(c[1648]), .CLK(clk), .RST(rst), .Q(sreg[1647]) );
  DFF \sreg_reg[1646]  ( .D(c[1647]), .CLK(clk), .RST(rst), .Q(sreg[1646]) );
  DFF \sreg_reg[1645]  ( .D(c[1646]), .CLK(clk), .RST(rst), .Q(sreg[1645]) );
  DFF \sreg_reg[1644]  ( .D(c[1645]), .CLK(clk), .RST(rst), .Q(sreg[1644]) );
  DFF \sreg_reg[1643]  ( .D(c[1644]), .CLK(clk), .RST(rst), .Q(sreg[1643]) );
  DFF \sreg_reg[1642]  ( .D(c[1643]), .CLK(clk), .RST(rst), .Q(sreg[1642]) );
  DFF \sreg_reg[1641]  ( .D(c[1642]), .CLK(clk), .RST(rst), .Q(sreg[1641]) );
  DFF \sreg_reg[1640]  ( .D(c[1641]), .CLK(clk), .RST(rst), .Q(sreg[1640]) );
  DFF \sreg_reg[1639]  ( .D(c[1640]), .CLK(clk), .RST(rst), .Q(sreg[1639]) );
  DFF \sreg_reg[1638]  ( .D(c[1639]), .CLK(clk), .RST(rst), .Q(sreg[1638]) );
  DFF \sreg_reg[1637]  ( .D(c[1638]), .CLK(clk), .RST(rst), .Q(sreg[1637]) );
  DFF \sreg_reg[1636]  ( .D(c[1637]), .CLK(clk), .RST(rst), .Q(sreg[1636]) );
  DFF \sreg_reg[1635]  ( .D(c[1636]), .CLK(clk), .RST(rst), .Q(sreg[1635]) );
  DFF \sreg_reg[1634]  ( .D(c[1635]), .CLK(clk), .RST(rst), .Q(sreg[1634]) );
  DFF \sreg_reg[1633]  ( .D(c[1634]), .CLK(clk), .RST(rst), .Q(sreg[1633]) );
  DFF \sreg_reg[1632]  ( .D(c[1633]), .CLK(clk), .RST(rst), .Q(sreg[1632]) );
  DFF \sreg_reg[1631]  ( .D(c[1632]), .CLK(clk), .RST(rst), .Q(sreg[1631]) );
  DFF \sreg_reg[1630]  ( .D(c[1631]), .CLK(clk), .RST(rst), .Q(sreg[1630]) );
  DFF \sreg_reg[1629]  ( .D(c[1630]), .CLK(clk), .RST(rst), .Q(sreg[1629]) );
  DFF \sreg_reg[1628]  ( .D(c[1629]), .CLK(clk), .RST(rst), .Q(sreg[1628]) );
  DFF \sreg_reg[1627]  ( .D(c[1628]), .CLK(clk), .RST(rst), .Q(sreg[1627]) );
  DFF \sreg_reg[1626]  ( .D(c[1627]), .CLK(clk), .RST(rst), .Q(sreg[1626]) );
  DFF \sreg_reg[1625]  ( .D(c[1626]), .CLK(clk), .RST(rst), .Q(sreg[1625]) );
  DFF \sreg_reg[1624]  ( .D(c[1625]), .CLK(clk), .RST(rst), .Q(sreg[1624]) );
  DFF \sreg_reg[1623]  ( .D(c[1624]), .CLK(clk), .RST(rst), .Q(sreg[1623]) );
  DFF \sreg_reg[1622]  ( .D(c[1623]), .CLK(clk), .RST(rst), .Q(sreg[1622]) );
  DFF \sreg_reg[1621]  ( .D(c[1622]), .CLK(clk), .RST(rst), .Q(sreg[1621]) );
  DFF \sreg_reg[1620]  ( .D(c[1621]), .CLK(clk), .RST(rst), .Q(sreg[1620]) );
  DFF \sreg_reg[1619]  ( .D(c[1620]), .CLK(clk), .RST(rst), .Q(sreg[1619]) );
  DFF \sreg_reg[1618]  ( .D(c[1619]), .CLK(clk), .RST(rst), .Q(sreg[1618]) );
  DFF \sreg_reg[1617]  ( .D(c[1618]), .CLK(clk), .RST(rst), .Q(sreg[1617]) );
  DFF \sreg_reg[1616]  ( .D(c[1617]), .CLK(clk), .RST(rst), .Q(sreg[1616]) );
  DFF \sreg_reg[1615]  ( .D(c[1616]), .CLK(clk), .RST(rst), .Q(sreg[1615]) );
  DFF \sreg_reg[1614]  ( .D(c[1615]), .CLK(clk), .RST(rst), .Q(sreg[1614]) );
  DFF \sreg_reg[1613]  ( .D(c[1614]), .CLK(clk), .RST(rst), .Q(sreg[1613]) );
  DFF \sreg_reg[1612]  ( .D(c[1613]), .CLK(clk), .RST(rst), .Q(sreg[1612]) );
  DFF \sreg_reg[1611]  ( .D(c[1612]), .CLK(clk), .RST(rst), .Q(sreg[1611]) );
  DFF \sreg_reg[1610]  ( .D(c[1611]), .CLK(clk), .RST(rst), .Q(sreg[1610]) );
  DFF \sreg_reg[1609]  ( .D(c[1610]), .CLK(clk), .RST(rst), .Q(sreg[1609]) );
  DFF \sreg_reg[1608]  ( .D(c[1609]), .CLK(clk), .RST(rst), .Q(sreg[1608]) );
  DFF \sreg_reg[1607]  ( .D(c[1608]), .CLK(clk), .RST(rst), .Q(sreg[1607]) );
  DFF \sreg_reg[1606]  ( .D(c[1607]), .CLK(clk), .RST(rst), .Q(sreg[1606]) );
  DFF \sreg_reg[1605]  ( .D(c[1606]), .CLK(clk), .RST(rst), .Q(sreg[1605]) );
  DFF \sreg_reg[1604]  ( .D(c[1605]), .CLK(clk), .RST(rst), .Q(sreg[1604]) );
  DFF \sreg_reg[1603]  ( .D(c[1604]), .CLK(clk), .RST(rst), .Q(sreg[1603]) );
  DFF \sreg_reg[1602]  ( .D(c[1603]), .CLK(clk), .RST(rst), .Q(sreg[1602]) );
  DFF \sreg_reg[1601]  ( .D(c[1602]), .CLK(clk), .RST(rst), .Q(sreg[1601]) );
  DFF \sreg_reg[1600]  ( .D(c[1601]), .CLK(clk), .RST(rst), .Q(sreg[1600]) );
  DFF \sreg_reg[1599]  ( .D(c[1600]), .CLK(clk), .RST(rst), .Q(sreg[1599]) );
  DFF \sreg_reg[1598]  ( .D(c[1599]), .CLK(clk), .RST(rst), .Q(sreg[1598]) );
  DFF \sreg_reg[1597]  ( .D(c[1598]), .CLK(clk), .RST(rst), .Q(sreg[1597]) );
  DFF \sreg_reg[1596]  ( .D(c[1597]), .CLK(clk), .RST(rst), .Q(sreg[1596]) );
  DFF \sreg_reg[1595]  ( .D(c[1596]), .CLK(clk), .RST(rst), .Q(sreg[1595]) );
  DFF \sreg_reg[1594]  ( .D(c[1595]), .CLK(clk), .RST(rst), .Q(sreg[1594]) );
  DFF \sreg_reg[1593]  ( .D(c[1594]), .CLK(clk), .RST(rst), .Q(sreg[1593]) );
  DFF \sreg_reg[1592]  ( .D(c[1593]), .CLK(clk), .RST(rst), .Q(sreg[1592]) );
  DFF \sreg_reg[1591]  ( .D(c[1592]), .CLK(clk), .RST(rst), .Q(sreg[1591]) );
  DFF \sreg_reg[1590]  ( .D(c[1591]), .CLK(clk), .RST(rst), .Q(sreg[1590]) );
  DFF \sreg_reg[1589]  ( .D(c[1590]), .CLK(clk), .RST(rst), .Q(sreg[1589]) );
  DFF \sreg_reg[1588]  ( .D(c[1589]), .CLK(clk), .RST(rst), .Q(sreg[1588]) );
  DFF \sreg_reg[1587]  ( .D(c[1588]), .CLK(clk), .RST(rst), .Q(sreg[1587]) );
  DFF \sreg_reg[1586]  ( .D(c[1587]), .CLK(clk), .RST(rst), .Q(sreg[1586]) );
  DFF \sreg_reg[1585]  ( .D(c[1586]), .CLK(clk), .RST(rst), .Q(sreg[1585]) );
  DFF \sreg_reg[1584]  ( .D(c[1585]), .CLK(clk), .RST(rst), .Q(sreg[1584]) );
  DFF \sreg_reg[1583]  ( .D(c[1584]), .CLK(clk), .RST(rst), .Q(sreg[1583]) );
  DFF \sreg_reg[1582]  ( .D(c[1583]), .CLK(clk), .RST(rst), .Q(sreg[1582]) );
  DFF \sreg_reg[1581]  ( .D(c[1582]), .CLK(clk), .RST(rst), .Q(sreg[1581]) );
  DFF \sreg_reg[1580]  ( .D(c[1581]), .CLK(clk), .RST(rst), .Q(sreg[1580]) );
  DFF \sreg_reg[1579]  ( .D(c[1580]), .CLK(clk), .RST(rst), .Q(sreg[1579]) );
  DFF \sreg_reg[1578]  ( .D(c[1579]), .CLK(clk), .RST(rst), .Q(sreg[1578]) );
  DFF \sreg_reg[1577]  ( .D(c[1578]), .CLK(clk), .RST(rst), .Q(sreg[1577]) );
  DFF \sreg_reg[1576]  ( .D(c[1577]), .CLK(clk), .RST(rst), .Q(sreg[1576]) );
  DFF \sreg_reg[1575]  ( .D(c[1576]), .CLK(clk), .RST(rst), .Q(sreg[1575]) );
  DFF \sreg_reg[1574]  ( .D(c[1575]), .CLK(clk), .RST(rst), .Q(sreg[1574]) );
  DFF \sreg_reg[1573]  ( .D(c[1574]), .CLK(clk), .RST(rst), .Q(sreg[1573]) );
  DFF \sreg_reg[1572]  ( .D(c[1573]), .CLK(clk), .RST(rst), .Q(sreg[1572]) );
  DFF \sreg_reg[1571]  ( .D(c[1572]), .CLK(clk), .RST(rst), .Q(sreg[1571]) );
  DFF \sreg_reg[1570]  ( .D(c[1571]), .CLK(clk), .RST(rst), .Q(sreg[1570]) );
  DFF \sreg_reg[1569]  ( .D(c[1570]), .CLK(clk), .RST(rst), .Q(sreg[1569]) );
  DFF \sreg_reg[1568]  ( .D(c[1569]), .CLK(clk), .RST(rst), .Q(sreg[1568]) );
  DFF \sreg_reg[1567]  ( .D(c[1568]), .CLK(clk), .RST(rst), .Q(sreg[1567]) );
  DFF \sreg_reg[1566]  ( .D(c[1567]), .CLK(clk), .RST(rst), .Q(sreg[1566]) );
  DFF \sreg_reg[1565]  ( .D(c[1566]), .CLK(clk), .RST(rst), .Q(sreg[1565]) );
  DFF \sreg_reg[1564]  ( .D(c[1565]), .CLK(clk), .RST(rst), .Q(sreg[1564]) );
  DFF \sreg_reg[1563]  ( .D(c[1564]), .CLK(clk), .RST(rst), .Q(sreg[1563]) );
  DFF \sreg_reg[1562]  ( .D(c[1563]), .CLK(clk), .RST(rst), .Q(sreg[1562]) );
  DFF \sreg_reg[1561]  ( .D(c[1562]), .CLK(clk), .RST(rst), .Q(sreg[1561]) );
  DFF \sreg_reg[1560]  ( .D(c[1561]), .CLK(clk), .RST(rst), .Q(sreg[1560]) );
  DFF \sreg_reg[1559]  ( .D(c[1560]), .CLK(clk), .RST(rst), .Q(sreg[1559]) );
  DFF \sreg_reg[1558]  ( .D(c[1559]), .CLK(clk), .RST(rst), .Q(sreg[1558]) );
  DFF \sreg_reg[1557]  ( .D(c[1558]), .CLK(clk), .RST(rst), .Q(sreg[1557]) );
  DFF \sreg_reg[1556]  ( .D(c[1557]), .CLK(clk), .RST(rst), .Q(sreg[1556]) );
  DFF \sreg_reg[1555]  ( .D(c[1556]), .CLK(clk), .RST(rst), .Q(sreg[1555]) );
  DFF \sreg_reg[1554]  ( .D(c[1555]), .CLK(clk), .RST(rst), .Q(sreg[1554]) );
  DFF \sreg_reg[1553]  ( .D(c[1554]), .CLK(clk), .RST(rst), .Q(sreg[1553]) );
  DFF \sreg_reg[1552]  ( .D(c[1553]), .CLK(clk), .RST(rst), .Q(sreg[1552]) );
  DFF \sreg_reg[1551]  ( .D(c[1552]), .CLK(clk), .RST(rst), .Q(sreg[1551]) );
  DFF \sreg_reg[1550]  ( .D(c[1551]), .CLK(clk), .RST(rst), .Q(sreg[1550]) );
  DFF \sreg_reg[1549]  ( .D(c[1550]), .CLK(clk), .RST(rst), .Q(sreg[1549]) );
  DFF \sreg_reg[1548]  ( .D(c[1549]), .CLK(clk), .RST(rst), .Q(sreg[1548]) );
  DFF \sreg_reg[1547]  ( .D(c[1548]), .CLK(clk), .RST(rst), .Q(sreg[1547]) );
  DFF \sreg_reg[1546]  ( .D(c[1547]), .CLK(clk), .RST(rst), .Q(sreg[1546]) );
  DFF \sreg_reg[1545]  ( .D(c[1546]), .CLK(clk), .RST(rst), .Q(sreg[1545]) );
  DFF \sreg_reg[1544]  ( .D(c[1545]), .CLK(clk), .RST(rst), .Q(sreg[1544]) );
  DFF \sreg_reg[1543]  ( .D(c[1544]), .CLK(clk), .RST(rst), .Q(sreg[1543]) );
  DFF \sreg_reg[1542]  ( .D(c[1543]), .CLK(clk), .RST(rst), .Q(sreg[1542]) );
  DFF \sreg_reg[1541]  ( .D(c[1542]), .CLK(clk), .RST(rst), .Q(sreg[1541]) );
  DFF \sreg_reg[1540]  ( .D(c[1541]), .CLK(clk), .RST(rst), .Q(sreg[1540]) );
  DFF \sreg_reg[1539]  ( .D(c[1540]), .CLK(clk), .RST(rst), .Q(sreg[1539]) );
  DFF \sreg_reg[1538]  ( .D(c[1539]), .CLK(clk), .RST(rst), .Q(sreg[1538]) );
  DFF \sreg_reg[1537]  ( .D(c[1538]), .CLK(clk), .RST(rst), .Q(sreg[1537]) );
  DFF \sreg_reg[1536]  ( .D(c[1537]), .CLK(clk), .RST(rst), .Q(sreg[1536]) );
  DFF \sreg_reg[1535]  ( .D(c[1536]), .CLK(clk), .RST(rst), .Q(sreg[1535]) );
  DFF \sreg_reg[1534]  ( .D(c[1535]), .CLK(clk), .RST(rst), .Q(sreg[1534]) );
  DFF \sreg_reg[1533]  ( .D(c[1534]), .CLK(clk), .RST(rst), .Q(sreg[1533]) );
  DFF \sreg_reg[1532]  ( .D(c[1533]), .CLK(clk), .RST(rst), .Q(sreg[1532]) );
  DFF \sreg_reg[1531]  ( .D(c[1532]), .CLK(clk), .RST(rst), .Q(sreg[1531]) );
  DFF \sreg_reg[1530]  ( .D(c[1531]), .CLK(clk), .RST(rst), .Q(sreg[1530]) );
  DFF \sreg_reg[1529]  ( .D(c[1530]), .CLK(clk), .RST(rst), .Q(sreg[1529]) );
  DFF \sreg_reg[1528]  ( .D(c[1529]), .CLK(clk), .RST(rst), .Q(sreg[1528]) );
  DFF \sreg_reg[1527]  ( .D(c[1528]), .CLK(clk), .RST(rst), .Q(sreg[1527]) );
  DFF \sreg_reg[1526]  ( .D(c[1527]), .CLK(clk), .RST(rst), .Q(sreg[1526]) );
  DFF \sreg_reg[1525]  ( .D(c[1526]), .CLK(clk), .RST(rst), .Q(sreg[1525]) );
  DFF \sreg_reg[1524]  ( .D(c[1525]), .CLK(clk), .RST(rst), .Q(sreg[1524]) );
  DFF \sreg_reg[1523]  ( .D(c[1524]), .CLK(clk), .RST(rst), .Q(sreg[1523]) );
  DFF \sreg_reg[1522]  ( .D(c[1523]), .CLK(clk), .RST(rst), .Q(sreg[1522]) );
  DFF \sreg_reg[1521]  ( .D(c[1522]), .CLK(clk), .RST(rst), .Q(sreg[1521]) );
  DFF \sreg_reg[1520]  ( .D(c[1521]), .CLK(clk), .RST(rst), .Q(sreg[1520]) );
  DFF \sreg_reg[1519]  ( .D(c[1520]), .CLK(clk), .RST(rst), .Q(sreg[1519]) );
  DFF \sreg_reg[1518]  ( .D(c[1519]), .CLK(clk), .RST(rst), .Q(sreg[1518]) );
  DFF \sreg_reg[1517]  ( .D(c[1518]), .CLK(clk), .RST(rst), .Q(sreg[1517]) );
  DFF \sreg_reg[1516]  ( .D(c[1517]), .CLK(clk), .RST(rst), .Q(sreg[1516]) );
  DFF \sreg_reg[1515]  ( .D(c[1516]), .CLK(clk), .RST(rst), .Q(sreg[1515]) );
  DFF \sreg_reg[1514]  ( .D(c[1515]), .CLK(clk), .RST(rst), .Q(sreg[1514]) );
  DFF \sreg_reg[1513]  ( .D(c[1514]), .CLK(clk), .RST(rst), .Q(sreg[1513]) );
  DFF \sreg_reg[1512]  ( .D(c[1513]), .CLK(clk), .RST(rst), .Q(sreg[1512]) );
  DFF \sreg_reg[1511]  ( .D(c[1512]), .CLK(clk), .RST(rst), .Q(sreg[1511]) );
  DFF \sreg_reg[1510]  ( .D(c[1511]), .CLK(clk), .RST(rst), .Q(sreg[1510]) );
  DFF \sreg_reg[1509]  ( .D(c[1510]), .CLK(clk), .RST(rst), .Q(sreg[1509]) );
  DFF \sreg_reg[1508]  ( .D(c[1509]), .CLK(clk), .RST(rst), .Q(sreg[1508]) );
  DFF \sreg_reg[1507]  ( .D(c[1508]), .CLK(clk), .RST(rst), .Q(sreg[1507]) );
  DFF \sreg_reg[1506]  ( .D(c[1507]), .CLK(clk), .RST(rst), .Q(sreg[1506]) );
  DFF \sreg_reg[1505]  ( .D(c[1506]), .CLK(clk), .RST(rst), .Q(sreg[1505]) );
  DFF \sreg_reg[1504]  ( .D(c[1505]), .CLK(clk), .RST(rst), .Q(sreg[1504]) );
  DFF \sreg_reg[1503]  ( .D(c[1504]), .CLK(clk), .RST(rst), .Q(sreg[1503]) );
  DFF \sreg_reg[1502]  ( .D(c[1503]), .CLK(clk), .RST(rst), .Q(sreg[1502]) );
  DFF \sreg_reg[1501]  ( .D(c[1502]), .CLK(clk), .RST(rst), .Q(sreg[1501]) );
  DFF \sreg_reg[1500]  ( .D(c[1501]), .CLK(clk), .RST(rst), .Q(sreg[1500]) );
  DFF \sreg_reg[1499]  ( .D(c[1500]), .CLK(clk), .RST(rst), .Q(sreg[1499]) );
  DFF \sreg_reg[1498]  ( .D(c[1499]), .CLK(clk), .RST(rst), .Q(sreg[1498]) );
  DFF \sreg_reg[1497]  ( .D(c[1498]), .CLK(clk), .RST(rst), .Q(sreg[1497]) );
  DFF \sreg_reg[1496]  ( .D(c[1497]), .CLK(clk), .RST(rst), .Q(sreg[1496]) );
  DFF \sreg_reg[1495]  ( .D(c[1496]), .CLK(clk), .RST(rst), .Q(sreg[1495]) );
  DFF \sreg_reg[1494]  ( .D(c[1495]), .CLK(clk), .RST(rst), .Q(sreg[1494]) );
  DFF \sreg_reg[1493]  ( .D(c[1494]), .CLK(clk), .RST(rst), .Q(sreg[1493]) );
  DFF \sreg_reg[1492]  ( .D(c[1493]), .CLK(clk), .RST(rst), .Q(sreg[1492]) );
  DFF \sreg_reg[1491]  ( .D(c[1492]), .CLK(clk), .RST(rst), .Q(sreg[1491]) );
  DFF \sreg_reg[1490]  ( .D(c[1491]), .CLK(clk), .RST(rst), .Q(sreg[1490]) );
  DFF \sreg_reg[1489]  ( .D(c[1490]), .CLK(clk), .RST(rst), .Q(sreg[1489]) );
  DFF \sreg_reg[1488]  ( .D(c[1489]), .CLK(clk), .RST(rst), .Q(sreg[1488]) );
  DFF \sreg_reg[1487]  ( .D(c[1488]), .CLK(clk), .RST(rst), .Q(sreg[1487]) );
  DFF \sreg_reg[1486]  ( .D(c[1487]), .CLK(clk), .RST(rst), .Q(sreg[1486]) );
  DFF \sreg_reg[1485]  ( .D(c[1486]), .CLK(clk), .RST(rst), .Q(sreg[1485]) );
  DFF \sreg_reg[1484]  ( .D(c[1485]), .CLK(clk), .RST(rst), .Q(sreg[1484]) );
  DFF \sreg_reg[1483]  ( .D(c[1484]), .CLK(clk), .RST(rst), .Q(sreg[1483]) );
  DFF \sreg_reg[1482]  ( .D(c[1483]), .CLK(clk), .RST(rst), .Q(sreg[1482]) );
  DFF \sreg_reg[1481]  ( .D(c[1482]), .CLK(clk), .RST(rst), .Q(sreg[1481]) );
  DFF \sreg_reg[1480]  ( .D(c[1481]), .CLK(clk), .RST(rst), .Q(sreg[1480]) );
  DFF \sreg_reg[1479]  ( .D(c[1480]), .CLK(clk), .RST(rst), .Q(sreg[1479]) );
  DFF \sreg_reg[1478]  ( .D(c[1479]), .CLK(clk), .RST(rst), .Q(sreg[1478]) );
  DFF \sreg_reg[1477]  ( .D(c[1478]), .CLK(clk), .RST(rst), .Q(sreg[1477]) );
  DFF \sreg_reg[1476]  ( .D(c[1477]), .CLK(clk), .RST(rst), .Q(sreg[1476]) );
  DFF \sreg_reg[1475]  ( .D(c[1476]), .CLK(clk), .RST(rst), .Q(sreg[1475]) );
  DFF \sreg_reg[1474]  ( .D(c[1475]), .CLK(clk), .RST(rst), .Q(sreg[1474]) );
  DFF \sreg_reg[1473]  ( .D(c[1474]), .CLK(clk), .RST(rst), .Q(sreg[1473]) );
  DFF \sreg_reg[1472]  ( .D(c[1473]), .CLK(clk), .RST(rst), .Q(sreg[1472]) );
  DFF \sreg_reg[1471]  ( .D(c[1472]), .CLK(clk), .RST(rst), .Q(sreg[1471]) );
  DFF \sreg_reg[1470]  ( .D(c[1471]), .CLK(clk), .RST(rst), .Q(sreg[1470]) );
  DFF \sreg_reg[1469]  ( .D(c[1470]), .CLK(clk), .RST(rst), .Q(sreg[1469]) );
  DFF \sreg_reg[1468]  ( .D(c[1469]), .CLK(clk), .RST(rst), .Q(sreg[1468]) );
  DFF \sreg_reg[1467]  ( .D(c[1468]), .CLK(clk), .RST(rst), .Q(sreg[1467]) );
  DFF \sreg_reg[1466]  ( .D(c[1467]), .CLK(clk), .RST(rst), .Q(sreg[1466]) );
  DFF \sreg_reg[1465]  ( .D(c[1466]), .CLK(clk), .RST(rst), .Q(sreg[1465]) );
  DFF \sreg_reg[1464]  ( .D(c[1465]), .CLK(clk), .RST(rst), .Q(sreg[1464]) );
  DFF \sreg_reg[1463]  ( .D(c[1464]), .CLK(clk), .RST(rst), .Q(sreg[1463]) );
  DFF \sreg_reg[1462]  ( .D(c[1463]), .CLK(clk), .RST(rst), .Q(sreg[1462]) );
  DFF \sreg_reg[1461]  ( .D(c[1462]), .CLK(clk), .RST(rst), .Q(sreg[1461]) );
  DFF \sreg_reg[1460]  ( .D(c[1461]), .CLK(clk), .RST(rst), .Q(sreg[1460]) );
  DFF \sreg_reg[1459]  ( .D(c[1460]), .CLK(clk), .RST(rst), .Q(sreg[1459]) );
  DFF \sreg_reg[1458]  ( .D(c[1459]), .CLK(clk), .RST(rst), .Q(sreg[1458]) );
  DFF \sreg_reg[1457]  ( .D(c[1458]), .CLK(clk), .RST(rst), .Q(sreg[1457]) );
  DFF \sreg_reg[1456]  ( .D(c[1457]), .CLK(clk), .RST(rst), .Q(sreg[1456]) );
  DFF \sreg_reg[1455]  ( .D(c[1456]), .CLK(clk), .RST(rst), .Q(sreg[1455]) );
  DFF \sreg_reg[1454]  ( .D(c[1455]), .CLK(clk), .RST(rst), .Q(sreg[1454]) );
  DFF \sreg_reg[1453]  ( .D(c[1454]), .CLK(clk), .RST(rst), .Q(sreg[1453]) );
  DFF \sreg_reg[1452]  ( .D(c[1453]), .CLK(clk), .RST(rst), .Q(sreg[1452]) );
  DFF \sreg_reg[1451]  ( .D(c[1452]), .CLK(clk), .RST(rst), .Q(sreg[1451]) );
  DFF \sreg_reg[1450]  ( .D(c[1451]), .CLK(clk), .RST(rst), .Q(sreg[1450]) );
  DFF \sreg_reg[1449]  ( .D(c[1450]), .CLK(clk), .RST(rst), .Q(sreg[1449]) );
  DFF \sreg_reg[1448]  ( .D(c[1449]), .CLK(clk), .RST(rst), .Q(sreg[1448]) );
  DFF \sreg_reg[1447]  ( .D(c[1448]), .CLK(clk), .RST(rst), .Q(sreg[1447]) );
  DFF \sreg_reg[1446]  ( .D(c[1447]), .CLK(clk), .RST(rst), .Q(sreg[1446]) );
  DFF \sreg_reg[1445]  ( .D(c[1446]), .CLK(clk), .RST(rst), .Q(sreg[1445]) );
  DFF \sreg_reg[1444]  ( .D(c[1445]), .CLK(clk), .RST(rst), .Q(sreg[1444]) );
  DFF \sreg_reg[1443]  ( .D(c[1444]), .CLK(clk), .RST(rst), .Q(sreg[1443]) );
  DFF \sreg_reg[1442]  ( .D(c[1443]), .CLK(clk), .RST(rst), .Q(sreg[1442]) );
  DFF \sreg_reg[1441]  ( .D(c[1442]), .CLK(clk), .RST(rst), .Q(sreg[1441]) );
  DFF \sreg_reg[1440]  ( .D(c[1441]), .CLK(clk), .RST(rst), .Q(sreg[1440]) );
  DFF \sreg_reg[1439]  ( .D(c[1440]), .CLK(clk), .RST(rst), .Q(sreg[1439]) );
  DFF \sreg_reg[1438]  ( .D(c[1439]), .CLK(clk), .RST(rst), .Q(sreg[1438]) );
  DFF \sreg_reg[1437]  ( .D(c[1438]), .CLK(clk), .RST(rst), .Q(sreg[1437]) );
  DFF \sreg_reg[1436]  ( .D(c[1437]), .CLK(clk), .RST(rst), .Q(sreg[1436]) );
  DFF \sreg_reg[1435]  ( .D(c[1436]), .CLK(clk), .RST(rst), .Q(sreg[1435]) );
  DFF \sreg_reg[1434]  ( .D(c[1435]), .CLK(clk), .RST(rst), .Q(sreg[1434]) );
  DFF \sreg_reg[1433]  ( .D(c[1434]), .CLK(clk), .RST(rst), .Q(sreg[1433]) );
  DFF \sreg_reg[1432]  ( .D(c[1433]), .CLK(clk), .RST(rst), .Q(sreg[1432]) );
  DFF \sreg_reg[1431]  ( .D(c[1432]), .CLK(clk), .RST(rst), .Q(sreg[1431]) );
  DFF \sreg_reg[1430]  ( .D(c[1431]), .CLK(clk), .RST(rst), .Q(sreg[1430]) );
  DFF \sreg_reg[1429]  ( .D(c[1430]), .CLK(clk), .RST(rst), .Q(sreg[1429]) );
  DFF \sreg_reg[1428]  ( .D(c[1429]), .CLK(clk), .RST(rst), .Q(sreg[1428]) );
  DFF \sreg_reg[1427]  ( .D(c[1428]), .CLK(clk), .RST(rst), .Q(sreg[1427]) );
  DFF \sreg_reg[1426]  ( .D(c[1427]), .CLK(clk), .RST(rst), .Q(sreg[1426]) );
  DFF \sreg_reg[1425]  ( .D(c[1426]), .CLK(clk), .RST(rst), .Q(sreg[1425]) );
  DFF \sreg_reg[1424]  ( .D(c[1425]), .CLK(clk), .RST(rst), .Q(sreg[1424]) );
  DFF \sreg_reg[1423]  ( .D(c[1424]), .CLK(clk), .RST(rst), .Q(sreg[1423]) );
  DFF \sreg_reg[1422]  ( .D(c[1423]), .CLK(clk), .RST(rst), .Q(sreg[1422]) );
  DFF \sreg_reg[1421]  ( .D(c[1422]), .CLK(clk), .RST(rst), .Q(sreg[1421]) );
  DFF \sreg_reg[1420]  ( .D(c[1421]), .CLK(clk), .RST(rst), .Q(sreg[1420]) );
  DFF \sreg_reg[1419]  ( .D(c[1420]), .CLK(clk), .RST(rst), .Q(sreg[1419]) );
  DFF \sreg_reg[1418]  ( .D(c[1419]), .CLK(clk), .RST(rst), .Q(sreg[1418]) );
  DFF \sreg_reg[1417]  ( .D(c[1418]), .CLK(clk), .RST(rst), .Q(sreg[1417]) );
  DFF \sreg_reg[1416]  ( .D(c[1417]), .CLK(clk), .RST(rst), .Q(sreg[1416]) );
  DFF \sreg_reg[1415]  ( .D(c[1416]), .CLK(clk), .RST(rst), .Q(sreg[1415]) );
  DFF \sreg_reg[1414]  ( .D(c[1415]), .CLK(clk), .RST(rst), .Q(sreg[1414]) );
  DFF \sreg_reg[1413]  ( .D(c[1414]), .CLK(clk), .RST(rst), .Q(sreg[1413]) );
  DFF \sreg_reg[1412]  ( .D(c[1413]), .CLK(clk), .RST(rst), .Q(sreg[1412]) );
  DFF \sreg_reg[1411]  ( .D(c[1412]), .CLK(clk), .RST(rst), .Q(sreg[1411]) );
  DFF \sreg_reg[1410]  ( .D(c[1411]), .CLK(clk), .RST(rst), .Q(sreg[1410]) );
  DFF \sreg_reg[1409]  ( .D(c[1410]), .CLK(clk), .RST(rst), .Q(sreg[1409]) );
  DFF \sreg_reg[1408]  ( .D(c[1409]), .CLK(clk), .RST(rst), .Q(sreg[1408]) );
  DFF \sreg_reg[1407]  ( .D(c[1408]), .CLK(clk), .RST(rst), .Q(sreg[1407]) );
  DFF \sreg_reg[1406]  ( .D(c[1407]), .CLK(clk), .RST(rst), .Q(sreg[1406]) );
  DFF \sreg_reg[1405]  ( .D(c[1406]), .CLK(clk), .RST(rst), .Q(sreg[1405]) );
  DFF \sreg_reg[1404]  ( .D(c[1405]), .CLK(clk), .RST(rst), .Q(sreg[1404]) );
  DFF \sreg_reg[1403]  ( .D(c[1404]), .CLK(clk), .RST(rst), .Q(sreg[1403]) );
  DFF \sreg_reg[1402]  ( .D(c[1403]), .CLK(clk), .RST(rst), .Q(sreg[1402]) );
  DFF \sreg_reg[1401]  ( .D(c[1402]), .CLK(clk), .RST(rst), .Q(sreg[1401]) );
  DFF \sreg_reg[1400]  ( .D(c[1401]), .CLK(clk), .RST(rst), .Q(sreg[1400]) );
  DFF \sreg_reg[1399]  ( .D(c[1400]), .CLK(clk), .RST(rst), .Q(sreg[1399]) );
  DFF \sreg_reg[1398]  ( .D(c[1399]), .CLK(clk), .RST(rst), .Q(sreg[1398]) );
  DFF \sreg_reg[1397]  ( .D(c[1398]), .CLK(clk), .RST(rst), .Q(sreg[1397]) );
  DFF \sreg_reg[1396]  ( .D(c[1397]), .CLK(clk), .RST(rst), .Q(sreg[1396]) );
  DFF \sreg_reg[1395]  ( .D(c[1396]), .CLK(clk), .RST(rst), .Q(sreg[1395]) );
  DFF \sreg_reg[1394]  ( .D(c[1395]), .CLK(clk), .RST(rst), .Q(sreg[1394]) );
  DFF \sreg_reg[1393]  ( .D(c[1394]), .CLK(clk), .RST(rst), .Q(sreg[1393]) );
  DFF \sreg_reg[1392]  ( .D(c[1393]), .CLK(clk), .RST(rst), .Q(sreg[1392]) );
  DFF \sreg_reg[1391]  ( .D(c[1392]), .CLK(clk), .RST(rst), .Q(sreg[1391]) );
  DFF \sreg_reg[1390]  ( .D(c[1391]), .CLK(clk), .RST(rst), .Q(sreg[1390]) );
  DFF \sreg_reg[1389]  ( .D(c[1390]), .CLK(clk), .RST(rst), .Q(sreg[1389]) );
  DFF \sreg_reg[1388]  ( .D(c[1389]), .CLK(clk), .RST(rst), .Q(sreg[1388]) );
  DFF \sreg_reg[1387]  ( .D(c[1388]), .CLK(clk), .RST(rst), .Q(sreg[1387]) );
  DFF \sreg_reg[1386]  ( .D(c[1387]), .CLK(clk), .RST(rst), .Q(sreg[1386]) );
  DFF \sreg_reg[1385]  ( .D(c[1386]), .CLK(clk), .RST(rst), .Q(sreg[1385]) );
  DFF \sreg_reg[1384]  ( .D(c[1385]), .CLK(clk), .RST(rst), .Q(sreg[1384]) );
  DFF \sreg_reg[1383]  ( .D(c[1384]), .CLK(clk), .RST(rst), .Q(sreg[1383]) );
  DFF \sreg_reg[1382]  ( .D(c[1383]), .CLK(clk), .RST(rst), .Q(sreg[1382]) );
  DFF \sreg_reg[1381]  ( .D(c[1382]), .CLK(clk), .RST(rst), .Q(sreg[1381]) );
  DFF \sreg_reg[1380]  ( .D(c[1381]), .CLK(clk), .RST(rst), .Q(sreg[1380]) );
  DFF \sreg_reg[1379]  ( .D(c[1380]), .CLK(clk), .RST(rst), .Q(sreg[1379]) );
  DFF \sreg_reg[1378]  ( .D(c[1379]), .CLK(clk), .RST(rst), .Q(sreg[1378]) );
  DFF \sreg_reg[1377]  ( .D(c[1378]), .CLK(clk), .RST(rst), .Q(sreg[1377]) );
  DFF \sreg_reg[1376]  ( .D(c[1377]), .CLK(clk), .RST(rst), .Q(sreg[1376]) );
  DFF \sreg_reg[1375]  ( .D(c[1376]), .CLK(clk), .RST(rst), .Q(sreg[1375]) );
  DFF \sreg_reg[1374]  ( .D(c[1375]), .CLK(clk), .RST(rst), .Q(sreg[1374]) );
  DFF \sreg_reg[1373]  ( .D(c[1374]), .CLK(clk), .RST(rst), .Q(sreg[1373]) );
  DFF \sreg_reg[1372]  ( .D(c[1373]), .CLK(clk), .RST(rst), .Q(sreg[1372]) );
  DFF \sreg_reg[1371]  ( .D(c[1372]), .CLK(clk), .RST(rst), .Q(sreg[1371]) );
  DFF \sreg_reg[1370]  ( .D(c[1371]), .CLK(clk), .RST(rst), .Q(sreg[1370]) );
  DFF \sreg_reg[1369]  ( .D(c[1370]), .CLK(clk), .RST(rst), .Q(sreg[1369]) );
  DFF \sreg_reg[1368]  ( .D(c[1369]), .CLK(clk), .RST(rst), .Q(sreg[1368]) );
  DFF \sreg_reg[1367]  ( .D(c[1368]), .CLK(clk), .RST(rst), .Q(sreg[1367]) );
  DFF \sreg_reg[1366]  ( .D(c[1367]), .CLK(clk), .RST(rst), .Q(sreg[1366]) );
  DFF \sreg_reg[1365]  ( .D(c[1366]), .CLK(clk), .RST(rst), .Q(sreg[1365]) );
  DFF \sreg_reg[1364]  ( .D(c[1365]), .CLK(clk), .RST(rst), .Q(sreg[1364]) );
  DFF \sreg_reg[1363]  ( .D(c[1364]), .CLK(clk), .RST(rst), .Q(sreg[1363]) );
  DFF \sreg_reg[1362]  ( .D(c[1363]), .CLK(clk), .RST(rst), .Q(sreg[1362]) );
  DFF \sreg_reg[1361]  ( .D(c[1362]), .CLK(clk), .RST(rst), .Q(sreg[1361]) );
  DFF \sreg_reg[1360]  ( .D(c[1361]), .CLK(clk), .RST(rst), .Q(sreg[1360]) );
  DFF \sreg_reg[1359]  ( .D(c[1360]), .CLK(clk), .RST(rst), .Q(sreg[1359]) );
  DFF \sreg_reg[1358]  ( .D(c[1359]), .CLK(clk), .RST(rst), .Q(sreg[1358]) );
  DFF \sreg_reg[1357]  ( .D(c[1358]), .CLK(clk), .RST(rst), .Q(sreg[1357]) );
  DFF \sreg_reg[1356]  ( .D(c[1357]), .CLK(clk), .RST(rst), .Q(sreg[1356]) );
  DFF \sreg_reg[1355]  ( .D(c[1356]), .CLK(clk), .RST(rst), .Q(sreg[1355]) );
  DFF \sreg_reg[1354]  ( .D(c[1355]), .CLK(clk), .RST(rst), .Q(sreg[1354]) );
  DFF \sreg_reg[1353]  ( .D(c[1354]), .CLK(clk), .RST(rst), .Q(sreg[1353]) );
  DFF \sreg_reg[1352]  ( .D(c[1353]), .CLK(clk), .RST(rst), .Q(sreg[1352]) );
  DFF \sreg_reg[1351]  ( .D(c[1352]), .CLK(clk), .RST(rst), .Q(sreg[1351]) );
  DFF \sreg_reg[1350]  ( .D(c[1351]), .CLK(clk), .RST(rst), .Q(sreg[1350]) );
  DFF \sreg_reg[1349]  ( .D(c[1350]), .CLK(clk), .RST(rst), .Q(sreg[1349]) );
  DFF \sreg_reg[1348]  ( .D(c[1349]), .CLK(clk), .RST(rst), .Q(sreg[1348]) );
  DFF \sreg_reg[1347]  ( .D(c[1348]), .CLK(clk), .RST(rst), .Q(sreg[1347]) );
  DFF \sreg_reg[1346]  ( .D(c[1347]), .CLK(clk), .RST(rst), .Q(sreg[1346]) );
  DFF \sreg_reg[1345]  ( .D(c[1346]), .CLK(clk), .RST(rst), .Q(sreg[1345]) );
  DFF \sreg_reg[1344]  ( .D(c[1345]), .CLK(clk), .RST(rst), .Q(sreg[1344]) );
  DFF \sreg_reg[1343]  ( .D(c[1344]), .CLK(clk), .RST(rst), .Q(sreg[1343]) );
  DFF \sreg_reg[1342]  ( .D(c[1343]), .CLK(clk), .RST(rst), .Q(sreg[1342]) );
  DFF \sreg_reg[1341]  ( .D(c[1342]), .CLK(clk), .RST(rst), .Q(sreg[1341]) );
  DFF \sreg_reg[1340]  ( .D(c[1341]), .CLK(clk), .RST(rst), .Q(sreg[1340]) );
  DFF \sreg_reg[1339]  ( .D(c[1340]), .CLK(clk), .RST(rst), .Q(sreg[1339]) );
  DFF \sreg_reg[1338]  ( .D(c[1339]), .CLK(clk), .RST(rst), .Q(sreg[1338]) );
  DFF \sreg_reg[1337]  ( .D(c[1338]), .CLK(clk), .RST(rst), .Q(sreg[1337]) );
  DFF \sreg_reg[1336]  ( .D(c[1337]), .CLK(clk), .RST(rst), .Q(sreg[1336]) );
  DFF \sreg_reg[1335]  ( .D(c[1336]), .CLK(clk), .RST(rst), .Q(sreg[1335]) );
  DFF \sreg_reg[1334]  ( .D(c[1335]), .CLK(clk), .RST(rst), .Q(sreg[1334]) );
  DFF \sreg_reg[1333]  ( .D(c[1334]), .CLK(clk), .RST(rst), .Q(sreg[1333]) );
  DFF \sreg_reg[1332]  ( .D(c[1333]), .CLK(clk), .RST(rst), .Q(sreg[1332]) );
  DFF \sreg_reg[1331]  ( .D(c[1332]), .CLK(clk), .RST(rst), .Q(sreg[1331]) );
  DFF \sreg_reg[1330]  ( .D(c[1331]), .CLK(clk), .RST(rst), .Q(sreg[1330]) );
  DFF \sreg_reg[1329]  ( .D(c[1330]), .CLK(clk), .RST(rst), .Q(sreg[1329]) );
  DFF \sreg_reg[1328]  ( .D(c[1329]), .CLK(clk), .RST(rst), .Q(sreg[1328]) );
  DFF \sreg_reg[1327]  ( .D(c[1328]), .CLK(clk), .RST(rst), .Q(sreg[1327]) );
  DFF \sreg_reg[1326]  ( .D(c[1327]), .CLK(clk), .RST(rst), .Q(sreg[1326]) );
  DFF \sreg_reg[1325]  ( .D(c[1326]), .CLK(clk), .RST(rst), .Q(sreg[1325]) );
  DFF \sreg_reg[1324]  ( .D(c[1325]), .CLK(clk), .RST(rst), .Q(sreg[1324]) );
  DFF \sreg_reg[1323]  ( .D(c[1324]), .CLK(clk), .RST(rst), .Q(sreg[1323]) );
  DFF \sreg_reg[1322]  ( .D(c[1323]), .CLK(clk), .RST(rst), .Q(sreg[1322]) );
  DFF \sreg_reg[1321]  ( .D(c[1322]), .CLK(clk), .RST(rst), .Q(sreg[1321]) );
  DFF \sreg_reg[1320]  ( .D(c[1321]), .CLK(clk), .RST(rst), .Q(sreg[1320]) );
  DFF \sreg_reg[1319]  ( .D(c[1320]), .CLK(clk), .RST(rst), .Q(sreg[1319]) );
  DFF \sreg_reg[1318]  ( .D(c[1319]), .CLK(clk), .RST(rst), .Q(sreg[1318]) );
  DFF \sreg_reg[1317]  ( .D(c[1318]), .CLK(clk), .RST(rst), .Q(sreg[1317]) );
  DFF \sreg_reg[1316]  ( .D(c[1317]), .CLK(clk), .RST(rst), .Q(sreg[1316]) );
  DFF \sreg_reg[1315]  ( .D(c[1316]), .CLK(clk), .RST(rst), .Q(sreg[1315]) );
  DFF \sreg_reg[1314]  ( .D(c[1315]), .CLK(clk), .RST(rst), .Q(sreg[1314]) );
  DFF \sreg_reg[1313]  ( .D(c[1314]), .CLK(clk), .RST(rst), .Q(sreg[1313]) );
  DFF \sreg_reg[1312]  ( .D(c[1313]), .CLK(clk), .RST(rst), .Q(sreg[1312]) );
  DFF \sreg_reg[1311]  ( .D(c[1312]), .CLK(clk), .RST(rst), .Q(sreg[1311]) );
  DFF \sreg_reg[1310]  ( .D(c[1311]), .CLK(clk), .RST(rst), .Q(sreg[1310]) );
  DFF \sreg_reg[1309]  ( .D(c[1310]), .CLK(clk), .RST(rst), .Q(sreg[1309]) );
  DFF \sreg_reg[1308]  ( .D(c[1309]), .CLK(clk), .RST(rst), .Q(sreg[1308]) );
  DFF \sreg_reg[1307]  ( .D(c[1308]), .CLK(clk), .RST(rst), .Q(sreg[1307]) );
  DFF \sreg_reg[1306]  ( .D(c[1307]), .CLK(clk), .RST(rst), .Q(sreg[1306]) );
  DFF \sreg_reg[1305]  ( .D(c[1306]), .CLK(clk), .RST(rst), .Q(sreg[1305]) );
  DFF \sreg_reg[1304]  ( .D(c[1305]), .CLK(clk), .RST(rst), .Q(sreg[1304]) );
  DFF \sreg_reg[1303]  ( .D(c[1304]), .CLK(clk), .RST(rst), .Q(sreg[1303]) );
  DFF \sreg_reg[1302]  ( .D(c[1303]), .CLK(clk), .RST(rst), .Q(sreg[1302]) );
  DFF \sreg_reg[1301]  ( .D(c[1302]), .CLK(clk), .RST(rst), .Q(sreg[1301]) );
  DFF \sreg_reg[1300]  ( .D(c[1301]), .CLK(clk), .RST(rst), .Q(sreg[1300]) );
  DFF \sreg_reg[1299]  ( .D(c[1300]), .CLK(clk), .RST(rst), .Q(sreg[1299]) );
  DFF \sreg_reg[1298]  ( .D(c[1299]), .CLK(clk), .RST(rst), .Q(sreg[1298]) );
  DFF \sreg_reg[1297]  ( .D(c[1298]), .CLK(clk), .RST(rst), .Q(sreg[1297]) );
  DFF \sreg_reg[1296]  ( .D(c[1297]), .CLK(clk), .RST(rst), .Q(sreg[1296]) );
  DFF \sreg_reg[1295]  ( .D(c[1296]), .CLK(clk), .RST(rst), .Q(sreg[1295]) );
  DFF \sreg_reg[1294]  ( .D(c[1295]), .CLK(clk), .RST(rst), .Q(sreg[1294]) );
  DFF \sreg_reg[1293]  ( .D(c[1294]), .CLK(clk), .RST(rst), .Q(sreg[1293]) );
  DFF \sreg_reg[1292]  ( .D(c[1293]), .CLK(clk), .RST(rst), .Q(sreg[1292]) );
  DFF \sreg_reg[1291]  ( .D(c[1292]), .CLK(clk), .RST(rst), .Q(sreg[1291]) );
  DFF \sreg_reg[1290]  ( .D(c[1291]), .CLK(clk), .RST(rst), .Q(sreg[1290]) );
  DFF \sreg_reg[1289]  ( .D(c[1290]), .CLK(clk), .RST(rst), .Q(sreg[1289]) );
  DFF \sreg_reg[1288]  ( .D(c[1289]), .CLK(clk), .RST(rst), .Q(sreg[1288]) );
  DFF \sreg_reg[1287]  ( .D(c[1288]), .CLK(clk), .RST(rst), .Q(sreg[1287]) );
  DFF \sreg_reg[1286]  ( .D(c[1287]), .CLK(clk), .RST(rst), .Q(sreg[1286]) );
  DFF \sreg_reg[1285]  ( .D(c[1286]), .CLK(clk), .RST(rst), .Q(sreg[1285]) );
  DFF \sreg_reg[1284]  ( .D(c[1285]), .CLK(clk), .RST(rst), .Q(sreg[1284]) );
  DFF \sreg_reg[1283]  ( .D(c[1284]), .CLK(clk), .RST(rst), .Q(sreg[1283]) );
  DFF \sreg_reg[1282]  ( .D(c[1283]), .CLK(clk), .RST(rst), .Q(sreg[1282]) );
  DFF \sreg_reg[1281]  ( .D(c[1282]), .CLK(clk), .RST(rst), .Q(sreg[1281]) );
  DFF \sreg_reg[1280]  ( .D(c[1281]), .CLK(clk), .RST(rst), .Q(sreg[1280]) );
  DFF \sreg_reg[1279]  ( .D(c[1280]), .CLK(clk), .RST(rst), .Q(sreg[1279]) );
  DFF \sreg_reg[1278]  ( .D(c[1279]), .CLK(clk), .RST(rst), .Q(sreg[1278]) );
  DFF \sreg_reg[1277]  ( .D(c[1278]), .CLK(clk), .RST(rst), .Q(sreg[1277]) );
  DFF \sreg_reg[1276]  ( .D(c[1277]), .CLK(clk), .RST(rst), .Q(sreg[1276]) );
  DFF \sreg_reg[1275]  ( .D(c[1276]), .CLK(clk), .RST(rst), .Q(sreg[1275]) );
  DFF \sreg_reg[1274]  ( .D(c[1275]), .CLK(clk), .RST(rst), .Q(sreg[1274]) );
  DFF \sreg_reg[1273]  ( .D(c[1274]), .CLK(clk), .RST(rst), .Q(sreg[1273]) );
  DFF \sreg_reg[1272]  ( .D(c[1273]), .CLK(clk), .RST(rst), .Q(sreg[1272]) );
  DFF \sreg_reg[1271]  ( .D(c[1272]), .CLK(clk), .RST(rst), .Q(sreg[1271]) );
  DFF \sreg_reg[1270]  ( .D(c[1271]), .CLK(clk), .RST(rst), .Q(sreg[1270]) );
  DFF \sreg_reg[1269]  ( .D(c[1270]), .CLK(clk), .RST(rst), .Q(sreg[1269]) );
  DFF \sreg_reg[1268]  ( .D(c[1269]), .CLK(clk), .RST(rst), .Q(sreg[1268]) );
  DFF \sreg_reg[1267]  ( .D(c[1268]), .CLK(clk), .RST(rst), .Q(sreg[1267]) );
  DFF \sreg_reg[1266]  ( .D(c[1267]), .CLK(clk), .RST(rst), .Q(sreg[1266]) );
  DFF \sreg_reg[1265]  ( .D(c[1266]), .CLK(clk), .RST(rst), .Q(sreg[1265]) );
  DFF \sreg_reg[1264]  ( .D(c[1265]), .CLK(clk), .RST(rst), .Q(sreg[1264]) );
  DFF \sreg_reg[1263]  ( .D(c[1264]), .CLK(clk), .RST(rst), .Q(sreg[1263]) );
  DFF \sreg_reg[1262]  ( .D(c[1263]), .CLK(clk), .RST(rst), .Q(sreg[1262]) );
  DFF \sreg_reg[1261]  ( .D(c[1262]), .CLK(clk), .RST(rst), .Q(sreg[1261]) );
  DFF \sreg_reg[1260]  ( .D(c[1261]), .CLK(clk), .RST(rst), .Q(sreg[1260]) );
  DFF \sreg_reg[1259]  ( .D(c[1260]), .CLK(clk), .RST(rst), .Q(sreg[1259]) );
  DFF \sreg_reg[1258]  ( .D(c[1259]), .CLK(clk), .RST(rst), .Q(sreg[1258]) );
  DFF \sreg_reg[1257]  ( .D(c[1258]), .CLK(clk), .RST(rst), .Q(sreg[1257]) );
  DFF \sreg_reg[1256]  ( .D(c[1257]), .CLK(clk), .RST(rst), .Q(sreg[1256]) );
  DFF \sreg_reg[1255]  ( .D(c[1256]), .CLK(clk), .RST(rst), .Q(sreg[1255]) );
  DFF \sreg_reg[1254]  ( .D(c[1255]), .CLK(clk), .RST(rst), .Q(sreg[1254]) );
  DFF \sreg_reg[1253]  ( .D(c[1254]), .CLK(clk), .RST(rst), .Q(sreg[1253]) );
  DFF \sreg_reg[1252]  ( .D(c[1253]), .CLK(clk), .RST(rst), .Q(sreg[1252]) );
  DFF \sreg_reg[1251]  ( .D(c[1252]), .CLK(clk), .RST(rst), .Q(sreg[1251]) );
  DFF \sreg_reg[1250]  ( .D(c[1251]), .CLK(clk), .RST(rst), .Q(sreg[1250]) );
  DFF \sreg_reg[1249]  ( .D(c[1250]), .CLK(clk), .RST(rst), .Q(sreg[1249]) );
  DFF \sreg_reg[1248]  ( .D(c[1249]), .CLK(clk), .RST(rst), .Q(sreg[1248]) );
  DFF \sreg_reg[1247]  ( .D(c[1248]), .CLK(clk), .RST(rst), .Q(sreg[1247]) );
  DFF \sreg_reg[1246]  ( .D(c[1247]), .CLK(clk), .RST(rst), .Q(sreg[1246]) );
  DFF \sreg_reg[1245]  ( .D(c[1246]), .CLK(clk), .RST(rst), .Q(sreg[1245]) );
  DFF \sreg_reg[1244]  ( .D(c[1245]), .CLK(clk), .RST(rst), .Q(sreg[1244]) );
  DFF \sreg_reg[1243]  ( .D(c[1244]), .CLK(clk), .RST(rst), .Q(sreg[1243]) );
  DFF \sreg_reg[1242]  ( .D(c[1243]), .CLK(clk), .RST(rst), .Q(sreg[1242]) );
  DFF \sreg_reg[1241]  ( .D(c[1242]), .CLK(clk), .RST(rst), .Q(sreg[1241]) );
  DFF \sreg_reg[1240]  ( .D(c[1241]), .CLK(clk), .RST(rst), .Q(sreg[1240]) );
  DFF \sreg_reg[1239]  ( .D(c[1240]), .CLK(clk), .RST(rst), .Q(sreg[1239]) );
  DFF \sreg_reg[1238]  ( .D(c[1239]), .CLK(clk), .RST(rst), .Q(sreg[1238]) );
  DFF \sreg_reg[1237]  ( .D(c[1238]), .CLK(clk), .RST(rst), .Q(sreg[1237]) );
  DFF \sreg_reg[1236]  ( .D(c[1237]), .CLK(clk), .RST(rst), .Q(sreg[1236]) );
  DFF \sreg_reg[1235]  ( .D(c[1236]), .CLK(clk), .RST(rst), .Q(sreg[1235]) );
  DFF \sreg_reg[1234]  ( .D(c[1235]), .CLK(clk), .RST(rst), .Q(sreg[1234]) );
  DFF \sreg_reg[1233]  ( .D(c[1234]), .CLK(clk), .RST(rst), .Q(sreg[1233]) );
  DFF \sreg_reg[1232]  ( .D(c[1233]), .CLK(clk), .RST(rst), .Q(sreg[1232]) );
  DFF \sreg_reg[1231]  ( .D(c[1232]), .CLK(clk), .RST(rst), .Q(sreg[1231]) );
  DFF \sreg_reg[1230]  ( .D(c[1231]), .CLK(clk), .RST(rst), .Q(sreg[1230]) );
  DFF \sreg_reg[1229]  ( .D(c[1230]), .CLK(clk), .RST(rst), .Q(sreg[1229]) );
  DFF \sreg_reg[1228]  ( .D(c[1229]), .CLK(clk), .RST(rst), .Q(sreg[1228]) );
  DFF \sreg_reg[1227]  ( .D(c[1228]), .CLK(clk), .RST(rst), .Q(sreg[1227]) );
  DFF \sreg_reg[1226]  ( .D(c[1227]), .CLK(clk), .RST(rst), .Q(sreg[1226]) );
  DFF \sreg_reg[1225]  ( .D(c[1226]), .CLK(clk), .RST(rst), .Q(sreg[1225]) );
  DFF \sreg_reg[1224]  ( .D(c[1225]), .CLK(clk), .RST(rst), .Q(sreg[1224]) );
  DFF \sreg_reg[1223]  ( .D(c[1224]), .CLK(clk), .RST(rst), .Q(sreg[1223]) );
  DFF \sreg_reg[1222]  ( .D(c[1223]), .CLK(clk), .RST(rst), .Q(sreg[1222]) );
  DFF \sreg_reg[1221]  ( .D(c[1222]), .CLK(clk), .RST(rst), .Q(sreg[1221]) );
  DFF \sreg_reg[1220]  ( .D(c[1221]), .CLK(clk), .RST(rst), .Q(sreg[1220]) );
  DFF \sreg_reg[1219]  ( .D(c[1220]), .CLK(clk), .RST(rst), .Q(sreg[1219]) );
  DFF \sreg_reg[1218]  ( .D(c[1219]), .CLK(clk), .RST(rst), .Q(sreg[1218]) );
  DFF \sreg_reg[1217]  ( .D(c[1218]), .CLK(clk), .RST(rst), .Q(sreg[1217]) );
  DFF \sreg_reg[1216]  ( .D(c[1217]), .CLK(clk), .RST(rst), .Q(sreg[1216]) );
  DFF \sreg_reg[1215]  ( .D(c[1216]), .CLK(clk), .RST(rst), .Q(sreg[1215]) );
  DFF \sreg_reg[1214]  ( .D(c[1215]), .CLK(clk), .RST(rst), .Q(sreg[1214]) );
  DFF \sreg_reg[1213]  ( .D(c[1214]), .CLK(clk), .RST(rst), .Q(sreg[1213]) );
  DFF \sreg_reg[1212]  ( .D(c[1213]), .CLK(clk), .RST(rst), .Q(sreg[1212]) );
  DFF \sreg_reg[1211]  ( .D(c[1212]), .CLK(clk), .RST(rst), .Q(sreg[1211]) );
  DFF \sreg_reg[1210]  ( .D(c[1211]), .CLK(clk), .RST(rst), .Q(sreg[1210]) );
  DFF \sreg_reg[1209]  ( .D(c[1210]), .CLK(clk), .RST(rst), .Q(sreg[1209]) );
  DFF \sreg_reg[1208]  ( .D(c[1209]), .CLK(clk), .RST(rst), .Q(sreg[1208]) );
  DFF \sreg_reg[1207]  ( .D(c[1208]), .CLK(clk), .RST(rst), .Q(sreg[1207]) );
  DFF \sreg_reg[1206]  ( .D(c[1207]), .CLK(clk), .RST(rst), .Q(sreg[1206]) );
  DFF \sreg_reg[1205]  ( .D(c[1206]), .CLK(clk), .RST(rst), .Q(sreg[1205]) );
  DFF \sreg_reg[1204]  ( .D(c[1205]), .CLK(clk), .RST(rst), .Q(sreg[1204]) );
  DFF \sreg_reg[1203]  ( .D(c[1204]), .CLK(clk), .RST(rst), .Q(sreg[1203]) );
  DFF \sreg_reg[1202]  ( .D(c[1203]), .CLK(clk), .RST(rst), .Q(sreg[1202]) );
  DFF \sreg_reg[1201]  ( .D(c[1202]), .CLK(clk), .RST(rst), .Q(sreg[1201]) );
  DFF \sreg_reg[1200]  ( .D(c[1201]), .CLK(clk), .RST(rst), .Q(sreg[1200]) );
  DFF \sreg_reg[1199]  ( .D(c[1200]), .CLK(clk), .RST(rst), .Q(sreg[1199]) );
  DFF \sreg_reg[1198]  ( .D(c[1199]), .CLK(clk), .RST(rst), .Q(sreg[1198]) );
  DFF \sreg_reg[1197]  ( .D(c[1198]), .CLK(clk), .RST(rst), .Q(sreg[1197]) );
  DFF \sreg_reg[1196]  ( .D(c[1197]), .CLK(clk), .RST(rst), .Q(sreg[1196]) );
  DFF \sreg_reg[1195]  ( .D(c[1196]), .CLK(clk), .RST(rst), .Q(sreg[1195]) );
  DFF \sreg_reg[1194]  ( .D(c[1195]), .CLK(clk), .RST(rst), .Q(sreg[1194]) );
  DFF \sreg_reg[1193]  ( .D(c[1194]), .CLK(clk), .RST(rst), .Q(sreg[1193]) );
  DFF \sreg_reg[1192]  ( .D(c[1193]), .CLK(clk), .RST(rst), .Q(sreg[1192]) );
  DFF \sreg_reg[1191]  ( .D(c[1192]), .CLK(clk), .RST(rst), .Q(sreg[1191]) );
  DFF \sreg_reg[1190]  ( .D(c[1191]), .CLK(clk), .RST(rst), .Q(sreg[1190]) );
  DFF \sreg_reg[1189]  ( .D(c[1190]), .CLK(clk), .RST(rst), .Q(sreg[1189]) );
  DFF \sreg_reg[1188]  ( .D(c[1189]), .CLK(clk), .RST(rst), .Q(sreg[1188]) );
  DFF \sreg_reg[1187]  ( .D(c[1188]), .CLK(clk), .RST(rst), .Q(sreg[1187]) );
  DFF \sreg_reg[1186]  ( .D(c[1187]), .CLK(clk), .RST(rst), .Q(sreg[1186]) );
  DFF \sreg_reg[1185]  ( .D(c[1186]), .CLK(clk), .RST(rst), .Q(sreg[1185]) );
  DFF \sreg_reg[1184]  ( .D(c[1185]), .CLK(clk), .RST(rst), .Q(sreg[1184]) );
  DFF \sreg_reg[1183]  ( .D(c[1184]), .CLK(clk), .RST(rst), .Q(sreg[1183]) );
  DFF \sreg_reg[1182]  ( .D(c[1183]), .CLK(clk), .RST(rst), .Q(sreg[1182]) );
  DFF \sreg_reg[1181]  ( .D(c[1182]), .CLK(clk), .RST(rst), .Q(sreg[1181]) );
  DFF \sreg_reg[1180]  ( .D(c[1181]), .CLK(clk), .RST(rst), .Q(sreg[1180]) );
  DFF \sreg_reg[1179]  ( .D(c[1180]), .CLK(clk), .RST(rst), .Q(sreg[1179]) );
  DFF \sreg_reg[1178]  ( .D(c[1179]), .CLK(clk), .RST(rst), .Q(sreg[1178]) );
  DFF \sreg_reg[1177]  ( .D(c[1178]), .CLK(clk), .RST(rst), .Q(sreg[1177]) );
  DFF \sreg_reg[1176]  ( .D(c[1177]), .CLK(clk), .RST(rst), .Q(sreg[1176]) );
  DFF \sreg_reg[1175]  ( .D(c[1176]), .CLK(clk), .RST(rst), .Q(sreg[1175]) );
  DFF \sreg_reg[1174]  ( .D(c[1175]), .CLK(clk), .RST(rst), .Q(sreg[1174]) );
  DFF \sreg_reg[1173]  ( .D(c[1174]), .CLK(clk), .RST(rst), .Q(sreg[1173]) );
  DFF \sreg_reg[1172]  ( .D(c[1173]), .CLK(clk), .RST(rst), .Q(sreg[1172]) );
  DFF \sreg_reg[1171]  ( .D(c[1172]), .CLK(clk), .RST(rst), .Q(sreg[1171]) );
  DFF \sreg_reg[1170]  ( .D(c[1171]), .CLK(clk), .RST(rst), .Q(sreg[1170]) );
  DFF \sreg_reg[1169]  ( .D(c[1170]), .CLK(clk), .RST(rst), .Q(sreg[1169]) );
  DFF \sreg_reg[1168]  ( .D(c[1169]), .CLK(clk), .RST(rst), .Q(sreg[1168]) );
  DFF \sreg_reg[1167]  ( .D(c[1168]), .CLK(clk), .RST(rst), .Q(sreg[1167]) );
  DFF \sreg_reg[1166]  ( .D(c[1167]), .CLK(clk), .RST(rst), .Q(sreg[1166]) );
  DFF \sreg_reg[1165]  ( .D(c[1166]), .CLK(clk), .RST(rst), .Q(sreg[1165]) );
  DFF \sreg_reg[1164]  ( .D(c[1165]), .CLK(clk), .RST(rst), .Q(sreg[1164]) );
  DFF \sreg_reg[1163]  ( .D(c[1164]), .CLK(clk), .RST(rst), .Q(sreg[1163]) );
  DFF \sreg_reg[1162]  ( .D(c[1163]), .CLK(clk), .RST(rst), .Q(sreg[1162]) );
  DFF \sreg_reg[1161]  ( .D(c[1162]), .CLK(clk), .RST(rst), .Q(sreg[1161]) );
  DFF \sreg_reg[1160]  ( .D(c[1161]), .CLK(clk), .RST(rst), .Q(sreg[1160]) );
  DFF \sreg_reg[1159]  ( .D(c[1160]), .CLK(clk), .RST(rst), .Q(sreg[1159]) );
  DFF \sreg_reg[1158]  ( .D(c[1159]), .CLK(clk), .RST(rst), .Q(sreg[1158]) );
  DFF \sreg_reg[1157]  ( .D(c[1158]), .CLK(clk), .RST(rst), .Q(sreg[1157]) );
  DFF \sreg_reg[1156]  ( .D(c[1157]), .CLK(clk), .RST(rst), .Q(sreg[1156]) );
  DFF \sreg_reg[1155]  ( .D(c[1156]), .CLK(clk), .RST(rst), .Q(sreg[1155]) );
  DFF \sreg_reg[1154]  ( .D(c[1155]), .CLK(clk), .RST(rst), .Q(sreg[1154]) );
  DFF \sreg_reg[1153]  ( .D(c[1154]), .CLK(clk), .RST(rst), .Q(sreg[1153]) );
  DFF \sreg_reg[1152]  ( .D(c[1153]), .CLK(clk), .RST(rst), .Q(sreg[1152]) );
  DFF \sreg_reg[1151]  ( .D(c[1152]), .CLK(clk), .RST(rst), .Q(sreg[1151]) );
  DFF \sreg_reg[1150]  ( .D(c[1151]), .CLK(clk), .RST(rst), .Q(sreg[1150]) );
  DFF \sreg_reg[1149]  ( .D(c[1150]), .CLK(clk), .RST(rst), .Q(sreg[1149]) );
  DFF \sreg_reg[1148]  ( .D(c[1149]), .CLK(clk), .RST(rst), .Q(sreg[1148]) );
  DFF \sreg_reg[1147]  ( .D(c[1148]), .CLK(clk), .RST(rst), .Q(sreg[1147]) );
  DFF \sreg_reg[1146]  ( .D(c[1147]), .CLK(clk), .RST(rst), .Q(sreg[1146]) );
  DFF \sreg_reg[1145]  ( .D(c[1146]), .CLK(clk), .RST(rst), .Q(sreg[1145]) );
  DFF \sreg_reg[1144]  ( .D(c[1145]), .CLK(clk), .RST(rst), .Q(sreg[1144]) );
  DFF \sreg_reg[1143]  ( .D(c[1144]), .CLK(clk), .RST(rst), .Q(sreg[1143]) );
  DFF \sreg_reg[1142]  ( .D(c[1143]), .CLK(clk), .RST(rst), .Q(sreg[1142]) );
  DFF \sreg_reg[1141]  ( .D(c[1142]), .CLK(clk), .RST(rst), .Q(sreg[1141]) );
  DFF \sreg_reg[1140]  ( .D(c[1141]), .CLK(clk), .RST(rst), .Q(sreg[1140]) );
  DFF \sreg_reg[1139]  ( .D(c[1140]), .CLK(clk), .RST(rst), .Q(sreg[1139]) );
  DFF \sreg_reg[1138]  ( .D(c[1139]), .CLK(clk), .RST(rst), .Q(sreg[1138]) );
  DFF \sreg_reg[1137]  ( .D(c[1138]), .CLK(clk), .RST(rst), .Q(sreg[1137]) );
  DFF \sreg_reg[1136]  ( .D(c[1137]), .CLK(clk), .RST(rst), .Q(sreg[1136]) );
  DFF \sreg_reg[1135]  ( .D(c[1136]), .CLK(clk), .RST(rst), .Q(sreg[1135]) );
  DFF \sreg_reg[1134]  ( .D(c[1135]), .CLK(clk), .RST(rst), .Q(sreg[1134]) );
  DFF \sreg_reg[1133]  ( .D(c[1134]), .CLK(clk), .RST(rst), .Q(sreg[1133]) );
  DFF \sreg_reg[1132]  ( .D(c[1133]), .CLK(clk), .RST(rst), .Q(sreg[1132]) );
  DFF \sreg_reg[1131]  ( .D(c[1132]), .CLK(clk), .RST(rst), .Q(sreg[1131]) );
  DFF \sreg_reg[1130]  ( .D(c[1131]), .CLK(clk), .RST(rst), .Q(sreg[1130]) );
  DFF \sreg_reg[1129]  ( .D(c[1130]), .CLK(clk), .RST(rst), .Q(sreg[1129]) );
  DFF \sreg_reg[1128]  ( .D(c[1129]), .CLK(clk), .RST(rst), .Q(sreg[1128]) );
  DFF \sreg_reg[1127]  ( .D(c[1128]), .CLK(clk), .RST(rst), .Q(sreg[1127]) );
  DFF \sreg_reg[1126]  ( .D(c[1127]), .CLK(clk), .RST(rst), .Q(sreg[1126]) );
  DFF \sreg_reg[1125]  ( .D(c[1126]), .CLK(clk), .RST(rst), .Q(sreg[1125]) );
  DFF \sreg_reg[1124]  ( .D(c[1125]), .CLK(clk), .RST(rst), .Q(sreg[1124]) );
  DFF \sreg_reg[1123]  ( .D(c[1124]), .CLK(clk), .RST(rst), .Q(sreg[1123]) );
  DFF \sreg_reg[1122]  ( .D(c[1123]), .CLK(clk), .RST(rst), .Q(sreg[1122]) );
  DFF \sreg_reg[1121]  ( .D(c[1122]), .CLK(clk), .RST(rst), .Q(sreg[1121]) );
  DFF \sreg_reg[1120]  ( .D(c[1121]), .CLK(clk), .RST(rst), .Q(sreg[1120]) );
  DFF \sreg_reg[1119]  ( .D(c[1120]), .CLK(clk), .RST(rst), .Q(sreg[1119]) );
  DFF \sreg_reg[1118]  ( .D(c[1119]), .CLK(clk), .RST(rst), .Q(sreg[1118]) );
  DFF \sreg_reg[1117]  ( .D(c[1118]), .CLK(clk), .RST(rst), .Q(sreg[1117]) );
  DFF \sreg_reg[1116]  ( .D(c[1117]), .CLK(clk), .RST(rst), .Q(sreg[1116]) );
  DFF \sreg_reg[1115]  ( .D(c[1116]), .CLK(clk), .RST(rst), .Q(sreg[1115]) );
  DFF \sreg_reg[1114]  ( .D(c[1115]), .CLK(clk), .RST(rst), .Q(sreg[1114]) );
  DFF \sreg_reg[1113]  ( .D(c[1114]), .CLK(clk), .RST(rst), .Q(sreg[1113]) );
  DFF \sreg_reg[1112]  ( .D(c[1113]), .CLK(clk), .RST(rst), .Q(sreg[1112]) );
  DFF \sreg_reg[1111]  ( .D(c[1112]), .CLK(clk), .RST(rst), .Q(sreg[1111]) );
  DFF \sreg_reg[1110]  ( .D(c[1111]), .CLK(clk), .RST(rst), .Q(sreg[1110]) );
  DFF \sreg_reg[1109]  ( .D(c[1110]), .CLK(clk), .RST(rst), .Q(sreg[1109]) );
  DFF \sreg_reg[1108]  ( .D(c[1109]), .CLK(clk), .RST(rst), .Q(sreg[1108]) );
  DFF \sreg_reg[1107]  ( .D(c[1108]), .CLK(clk), .RST(rst), .Q(sreg[1107]) );
  DFF \sreg_reg[1106]  ( .D(c[1107]), .CLK(clk), .RST(rst), .Q(sreg[1106]) );
  DFF \sreg_reg[1105]  ( .D(c[1106]), .CLK(clk), .RST(rst), .Q(sreg[1105]) );
  DFF \sreg_reg[1104]  ( .D(c[1105]), .CLK(clk), .RST(rst), .Q(sreg[1104]) );
  DFF \sreg_reg[1103]  ( .D(c[1104]), .CLK(clk), .RST(rst), .Q(sreg[1103]) );
  DFF \sreg_reg[1102]  ( .D(c[1103]), .CLK(clk), .RST(rst), .Q(sreg[1102]) );
  DFF \sreg_reg[1101]  ( .D(c[1102]), .CLK(clk), .RST(rst), .Q(sreg[1101]) );
  DFF \sreg_reg[1100]  ( .D(c[1101]), .CLK(clk), .RST(rst), .Q(sreg[1100]) );
  DFF \sreg_reg[1099]  ( .D(c[1100]), .CLK(clk), .RST(rst), .Q(sreg[1099]) );
  DFF \sreg_reg[1098]  ( .D(c[1099]), .CLK(clk), .RST(rst), .Q(sreg[1098]) );
  DFF \sreg_reg[1097]  ( .D(c[1098]), .CLK(clk), .RST(rst), .Q(sreg[1097]) );
  DFF \sreg_reg[1096]  ( .D(c[1097]), .CLK(clk), .RST(rst), .Q(sreg[1096]) );
  DFF \sreg_reg[1095]  ( .D(c[1096]), .CLK(clk), .RST(rst), .Q(sreg[1095]) );
  DFF \sreg_reg[1094]  ( .D(c[1095]), .CLK(clk), .RST(rst), .Q(sreg[1094]) );
  DFF \sreg_reg[1093]  ( .D(c[1094]), .CLK(clk), .RST(rst), .Q(sreg[1093]) );
  DFF \sreg_reg[1092]  ( .D(c[1093]), .CLK(clk), .RST(rst), .Q(sreg[1092]) );
  DFF \sreg_reg[1091]  ( .D(c[1092]), .CLK(clk), .RST(rst), .Q(sreg[1091]) );
  DFF \sreg_reg[1090]  ( .D(c[1091]), .CLK(clk), .RST(rst), .Q(sreg[1090]) );
  DFF \sreg_reg[1089]  ( .D(c[1090]), .CLK(clk), .RST(rst), .Q(sreg[1089]) );
  DFF \sreg_reg[1088]  ( .D(c[1089]), .CLK(clk), .RST(rst), .Q(sreg[1088]) );
  DFF \sreg_reg[1087]  ( .D(c[1088]), .CLK(clk), .RST(rst), .Q(sreg[1087]) );
  DFF \sreg_reg[1086]  ( .D(c[1087]), .CLK(clk), .RST(rst), .Q(sreg[1086]) );
  DFF \sreg_reg[1085]  ( .D(c[1086]), .CLK(clk), .RST(rst), .Q(sreg[1085]) );
  DFF \sreg_reg[1084]  ( .D(c[1085]), .CLK(clk), .RST(rst), .Q(sreg[1084]) );
  DFF \sreg_reg[1083]  ( .D(c[1084]), .CLK(clk), .RST(rst), .Q(sreg[1083]) );
  DFF \sreg_reg[1082]  ( .D(c[1083]), .CLK(clk), .RST(rst), .Q(sreg[1082]) );
  DFF \sreg_reg[1081]  ( .D(c[1082]), .CLK(clk), .RST(rst), .Q(sreg[1081]) );
  DFF \sreg_reg[1080]  ( .D(c[1081]), .CLK(clk), .RST(rst), .Q(sreg[1080]) );
  DFF \sreg_reg[1079]  ( .D(c[1080]), .CLK(clk), .RST(rst), .Q(sreg[1079]) );
  DFF \sreg_reg[1078]  ( .D(c[1079]), .CLK(clk), .RST(rst), .Q(sreg[1078]) );
  DFF \sreg_reg[1077]  ( .D(c[1078]), .CLK(clk), .RST(rst), .Q(sreg[1077]) );
  DFF \sreg_reg[1076]  ( .D(c[1077]), .CLK(clk), .RST(rst), .Q(sreg[1076]) );
  DFF \sreg_reg[1075]  ( .D(c[1076]), .CLK(clk), .RST(rst), .Q(sreg[1075]) );
  DFF \sreg_reg[1074]  ( .D(c[1075]), .CLK(clk), .RST(rst), .Q(sreg[1074]) );
  DFF \sreg_reg[1073]  ( .D(c[1074]), .CLK(clk), .RST(rst), .Q(sreg[1073]) );
  DFF \sreg_reg[1072]  ( .D(c[1073]), .CLK(clk), .RST(rst), .Q(sreg[1072]) );
  DFF \sreg_reg[1071]  ( .D(c[1072]), .CLK(clk), .RST(rst), .Q(sreg[1071]) );
  DFF \sreg_reg[1070]  ( .D(c[1071]), .CLK(clk), .RST(rst), .Q(sreg[1070]) );
  DFF \sreg_reg[1069]  ( .D(c[1070]), .CLK(clk), .RST(rst), .Q(sreg[1069]) );
  DFF \sreg_reg[1068]  ( .D(c[1069]), .CLK(clk), .RST(rst), .Q(sreg[1068]) );
  DFF \sreg_reg[1067]  ( .D(c[1068]), .CLK(clk), .RST(rst), .Q(sreg[1067]) );
  DFF \sreg_reg[1066]  ( .D(c[1067]), .CLK(clk), .RST(rst), .Q(sreg[1066]) );
  DFF \sreg_reg[1065]  ( .D(c[1066]), .CLK(clk), .RST(rst), .Q(sreg[1065]) );
  DFF \sreg_reg[1064]  ( .D(c[1065]), .CLK(clk), .RST(rst), .Q(sreg[1064]) );
  DFF \sreg_reg[1063]  ( .D(c[1064]), .CLK(clk), .RST(rst), .Q(sreg[1063]) );
  DFF \sreg_reg[1062]  ( .D(c[1063]), .CLK(clk), .RST(rst), .Q(sreg[1062]) );
  DFF \sreg_reg[1061]  ( .D(c[1062]), .CLK(clk), .RST(rst), .Q(sreg[1061]) );
  DFF \sreg_reg[1060]  ( .D(c[1061]), .CLK(clk), .RST(rst), .Q(sreg[1060]) );
  DFF \sreg_reg[1059]  ( .D(c[1060]), .CLK(clk), .RST(rst), .Q(sreg[1059]) );
  DFF \sreg_reg[1058]  ( .D(c[1059]), .CLK(clk), .RST(rst), .Q(sreg[1058]) );
  DFF \sreg_reg[1057]  ( .D(c[1058]), .CLK(clk), .RST(rst), .Q(sreg[1057]) );
  DFF \sreg_reg[1056]  ( .D(c[1057]), .CLK(clk), .RST(rst), .Q(sreg[1056]) );
  DFF \sreg_reg[1055]  ( .D(c[1056]), .CLK(clk), .RST(rst), .Q(sreg[1055]) );
  DFF \sreg_reg[1054]  ( .D(c[1055]), .CLK(clk), .RST(rst), .Q(sreg[1054]) );
  DFF \sreg_reg[1053]  ( .D(c[1054]), .CLK(clk), .RST(rst), .Q(sreg[1053]) );
  DFF \sreg_reg[1052]  ( .D(c[1053]), .CLK(clk), .RST(rst), .Q(sreg[1052]) );
  DFF \sreg_reg[1051]  ( .D(c[1052]), .CLK(clk), .RST(rst), .Q(sreg[1051]) );
  DFF \sreg_reg[1050]  ( .D(c[1051]), .CLK(clk), .RST(rst), .Q(sreg[1050]) );
  DFF \sreg_reg[1049]  ( .D(c[1050]), .CLK(clk), .RST(rst), .Q(sreg[1049]) );
  DFF \sreg_reg[1048]  ( .D(c[1049]), .CLK(clk), .RST(rst), .Q(sreg[1048]) );
  DFF \sreg_reg[1047]  ( .D(c[1048]), .CLK(clk), .RST(rst), .Q(sreg[1047]) );
  DFF \sreg_reg[1046]  ( .D(c[1047]), .CLK(clk), .RST(rst), .Q(sreg[1046]) );
  DFF \sreg_reg[1045]  ( .D(c[1046]), .CLK(clk), .RST(rst), .Q(sreg[1045]) );
  DFF \sreg_reg[1044]  ( .D(c[1045]), .CLK(clk), .RST(rst), .Q(sreg[1044]) );
  DFF \sreg_reg[1043]  ( .D(c[1044]), .CLK(clk), .RST(rst), .Q(sreg[1043]) );
  DFF \sreg_reg[1042]  ( .D(c[1043]), .CLK(clk), .RST(rst), .Q(sreg[1042]) );
  DFF \sreg_reg[1041]  ( .D(c[1042]), .CLK(clk), .RST(rst), .Q(sreg[1041]) );
  DFF \sreg_reg[1040]  ( .D(c[1041]), .CLK(clk), .RST(rst), .Q(sreg[1040]) );
  DFF \sreg_reg[1039]  ( .D(c[1040]), .CLK(clk), .RST(rst), .Q(sreg[1039]) );
  DFF \sreg_reg[1038]  ( .D(c[1039]), .CLK(clk), .RST(rst), .Q(sreg[1038]) );
  DFF \sreg_reg[1037]  ( .D(c[1038]), .CLK(clk), .RST(rst), .Q(sreg[1037]) );
  DFF \sreg_reg[1036]  ( .D(c[1037]), .CLK(clk), .RST(rst), .Q(sreg[1036]) );
  DFF \sreg_reg[1035]  ( .D(c[1036]), .CLK(clk), .RST(rst), .Q(sreg[1035]) );
  DFF \sreg_reg[1034]  ( .D(c[1035]), .CLK(clk), .RST(rst), .Q(sreg[1034]) );
  DFF \sreg_reg[1033]  ( .D(c[1034]), .CLK(clk), .RST(rst), .Q(sreg[1033]) );
  DFF \sreg_reg[1032]  ( .D(c[1033]), .CLK(clk), .RST(rst), .Q(sreg[1032]) );
  DFF \sreg_reg[1031]  ( .D(c[1032]), .CLK(clk), .RST(rst), .Q(sreg[1031]) );
  DFF \sreg_reg[1030]  ( .D(c[1031]), .CLK(clk), .RST(rst), .Q(sreg[1030]) );
  DFF \sreg_reg[1029]  ( .D(c[1030]), .CLK(clk), .RST(rst), .Q(sreg[1029]) );
  DFF \sreg_reg[1028]  ( .D(c[1029]), .CLK(clk), .RST(rst), .Q(sreg[1028]) );
  DFF \sreg_reg[1027]  ( .D(c[1028]), .CLK(clk), .RST(rst), .Q(sreg[1027]) );
  DFF \sreg_reg[1026]  ( .D(c[1027]), .CLK(clk), .RST(rst), .Q(sreg[1026]) );
  DFF \sreg_reg[1025]  ( .D(c[1026]), .CLK(clk), .RST(rst), .Q(sreg[1025]) );
  DFF \sreg_reg[1024]  ( .D(c[1025]), .CLK(clk), .RST(rst), .Q(sreg[1024]) );
  DFF \sreg_reg[1023]  ( .D(c[1024]), .CLK(clk), .RST(rst), .Q(sreg[1023]) );
  DFF \sreg_reg[1022]  ( .D(c[1023]), .CLK(clk), .RST(rst), .Q(c[1022]) );
  DFF \sreg_reg[1021]  ( .D(c[1022]), .CLK(clk), .RST(rst), .Q(c[1021]) );
  DFF \sreg_reg[1020]  ( .D(c[1021]), .CLK(clk), .RST(rst), .Q(c[1020]) );
  DFF \sreg_reg[1019]  ( .D(c[1020]), .CLK(clk), .RST(rst), .Q(c[1019]) );
  DFF \sreg_reg[1018]  ( .D(c[1019]), .CLK(clk), .RST(rst), .Q(c[1018]) );
  DFF \sreg_reg[1017]  ( .D(c[1018]), .CLK(clk), .RST(rst), .Q(c[1017]) );
  DFF \sreg_reg[1016]  ( .D(c[1017]), .CLK(clk), .RST(rst), .Q(c[1016]) );
  DFF \sreg_reg[1015]  ( .D(c[1016]), .CLK(clk), .RST(rst), .Q(c[1015]) );
  DFF \sreg_reg[1014]  ( .D(c[1015]), .CLK(clk), .RST(rst), .Q(c[1014]) );
  DFF \sreg_reg[1013]  ( .D(c[1014]), .CLK(clk), .RST(rst), .Q(c[1013]) );
  DFF \sreg_reg[1012]  ( .D(c[1013]), .CLK(clk), .RST(rst), .Q(c[1012]) );
  DFF \sreg_reg[1011]  ( .D(c[1012]), .CLK(clk), .RST(rst), .Q(c[1011]) );
  DFF \sreg_reg[1010]  ( .D(c[1011]), .CLK(clk), .RST(rst), .Q(c[1010]) );
  DFF \sreg_reg[1009]  ( .D(c[1010]), .CLK(clk), .RST(rst), .Q(c[1009]) );
  DFF \sreg_reg[1008]  ( .D(c[1009]), .CLK(clk), .RST(rst), .Q(c[1008]) );
  DFF \sreg_reg[1007]  ( .D(c[1008]), .CLK(clk), .RST(rst), .Q(c[1007]) );
  DFF \sreg_reg[1006]  ( .D(c[1007]), .CLK(clk), .RST(rst), .Q(c[1006]) );
  DFF \sreg_reg[1005]  ( .D(c[1006]), .CLK(clk), .RST(rst), .Q(c[1005]) );
  DFF \sreg_reg[1004]  ( .D(c[1005]), .CLK(clk), .RST(rst), .Q(c[1004]) );
  DFF \sreg_reg[1003]  ( .D(c[1004]), .CLK(clk), .RST(rst), .Q(c[1003]) );
  DFF \sreg_reg[1002]  ( .D(c[1003]), .CLK(clk), .RST(rst), .Q(c[1002]) );
  DFF \sreg_reg[1001]  ( .D(c[1002]), .CLK(clk), .RST(rst), .Q(c[1001]) );
  DFF \sreg_reg[1000]  ( .D(c[1001]), .CLK(clk), .RST(rst), .Q(c[1000]) );
  DFF \sreg_reg[999]  ( .D(c[1000]), .CLK(clk), .RST(rst), .Q(c[999]) );
  DFF \sreg_reg[998]  ( .D(c[999]), .CLK(clk), .RST(rst), .Q(c[998]) );
  DFF \sreg_reg[997]  ( .D(c[998]), .CLK(clk), .RST(rst), .Q(c[997]) );
  DFF \sreg_reg[996]  ( .D(c[997]), .CLK(clk), .RST(rst), .Q(c[996]) );
  DFF \sreg_reg[995]  ( .D(c[996]), .CLK(clk), .RST(rst), .Q(c[995]) );
  DFF \sreg_reg[994]  ( .D(c[995]), .CLK(clk), .RST(rst), .Q(c[994]) );
  DFF \sreg_reg[993]  ( .D(c[994]), .CLK(clk), .RST(rst), .Q(c[993]) );
  DFF \sreg_reg[992]  ( .D(c[993]), .CLK(clk), .RST(rst), .Q(c[992]) );
  DFF \sreg_reg[991]  ( .D(c[992]), .CLK(clk), .RST(rst), .Q(c[991]) );
  DFF \sreg_reg[990]  ( .D(c[991]), .CLK(clk), .RST(rst), .Q(c[990]) );
  DFF \sreg_reg[989]  ( .D(c[990]), .CLK(clk), .RST(rst), .Q(c[989]) );
  DFF \sreg_reg[988]  ( .D(c[989]), .CLK(clk), .RST(rst), .Q(c[988]) );
  DFF \sreg_reg[987]  ( .D(c[988]), .CLK(clk), .RST(rst), .Q(c[987]) );
  DFF \sreg_reg[986]  ( .D(c[987]), .CLK(clk), .RST(rst), .Q(c[986]) );
  DFF \sreg_reg[985]  ( .D(c[986]), .CLK(clk), .RST(rst), .Q(c[985]) );
  DFF \sreg_reg[984]  ( .D(c[985]), .CLK(clk), .RST(rst), .Q(c[984]) );
  DFF \sreg_reg[983]  ( .D(c[984]), .CLK(clk), .RST(rst), .Q(c[983]) );
  DFF \sreg_reg[982]  ( .D(c[983]), .CLK(clk), .RST(rst), .Q(c[982]) );
  DFF \sreg_reg[981]  ( .D(c[982]), .CLK(clk), .RST(rst), .Q(c[981]) );
  DFF \sreg_reg[980]  ( .D(c[981]), .CLK(clk), .RST(rst), .Q(c[980]) );
  DFF \sreg_reg[979]  ( .D(c[980]), .CLK(clk), .RST(rst), .Q(c[979]) );
  DFF \sreg_reg[978]  ( .D(c[979]), .CLK(clk), .RST(rst), .Q(c[978]) );
  DFF \sreg_reg[977]  ( .D(c[978]), .CLK(clk), .RST(rst), .Q(c[977]) );
  DFF \sreg_reg[976]  ( .D(c[977]), .CLK(clk), .RST(rst), .Q(c[976]) );
  DFF \sreg_reg[975]  ( .D(c[976]), .CLK(clk), .RST(rst), .Q(c[975]) );
  DFF \sreg_reg[974]  ( .D(c[975]), .CLK(clk), .RST(rst), .Q(c[974]) );
  DFF \sreg_reg[973]  ( .D(c[974]), .CLK(clk), .RST(rst), .Q(c[973]) );
  DFF \sreg_reg[972]  ( .D(c[973]), .CLK(clk), .RST(rst), .Q(c[972]) );
  DFF \sreg_reg[971]  ( .D(c[972]), .CLK(clk), .RST(rst), .Q(c[971]) );
  DFF \sreg_reg[970]  ( .D(c[971]), .CLK(clk), .RST(rst), .Q(c[970]) );
  DFF \sreg_reg[969]  ( .D(c[970]), .CLK(clk), .RST(rst), .Q(c[969]) );
  DFF \sreg_reg[968]  ( .D(c[969]), .CLK(clk), .RST(rst), .Q(c[968]) );
  DFF \sreg_reg[967]  ( .D(c[968]), .CLK(clk), .RST(rst), .Q(c[967]) );
  DFF \sreg_reg[966]  ( .D(c[967]), .CLK(clk), .RST(rst), .Q(c[966]) );
  DFF \sreg_reg[965]  ( .D(c[966]), .CLK(clk), .RST(rst), .Q(c[965]) );
  DFF \sreg_reg[964]  ( .D(c[965]), .CLK(clk), .RST(rst), .Q(c[964]) );
  DFF \sreg_reg[963]  ( .D(c[964]), .CLK(clk), .RST(rst), .Q(c[963]) );
  DFF \sreg_reg[962]  ( .D(c[963]), .CLK(clk), .RST(rst), .Q(c[962]) );
  DFF \sreg_reg[961]  ( .D(c[962]), .CLK(clk), .RST(rst), .Q(c[961]) );
  DFF \sreg_reg[960]  ( .D(c[961]), .CLK(clk), .RST(rst), .Q(c[960]) );
  DFF \sreg_reg[959]  ( .D(c[960]), .CLK(clk), .RST(rst), .Q(c[959]) );
  DFF \sreg_reg[958]  ( .D(c[959]), .CLK(clk), .RST(rst), .Q(c[958]) );
  DFF \sreg_reg[957]  ( .D(c[958]), .CLK(clk), .RST(rst), .Q(c[957]) );
  DFF \sreg_reg[956]  ( .D(c[957]), .CLK(clk), .RST(rst), .Q(c[956]) );
  DFF \sreg_reg[955]  ( .D(c[956]), .CLK(clk), .RST(rst), .Q(c[955]) );
  DFF \sreg_reg[954]  ( .D(c[955]), .CLK(clk), .RST(rst), .Q(c[954]) );
  DFF \sreg_reg[953]  ( .D(c[954]), .CLK(clk), .RST(rst), .Q(c[953]) );
  DFF \sreg_reg[952]  ( .D(c[953]), .CLK(clk), .RST(rst), .Q(c[952]) );
  DFF \sreg_reg[951]  ( .D(c[952]), .CLK(clk), .RST(rst), .Q(c[951]) );
  DFF \sreg_reg[950]  ( .D(c[951]), .CLK(clk), .RST(rst), .Q(c[950]) );
  DFF \sreg_reg[949]  ( .D(c[950]), .CLK(clk), .RST(rst), .Q(c[949]) );
  DFF \sreg_reg[948]  ( .D(c[949]), .CLK(clk), .RST(rst), .Q(c[948]) );
  DFF \sreg_reg[947]  ( .D(c[948]), .CLK(clk), .RST(rst), .Q(c[947]) );
  DFF \sreg_reg[946]  ( .D(c[947]), .CLK(clk), .RST(rst), .Q(c[946]) );
  DFF \sreg_reg[945]  ( .D(c[946]), .CLK(clk), .RST(rst), .Q(c[945]) );
  DFF \sreg_reg[944]  ( .D(c[945]), .CLK(clk), .RST(rst), .Q(c[944]) );
  DFF \sreg_reg[943]  ( .D(c[944]), .CLK(clk), .RST(rst), .Q(c[943]) );
  DFF \sreg_reg[942]  ( .D(c[943]), .CLK(clk), .RST(rst), .Q(c[942]) );
  DFF \sreg_reg[941]  ( .D(c[942]), .CLK(clk), .RST(rst), .Q(c[941]) );
  DFF \sreg_reg[940]  ( .D(c[941]), .CLK(clk), .RST(rst), .Q(c[940]) );
  DFF \sreg_reg[939]  ( .D(c[940]), .CLK(clk), .RST(rst), .Q(c[939]) );
  DFF \sreg_reg[938]  ( .D(c[939]), .CLK(clk), .RST(rst), .Q(c[938]) );
  DFF \sreg_reg[937]  ( .D(c[938]), .CLK(clk), .RST(rst), .Q(c[937]) );
  DFF \sreg_reg[936]  ( .D(c[937]), .CLK(clk), .RST(rst), .Q(c[936]) );
  DFF \sreg_reg[935]  ( .D(c[936]), .CLK(clk), .RST(rst), .Q(c[935]) );
  DFF \sreg_reg[934]  ( .D(c[935]), .CLK(clk), .RST(rst), .Q(c[934]) );
  DFF \sreg_reg[933]  ( .D(c[934]), .CLK(clk), .RST(rst), .Q(c[933]) );
  DFF \sreg_reg[932]  ( .D(c[933]), .CLK(clk), .RST(rst), .Q(c[932]) );
  DFF \sreg_reg[931]  ( .D(c[932]), .CLK(clk), .RST(rst), .Q(c[931]) );
  DFF \sreg_reg[930]  ( .D(c[931]), .CLK(clk), .RST(rst), .Q(c[930]) );
  DFF \sreg_reg[929]  ( .D(c[930]), .CLK(clk), .RST(rst), .Q(c[929]) );
  DFF \sreg_reg[928]  ( .D(c[929]), .CLK(clk), .RST(rst), .Q(c[928]) );
  DFF \sreg_reg[927]  ( .D(c[928]), .CLK(clk), .RST(rst), .Q(c[927]) );
  DFF \sreg_reg[926]  ( .D(c[927]), .CLK(clk), .RST(rst), .Q(c[926]) );
  DFF \sreg_reg[925]  ( .D(c[926]), .CLK(clk), .RST(rst), .Q(c[925]) );
  DFF \sreg_reg[924]  ( .D(c[925]), .CLK(clk), .RST(rst), .Q(c[924]) );
  DFF \sreg_reg[923]  ( .D(c[924]), .CLK(clk), .RST(rst), .Q(c[923]) );
  DFF \sreg_reg[922]  ( .D(c[923]), .CLK(clk), .RST(rst), .Q(c[922]) );
  DFF \sreg_reg[921]  ( .D(c[922]), .CLK(clk), .RST(rst), .Q(c[921]) );
  DFF \sreg_reg[920]  ( .D(c[921]), .CLK(clk), .RST(rst), .Q(c[920]) );
  DFF \sreg_reg[919]  ( .D(c[920]), .CLK(clk), .RST(rst), .Q(c[919]) );
  DFF \sreg_reg[918]  ( .D(c[919]), .CLK(clk), .RST(rst), .Q(c[918]) );
  DFF \sreg_reg[917]  ( .D(c[918]), .CLK(clk), .RST(rst), .Q(c[917]) );
  DFF \sreg_reg[916]  ( .D(c[917]), .CLK(clk), .RST(rst), .Q(c[916]) );
  DFF \sreg_reg[915]  ( .D(c[916]), .CLK(clk), .RST(rst), .Q(c[915]) );
  DFF \sreg_reg[914]  ( .D(c[915]), .CLK(clk), .RST(rst), .Q(c[914]) );
  DFF \sreg_reg[913]  ( .D(c[914]), .CLK(clk), .RST(rst), .Q(c[913]) );
  DFF \sreg_reg[912]  ( .D(c[913]), .CLK(clk), .RST(rst), .Q(c[912]) );
  DFF \sreg_reg[911]  ( .D(c[912]), .CLK(clk), .RST(rst), .Q(c[911]) );
  DFF \sreg_reg[910]  ( .D(c[911]), .CLK(clk), .RST(rst), .Q(c[910]) );
  DFF \sreg_reg[909]  ( .D(c[910]), .CLK(clk), .RST(rst), .Q(c[909]) );
  DFF \sreg_reg[908]  ( .D(c[909]), .CLK(clk), .RST(rst), .Q(c[908]) );
  DFF \sreg_reg[907]  ( .D(c[908]), .CLK(clk), .RST(rst), .Q(c[907]) );
  DFF \sreg_reg[906]  ( .D(c[907]), .CLK(clk), .RST(rst), .Q(c[906]) );
  DFF \sreg_reg[905]  ( .D(c[906]), .CLK(clk), .RST(rst), .Q(c[905]) );
  DFF \sreg_reg[904]  ( .D(c[905]), .CLK(clk), .RST(rst), .Q(c[904]) );
  DFF \sreg_reg[903]  ( .D(c[904]), .CLK(clk), .RST(rst), .Q(c[903]) );
  DFF \sreg_reg[902]  ( .D(c[903]), .CLK(clk), .RST(rst), .Q(c[902]) );
  DFF \sreg_reg[901]  ( .D(c[902]), .CLK(clk), .RST(rst), .Q(c[901]) );
  DFF \sreg_reg[900]  ( .D(c[901]), .CLK(clk), .RST(rst), .Q(c[900]) );
  DFF \sreg_reg[899]  ( .D(c[900]), .CLK(clk), .RST(rst), .Q(c[899]) );
  DFF \sreg_reg[898]  ( .D(c[899]), .CLK(clk), .RST(rst), .Q(c[898]) );
  DFF \sreg_reg[897]  ( .D(c[898]), .CLK(clk), .RST(rst), .Q(c[897]) );
  DFF \sreg_reg[896]  ( .D(c[897]), .CLK(clk), .RST(rst), .Q(c[896]) );
  DFF \sreg_reg[895]  ( .D(c[896]), .CLK(clk), .RST(rst), .Q(c[895]) );
  DFF \sreg_reg[894]  ( .D(c[895]), .CLK(clk), .RST(rst), .Q(c[894]) );
  DFF \sreg_reg[893]  ( .D(c[894]), .CLK(clk), .RST(rst), .Q(c[893]) );
  DFF \sreg_reg[892]  ( .D(c[893]), .CLK(clk), .RST(rst), .Q(c[892]) );
  DFF \sreg_reg[891]  ( .D(c[892]), .CLK(clk), .RST(rst), .Q(c[891]) );
  DFF \sreg_reg[890]  ( .D(c[891]), .CLK(clk), .RST(rst), .Q(c[890]) );
  DFF \sreg_reg[889]  ( .D(c[890]), .CLK(clk), .RST(rst), .Q(c[889]) );
  DFF \sreg_reg[888]  ( .D(c[889]), .CLK(clk), .RST(rst), .Q(c[888]) );
  DFF \sreg_reg[887]  ( .D(c[888]), .CLK(clk), .RST(rst), .Q(c[887]) );
  DFF \sreg_reg[886]  ( .D(c[887]), .CLK(clk), .RST(rst), .Q(c[886]) );
  DFF \sreg_reg[885]  ( .D(c[886]), .CLK(clk), .RST(rst), .Q(c[885]) );
  DFF \sreg_reg[884]  ( .D(c[885]), .CLK(clk), .RST(rst), .Q(c[884]) );
  DFF \sreg_reg[883]  ( .D(c[884]), .CLK(clk), .RST(rst), .Q(c[883]) );
  DFF \sreg_reg[882]  ( .D(c[883]), .CLK(clk), .RST(rst), .Q(c[882]) );
  DFF \sreg_reg[881]  ( .D(c[882]), .CLK(clk), .RST(rst), .Q(c[881]) );
  DFF \sreg_reg[880]  ( .D(c[881]), .CLK(clk), .RST(rst), .Q(c[880]) );
  DFF \sreg_reg[879]  ( .D(c[880]), .CLK(clk), .RST(rst), .Q(c[879]) );
  DFF \sreg_reg[878]  ( .D(c[879]), .CLK(clk), .RST(rst), .Q(c[878]) );
  DFF \sreg_reg[877]  ( .D(c[878]), .CLK(clk), .RST(rst), .Q(c[877]) );
  DFF \sreg_reg[876]  ( .D(c[877]), .CLK(clk), .RST(rst), .Q(c[876]) );
  DFF \sreg_reg[875]  ( .D(c[876]), .CLK(clk), .RST(rst), .Q(c[875]) );
  DFF \sreg_reg[874]  ( .D(c[875]), .CLK(clk), .RST(rst), .Q(c[874]) );
  DFF \sreg_reg[873]  ( .D(c[874]), .CLK(clk), .RST(rst), .Q(c[873]) );
  DFF \sreg_reg[872]  ( .D(c[873]), .CLK(clk), .RST(rst), .Q(c[872]) );
  DFF \sreg_reg[871]  ( .D(c[872]), .CLK(clk), .RST(rst), .Q(c[871]) );
  DFF \sreg_reg[870]  ( .D(c[871]), .CLK(clk), .RST(rst), .Q(c[870]) );
  DFF \sreg_reg[869]  ( .D(c[870]), .CLK(clk), .RST(rst), .Q(c[869]) );
  DFF \sreg_reg[868]  ( .D(c[869]), .CLK(clk), .RST(rst), .Q(c[868]) );
  DFF \sreg_reg[867]  ( .D(c[868]), .CLK(clk), .RST(rst), .Q(c[867]) );
  DFF \sreg_reg[866]  ( .D(c[867]), .CLK(clk), .RST(rst), .Q(c[866]) );
  DFF \sreg_reg[865]  ( .D(c[866]), .CLK(clk), .RST(rst), .Q(c[865]) );
  DFF \sreg_reg[864]  ( .D(c[865]), .CLK(clk), .RST(rst), .Q(c[864]) );
  DFF \sreg_reg[863]  ( .D(c[864]), .CLK(clk), .RST(rst), .Q(c[863]) );
  DFF \sreg_reg[862]  ( .D(c[863]), .CLK(clk), .RST(rst), .Q(c[862]) );
  DFF \sreg_reg[861]  ( .D(c[862]), .CLK(clk), .RST(rst), .Q(c[861]) );
  DFF \sreg_reg[860]  ( .D(c[861]), .CLK(clk), .RST(rst), .Q(c[860]) );
  DFF \sreg_reg[859]  ( .D(c[860]), .CLK(clk), .RST(rst), .Q(c[859]) );
  DFF \sreg_reg[858]  ( .D(c[859]), .CLK(clk), .RST(rst), .Q(c[858]) );
  DFF \sreg_reg[857]  ( .D(c[858]), .CLK(clk), .RST(rst), .Q(c[857]) );
  DFF \sreg_reg[856]  ( .D(c[857]), .CLK(clk), .RST(rst), .Q(c[856]) );
  DFF \sreg_reg[855]  ( .D(c[856]), .CLK(clk), .RST(rst), .Q(c[855]) );
  DFF \sreg_reg[854]  ( .D(c[855]), .CLK(clk), .RST(rst), .Q(c[854]) );
  DFF \sreg_reg[853]  ( .D(c[854]), .CLK(clk), .RST(rst), .Q(c[853]) );
  DFF \sreg_reg[852]  ( .D(c[853]), .CLK(clk), .RST(rst), .Q(c[852]) );
  DFF \sreg_reg[851]  ( .D(c[852]), .CLK(clk), .RST(rst), .Q(c[851]) );
  DFF \sreg_reg[850]  ( .D(c[851]), .CLK(clk), .RST(rst), .Q(c[850]) );
  DFF \sreg_reg[849]  ( .D(c[850]), .CLK(clk), .RST(rst), .Q(c[849]) );
  DFF \sreg_reg[848]  ( .D(c[849]), .CLK(clk), .RST(rst), .Q(c[848]) );
  DFF \sreg_reg[847]  ( .D(c[848]), .CLK(clk), .RST(rst), .Q(c[847]) );
  DFF \sreg_reg[846]  ( .D(c[847]), .CLK(clk), .RST(rst), .Q(c[846]) );
  DFF \sreg_reg[845]  ( .D(c[846]), .CLK(clk), .RST(rst), .Q(c[845]) );
  DFF \sreg_reg[844]  ( .D(c[845]), .CLK(clk), .RST(rst), .Q(c[844]) );
  DFF \sreg_reg[843]  ( .D(c[844]), .CLK(clk), .RST(rst), .Q(c[843]) );
  DFF \sreg_reg[842]  ( .D(c[843]), .CLK(clk), .RST(rst), .Q(c[842]) );
  DFF \sreg_reg[841]  ( .D(c[842]), .CLK(clk), .RST(rst), .Q(c[841]) );
  DFF \sreg_reg[840]  ( .D(c[841]), .CLK(clk), .RST(rst), .Q(c[840]) );
  DFF \sreg_reg[839]  ( .D(c[840]), .CLK(clk), .RST(rst), .Q(c[839]) );
  DFF \sreg_reg[838]  ( .D(c[839]), .CLK(clk), .RST(rst), .Q(c[838]) );
  DFF \sreg_reg[837]  ( .D(c[838]), .CLK(clk), .RST(rst), .Q(c[837]) );
  DFF \sreg_reg[836]  ( .D(c[837]), .CLK(clk), .RST(rst), .Q(c[836]) );
  DFF \sreg_reg[835]  ( .D(c[836]), .CLK(clk), .RST(rst), .Q(c[835]) );
  DFF \sreg_reg[834]  ( .D(c[835]), .CLK(clk), .RST(rst), .Q(c[834]) );
  DFF \sreg_reg[833]  ( .D(c[834]), .CLK(clk), .RST(rst), .Q(c[833]) );
  DFF \sreg_reg[832]  ( .D(c[833]), .CLK(clk), .RST(rst), .Q(c[832]) );
  DFF \sreg_reg[831]  ( .D(c[832]), .CLK(clk), .RST(rst), .Q(c[831]) );
  DFF \sreg_reg[830]  ( .D(c[831]), .CLK(clk), .RST(rst), .Q(c[830]) );
  DFF \sreg_reg[829]  ( .D(c[830]), .CLK(clk), .RST(rst), .Q(c[829]) );
  DFF \sreg_reg[828]  ( .D(c[829]), .CLK(clk), .RST(rst), .Q(c[828]) );
  DFF \sreg_reg[827]  ( .D(c[828]), .CLK(clk), .RST(rst), .Q(c[827]) );
  DFF \sreg_reg[826]  ( .D(c[827]), .CLK(clk), .RST(rst), .Q(c[826]) );
  DFF \sreg_reg[825]  ( .D(c[826]), .CLK(clk), .RST(rst), .Q(c[825]) );
  DFF \sreg_reg[824]  ( .D(c[825]), .CLK(clk), .RST(rst), .Q(c[824]) );
  DFF \sreg_reg[823]  ( .D(c[824]), .CLK(clk), .RST(rst), .Q(c[823]) );
  DFF \sreg_reg[822]  ( .D(c[823]), .CLK(clk), .RST(rst), .Q(c[822]) );
  DFF \sreg_reg[821]  ( .D(c[822]), .CLK(clk), .RST(rst), .Q(c[821]) );
  DFF \sreg_reg[820]  ( .D(c[821]), .CLK(clk), .RST(rst), .Q(c[820]) );
  DFF \sreg_reg[819]  ( .D(c[820]), .CLK(clk), .RST(rst), .Q(c[819]) );
  DFF \sreg_reg[818]  ( .D(c[819]), .CLK(clk), .RST(rst), .Q(c[818]) );
  DFF \sreg_reg[817]  ( .D(c[818]), .CLK(clk), .RST(rst), .Q(c[817]) );
  DFF \sreg_reg[816]  ( .D(c[817]), .CLK(clk), .RST(rst), .Q(c[816]) );
  DFF \sreg_reg[815]  ( .D(c[816]), .CLK(clk), .RST(rst), .Q(c[815]) );
  DFF \sreg_reg[814]  ( .D(c[815]), .CLK(clk), .RST(rst), .Q(c[814]) );
  DFF \sreg_reg[813]  ( .D(c[814]), .CLK(clk), .RST(rst), .Q(c[813]) );
  DFF \sreg_reg[812]  ( .D(c[813]), .CLK(clk), .RST(rst), .Q(c[812]) );
  DFF \sreg_reg[811]  ( .D(c[812]), .CLK(clk), .RST(rst), .Q(c[811]) );
  DFF \sreg_reg[810]  ( .D(c[811]), .CLK(clk), .RST(rst), .Q(c[810]) );
  DFF \sreg_reg[809]  ( .D(c[810]), .CLK(clk), .RST(rst), .Q(c[809]) );
  DFF \sreg_reg[808]  ( .D(c[809]), .CLK(clk), .RST(rst), .Q(c[808]) );
  DFF \sreg_reg[807]  ( .D(c[808]), .CLK(clk), .RST(rst), .Q(c[807]) );
  DFF \sreg_reg[806]  ( .D(c[807]), .CLK(clk), .RST(rst), .Q(c[806]) );
  DFF \sreg_reg[805]  ( .D(c[806]), .CLK(clk), .RST(rst), .Q(c[805]) );
  DFF \sreg_reg[804]  ( .D(c[805]), .CLK(clk), .RST(rst), .Q(c[804]) );
  DFF \sreg_reg[803]  ( .D(c[804]), .CLK(clk), .RST(rst), .Q(c[803]) );
  DFF \sreg_reg[802]  ( .D(c[803]), .CLK(clk), .RST(rst), .Q(c[802]) );
  DFF \sreg_reg[801]  ( .D(c[802]), .CLK(clk), .RST(rst), .Q(c[801]) );
  DFF \sreg_reg[800]  ( .D(c[801]), .CLK(clk), .RST(rst), .Q(c[800]) );
  DFF \sreg_reg[799]  ( .D(c[800]), .CLK(clk), .RST(rst), .Q(c[799]) );
  DFF \sreg_reg[798]  ( .D(c[799]), .CLK(clk), .RST(rst), .Q(c[798]) );
  DFF \sreg_reg[797]  ( .D(c[798]), .CLK(clk), .RST(rst), .Q(c[797]) );
  DFF \sreg_reg[796]  ( .D(c[797]), .CLK(clk), .RST(rst), .Q(c[796]) );
  DFF \sreg_reg[795]  ( .D(c[796]), .CLK(clk), .RST(rst), .Q(c[795]) );
  DFF \sreg_reg[794]  ( .D(c[795]), .CLK(clk), .RST(rst), .Q(c[794]) );
  DFF \sreg_reg[793]  ( .D(c[794]), .CLK(clk), .RST(rst), .Q(c[793]) );
  DFF \sreg_reg[792]  ( .D(c[793]), .CLK(clk), .RST(rst), .Q(c[792]) );
  DFF \sreg_reg[791]  ( .D(c[792]), .CLK(clk), .RST(rst), .Q(c[791]) );
  DFF \sreg_reg[790]  ( .D(c[791]), .CLK(clk), .RST(rst), .Q(c[790]) );
  DFF \sreg_reg[789]  ( .D(c[790]), .CLK(clk), .RST(rst), .Q(c[789]) );
  DFF \sreg_reg[788]  ( .D(c[789]), .CLK(clk), .RST(rst), .Q(c[788]) );
  DFF \sreg_reg[787]  ( .D(c[788]), .CLK(clk), .RST(rst), .Q(c[787]) );
  DFF \sreg_reg[786]  ( .D(c[787]), .CLK(clk), .RST(rst), .Q(c[786]) );
  DFF \sreg_reg[785]  ( .D(c[786]), .CLK(clk), .RST(rst), .Q(c[785]) );
  DFF \sreg_reg[784]  ( .D(c[785]), .CLK(clk), .RST(rst), .Q(c[784]) );
  DFF \sreg_reg[783]  ( .D(c[784]), .CLK(clk), .RST(rst), .Q(c[783]) );
  DFF \sreg_reg[782]  ( .D(c[783]), .CLK(clk), .RST(rst), .Q(c[782]) );
  DFF \sreg_reg[781]  ( .D(c[782]), .CLK(clk), .RST(rst), .Q(c[781]) );
  DFF \sreg_reg[780]  ( .D(c[781]), .CLK(clk), .RST(rst), .Q(c[780]) );
  DFF \sreg_reg[779]  ( .D(c[780]), .CLK(clk), .RST(rst), .Q(c[779]) );
  DFF \sreg_reg[778]  ( .D(c[779]), .CLK(clk), .RST(rst), .Q(c[778]) );
  DFF \sreg_reg[777]  ( .D(c[778]), .CLK(clk), .RST(rst), .Q(c[777]) );
  DFF \sreg_reg[776]  ( .D(c[777]), .CLK(clk), .RST(rst), .Q(c[776]) );
  DFF \sreg_reg[775]  ( .D(c[776]), .CLK(clk), .RST(rst), .Q(c[775]) );
  DFF \sreg_reg[774]  ( .D(c[775]), .CLK(clk), .RST(rst), .Q(c[774]) );
  DFF \sreg_reg[773]  ( .D(c[774]), .CLK(clk), .RST(rst), .Q(c[773]) );
  DFF \sreg_reg[772]  ( .D(c[773]), .CLK(clk), .RST(rst), .Q(c[772]) );
  DFF \sreg_reg[771]  ( .D(c[772]), .CLK(clk), .RST(rst), .Q(c[771]) );
  DFF \sreg_reg[770]  ( .D(c[771]), .CLK(clk), .RST(rst), .Q(c[770]) );
  DFF \sreg_reg[769]  ( .D(c[770]), .CLK(clk), .RST(rst), .Q(c[769]) );
  DFF \sreg_reg[768]  ( .D(c[769]), .CLK(clk), .RST(rst), .Q(c[768]) );
  DFF \sreg_reg[767]  ( .D(c[768]), .CLK(clk), .RST(rst), .Q(c[767]) );
  DFF \sreg_reg[766]  ( .D(c[767]), .CLK(clk), .RST(rst), .Q(c[766]) );
  DFF \sreg_reg[765]  ( .D(c[766]), .CLK(clk), .RST(rst), .Q(c[765]) );
  DFF \sreg_reg[764]  ( .D(c[765]), .CLK(clk), .RST(rst), .Q(c[764]) );
  DFF \sreg_reg[763]  ( .D(c[764]), .CLK(clk), .RST(rst), .Q(c[763]) );
  DFF \sreg_reg[762]  ( .D(c[763]), .CLK(clk), .RST(rst), .Q(c[762]) );
  DFF \sreg_reg[761]  ( .D(c[762]), .CLK(clk), .RST(rst), .Q(c[761]) );
  DFF \sreg_reg[760]  ( .D(c[761]), .CLK(clk), .RST(rst), .Q(c[760]) );
  DFF \sreg_reg[759]  ( .D(c[760]), .CLK(clk), .RST(rst), .Q(c[759]) );
  DFF \sreg_reg[758]  ( .D(c[759]), .CLK(clk), .RST(rst), .Q(c[758]) );
  DFF \sreg_reg[757]  ( .D(c[758]), .CLK(clk), .RST(rst), .Q(c[757]) );
  DFF \sreg_reg[756]  ( .D(c[757]), .CLK(clk), .RST(rst), .Q(c[756]) );
  DFF \sreg_reg[755]  ( .D(c[756]), .CLK(clk), .RST(rst), .Q(c[755]) );
  DFF \sreg_reg[754]  ( .D(c[755]), .CLK(clk), .RST(rst), .Q(c[754]) );
  DFF \sreg_reg[753]  ( .D(c[754]), .CLK(clk), .RST(rst), .Q(c[753]) );
  DFF \sreg_reg[752]  ( .D(c[753]), .CLK(clk), .RST(rst), .Q(c[752]) );
  DFF \sreg_reg[751]  ( .D(c[752]), .CLK(clk), .RST(rst), .Q(c[751]) );
  DFF \sreg_reg[750]  ( .D(c[751]), .CLK(clk), .RST(rst), .Q(c[750]) );
  DFF \sreg_reg[749]  ( .D(c[750]), .CLK(clk), .RST(rst), .Q(c[749]) );
  DFF \sreg_reg[748]  ( .D(c[749]), .CLK(clk), .RST(rst), .Q(c[748]) );
  DFF \sreg_reg[747]  ( .D(c[748]), .CLK(clk), .RST(rst), .Q(c[747]) );
  DFF \sreg_reg[746]  ( .D(c[747]), .CLK(clk), .RST(rst), .Q(c[746]) );
  DFF \sreg_reg[745]  ( .D(c[746]), .CLK(clk), .RST(rst), .Q(c[745]) );
  DFF \sreg_reg[744]  ( .D(c[745]), .CLK(clk), .RST(rst), .Q(c[744]) );
  DFF \sreg_reg[743]  ( .D(c[744]), .CLK(clk), .RST(rst), .Q(c[743]) );
  DFF \sreg_reg[742]  ( .D(c[743]), .CLK(clk), .RST(rst), .Q(c[742]) );
  DFF \sreg_reg[741]  ( .D(c[742]), .CLK(clk), .RST(rst), .Q(c[741]) );
  DFF \sreg_reg[740]  ( .D(c[741]), .CLK(clk), .RST(rst), .Q(c[740]) );
  DFF \sreg_reg[739]  ( .D(c[740]), .CLK(clk), .RST(rst), .Q(c[739]) );
  DFF \sreg_reg[738]  ( .D(c[739]), .CLK(clk), .RST(rst), .Q(c[738]) );
  DFF \sreg_reg[737]  ( .D(c[738]), .CLK(clk), .RST(rst), .Q(c[737]) );
  DFF \sreg_reg[736]  ( .D(c[737]), .CLK(clk), .RST(rst), .Q(c[736]) );
  DFF \sreg_reg[735]  ( .D(c[736]), .CLK(clk), .RST(rst), .Q(c[735]) );
  DFF \sreg_reg[734]  ( .D(c[735]), .CLK(clk), .RST(rst), .Q(c[734]) );
  DFF \sreg_reg[733]  ( .D(c[734]), .CLK(clk), .RST(rst), .Q(c[733]) );
  DFF \sreg_reg[732]  ( .D(c[733]), .CLK(clk), .RST(rst), .Q(c[732]) );
  DFF \sreg_reg[731]  ( .D(c[732]), .CLK(clk), .RST(rst), .Q(c[731]) );
  DFF \sreg_reg[730]  ( .D(c[731]), .CLK(clk), .RST(rst), .Q(c[730]) );
  DFF \sreg_reg[729]  ( .D(c[730]), .CLK(clk), .RST(rst), .Q(c[729]) );
  DFF \sreg_reg[728]  ( .D(c[729]), .CLK(clk), .RST(rst), .Q(c[728]) );
  DFF \sreg_reg[727]  ( .D(c[728]), .CLK(clk), .RST(rst), .Q(c[727]) );
  DFF \sreg_reg[726]  ( .D(c[727]), .CLK(clk), .RST(rst), .Q(c[726]) );
  DFF \sreg_reg[725]  ( .D(c[726]), .CLK(clk), .RST(rst), .Q(c[725]) );
  DFF \sreg_reg[724]  ( .D(c[725]), .CLK(clk), .RST(rst), .Q(c[724]) );
  DFF \sreg_reg[723]  ( .D(c[724]), .CLK(clk), .RST(rst), .Q(c[723]) );
  DFF \sreg_reg[722]  ( .D(c[723]), .CLK(clk), .RST(rst), .Q(c[722]) );
  DFF \sreg_reg[721]  ( .D(c[722]), .CLK(clk), .RST(rst), .Q(c[721]) );
  DFF \sreg_reg[720]  ( .D(c[721]), .CLK(clk), .RST(rst), .Q(c[720]) );
  DFF \sreg_reg[719]  ( .D(c[720]), .CLK(clk), .RST(rst), .Q(c[719]) );
  DFF \sreg_reg[718]  ( .D(c[719]), .CLK(clk), .RST(rst), .Q(c[718]) );
  DFF \sreg_reg[717]  ( .D(c[718]), .CLK(clk), .RST(rst), .Q(c[717]) );
  DFF \sreg_reg[716]  ( .D(c[717]), .CLK(clk), .RST(rst), .Q(c[716]) );
  DFF \sreg_reg[715]  ( .D(c[716]), .CLK(clk), .RST(rst), .Q(c[715]) );
  DFF \sreg_reg[714]  ( .D(c[715]), .CLK(clk), .RST(rst), .Q(c[714]) );
  DFF \sreg_reg[713]  ( .D(c[714]), .CLK(clk), .RST(rst), .Q(c[713]) );
  DFF \sreg_reg[712]  ( .D(c[713]), .CLK(clk), .RST(rst), .Q(c[712]) );
  DFF \sreg_reg[711]  ( .D(c[712]), .CLK(clk), .RST(rst), .Q(c[711]) );
  DFF \sreg_reg[710]  ( .D(c[711]), .CLK(clk), .RST(rst), .Q(c[710]) );
  DFF \sreg_reg[709]  ( .D(c[710]), .CLK(clk), .RST(rst), .Q(c[709]) );
  DFF \sreg_reg[708]  ( .D(c[709]), .CLK(clk), .RST(rst), .Q(c[708]) );
  DFF \sreg_reg[707]  ( .D(c[708]), .CLK(clk), .RST(rst), .Q(c[707]) );
  DFF \sreg_reg[706]  ( .D(c[707]), .CLK(clk), .RST(rst), .Q(c[706]) );
  DFF \sreg_reg[705]  ( .D(c[706]), .CLK(clk), .RST(rst), .Q(c[705]) );
  DFF \sreg_reg[704]  ( .D(c[705]), .CLK(clk), .RST(rst), .Q(c[704]) );
  DFF \sreg_reg[703]  ( .D(c[704]), .CLK(clk), .RST(rst), .Q(c[703]) );
  DFF \sreg_reg[702]  ( .D(c[703]), .CLK(clk), .RST(rst), .Q(c[702]) );
  DFF \sreg_reg[701]  ( .D(c[702]), .CLK(clk), .RST(rst), .Q(c[701]) );
  DFF \sreg_reg[700]  ( .D(c[701]), .CLK(clk), .RST(rst), .Q(c[700]) );
  DFF \sreg_reg[699]  ( .D(c[700]), .CLK(clk), .RST(rst), .Q(c[699]) );
  DFF \sreg_reg[698]  ( .D(c[699]), .CLK(clk), .RST(rst), .Q(c[698]) );
  DFF \sreg_reg[697]  ( .D(c[698]), .CLK(clk), .RST(rst), .Q(c[697]) );
  DFF \sreg_reg[696]  ( .D(c[697]), .CLK(clk), .RST(rst), .Q(c[696]) );
  DFF \sreg_reg[695]  ( .D(c[696]), .CLK(clk), .RST(rst), .Q(c[695]) );
  DFF \sreg_reg[694]  ( .D(c[695]), .CLK(clk), .RST(rst), .Q(c[694]) );
  DFF \sreg_reg[693]  ( .D(c[694]), .CLK(clk), .RST(rst), .Q(c[693]) );
  DFF \sreg_reg[692]  ( .D(c[693]), .CLK(clk), .RST(rst), .Q(c[692]) );
  DFF \sreg_reg[691]  ( .D(c[692]), .CLK(clk), .RST(rst), .Q(c[691]) );
  DFF \sreg_reg[690]  ( .D(c[691]), .CLK(clk), .RST(rst), .Q(c[690]) );
  DFF \sreg_reg[689]  ( .D(c[690]), .CLK(clk), .RST(rst), .Q(c[689]) );
  DFF \sreg_reg[688]  ( .D(c[689]), .CLK(clk), .RST(rst), .Q(c[688]) );
  DFF \sreg_reg[687]  ( .D(c[688]), .CLK(clk), .RST(rst), .Q(c[687]) );
  DFF \sreg_reg[686]  ( .D(c[687]), .CLK(clk), .RST(rst), .Q(c[686]) );
  DFF \sreg_reg[685]  ( .D(c[686]), .CLK(clk), .RST(rst), .Q(c[685]) );
  DFF \sreg_reg[684]  ( .D(c[685]), .CLK(clk), .RST(rst), .Q(c[684]) );
  DFF \sreg_reg[683]  ( .D(c[684]), .CLK(clk), .RST(rst), .Q(c[683]) );
  DFF \sreg_reg[682]  ( .D(c[683]), .CLK(clk), .RST(rst), .Q(c[682]) );
  DFF \sreg_reg[681]  ( .D(c[682]), .CLK(clk), .RST(rst), .Q(c[681]) );
  DFF \sreg_reg[680]  ( .D(c[681]), .CLK(clk), .RST(rst), .Q(c[680]) );
  DFF \sreg_reg[679]  ( .D(c[680]), .CLK(clk), .RST(rst), .Q(c[679]) );
  DFF \sreg_reg[678]  ( .D(c[679]), .CLK(clk), .RST(rst), .Q(c[678]) );
  DFF \sreg_reg[677]  ( .D(c[678]), .CLK(clk), .RST(rst), .Q(c[677]) );
  DFF \sreg_reg[676]  ( .D(c[677]), .CLK(clk), .RST(rst), .Q(c[676]) );
  DFF \sreg_reg[675]  ( .D(c[676]), .CLK(clk), .RST(rst), .Q(c[675]) );
  DFF \sreg_reg[674]  ( .D(c[675]), .CLK(clk), .RST(rst), .Q(c[674]) );
  DFF \sreg_reg[673]  ( .D(c[674]), .CLK(clk), .RST(rst), .Q(c[673]) );
  DFF \sreg_reg[672]  ( .D(c[673]), .CLK(clk), .RST(rst), .Q(c[672]) );
  DFF \sreg_reg[671]  ( .D(c[672]), .CLK(clk), .RST(rst), .Q(c[671]) );
  DFF \sreg_reg[670]  ( .D(c[671]), .CLK(clk), .RST(rst), .Q(c[670]) );
  DFF \sreg_reg[669]  ( .D(c[670]), .CLK(clk), .RST(rst), .Q(c[669]) );
  DFF \sreg_reg[668]  ( .D(c[669]), .CLK(clk), .RST(rst), .Q(c[668]) );
  DFF \sreg_reg[667]  ( .D(c[668]), .CLK(clk), .RST(rst), .Q(c[667]) );
  DFF \sreg_reg[666]  ( .D(c[667]), .CLK(clk), .RST(rst), .Q(c[666]) );
  DFF \sreg_reg[665]  ( .D(c[666]), .CLK(clk), .RST(rst), .Q(c[665]) );
  DFF \sreg_reg[664]  ( .D(c[665]), .CLK(clk), .RST(rst), .Q(c[664]) );
  DFF \sreg_reg[663]  ( .D(c[664]), .CLK(clk), .RST(rst), .Q(c[663]) );
  DFF \sreg_reg[662]  ( .D(c[663]), .CLK(clk), .RST(rst), .Q(c[662]) );
  DFF \sreg_reg[661]  ( .D(c[662]), .CLK(clk), .RST(rst), .Q(c[661]) );
  DFF \sreg_reg[660]  ( .D(c[661]), .CLK(clk), .RST(rst), .Q(c[660]) );
  DFF \sreg_reg[659]  ( .D(c[660]), .CLK(clk), .RST(rst), .Q(c[659]) );
  DFF \sreg_reg[658]  ( .D(c[659]), .CLK(clk), .RST(rst), .Q(c[658]) );
  DFF \sreg_reg[657]  ( .D(c[658]), .CLK(clk), .RST(rst), .Q(c[657]) );
  DFF \sreg_reg[656]  ( .D(c[657]), .CLK(clk), .RST(rst), .Q(c[656]) );
  DFF \sreg_reg[655]  ( .D(c[656]), .CLK(clk), .RST(rst), .Q(c[655]) );
  DFF \sreg_reg[654]  ( .D(c[655]), .CLK(clk), .RST(rst), .Q(c[654]) );
  DFF \sreg_reg[653]  ( .D(c[654]), .CLK(clk), .RST(rst), .Q(c[653]) );
  DFF \sreg_reg[652]  ( .D(c[653]), .CLK(clk), .RST(rst), .Q(c[652]) );
  DFF \sreg_reg[651]  ( .D(c[652]), .CLK(clk), .RST(rst), .Q(c[651]) );
  DFF \sreg_reg[650]  ( .D(c[651]), .CLK(clk), .RST(rst), .Q(c[650]) );
  DFF \sreg_reg[649]  ( .D(c[650]), .CLK(clk), .RST(rst), .Q(c[649]) );
  DFF \sreg_reg[648]  ( .D(c[649]), .CLK(clk), .RST(rst), .Q(c[648]) );
  DFF \sreg_reg[647]  ( .D(c[648]), .CLK(clk), .RST(rst), .Q(c[647]) );
  DFF \sreg_reg[646]  ( .D(c[647]), .CLK(clk), .RST(rst), .Q(c[646]) );
  DFF \sreg_reg[645]  ( .D(c[646]), .CLK(clk), .RST(rst), .Q(c[645]) );
  DFF \sreg_reg[644]  ( .D(c[645]), .CLK(clk), .RST(rst), .Q(c[644]) );
  DFF \sreg_reg[643]  ( .D(c[644]), .CLK(clk), .RST(rst), .Q(c[643]) );
  DFF \sreg_reg[642]  ( .D(c[643]), .CLK(clk), .RST(rst), .Q(c[642]) );
  DFF \sreg_reg[641]  ( .D(c[642]), .CLK(clk), .RST(rst), .Q(c[641]) );
  DFF \sreg_reg[640]  ( .D(c[641]), .CLK(clk), .RST(rst), .Q(c[640]) );
  DFF \sreg_reg[639]  ( .D(c[640]), .CLK(clk), .RST(rst), .Q(c[639]) );
  DFF \sreg_reg[638]  ( .D(c[639]), .CLK(clk), .RST(rst), .Q(c[638]) );
  DFF \sreg_reg[637]  ( .D(c[638]), .CLK(clk), .RST(rst), .Q(c[637]) );
  DFF \sreg_reg[636]  ( .D(c[637]), .CLK(clk), .RST(rst), .Q(c[636]) );
  DFF \sreg_reg[635]  ( .D(c[636]), .CLK(clk), .RST(rst), .Q(c[635]) );
  DFF \sreg_reg[634]  ( .D(c[635]), .CLK(clk), .RST(rst), .Q(c[634]) );
  DFF \sreg_reg[633]  ( .D(c[634]), .CLK(clk), .RST(rst), .Q(c[633]) );
  DFF \sreg_reg[632]  ( .D(c[633]), .CLK(clk), .RST(rst), .Q(c[632]) );
  DFF \sreg_reg[631]  ( .D(c[632]), .CLK(clk), .RST(rst), .Q(c[631]) );
  DFF \sreg_reg[630]  ( .D(c[631]), .CLK(clk), .RST(rst), .Q(c[630]) );
  DFF \sreg_reg[629]  ( .D(c[630]), .CLK(clk), .RST(rst), .Q(c[629]) );
  DFF \sreg_reg[628]  ( .D(c[629]), .CLK(clk), .RST(rst), .Q(c[628]) );
  DFF \sreg_reg[627]  ( .D(c[628]), .CLK(clk), .RST(rst), .Q(c[627]) );
  DFF \sreg_reg[626]  ( .D(c[627]), .CLK(clk), .RST(rst), .Q(c[626]) );
  DFF \sreg_reg[625]  ( .D(c[626]), .CLK(clk), .RST(rst), .Q(c[625]) );
  DFF \sreg_reg[624]  ( .D(c[625]), .CLK(clk), .RST(rst), .Q(c[624]) );
  DFF \sreg_reg[623]  ( .D(c[624]), .CLK(clk), .RST(rst), .Q(c[623]) );
  DFF \sreg_reg[622]  ( .D(c[623]), .CLK(clk), .RST(rst), .Q(c[622]) );
  DFF \sreg_reg[621]  ( .D(c[622]), .CLK(clk), .RST(rst), .Q(c[621]) );
  DFF \sreg_reg[620]  ( .D(c[621]), .CLK(clk), .RST(rst), .Q(c[620]) );
  DFF \sreg_reg[619]  ( .D(c[620]), .CLK(clk), .RST(rst), .Q(c[619]) );
  DFF \sreg_reg[618]  ( .D(c[619]), .CLK(clk), .RST(rst), .Q(c[618]) );
  DFF \sreg_reg[617]  ( .D(c[618]), .CLK(clk), .RST(rst), .Q(c[617]) );
  DFF \sreg_reg[616]  ( .D(c[617]), .CLK(clk), .RST(rst), .Q(c[616]) );
  DFF \sreg_reg[615]  ( .D(c[616]), .CLK(clk), .RST(rst), .Q(c[615]) );
  DFF \sreg_reg[614]  ( .D(c[615]), .CLK(clk), .RST(rst), .Q(c[614]) );
  DFF \sreg_reg[613]  ( .D(c[614]), .CLK(clk), .RST(rst), .Q(c[613]) );
  DFF \sreg_reg[612]  ( .D(c[613]), .CLK(clk), .RST(rst), .Q(c[612]) );
  DFF \sreg_reg[611]  ( .D(c[612]), .CLK(clk), .RST(rst), .Q(c[611]) );
  DFF \sreg_reg[610]  ( .D(c[611]), .CLK(clk), .RST(rst), .Q(c[610]) );
  DFF \sreg_reg[609]  ( .D(c[610]), .CLK(clk), .RST(rst), .Q(c[609]) );
  DFF \sreg_reg[608]  ( .D(c[609]), .CLK(clk), .RST(rst), .Q(c[608]) );
  DFF \sreg_reg[607]  ( .D(c[608]), .CLK(clk), .RST(rst), .Q(c[607]) );
  DFF \sreg_reg[606]  ( .D(c[607]), .CLK(clk), .RST(rst), .Q(c[606]) );
  DFF \sreg_reg[605]  ( .D(c[606]), .CLK(clk), .RST(rst), .Q(c[605]) );
  DFF \sreg_reg[604]  ( .D(c[605]), .CLK(clk), .RST(rst), .Q(c[604]) );
  DFF \sreg_reg[603]  ( .D(c[604]), .CLK(clk), .RST(rst), .Q(c[603]) );
  DFF \sreg_reg[602]  ( .D(c[603]), .CLK(clk), .RST(rst), .Q(c[602]) );
  DFF \sreg_reg[601]  ( .D(c[602]), .CLK(clk), .RST(rst), .Q(c[601]) );
  DFF \sreg_reg[600]  ( .D(c[601]), .CLK(clk), .RST(rst), .Q(c[600]) );
  DFF \sreg_reg[599]  ( .D(c[600]), .CLK(clk), .RST(rst), .Q(c[599]) );
  DFF \sreg_reg[598]  ( .D(c[599]), .CLK(clk), .RST(rst), .Q(c[598]) );
  DFF \sreg_reg[597]  ( .D(c[598]), .CLK(clk), .RST(rst), .Q(c[597]) );
  DFF \sreg_reg[596]  ( .D(c[597]), .CLK(clk), .RST(rst), .Q(c[596]) );
  DFF \sreg_reg[595]  ( .D(c[596]), .CLK(clk), .RST(rst), .Q(c[595]) );
  DFF \sreg_reg[594]  ( .D(c[595]), .CLK(clk), .RST(rst), .Q(c[594]) );
  DFF \sreg_reg[593]  ( .D(c[594]), .CLK(clk), .RST(rst), .Q(c[593]) );
  DFF \sreg_reg[592]  ( .D(c[593]), .CLK(clk), .RST(rst), .Q(c[592]) );
  DFF \sreg_reg[591]  ( .D(c[592]), .CLK(clk), .RST(rst), .Q(c[591]) );
  DFF \sreg_reg[590]  ( .D(c[591]), .CLK(clk), .RST(rst), .Q(c[590]) );
  DFF \sreg_reg[589]  ( .D(c[590]), .CLK(clk), .RST(rst), .Q(c[589]) );
  DFF \sreg_reg[588]  ( .D(c[589]), .CLK(clk), .RST(rst), .Q(c[588]) );
  DFF \sreg_reg[587]  ( .D(c[588]), .CLK(clk), .RST(rst), .Q(c[587]) );
  DFF \sreg_reg[586]  ( .D(c[587]), .CLK(clk), .RST(rst), .Q(c[586]) );
  DFF \sreg_reg[585]  ( .D(c[586]), .CLK(clk), .RST(rst), .Q(c[585]) );
  DFF \sreg_reg[584]  ( .D(c[585]), .CLK(clk), .RST(rst), .Q(c[584]) );
  DFF \sreg_reg[583]  ( .D(c[584]), .CLK(clk), .RST(rst), .Q(c[583]) );
  DFF \sreg_reg[582]  ( .D(c[583]), .CLK(clk), .RST(rst), .Q(c[582]) );
  DFF \sreg_reg[581]  ( .D(c[582]), .CLK(clk), .RST(rst), .Q(c[581]) );
  DFF \sreg_reg[580]  ( .D(c[581]), .CLK(clk), .RST(rst), .Q(c[580]) );
  DFF \sreg_reg[579]  ( .D(c[580]), .CLK(clk), .RST(rst), .Q(c[579]) );
  DFF \sreg_reg[578]  ( .D(c[579]), .CLK(clk), .RST(rst), .Q(c[578]) );
  DFF \sreg_reg[577]  ( .D(c[578]), .CLK(clk), .RST(rst), .Q(c[577]) );
  DFF \sreg_reg[576]  ( .D(c[577]), .CLK(clk), .RST(rst), .Q(c[576]) );
  DFF \sreg_reg[575]  ( .D(c[576]), .CLK(clk), .RST(rst), .Q(c[575]) );
  DFF \sreg_reg[574]  ( .D(c[575]), .CLK(clk), .RST(rst), .Q(c[574]) );
  DFF \sreg_reg[573]  ( .D(c[574]), .CLK(clk), .RST(rst), .Q(c[573]) );
  DFF \sreg_reg[572]  ( .D(c[573]), .CLK(clk), .RST(rst), .Q(c[572]) );
  DFF \sreg_reg[571]  ( .D(c[572]), .CLK(clk), .RST(rst), .Q(c[571]) );
  DFF \sreg_reg[570]  ( .D(c[571]), .CLK(clk), .RST(rst), .Q(c[570]) );
  DFF \sreg_reg[569]  ( .D(c[570]), .CLK(clk), .RST(rst), .Q(c[569]) );
  DFF \sreg_reg[568]  ( .D(c[569]), .CLK(clk), .RST(rst), .Q(c[568]) );
  DFF \sreg_reg[567]  ( .D(c[568]), .CLK(clk), .RST(rst), .Q(c[567]) );
  DFF \sreg_reg[566]  ( .D(c[567]), .CLK(clk), .RST(rst), .Q(c[566]) );
  DFF \sreg_reg[565]  ( .D(c[566]), .CLK(clk), .RST(rst), .Q(c[565]) );
  DFF \sreg_reg[564]  ( .D(c[565]), .CLK(clk), .RST(rst), .Q(c[564]) );
  DFF \sreg_reg[563]  ( .D(c[564]), .CLK(clk), .RST(rst), .Q(c[563]) );
  DFF \sreg_reg[562]  ( .D(c[563]), .CLK(clk), .RST(rst), .Q(c[562]) );
  DFF \sreg_reg[561]  ( .D(c[562]), .CLK(clk), .RST(rst), .Q(c[561]) );
  DFF \sreg_reg[560]  ( .D(c[561]), .CLK(clk), .RST(rst), .Q(c[560]) );
  DFF \sreg_reg[559]  ( .D(c[560]), .CLK(clk), .RST(rst), .Q(c[559]) );
  DFF \sreg_reg[558]  ( .D(c[559]), .CLK(clk), .RST(rst), .Q(c[558]) );
  DFF \sreg_reg[557]  ( .D(c[558]), .CLK(clk), .RST(rst), .Q(c[557]) );
  DFF \sreg_reg[556]  ( .D(c[557]), .CLK(clk), .RST(rst), .Q(c[556]) );
  DFF \sreg_reg[555]  ( .D(c[556]), .CLK(clk), .RST(rst), .Q(c[555]) );
  DFF \sreg_reg[554]  ( .D(c[555]), .CLK(clk), .RST(rst), .Q(c[554]) );
  DFF \sreg_reg[553]  ( .D(c[554]), .CLK(clk), .RST(rst), .Q(c[553]) );
  DFF \sreg_reg[552]  ( .D(c[553]), .CLK(clk), .RST(rst), .Q(c[552]) );
  DFF \sreg_reg[551]  ( .D(c[552]), .CLK(clk), .RST(rst), .Q(c[551]) );
  DFF \sreg_reg[550]  ( .D(c[551]), .CLK(clk), .RST(rst), .Q(c[550]) );
  DFF \sreg_reg[549]  ( .D(c[550]), .CLK(clk), .RST(rst), .Q(c[549]) );
  DFF \sreg_reg[548]  ( .D(c[549]), .CLK(clk), .RST(rst), .Q(c[548]) );
  DFF \sreg_reg[547]  ( .D(c[548]), .CLK(clk), .RST(rst), .Q(c[547]) );
  DFF \sreg_reg[546]  ( .D(c[547]), .CLK(clk), .RST(rst), .Q(c[546]) );
  DFF \sreg_reg[545]  ( .D(c[546]), .CLK(clk), .RST(rst), .Q(c[545]) );
  DFF \sreg_reg[544]  ( .D(c[545]), .CLK(clk), .RST(rst), .Q(c[544]) );
  DFF \sreg_reg[543]  ( .D(c[544]), .CLK(clk), .RST(rst), .Q(c[543]) );
  DFF \sreg_reg[542]  ( .D(c[543]), .CLK(clk), .RST(rst), .Q(c[542]) );
  DFF \sreg_reg[541]  ( .D(c[542]), .CLK(clk), .RST(rst), .Q(c[541]) );
  DFF \sreg_reg[540]  ( .D(c[541]), .CLK(clk), .RST(rst), .Q(c[540]) );
  DFF \sreg_reg[539]  ( .D(c[540]), .CLK(clk), .RST(rst), .Q(c[539]) );
  DFF \sreg_reg[538]  ( .D(c[539]), .CLK(clk), .RST(rst), .Q(c[538]) );
  DFF \sreg_reg[537]  ( .D(c[538]), .CLK(clk), .RST(rst), .Q(c[537]) );
  DFF \sreg_reg[536]  ( .D(c[537]), .CLK(clk), .RST(rst), .Q(c[536]) );
  DFF \sreg_reg[535]  ( .D(c[536]), .CLK(clk), .RST(rst), .Q(c[535]) );
  DFF \sreg_reg[534]  ( .D(c[535]), .CLK(clk), .RST(rst), .Q(c[534]) );
  DFF \sreg_reg[533]  ( .D(c[534]), .CLK(clk), .RST(rst), .Q(c[533]) );
  DFF \sreg_reg[532]  ( .D(c[533]), .CLK(clk), .RST(rst), .Q(c[532]) );
  DFF \sreg_reg[531]  ( .D(c[532]), .CLK(clk), .RST(rst), .Q(c[531]) );
  DFF \sreg_reg[530]  ( .D(c[531]), .CLK(clk), .RST(rst), .Q(c[530]) );
  DFF \sreg_reg[529]  ( .D(c[530]), .CLK(clk), .RST(rst), .Q(c[529]) );
  DFF \sreg_reg[528]  ( .D(c[529]), .CLK(clk), .RST(rst), .Q(c[528]) );
  DFF \sreg_reg[527]  ( .D(c[528]), .CLK(clk), .RST(rst), .Q(c[527]) );
  DFF \sreg_reg[526]  ( .D(c[527]), .CLK(clk), .RST(rst), .Q(c[526]) );
  DFF \sreg_reg[525]  ( .D(c[526]), .CLK(clk), .RST(rst), .Q(c[525]) );
  DFF \sreg_reg[524]  ( .D(c[525]), .CLK(clk), .RST(rst), .Q(c[524]) );
  DFF \sreg_reg[523]  ( .D(c[524]), .CLK(clk), .RST(rst), .Q(c[523]) );
  DFF \sreg_reg[522]  ( .D(c[523]), .CLK(clk), .RST(rst), .Q(c[522]) );
  DFF \sreg_reg[521]  ( .D(c[522]), .CLK(clk), .RST(rst), .Q(c[521]) );
  DFF \sreg_reg[520]  ( .D(c[521]), .CLK(clk), .RST(rst), .Q(c[520]) );
  DFF \sreg_reg[519]  ( .D(c[520]), .CLK(clk), .RST(rst), .Q(c[519]) );
  DFF \sreg_reg[518]  ( .D(c[519]), .CLK(clk), .RST(rst), .Q(c[518]) );
  DFF \sreg_reg[517]  ( .D(c[518]), .CLK(clk), .RST(rst), .Q(c[517]) );
  DFF \sreg_reg[516]  ( .D(c[517]), .CLK(clk), .RST(rst), .Q(c[516]) );
  DFF \sreg_reg[515]  ( .D(c[516]), .CLK(clk), .RST(rst), .Q(c[515]) );
  DFF \sreg_reg[514]  ( .D(c[515]), .CLK(clk), .RST(rst), .Q(c[514]) );
  DFF \sreg_reg[513]  ( .D(c[514]), .CLK(clk), .RST(rst), .Q(c[513]) );
  DFF \sreg_reg[512]  ( .D(c[513]), .CLK(clk), .RST(rst), .Q(c[512]) );
  DFF \sreg_reg[511]  ( .D(c[512]), .CLK(clk), .RST(rst), .Q(c[511]) );
  DFF \sreg_reg[510]  ( .D(c[511]), .CLK(clk), .RST(rst), .Q(c[510]) );
  DFF \sreg_reg[509]  ( .D(c[510]), .CLK(clk), .RST(rst), .Q(c[509]) );
  DFF \sreg_reg[508]  ( .D(c[509]), .CLK(clk), .RST(rst), .Q(c[508]) );
  DFF \sreg_reg[507]  ( .D(c[508]), .CLK(clk), .RST(rst), .Q(c[507]) );
  DFF \sreg_reg[506]  ( .D(c[507]), .CLK(clk), .RST(rst), .Q(c[506]) );
  DFF \sreg_reg[505]  ( .D(c[506]), .CLK(clk), .RST(rst), .Q(c[505]) );
  DFF \sreg_reg[504]  ( .D(c[505]), .CLK(clk), .RST(rst), .Q(c[504]) );
  DFF \sreg_reg[503]  ( .D(c[504]), .CLK(clk), .RST(rst), .Q(c[503]) );
  DFF \sreg_reg[502]  ( .D(c[503]), .CLK(clk), .RST(rst), .Q(c[502]) );
  DFF \sreg_reg[501]  ( .D(c[502]), .CLK(clk), .RST(rst), .Q(c[501]) );
  DFF \sreg_reg[500]  ( .D(c[501]), .CLK(clk), .RST(rst), .Q(c[500]) );
  DFF \sreg_reg[499]  ( .D(c[500]), .CLK(clk), .RST(rst), .Q(c[499]) );
  DFF \sreg_reg[498]  ( .D(c[499]), .CLK(clk), .RST(rst), .Q(c[498]) );
  DFF \sreg_reg[497]  ( .D(c[498]), .CLK(clk), .RST(rst), .Q(c[497]) );
  DFF \sreg_reg[496]  ( .D(c[497]), .CLK(clk), .RST(rst), .Q(c[496]) );
  DFF \sreg_reg[495]  ( .D(c[496]), .CLK(clk), .RST(rst), .Q(c[495]) );
  DFF \sreg_reg[494]  ( .D(c[495]), .CLK(clk), .RST(rst), .Q(c[494]) );
  DFF \sreg_reg[493]  ( .D(c[494]), .CLK(clk), .RST(rst), .Q(c[493]) );
  DFF \sreg_reg[492]  ( .D(c[493]), .CLK(clk), .RST(rst), .Q(c[492]) );
  DFF \sreg_reg[491]  ( .D(c[492]), .CLK(clk), .RST(rst), .Q(c[491]) );
  DFF \sreg_reg[490]  ( .D(c[491]), .CLK(clk), .RST(rst), .Q(c[490]) );
  DFF \sreg_reg[489]  ( .D(c[490]), .CLK(clk), .RST(rst), .Q(c[489]) );
  DFF \sreg_reg[488]  ( .D(c[489]), .CLK(clk), .RST(rst), .Q(c[488]) );
  DFF \sreg_reg[487]  ( .D(c[488]), .CLK(clk), .RST(rst), .Q(c[487]) );
  DFF \sreg_reg[486]  ( .D(c[487]), .CLK(clk), .RST(rst), .Q(c[486]) );
  DFF \sreg_reg[485]  ( .D(c[486]), .CLK(clk), .RST(rst), .Q(c[485]) );
  DFF \sreg_reg[484]  ( .D(c[485]), .CLK(clk), .RST(rst), .Q(c[484]) );
  DFF \sreg_reg[483]  ( .D(c[484]), .CLK(clk), .RST(rst), .Q(c[483]) );
  DFF \sreg_reg[482]  ( .D(c[483]), .CLK(clk), .RST(rst), .Q(c[482]) );
  DFF \sreg_reg[481]  ( .D(c[482]), .CLK(clk), .RST(rst), .Q(c[481]) );
  DFF \sreg_reg[480]  ( .D(c[481]), .CLK(clk), .RST(rst), .Q(c[480]) );
  DFF \sreg_reg[479]  ( .D(c[480]), .CLK(clk), .RST(rst), .Q(c[479]) );
  DFF \sreg_reg[478]  ( .D(c[479]), .CLK(clk), .RST(rst), .Q(c[478]) );
  DFF \sreg_reg[477]  ( .D(c[478]), .CLK(clk), .RST(rst), .Q(c[477]) );
  DFF \sreg_reg[476]  ( .D(c[477]), .CLK(clk), .RST(rst), .Q(c[476]) );
  DFF \sreg_reg[475]  ( .D(c[476]), .CLK(clk), .RST(rst), .Q(c[475]) );
  DFF \sreg_reg[474]  ( .D(c[475]), .CLK(clk), .RST(rst), .Q(c[474]) );
  DFF \sreg_reg[473]  ( .D(c[474]), .CLK(clk), .RST(rst), .Q(c[473]) );
  DFF \sreg_reg[472]  ( .D(c[473]), .CLK(clk), .RST(rst), .Q(c[472]) );
  DFF \sreg_reg[471]  ( .D(c[472]), .CLK(clk), .RST(rst), .Q(c[471]) );
  DFF \sreg_reg[470]  ( .D(c[471]), .CLK(clk), .RST(rst), .Q(c[470]) );
  DFF \sreg_reg[469]  ( .D(c[470]), .CLK(clk), .RST(rst), .Q(c[469]) );
  DFF \sreg_reg[468]  ( .D(c[469]), .CLK(clk), .RST(rst), .Q(c[468]) );
  DFF \sreg_reg[467]  ( .D(c[468]), .CLK(clk), .RST(rst), .Q(c[467]) );
  DFF \sreg_reg[466]  ( .D(c[467]), .CLK(clk), .RST(rst), .Q(c[466]) );
  DFF \sreg_reg[465]  ( .D(c[466]), .CLK(clk), .RST(rst), .Q(c[465]) );
  DFF \sreg_reg[464]  ( .D(c[465]), .CLK(clk), .RST(rst), .Q(c[464]) );
  DFF \sreg_reg[463]  ( .D(c[464]), .CLK(clk), .RST(rst), .Q(c[463]) );
  DFF \sreg_reg[462]  ( .D(c[463]), .CLK(clk), .RST(rst), .Q(c[462]) );
  DFF \sreg_reg[461]  ( .D(c[462]), .CLK(clk), .RST(rst), .Q(c[461]) );
  DFF \sreg_reg[460]  ( .D(c[461]), .CLK(clk), .RST(rst), .Q(c[460]) );
  DFF \sreg_reg[459]  ( .D(c[460]), .CLK(clk), .RST(rst), .Q(c[459]) );
  DFF \sreg_reg[458]  ( .D(c[459]), .CLK(clk), .RST(rst), .Q(c[458]) );
  DFF \sreg_reg[457]  ( .D(c[458]), .CLK(clk), .RST(rst), .Q(c[457]) );
  DFF \sreg_reg[456]  ( .D(c[457]), .CLK(clk), .RST(rst), .Q(c[456]) );
  DFF \sreg_reg[455]  ( .D(c[456]), .CLK(clk), .RST(rst), .Q(c[455]) );
  DFF \sreg_reg[454]  ( .D(c[455]), .CLK(clk), .RST(rst), .Q(c[454]) );
  DFF \sreg_reg[453]  ( .D(c[454]), .CLK(clk), .RST(rst), .Q(c[453]) );
  DFF \sreg_reg[452]  ( .D(c[453]), .CLK(clk), .RST(rst), .Q(c[452]) );
  DFF \sreg_reg[451]  ( .D(c[452]), .CLK(clk), .RST(rst), .Q(c[451]) );
  DFF \sreg_reg[450]  ( .D(c[451]), .CLK(clk), .RST(rst), .Q(c[450]) );
  DFF \sreg_reg[449]  ( .D(c[450]), .CLK(clk), .RST(rst), .Q(c[449]) );
  DFF \sreg_reg[448]  ( .D(c[449]), .CLK(clk), .RST(rst), .Q(c[448]) );
  DFF \sreg_reg[447]  ( .D(c[448]), .CLK(clk), .RST(rst), .Q(c[447]) );
  DFF \sreg_reg[446]  ( .D(c[447]), .CLK(clk), .RST(rst), .Q(c[446]) );
  DFF \sreg_reg[445]  ( .D(c[446]), .CLK(clk), .RST(rst), .Q(c[445]) );
  DFF \sreg_reg[444]  ( .D(c[445]), .CLK(clk), .RST(rst), .Q(c[444]) );
  DFF \sreg_reg[443]  ( .D(c[444]), .CLK(clk), .RST(rst), .Q(c[443]) );
  DFF \sreg_reg[442]  ( .D(c[443]), .CLK(clk), .RST(rst), .Q(c[442]) );
  DFF \sreg_reg[441]  ( .D(c[442]), .CLK(clk), .RST(rst), .Q(c[441]) );
  DFF \sreg_reg[440]  ( .D(c[441]), .CLK(clk), .RST(rst), .Q(c[440]) );
  DFF \sreg_reg[439]  ( .D(c[440]), .CLK(clk), .RST(rst), .Q(c[439]) );
  DFF \sreg_reg[438]  ( .D(c[439]), .CLK(clk), .RST(rst), .Q(c[438]) );
  DFF \sreg_reg[437]  ( .D(c[438]), .CLK(clk), .RST(rst), .Q(c[437]) );
  DFF \sreg_reg[436]  ( .D(c[437]), .CLK(clk), .RST(rst), .Q(c[436]) );
  DFF \sreg_reg[435]  ( .D(c[436]), .CLK(clk), .RST(rst), .Q(c[435]) );
  DFF \sreg_reg[434]  ( .D(c[435]), .CLK(clk), .RST(rst), .Q(c[434]) );
  DFF \sreg_reg[433]  ( .D(c[434]), .CLK(clk), .RST(rst), .Q(c[433]) );
  DFF \sreg_reg[432]  ( .D(c[433]), .CLK(clk), .RST(rst), .Q(c[432]) );
  DFF \sreg_reg[431]  ( .D(c[432]), .CLK(clk), .RST(rst), .Q(c[431]) );
  DFF \sreg_reg[430]  ( .D(c[431]), .CLK(clk), .RST(rst), .Q(c[430]) );
  DFF \sreg_reg[429]  ( .D(c[430]), .CLK(clk), .RST(rst), .Q(c[429]) );
  DFF \sreg_reg[428]  ( .D(c[429]), .CLK(clk), .RST(rst), .Q(c[428]) );
  DFF \sreg_reg[427]  ( .D(c[428]), .CLK(clk), .RST(rst), .Q(c[427]) );
  DFF \sreg_reg[426]  ( .D(c[427]), .CLK(clk), .RST(rst), .Q(c[426]) );
  DFF \sreg_reg[425]  ( .D(c[426]), .CLK(clk), .RST(rst), .Q(c[425]) );
  DFF \sreg_reg[424]  ( .D(c[425]), .CLK(clk), .RST(rst), .Q(c[424]) );
  DFF \sreg_reg[423]  ( .D(c[424]), .CLK(clk), .RST(rst), .Q(c[423]) );
  DFF \sreg_reg[422]  ( .D(c[423]), .CLK(clk), .RST(rst), .Q(c[422]) );
  DFF \sreg_reg[421]  ( .D(c[422]), .CLK(clk), .RST(rst), .Q(c[421]) );
  DFF \sreg_reg[420]  ( .D(c[421]), .CLK(clk), .RST(rst), .Q(c[420]) );
  DFF \sreg_reg[419]  ( .D(c[420]), .CLK(clk), .RST(rst), .Q(c[419]) );
  DFF \sreg_reg[418]  ( .D(c[419]), .CLK(clk), .RST(rst), .Q(c[418]) );
  DFF \sreg_reg[417]  ( .D(c[418]), .CLK(clk), .RST(rst), .Q(c[417]) );
  DFF \sreg_reg[416]  ( .D(c[417]), .CLK(clk), .RST(rst), .Q(c[416]) );
  DFF \sreg_reg[415]  ( .D(c[416]), .CLK(clk), .RST(rst), .Q(c[415]) );
  DFF \sreg_reg[414]  ( .D(c[415]), .CLK(clk), .RST(rst), .Q(c[414]) );
  DFF \sreg_reg[413]  ( .D(c[414]), .CLK(clk), .RST(rst), .Q(c[413]) );
  DFF \sreg_reg[412]  ( .D(c[413]), .CLK(clk), .RST(rst), .Q(c[412]) );
  DFF \sreg_reg[411]  ( .D(c[412]), .CLK(clk), .RST(rst), .Q(c[411]) );
  DFF \sreg_reg[410]  ( .D(c[411]), .CLK(clk), .RST(rst), .Q(c[410]) );
  DFF \sreg_reg[409]  ( .D(c[410]), .CLK(clk), .RST(rst), .Q(c[409]) );
  DFF \sreg_reg[408]  ( .D(c[409]), .CLK(clk), .RST(rst), .Q(c[408]) );
  DFF \sreg_reg[407]  ( .D(c[408]), .CLK(clk), .RST(rst), .Q(c[407]) );
  DFF \sreg_reg[406]  ( .D(c[407]), .CLK(clk), .RST(rst), .Q(c[406]) );
  DFF \sreg_reg[405]  ( .D(c[406]), .CLK(clk), .RST(rst), .Q(c[405]) );
  DFF \sreg_reg[404]  ( .D(c[405]), .CLK(clk), .RST(rst), .Q(c[404]) );
  DFF \sreg_reg[403]  ( .D(c[404]), .CLK(clk), .RST(rst), .Q(c[403]) );
  DFF \sreg_reg[402]  ( .D(c[403]), .CLK(clk), .RST(rst), .Q(c[402]) );
  DFF \sreg_reg[401]  ( .D(c[402]), .CLK(clk), .RST(rst), .Q(c[401]) );
  DFF \sreg_reg[400]  ( .D(c[401]), .CLK(clk), .RST(rst), .Q(c[400]) );
  DFF \sreg_reg[399]  ( .D(c[400]), .CLK(clk), .RST(rst), .Q(c[399]) );
  DFF \sreg_reg[398]  ( .D(c[399]), .CLK(clk), .RST(rst), .Q(c[398]) );
  DFF \sreg_reg[397]  ( .D(c[398]), .CLK(clk), .RST(rst), .Q(c[397]) );
  DFF \sreg_reg[396]  ( .D(c[397]), .CLK(clk), .RST(rst), .Q(c[396]) );
  DFF \sreg_reg[395]  ( .D(c[396]), .CLK(clk), .RST(rst), .Q(c[395]) );
  DFF \sreg_reg[394]  ( .D(c[395]), .CLK(clk), .RST(rst), .Q(c[394]) );
  DFF \sreg_reg[393]  ( .D(c[394]), .CLK(clk), .RST(rst), .Q(c[393]) );
  DFF \sreg_reg[392]  ( .D(c[393]), .CLK(clk), .RST(rst), .Q(c[392]) );
  DFF \sreg_reg[391]  ( .D(c[392]), .CLK(clk), .RST(rst), .Q(c[391]) );
  DFF \sreg_reg[390]  ( .D(c[391]), .CLK(clk), .RST(rst), .Q(c[390]) );
  DFF \sreg_reg[389]  ( .D(c[390]), .CLK(clk), .RST(rst), .Q(c[389]) );
  DFF \sreg_reg[388]  ( .D(c[389]), .CLK(clk), .RST(rst), .Q(c[388]) );
  DFF \sreg_reg[387]  ( .D(c[388]), .CLK(clk), .RST(rst), .Q(c[387]) );
  DFF \sreg_reg[386]  ( .D(c[387]), .CLK(clk), .RST(rst), .Q(c[386]) );
  DFF \sreg_reg[385]  ( .D(c[386]), .CLK(clk), .RST(rst), .Q(c[385]) );
  DFF \sreg_reg[384]  ( .D(c[385]), .CLK(clk), .RST(rst), .Q(c[384]) );
  DFF \sreg_reg[383]  ( .D(c[384]), .CLK(clk), .RST(rst), .Q(c[383]) );
  DFF \sreg_reg[382]  ( .D(c[383]), .CLK(clk), .RST(rst), .Q(c[382]) );
  DFF \sreg_reg[381]  ( .D(c[382]), .CLK(clk), .RST(rst), .Q(c[381]) );
  DFF \sreg_reg[380]  ( .D(c[381]), .CLK(clk), .RST(rst), .Q(c[380]) );
  DFF \sreg_reg[379]  ( .D(c[380]), .CLK(clk), .RST(rst), .Q(c[379]) );
  DFF \sreg_reg[378]  ( .D(c[379]), .CLK(clk), .RST(rst), .Q(c[378]) );
  DFF \sreg_reg[377]  ( .D(c[378]), .CLK(clk), .RST(rst), .Q(c[377]) );
  DFF \sreg_reg[376]  ( .D(c[377]), .CLK(clk), .RST(rst), .Q(c[376]) );
  DFF \sreg_reg[375]  ( .D(c[376]), .CLK(clk), .RST(rst), .Q(c[375]) );
  DFF \sreg_reg[374]  ( .D(c[375]), .CLK(clk), .RST(rst), .Q(c[374]) );
  DFF \sreg_reg[373]  ( .D(c[374]), .CLK(clk), .RST(rst), .Q(c[373]) );
  DFF \sreg_reg[372]  ( .D(c[373]), .CLK(clk), .RST(rst), .Q(c[372]) );
  DFF \sreg_reg[371]  ( .D(c[372]), .CLK(clk), .RST(rst), .Q(c[371]) );
  DFF \sreg_reg[370]  ( .D(c[371]), .CLK(clk), .RST(rst), .Q(c[370]) );
  DFF \sreg_reg[369]  ( .D(c[370]), .CLK(clk), .RST(rst), .Q(c[369]) );
  DFF \sreg_reg[368]  ( .D(c[369]), .CLK(clk), .RST(rst), .Q(c[368]) );
  DFF \sreg_reg[367]  ( .D(c[368]), .CLK(clk), .RST(rst), .Q(c[367]) );
  DFF \sreg_reg[366]  ( .D(c[367]), .CLK(clk), .RST(rst), .Q(c[366]) );
  DFF \sreg_reg[365]  ( .D(c[366]), .CLK(clk), .RST(rst), .Q(c[365]) );
  DFF \sreg_reg[364]  ( .D(c[365]), .CLK(clk), .RST(rst), .Q(c[364]) );
  DFF \sreg_reg[363]  ( .D(c[364]), .CLK(clk), .RST(rst), .Q(c[363]) );
  DFF \sreg_reg[362]  ( .D(c[363]), .CLK(clk), .RST(rst), .Q(c[362]) );
  DFF \sreg_reg[361]  ( .D(c[362]), .CLK(clk), .RST(rst), .Q(c[361]) );
  DFF \sreg_reg[360]  ( .D(c[361]), .CLK(clk), .RST(rst), .Q(c[360]) );
  DFF \sreg_reg[359]  ( .D(c[360]), .CLK(clk), .RST(rst), .Q(c[359]) );
  DFF \sreg_reg[358]  ( .D(c[359]), .CLK(clk), .RST(rst), .Q(c[358]) );
  DFF \sreg_reg[357]  ( .D(c[358]), .CLK(clk), .RST(rst), .Q(c[357]) );
  DFF \sreg_reg[356]  ( .D(c[357]), .CLK(clk), .RST(rst), .Q(c[356]) );
  DFF \sreg_reg[355]  ( .D(c[356]), .CLK(clk), .RST(rst), .Q(c[355]) );
  DFF \sreg_reg[354]  ( .D(c[355]), .CLK(clk), .RST(rst), .Q(c[354]) );
  DFF \sreg_reg[353]  ( .D(c[354]), .CLK(clk), .RST(rst), .Q(c[353]) );
  DFF \sreg_reg[352]  ( .D(c[353]), .CLK(clk), .RST(rst), .Q(c[352]) );
  DFF \sreg_reg[351]  ( .D(c[352]), .CLK(clk), .RST(rst), .Q(c[351]) );
  DFF \sreg_reg[350]  ( .D(c[351]), .CLK(clk), .RST(rst), .Q(c[350]) );
  DFF \sreg_reg[349]  ( .D(c[350]), .CLK(clk), .RST(rst), .Q(c[349]) );
  DFF \sreg_reg[348]  ( .D(c[349]), .CLK(clk), .RST(rst), .Q(c[348]) );
  DFF \sreg_reg[347]  ( .D(c[348]), .CLK(clk), .RST(rst), .Q(c[347]) );
  DFF \sreg_reg[346]  ( .D(c[347]), .CLK(clk), .RST(rst), .Q(c[346]) );
  DFF \sreg_reg[345]  ( .D(c[346]), .CLK(clk), .RST(rst), .Q(c[345]) );
  DFF \sreg_reg[344]  ( .D(c[345]), .CLK(clk), .RST(rst), .Q(c[344]) );
  DFF \sreg_reg[343]  ( .D(c[344]), .CLK(clk), .RST(rst), .Q(c[343]) );
  DFF \sreg_reg[342]  ( .D(c[343]), .CLK(clk), .RST(rst), .Q(c[342]) );
  DFF \sreg_reg[341]  ( .D(c[342]), .CLK(clk), .RST(rst), .Q(c[341]) );
  DFF \sreg_reg[340]  ( .D(c[341]), .CLK(clk), .RST(rst), .Q(c[340]) );
  DFF \sreg_reg[339]  ( .D(c[340]), .CLK(clk), .RST(rst), .Q(c[339]) );
  DFF \sreg_reg[338]  ( .D(c[339]), .CLK(clk), .RST(rst), .Q(c[338]) );
  DFF \sreg_reg[337]  ( .D(c[338]), .CLK(clk), .RST(rst), .Q(c[337]) );
  DFF \sreg_reg[336]  ( .D(c[337]), .CLK(clk), .RST(rst), .Q(c[336]) );
  DFF \sreg_reg[335]  ( .D(c[336]), .CLK(clk), .RST(rst), .Q(c[335]) );
  DFF \sreg_reg[334]  ( .D(c[335]), .CLK(clk), .RST(rst), .Q(c[334]) );
  DFF \sreg_reg[333]  ( .D(c[334]), .CLK(clk), .RST(rst), .Q(c[333]) );
  DFF \sreg_reg[332]  ( .D(c[333]), .CLK(clk), .RST(rst), .Q(c[332]) );
  DFF \sreg_reg[331]  ( .D(c[332]), .CLK(clk), .RST(rst), .Q(c[331]) );
  DFF \sreg_reg[330]  ( .D(c[331]), .CLK(clk), .RST(rst), .Q(c[330]) );
  DFF \sreg_reg[329]  ( .D(c[330]), .CLK(clk), .RST(rst), .Q(c[329]) );
  DFF \sreg_reg[328]  ( .D(c[329]), .CLK(clk), .RST(rst), .Q(c[328]) );
  DFF \sreg_reg[327]  ( .D(c[328]), .CLK(clk), .RST(rst), .Q(c[327]) );
  DFF \sreg_reg[326]  ( .D(c[327]), .CLK(clk), .RST(rst), .Q(c[326]) );
  DFF \sreg_reg[325]  ( .D(c[326]), .CLK(clk), .RST(rst), .Q(c[325]) );
  DFF \sreg_reg[324]  ( .D(c[325]), .CLK(clk), .RST(rst), .Q(c[324]) );
  DFF \sreg_reg[323]  ( .D(c[324]), .CLK(clk), .RST(rst), .Q(c[323]) );
  DFF \sreg_reg[322]  ( .D(c[323]), .CLK(clk), .RST(rst), .Q(c[322]) );
  DFF \sreg_reg[321]  ( .D(c[322]), .CLK(clk), .RST(rst), .Q(c[321]) );
  DFF \sreg_reg[320]  ( .D(c[321]), .CLK(clk), .RST(rst), .Q(c[320]) );
  DFF \sreg_reg[319]  ( .D(c[320]), .CLK(clk), .RST(rst), .Q(c[319]) );
  DFF \sreg_reg[318]  ( .D(c[319]), .CLK(clk), .RST(rst), .Q(c[318]) );
  DFF \sreg_reg[317]  ( .D(c[318]), .CLK(clk), .RST(rst), .Q(c[317]) );
  DFF \sreg_reg[316]  ( .D(c[317]), .CLK(clk), .RST(rst), .Q(c[316]) );
  DFF \sreg_reg[315]  ( .D(c[316]), .CLK(clk), .RST(rst), .Q(c[315]) );
  DFF \sreg_reg[314]  ( .D(c[315]), .CLK(clk), .RST(rst), .Q(c[314]) );
  DFF \sreg_reg[313]  ( .D(c[314]), .CLK(clk), .RST(rst), .Q(c[313]) );
  DFF \sreg_reg[312]  ( .D(c[313]), .CLK(clk), .RST(rst), .Q(c[312]) );
  DFF \sreg_reg[311]  ( .D(c[312]), .CLK(clk), .RST(rst), .Q(c[311]) );
  DFF \sreg_reg[310]  ( .D(c[311]), .CLK(clk), .RST(rst), .Q(c[310]) );
  DFF \sreg_reg[309]  ( .D(c[310]), .CLK(clk), .RST(rst), .Q(c[309]) );
  DFF \sreg_reg[308]  ( .D(c[309]), .CLK(clk), .RST(rst), .Q(c[308]) );
  DFF \sreg_reg[307]  ( .D(c[308]), .CLK(clk), .RST(rst), .Q(c[307]) );
  DFF \sreg_reg[306]  ( .D(c[307]), .CLK(clk), .RST(rst), .Q(c[306]) );
  DFF \sreg_reg[305]  ( .D(c[306]), .CLK(clk), .RST(rst), .Q(c[305]) );
  DFF \sreg_reg[304]  ( .D(c[305]), .CLK(clk), .RST(rst), .Q(c[304]) );
  DFF \sreg_reg[303]  ( .D(c[304]), .CLK(clk), .RST(rst), .Q(c[303]) );
  DFF \sreg_reg[302]  ( .D(c[303]), .CLK(clk), .RST(rst), .Q(c[302]) );
  DFF \sreg_reg[301]  ( .D(c[302]), .CLK(clk), .RST(rst), .Q(c[301]) );
  DFF \sreg_reg[300]  ( .D(c[301]), .CLK(clk), .RST(rst), .Q(c[300]) );
  DFF \sreg_reg[299]  ( .D(c[300]), .CLK(clk), .RST(rst), .Q(c[299]) );
  DFF \sreg_reg[298]  ( .D(c[299]), .CLK(clk), .RST(rst), .Q(c[298]) );
  DFF \sreg_reg[297]  ( .D(c[298]), .CLK(clk), .RST(rst), .Q(c[297]) );
  DFF \sreg_reg[296]  ( .D(c[297]), .CLK(clk), .RST(rst), .Q(c[296]) );
  DFF \sreg_reg[295]  ( .D(c[296]), .CLK(clk), .RST(rst), .Q(c[295]) );
  DFF \sreg_reg[294]  ( .D(c[295]), .CLK(clk), .RST(rst), .Q(c[294]) );
  DFF \sreg_reg[293]  ( .D(c[294]), .CLK(clk), .RST(rst), .Q(c[293]) );
  DFF \sreg_reg[292]  ( .D(c[293]), .CLK(clk), .RST(rst), .Q(c[292]) );
  DFF \sreg_reg[291]  ( .D(c[292]), .CLK(clk), .RST(rst), .Q(c[291]) );
  DFF \sreg_reg[290]  ( .D(c[291]), .CLK(clk), .RST(rst), .Q(c[290]) );
  DFF \sreg_reg[289]  ( .D(c[290]), .CLK(clk), .RST(rst), .Q(c[289]) );
  DFF \sreg_reg[288]  ( .D(c[289]), .CLK(clk), .RST(rst), .Q(c[288]) );
  DFF \sreg_reg[287]  ( .D(c[288]), .CLK(clk), .RST(rst), .Q(c[287]) );
  DFF \sreg_reg[286]  ( .D(c[287]), .CLK(clk), .RST(rst), .Q(c[286]) );
  DFF \sreg_reg[285]  ( .D(c[286]), .CLK(clk), .RST(rst), .Q(c[285]) );
  DFF \sreg_reg[284]  ( .D(c[285]), .CLK(clk), .RST(rst), .Q(c[284]) );
  DFF \sreg_reg[283]  ( .D(c[284]), .CLK(clk), .RST(rst), .Q(c[283]) );
  DFF \sreg_reg[282]  ( .D(c[283]), .CLK(clk), .RST(rst), .Q(c[282]) );
  DFF \sreg_reg[281]  ( .D(c[282]), .CLK(clk), .RST(rst), .Q(c[281]) );
  DFF \sreg_reg[280]  ( .D(c[281]), .CLK(clk), .RST(rst), .Q(c[280]) );
  DFF \sreg_reg[279]  ( .D(c[280]), .CLK(clk), .RST(rst), .Q(c[279]) );
  DFF \sreg_reg[278]  ( .D(c[279]), .CLK(clk), .RST(rst), .Q(c[278]) );
  DFF \sreg_reg[277]  ( .D(c[278]), .CLK(clk), .RST(rst), .Q(c[277]) );
  DFF \sreg_reg[276]  ( .D(c[277]), .CLK(clk), .RST(rst), .Q(c[276]) );
  DFF \sreg_reg[275]  ( .D(c[276]), .CLK(clk), .RST(rst), .Q(c[275]) );
  DFF \sreg_reg[274]  ( .D(c[275]), .CLK(clk), .RST(rst), .Q(c[274]) );
  DFF \sreg_reg[273]  ( .D(c[274]), .CLK(clk), .RST(rst), .Q(c[273]) );
  DFF \sreg_reg[272]  ( .D(c[273]), .CLK(clk), .RST(rst), .Q(c[272]) );
  DFF \sreg_reg[271]  ( .D(c[272]), .CLK(clk), .RST(rst), .Q(c[271]) );
  DFF \sreg_reg[270]  ( .D(c[271]), .CLK(clk), .RST(rst), .Q(c[270]) );
  DFF \sreg_reg[269]  ( .D(c[270]), .CLK(clk), .RST(rst), .Q(c[269]) );
  DFF \sreg_reg[268]  ( .D(c[269]), .CLK(clk), .RST(rst), .Q(c[268]) );
  DFF \sreg_reg[267]  ( .D(c[268]), .CLK(clk), .RST(rst), .Q(c[267]) );
  DFF \sreg_reg[266]  ( .D(c[267]), .CLK(clk), .RST(rst), .Q(c[266]) );
  DFF \sreg_reg[265]  ( .D(c[266]), .CLK(clk), .RST(rst), .Q(c[265]) );
  DFF \sreg_reg[264]  ( .D(c[265]), .CLK(clk), .RST(rst), .Q(c[264]) );
  DFF \sreg_reg[263]  ( .D(c[264]), .CLK(clk), .RST(rst), .Q(c[263]) );
  DFF \sreg_reg[262]  ( .D(c[263]), .CLK(clk), .RST(rst), .Q(c[262]) );
  DFF \sreg_reg[261]  ( .D(c[262]), .CLK(clk), .RST(rst), .Q(c[261]) );
  DFF \sreg_reg[260]  ( .D(c[261]), .CLK(clk), .RST(rst), .Q(c[260]) );
  DFF \sreg_reg[259]  ( .D(c[260]), .CLK(clk), .RST(rst), .Q(c[259]) );
  DFF \sreg_reg[258]  ( .D(c[259]), .CLK(clk), .RST(rst), .Q(c[258]) );
  DFF \sreg_reg[257]  ( .D(c[258]), .CLK(clk), .RST(rst), .Q(c[257]) );
  DFF \sreg_reg[256]  ( .D(c[257]), .CLK(clk), .RST(rst), .Q(c[256]) );
  DFF \sreg_reg[255]  ( .D(c[256]), .CLK(clk), .RST(rst), .Q(c[255]) );
  DFF \sreg_reg[254]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(c[254]) );
  DFF \sreg_reg[253]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(c[253]) );
  DFF \sreg_reg[252]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(c[252]) );
  DFF \sreg_reg[251]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(c[251]) );
  DFF \sreg_reg[250]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(c[250]) );
  DFF \sreg_reg[249]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(c[249]) );
  DFF \sreg_reg[248]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(c[248]) );
  DFF \sreg_reg[247]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(c[247]) );
  DFF \sreg_reg[246]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(c[246]) );
  DFF \sreg_reg[245]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(c[245]) );
  DFF \sreg_reg[244]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(c[244]) );
  DFF \sreg_reg[243]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(c[243]) );
  DFF \sreg_reg[242]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(c[242]) );
  DFF \sreg_reg[241]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(c[241]) );
  DFF \sreg_reg[240]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(c[240]) );
  DFF \sreg_reg[239]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(c[239]) );
  DFF \sreg_reg[238]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(c[238]) );
  DFF \sreg_reg[237]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(c[237]) );
  DFF \sreg_reg[236]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(c[236]) );
  DFF \sreg_reg[235]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(c[235]) );
  DFF \sreg_reg[234]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(c[234]) );
  DFF \sreg_reg[233]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(c[233]) );
  DFF \sreg_reg[232]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(c[232]) );
  DFF \sreg_reg[231]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(c[231]) );
  DFF \sreg_reg[230]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(c[230]) );
  DFF \sreg_reg[229]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(c[229]) );
  DFF \sreg_reg[228]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(c[228]) );
  DFF \sreg_reg[227]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(c[227]) );
  DFF \sreg_reg[226]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(c[226]) );
  DFF \sreg_reg[225]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(c[225]) );
  DFF \sreg_reg[224]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(c[224]) );
  DFF \sreg_reg[223]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(c[223]) );
  DFF \sreg_reg[222]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(c[222]) );
  DFF \sreg_reg[221]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(c[221]) );
  DFF \sreg_reg[220]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(c[220]) );
  DFF \sreg_reg[219]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(c[219]) );
  DFF \sreg_reg[218]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(c[218]) );
  DFF \sreg_reg[217]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(c[217]) );
  DFF \sreg_reg[216]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(c[216]) );
  DFF \sreg_reg[215]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(c[215]) );
  DFF \sreg_reg[214]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(c[214]) );
  DFF \sreg_reg[213]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(c[213]) );
  DFF \sreg_reg[212]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(c[212]) );
  DFF \sreg_reg[211]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(c[211]) );
  DFF \sreg_reg[210]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(c[210]) );
  DFF \sreg_reg[209]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(c[209]) );
  DFF \sreg_reg[208]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(c[208]) );
  DFF \sreg_reg[207]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(c[207]) );
  DFF \sreg_reg[206]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(c[206]) );
  DFF \sreg_reg[205]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(c[205]) );
  DFF \sreg_reg[204]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(c[204]) );
  DFF \sreg_reg[203]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(c[203]) );
  DFF \sreg_reg[202]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(c[202]) );
  DFF \sreg_reg[201]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(c[201]) );
  DFF \sreg_reg[200]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(c[200]) );
  DFF \sreg_reg[199]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(c[199]) );
  DFF \sreg_reg[198]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(c[198]) );
  DFF \sreg_reg[197]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(c[197]) );
  DFF \sreg_reg[196]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(c[196]) );
  DFF \sreg_reg[195]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(c[195]) );
  DFF \sreg_reg[194]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(c[194]) );
  DFF \sreg_reg[193]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(c[193]) );
  DFF \sreg_reg[192]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(c[192]) );
  DFF \sreg_reg[191]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(c[191]) );
  DFF \sreg_reg[190]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(c[190]) );
  DFF \sreg_reg[189]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(c[189]) );
  DFF \sreg_reg[188]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(c[188]) );
  DFF \sreg_reg[187]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(c[187]) );
  DFF \sreg_reg[186]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(c[186]) );
  DFF \sreg_reg[185]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(c[185]) );
  DFF \sreg_reg[184]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(c[184]) );
  DFF \sreg_reg[183]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(c[183]) );
  DFF \sreg_reg[182]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(c[182]) );
  DFF \sreg_reg[181]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(c[181]) );
  DFF \sreg_reg[180]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(c[180]) );
  DFF \sreg_reg[179]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(c[179]) );
  DFF \sreg_reg[178]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(c[178]) );
  DFF \sreg_reg[177]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(c[177]) );
  DFF \sreg_reg[176]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(c[176]) );
  DFF \sreg_reg[175]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(c[175]) );
  DFF \sreg_reg[174]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(c[174]) );
  DFF \sreg_reg[173]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(c[173]) );
  DFF \sreg_reg[172]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(c[172]) );
  DFF \sreg_reg[171]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(c[171]) );
  DFF \sreg_reg[170]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(c[170]) );
  DFF \sreg_reg[169]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(c[169]) );
  DFF \sreg_reg[168]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(c[168]) );
  DFF \sreg_reg[167]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(c[167]) );
  DFF \sreg_reg[166]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(c[166]) );
  DFF \sreg_reg[165]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(c[165]) );
  DFF \sreg_reg[164]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(c[164]) );
  DFF \sreg_reg[163]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(c[163]) );
  DFF \sreg_reg[162]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(c[162]) );
  DFF \sreg_reg[161]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(c[161]) );
  DFF \sreg_reg[160]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(c[160]) );
  DFF \sreg_reg[159]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(c[159]) );
  DFF \sreg_reg[158]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(c[158]) );
  DFF \sreg_reg[157]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(c[157]) );
  DFF \sreg_reg[156]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(c[156]) );
  DFF \sreg_reg[155]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(c[155]) );
  DFF \sreg_reg[154]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(c[154]) );
  DFF \sreg_reg[153]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(c[153]) );
  DFF \sreg_reg[152]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(c[152]) );
  DFF \sreg_reg[151]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(c[151]) );
  DFF \sreg_reg[150]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(c[150]) );
  DFF \sreg_reg[149]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(c[149]) );
  DFF \sreg_reg[148]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(c[148]) );
  DFF \sreg_reg[147]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(c[147]) );
  DFF \sreg_reg[146]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(c[146]) );
  DFF \sreg_reg[145]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(c[145]) );
  DFF \sreg_reg[144]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(c[144]) );
  DFF \sreg_reg[143]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(c[143]) );
  DFF \sreg_reg[142]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(c[142]) );
  DFF \sreg_reg[141]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(c[141]) );
  DFF \sreg_reg[140]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(c[140]) );
  DFF \sreg_reg[139]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(c[139]) );
  DFF \sreg_reg[138]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(c[138]) );
  DFF \sreg_reg[137]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(c[137]) );
  DFF \sreg_reg[136]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(c[136]) );
  DFF \sreg_reg[135]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(c[135]) );
  DFF \sreg_reg[134]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(c[134]) );
  DFF \sreg_reg[133]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(c[133]) );
  DFF \sreg_reg[132]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(c[132]) );
  DFF \sreg_reg[131]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(c[131]) );
  DFF \sreg_reg[130]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(c[130]) );
  DFF \sreg_reg[129]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(c[129]) );
  DFF \sreg_reg[128]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(c[128]) );
  DFF \sreg_reg[127]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(c[127]) );
  DFF \sreg_reg[126]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[125]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[124]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[123]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[3]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[2]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[1]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NAND U4 ( .A(n422), .B(sreg[1069]), .Z(n1) );
  XOR U5 ( .A(n422), .B(sreg[1069]), .Z(n2) );
  NANDN U6 ( .A(n421), .B(n2), .Z(n3) );
  NAND U7 ( .A(n1), .B(n3), .Z(n424) );
  XOR U8 ( .A(n621), .B(sreg[1111]), .Z(n4) );
  NANDN U9 ( .A(n622), .B(n4), .Z(n5) );
  NAND U10 ( .A(n621), .B(sreg[1111]), .Z(n6) );
  AND U11 ( .A(n5), .B(n6), .Z(n625) );
  NAND U12 ( .A(sreg[1135]), .B(n736), .Z(n7) );
  XOR U13 ( .A(sreg[1135]), .B(n736), .Z(n8) );
  NANDN U14 ( .A(n735), .B(n8), .Z(n9) );
  NAND U15 ( .A(n7), .B(n9), .Z(n739) );
  XOR U16 ( .A(n1303), .B(sreg[1253]), .Z(n10) );
  NANDN U17 ( .A(n1304), .B(n10), .Z(n11) );
  NAND U18 ( .A(n1303), .B(sreg[1253]), .Z(n12) );
  AND U19 ( .A(n11), .B(n12), .Z(n1307) );
  NAND U20 ( .A(n2126), .B(sreg[1421]), .Z(n13) );
  XOR U21 ( .A(n2126), .B(sreg[1421]), .Z(n14) );
  NANDN U22 ( .A(n2125), .B(n14), .Z(n15) );
  NAND U23 ( .A(n13), .B(n15), .Z(n2128) );
  NAND U24 ( .A(n4492), .B(sreg[1901]), .Z(n16) );
  XOR U25 ( .A(n4492), .B(sreg[1901]), .Z(n17) );
  NANDN U26 ( .A(n4491), .B(n17), .Z(n18) );
  NAND U27 ( .A(n16), .B(n18), .Z(n4494) );
  NAND U28 ( .A(sreg[1913]), .B(n4548), .Z(n19) );
  XOR U29 ( .A(sreg[1913]), .B(n4548), .Z(n20) );
  NANDN U30 ( .A(n4547), .B(n20), .Z(n21) );
  NAND U31 ( .A(n19), .B(n21), .Z(n4550) );
  NAND U32 ( .A(sreg[1959]), .B(n4771), .Z(n22) );
  XOR U33 ( .A(sreg[1959]), .B(n4771), .Z(n23) );
  NANDN U34 ( .A(n4772), .B(n23), .Z(n24) );
  NAND U35 ( .A(n22), .B(n24), .Z(n4775) );
  NAND U36 ( .A(sreg[2013]), .B(n5026), .Z(n25) );
  XOR U37 ( .A(sreg[2013]), .B(n5026), .Z(n26) );
  NANDN U38 ( .A(n5025), .B(n26), .Z(n27) );
  NAND U39 ( .A(n25), .B(n27), .Z(n5029) );
  XOR U40 ( .A(n5036), .B(sreg[2016]), .Z(n28) );
  NANDN U41 ( .A(n5037), .B(n28), .Z(n29) );
  NAND U42 ( .A(n5036), .B(sreg[2016]), .Z(n30) );
  AND U43 ( .A(n29), .B(n30), .Z(n5040) );
  NAND U44 ( .A(sreg[1024]), .B(n199), .Z(n31) );
  XOR U45 ( .A(sreg[1024]), .B(n199), .Z(n32) );
  NANDN U46 ( .A(n198), .B(n32), .Z(n33) );
  NAND U47 ( .A(n31), .B(n33), .Z(n202) );
  XOR U48 ( .A(n429), .B(sreg[1071]), .Z(n34) );
  NANDN U49 ( .A(n430), .B(n34), .Z(n35) );
  NAND U50 ( .A(n429), .B(sreg[1071]), .Z(n36) );
  AND U51 ( .A(n35), .B(n36), .Z(n433) );
  NAND U52 ( .A(sreg[1074]), .B(n443), .Z(n37) );
  XOR U53 ( .A(sreg[1074]), .B(n443), .Z(n38) );
  NANDN U54 ( .A(n442), .B(n38), .Z(n39) );
  NAND U55 ( .A(n37), .B(n39), .Z(n446) );
  XOR U56 ( .A(n455), .B(sreg[1077]), .Z(n40) );
  NANDN U57 ( .A(n456), .B(n40), .Z(n41) );
  NAND U58 ( .A(n455), .B(sreg[1077]), .Z(n42) );
  AND U59 ( .A(n41), .B(n42), .Z(n459) );
  NAND U60 ( .A(sreg[1080]), .B(n469), .Z(n43) );
  XOR U61 ( .A(sreg[1080]), .B(n469), .Z(n44) );
  NANDN U62 ( .A(n468), .B(n44), .Z(n45) );
  NAND U63 ( .A(n43), .B(n45), .Z(n472) );
  XOR U64 ( .A(n629), .B(sreg[1113]), .Z(n46) );
  NANDN U65 ( .A(n630), .B(n46), .Z(n47) );
  NAND U66 ( .A(n629), .B(sreg[1113]), .Z(n48) );
  AND U67 ( .A(n47), .B(n48), .Z(n633) );
  NAND U68 ( .A(sreg[1133]), .B(n728), .Z(n49) );
  XOR U69 ( .A(sreg[1133]), .B(n728), .Z(n50) );
  NANDN U70 ( .A(n727), .B(n50), .Z(n51) );
  NAND U71 ( .A(n49), .B(n51), .Z(n731) );
  NAND U72 ( .A(sreg[1136]), .B(n739), .Z(n52) );
  XOR U73 ( .A(sreg[1136]), .B(n739), .Z(n53) );
  NANDN U74 ( .A(n738), .B(n53), .Z(n54) );
  NAND U75 ( .A(n52), .B(n54), .Z(n742) );
  NAND U76 ( .A(sreg[1167]), .B(n891), .Z(n55) );
  XOR U77 ( .A(sreg[1167]), .B(n891), .Z(n56) );
  NANDN U78 ( .A(n892), .B(n56), .Z(n57) );
  NAND U79 ( .A(n55), .B(n57), .Z(n895) );
  XOR U80 ( .A(n904), .B(sreg[1170]), .Z(n58) );
  NANDN U81 ( .A(n905), .B(n58), .Z(n59) );
  NAND U82 ( .A(n904), .B(sreg[1170]), .Z(n60) );
  AND U83 ( .A(n59), .B(n60), .Z(n908) );
  NAND U84 ( .A(sreg[1173]), .B(n918), .Z(n61) );
  XOR U85 ( .A(sreg[1173]), .B(n918), .Z(n62) );
  NANDN U86 ( .A(n917), .B(n62), .Z(n63) );
  NAND U87 ( .A(n61), .B(n63), .Z(n921) );
  XOR U88 ( .A(n930), .B(sreg[1176]), .Z(n64) );
  NANDN U89 ( .A(n931), .B(n64), .Z(n65) );
  NAND U90 ( .A(n930), .B(sreg[1176]), .Z(n66) );
  AND U91 ( .A(n65), .B(n66), .Z(n934) );
  NAND U92 ( .A(sreg[1231]), .B(n1203), .Z(n67) );
  XOR U93 ( .A(sreg[1231]), .B(n1203), .Z(n68) );
  NANDN U94 ( .A(n1204), .B(n68), .Z(n69) );
  NAND U95 ( .A(n67), .B(n69), .Z(n1207) );
  XOR U96 ( .A(n1251), .B(sreg[1241]), .Z(n70) );
  NANDN U97 ( .A(n1252), .B(n70), .Z(n71) );
  NAND U98 ( .A(n1251), .B(sreg[1241]), .Z(n72) );
  AND U99 ( .A(n71), .B(n72), .Z(n1255) );
  NAND U100 ( .A(sreg[1244]), .B(n1265), .Z(n73) );
  XOR U101 ( .A(sreg[1244]), .B(n1265), .Z(n74) );
  NANDN U102 ( .A(n1264), .B(n74), .Z(n75) );
  NAND U103 ( .A(n73), .B(n75), .Z(n1268) );
  XOR U104 ( .A(n1277), .B(sreg[1247]), .Z(n76) );
  NANDN U105 ( .A(n1278), .B(n76), .Z(n77) );
  NAND U106 ( .A(n1277), .B(sreg[1247]), .Z(n78) );
  AND U107 ( .A(n77), .B(n78), .Z(n1281) );
  NAND U108 ( .A(sreg[1250]), .B(n1291), .Z(n79) );
  XOR U109 ( .A(sreg[1250]), .B(n1291), .Z(n80) );
  NANDN U110 ( .A(n1290), .B(n80), .Z(n81) );
  NAND U111 ( .A(n79), .B(n81), .Z(n1294) );
  NAND U112 ( .A(sreg[1255]), .B(n1312), .Z(n82) );
  XOR U113 ( .A(sreg[1255]), .B(n1312), .Z(n83) );
  NANDN U114 ( .A(n1311), .B(n83), .Z(n84) );
  NAND U115 ( .A(n82), .B(n84), .Z(n1315) );
  NAND U116 ( .A(sreg[1287]), .B(n1469), .Z(n85) );
  XOR U117 ( .A(sreg[1287]), .B(n1469), .Z(n86) );
  NANDN U118 ( .A(n1470), .B(n86), .Z(n87) );
  NAND U119 ( .A(n85), .B(n87), .Z(n1473) );
  XOR U120 ( .A(n1508), .B(n1507), .Z(n88) );
  NANDN U121 ( .A(sreg[1295]), .B(n88), .Z(n89) );
  NAND U122 ( .A(n1508), .B(n1507), .Z(n90) );
  AND U123 ( .A(n89), .B(n90), .Z(n1511) );
  NAND U124 ( .A(n1666), .B(sreg[1327]), .Z(n91) );
  XOR U125 ( .A(n1666), .B(sreg[1327]), .Z(n92) );
  NANDN U126 ( .A(n1665), .B(n92), .Z(n93) );
  NAND U127 ( .A(n91), .B(n93), .Z(n1668) );
  NAND U128 ( .A(sreg[1330]), .B(n1679), .Z(n94) );
  XOR U129 ( .A(sreg[1330]), .B(n1679), .Z(n95) );
  NANDN U130 ( .A(n1678), .B(n95), .Z(n96) );
  NAND U131 ( .A(n94), .B(n96), .Z(n1682) );
  NAND U132 ( .A(sreg[1338]), .B(n1717), .Z(n97) );
  XOR U133 ( .A(sreg[1338]), .B(n1717), .Z(n98) );
  NANDN U134 ( .A(n1716), .B(n98), .Z(n99) );
  NAND U135 ( .A(n97), .B(n99), .Z(n1720) );
  XOR U136 ( .A(n1759), .B(sreg[1347]), .Z(n100) );
  NANDN U137 ( .A(n1760), .B(n100), .Z(n101) );
  NAND U138 ( .A(n1759), .B(sreg[1347]), .Z(n102) );
  AND U139 ( .A(n101), .B(n102), .Z(n1763) );
  NAND U140 ( .A(n1978), .B(sreg[1391]), .Z(n103) );
  XOR U141 ( .A(n1978), .B(sreg[1391]), .Z(n104) );
  NANDN U142 ( .A(n1977), .B(n104), .Z(n105) );
  NAND U143 ( .A(n103), .B(n105), .Z(n1980) );
  XOR U144 ( .A(n2133), .B(sreg[1423]), .Z(n106) );
  NANDN U145 ( .A(n2134), .B(n106), .Z(n107) );
  NAND U146 ( .A(n2133), .B(sreg[1423]), .Z(n108) );
  AND U147 ( .A(n107), .B(n108), .Z(n2137) );
  NAND U148 ( .A(n2292), .B(sreg[1455]), .Z(n109) );
  XOR U149 ( .A(n2292), .B(sreg[1455]), .Z(n110) );
  NANDN U150 ( .A(n2291), .B(n110), .Z(n111) );
  NAND U151 ( .A(n109), .B(n111), .Z(n2294) );
  NAND U152 ( .A(sreg[1481]), .B(n2419), .Z(n112) );
  XOR U153 ( .A(sreg[1481]), .B(n2419), .Z(n113) );
  NANDN U154 ( .A(n2420), .B(n113), .Z(n114) );
  NAND U155 ( .A(n112), .B(n114), .Z(n2423) );
  NAND U156 ( .A(n2568), .B(sreg[1511]), .Z(n115) );
  XOR U157 ( .A(n2568), .B(sreg[1511]), .Z(n116) );
  NANDN U158 ( .A(n2567), .B(n116), .Z(n117) );
  NAND U159 ( .A(n115), .B(n117), .Z(n2570) );
  NAND U160 ( .A(sreg[1514]), .B(n2581), .Z(n118) );
  XOR U161 ( .A(sreg[1514]), .B(n2581), .Z(n119) );
  NANDN U162 ( .A(n2580), .B(n119), .Z(n120) );
  NAND U163 ( .A(n118), .B(n120), .Z(n2584) );
  NAND U164 ( .A(n2819), .B(sreg[1562]), .Z(n121) );
  XOR U165 ( .A(n2819), .B(sreg[1562]), .Z(n122) );
  NAND U166 ( .A(n122), .B(n2818), .Z(n123) );
  NAND U167 ( .A(n121), .B(n123), .Z(n2822) );
  NAND U168 ( .A(sreg[1615]), .B(n3081), .Z(n124) );
  XOR U169 ( .A(sreg[1615]), .B(n3081), .Z(n125) );
  NANDN U170 ( .A(n3082), .B(n125), .Z(n126) );
  NAND U171 ( .A(n124), .B(n126), .Z(n3085) );
  NAND U172 ( .A(sreg[1658]), .B(n3294), .Z(n127) );
  XOR U173 ( .A(sreg[1658]), .B(n3294), .Z(n128) );
  NANDN U174 ( .A(n3295), .B(n128), .Z(n129) );
  NAND U175 ( .A(n127), .B(n129), .Z(n3298) );
  NAND U176 ( .A(sreg[1679]), .B(n3398), .Z(n130) );
  XOR U177 ( .A(sreg[1679]), .B(n3398), .Z(n131) );
  NANDN U178 ( .A(n3397), .B(n131), .Z(n132) );
  NAND U179 ( .A(n130), .B(n132), .Z(n3402) );
  NAND U180 ( .A(n3548), .B(sreg[1709]), .Z(n133) );
  XOR U181 ( .A(n3548), .B(sreg[1709]), .Z(n134) );
  NANDN U182 ( .A(n3547), .B(n134), .Z(n135) );
  NAND U183 ( .A(n133), .B(n135), .Z(n3550) );
  NAND U184 ( .A(sreg[1712]), .B(n3561), .Z(n136) );
  XOR U185 ( .A(sreg[1712]), .B(n3561), .Z(n137) );
  NANDN U186 ( .A(n3560), .B(n137), .Z(n138) );
  NAND U187 ( .A(n136), .B(n138), .Z(n3564) );
  XOR U188 ( .A(n3828), .B(sreg[1766]), .Z(n139) );
  NANDN U189 ( .A(n3829), .B(n139), .Z(n140) );
  NAND U190 ( .A(n3828), .B(sreg[1766]), .Z(n141) );
  AND U191 ( .A(n140), .B(n141), .Z(n3832) );
  NAND U192 ( .A(sreg[1769]), .B(n3842), .Z(n142) );
  XOR U193 ( .A(sreg[1769]), .B(n3842), .Z(n143) );
  NANDN U194 ( .A(n3841), .B(n143), .Z(n144) );
  NAND U195 ( .A(n142), .B(n144), .Z(n3845) );
  XOR U196 ( .A(n3854), .B(sreg[1772]), .Z(n145) );
  NANDN U197 ( .A(n3855), .B(n145), .Z(n146) );
  NAND U198 ( .A(n3854), .B(sreg[1772]), .Z(n147) );
  AND U199 ( .A(n146), .B(n147), .Z(n3858) );
  XOR U200 ( .A(n3867), .B(sreg[1775]), .Z(n148) );
  NANDN U201 ( .A(n3868), .B(n148), .Z(n149) );
  NAND U202 ( .A(n3867), .B(sreg[1775]), .Z(n150) );
  AND U203 ( .A(n149), .B(n150), .Z(n3871) );
  XOR U204 ( .A(n4241), .B(n4240), .Z(n151) );
  NANDN U205 ( .A(sreg[1850]), .B(n151), .Z(n152) );
  NAND U206 ( .A(n4241), .B(n4240), .Z(n153) );
  AND U207 ( .A(n152), .B(n153), .Z(n4243) );
  NAND U208 ( .A(sreg[1871]), .B(n4343), .Z(n154) );
  XOR U209 ( .A(sreg[1871]), .B(n4343), .Z(n155) );
  NANDN U210 ( .A(n4344), .B(n155), .Z(n156) );
  NAND U211 ( .A(n154), .B(n156), .Z(n4347) );
  XOR U212 ( .A(n4499), .B(sreg[1903]), .Z(n157) );
  NANDN U213 ( .A(n4500), .B(n157), .Z(n158) );
  NAND U214 ( .A(n4499), .B(sreg[1903]), .Z(n159) );
  AND U215 ( .A(n158), .B(n159), .Z(n4503) );
  NAND U216 ( .A(n4550), .B(n4551), .Z(n160) );
  XOR U217 ( .A(n4550), .B(n4551), .Z(n161) );
  NAND U218 ( .A(n161), .B(sreg[1914]), .Z(n162) );
  NAND U219 ( .A(n160), .B(n162), .Z(n4554) );
  NAND U220 ( .A(n4654), .B(sreg[1935]), .Z(n163) );
  XOR U221 ( .A(n4654), .B(sreg[1935]), .Z(n164) );
  NANDN U222 ( .A(n4653), .B(n164), .Z(n165) );
  NAND U223 ( .A(n163), .B(n165), .Z(n4656) );
  NAND U224 ( .A(sreg[1961]), .B(n4780), .Z(n166) );
  XOR U225 ( .A(sreg[1961]), .B(n4780), .Z(n167) );
  NANDN U226 ( .A(n4779), .B(n167), .Z(n168) );
  NAND U227 ( .A(n166), .B(n168), .Z(n4783) );
  XOR U228 ( .A(n4807), .B(sreg[1967]), .Z(n169) );
  NANDN U229 ( .A(n4808), .B(n169), .Z(n170) );
  NAND U230 ( .A(n4807), .B(sreg[1967]), .Z(n171) );
  AND U231 ( .A(n170), .B(n171), .Z(n4811) );
  NAND U232 ( .A(sreg[1970]), .B(n4821), .Z(n172) );
  XOR U233 ( .A(sreg[1970]), .B(n4821), .Z(n173) );
  NANDN U234 ( .A(n4820), .B(n173), .Z(n174) );
  NAND U235 ( .A(n172), .B(n174), .Z(n4824) );
  NAND U236 ( .A(n4964), .B(sreg[1999]), .Z(n175) );
  XOR U237 ( .A(n4964), .B(sreg[1999]), .Z(n176) );
  NANDN U238 ( .A(n4963), .B(n176), .Z(n177) );
  NAND U239 ( .A(n175), .B(n177), .Z(n4966) );
  NAND U240 ( .A(sreg[2002]), .B(n4977), .Z(n178) );
  XOR U241 ( .A(sreg[2002]), .B(n4977), .Z(n179) );
  NANDN U242 ( .A(n4976), .B(n179), .Z(n180) );
  NAND U243 ( .A(n178), .B(n180), .Z(n4980) );
  XOR U244 ( .A(n4989), .B(sreg[2005]), .Z(n181) );
  NANDN U245 ( .A(n4990), .B(n181), .Z(n182) );
  NAND U246 ( .A(n4989), .B(sreg[2005]), .Z(n183) );
  AND U247 ( .A(n182), .B(n183), .Z(n4993) );
  XOR U248 ( .A(n5012), .B(sreg[2010]), .Z(n184) );
  NANDN U249 ( .A(n5013), .B(n184), .Z(n185) );
  NAND U250 ( .A(n5012), .B(sreg[2010]), .Z(n186) );
  AND U251 ( .A(n185), .B(n186), .Z(n5016) );
  NAND U252 ( .A(sreg[2014]), .B(n5029), .Z(n187) );
  XOR U253 ( .A(sreg[2014]), .B(n5029), .Z(n188) );
  NANDN U254 ( .A(n5028), .B(n188), .Z(n189) );
  NAND U255 ( .A(n187), .B(n189), .Z(n5032) );
  XOR U256 ( .A(n5039), .B(sreg[2017]), .Z(n190) );
  NANDN U257 ( .A(n5040), .B(n190), .Z(n191) );
  NAND U258 ( .A(n5039), .B(sreg[2017]), .Z(n192) );
  AND U259 ( .A(n191), .B(n192), .Z(n5043) );
  NAND U260 ( .A(n5183), .B(sreg[2046]), .Z(n193) );
  XOR U261 ( .A(n5183), .B(sreg[2046]), .Z(n194) );
  NANDN U262 ( .A(n5182), .B(n194), .Z(n195) );
  NAND U263 ( .A(n193), .B(n195), .Z(c[2047]) );
  AND U264 ( .A(b[0]), .B(a[0]), .Z(n196) );
  XOR U265 ( .A(n196), .B(sreg[1023]), .Z(c[1023]) );
  AND U266 ( .A(n196), .B(sreg[1023]), .Z(n199) );
  NAND U267 ( .A(b[0]), .B(a[1]), .Z(n198) );
  XOR U268 ( .A(sreg[1024]), .B(n198), .Z(n197) );
  XNOR U269 ( .A(n199), .B(n197), .Z(c[1024]) );
  NAND U270 ( .A(b[0]), .B(a[2]), .Z(n200) );
  XNOR U271 ( .A(sreg[1025]), .B(n200), .Z(n201) );
  XOR U272 ( .A(n202), .B(n201), .Z(c[1025]) );
  NAND U273 ( .A(b[0]), .B(a[3]), .Z(n205) );
  XNOR U274 ( .A(sreg[1026]), .B(n205), .Z(n207) );
  NANDN U275 ( .A(n200), .B(sreg[1025]), .Z(n204) );
  NAND U276 ( .A(n202), .B(n201), .Z(n203) );
  NAND U277 ( .A(n204), .B(n203), .Z(n206) );
  XOR U278 ( .A(n207), .B(n206), .Z(c[1026]) );
  NANDN U279 ( .A(n205), .B(sreg[1026]), .Z(n209) );
  NAND U280 ( .A(n207), .B(n206), .Z(n208) );
  AND U281 ( .A(n209), .B(n208), .Z(n212) );
  NAND U282 ( .A(b[0]), .B(a[4]), .Z(n210) );
  XNOR U283 ( .A(sreg[1027]), .B(n210), .Z(n211) );
  XNOR U284 ( .A(n212), .B(n211), .Z(c[1027]) );
  NAND U285 ( .A(b[0]), .B(a[5]), .Z(n215) );
  XNOR U286 ( .A(sreg[1028]), .B(n215), .Z(n217) );
  NANDN U287 ( .A(sreg[1027]), .B(n210), .Z(n214) );
  NAND U288 ( .A(n212), .B(n211), .Z(n213) );
  NAND U289 ( .A(n214), .B(n213), .Z(n216) );
  XNOR U290 ( .A(n217), .B(n216), .Z(c[1028]) );
  NAND U291 ( .A(b[0]), .B(a[6]), .Z(n220) );
  XNOR U292 ( .A(sreg[1029]), .B(n220), .Z(n222) );
  NANDN U293 ( .A(sreg[1028]), .B(n215), .Z(n219) );
  NAND U294 ( .A(n217), .B(n216), .Z(n218) );
  NAND U295 ( .A(n219), .B(n218), .Z(n221) );
  XNOR U296 ( .A(n222), .B(n221), .Z(c[1029]) );
  NAND U297 ( .A(b[0]), .B(a[7]), .Z(n225) );
  XNOR U298 ( .A(sreg[1030]), .B(n225), .Z(n227) );
  NANDN U299 ( .A(sreg[1029]), .B(n220), .Z(n224) );
  NAND U300 ( .A(n222), .B(n221), .Z(n223) );
  NAND U301 ( .A(n224), .B(n223), .Z(n226) );
  XNOR U302 ( .A(n227), .B(n226), .Z(c[1030]) );
  NAND U303 ( .A(b[0]), .B(a[8]), .Z(n230) );
  XNOR U304 ( .A(sreg[1031]), .B(n230), .Z(n232) );
  NANDN U305 ( .A(sreg[1030]), .B(n225), .Z(n229) );
  NAND U306 ( .A(n227), .B(n226), .Z(n228) );
  NAND U307 ( .A(n229), .B(n228), .Z(n231) );
  XNOR U308 ( .A(n232), .B(n231), .Z(c[1031]) );
  NAND U309 ( .A(b[0]), .B(a[9]), .Z(n235) );
  XNOR U310 ( .A(sreg[1032]), .B(n235), .Z(n237) );
  NANDN U311 ( .A(sreg[1031]), .B(n230), .Z(n234) );
  NAND U312 ( .A(n232), .B(n231), .Z(n233) );
  NAND U313 ( .A(n234), .B(n233), .Z(n236) );
  XNOR U314 ( .A(n237), .B(n236), .Z(c[1032]) );
  NAND U315 ( .A(b[0]), .B(a[10]), .Z(n240) );
  XNOR U316 ( .A(sreg[1033]), .B(n240), .Z(n242) );
  NANDN U317 ( .A(sreg[1032]), .B(n235), .Z(n239) );
  NAND U318 ( .A(n237), .B(n236), .Z(n238) );
  NAND U319 ( .A(n239), .B(n238), .Z(n241) );
  XNOR U320 ( .A(n242), .B(n241), .Z(c[1033]) );
  NAND U321 ( .A(b[0]), .B(a[11]), .Z(n245) );
  XNOR U322 ( .A(sreg[1034]), .B(n245), .Z(n247) );
  NANDN U323 ( .A(sreg[1033]), .B(n240), .Z(n244) );
  NAND U324 ( .A(n242), .B(n241), .Z(n243) );
  NAND U325 ( .A(n244), .B(n243), .Z(n246) );
  XNOR U326 ( .A(n247), .B(n246), .Z(c[1034]) );
  NAND U327 ( .A(b[0]), .B(a[12]), .Z(n250) );
  XNOR U328 ( .A(sreg[1035]), .B(n250), .Z(n252) );
  NANDN U329 ( .A(sreg[1034]), .B(n245), .Z(n249) );
  NAND U330 ( .A(n247), .B(n246), .Z(n248) );
  NAND U331 ( .A(n249), .B(n248), .Z(n251) );
  XNOR U332 ( .A(n252), .B(n251), .Z(c[1035]) );
  NAND U333 ( .A(b[0]), .B(a[13]), .Z(n255) );
  XNOR U334 ( .A(sreg[1036]), .B(n255), .Z(n257) );
  NANDN U335 ( .A(sreg[1035]), .B(n250), .Z(n254) );
  NAND U336 ( .A(n252), .B(n251), .Z(n253) );
  NAND U337 ( .A(n254), .B(n253), .Z(n256) );
  XNOR U338 ( .A(n257), .B(n256), .Z(c[1036]) );
  NANDN U339 ( .A(sreg[1036]), .B(n255), .Z(n259) );
  NAND U340 ( .A(n257), .B(n256), .Z(n258) );
  AND U341 ( .A(n259), .B(n258), .Z(n262) );
  NAND U342 ( .A(b[0]), .B(a[14]), .Z(n260) );
  XNOR U343 ( .A(sreg[1037]), .B(n260), .Z(n261) );
  XOR U344 ( .A(n262), .B(n261), .Z(c[1037]) );
  NAND U345 ( .A(b[0]), .B(a[15]), .Z(n265) );
  XNOR U346 ( .A(sreg[1038]), .B(n265), .Z(n267) );
  NANDN U347 ( .A(n260), .B(sreg[1037]), .Z(n264) );
  NAND U348 ( .A(n262), .B(n261), .Z(n263) );
  AND U349 ( .A(n264), .B(n263), .Z(n266) );
  XNOR U350 ( .A(n267), .B(n266), .Z(c[1038]) );
  NANDN U351 ( .A(sreg[1038]), .B(n265), .Z(n269) );
  NAND U352 ( .A(n267), .B(n266), .Z(n268) );
  AND U353 ( .A(n269), .B(n268), .Z(n272) );
  NAND U354 ( .A(b[0]), .B(a[16]), .Z(n270) );
  XNOR U355 ( .A(sreg[1039]), .B(n270), .Z(n271) );
  XOR U356 ( .A(n272), .B(n271), .Z(c[1039]) );
  NAND U357 ( .A(b[0]), .B(a[17]), .Z(n275) );
  XNOR U358 ( .A(sreg[1040]), .B(n275), .Z(n277) );
  NANDN U359 ( .A(n270), .B(sreg[1039]), .Z(n274) );
  NAND U360 ( .A(n272), .B(n271), .Z(n273) );
  NAND U361 ( .A(n274), .B(n273), .Z(n276) );
  XOR U362 ( .A(n277), .B(n276), .Z(c[1040]) );
  NAND U363 ( .A(b[0]), .B(a[18]), .Z(n280) );
  XNOR U364 ( .A(sreg[1041]), .B(n280), .Z(n282) );
  NANDN U365 ( .A(n275), .B(sreg[1040]), .Z(n279) );
  NAND U366 ( .A(n277), .B(n276), .Z(n278) );
  NAND U367 ( .A(n279), .B(n278), .Z(n281) );
  XOR U368 ( .A(n282), .B(n281), .Z(c[1041]) );
  NAND U369 ( .A(b[0]), .B(a[19]), .Z(n285) );
  XNOR U370 ( .A(sreg[1042]), .B(n285), .Z(n287) );
  NANDN U371 ( .A(n280), .B(sreg[1041]), .Z(n284) );
  NAND U372 ( .A(n282), .B(n281), .Z(n283) );
  NAND U373 ( .A(n284), .B(n283), .Z(n286) );
  XOR U374 ( .A(n287), .B(n286), .Z(c[1042]) );
  NAND U375 ( .A(b[0]), .B(a[20]), .Z(n290) );
  XNOR U376 ( .A(sreg[1043]), .B(n290), .Z(n292) );
  NANDN U377 ( .A(n285), .B(sreg[1042]), .Z(n289) );
  NAND U378 ( .A(n287), .B(n286), .Z(n288) );
  NAND U379 ( .A(n289), .B(n288), .Z(n291) );
  XOR U380 ( .A(n292), .B(n291), .Z(c[1043]) );
  NAND U381 ( .A(b[0]), .B(a[21]), .Z(n295) );
  XNOR U382 ( .A(sreg[1044]), .B(n295), .Z(n297) );
  NANDN U383 ( .A(n290), .B(sreg[1043]), .Z(n294) );
  NAND U384 ( .A(n292), .B(n291), .Z(n293) );
  NAND U385 ( .A(n294), .B(n293), .Z(n296) );
  XOR U386 ( .A(n297), .B(n296), .Z(c[1044]) );
  NANDN U387 ( .A(n295), .B(sreg[1044]), .Z(n299) );
  NAND U388 ( .A(n297), .B(n296), .Z(n298) );
  AND U389 ( .A(n299), .B(n298), .Z(n302) );
  NAND U390 ( .A(b[0]), .B(a[22]), .Z(n300) );
  XNOR U391 ( .A(sreg[1045]), .B(n300), .Z(n301) );
  XNOR U392 ( .A(n302), .B(n301), .Z(c[1045]) );
  NAND U393 ( .A(b[0]), .B(a[23]), .Z(n305) );
  XNOR U394 ( .A(sreg[1046]), .B(n305), .Z(n307) );
  NANDN U395 ( .A(sreg[1045]), .B(n300), .Z(n304) );
  NAND U396 ( .A(n302), .B(n301), .Z(n303) );
  NAND U397 ( .A(n304), .B(n303), .Z(n306) );
  XNOR U398 ( .A(n307), .B(n306), .Z(c[1046]) );
  NAND U399 ( .A(b[0]), .B(a[24]), .Z(n310) );
  XNOR U400 ( .A(sreg[1047]), .B(n310), .Z(n312) );
  NANDN U401 ( .A(sreg[1046]), .B(n305), .Z(n309) );
  NAND U402 ( .A(n307), .B(n306), .Z(n308) );
  AND U403 ( .A(n309), .B(n308), .Z(n311) );
  XOR U404 ( .A(n312), .B(n311), .Z(c[1047]) );
  NAND U405 ( .A(b[0]), .B(a[25]), .Z(n315) );
  XNOR U406 ( .A(sreg[1048]), .B(n315), .Z(n317) );
  NANDN U407 ( .A(n310), .B(sreg[1047]), .Z(n314) );
  NAND U408 ( .A(n312), .B(n311), .Z(n313) );
  AND U409 ( .A(n314), .B(n313), .Z(n316) );
  XNOR U410 ( .A(n317), .B(n316), .Z(c[1048]) );
  NAND U411 ( .A(b[0]), .B(a[26]), .Z(n320) );
  XNOR U412 ( .A(sreg[1049]), .B(n320), .Z(n322) );
  NANDN U413 ( .A(sreg[1048]), .B(n315), .Z(n319) );
  NAND U414 ( .A(n317), .B(n316), .Z(n318) );
  NAND U415 ( .A(n319), .B(n318), .Z(n321) );
  XNOR U416 ( .A(n322), .B(n321), .Z(c[1049]) );
  NANDN U417 ( .A(sreg[1049]), .B(n320), .Z(n324) );
  NAND U418 ( .A(n322), .B(n321), .Z(n323) );
  AND U419 ( .A(n324), .B(n323), .Z(n327) );
  NAND U420 ( .A(b[0]), .B(a[27]), .Z(n325) );
  XNOR U421 ( .A(sreg[1050]), .B(n325), .Z(n326) );
  XOR U422 ( .A(n327), .B(n326), .Z(c[1050]) );
  NANDN U423 ( .A(n325), .B(sreg[1050]), .Z(n329) );
  NAND U424 ( .A(n327), .B(n326), .Z(n328) );
  AND U425 ( .A(n329), .B(n328), .Z(n332) );
  NAND U426 ( .A(b[0]), .B(a[28]), .Z(n330) );
  XNOR U427 ( .A(sreg[1051]), .B(n330), .Z(n331) );
  XNOR U428 ( .A(n332), .B(n331), .Z(c[1051]) );
  NAND U429 ( .A(b[0]), .B(a[29]), .Z(n335) );
  XNOR U430 ( .A(sreg[1052]), .B(n335), .Z(n337) );
  NANDN U431 ( .A(sreg[1051]), .B(n330), .Z(n334) );
  NAND U432 ( .A(n332), .B(n331), .Z(n333) );
  AND U433 ( .A(n334), .B(n333), .Z(n336) );
  XOR U434 ( .A(n337), .B(n336), .Z(c[1052]) );
  NAND U435 ( .A(b[0]), .B(a[30]), .Z(n340) );
  XNOR U436 ( .A(sreg[1053]), .B(n340), .Z(n342) );
  NANDN U437 ( .A(n335), .B(sreg[1052]), .Z(n339) );
  NAND U438 ( .A(n337), .B(n336), .Z(n338) );
  NAND U439 ( .A(n339), .B(n338), .Z(n341) );
  XOR U440 ( .A(n342), .B(n341), .Z(c[1053]) );
  NAND U441 ( .A(b[0]), .B(a[31]), .Z(n345) );
  XNOR U442 ( .A(sreg[1054]), .B(n345), .Z(n347) );
  NANDN U443 ( .A(n340), .B(sreg[1053]), .Z(n344) );
  NAND U444 ( .A(n342), .B(n341), .Z(n343) );
  AND U445 ( .A(n344), .B(n343), .Z(n346) );
  XNOR U446 ( .A(n347), .B(n346), .Z(c[1054]) );
  NAND U447 ( .A(b[0]), .B(a[32]), .Z(n350) );
  XNOR U448 ( .A(sreg[1055]), .B(n350), .Z(n352) );
  NANDN U449 ( .A(sreg[1054]), .B(n345), .Z(n349) );
  NAND U450 ( .A(n347), .B(n346), .Z(n348) );
  NAND U451 ( .A(n349), .B(n348), .Z(n351) );
  XNOR U452 ( .A(n352), .B(n351), .Z(c[1055]) );
  NAND U453 ( .A(b[0]), .B(a[33]), .Z(n355) );
  XNOR U454 ( .A(sreg[1056]), .B(n355), .Z(n357) );
  NANDN U455 ( .A(sreg[1055]), .B(n350), .Z(n354) );
  NAND U456 ( .A(n352), .B(n351), .Z(n353) );
  AND U457 ( .A(n354), .B(n353), .Z(n356) );
  XOR U458 ( .A(n357), .B(n356), .Z(c[1056]) );
  NANDN U459 ( .A(n355), .B(sreg[1056]), .Z(n359) );
  NAND U460 ( .A(n357), .B(n356), .Z(n358) );
  AND U461 ( .A(n359), .B(n358), .Z(n362) );
  NAND U462 ( .A(b[0]), .B(a[34]), .Z(n360) );
  XNOR U463 ( .A(sreg[1057]), .B(n360), .Z(n361) );
  XNOR U464 ( .A(n362), .B(n361), .Z(c[1057]) );
  NAND U465 ( .A(b[0]), .B(a[35]), .Z(n365) );
  XNOR U466 ( .A(sreg[1058]), .B(n365), .Z(n367) );
  NANDN U467 ( .A(sreg[1057]), .B(n360), .Z(n364) );
  NAND U468 ( .A(n362), .B(n361), .Z(n363) );
  NAND U469 ( .A(n364), .B(n363), .Z(n366) );
  XNOR U470 ( .A(n367), .B(n366), .Z(c[1058]) );
  NAND U471 ( .A(b[0]), .B(a[36]), .Z(n370) );
  XNOR U472 ( .A(sreg[1059]), .B(n370), .Z(n372) );
  NANDN U473 ( .A(sreg[1058]), .B(n365), .Z(n369) );
  NAND U474 ( .A(n367), .B(n366), .Z(n368) );
  AND U475 ( .A(n369), .B(n368), .Z(n371) );
  XOR U476 ( .A(n372), .B(n371), .Z(c[1059]) );
  NAND U477 ( .A(b[0]), .B(a[37]), .Z(n375) );
  XNOR U478 ( .A(sreg[1060]), .B(n375), .Z(n377) );
  NANDN U479 ( .A(n370), .B(sreg[1059]), .Z(n374) );
  NAND U480 ( .A(n372), .B(n371), .Z(n373) );
  AND U481 ( .A(n374), .B(n373), .Z(n376) );
  XNOR U482 ( .A(n377), .B(n376), .Z(c[1060]) );
  NAND U483 ( .A(b[0]), .B(a[38]), .Z(n380) );
  XNOR U484 ( .A(sreg[1061]), .B(n380), .Z(n382) );
  NANDN U485 ( .A(sreg[1060]), .B(n375), .Z(n379) );
  NAND U486 ( .A(n377), .B(n376), .Z(n378) );
  NAND U487 ( .A(n379), .B(n378), .Z(n381) );
  XNOR U488 ( .A(n382), .B(n381), .Z(c[1061]) );
  NAND U489 ( .A(b[0]), .B(a[39]), .Z(n385) );
  XNOR U490 ( .A(sreg[1062]), .B(n385), .Z(n387) );
  NANDN U491 ( .A(sreg[1061]), .B(n380), .Z(n384) );
  NAND U492 ( .A(n382), .B(n381), .Z(n383) );
  AND U493 ( .A(n384), .B(n383), .Z(n386) );
  XOR U494 ( .A(n387), .B(n386), .Z(c[1062]) );
  NANDN U495 ( .A(n385), .B(sreg[1062]), .Z(n389) );
  NAND U496 ( .A(n387), .B(n386), .Z(n388) );
  AND U497 ( .A(n389), .B(n388), .Z(n392) );
  NAND U498 ( .A(b[0]), .B(a[40]), .Z(n390) );
  XNOR U499 ( .A(sreg[1063]), .B(n390), .Z(n391) );
  XNOR U500 ( .A(n392), .B(n391), .Z(c[1063]) );
  NAND U501 ( .A(b[0]), .B(a[41]), .Z(n395) );
  XNOR U502 ( .A(sreg[1064]), .B(n395), .Z(n397) );
  NANDN U503 ( .A(sreg[1063]), .B(n390), .Z(n394) );
  NAND U504 ( .A(n392), .B(n391), .Z(n393) );
  NAND U505 ( .A(n394), .B(n393), .Z(n396) );
  XNOR U506 ( .A(n397), .B(n396), .Z(c[1064]) );
  NAND U507 ( .A(b[0]), .B(a[42]), .Z(n400) );
  XNOR U508 ( .A(sreg[1065]), .B(n400), .Z(n402) );
  NANDN U509 ( .A(sreg[1064]), .B(n395), .Z(n399) );
  NAND U510 ( .A(n397), .B(n396), .Z(n398) );
  AND U511 ( .A(n399), .B(n398), .Z(n401) );
  XOR U512 ( .A(n402), .B(n401), .Z(c[1065]) );
  NANDN U513 ( .A(n400), .B(sreg[1065]), .Z(n404) );
  NAND U514 ( .A(n402), .B(n401), .Z(n403) );
  AND U515 ( .A(n404), .B(n403), .Z(n407) );
  NAND U516 ( .A(b[0]), .B(a[43]), .Z(n405) );
  XNOR U517 ( .A(sreg[1066]), .B(n405), .Z(n406) );
  XNOR U518 ( .A(n407), .B(n406), .Z(c[1066]) );
  NAND U519 ( .A(b[0]), .B(a[44]), .Z(n410) );
  XNOR U520 ( .A(sreg[1067]), .B(n410), .Z(n412) );
  NANDN U521 ( .A(sreg[1066]), .B(n405), .Z(n409) );
  NAND U522 ( .A(n407), .B(n406), .Z(n408) );
  NAND U523 ( .A(n409), .B(n408), .Z(n411) );
  XNOR U524 ( .A(n412), .B(n411), .Z(c[1067]) );
  NANDN U525 ( .A(sreg[1067]), .B(n410), .Z(n414) );
  NAND U526 ( .A(n412), .B(n411), .Z(n413) );
  AND U527 ( .A(n414), .B(n413), .Z(n417) );
  NAND U528 ( .A(b[0]), .B(a[45]), .Z(n415) );
  XNOR U529 ( .A(sreg[1068]), .B(n415), .Z(n416) );
  XOR U530 ( .A(n417), .B(n416), .Z(c[1068]) );
  NANDN U531 ( .A(n415), .B(sreg[1068]), .Z(n419) );
  NAND U532 ( .A(n417), .B(n416), .Z(n418) );
  AND U533 ( .A(n419), .B(n418), .Z(n421) );
  AND U534 ( .A(b[0]), .B(a[46]), .Z(n422) );
  XNOR U535 ( .A(sreg[1069]), .B(n422), .Z(n420) );
  XOR U536 ( .A(n421), .B(n420), .Z(c[1069]) );
  NAND U537 ( .A(b[0]), .B(a[47]), .Z(n423) );
  XNOR U538 ( .A(sreg[1070]), .B(n423), .Z(n425) );
  XOR U539 ( .A(n425), .B(n424), .Z(c[1070]) );
  NAND U540 ( .A(b[0]), .B(a[48]), .Z(n430) );
  NANDN U541 ( .A(n423), .B(sreg[1070]), .Z(n427) );
  NAND U542 ( .A(n425), .B(n424), .Z(n426) );
  NAND U543 ( .A(n427), .B(n426), .Z(n429) );
  XOR U544 ( .A(n429), .B(sreg[1071]), .Z(n428) );
  XNOR U545 ( .A(n430), .B(n428), .Z(c[1071]) );
  NAND U546 ( .A(b[0]), .B(a[49]), .Z(n431) );
  XNOR U547 ( .A(sreg[1072]), .B(n431), .Z(n432) );
  XNOR U548 ( .A(n433), .B(n432), .Z(c[1072]) );
  NAND U549 ( .A(b[0]), .B(a[50]), .Z(n436) );
  XNOR U550 ( .A(sreg[1073]), .B(n436), .Z(n438) );
  NANDN U551 ( .A(n431), .B(sreg[1072]), .Z(n435) );
  NANDN U552 ( .A(n433), .B(n432), .Z(n434) );
  NAND U553 ( .A(n435), .B(n434), .Z(n437) );
  XOR U554 ( .A(n438), .B(n437), .Z(c[1073]) );
  NANDN U555 ( .A(n436), .B(sreg[1073]), .Z(n440) );
  NAND U556 ( .A(n438), .B(n437), .Z(n439) );
  NAND U557 ( .A(n440), .B(n439), .Z(n443) );
  NAND U558 ( .A(b[0]), .B(a[51]), .Z(n442) );
  XOR U559 ( .A(sreg[1074]), .B(n442), .Z(n441) );
  XNOR U560 ( .A(n443), .B(n441), .Z(c[1074]) );
  NAND U561 ( .A(b[0]), .B(a[52]), .Z(n444) );
  XNOR U562 ( .A(sreg[1075]), .B(n444), .Z(n445) );
  XOR U563 ( .A(n446), .B(n445), .Z(c[1075]) );
  NAND U564 ( .A(b[0]), .B(a[53]), .Z(n449) );
  XNOR U565 ( .A(sreg[1076]), .B(n449), .Z(n451) );
  NANDN U566 ( .A(n444), .B(sreg[1075]), .Z(n448) );
  NAND U567 ( .A(n446), .B(n445), .Z(n447) );
  NAND U568 ( .A(n448), .B(n447), .Z(n450) );
  XOR U569 ( .A(n451), .B(n450), .Z(c[1076]) );
  AND U570 ( .A(b[0]), .B(a[54]), .Z(n455) );
  NANDN U571 ( .A(n449), .B(sreg[1076]), .Z(n453) );
  NAND U572 ( .A(n451), .B(n450), .Z(n452) );
  AND U573 ( .A(n453), .B(n452), .Z(n456) );
  XNOR U574 ( .A(sreg[1077]), .B(n456), .Z(n454) );
  XOR U575 ( .A(n455), .B(n454), .Z(c[1077]) );
  NAND U576 ( .A(b[0]), .B(a[55]), .Z(n457) );
  XNOR U577 ( .A(sreg[1078]), .B(n457), .Z(n458) );
  XNOR U578 ( .A(n459), .B(n458), .Z(c[1078]) );
  NAND U579 ( .A(b[0]), .B(a[56]), .Z(n462) );
  XNOR U580 ( .A(sreg[1079]), .B(n462), .Z(n464) );
  NANDN U581 ( .A(sreg[1078]), .B(n457), .Z(n461) );
  NAND U582 ( .A(n459), .B(n458), .Z(n460) );
  AND U583 ( .A(n461), .B(n460), .Z(n463) );
  XOR U584 ( .A(n464), .B(n463), .Z(c[1079]) );
  NANDN U585 ( .A(n462), .B(sreg[1079]), .Z(n466) );
  NAND U586 ( .A(n464), .B(n463), .Z(n465) );
  NAND U587 ( .A(n466), .B(n465), .Z(n469) );
  NAND U588 ( .A(b[0]), .B(a[57]), .Z(n468) );
  XOR U589 ( .A(sreg[1080]), .B(n468), .Z(n467) );
  XNOR U590 ( .A(n469), .B(n467), .Z(c[1080]) );
  NAND U591 ( .A(b[0]), .B(a[58]), .Z(n470) );
  XNOR U592 ( .A(sreg[1081]), .B(n470), .Z(n471) );
  XOR U593 ( .A(n472), .B(n471), .Z(c[1081]) );
  NANDN U594 ( .A(sreg[1081]), .B(n470), .Z(n474) );
  NANDN U595 ( .A(n472), .B(n471), .Z(n473) );
  AND U596 ( .A(n474), .B(n473), .Z(n477) );
  NAND U597 ( .A(b[0]), .B(a[59]), .Z(n475) );
  XNOR U598 ( .A(sreg[1082]), .B(n475), .Z(n476) );
  XOR U599 ( .A(n477), .B(n476), .Z(c[1082]) );
  NANDN U600 ( .A(n475), .B(sreg[1082]), .Z(n479) );
  NAND U601 ( .A(n477), .B(n476), .Z(n478) );
  AND U602 ( .A(n479), .B(n478), .Z(n482) );
  NAND U603 ( .A(b[0]), .B(a[60]), .Z(n480) );
  XNOR U604 ( .A(sreg[1083]), .B(n480), .Z(n481) );
  XNOR U605 ( .A(n482), .B(n481), .Z(c[1083]) );
  NANDN U606 ( .A(sreg[1083]), .B(n480), .Z(n484) );
  NAND U607 ( .A(n482), .B(n481), .Z(n483) );
  AND U608 ( .A(n484), .B(n483), .Z(n487) );
  NAND U609 ( .A(b[0]), .B(a[61]), .Z(n485) );
  XNOR U610 ( .A(sreg[1084]), .B(n485), .Z(n486) );
  XOR U611 ( .A(n487), .B(n486), .Z(c[1084]) );
  NAND U612 ( .A(b[0]), .B(a[62]), .Z(n490) );
  XNOR U613 ( .A(sreg[1085]), .B(n490), .Z(n492) );
  NANDN U614 ( .A(n485), .B(sreg[1084]), .Z(n489) );
  NAND U615 ( .A(n487), .B(n486), .Z(n488) );
  NAND U616 ( .A(n489), .B(n488), .Z(n491) );
  XOR U617 ( .A(n492), .B(n491), .Z(c[1085]) );
  NAND U618 ( .A(b[0]), .B(a[63]), .Z(n495) );
  XNOR U619 ( .A(sreg[1086]), .B(n495), .Z(n497) );
  NANDN U620 ( .A(n490), .B(sreg[1085]), .Z(n494) );
  NAND U621 ( .A(n492), .B(n491), .Z(n493) );
  AND U622 ( .A(n494), .B(n493), .Z(n496) );
  XNOR U623 ( .A(n497), .B(n496), .Z(c[1086]) );
  NANDN U624 ( .A(sreg[1086]), .B(n495), .Z(n499) );
  NAND U625 ( .A(n497), .B(n496), .Z(n498) );
  AND U626 ( .A(n499), .B(n498), .Z(n502) );
  NAND U627 ( .A(b[0]), .B(a[64]), .Z(n500) );
  XNOR U628 ( .A(sreg[1087]), .B(n500), .Z(n501) );
  XOR U629 ( .A(n502), .B(n501), .Z(c[1087]) );
  NAND U630 ( .A(b[0]), .B(a[65]), .Z(n505) );
  XNOR U631 ( .A(sreg[1088]), .B(n505), .Z(n507) );
  NANDN U632 ( .A(n500), .B(sreg[1087]), .Z(n504) );
  NAND U633 ( .A(n502), .B(n501), .Z(n503) );
  NAND U634 ( .A(n504), .B(n503), .Z(n506) );
  XOR U635 ( .A(n507), .B(n506), .Z(c[1088]) );
  NAND U636 ( .A(b[0]), .B(a[66]), .Z(n510) );
  XNOR U637 ( .A(sreg[1089]), .B(n510), .Z(n512) );
  NANDN U638 ( .A(n505), .B(sreg[1088]), .Z(n509) );
  NAND U639 ( .A(n507), .B(n506), .Z(n508) );
  AND U640 ( .A(n509), .B(n508), .Z(n511) );
  XNOR U641 ( .A(n512), .B(n511), .Z(c[1089]) );
  NAND U642 ( .A(b[0]), .B(a[67]), .Z(n515) );
  XNOR U643 ( .A(sreg[1090]), .B(n515), .Z(n517) );
  NANDN U644 ( .A(sreg[1089]), .B(n510), .Z(n514) );
  NAND U645 ( .A(n512), .B(n511), .Z(n513) );
  AND U646 ( .A(n514), .B(n513), .Z(n516) );
  XOR U647 ( .A(n517), .B(n516), .Z(c[1090]) );
  NAND U648 ( .A(b[0]), .B(a[68]), .Z(n520) );
  XNOR U649 ( .A(sreg[1091]), .B(n520), .Z(n522) );
  NANDN U650 ( .A(n515), .B(sreg[1090]), .Z(n519) );
  NAND U651 ( .A(n517), .B(n516), .Z(n518) );
  NAND U652 ( .A(n519), .B(n518), .Z(n521) );
  XOR U653 ( .A(n522), .B(n521), .Z(c[1091]) );
  NANDN U654 ( .A(n520), .B(sreg[1091]), .Z(n524) );
  NAND U655 ( .A(n522), .B(n521), .Z(n523) );
  AND U656 ( .A(n524), .B(n523), .Z(n527) );
  NAND U657 ( .A(b[0]), .B(a[69]), .Z(n525) );
  XNOR U658 ( .A(sreg[1092]), .B(n525), .Z(n526) );
  XNOR U659 ( .A(n527), .B(n526), .Z(c[1092]) );
  NAND U660 ( .A(b[0]), .B(a[70]), .Z(n530) );
  XNOR U661 ( .A(sreg[1093]), .B(n530), .Z(n532) );
  NANDN U662 ( .A(sreg[1092]), .B(n525), .Z(n529) );
  NAND U663 ( .A(n527), .B(n526), .Z(n528) );
  NAND U664 ( .A(n529), .B(n528), .Z(n531) );
  XNOR U665 ( .A(n532), .B(n531), .Z(c[1093]) );
  NAND U666 ( .A(b[0]), .B(a[71]), .Z(n535) );
  XNOR U667 ( .A(sreg[1094]), .B(n535), .Z(n537) );
  NANDN U668 ( .A(sreg[1093]), .B(n530), .Z(n534) );
  NAND U669 ( .A(n532), .B(n531), .Z(n533) );
  NAND U670 ( .A(n534), .B(n533), .Z(n536) );
  XNOR U671 ( .A(n537), .B(n536), .Z(c[1094]) );
  NAND U672 ( .A(b[0]), .B(a[72]), .Z(n540) );
  XNOR U673 ( .A(sreg[1095]), .B(n540), .Z(n542) );
  NANDN U674 ( .A(sreg[1094]), .B(n535), .Z(n539) );
  NAND U675 ( .A(n537), .B(n536), .Z(n538) );
  NAND U676 ( .A(n539), .B(n538), .Z(n541) );
  XNOR U677 ( .A(n542), .B(n541), .Z(c[1095]) );
  NAND U678 ( .A(b[0]), .B(a[73]), .Z(n545) );
  XNOR U679 ( .A(sreg[1096]), .B(n545), .Z(n547) );
  NANDN U680 ( .A(sreg[1095]), .B(n540), .Z(n544) );
  NAND U681 ( .A(n542), .B(n541), .Z(n543) );
  NAND U682 ( .A(n544), .B(n543), .Z(n546) );
  XNOR U683 ( .A(n547), .B(n546), .Z(c[1096]) );
  NAND U684 ( .A(b[0]), .B(a[74]), .Z(n550) );
  XNOR U685 ( .A(sreg[1097]), .B(n550), .Z(n552) );
  NANDN U686 ( .A(sreg[1096]), .B(n545), .Z(n549) );
  NAND U687 ( .A(n547), .B(n546), .Z(n548) );
  NAND U688 ( .A(n549), .B(n548), .Z(n551) );
  XNOR U689 ( .A(n552), .B(n551), .Z(c[1097]) );
  NAND U690 ( .A(b[0]), .B(a[75]), .Z(n555) );
  XNOR U691 ( .A(sreg[1098]), .B(n555), .Z(n557) );
  NANDN U692 ( .A(sreg[1097]), .B(n550), .Z(n554) );
  NAND U693 ( .A(n552), .B(n551), .Z(n553) );
  NAND U694 ( .A(n554), .B(n553), .Z(n556) );
  XNOR U695 ( .A(n557), .B(n556), .Z(c[1098]) );
  NANDN U696 ( .A(sreg[1098]), .B(n555), .Z(n559) );
  NAND U697 ( .A(n557), .B(n556), .Z(n558) );
  AND U698 ( .A(n559), .B(n558), .Z(n562) );
  NAND U699 ( .A(b[0]), .B(a[76]), .Z(n560) );
  XNOR U700 ( .A(sreg[1099]), .B(n560), .Z(n561) );
  XOR U701 ( .A(n562), .B(n561), .Z(c[1099]) );
  NANDN U702 ( .A(n560), .B(sreg[1099]), .Z(n564) );
  NAND U703 ( .A(n562), .B(n561), .Z(n563) );
  AND U704 ( .A(n564), .B(n563), .Z(n567) );
  NAND U705 ( .A(b[0]), .B(a[77]), .Z(n565) );
  XNOR U706 ( .A(sreg[1100]), .B(n565), .Z(n566) );
  XNOR U707 ( .A(n567), .B(n566), .Z(c[1100]) );
  NANDN U708 ( .A(sreg[1100]), .B(n565), .Z(n569) );
  NAND U709 ( .A(n567), .B(n566), .Z(n568) );
  AND U710 ( .A(n569), .B(n568), .Z(n572) );
  NAND U711 ( .A(b[0]), .B(a[78]), .Z(n570) );
  XNOR U712 ( .A(sreg[1101]), .B(n570), .Z(n571) );
  XOR U713 ( .A(n572), .B(n571), .Z(c[1101]) );
  NAND U714 ( .A(b[0]), .B(a[79]), .Z(n575) );
  XNOR U715 ( .A(sreg[1102]), .B(n575), .Z(n577) );
  NANDN U716 ( .A(n570), .B(sreg[1101]), .Z(n574) );
  NAND U717 ( .A(n572), .B(n571), .Z(n573) );
  NAND U718 ( .A(n574), .B(n573), .Z(n576) );
  XOR U719 ( .A(n577), .B(n576), .Z(c[1102]) );
  NAND U720 ( .A(b[0]), .B(a[80]), .Z(n580) );
  XNOR U721 ( .A(sreg[1103]), .B(n580), .Z(n582) );
  NANDN U722 ( .A(n575), .B(sreg[1102]), .Z(n579) );
  NAND U723 ( .A(n577), .B(n576), .Z(n578) );
  NAND U724 ( .A(n579), .B(n578), .Z(n581) );
  XOR U725 ( .A(n582), .B(n581), .Z(c[1103]) );
  NAND U726 ( .A(b[0]), .B(a[81]), .Z(n585) );
  XNOR U727 ( .A(sreg[1104]), .B(n585), .Z(n587) );
  NANDN U728 ( .A(n580), .B(sreg[1103]), .Z(n584) );
  NAND U729 ( .A(n582), .B(n581), .Z(n583) );
  NAND U730 ( .A(n584), .B(n583), .Z(n586) );
  XOR U731 ( .A(n587), .B(n586), .Z(c[1104]) );
  NAND U732 ( .A(b[0]), .B(a[82]), .Z(n590) );
  XNOR U733 ( .A(sreg[1105]), .B(n590), .Z(n592) );
  NANDN U734 ( .A(n585), .B(sreg[1104]), .Z(n589) );
  NAND U735 ( .A(n587), .B(n586), .Z(n588) );
  NAND U736 ( .A(n589), .B(n588), .Z(n591) );
  XOR U737 ( .A(n592), .B(n591), .Z(c[1105]) );
  NAND U738 ( .A(b[0]), .B(a[83]), .Z(n595) );
  XNOR U739 ( .A(sreg[1106]), .B(n595), .Z(n597) );
  NANDN U740 ( .A(n590), .B(sreg[1105]), .Z(n594) );
  NAND U741 ( .A(n592), .B(n591), .Z(n593) );
  NAND U742 ( .A(n594), .B(n593), .Z(n596) );
  XOR U743 ( .A(n597), .B(n596), .Z(c[1106]) );
  NAND U744 ( .A(b[0]), .B(a[84]), .Z(n600) );
  XNOR U745 ( .A(sreg[1107]), .B(n600), .Z(n602) );
  NANDN U746 ( .A(n595), .B(sreg[1106]), .Z(n599) );
  NAND U747 ( .A(n597), .B(n596), .Z(n598) );
  NAND U748 ( .A(n599), .B(n598), .Z(n601) );
  XOR U749 ( .A(n602), .B(n601), .Z(c[1107]) );
  NANDN U750 ( .A(n600), .B(sreg[1107]), .Z(n604) );
  NAND U751 ( .A(n602), .B(n601), .Z(n603) );
  AND U752 ( .A(n604), .B(n603), .Z(n607) );
  NAND U753 ( .A(b[0]), .B(a[85]), .Z(n605) );
  XNOR U754 ( .A(sreg[1108]), .B(n605), .Z(n606) );
  XNOR U755 ( .A(n607), .B(n606), .Z(c[1108]) );
  NAND U756 ( .A(b[0]), .B(a[86]), .Z(n610) );
  XNOR U757 ( .A(sreg[1109]), .B(n610), .Z(n612) );
  NANDN U758 ( .A(sreg[1108]), .B(n605), .Z(n609) );
  NAND U759 ( .A(n607), .B(n606), .Z(n608) );
  AND U760 ( .A(n609), .B(n608), .Z(n611) );
  XOR U761 ( .A(n612), .B(n611), .Z(c[1109]) );
  NAND U762 ( .A(b[0]), .B(a[87]), .Z(n615) );
  XNOR U763 ( .A(sreg[1110]), .B(n615), .Z(n617) );
  NANDN U764 ( .A(n610), .B(sreg[1109]), .Z(n614) );
  NAND U765 ( .A(n612), .B(n611), .Z(n613) );
  NAND U766 ( .A(n614), .B(n613), .Z(n616) );
  XOR U767 ( .A(n617), .B(n616), .Z(c[1110]) );
  AND U768 ( .A(b[0]), .B(a[88]), .Z(n621) );
  NANDN U769 ( .A(n615), .B(sreg[1110]), .Z(n619) );
  NAND U770 ( .A(n617), .B(n616), .Z(n618) );
  AND U771 ( .A(n619), .B(n618), .Z(n622) );
  XNOR U772 ( .A(sreg[1111]), .B(n622), .Z(n620) );
  XOR U773 ( .A(n621), .B(n620), .Z(c[1111]) );
  NAND U774 ( .A(b[0]), .B(a[89]), .Z(n623) );
  XNOR U775 ( .A(sreg[1112]), .B(n623), .Z(n624) );
  XNOR U776 ( .A(n625), .B(n624), .Z(c[1112]) );
  NAND U777 ( .A(b[0]), .B(a[90]), .Z(n630) );
  NANDN U778 ( .A(n623), .B(sreg[1112]), .Z(n627) );
  NANDN U779 ( .A(n625), .B(n624), .Z(n626) );
  NAND U780 ( .A(n627), .B(n626), .Z(n629) );
  XOR U781 ( .A(n629), .B(sreg[1113]), .Z(n628) );
  XNOR U782 ( .A(n630), .B(n628), .Z(c[1113]) );
  NAND U783 ( .A(b[0]), .B(a[91]), .Z(n631) );
  XNOR U784 ( .A(sreg[1114]), .B(n631), .Z(n632) );
  XNOR U785 ( .A(n633), .B(n632), .Z(c[1114]) );
  NAND U786 ( .A(b[0]), .B(a[92]), .Z(n636) );
  XNOR U787 ( .A(sreg[1115]), .B(n636), .Z(n638) );
  NANDN U788 ( .A(n631), .B(sreg[1114]), .Z(n635) );
  NANDN U789 ( .A(n633), .B(n632), .Z(n634) );
  NAND U790 ( .A(n635), .B(n634), .Z(n637) );
  XOR U791 ( .A(n638), .B(n637), .Z(c[1115]) );
  NAND U792 ( .A(b[0]), .B(a[93]), .Z(n641) );
  XNOR U793 ( .A(sreg[1116]), .B(n641), .Z(n643) );
  NANDN U794 ( .A(n636), .B(sreg[1115]), .Z(n640) );
  NAND U795 ( .A(n638), .B(n637), .Z(n639) );
  AND U796 ( .A(n640), .B(n639), .Z(n642) );
  XNOR U797 ( .A(n643), .B(n642), .Z(c[1116]) );
  NANDN U798 ( .A(sreg[1116]), .B(n641), .Z(n645) );
  NAND U799 ( .A(n643), .B(n642), .Z(n644) );
  AND U800 ( .A(n645), .B(n644), .Z(n648) );
  NAND U801 ( .A(b[0]), .B(a[94]), .Z(n646) );
  XNOR U802 ( .A(sreg[1117]), .B(n646), .Z(n647) );
  XOR U803 ( .A(n648), .B(n647), .Z(c[1117]) );
  NAND U804 ( .A(b[0]), .B(a[95]), .Z(n651) );
  XNOR U805 ( .A(sreg[1118]), .B(n651), .Z(n653) );
  NANDN U806 ( .A(n646), .B(sreg[1117]), .Z(n650) );
  NAND U807 ( .A(n648), .B(n647), .Z(n649) );
  NAND U808 ( .A(n650), .B(n649), .Z(n652) );
  XOR U809 ( .A(n653), .B(n652), .Z(c[1118]) );
  NAND U810 ( .A(b[0]), .B(a[96]), .Z(n656) );
  XNOR U811 ( .A(sreg[1119]), .B(n656), .Z(n658) );
  NANDN U812 ( .A(n651), .B(sreg[1118]), .Z(n655) );
  NAND U813 ( .A(n653), .B(n652), .Z(n654) );
  NAND U814 ( .A(n655), .B(n654), .Z(n657) );
  XOR U815 ( .A(n658), .B(n657), .Z(c[1119]) );
  NAND U816 ( .A(b[0]), .B(a[97]), .Z(n661) );
  XNOR U817 ( .A(sreg[1120]), .B(n661), .Z(n663) );
  NANDN U818 ( .A(n656), .B(sreg[1119]), .Z(n660) );
  NAND U819 ( .A(n658), .B(n657), .Z(n659) );
  NAND U820 ( .A(n660), .B(n659), .Z(n662) );
  XOR U821 ( .A(n663), .B(n662), .Z(c[1120]) );
  NAND U822 ( .A(b[0]), .B(a[98]), .Z(n666) );
  XNOR U823 ( .A(sreg[1121]), .B(n666), .Z(n668) );
  NANDN U824 ( .A(n661), .B(sreg[1120]), .Z(n665) );
  NAND U825 ( .A(n663), .B(n662), .Z(n664) );
  NAND U826 ( .A(n665), .B(n664), .Z(n667) );
  XOR U827 ( .A(n668), .B(n667), .Z(c[1121]) );
  NAND U828 ( .A(b[0]), .B(a[99]), .Z(n671) );
  XNOR U829 ( .A(sreg[1122]), .B(n671), .Z(n673) );
  NANDN U830 ( .A(n666), .B(sreg[1121]), .Z(n670) );
  NAND U831 ( .A(n668), .B(n667), .Z(n669) );
  NAND U832 ( .A(n670), .B(n669), .Z(n672) );
  XOR U833 ( .A(n673), .B(n672), .Z(c[1122]) );
  NANDN U834 ( .A(n671), .B(sreg[1122]), .Z(n675) );
  NAND U835 ( .A(n673), .B(n672), .Z(n674) );
  AND U836 ( .A(n675), .B(n674), .Z(n678) );
  NAND U837 ( .A(b[0]), .B(a[100]), .Z(n676) );
  XNOR U838 ( .A(sreg[1123]), .B(n676), .Z(n677) );
  XNOR U839 ( .A(n678), .B(n677), .Z(c[1123]) );
  NAND U840 ( .A(b[0]), .B(a[101]), .Z(n681) );
  XNOR U841 ( .A(sreg[1124]), .B(n681), .Z(n683) );
  NANDN U842 ( .A(sreg[1123]), .B(n676), .Z(n680) );
  NAND U843 ( .A(n678), .B(n677), .Z(n679) );
  AND U844 ( .A(n680), .B(n679), .Z(n682) );
  XOR U845 ( .A(n683), .B(n682), .Z(c[1124]) );
  NANDN U846 ( .A(n681), .B(sreg[1124]), .Z(n685) );
  NAND U847 ( .A(n683), .B(n682), .Z(n684) );
  AND U848 ( .A(n685), .B(n684), .Z(n688) );
  NAND U849 ( .A(b[0]), .B(a[102]), .Z(n686) );
  XNOR U850 ( .A(sreg[1125]), .B(n686), .Z(n687) );
  XNOR U851 ( .A(n688), .B(n687), .Z(c[1125]) );
  NAND U852 ( .A(b[0]), .B(a[103]), .Z(n691) );
  XNOR U853 ( .A(sreg[1126]), .B(n691), .Z(n693) );
  NANDN U854 ( .A(sreg[1125]), .B(n686), .Z(n690) );
  NAND U855 ( .A(n688), .B(n687), .Z(n689) );
  NAND U856 ( .A(n690), .B(n689), .Z(n692) );
  XNOR U857 ( .A(n693), .B(n692), .Z(c[1126]) );
  NAND U858 ( .A(b[0]), .B(a[104]), .Z(n696) );
  XNOR U859 ( .A(sreg[1127]), .B(n696), .Z(n698) );
  NANDN U860 ( .A(sreg[1126]), .B(n691), .Z(n695) );
  NAND U861 ( .A(n693), .B(n692), .Z(n694) );
  AND U862 ( .A(n695), .B(n694), .Z(n697) );
  XOR U863 ( .A(n698), .B(n697), .Z(c[1127]) );
  NANDN U864 ( .A(n696), .B(sreg[1127]), .Z(n700) );
  NAND U865 ( .A(n698), .B(n697), .Z(n699) );
  AND U866 ( .A(n700), .B(n699), .Z(n703) );
  NAND U867 ( .A(b[0]), .B(a[105]), .Z(n701) );
  XNOR U868 ( .A(sreg[1128]), .B(n701), .Z(n702) );
  XNOR U869 ( .A(n703), .B(n702), .Z(c[1128]) );
  NAND U870 ( .A(b[0]), .B(a[106]), .Z(n706) );
  XNOR U871 ( .A(sreg[1129]), .B(n706), .Z(n708) );
  NANDN U872 ( .A(sreg[1128]), .B(n701), .Z(n705) );
  NAND U873 ( .A(n703), .B(n702), .Z(n704) );
  NAND U874 ( .A(n705), .B(n704), .Z(n707) );
  XNOR U875 ( .A(n708), .B(n707), .Z(c[1129]) );
  NAND U876 ( .A(b[0]), .B(a[107]), .Z(n711) );
  XNOR U877 ( .A(sreg[1130]), .B(n711), .Z(n713) );
  NANDN U878 ( .A(sreg[1129]), .B(n706), .Z(n710) );
  NAND U879 ( .A(n708), .B(n707), .Z(n709) );
  AND U880 ( .A(n710), .B(n709), .Z(n712) );
  XOR U881 ( .A(n713), .B(n712), .Z(c[1130]) );
  NANDN U882 ( .A(n711), .B(sreg[1130]), .Z(n715) );
  NAND U883 ( .A(n713), .B(n712), .Z(n714) );
  AND U884 ( .A(n715), .B(n714), .Z(n718) );
  NAND U885 ( .A(b[0]), .B(a[108]), .Z(n716) );
  XNOR U886 ( .A(sreg[1131]), .B(n716), .Z(n717) );
  XNOR U887 ( .A(n718), .B(n717), .Z(c[1131]) );
  NAND U888 ( .A(b[0]), .B(a[109]), .Z(n721) );
  XNOR U889 ( .A(sreg[1132]), .B(n721), .Z(n723) );
  NANDN U890 ( .A(sreg[1131]), .B(n716), .Z(n720) );
  NAND U891 ( .A(n718), .B(n717), .Z(n719) );
  NAND U892 ( .A(n720), .B(n719), .Z(n722) );
  XNOR U893 ( .A(n723), .B(n722), .Z(c[1132]) );
  NANDN U894 ( .A(sreg[1132]), .B(n721), .Z(n725) );
  NAND U895 ( .A(n723), .B(n722), .Z(n724) );
  AND U896 ( .A(n725), .B(n724), .Z(n728) );
  NAND U897 ( .A(b[0]), .B(a[110]), .Z(n727) );
  XOR U898 ( .A(sreg[1133]), .B(n727), .Z(n726) );
  XNOR U899 ( .A(n728), .B(n726), .Z(c[1133]) );
  NAND U900 ( .A(b[0]), .B(a[111]), .Z(n729) );
  XNOR U901 ( .A(sreg[1134]), .B(n729), .Z(n730) );
  XOR U902 ( .A(n731), .B(n730), .Z(c[1134]) );
  NANDN U903 ( .A(sreg[1134]), .B(n729), .Z(n733) );
  NANDN U904 ( .A(n731), .B(n730), .Z(n732) );
  AND U905 ( .A(n733), .B(n732), .Z(n736) );
  NAND U906 ( .A(b[0]), .B(a[112]), .Z(n735) );
  XOR U907 ( .A(sreg[1135]), .B(n735), .Z(n734) );
  XNOR U908 ( .A(n736), .B(n734), .Z(c[1135]) );
  NAND U909 ( .A(b[0]), .B(a[113]), .Z(n738) );
  XOR U910 ( .A(sreg[1136]), .B(n738), .Z(n737) );
  XNOR U911 ( .A(n739), .B(n737), .Z(c[1136]) );
  NAND U912 ( .A(b[0]), .B(a[114]), .Z(n740) );
  XNOR U913 ( .A(sreg[1137]), .B(n740), .Z(n741) );
  XOR U914 ( .A(n742), .B(n741), .Z(c[1137]) );
  NAND U915 ( .A(b[0]), .B(a[115]), .Z(n745) );
  XNOR U916 ( .A(sreg[1138]), .B(n745), .Z(n747) );
  NANDN U917 ( .A(n740), .B(sreg[1137]), .Z(n744) );
  NAND U918 ( .A(n742), .B(n741), .Z(n743) );
  AND U919 ( .A(n744), .B(n743), .Z(n746) );
  XNOR U920 ( .A(n747), .B(n746), .Z(c[1138]) );
  NAND U921 ( .A(b[0]), .B(a[116]), .Z(n750) );
  XNOR U922 ( .A(sreg[1139]), .B(n750), .Z(n752) );
  NANDN U923 ( .A(sreg[1138]), .B(n745), .Z(n749) );
  NAND U924 ( .A(n747), .B(n746), .Z(n748) );
  NAND U925 ( .A(n749), .B(n748), .Z(n751) );
  XNOR U926 ( .A(n752), .B(n751), .Z(c[1139]) );
  NAND U927 ( .A(b[0]), .B(a[117]), .Z(n755) );
  XNOR U928 ( .A(sreg[1140]), .B(n755), .Z(n757) );
  NANDN U929 ( .A(sreg[1139]), .B(n750), .Z(n754) );
  NAND U930 ( .A(n752), .B(n751), .Z(n753) );
  AND U931 ( .A(n754), .B(n753), .Z(n756) );
  XOR U932 ( .A(n757), .B(n756), .Z(c[1140]) );
  NAND U933 ( .A(b[0]), .B(a[118]), .Z(n760) );
  XNOR U934 ( .A(sreg[1141]), .B(n760), .Z(n762) );
  NANDN U935 ( .A(n755), .B(sreg[1140]), .Z(n759) );
  NAND U936 ( .A(n757), .B(n756), .Z(n758) );
  NAND U937 ( .A(n759), .B(n758), .Z(n761) );
  XOR U938 ( .A(n762), .B(n761), .Z(c[1141]) );
  NANDN U939 ( .A(n760), .B(sreg[1141]), .Z(n764) );
  NAND U940 ( .A(n762), .B(n761), .Z(n763) );
  AND U941 ( .A(n764), .B(n763), .Z(n767) );
  NAND U942 ( .A(b[0]), .B(a[119]), .Z(n765) );
  XNOR U943 ( .A(sreg[1142]), .B(n765), .Z(n766) );
  XNOR U944 ( .A(n767), .B(n766), .Z(c[1142]) );
  NAND U945 ( .A(b[0]), .B(a[120]), .Z(n770) );
  XNOR U946 ( .A(sreg[1143]), .B(n770), .Z(n772) );
  NANDN U947 ( .A(sreg[1142]), .B(n765), .Z(n769) );
  NAND U948 ( .A(n767), .B(n766), .Z(n768) );
  NAND U949 ( .A(n769), .B(n768), .Z(n771) );
  XNOR U950 ( .A(n772), .B(n771), .Z(c[1143]) );
  NAND U951 ( .A(b[0]), .B(a[121]), .Z(n775) );
  XNOR U952 ( .A(sreg[1144]), .B(n775), .Z(n777) );
  NANDN U953 ( .A(sreg[1143]), .B(n770), .Z(n774) );
  NAND U954 ( .A(n772), .B(n771), .Z(n773) );
  AND U955 ( .A(n774), .B(n773), .Z(n776) );
  XOR U956 ( .A(n777), .B(n776), .Z(c[1144]) );
  NANDN U957 ( .A(n775), .B(sreg[1144]), .Z(n779) );
  NAND U958 ( .A(n777), .B(n776), .Z(n778) );
  AND U959 ( .A(n779), .B(n778), .Z(n782) );
  NAND U960 ( .A(b[0]), .B(a[122]), .Z(n780) );
  XNOR U961 ( .A(sreg[1145]), .B(n780), .Z(n781) );
  XNOR U962 ( .A(n782), .B(n781), .Z(c[1145]) );
  NAND U963 ( .A(b[0]), .B(a[123]), .Z(n785) );
  XNOR U964 ( .A(sreg[1146]), .B(n785), .Z(n787) );
  NANDN U965 ( .A(sreg[1145]), .B(n780), .Z(n784) );
  NAND U966 ( .A(n782), .B(n781), .Z(n783) );
  NAND U967 ( .A(n784), .B(n783), .Z(n786) );
  XNOR U968 ( .A(n787), .B(n786), .Z(c[1146]) );
  NAND U969 ( .A(b[0]), .B(a[124]), .Z(n790) );
  XNOR U970 ( .A(sreg[1147]), .B(n790), .Z(n792) );
  NANDN U971 ( .A(sreg[1146]), .B(n785), .Z(n789) );
  NAND U972 ( .A(n787), .B(n786), .Z(n788) );
  AND U973 ( .A(n789), .B(n788), .Z(n791) );
  XOR U974 ( .A(n792), .B(n791), .Z(c[1147]) );
  NANDN U975 ( .A(n790), .B(sreg[1147]), .Z(n794) );
  NAND U976 ( .A(n792), .B(n791), .Z(n793) );
  AND U977 ( .A(n794), .B(n793), .Z(n797) );
  NAND U978 ( .A(b[0]), .B(a[125]), .Z(n795) );
  XNOR U979 ( .A(sreg[1148]), .B(n795), .Z(n796) );
  XNOR U980 ( .A(n797), .B(n796), .Z(c[1148]) );
  NAND U981 ( .A(b[0]), .B(a[126]), .Z(n800) );
  XNOR U982 ( .A(sreg[1149]), .B(n800), .Z(n802) );
  NANDN U983 ( .A(sreg[1148]), .B(n795), .Z(n799) );
  NAND U984 ( .A(n797), .B(n796), .Z(n798) );
  NAND U985 ( .A(n799), .B(n798), .Z(n801) );
  XNOR U986 ( .A(n802), .B(n801), .Z(c[1149]) );
  NAND U987 ( .A(b[0]), .B(a[127]), .Z(n805) );
  XNOR U988 ( .A(sreg[1150]), .B(n805), .Z(n807) );
  NANDN U989 ( .A(sreg[1149]), .B(n800), .Z(n804) );
  NAND U990 ( .A(n802), .B(n801), .Z(n803) );
  NAND U991 ( .A(n804), .B(n803), .Z(n806) );
  XNOR U992 ( .A(n807), .B(n806), .Z(c[1150]) );
  NAND U993 ( .A(b[0]), .B(a[128]), .Z(n810) );
  XNOR U994 ( .A(sreg[1151]), .B(n810), .Z(n812) );
  NANDN U995 ( .A(sreg[1150]), .B(n805), .Z(n809) );
  NAND U996 ( .A(n807), .B(n806), .Z(n808) );
  NAND U997 ( .A(n809), .B(n808), .Z(n811) );
  XNOR U998 ( .A(n812), .B(n811), .Z(c[1151]) );
  NAND U999 ( .A(b[0]), .B(a[129]), .Z(n815) );
  XNOR U1000 ( .A(sreg[1152]), .B(n815), .Z(n817) );
  NANDN U1001 ( .A(sreg[1151]), .B(n810), .Z(n814) );
  NAND U1002 ( .A(n812), .B(n811), .Z(n813) );
  NAND U1003 ( .A(n814), .B(n813), .Z(n816) );
  XNOR U1004 ( .A(n817), .B(n816), .Z(c[1152]) );
  NAND U1005 ( .A(b[0]), .B(a[130]), .Z(n820) );
  XNOR U1006 ( .A(sreg[1153]), .B(n820), .Z(n822) );
  NANDN U1007 ( .A(sreg[1152]), .B(n815), .Z(n819) );
  NAND U1008 ( .A(n817), .B(n816), .Z(n818) );
  NAND U1009 ( .A(n819), .B(n818), .Z(n821) );
  XNOR U1010 ( .A(n822), .B(n821), .Z(c[1153]) );
  NAND U1011 ( .A(b[0]), .B(a[131]), .Z(n825) );
  XNOR U1012 ( .A(sreg[1154]), .B(n825), .Z(n827) );
  NANDN U1013 ( .A(sreg[1153]), .B(n820), .Z(n824) );
  NAND U1014 ( .A(n822), .B(n821), .Z(n823) );
  NAND U1015 ( .A(n824), .B(n823), .Z(n826) );
  XNOR U1016 ( .A(n827), .B(n826), .Z(c[1154]) );
  NAND U1017 ( .A(b[0]), .B(a[132]), .Z(n830) );
  XNOR U1018 ( .A(sreg[1155]), .B(n830), .Z(n832) );
  NANDN U1019 ( .A(sreg[1154]), .B(n825), .Z(n829) );
  NAND U1020 ( .A(n827), .B(n826), .Z(n828) );
  NAND U1021 ( .A(n829), .B(n828), .Z(n831) );
  XNOR U1022 ( .A(n832), .B(n831), .Z(c[1155]) );
  NAND U1023 ( .A(b[0]), .B(a[133]), .Z(n835) );
  XNOR U1024 ( .A(sreg[1156]), .B(n835), .Z(n837) );
  NANDN U1025 ( .A(sreg[1155]), .B(n830), .Z(n834) );
  NAND U1026 ( .A(n832), .B(n831), .Z(n833) );
  NAND U1027 ( .A(n834), .B(n833), .Z(n836) );
  XNOR U1028 ( .A(n837), .B(n836), .Z(c[1156]) );
  NAND U1029 ( .A(b[0]), .B(a[134]), .Z(n840) );
  XNOR U1030 ( .A(sreg[1157]), .B(n840), .Z(n842) );
  NANDN U1031 ( .A(sreg[1156]), .B(n835), .Z(n839) );
  NAND U1032 ( .A(n837), .B(n836), .Z(n838) );
  NAND U1033 ( .A(n839), .B(n838), .Z(n841) );
  XNOR U1034 ( .A(n842), .B(n841), .Z(c[1157]) );
  NAND U1035 ( .A(b[0]), .B(a[135]), .Z(n845) );
  XNOR U1036 ( .A(sreg[1158]), .B(n845), .Z(n847) );
  NANDN U1037 ( .A(sreg[1157]), .B(n840), .Z(n844) );
  NAND U1038 ( .A(n842), .B(n841), .Z(n843) );
  NAND U1039 ( .A(n844), .B(n843), .Z(n846) );
  XNOR U1040 ( .A(n847), .B(n846), .Z(c[1158]) );
  NAND U1041 ( .A(b[0]), .B(a[136]), .Z(n850) );
  XNOR U1042 ( .A(sreg[1159]), .B(n850), .Z(n852) );
  NANDN U1043 ( .A(sreg[1158]), .B(n845), .Z(n849) );
  NAND U1044 ( .A(n847), .B(n846), .Z(n848) );
  NAND U1045 ( .A(n849), .B(n848), .Z(n851) );
  XNOR U1046 ( .A(n852), .B(n851), .Z(c[1159]) );
  NAND U1047 ( .A(b[0]), .B(a[137]), .Z(n855) );
  XNOR U1048 ( .A(sreg[1160]), .B(n855), .Z(n857) );
  NANDN U1049 ( .A(sreg[1159]), .B(n850), .Z(n854) );
  NAND U1050 ( .A(n852), .B(n851), .Z(n853) );
  NAND U1051 ( .A(n854), .B(n853), .Z(n856) );
  XNOR U1052 ( .A(n857), .B(n856), .Z(c[1160]) );
  NAND U1053 ( .A(b[0]), .B(a[138]), .Z(n860) );
  XNOR U1054 ( .A(sreg[1161]), .B(n860), .Z(n862) );
  NANDN U1055 ( .A(sreg[1160]), .B(n855), .Z(n859) );
  NAND U1056 ( .A(n857), .B(n856), .Z(n858) );
  AND U1057 ( .A(n859), .B(n858), .Z(n861) );
  XOR U1058 ( .A(n862), .B(n861), .Z(c[1161]) );
  NANDN U1059 ( .A(n860), .B(sreg[1161]), .Z(n864) );
  NAND U1060 ( .A(n862), .B(n861), .Z(n863) );
  AND U1061 ( .A(n864), .B(n863), .Z(n867) );
  NAND U1062 ( .A(b[0]), .B(a[139]), .Z(n865) );
  XNOR U1063 ( .A(sreg[1162]), .B(n865), .Z(n866) );
  XNOR U1064 ( .A(n867), .B(n866), .Z(c[1162]) );
  NAND U1065 ( .A(b[0]), .B(a[140]), .Z(n870) );
  XNOR U1066 ( .A(sreg[1163]), .B(n870), .Z(n872) );
  NANDN U1067 ( .A(sreg[1162]), .B(n865), .Z(n869) );
  NAND U1068 ( .A(n867), .B(n866), .Z(n868) );
  NAND U1069 ( .A(n869), .B(n868), .Z(n871) );
  XNOR U1070 ( .A(n872), .B(n871), .Z(c[1163]) );
  NAND U1071 ( .A(b[0]), .B(a[141]), .Z(n875) );
  XNOR U1072 ( .A(sreg[1164]), .B(n875), .Z(n877) );
  NANDN U1073 ( .A(sreg[1163]), .B(n870), .Z(n874) );
  NAND U1074 ( .A(n872), .B(n871), .Z(n873) );
  NAND U1075 ( .A(n874), .B(n873), .Z(n876) );
  XNOR U1076 ( .A(n877), .B(n876), .Z(c[1164]) );
  NANDN U1077 ( .A(sreg[1164]), .B(n875), .Z(n879) );
  NAND U1078 ( .A(n877), .B(n876), .Z(n878) );
  AND U1079 ( .A(n879), .B(n878), .Z(n882) );
  NAND U1080 ( .A(b[0]), .B(a[142]), .Z(n880) );
  XNOR U1081 ( .A(sreg[1165]), .B(n880), .Z(n881) );
  XOR U1082 ( .A(n882), .B(n881), .Z(c[1165]) );
  NAND U1083 ( .A(b[0]), .B(a[143]), .Z(n885) );
  XNOR U1084 ( .A(sreg[1166]), .B(n885), .Z(n887) );
  NANDN U1085 ( .A(n880), .B(sreg[1165]), .Z(n884) );
  NAND U1086 ( .A(n882), .B(n881), .Z(n883) );
  AND U1087 ( .A(n884), .B(n883), .Z(n886) );
  XNOR U1088 ( .A(n887), .B(n886), .Z(c[1166]) );
  NAND U1089 ( .A(b[0]), .B(a[144]), .Z(n892) );
  NANDN U1090 ( .A(sreg[1166]), .B(n885), .Z(n889) );
  NAND U1091 ( .A(n887), .B(n886), .Z(n888) );
  AND U1092 ( .A(n889), .B(n888), .Z(n891) );
  XOR U1093 ( .A(sreg[1167]), .B(n891), .Z(n890) );
  XNOR U1094 ( .A(n892), .B(n890), .Z(c[1167]) );
  NAND U1095 ( .A(b[0]), .B(a[145]), .Z(n893) );
  XNOR U1096 ( .A(sreg[1168]), .B(n893), .Z(n894) );
  XOR U1097 ( .A(n895), .B(n894), .Z(c[1168]) );
  NAND U1098 ( .A(b[0]), .B(a[146]), .Z(n898) );
  XNOR U1099 ( .A(sreg[1169]), .B(n898), .Z(n900) );
  NANDN U1100 ( .A(n893), .B(sreg[1168]), .Z(n897) );
  NAND U1101 ( .A(n895), .B(n894), .Z(n896) );
  NAND U1102 ( .A(n897), .B(n896), .Z(n899) );
  XOR U1103 ( .A(n900), .B(n899), .Z(c[1169]) );
  AND U1104 ( .A(b[0]), .B(a[147]), .Z(n904) );
  NANDN U1105 ( .A(n898), .B(sreg[1169]), .Z(n902) );
  NAND U1106 ( .A(n900), .B(n899), .Z(n901) );
  AND U1107 ( .A(n902), .B(n901), .Z(n905) );
  XNOR U1108 ( .A(sreg[1170]), .B(n905), .Z(n903) );
  XOR U1109 ( .A(n904), .B(n903), .Z(c[1170]) );
  NAND U1110 ( .A(b[0]), .B(a[148]), .Z(n906) );
  XNOR U1111 ( .A(sreg[1171]), .B(n906), .Z(n907) );
  XNOR U1112 ( .A(n908), .B(n907), .Z(c[1171]) );
  NAND U1113 ( .A(b[0]), .B(a[149]), .Z(n911) );
  XNOR U1114 ( .A(sreg[1172]), .B(n911), .Z(n913) );
  NANDN U1115 ( .A(n906), .B(sreg[1171]), .Z(n910) );
  NANDN U1116 ( .A(n908), .B(n907), .Z(n909) );
  NAND U1117 ( .A(n910), .B(n909), .Z(n912) );
  XOR U1118 ( .A(n913), .B(n912), .Z(c[1172]) );
  NANDN U1119 ( .A(n911), .B(sreg[1172]), .Z(n915) );
  NAND U1120 ( .A(n913), .B(n912), .Z(n914) );
  NAND U1121 ( .A(n915), .B(n914), .Z(n918) );
  NAND U1122 ( .A(b[0]), .B(a[150]), .Z(n917) );
  XOR U1123 ( .A(sreg[1173]), .B(n917), .Z(n916) );
  XNOR U1124 ( .A(n918), .B(n916), .Z(c[1173]) );
  NAND U1125 ( .A(b[0]), .B(a[151]), .Z(n919) );
  XNOR U1126 ( .A(sreg[1174]), .B(n919), .Z(n920) );
  XOR U1127 ( .A(n921), .B(n920), .Z(c[1174]) );
  NAND U1128 ( .A(b[0]), .B(a[152]), .Z(n924) );
  XNOR U1129 ( .A(sreg[1175]), .B(n924), .Z(n926) );
  NANDN U1130 ( .A(n919), .B(sreg[1174]), .Z(n923) );
  NAND U1131 ( .A(n921), .B(n920), .Z(n922) );
  NAND U1132 ( .A(n923), .B(n922), .Z(n925) );
  XOR U1133 ( .A(n926), .B(n925), .Z(c[1175]) );
  AND U1134 ( .A(b[0]), .B(a[153]), .Z(n930) );
  NANDN U1135 ( .A(n924), .B(sreg[1175]), .Z(n928) );
  NAND U1136 ( .A(n926), .B(n925), .Z(n927) );
  AND U1137 ( .A(n928), .B(n927), .Z(n931) );
  XNOR U1138 ( .A(sreg[1176]), .B(n931), .Z(n929) );
  XOR U1139 ( .A(n930), .B(n929), .Z(c[1176]) );
  NAND U1140 ( .A(b[0]), .B(a[154]), .Z(n932) );
  XNOR U1141 ( .A(sreg[1177]), .B(n932), .Z(n933) );
  XNOR U1142 ( .A(n934), .B(n933), .Z(c[1177]) );
  NAND U1143 ( .A(b[0]), .B(a[155]), .Z(n937) );
  XNOR U1144 ( .A(sreg[1178]), .B(n937), .Z(n939) );
  NANDN U1145 ( .A(n932), .B(sreg[1177]), .Z(n936) );
  NANDN U1146 ( .A(n934), .B(n933), .Z(n935) );
  NAND U1147 ( .A(n936), .B(n935), .Z(n938) );
  XOR U1148 ( .A(n939), .B(n938), .Z(c[1178]) );
  NANDN U1149 ( .A(n937), .B(sreg[1178]), .Z(n941) );
  NAND U1150 ( .A(n939), .B(n938), .Z(n940) );
  AND U1151 ( .A(n941), .B(n940), .Z(n944) );
  NAND U1152 ( .A(b[0]), .B(a[156]), .Z(n942) );
  XNOR U1153 ( .A(sreg[1179]), .B(n942), .Z(n943) );
  XNOR U1154 ( .A(n944), .B(n943), .Z(c[1179]) );
  NAND U1155 ( .A(b[0]), .B(a[157]), .Z(n947) );
  XNOR U1156 ( .A(sreg[1180]), .B(n947), .Z(n949) );
  NANDN U1157 ( .A(sreg[1179]), .B(n942), .Z(n946) );
  NAND U1158 ( .A(n944), .B(n943), .Z(n945) );
  AND U1159 ( .A(n946), .B(n945), .Z(n948) );
  XOR U1160 ( .A(n949), .B(n948), .Z(c[1180]) );
  NAND U1161 ( .A(b[0]), .B(a[158]), .Z(n952) );
  XNOR U1162 ( .A(sreg[1181]), .B(n952), .Z(n954) );
  NANDN U1163 ( .A(n947), .B(sreg[1180]), .Z(n951) );
  NAND U1164 ( .A(n949), .B(n948), .Z(n950) );
  NAND U1165 ( .A(n951), .B(n950), .Z(n953) );
  XOR U1166 ( .A(n954), .B(n953), .Z(c[1181]) );
  NAND U1167 ( .A(b[0]), .B(a[159]), .Z(n957) );
  XNOR U1168 ( .A(sreg[1182]), .B(n957), .Z(n959) );
  NANDN U1169 ( .A(n952), .B(sreg[1181]), .Z(n956) );
  NAND U1170 ( .A(n954), .B(n953), .Z(n955) );
  AND U1171 ( .A(n956), .B(n955), .Z(n958) );
  XNOR U1172 ( .A(n959), .B(n958), .Z(c[1182]) );
  NAND U1173 ( .A(b[0]), .B(a[160]), .Z(n962) );
  XNOR U1174 ( .A(sreg[1183]), .B(n962), .Z(n964) );
  NANDN U1175 ( .A(sreg[1182]), .B(n957), .Z(n961) );
  NAND U1176 ( .A(n959), .B(n958), .Z(n960) );
  AND U1177 ( .A(n961), .B(n960), .Z(n963) );
  XOR U1178 ( .A(n964), .B(n963), .Z(c[1183]) );
  NAND U1179 ( .A(b[0]), .B(a[161]), .Z(n967) );
  XNOR U1180 ( .A(sreg[1184]), .B(n967), .Z(n969) );
  NANDN U1181 ( .A(n962), .B(sreg[1183]), .Z(n966) );
  NAND U1182 ( .A(n964), .B(n963), .Z(n965) );
  NAND U1183 ( .A(n966), .B(n965), .Z(n968) );
  XOR U1184 ( .A(n969), .B(n968), .Z(c[1184]) );
  NAND U1185 ( .A(b[0]), .B(a[162]), .Z(n972) );
  XNOR U1186 ( .A(sreg[1185]), .B(n972), .Z(n974) );
  NANDN U1187 ( .A(n967), .B(sreg[1184]), .Z(n971) );
  NAND U1188 ( .A(n969), .B(n968), .Z(n970) );
  NAND U1189 ( .A(n971), .B(n970), .Z(n973) );
  XOR U1190 ( .A(n974), .B(n973), .Z(c[1185]) );
  NAND U1191 ( .A(b[0]), .B(a[163]), .Z(n977) );
  XNOR U1192 ( .A(sreg[1186]), .B(n977), .Z(n979) );
  NANDN U1193 ( .A(n972), .B(sreg[1185]), .Z(n976) );
  NAND U1194 ( .A(n974), .B(n973), .Z(n975) );
  AND U1195 ( .A(n976), .B(n975), .Z(n978) );
  XNOR U1196 ( .A(n979), .B(n978), .Z(c[1186]) );
  NANDN U1197 ( .A(sreg[1186]), .B(n977), .Z(n981) );
  NAND U1198 ( .A(n979), .B(n978), .Z(n980) );
  AND U1199 ( .A(n981), .B(n980), .Z(n984) );
  NAND U1200 ( .A(b[0]), .B(a[164]), .Z(n982) );
  XNOR U1201 ( .A(sreg[1187]), .B(n982), .Z(n983) );
  XOR U1202 ( .A(n984), .B(n983), .Z(c[1187]) );
  NAND U1203 ( .A(b[0]), .B(a[165]), .Z(n987) );
  XNOR U1204 ( .A(sreg[1188]), .B(n987), .Z(n989) );
  NANDN U1205 ( .A(n982), .B(sreg[1187]), .Z(n986) );
  NAND U1206 ( .A(n984), .B(n983), .Z(n985) );
  NAND U1207 ( .A(n986), .B(n985), .Z(n988) );
  XOR U1208 ( .A(n989), .B(n988), .Z(c[1188]) );
  NAND U1209 ( .A(b[0]), .B(a[166]), .Z(n992) );
  XNOR U1210 ( .A(sreg[1189]), .B(n992), .Z(n994) );
  NANDN U1211 ( .A(n987), .B(sreg[1188]), .Z(n991) );
  NAND U1212 ( .A(n989), .B(n988), .Z(n990) );
  AND U1213 ( .A(n991), .B(n990), .Z(n993) );
  XNOR U1214 ( .A(n994), .B(n993), .Z(c[1189]) );
  NANDN U1215 ( .A(sreg[1189]), .B(n992), .Z(n996) );
  NAND U1216 ( .A(n994), .B(n993), .Z(n995) );
  AND U1217 ( .A(n996), .B(n995), .Z(n999) );
  NAND U1218 ( .A(b[0]), .B(a[167]), .Z(n997) );
  XNOR U1219 ( .A(sreg[1190]), .B(n997), .Z(n998) );
  XOR U1220 ( .A(n999), .B(n998), .Z(c[1190]) );
  NAND U1221 ( .A(b[0]), .B(a[168]), .Z(n1002) );
  XNOR U1222 ( .A(sreg[1191]), .B(n1002), .Z(n1004) );
  NANDN U1223 ( .A(n997), .B(sreg[1190]), .Z(n1001) );
  NAND U1224 ( .A(n999), .B(n998), .Z(n1000) );
  NAND U1225 ( .A(n1001), .B(n1000), .Z(n1003) );
  XOR U1226 ( .A(n1004), .B(n1003), .Z(c[1191]) );
  NANDN U1227 ( .A(n1002), .B(sreg[1191]), .Z(n1006) );
  NAND U1228 ( .A(n1004), .B(n1003), .Z(n1005) );
  AND U1229 ( .A(n1006), .B(n1005), .Z(n1009) );
  NAND U1230 ( .A(b[0]), .B(a[169]), .Z(n1007) );
  XNOR U1231 ( .A(sreg[1192]), .B(n1007), .Z(n1008) );
  XNOR U1232 ( .A(n1009), .B(n1008), .Z(c[1192]) );
  NAND U1233 ( .A(b[0]), .B(a[170]), .Z(n1012) );
  XNOR U1234 ( .A(sreg[1193]), .B(n1012), .Z(n1014) );
  NANDN U1235 ( .A(sreg[1192]), .B(n1007), .Z(n1011) );
  NAND U1236 ( .A(n1009), .B(n1008), .Z(n1010) );
  NAND U1237 ( .A(n1011), .B(n1010), .Z(n1013) );
  XNOR U1238 ( .A(n1014), .B(n1013), .Z(c[1193]) );
  NANDN U1239 ( .A(sreg[1193]), .B(n1012), .Z(n1016) );
  NAND U1240 ( .A(n1014), .B(n1013), .Z(n1015) );
  AND U1241 ( .A(n1016), .B(n1015), .Z(n1019) );
  NAND U1242 ( .A(b[0]), .B(a[171]), .Z(n1017) );
  XNOR U1243 ( .A(sreg[1194]), .B(n1017), .Z(n1018) );
  XOR U1244 ( .A(n1019), .B(n1018), .Z(c[1194]) );
  NANDN U1245 ( .A(n1017), .B(sreg[1194]), .Z(n1021) );
  NAND U1246 ( .A(n1019), .B(n1018), .Z(n1020) );
  AND U1247 ( .A(n1021), .B(n1020), .Z(n1024) );
  NAND U1248 ( .A(b[0]), .B(a[172]), .Z(n1022) );
  XNOR U1249 ( .A(sreg[1195]), .B(n1022), .Z(n1023) );
  XNOR U1250 ( .A(n1024), .B(n1023), .Z(c[1195]) );
  NAND U1251 ( .A(b[0]), .B(a[173]), .Z(n1027) );
  XNOR U1252 ( .A(sreg[1196]), .B(n1027), .Z(n1029) );
  NANDN U1253 ( .A(sreg[1195]), .B(n1022), .Z(n1026) );
  NAND U1254 ( .A(n1024), .B(n1023), .Z(n1025) );
  NAND U1255 ( .A(n1026), .B(n1025), .Z(n1028) );
  XNOR U1256 ( .A(n1029), .B(n1028), .Z(c[1196]) );
  NANDN U1257 ( .A(sreg[1196]), .B(n1027), .Z(n1031) );
  NAND U1258 ( .A(n1029), .B(n1028), .Z(n1030) );
  AND U1259 ( .A(n1031), .B(n1030), .Z(n1034) );
  NAND U1260 ( .A(b[0]), .B(a[174]), .Z(n1032) );
  XNOR U1261 ( .A(sreg[1197]), .B(n1032), .Z(n1033) );
  XOR U1262 ( .A(n1034), .B(n1033), .Z(c[1197]) );
  NANDN U1263 ( .A(n1032), .B(sreg[1197]), .Z(n1036) );
  NAND U1264 ( .A(n1034), .B(n1033), .Z(n1035) );
  AND U1265 ( .A(n1036), .B(n1035), .Z(n1039) );
  NAND U1266 ( .A(b[0]), .B(a[175]), .Z(n1037) );
  XNOR U1267 ( .A(sreg[1198]), .B(n1037), .Z(n1038) );
  XNOR U1268 ( .A(n1039), .B(n1038), .Z(c[1198]) );
  NAND U1269 ( .A(b[0]), .B(a[176]), .Z(n1042) );
  XNOR U1270 ( .A(sreg[1199]), .B(n1042), .Z(n1044) );
  NANDN U1271 ( .A(sreg[1198]), .B(n1037), .Z(n1041) );
  NAND U1272 ( .A(n1039), .B(n1038), .Z(n1040) );
  AND U1273 ( .A(n1041), .B(n1040), .Z(n1043) );
  XOR U1274 ( .A(n1044), .B(n1043), .Z(c[1199]) );
  NAND U1275 ( .A(b[0]), .B(a[177]), .Z(n1047) );
  XNOR U1276 ( .A(sreg[1200]), .B(n1047), .Z(n1049) );
  NANDN U1277 ( .A(n1042), .B(sreg[1199]), .Z(n1046) );
  NAND U1278 ( .A(n1044), .B(n1043), .Z(n1045) );
  NAND U1279 ( .A(n1046), .B(n1045), .Z(n1048) );
  XOR U1280 ( .A(n1049), .B(n1048), .Z(c[1200]) );
  NAND U1281 ( .A(b[0]), .B(a[178]), .Z(n1052) );
  XNOR U1282 ( .A(sreg[1201]), .B(n1052), .Z(n1054) );
  NANDN U1283 ( .A(n1047), .B(sreg[1200]), .Z(n1051) );
  NAND U1284 ( .A(n1049), .B(n1048), .Z(n1050) );
  AND U1285 ( .A(n1051), .B(n1050), .Z(n1053) );
  XNOR U1286 ( .A(n1054), .B(n1053), .Z(c[1201]) );
  NAND U1287 ( .A(b[0]), .B(a[179]), .Z(n1057) );
  XNOR U1288 ( .A(sreg[1202]), .B(n1057), .Z(n1059) );
  NANDN U1289 ( .A(sreg[1201]), .B(n1052), .Z(n1056) );
  NAND U1290 ( .A(n1054), .B(n1053), .Z(n1055) );
  NAND U1291 ( .A(n1056), .B(n1055), .Z(n1058) );
  XNOR U1292 ( .A(n1059), .B(n1058), .Z(c[1202]) );
  NAND U1293 ( .A(b[0]), .B(a[180]), .Z(n1062) );
  XNOR U1294 ( .A(sreg[1203]), .B(n1062), .Z(n1064) );
  NANDN U1295 ( .A(sreg[1202]), .B(n1057), .Z(n1061) );
  NAND U1296 ( .A(n1059), .B(n1058), .Z(n1060) );
  AND U1297 ( .A(n1061), .B(n1060), .Z(n1063) );
  XOR U1298 ( .A(n1064), .B(n1063), .Z(c[1203]) );
  NANDN U1299 ( .A(n1062), .B(sreg[1203]), .Z(n1066) );
  NAND U1300 ( .A(n1064), .B(n1063), .Z(n1065) );
  AND U1301 ( .A(n1066), .B(n1065), .Z(n1069) );
  NAND U1302 ( .A(b[0]), .B(a[181]), .Z(n1067) );
  XNOR U1303 ( .A(sreg[1204]), .B(n1067), .Z(n1068) );
  XNOR U1304 ( .A(n1069), .B(n1068), .Z(c[1204]) );
  NAND U1305 ( .A(b[0]), .B(a[182]), .Z(n1072) );
  XNOR U1306 ( .A(sreg[1205]), .B(n1072), .Z(n1074) );
  NANDN U1307 ( .A(sreg[1204]), .B(n1067), .Z(n1071) );
  NAND U1308 ( .A(n1069), .B(n1068), .Z(n1070) );
  NAND U1309 ( .A(n1071), .B(n1070), .Z(n1073) );
  XNOR U1310 ( .A(n1074), .B(n1073), .Z(c[1205]) );
  NAND U1311 ( .A(b[0]), .B(a[183]), .Z(n1077) );
  XNOR U1312 ( .A(sreg[1206]), .B(n1077), .Z(n1079) );
  NANDN U1313 ( .A(sreg[1205]), .B(n1072), .Z(n1076) );
  NAND U1314 ( .A(n1074), .B(n1073), .Z(n1075) );
  NAND U1315 ( .A(n1076), .B(n1075), .Z(n1078) );
  XNOR U1316 ( .A(n1079), .B(n1078), .Z(c[1206]) );
  NANDN U1317 ( .A(sreg[1206]), .B(n1077), .Z(n1081) );
  NAND U1318 ( .A(n1079), .B(n1078), .Z(n1080) );
  AND U1319 ( .A(n1081), .B(n1080), .Z(n1084) );
  NAND U1320 ( .A(b[0]), .B(a[184]), .Z(n1082) );
  XNOR U1321 ( .A(sreg[1207]), .B(n1082), .Z(n1083) );
  XOR U1322 ( .A(n1084), .B(n1083), .Z(c[1207]) );
  NAND U1323 ( .A(b[0]), .B(a[185]), .Z(n1087) );
  XNOR U1324 ( .A(sreg[1208]), .B(n1087), .Z(n1089) );
  NANDN U1325 ( .A(n1082), .B(sreg[1207]), .Z(n1086) );
  NAND U1326 ( .A(n1084), .B(n1083), .Z(n1085) );
  NAND U1327 ( .A(n1086), .B(n1085), .Z(n1088) );
  XOR U1328 ( .A(n1089), .B(n1088), .Z(c[1208]) );
  NAND U1329 ( .A(b[0]), .B(a[186]), .Z(n1092) );
  XNOR U1330 ( .A(sreg[1209]), .B(n1092), .Z(n1094) );
  NANDN U1331 ( .A(n1087), .B(sreg[1208]), .Z(n1091) );
  NAND U1332 ( .A(n1089), .B(n1088), .Z(n1090) );
  NAND U1333 ( .A(n1091), .B(n1090), .Z(n1093) );
  XOR U1334 ( .A(n1094), .B(n1093), .Z(c[1209]) );
  NAND U1335 ( .A(b[0]), .B(a[187]), .Z(n1097) );
  XNOR U1336 ( .A(sreg[1210]), .B(n1097), .Z(n1099) );
  NANDN U1337 ( .A(n1092), .B(sreg[1209]), .Z(n1096) );
  NAND U1338 ( .A(n1094), .B(n1093), .Z(n1095) );
  NAND U1339 ( .A(n1096), .B(n1095), .Z(n1098) );
  XOR U1340 ( .A(n1099), .B(n1098), .Z(c[1210]) );
  NANDN U1341 ( .A(n1097), .B(sreg[1210]), .Z(n1101) );
  NAND U1342 ( .A(n1099), .B(n1098), .Z(n1100) );
  AND U1343 ( .A(n1101), .B(n1100), .Z(n1104) );
  NAND U1344 ( .A(b[0]), .B(a[188]), .Z(n1102) );
  XNOR U1345 ( .A(sreg[1211]), .B(n1102), .Z(n1103) );
  XNOR U1346 ( .A(n1104), .B(n1103), .Z(c[1211]) );
  NAND U1347 ( .A(b[0]), .B(a[189]), .Z(n1107) );
  XNOR U1348 ( .A(sreg[1212]), .B(n1107), .Z(n1109) );
  NANDN U1349 ( .A(sreg[1211]), .B(n1102), .Z(n1106) );
  NAND U1350 ( .A(n1104), .B(n1103), .Z(n1105) );
  AND U1351 ( .A(n1106), .B(n1105), .Z(n1108) );
  XOR U1352 ( .A(n1109), .B(n1108), .Z(c[1212]) );
  NAND U1353 ( .A(b[0]), .B(a[190]), .Z(n1112) );
  XNOR U1354 ( .A(sreg[1213]), .B(n1112), .Z(n1114) );
  NANDN U1355 ( .A(n1107), .B(sreg[1212]), .Z(n1111) );
  NAND U1356 ( .A(n1109), .B(n1108), .Z(n1110) );
  NAND U1357 ( .A(n1111), .B(n1110), .Z(n1113) );
  XOR U1358 ( .A(n1114), .B(n1113), .Z(c[1213]) );
  NANDN U1359 ( .A(n1112), .B(sreg[1213]), .Z(n1116) );
  NAND U1360 ( .A(n1114), .B(n1113), .Z(n1115) );
  AND U1361 ( .A(n1116), .B(n1115), .Z(n1119) );
  NAND U1362 ( .A(b[0]), .B(a[191]), .Z(n1117) );
  XNOR U1363 ( .A(sreg[1214]), .B(n1117), .Z(n1118) );
  XNOR U1364 ( .A(n1119), .B(n1118), .Z(c[1214]) );
  NAND U1365 ( .A(b[0]), .B(a[192]), .Z(n1122) );
  XNOR U1366 ( .A(sreg[1215]), .B(n1122), .Z(n1124) );
  NANDN U1367 ( .A(sreg[1214]), .B(n1117), .Z(n1121) );
  NAND U1368 ( .A(n1119), .B(n1118), .Z(n1120) );
  AND U1369 ( .A(n1121), .B(n1120), .Z(n1123) );
  XOR U1370 ( .A(n1124), .B(n1123), .Z(c[1215]) );
  NAND U1371 ( .A(b[0]), .B(a[193]), .Z(n1127) );
  XNOR U1372 ( .A(sreg[1216]), .B(n1127), .Z(n1129) );
  NANDN U1373 ( .A(n1122), .B(sreg[1215]), .Z(n1126) );
  NAND U1374 ( .A(n1124), .B(n1123), .Z(n1125) );
  NAND U1375 ( .A(n1126), .B(n1125), .Z(n1128) );
  XOR U1376 ( .A(n1129), .B(n1128), .Z(c[1216]) );
  NAND U1377 ( .A(b[0]), .B(a[194]), .Z(n1132) );
  XNOR U1378 ( .A(sreg[1217]), .B(n1132), .Z(n1134) );
  NANDN U1379 ( .A(n1127), .B(sreg[1216]), .Z(n1131) );
  NAND U1380 ( .A(n1129), .B(n1128), .Z(n1130) );
  NAND U1381 ( .A(n1131), .B(n1130), .Z(n1133) );
  XOR U1382 ( .A(n1134), .B(n1133), .Z(c[1217]) );
  NAND U1383 ( .A(b[0]), .B(a[195]), .Z(n1137) );
  XNOR U1384 ( .A(sreg[1218]), .B(n1137), .Z(n1139) );
  NANDN U1385 ( .A(n1132), .B(sreg[1217]), .Z(n1136) );
  NAND U1386 ( .A(n1134), .B(n1133), .Z(n1135) );
  AND U1387 ( .A(n1136), .B(n1135), .Z(n1138) );
  XNOR U1388 ( .A(n1139), .B(n1138), .Z(c[1218]) );
  NANDN U1389 ( .A(sreg[1218]), .B(n1137), .Z(n1141) );
  NAND U1390 ( .A(n1139), .B(n1138), .Z(n1140) );
  AND U1391 ( .A(n1141), .B(n1140), .Z(n1144) );
  NAND U1392 ( .A(b[0]), .B(a[196]), .Z(n1142) );
  XNOR U1393 ( .A(sreg[1219]), .B(n1142), .Z(n1143) );
  XOR U1394 ( .A(n1144), .B(n1143), .Z(c[1219]) );
  NAND U1395 ( .A(b[0]), .B(a[197]), .Z(n1147) );
  XNOR U1396 ( .A(sreg[1220]), .B(n1147), .Z(n1149) );
  NANDN U1397 ( .A(n1142), .B(sreg[1219]), .Z(n1146) );
  NAND U1398 ( .A(n1144), .B(n1143), .Z(n1145) );
  NAND U1399 ( .A(n1146), .B(n1145), .Z(n1148) );
  XOR U1400 ( .A(n1149), .B(n1148), .Z(c[1220]) );
  NAND U1401 ( .A(b[0]), .B(a[198]), .Z(n1152) );
  XNOR U1402 ( .A(sreg[1221]), .B(n1152), .Z(n1154) );
  NANDN U1403 ( .A(n1147), .B(sreg[1220]), .Z(n1151) );
  NAND U1404 ( .A(n1149), .B(n1148), .Z(n1150) );
  AND U1405 ( .A(n1151), .B(n1150), .Z(n1153) );
  XNOR U1406 ( .A(n1154), .B(n1153), .Z(c[1221]) );
  NANDN U1407 ( .A(sreg[1221]), .B(n1152), .Z(n1156) );
  NAND U1408 ( .A(n1154), .B(n1153), .Z(n1155) );
  AND U1409 ( .A(n1156), .B(n1155), .Z(n1159) );
  NAND U1410 ( .A(b[0]), .B(a[199]), .Z(n1157) );
  XNOR U1411 ( .A(sreg[1222]), .B(n1157), .Z(n1158) );
  XOR U1412 ( .A(n1159), .B(n1158), .Z(c[1222]) );
  NAND U1413 ( .A(b[0]), .B(a[200]), .Z(n1162) );
  XNOR U1414 ( .A(sreg[1223]), .B(n1162), .Z(n1164) );
  NANDN U1415 ( .A(n1157), .B(sreg[1222]), .Z(n1161) );
  NAND U1416 ( .A(n1159), .B(n1158), .Z(n1160) );
  NAND U1417 ( .A(n1161), .B(n1160), .Z(n1163) );
  XOR U1418 ( .A(n1164), .B(n1163), .Z(c[1223]) );
  NANDN U1419 ( .A(n1162), .B(sreg[1223]), .Z(n1166) );
  NAND U1420 ( .A(n1164), .B(n1163), .Z(n1165) );
  AND U1421 ( .A(n1166), .B(n1165), .Z(n1169) );
  NAND U1422 ( .A(b[0]), .B(a[201]), .Z(n1167) );
  XNOR U1423 ( .A(sreg[1224]), .B(n1167), .Z(n1168) );
  XNOR U1424 ( .A(n1169), .B(n1168), .Z(c[1224]) );
  NAND U1425 ( .A(b[0]), .B(a[202]), .Z(n1172) );
  XNOR U1426 ( .A(sreg[1225]), .B(n1172), .Z(n1174) );
  NANDN U1427 ( .A(sreg[1224]), .B(n1167), .Z(n1171) );
  NAND U1428 ( .A(n1169), .B(n1168), .Z(n1170) );
  NAND U1429 ( .A(n1171), .B(n1170), .Z(n1173) );
  XNOR U1430 ( .A(n1174), .B(n1173), .Z(c[1225]) );
  NAND U1431 ( .A(b[0]), .B(a[203]), .Z(n1177) );
  XNOR U1432 ( .A(sreg[1226]), .B(n1177), .Z(n1179) );
  NANDN U1433 ( .A(sreg[1225]), .B(n1172), .Z(n1176) );
  NAND U1434 ( .A(n1174), .B(n1173), .Z(n1175) );
  NAND U1435 ( .A(n1176), .B(n1175), .Z(n1178) );
  XNOR U1436 ( .A(n1179), .B(n1178), .Z(c[1226]) );
  NAND U1437 ( .A(b[0]), .B(a[204]), .Z(n1182) );
  XNOR U1438 ( .A(sreg[1227]), .B(n1182), .Z(n1184) );
  NANDN U1439 ( .A(sreg[1226]), .B(n1177), .Z(n1181) );
  NAND U1440 ( .A(n1179), .B(n1178), .Z(n1180) );
  NAND U1441 ( .A(n1181), .B(n1180), .Z(n1183) );
  XNOR U1442 ( .A(n1184), .B(n1183), .Z(c[1227]) );
  NAND U1443 ( .A(b[0]), .B(a[205]), .Z(n1187) );
  XNOR U1444 ( .A(sreg[1228]), .B(n1187), .Z(n1189) );
  NANDN U1445 ( .A(sreg[1227]), .B(n1182), .Z(n1186) );
  NAND U1446 ( .A(n1184), .B(n1183), .Z(n1185) );
  NAND U1447 ( .A(n1186), .B(n1185), .Z(n1188) );
  XNOR U1448 ( .A(n1189), .B(n1188), .Z(c[1228]) );
  NAND U1449 ( .A(b[0]), .B(a[206]), .Z(n1192) );
  XNOR U1450 ( .A(sreg[1229]), .B(n1192), .Z(n1194) );
  NANDN U1451 ( .A(sreg[1228]), .B(n1187), .Z(n1191) );
  NAND U1452 ( .A(n1189), .B(n1188), .Z(n1190) );
  NAND U1453 ( .A(n1191), .B(n1190), .Z(n1193) );
  XNOR U1454 ( .A(n1194), .B(n1193), .Z(c[1229]) );
  NAND U1455 ( .A(b[0]), .B(a[207]), .Z(n1197) );
  XNOR U1456 ( .A(sreg[1230]), .B(n1197), .Z(n1199) );
  NANDN U1457 ( .A(sreg[1229]), .B(n1192), .Z(n1196) );
  NAND U1458 ( .A(n1194), .B(n1193), .Z(n1195) );
  NAND U1459 ( .A(n1196), .B(n1195), .Z(n1198) );
  XNOR U1460 ( .A(n1199), .B(n1198), .Z(c[1230]) );
  NAND U1461 ( .A(b[0]), .B(a[208]), .Z(n1204) );
  NANDN U1462 ( .A(sreg[1230]), .B(n1197), .Z(n1201) );
  NAND U1463 ( .A(n1199), .B(n1198), .Z(n1200) );
  AND U1464 ( .A(n1201), .B(n1200), .Z(n1203) );
  XOR U1465 ( .A(sreg[1231]), .B(n1203), .Z(n1202) );
  XNOR U1466 ( .A(n1204), .B(n1202), .Z(c[1231]) );
  NAND U1467 ( .A(b[0]), .B(a[209]), .Z(n1205) );
  XNOR U1468 ( .A(sreg[1232]), .B(n1205), .Z(n1206) );
  XOR U1469 ( .A(n1207), .B(n1206), .Z(c[1232]) );
  NAND U1470 ( .A(b[0]), .B(a[210]), .Z(n1210) );
  XNOR U1471 ( .A(sreg[1233]), .B(n1210), .Z(n1212) );
  NANDN U1472 ( .A(n1205), .B(sreg[1232]), .Z(n1209) );
  NAND U1473 ( .A(n1207), .B(n1206), .Z(n1208) );
  NAND U1474 ( .A(n1209), .B(n1208), .Z(n1211) );
  XOR U1475 ( .A(n1212), .B(n1211), .Z(c[1233]) );
  NAND U1476 ( .A(b[0]), .B(a[211]), .Z(n1215) );
  XNOR U1477 ( .A(sreg[1234]), .B(n1215), .Z(n1217) );
  NANDN U1478 ( .A(n1210), .B(sreg[1233]), .Z(n1214) );
  NAND U1479 ( .A(n1212), .B(n1211), .Z(n1213) );
  NAND U1480 ( .A(n1214), .B(n1213), .Z(n1216) );
  XOR U1481 ( .A(n1217), .B(n1216), .Z(c[1234]) );
  NAND U1482 ( .A(b[0]), .B(a[212]), .Z(n1220) );
  XNOR U1483 ( .A(sreg[1235]), .B(n1220), .Z(n1222) );
  NANDN U1484 ( .A(n1215), .B(sreg[1234]), .Z(n1219) );
  NAND U1485 ( .A(n1217), .B(n1216), .Z(n1218) );
  NAND U1486 ( .A(n1219), .B(n1218), .Z(n1221) );
  XOR U1487 ( .A(n1222), .B(n1221), .Z(c[1235]) );
  NAND U1488 ( .A(b[0]), .B(a[213]), .Z(n1225) );
  XNOR U1489 ( .A(sreg[1236]), .B(n1225), .Z(n1227) );
  NANDN U1490 ( .A(n1220), .B(sreg[1235]), .Z(n1224) );
  NAND U1491 ( .A(n1222), .B(n1221), .Z(n1223) );
  NAND U1492 ( .A(n1224), .B(n1223), .Z(n1226) );
  XOR U1493 ( .A(n1227), .B(n1226), .Z(c[1236]) );
  NAND U1494 ( .A(b[0]), .B(a[214]), .Z(n1230) );
  XNOR U1495 ( .A(sreg[1237]), .B(n1230), .Z(n1232) );
  NANDN U1496 ( .A(n1225), .B(sreg[1236]), .Z(n1229) );
  NAND U1497 ( .A(n1227), .B(n1226), .Z(n1228) );
  NAND U1498 ( .A(n1229), .B(n1228), .Z(n1231) );
  XOR U1499 ( .A(n1232), .B(n1231), .Z(c[1237]) );
  NAND U1500 ( .A(b[0]), .B(a[215]), .Z(n1235) );
  XNOR U1501 ( .A(sreg[1238]), .B(n1235), .Z(n1237) );
  NANDN U1502 ( .A(n1230), .B(sreg[1237]), .Z(n1234) );
  NAND U1503 ( .A(n1232), .B(n1231), .Z(n1233) );
  AND U1504 ( .A(n1234), .B(n1233), .Z(n1236) );
  XNOR U1505 ( .A(n1237), .B(n1236), .Z(c[1238]) );
  NANDN U1506 ( .A(sreg[1238]), .B(n1235), .Z(n1239) );
  NAND U1507 ( .A(n1237), .B(n1236), .Z(n1238) );
  AND U1508 ( .A(n1239), .B(n1238), .Z(n1242) );
  NAND U1509 ( .A(b[0]), .B(a[216]), .Z(n1240) );
  XNOR U1510 ( .A(sreg[1239]), .B(n1240), .Z(n1241) );
  XOR U1511 ( .A(n1242), .B(n1241), .Z(c[1239]) );
  NAND U1512 ( .A(b[0]), .B(a[217]), .Z(n1245) );
  XNOR U1513 ( .A(sreg[1240]), .B(n1245), .Z(n1247) );
  NANDN U1514 ( .A(n1240), .B(sreg[1239]), .Z(n1244) );
  NAND U1515 ( .A(n1242), .B(n1241), .Z(n1243) );
  NAND U1516 ( .A(n1244), .B(n1243), .Z(n1246) );
  XOR U1517 ( .A(n1247), .B(n1246), .Z(c[1240]) );
  NAND U1518 ( .A(b[0]), .B(a[218]), .Z(n1252) );
  NANDN U1519 ( .A(n1245), .B(sreg[1240]), .Z(n1249) );
  NAND U1520 ( .A(n1247), .B(n1246), .Z(n1248) );
  NAND U1521 ( .A(n1249), .B(n1248), .Z(n1251) );
  XOR U1522 ( .A(n1251), .B(sreg[1241]), .Z(n1250) );
  XNOR U1523 ( .A(n1252), .B(n1250), .Z(c[1241]) );
  NAND U1524 ( .A(b[0]), .B(a[219]), .Z(n1253) );
  XNOR U1525 ( .A(sreg[1242]), .B(n1253), .Z(n1254) );
  XNOR U1526 ( .A(n1255), .B(n1254), .Z(c[1242]) );
  NAND U1527 ( .A(b[0]), .B(a[220]), .Z(n1258) );
  XNOR U1528 ( .A(sreg[1243]), .B(n1258), .Z(n1260) );
  NANDN U1529 ( .A(n1253), .B(sreg[1242]), .Z(n1257) );
  NANDN U1530 ( .A(n1255), .B(n1254), .Z(n1256) );
  NAND U1531 ( .A(n1257), .B(n1256), .Z(n1259) );
  XOR U1532 ( .A(n1260), .B(n1259), .Z(c[1243]) );
  NANDN U1533 ( .A(n1258), .B(sreg[1243]), .Z(n1262) );
  NAND U1534 ( .A(n1260), .B(n1259), .Z(n1261) );
  NAND U1535 ( .A(n1262), .B(n1261), .Z(n1265) );
  NAND U1536 ( .A(b[0]), .B(a[221]), .Z(n1264) );
  XOR U1537 ( .A(sreg[1244]), .B(n1264), .Z(n1263) );
  XNOR U1538 ( .A(n1265), .B(n1263), .Z(c[1244]) );
  NAND U1539 ( .A(b[0]), .B(a[222]), .Z(n1266) );
  XNOR U1540 ( .A(sreg[1245]), .B(n1266), .Z(n1267) );
  XOR U1541 ( .A(n1268), .B(n1267), .Z(c[1245]) );
  NAND U1542 ( .A(b[0]), .B(a[223]), .Z(n1271) );
  XNOR U1543 ( .A(sreg[1246]), .B(n1271), .Z(n1273) );
  NANDN U1544 ( .A(n1266), .B(sreg[1245]), .Z(n1270) );
  NAND U1545 ( .A(n1268), .B(n1267), .Z(n1269) );
  NAND U1546 ( .A(n1270), .B(n1269), .Z(n1272) );
  XOR U1547 ( .A(n1273), .B(n1272), .Z(c[1246]) );
  AND U1548 ( .A(b[0]), .B(a[224]), .Z(n1277) );
  NANDN U1549 ( .A(n1271), .B(sreg[1246]), .Z(n1275) );
  NAND U1550 ( .A(n1273), .B(n1272), .Z(n1274) );
  AND U1551 ( .A(n1275), .B(n1274), .Z(n1278) );
  XNOR U1552 ( .A(sreg[1247]), .B(n1278), .Z(n1276) );
  XOR U1553 ( .A(n1277), .B(n1276), .Z(c[1247]) );
  NAND U1554 ( .A(b[0]), .B(a[225]), .Z(n1279) );
  XNOR U1555 ( .A(sreg[1248]), .B(n1279), .Z(n1280) );
  XNOR U1556 ( .A(n1281), .B(n1280), .Z(c[1248]) );
  NAND U1557 ( .A(b[0]), .B(a[226]), .Z(n1284) );
  XNOR U1558 ( .A(sreg[1249]), .B(n1284), .Z(n1286) );
  NANDN U1559 ( .A(n1279), .B(sreg[1248]), .Z(n1283) );
  NANDN U1560 ( .A(n1281), .B(n1280), .Z(n1282) );
  NAND U1561 ( .A(n1283), .B(n1282), .Z(n1285) );
  XOR U1562 ( .A(n1286), .B(n1285), .Z(c[1249]) );
  NANDN U1563 ( .A(n1284), .B(sreg[1249]), .Z(n1288) );
  NAND U1564 ( .A(n1286), .B(n1285), .Z(n1287) );
  NAND U1565 ( .A(n1288), .B(n1287), .Z(n1291) );
  NAND U1566 ( .A(b[0]), .B(a[227]), .Z(n1290) );
  XOR U1567 ( .A(sreg[1250]), .B(n1290), .Z(n1289) );
  XNOR U1568 ( .A(n1291), .B(n1289), .Z(c[1250]) );
  NAND U1569 ( .A(b[0]), .B(a[228]), .Z(n1292) );
  XNOR U1570 ( .A(sreg[1251]), .B(n1292), .Z(n1293) );
  XOR U1571 ( .A(n1294), .B(n1293), .Z(c[1251]) );
  NAND U1572 ( .A(b[0]), .B(a[229]), .Z(n1297) );
  XNOR U1573 ( .A(sreg[1252]), .B(n1297), .Z(n1299) );
  NANDN U1574 ( .A(n1292), .B(sreg[1251]), .Z(n1296) );
  NAND U1575 ( .A(n1294), .B(n1293), .Z(n1295) );
  NAND U1576 ( .A(n1296), .B(n1295), .Z(n1298) );
  XOR U1577 ( .A(n1299), .B(n1298), .Z(c[1252]) );
  AND U1578 ( .A(b[0]), .B(a[230]), .Z(n1303) );
  NANDN U1579 ( .A(n1297), .B(sreg[1252]), .Z(n1301) );
  NAND U1580 ( .A(n1299), .B(n1298), .Z(n1300) );
  AND U1581 ( .A(n1301), .B(n1300), .Z(n1304) );
  XNOR U1582 ( .A(sreg[1253]), .B(n1304), .Z(n1302) );
  XOR U1583 ( .A(n1303), .B(n1302), .Z(c[1253]) );
  NAND U1584 ( .A(b[0]), .B(a[231]), .Z(n1305) );
  XNOR U1585 ( .A(sreg[1254]), .B(n1305), .Z(n1306) );
  XNOR U1586 ( .A(n1307), .B(n1306), .Z(c[1254]) );
  AND U1587 ( .A(b[0]), .B(a[232]), .Z(n1312) );
  NANDN U1588 ( .A(sreg[1254]), .B(n1305), .Z(n1309) );
  NAND U1589 ( .A(n1307), .B(n1306), .Z(n1308) );
  NAND U1590 ( .A(n1309), .B(n1308), .Z(n1311) );
  XOR U1591 ( .A(sreg[1255]), .B(n1311), .Z(n1310) );
  XNOR U1592 ( .A(n1312), .B(n1310), .Z(c[1255]) );
  NAND U1593 ( .A(b[0]), .B(a[233]), .Z(n1313) );
  XNOR U1594 ( .A(sreg[1256]), .B(n1313), .Z(n1314) );
  XOR U1595 ( .A(n1315), .B(n1314), .Z(c[1256]) );
  NAND U1596 ( .A(b[0]), .B(a[234]), .Z(n1318) );
  XNOR U1597 ( .A(sreg[1257]), .B(n1318), .Z(n1320) );
  NANDN U1598 ( .A(n1313), .B(sreg[1256]), .Z(n1317) );
  NAND U1599 ( .A(n1315), .B(n1314), .Z(n1316) );
  NAND U1600 ( .A(n1317), .B(n1316), .Z(n1319) );
  XOR U1601 ( .A(n1320), .B(n1319), .Z(c[1257]) );
  NANDN U1602 ( .A(n1318), .B(sreg[1257]), .Z(n1322) );
  NAND U1603 ( .A(n1320), .B(n1319), .Z(n1321) );
  AND U1604 ( .A(n1322), .B(n1321), .Z(n1325) );
  NAND U1605 ( .A(b[0]), .B(a[235]), .Z(n1323) );
  XNOR U1606 ( .A(sreg[1258]), .B(n1323), .Z(n1324) );
  XNOR U1607 ( .A(n1325), .B(n1324), .Z(c[1258]) );
  NAND U1608 ( .A(b[0]), .B(a[236]), .Z(n1328) );
  XNOR U1609 ( .A(sreg[1259]), .B(n1328), .Z(n1330) );
  NANDN U1610 ( .A(sreg[1258]), .B(n1323), .Z(n1327) );
  NAND U1611 ( .A(n1325), .B(n1324), .Z(n1326) );
  NAND U1612 ( .A(n1327), .B(n1326), .Z(n1329) );
  XNOR U1613 ( .A(n1330), .B(n1329), .Z(c[1259]) );
  NAND U1614 ( .A(b[0]), .B(a[237]), .Z(n1333) );
  XNOR U1615 ( .A(sreg[1260]), .B(n1333), .Z(n1335) );
  NANDN U1616 ( .A(sreg[1259]), .B(n1328), .Z(n1332) );
  NAND U1617 ( .A(n1330), .B(n1329), .Z(n1331) );
  NAND U1618 ( .A(n1332), .B(n1331), .Z(n1334) );
  XNOR U1619 ( .A(n1335), .B(n1334), .Z(c[1260]) );
  NAND U1620 ( .A(b[0]), .B(a[238]), .Z(n1338) );
  XNOR U1621 ( .A(sreg[1261]), .B(n1338), .Z(n1340) );
  NANDN U1622 ( .A(sreg[1260]), .B(n1333), .Z(n1337) );
  NAND U1623 ( .A(n1335), .B(n1334), .Z(n1336) );
  NAND U1624 ( .A(n1337), .B(n1336), .Z(n1339) );
  XNOR U1625 ( .A(n1340), .B(n1339), .Z(c[1261]) );
  NAND U1626 ( .A(b[0]), .B(a[239]), .Z(n1343) );
  XNOR U1627 ( .A(sreg[1262]), .B(n1343), .Z(n1345) );
  NANDN U1628 ( .A(sreg[1261]), .B(n1338), .Z(n1342) );
  NAND U1629 ( .A(n1340), .B(n1339), .Z(n1341) );
  NAND U1630 ( .A(n1342), .B(n1341), .Z(n1344) );
  XNOR U1631 ( .A(n1345), .B(n1344), .Z(c[1262]) );
  NAND U1632 ( .A(b[0]), .B(a[240]), .Z(n1348) );
  XNOR U1633 ( .A(sreg[1263]), .B(n1348), .Z(n1350) );
  NANDN U1634 ( .A(sreg[1262]), .B(n1343), .Z(n1347) );
  NAND U1635 ( .A(n1345), .B(n1344), .Z(n1346) );
  NAND U1636 ( .A(n1347), .B(n1346), .Z(n1349) );
  XNOR U1637 ( .A(n1350), .B(n1349), .Z(c[1263]) );
  NAND U1638 ( .A(b[0]), .B(a[241]), .Z(n1353) );
  XNOR U1639 ( .A(sreg[1264]), .B(n1353), .Z(n1355) );
  NANDN U1640 ( .A(sreg[1263]), .B(n1348), .Z(n1352) );
  NAND U1641 ( .A(n1350), .B(n1349), .Z(n1351) );
  NAND U1642 ( .A(n1352), .B(n1351), .Z(n1354) );
  XNOR U1643 ( .A(n1355), .B(n1354), .Z(c[1264]) );
  NAND U1644 ( .A(b[0]), .B(a[242]), .Z(n1358) );
  XNOR U1645 ( .A(sreg[1265]), .B(n1358), .Z(n1360) );
  NANDN U1646 ( .A(sreg[1264]), .B(n1353), .Z(n1357) );
  NAND U1647 ( .A(n1355), .B(n1354), .Z(n1356) );
  AND U1648 ( .A(n1357), .B(n1356), .Z(n1359) );
  XOR U1649 ( .A(n1360), .B(n1359), .Z(c[1265]) );
  NAND U1650 ( .A(b[0]), .B(a[243]), .Z(n1363) );
  XNOR U1651 ( .A(sreg[1266]), .B(n1363), .Z(n1365) );
  NANDN U1652 ( .A(n1358), .B(sreg[1265]), .Z(n1362) );
  NAND U1653 ( .A(n1360), .B(n1359), .Z(n1361) );
  NAND U1654 ( .A(n1362), .B(n1361), .Z(n1364) );
  XOR U1655 ( .A(n1365), .B(n1364), .Z(c[1266]) );
  NAND U1656 ( .A(b[0]), .B(a[244]), .Z(n1368) );
  XNOR U1657 ( .A(sreg[1267]), .B(n1368), .Z(n1370) );
  NANDN U1658 ( .A(n1363), .B(sreg[1266]), .Z(n1367) );
  NAND U1659 ( .A(n1365), .B(n1364), .Z(n1366) );
  AND U1660 ( .A(n1367), .B(n1366), .Z(n1369) );
  XNOR U1661 ( .A(n1370), .B(n1369), .Z(c[1267]) );
  NAND U1662 ( .A(b[0]), .B(a[245]), .Z(n1373) );
  XNOR U1663 ( .A(sreg[1268]), .B(n1373), .Z(n1375) );
  NANDN U1664 ( .A(sreg[1267]), .B(n1368), .Z(n1372) );
  NAND U1665 ( .A(n1370), .B(n1369), .Z(n1371) );
  AND U1666 ( .A(n1372), .B(n1371), .Z(n1374) );
  XOR U1667 ( .A(n1375), .B(n1374), .Z(c[1268]) );
  NAND U1668 ( .A(b[0]), .B(a[246]), .Z(n1378) );
  XNOR U1669 ( .A(sreg[1269]), .B(n1378), .Z(n1380) );
  NANDN U1670 ( .A(n1373), .B(sreg[1268]), .Z(n1377) );
  NAND U1671 ( .A(n1375), .B(n1374), .Z(n1376) );
  NAND U1672 ( .A(n1377), .B(n1376), .Z(n1379) );
  XOR U1673 ( .A(n1380), .B(n1379), .Z(c[1269]) );
  NANDN U1674 ( .A(n1378), .B(sreg[1269]), .Z(n1382) );
  NAND U1675 ( .A(n1380), .B(n1379), .Z(n1381) );
  AND U1676 ( .A(n1382), .B(n1381), .Z(n1385) );
  NAND U1677 ( .A(b[0]), .B(a[247]), .Z(n1383) );
  XNOR U1678 ( .A(sreg[1270]), .B(n1383), .Z(n1384) );
  XNOR U1679 ( .A(n1385), .B(n1384), .Z(c[1270]) );
  NAND U1680 ( .A(b[0]), .B(a[248]), .Z(n1388) );
  XNOR U1681 ( .A(sreg[1271]), .B(n1388), .Z(n1390) );
  NANDN U1682 ( .A(sreg[1270]), .B(n1383), .Z(n1387) );
  NAND U1683 ( .A(n1385), .B(n1384), .Z(n1386) );
  AND U1684 ( .A(n1387), .B(n1386), .Z(n1389) );
  XOR U1685 ( .A(n1390), .B(n1389), .Z(c[1271]) );
  NAND U1686 ( .A(b[0]), .B(a[249]), .Z(n1393) );
  XNOR U1687 ( .A(sreg[1272]), .B(n1393), .Z(n1395) );
  NANDN U1688 ( .A(n1388), .B(sreg[1271]), .Z(n1392) );
  NAND U1689 ( .A(n1390), .B(n1389), .Z(n1391) );
  NAND U1690 ( .A(n1392), .B(n1391), .Z(n1394) );
  XOR U1691 ( .A(n1395), .B(n1394), .Z(c[1272]) );
  NANDN U1692 ( .A(n1393), .B(sreg[1272]), .Z(n1397) );
  NAND U1693 ( .A(n1395), .B(n1394), .Z(n1396) );
  AND U1694 ( .A(n1397), .B(n1396), .Z(n1400) );
  NAND U1695 ( .A(b[0]), .B(a[250]), .Z(n1398) );
  XNOR U1696 ( .A(sreg[1273]), .B(n1398), .Z(n1399) );
  XNOR U1697 ( .A(n1400), .B(n1399), .Z(c[1273]) );
  NAND U1698 ( .A(b[0]), .B(a[251]), .Z(n1403) );
  XNOR U1699 ( .A(sreg[1274]), .B(n1403), .Z(n1405) );
  NANDN U1700 ( .A(sreg[1273]), .B(n1398), .Z(n1402) );
  NAND U1701 ( .A(n1400), .B(n1399), .Z(n1401) );
  NAND U1702 ( .A(n1402), .B(n1401), .Z(n1404) );
  XNOR U1703 ( .A(n1405), .B(n1404), .Z(c[1274]) );
  NAND U1704 ( .A(b[0]), .B(a[252]), .Z(n1408) );
  XNOR U1705 ( .A(sreg[1275]), .B(n1408), .Z(n1410) );
  NANDN U1706 ( .A(sreg[1274]), .B(n1403), .Z(n1407) );
  NAND U1707 ( .A(n1405), .B(n1404), .Z(n1406) );
  NAND U1708 ( .A(n1407), .B(n1406), .Z(n1409) );
  XNOR U1709 ( .A(n1410), .B(n1409), .Z(c[1275]) );
  NAND U1710 ( .A(b[0]), .B(a[253]), .Z(n1413) );
  XNOR U1711 ( .A(sreg[1276]), .B(n1413), .Z(n1415) );
  NANDN U1712 ( .A(sreg[1275]), .B(n1408), .Z(n1412) );
  NAND U1713 ( .A(n1410), .B(n1409), .Z(n1411) );
  NAND U1714 ( .A(n1412), .B(n1411), .Z(n1414) );
  XNOR U1715 ( .A(n1415), .B(n1414), .Z(c[1276]) );
  NAND U1716 ( .A(b[0]), .B(a[254]), .Z(n1418) );
  XNOR U1717 ( .A(sreg[1277]), .B(n1418), .Z(n1420) );
  NANDN U1718 ( .A(sreg[1276]), .B(n1413), .Z(n1417) );
  NAND U1719 ( .A(n1415), .B(n1414), .Z(n1416) );
  NAND U1720 ( .A(n1417), .B(n1416), .Z(n1419) );
  XNOR U1721 ( .A(n1420), .B(n1419), .Z(c[1277]) );
  NAND U1722 ( .A(b[0]), .B(a[255]), .Z(n1423) );
  XNOR U1723 ( .A(sreg[1278]), .B(n1423), .Z(n1425) );
  NANDN U1724 ( .A(sreg[1277]), .B(n1418), .Z(n1422) );
  NAND U1725 ( .A(n1420), .B(n1419), .Z(n1421) );
  NAND U1726 ( .A(n1422), .B(n1421), .Z(n1424) );
  XNOR U1727 ( .A(n1425), .B(n1424), .Z(c[1278]) );
  NAND U1728 ( .A(b[0]), .B(a[256]), .Z(n1428) );
  XNOR U1729 ( .A(sreg[1279]), .B(n1428), .Z(n1430) );
  NANDN U1730 ( .A(sreg[1278]), .B(n1423), .Z(n1427) );
  NAND U1731 ( .A(n1425), .B(n1424), .Z(n1426) );
  NAND U1732 ( .A(n1427), .B(n1426), .Z(n1429) );
  XNOR U1733 ( .A(n1430), .B(n1429), .Z(c[1279]) );
  NAND U1734 ( .A(b[0]), .B(a[257]), .Z(n1433) );
  XNOR U1735 ( .A(sreg[1280]), .B(n1433), .Z(n1435) );
  NANDN U1736 ( .A(sreg[1279]), .B(n1428), .Z(n1432) );
  NAND U1737 ( .A(n1430), .B(n1429), .Z(n1431) );
  NAND U1738 ( .A(n1432), .B(n1431), .Z(n1434) );
  XNOR U1739 ( .A(n1435), .B(n1434), .Z(c[1280]) );
  NAND U1740 ( .A(b[0]), .B(a[258]), .Z(n1438) );
  XNOR U1741 ( .A(sreg[1281]), .B(n1438), .Z(n1440) );
  NANDN U1742 ( .A(sreg[1280]), .B(n1433), .Z(n1437) );
  NAND U1743 ( .A(n1435), .B(n1434), .Z(n1436) );
  NAND U1744 ( .A(n1437), .B(n1436), .Z(n1439) );
  XNOR U1745 ( .A(n1440), .B(n1439), .Z(c[1281]) );
  NANDN U1746 ( .A(sreg[1281]), .B(n1438), .Z(n1442) );
  NAND U1747 ( .A(n1440), .B(n1439), .Z(n1441) );
  AND U1748 ( .A(n1442), .B(n1441), .Z(n1445) );
  NAND U1749 ( .A(b[0]), .B(a[259]), .Z(n1443) );
  XNOR U1750 ( .A(sreg[1282]), .B(n1443), .Z(n1444) );
  XOR U1751 ( .A(n1445), .B(n1444), .Z(c[1282]) );
  NAND U1752 ( .A(b[0]), .B(a[260]), .Z(n1448) );
  XNOR U1753 ( .A(sreg[1283]), .B(n1448), .Z(n1450) );
  NANDN U1754 ( .A(n1443), .B(sreg[1282]), .Z(n1447) );
  NAND U1755 ( .A(n1445), .B(n1444), .Z(n1446) );
  AND U1756 ( .A(n1447), .B(n1446), .Z(n1449) );
  XNOR U1757 ( .A(n1450), .B(n1449), .Z(c[1283]) );
  NAND U1758 ( .A(b[0]), .B(a[261]), .Z(n1453) );
  XNOR U1759 ( .A(sreg[1284]), .B(n1453), .Z(n1455) );
  NANDN U1760 ( .A(sreg[1283]), .B(n1448), .Z(n1452) );
  NAND U1761 ( .A(n1450), .B(n1449), .Z(n1451) );
  NAND U1762 ( .A(n1452), .B(n1451), .Z(n1454) );
  XNOR U1763 ( .A(n1455), .B(n1454), .Z(c[1284]) );
  NANDN U1764 ( .A(sreg[1284]), .B(n1453), .Z(n1457) );
  NAND U1765 ( .A(n1455), .B(n1454), .Z(n1456) );
  AND U1766 ( .A(n1457), .B(n1456), .Z(n1460) );
  NAND U1767 ( .A(b[0]), .B(a[262]), .Z(n1458) );
  XNOR U1768 ( .A(sreg[1285]), .B(n1458), .Z(n1459) );
  XOR U1769 ( .A(n1460), .B(n1459), .Z(c[1285]) );
  NAND U1770 ( .A(b[0]), .B(a[263]), .Z(n1463) );
  XNOR U1771 ( .A(sreg[1286]), .B(n1463), .Z(n1465) );
  NANDN U1772 ( .A(n1458), .B(sreg[1285]), .Z(n1462) );
  NAND U1773 ( .A(n1460), .B(n1459), .Z(n1461) );
  NAND U1774 ( .A(n1462), .B(n1461), .Z(n1464) );
  XOR U1775 ( .A(n1465), .B(n1464), .Z(c[1286]) );
  NAND U1776 ( .A(b[0]), .B(a[264]), .Z(n1470) );
  NANDN U1777 ( .A(n1463), .B(sreg[1286]), .Z(n1467) );
  NAND U1778 ( .A(n1465), .B(n1464), .Z(n1466) );
  NAND U1779 ( .A(n1467), .B(n1466), .Z(n1469) );
  XOR U1780 ( .A(sreg[1287]), .B(n1469), .Z(n1468) );
  XNOR U1781 ( .A(n1470), .B(n1468), .Z(c[1287]) );
  NAND U1782 ( .A(b[0]), .B(a[265]), .Z(n1471) );
  XNOR U1783 ( .A(sreg[1288]), .B(n1471), .Z(n1472) );
  XOR U1784 ( .A(n1473), .B(n1472), .Z(c[1288]) );
  NAND U1785 ( .A(b[0]), .B(a[266]), .Z(n1476) );
  XNOR U1786 ( .A(sreg[1289]), .B(n1476), .Z(n1478) );
  NANDN U1787 ( .A(n1471), .B(sreg[1288]), .Z(n1475) );
  NAND U1788 ( .A(n1473), .B(n1472), .Z(n1474) );
  NAND U1789 ( .A(n1475), .B(n1474), .Z(n1477) );
  XOR U1790 ( .A(n1478), .B(n1477), .Z(c[1289]) );
  NAND U1791 ( .A(b[0]), .B(a[267]), .Z(n1481) );
  XNOR U1792 ( .A(sreg[1290]), .B(n1481), .Z(n1483) );
  NANDN U1793 ( .A(n1476), .B(sreg[1289]), .Z(n1480) );
  NAND U1794 ( .A(n1478), .B(n1477), .Z(n1479) );
  NAND U1795 ( .A(n1480), .B(n1479), .Z(n1482) );
  XOR U1796 ( .A(n1483), .B(n1482), .Z(c[1290]) );
  NAND U1797 ( .A(b[0]), .B(a[268]), .Z(n1486) );
  XNOR U1798 ( .A(sreg[1291]), .B(n1486), .Z(n1488) );
  NANDN U1799 ( .A(n1481), .B(sreg[1290]), .Z(n1485) );
  NAND U1800 ( .A(n1483), .B(n1482), .Z(n1484) );
  NAND U1801 ( .A(n1485), .B(n1484), .Z(n1487) );
  XOR U1802 ( .A(n1488), .B(n1487), .Z(c[1291]) );
  NAND U1803 ( .A(b[0]), .B(a[269]), .Z(n1491) );
  XNOR U1804 ( .A(sreg[1292]), .B(n1491), .Z(n1493) );
  NANDN U1805 ( .A(n1486), .B(sreg[1291]), .Z(n1490) );
  NAND U1806 ( .A(n1488), .B(n1487), .Z(n1489) );
  NAND U1807 ( .A(n1490), .B(n1489), .Z(n1492) );
  XOR U1808 ( .A(n1493), .B(n1492), .Z(c[1292]) );
  NANDN U1809 ( .A(n1491), .B(sreg[1292]), .Z(n1495) );
  NAND U1810 ( .A(n1493), .B(n1492), .Z(n1494) );
  AND U1811 ( .A(n1495), .B(n1494), .Z(n1498) );
  NAND U1812 ( .A(b[0]), .B(a[270]), .Z(n1496) );
  XNOR U1813 ( .A(sreg[1293]), .B(n1496), .Z(n1497) );
  XNOR U1814 ( .A(n1498), .B(n1497), .Z(c[1293]) );
  NANDN U1815 ( .A(sreg[1293]), .B(n1496), .Z(n1500) );
  NAND U1816 ( .A(n1498), .B(n1497), .Z(n1499) );
  AND U1817 ( .A(n1500), .B(n1499), .Z(n1503) );
  NAND U1818 ( .A(b[0]), .B(a[271]), .Z(n1501) );
  XNOR U1819 ( .A(sreg[1294]), .B(n1501), .Z(n1502) );
  XOR U1820 ( .A(n1503), .B(n1502), .Z(c[1294]) );
  NANDN U1821 ( .A(n1501), .B(sreg[1294]), .Z(n1505) );
  NAND U1822 ( .A(n1503), .B(n1502), .Z(n1504) );
  AND U1823 ( .A(n1505), .B(n1504), .Z(n1508) );
  NAND U1824 ( .A(b[0]), .B(a[272]), .Z(n1507) );
  XOR U1825 ( .A(n1507), .B(sreg[1295]), .Z(n1506) );
  XOR U1826 ( .A(n1508), .B(n1506), .Z(c[1295]) );
  NAND U1827 ( .A(b[0]), .B(a[273]), .Z(n1509) );
  XNOR U1828 ( .A(sreg[1296]), .B(n1509), .Z(n1510) );
  XOR U1829 ( .A(n1511), .B(n1510), .Z(c[1296]) );
  NAND U1830 ( .A(b[0]), .B(a[274]), .Z(n1514) );
  XNOR U1831 ( .A(sreg[1297]), .B(n1514), .Z(n1516) );
  NANDN U1832 ( .A(n1509), .B(sreg[1296]), .Z(n1513) );
  NAND U1833 ( .A(n1511), .B(n1510), .Z(n1512) );
  NAND U1834 ( .A(n1513), .B(n1512), .Z(n1515) );
  XOR U1835 ( .A(n1516), .B(n1515), .Z(c[1297]) );
  NANDN U1836 ( .A(n1514), .B(sreg[1297]), .Z(n1518) );
  NAND U1837 ( .A(n1516), .B(n1515), .Z(n1517) );
  AND U1838 ( .A(n1518), .B(n1517), .Z(n1521) );
  NAND U1839 ( .A(b[0]), .B(a[275]), .Z(n1519) );
  XNOR U1840 ( .A(sreg[1298]), .B(n1519), .Z(n1520) );
  XNOR U1841 ( .A(n1521), .B(n1520), .Z(c[1298]) );
  NAND U1842 ( .A(b[0]), .B(a[276]), .Z(n1524) );
  XNOR U1843 ( .A(sreg[1299]), .B(n1524), .Z(n1526) );
  NANDN U1844 ( .A(sreg[1298]), .B(n1519), .Z(n1523) );
  NAND U1845 ( .A(n1521), .B(n1520), .Z(n1522) );
  AND U1846 ( .A(n1523), .B(n1522), .Z(n1525) );
  XOR U1847 ( .A(n1526), .B(n1525), .Z(c[1299]) );
  NANDN U1848 ( .A(n1524), .B(sreg[1299]), .Z(n1528) );
  NAND U1849 ( .A(n1526), .B(n1525), .Z(n1527) );
  AND U1850 ( .A(n1528), .B(n1527), .Z(n1531) );
  NAND U1851 ( .A(b[0]), .B(a[277]), .Z(n1529) );
  XNOR U1852 ( .A(sreg[1300]), .B(n1529), .Z(n1530) );
  XNOR U1853 ( .A(n1531), .B(n1530), .Z(c[1300]) );
  NAND U1854 ( .A(b[0]), .B(a[278]), .Z(n1534) );
  XNOR U1855 ( .A(sreg[1301]), .B(n1534), .Z(n1536) );
  NANDN U1856 ( .A(sreg[1300]), .B(n1529), .Z(n1533) );
  NAND U1857 ( .A(n1531), .B(n1530), .Z(n1532) );
  NAND U1858 ( .A(n1533), .B(n1532), .Z(n1535) );
  XNOR U1859 ( .A(n1536), .B(n1535), .Z(c[1301]) );
  NAND U1860 ( .A(b[0]), .B(a[279]), .Z(n1539) );
  XNOR U1861 ( .A(sreg[1302]), .B(n1539), .Z(n1541) );
  NANDN U1862 ( .A(sreg[1301]), .B(n1534), .Z(n1538) );
  NAND U1863 ( .A(n1536), .B(n1535), .Z(n1537) );
  AND U1864 ( .A(n1538), .B(n1537), .Z(n1540) );
  XOR U1865 ( .A(n1541), .B(n1540), .Z(c[1302]) );
  NANDN U1866 ( .A(n1539), .B(sreg[1302]), .Z(n1543) );
  NAND U1867 ( .A(n1541), .B(n1540), .Z(n1542) );
  AND U1868 ( .A(n1543), .B(n1542), .Z(n1546) );
  NAND U1869 ( .A(b[0]), .B(a[280]), .Z(n1544) );
  XNOR U1870 ( .A(sreg[1303]), .B(n1544), .Z(n1545) );
  XNOR U1871 ( .A(n1546), .B(n1545), .Z(c[1303]) );
  NAND U1872 ( .A(b[0]), .B(a[281]), .Z(n1549) );
  XNOR U1873 ( .A(sreg[1304]), .B(n1549), .Z(n1551) );
  NANDN U1874 ( .A(sreg[1303]), .B(n1544), .Z(n1548) );
  NAND U1875 ( .A(n1546), .B(n1545), .Z(n1547) );
  NAND U1876 ( .A(n1548), .B(n1547), .Z(n1550) );
  XNOR U1877 ( .A(n1551), .B(n1550), .Z(c[1304]) );
  NAND U1878 ( .A(b[0]), .B(a[282]), .Z(n1554) );
  XNOR U1879 ( .A(sreg[1305]), .B(n1554), .Z(n1556) );
  NANDN U1880 ( .A(sreg[1304]), .B(n1549), .Z(n1553) );
  NAND U1881 ( .A(n1551), .B(n1550), .Z(n1552) );
  AND U1882 ( .A(n1553), .B(n1552), .Z(n1555) );
  XOR U1883 ( .A(n1556), .B(n1555), .Z(c[1305]) );
  NANDN U1884 ( .A(n1554), .B(sreg[1305]), .Z(n1558) );
  NAND U1885 ( .A(n1556), .B(n1555), .Z(n1557) );
  AND U1886 ( .A(n1558), .B(n1557), .Z(n1561) );
  NAND U1887 ( .A(b[0]), .B(a[283]), .Z(n1559) );
  XNOR U1888 ( .A(sreg[1306]), .B(n1559), .Z(n1560) );
  XNOR U1889 ( .A(n1561), .B(n1560), .Z(c[1306]) );
  NANDN U1890 ( .A(sreg[1306]), .B(n1559), .Z(n1563) );
  NAND U1891 ( .A(n1561), .B(n1560), .Z(n1562) );
  AND U1892 ( .A(n1563), .B(n1562), .Z(n1566) );
  NAND U1893 ( .A(b[0]), .B(a[284]), .Z(n1564) );
  XNOR U1894 ( .A(sreg[1307]), .B(n1564), .Z(n1565) );
  XOR U1895 ( .A(n1566), .B(n1565), .Z(c[1307]) );
  NAND U1896 ( .A(b[0]), .B(a[285]), .Z(n1569) );
  XNOR U1897 ( .A(sreg[1308]), .B(n1569), .Z(n1571) );
  NANDN U1898 ( .A(n1564), .B(sreg[1307]), .Z(n1568) );
  NAND U1899 ( .A(n1566), .B(n1565), .Z(n1567) );
  NAND U1900 ( .A(n1568), .B(n1567), .Z(n1570) );
  XOR U1901 ( .A(n1571), .B(n1570), .Z(c[1308]) );
  NAND U1902 ( .A(b[0]), .B(a[286]), .Z(n1574) );
  XNOR U1903 ( .A(sreg[1309]), .B(n1574), .Z(n1576) );
  NANDN U1904 ( .A(n1569), .B(sreg[1308]), .Z(n1573) );
  NAND U1905 ( .A(n1571), .B(n1570), .Z(n1572) );
  AND U1906 ( .A(n1573), .B(n1572), .Z(n1575) );
  XNOR U1907 ( .A(n1576), .B(n1575), .Z(c[1309]) );
  NAND U1908 ( .A(b[0]), .B(a[287]), .Z(n1579) );
  XNOR U1909 ( .A(sreg[1310]), .B(n1579), .Z(n1581) );
  NANDN U1910 ( .A(sreg[1309]), .B(n1574), .Z(n1578) );
  NAND U1911 ( .A(n1576), .B(n1575), .Z(n1577) );
  AND U1912 ( .A(n1578), .B(n1577), .Z(n1580) );
  XOR U1913 ( .A(n1581), .B(n1580), .Z(c[1310]) );
  NAND U1914 ( .A(b[0]), .B(a[288]), .Z(n1584) );
  XNOR U1915 ( .A(sreg[1311]), .B(n1584), .Z(n1586) );
  NANDN U1916 ( .A(n1579), .B(sreg[1310]), .Z(n1583) );
  NAND U1917 ( .A(n1581), .B(n1580), .Z(n1582) );
  NAND U1918 ( .A(n1583), .B(n1582), .Z(n1585) );
  XOR U1919 ( .A(n1586), .B(n1585), .Z(c[1311]) );
  NAND U1920 ( .A(b[0]), .B(a[289]), .Z(n1589) );
  XNOR U1921 ( .A(sreg[1312]), .B(n1589), .Z(n1591) );
  NANDN U1922 ( .A(n1584), .B(sreg[1311]), .Z(n1588) );
  NAND U1923 ( .A(n1586), .B(n1585), .Z(n1587) );
  NAND U1924 ( .A(n1588), .B(n1587), .Z(n1590) );
  XOR U1925 ( .A(n1591), .B(n1590), .Z(c[1312]) );
  NAND U1926 ( .A(b[0]), .B(a[290]), .Z(n1594) );
  XNOR U1927 ( .A(sreg[1313]), .B(n1594), .Z(n1596) );
  NANDN U1928 ( .A(n1589), .B(sreg[1312]), .Z(n1593) );
  NAND U1929 ( .A(n1591), .B(n1590), .Z(n1592) );
  AND U1930 ( .A(n1593), .B(n1592), .Z(n1595) );
  XNOR U1931 ( .A(n1596), .B(n1595), .Z(c[1313]) );
  NANDN U1932 ( .A(sreg[1313]), .B(n1594), .Z(n1598) );
  NAND U1933 ( .A(n1596), .B(n1595), .Z(n1597) );
  AND U1934 ( .A(n1598), .B(n1597), .Z(n1601) );
  NAND U1935 ( .A(b[0]), .B(a[291]), .Z(n1599) );
  XNOR U1936 ( .A(sreg[1314]), .B(n1599), .Z(n1600) );
  XOR U1937 ( .A(n1601), .B(n1600), .Z(c[1314]) );
  NAND U1938 ( .A(b[0]), .B(a[292]), .Z(n1604) );
  XNOR U1939 ( .A(sreg[1315]), .B(n1604), .Z(n1606) );
  NANDN U1940 ( .A(n1599), .B(sreg[1314]), .Z(n1603) );
  NAND U1941 ( .A(n1601), .B(n1600), .Z(n1602) );
  NAND U1942 ( .A(n1603), .B(n1602), .Z(n1605) );
  XOR U1943 ( .A(n1606), .B(n1605), .Z(c[1315]) );
  NAND U1944 ( .A(b[0]), .B(a[293]), .Z(n1609) );
  XNOR U1945 ( .A(sreg[1316]), .B(n1609), .Z(n1611) );
  NANDN U1946 ( .A(n1604), .B(sreg[1315]), .Z(n1608) );
  NAND U1947 ( .A(n1606), .B(n1605), .Z(n1607) );
  NAND U1948 ( .A(n1608), .B(n1607), .Z(n1610) );
  XOR U1949 ( .A(n1611), .B(n1610), .Z(c[1316]) );
  NAND U1950 ( .A(b[0]), .B(a[294]), .Z(n1614) );
  XNOR U1951 ( .A(sreg[1317]), .B(n1614), .Z(n1616) );
  NANDN U1952 ( .A(n1609), .B(sreg[1316]), .Z(n1613) );
  NAND U1953 ( .A(n1611), .B(n1610), .Z(n1612) );
  NAND U1954 ( .A(n1613), .B(n1612), .Z(n1615) );
  XOR U1955 ( .A(n1616), .B(n1615), .Z(c[1317]) );
  NAND U1956 ( .A(b[0]), .B(a[295]), .Z(n1619) );
  XNOR U1957 ( .A(sreg[1318]), .B(n1619), .Z(n1621) );
  NANDN U1958 ( .A(n1614), .B(sreg[1317]), .Z(n1618) );
  NAND U1959 ( .A(n1616), .B(n1615), .Z(n1617) );
  NAND U1960 ( .A(n1618), .B(n1617), .Z(n1620) );
  XOR U1961 ( .A(n1621), .B(n1620), .Z(c[1318]) );
  NAND U1962 ( .A(b[0]), .B(a[296]), .Z(n1624) );
  XNOR U1963 ( .A(sreg[1319]), .B(n1624), .Z(n1626) );
  NANDN U1964 ( .A(n1619), .B(sreg[1318]), .Z(n1623) );
  NAND U1965 ( .A(n1621), .B(n1620), .Z(n1622) );
  NAND U1966 ( .A(n1623), .B(n1622), .Z(n1625) );
  XOR U1967 ( .A(n1626), .B(n1625), .Z(c[1319]) );
  NAND U1968 ( .A(b[0]), .B(a[297]), .Z(n1629) );
  XNOR U1969 ( .A(sreg[1320]), .B(n1629), .Z(n1631) );
  NANDN U1970 ( .A(n1624), .B(sreg[1319]), .Z(n1628) );
  NAND U1971 ( .A(n1626), .B(n1625), .Z(n1627) );
  NAND U1972 ( .A(n1628), .B(n1627), .Z(n1630) );
  XOR U1973 ( .A(n1631), .B(n1630), .Z(c[1320]) );
  NAND U1974 ( .A(b[0]), .B(a[298]), .Z(n1634) );
  XNOR U1975 ( .A(sreg[1321]), .B(n1634), .Z(n1636) );
  NANDN U1976 ( .A(n1629), .B(sreg[1320]), .Z(n1633) );
  NAND U1977 ( .A(n1631), .B(n1630), .Z(n1632) );
  NAND U1978 ( .A(n1633), .B(n1632), .Z(n1635) );
  XOR U1979 ( .A(n1636), .B(n1635), .Z(c[1321]) );
  NAND U1980 ( .A(b[0]), .B(a[299]), .Z(n1639) );
  XNOR U1981 ( .A(sreg[1322]), .B(n1639), .Z(n1641) );
  NANDN U1982 ( .A(n1634), .B(sreg[1321]), .Z(n1638) );
  NAND U1983 ( .A(n1636), .B(n1635), .Z(n1637) );
  NAND U1984 ( .A(n1638), .B(n1637), .Z(n1640) );
  XOR U1985 ( .A(n1641), .B(n1640), .Z(c[1322]) );
  NAND U1986 ( .A(b[0]), .B(a[300]), .Z(n1644) );
  XNOR U1987 ( .A(sreg[1323]), .B(n1644), .Z(n1646) );
  NANDN U1988 ( .A(n1639), .B(sreg[1322]), .Z(n1643) );
  NAND U1989 ( .A(n1641), .B(n1640), .Z(n1642) );
  AND U1990 ( .A(n1643), .B(n1642), .Z(n1645) );
  XNOR U1991 ( .A(n1646), .B(n1645), .Z(c[1323]) );
  NAND U1992 ( .A(b[0]), .B(a[301]), .Z(n1649) );
  XNOR U1993 ( .A(sreg[1324]), .B(n1649), .Z(n1651) );
  NANDN U1994 ( .A(sreg[1323]), .B(n1644), .Z(n1648) );
  NAND U1995 ( .A(n1646), .B(n1645), .Z(n1647) );
  AND U1996 ( .A(n1648), .B(n1647), .Z(n1650) );
  XOR U1997 ( .A(n1651), .B(n1650), .Z(c[1324]) );
  NANDN U1998 ( .A(n1649), .B(sreg[1324]), .Z(n1653) );
  NAND U1999 ( .A(n1651), .B(n1650), .Z(n1652) );
  AND U2000 ( .A(n1653), .B(n1652), .Z(n1656) );
  NAND U2001 ( .A(b[0]), .B(a[302]), .Z(n1654) );
  XNOR U2002 ( .A(sreg[1325]), .B(n1654), .Z(n1655) );
  XNOR U2003 ( .A(n1656), .B(n1655), .Z(c[1325]) );
  NANDN U2004 ( .A(sreg[1325]), .B(n1654), .Z(n1658) );
  NAND U2005 ( .A(n1656), .B(n1655), .Z(n1657) );
  AND U2006 ( .A(n1658), .B(n1657), .Z(n1661) );
  NAND U2007 ( .A(b[0]), .B(a[303]), .Z(n1659) );
  XNOR U2008 ( .A(sreg[1326]), .B(n1659), .Z(n1660) );
  XOR U2009 ( .A(n1661), .B(n1660), .Z(c[1326]) );
  NANDN U2010 ( .A(n1659), .B(sreg[1326]), .Z(n1663) );
  NAND U2011 ( .A(n1661), .B(n1660), .Z(n1662) );
  AND U2012 ( .A(n1663), .B(n1662), .Z(n1665) );
  AND U2013 ( .A(b[0]), .B(a[304]), .Z(n1666) );
  XNOR U2014 ( .A(sreg[1327]), .B(n1666), .Z(n1664) );
  XOR U2015 ( .A(n1665), .B(n1664), .Z(c[1327]) );
  NAND U2016 ( .A(b[0]), .B(a[305]), .Z(n1667) );
  XNOR U2017 ( .A(sreg[1328]), .B(n1667), .Z(n1669) );
  XOR U2018 ( .A(n1669), .B(n1668), .Z(c[1328]) );
  NAND U2019 ( .A(b[0]), .B(a[306]), .Z(n1672) );
  XNOR U2020 ( .A(sreg[1329]), .B(n1672), .Z(n1674) );
  NANDN U2021 ( .A(n1667), .B(sreg[1328]), .Z(n1671) );
  NAND U2022 ( .A(n1669), .B(n1668), .Z(n1670) );
  NAND U2023 ( .A(n1671), .B(n1670), .Z(n1673) );
  XOR U2024 ( .A(n1674), .B(n1673), .Z(c[1329]) );
  NANDN U2025 ( .A(n1672), .B(sreg[1329]), .Z(n1676) );
  NAND U2026 ( .A(n1674), .B(n1673), .Z(n1675) );
  NAND U2027 ( .A(n1676), .B(n1675), .Z(n1679) );
  NAND U2028 ( .A(b[0]), .B(a[307]), .Z(n1678) );
  XOR U2029 ( .A(sreg[1330]), .B(n1678), .Z(n1677) );
  XNOR U2030 ( .A(n1679), .B(n1677), .Z(c[1330]) );
  NAND U2031 ( .A(b[0]), .B(a[308]), .Z(n1680) );
  XNOR U2032 ( .A(sreg[1331]), .B(n1680), .Z(n1681) );
  XOR U2033 ( .A(n1682), .B(n1681), .Z(c[1331]) );
  NAND U2034 ( .A(b[0]), .B(a[309]), .Z(n1685) );
  XNOR U2035 ( .A(sreg[1332]), .B(n1685), .Z(n1687) );
  NANDN U2036 ( .A(sreg[1331]), .B(n1680), .Z(n1684) );
  NANDN U2037 ( .A(n1682), .B(n1681), .Z(n1683) );
  NAND U2038 ( .A(n1684), .B(n1683), .Z(n1686) );
  XNOR U2039 ( .A(n1687), .B(n1686), .Z(c[1332]) );
  NAND U2040 ( .A(b[0]), .B(a[310]), .Z(n1690) );
  XNOR U2041 ( .A(sreg[1333]), .B(n1690), .Z(n1692) );
  NANDN U2042 ( .A(sreg[1332]), .B(n1685), .Z(n1689) );
  NAND U2043 ( .A(n1687), .B(n1686), .Z(n1688) );
  NAND U2044 ( .A(n1689), .B(n1688), .Z(n1691) );
  XNOR U2045 ( .A(n1692), .B(n1691), .Z(c[1333]) );
  NAND U2046 ( .A(b[0]), .B(a[311]), .Z(n1695) );
  XNOR U2047 ( .A(sreg[1334]), .B(n1695), .Z(n1697) );
  NANDN U2048 ( .A(sreg[1333]), .B(n1690), .Z(n1694) );
  NAND U2049 ( .A(n1692), .B(n1691), .Z(n1693) );
  NAND U2050 ( .A(n1694), .B(n1693), .Z(n1696) );
  XNOR U2051 ( .A(n1697), .B(n1696), .Z(c[1334]) );
  NAND U2052 ( .A(b[0]), .B(a[312]), .Z(n1700) );
  XNOR U2053 ( .A(sreg[1335]), .B(n1700), .Z(n1702) );
  NANDN U2054 ( .A(sreg[1334]), .B(n1695), .Z(n1699) );
  NAND U2055 ( .A(n1697), .B(n1696), .Z(n1698) );
  NAND U2056 ( .A(n1699), .B(n1698), .Z(n1701) );
  XNOR U2057 ( .A(n1702), .B(n1701), .Z(c[1335]) );
  NAND U2058 ( .A(b[0]), .B(a[313]), .Z(n1705) );
  XNOR U2059 ( .A(sreg[1336]), .B(n1705), .Z(n1707) );
  NANDN U2060 ( .A(sreg[1335]), .B(n1700), .Z(n1704) );
  NAND U2061 ( .A(n1702), .B(n1701), .Z(n1703) );
  NAND U2062 ( .A(n1704), .B(n1703), .Z(n1706) );
  XNOR U2063 ( .A(n1707), .B(n1706), .Z(c[1336]) );
  NAND U2064 ( .A(b[0]), .B(a[314]), .Z(n1710) );
  XNOR U2065 ( .A(sreg[1337]), .B(n1710), .Z(n1712) );
  NANDN U2066 ( .A(sreg[1336]), .B(n1705), .Z(n1709) );
  NAND U2067 ( .A(n1707), .B(n1706), .Z(n1708) );
  NAND U2068 ( .A(n1709), .B(n1708), .Z(n1711) );
  XNOR U2069 ( .A(n1712), .B(n1711), .Z(c[1337]) );
  AND U2070 ( .A(b[0]), .B(a[315]), .Z(n1717) );
  NANDN U2071 ( .A(sreg[1337]), .B(n1710), .Z(n1714) );
  NAND U2072 ( .A(n1712), .B(n1711), .Z(n1713) );
  NAND U2073 ( .A(n1714), .B(n1713), .Z(n1716) );
  XOR U2074 ( .A(sreg[1338]), .B(n1716), .Z(n1715) );
  XNOR U2075 ( .A(n1717), .B(n1715), .Z(c[1338]) );
  NAND U2076 ( .A(b[0]), .B(a[316]), .Z(n1718) );
  XNOR U2077 ( .A(sreg[1339]), .B(n1718), .Z(n1719) );
  XOR U2078 ( .A(n1720), .B(n1719), .Z(c[1339]) );
  NAND U2079 ( .A(b[0]), .B(a[317]), .Z(n1723) );
  XNOR U2080 ( .A(sreg[1340]), .B(n1723), .Z(n1725) );
  NANDN U2081 ( .A(n1718), .B(sreg[1339]), .Z(n1722) );
  NAND U2082 ( .A(n1720), .B(n1719), .Z(n1721) );
  NAND U2083 ( .A(n1722), .B(n1721), .Z(n1724) );
  XOR U2084 ( .A(n1725), .B(n1724), .Z(c[1340]) );
  NANDN U2085 ( .A(n1723), .B(sreg[1340]), .Z(n1727) );
  NAND U2086 ( .A(n1725), .B(n1724), .Z(n1726) );
  AND U2087 ( .A(n1727), .B(n1726), .Z(n1730) );
  NAND U2088 ( .A(b[0]), .B(a[318]), .Z(n1728) );
  XNOR U2089 ( .A(sreg[1341]), .B(n1728), .Z(n1729) );
  XNOR U2090 ( .A(n1730), .B(n1729), .Z(c[1341]) );
  NAND U2091 ( .A(b[0]), .B(a[319]), .Z(n1733) );
  XNOR U2092 ( .A(sreg[1342]), .B(n1733), .Z(n1735) );
  NANDN U2093 ( .A(sreg[1341]), .B(n1728), .Z(n1732) );
  NAND U2094 ( .A(n1730), .B(n1729), .Z(n1731) );
  AND U2095 ( .A(n1732), .B(n1731), .Z(n1734) );
  XOR U2096 ( .A(n1735), .B(n1734), .Z(c[1342]) );
  NAND U2097 ( .A(b[0]), .B(a[320]), .Z(n1738) );
  XNOR U2098 ( .A(sreg[1343]), .B(n1738), .Z(n1740) );
  NANDN U2099 ( .A(n1733), .B(sreg[1342]), .Z(n1737) );
  NAND U2100 ( .A(n1735), .B(n1734), .Z(n1736) );
  NAND U2101 ( .A(n1737), .B(n1736), .Z(n1739) );
  XOR U2102 ( .A(n1740), .B(n1739), .Z(c[1343]) );
  NANDN U2103 ( .A(n1738), .B(sreg[1343]), .Z(n1742) );
  NAND U2104 ( .A(n1740), .B(n1739), .Z(n1741) );
  AND U2105 ( .A(n1742), .B(n1741), .Z(n1745) );
  NAND U2106 ( .A(b[0]), .B(a[321]), .Z(n1743) );
  XNOR U2107 ( .A(sreg[1344]), .B(n1743), .Z(n1744) );
  XNOR U2108 ( .A(n1745), .B(n1744), .Z(c[1344]) );
  NAND U2109 ( .A(b[0]), .B(a[322]), .Z(n1748) );
  XNOR U2110 ( .A(sreg[1345]), .B(n1748), .Z(n1750) );
  NANDN U2111 ( .A(sreg[1344]), .B(n1743), .Z(n1747) );
  NAND U2112 ( .A(n1745), .B(n1744), .Z(n1746) );
  AND U2113 ( .A(n1747), .B(n1746), .Z(n1749) );
  XOR U2114 ( .A(n1750), .B(n1749), .Z(c[1345]) );
  NAND U2115 ( .A(b[0]), .B(a[323]), .Z(n1753) );
  XNOR U2116 ( .A(sreg[1346]), .B(n1753), .Z(n1755) );
  NANDN U2117 ( .A(n1748), .B(sreg[1345]), .Z(n1752) );
  NAND U2118 ( .A(n1750), .B(n1749), .Z(n1751) );
  NAND U2119 ( .A(n1752), .B(n1751), .Z(n1754) );
  XOR U2120 ( .A(n1755), .B(n1754), .Z(c[1346]) );
  AND U2121 ( .A(b[0]), .B(a[324]), .Z(n1759) );
  NANDN U2122 ( .A(n1753), .B(sreg[1346]), .Z(n1757) );
  NAND U2123 ( .A(n1755), .B(n1754), .Z(n1756) );
  AND U2124 ( .A(n1757), .B(n1756), .Z(n1760) );
  XNOR U2125 ( .A(sreg[1347]), .B(n1760), .Z(n1758) );
  XOR U2126 ( .A(n1759), .B(n1758), .Z(c[1347]) );
  NAND U2127 ( .A(b[0]), .B(a[325]), .Z(n1761) );
  XNOR U2128 ( .A(sreg[1348]), .B(n1761), .Z(n1762) );
  XNOR U2129 ( .A(n1763), .B(n1762), .Z(c[1348]) );
  NAND U2130 ( .A(b[0]), .B(a[326]), .Z(n1766) );
  XNOR U2131 ( .A(sreg[1349]), .B(n1766), .Z(n1768) );
  NANDN U2132 ( .A(n1761), .B(sreg[1348]), .Z(n1765) );
  NANDN U2133 ( .A(n1763), .B(n1762), .Z(n1764) );
  NAND U2134 ( .A(n1765), .B(n1764), .Z(n1767) );
  XOR U2135 ( .A(n1768), .B(n1767), .Z(c[1349]) );
  NAND U2136 ( .A(b[0]), .B(a[327]), .Z(n1771) );
  XNOR U2137 ( .A(sreg[1350]), .B(n1771), .Z(n1773) );
  NANDN U2138 ( .A(n1766), .B(sreg[1349]), .Z(n1770) );
  NAND U2139 ( .A(n1768), .B(n1767), .Z(n1769) );
  NAND U2140 ( .A(n1770), .B(n1769), .Z(n1772) );
  XOR U2141 ( .A(n1773), .B(n1772), .Z(c[1350]) );
  NAND U2142 ( .A(b[0]), .B(a[328]), .Z(n1776) );
  XNOR U2143 ( .A(sreg[1351]), .B(n1776), .Z(n1778) );
  NANDN U2144 ( .A(n1771), .B(sreg[1350]), .Z(n1775) );
  NAND U2145 ( .A(n1773), .B(n1772), .Z(n1774) );
  NAND U2146 ( .A(n1775), .B(n1774), .Z(n1777) );
  XOR U2147 ( .A(n1778), .B(n1777), .Z(c[1351]) );
  NAND U2148 ( .A(b[0]), .B(a[329]), .Z(n1781) );
  XNOR U2149 ( .A(sreg[1352]), .B(n1781), .Z(n1783) );
  NANDN U2150 ( .A(n1776), .B(sreg[1351]), .Z(n1780) );
  NAND U2151 ( .A(n1778), .B(n1777), .Z(n1779) );
  NAND U2152 ( .A(n1780), .B(n1779), .Z(n1782) );
  XOR U2153 ( .A(n1783), .B(n1782), .Z(c[1352]) );
  NAND U2154 ( .A(b[0]), .B(a[330]), .Z(n1786) );
  XNOR U2155 ( .A(sreg[1353]), .B(n1786), .Z(n1788) );
  NANDN U2156 ( .A(n1781), .B(sreg[1352]), .Z(n1785) );
  NAND U2157 ( .A(n1783), .B(n1782), .Z(n1784) );
  NAND U2158 ( .A(n1785), .B(n1784), .Z(n1787) );
  XOR U2159 ( .A(n1788), .B(n1787), .Z(c[1353]) );
  NAND U2160 ( .A(b[0]), .B(a[331]), .Z(n1791) );
  XNOR U2161 ( .A(sreg[1354]), .B(n1791), .Z(n1793) );
  NANDN U2162 ( .A(n1786), .B(sreg[1353]), .Z(n1790) );
  NAND U2163 ( .A(n1788), .B(n1787), .Z(n1789) );
  NAND U2164 ( .A(n1790), .B(n1789), .Z(n1792) );
  XOR U2165 ( .A(n1793), .B(n1792), .Z(c[1354]) );
  NAND U2166 ( .A(b[0]), .B(a[332]), .Z(n1796) );
  XNOR U2167 ( .A(sreg[1355]), .B(n1796), .Z(n1798) );
  NANDN U2168 ( .A(n1791), .B(sreg[1354]), .Z(n1795) );
  NAND U2169 ( .A(n1793), .B(n1792), .Z(n1794) );
  NAND U2170 ( .A(n1795), .B(n1794), .Z(n1797) );
  XOR U2171 ( .A(n1798), .B(n1797), .Z(c[1355]) );
  NAND U2172 ( .A(b[0]), .B(a[333]), .Z(n1801) );
  XNOR U2173 ( .A(sreg[1356]), .B(n1801), .Z(n1803) );
  NANDN U2174 ( .A(n1796), .B(sreg[1355]), .Z(n1800) );
  NAND U2175 ( .A(n1798), .B(n1797), .Z(n1799) );
  NAND U2176 ( .A(n1800), .B(n1799), .Z(n1802) );
  XOR U2177 ( .A(n1803), .B(n1802), .Z(c[1356]) );
  NAND U2178 ( .A(b[0]), .B(a[334]), .Z(n1806) );
  XNOR U2179 ( .A(sreg[1357]), .B(n1806), .Z(n1808) );
  NANDN U2180 ( .A(n1801), .B(sreg[1356]), .Z(n1805) );
  NAND U2181 ( .A(n1803), .B(n1802), .Z(n1804) );
  NAND U2182 ( .A(n1805), .B(n1804), .Z(n1807) );
  XOR U2183 ( .A(n1808), .B(n1807), .Z(c[1357]) );
  NAND U2184 ( .A(b[0]), .B(a[335]), .Z(n1811) );
  XNOR U2185 ( .A(sreg[1358]), .B(n1811), .Z(n1813) );
  NANDN U2186 ( .A(n1806), .B(sreg[1357]), .Z(n1810) );
  NAND U2187 ( .A(n1808), .B(n1807), .Z(n1809) );
  NAND U2188 ( .A(n1810), .B(n1809), .Z(n1812) );
  XOR U2189 ( .A(n1813), .B(n1812), .Z(c[1358]) );
  NAND U2190 ( .A(b[0]), .B(a[336]), .Z(n1816) );
  XNOR U2191 ( .A(sreg[1359]), .B(n1816), .Z(n1818) );
  NANDN U2192 ( .A(n1811), .B(sreg[1358]), .Z(n1815) );
  NAND U2193 ( .A(n1813), .B(n1812), .Z(n1814) );
  NAND U2194 ( .A(n1815), .B(n1814), .Z(n1817) );
  XOR U2195 ( .A(n1818), .B(n1817), .Z(c[1359]) );
  NANDN U2196 ( .A(n1816), .B(sreg[1359]), .Z(n1820) );
  NAND U2197 ( .A(n1818), .B(n1817), .Z(n1819) );
  AND U2198 ( .A(n1820), .B(n1819), .Z(n1823) );
  NAND U2199 ( .A(b[0]), .B(a[337]), .Z(n1821) );
  XNOR U2200 ( .A(sreg[1360]), .B(n1821), .Z(n1822) );
  XNOR U2201 ( .A(n1823), .B(n1822), .Z(c[1360]) );
  NAND U2202 ( .A(b[0]), .B(a[338]), .Z(n1826) );
  XNOR U2203 ( .A(sreg[1361]), .B(n1826), .Z(n1828) );
  NANDN U2204 ( .A(sreg[1360]), .B(n1821), .Z(n1825) );
  NAND U2205 ( .A(n1823), .B(n1822), .Z(n1824) );
  NAND U2206 ( .A(n1825), .B(n1824), .Z(n1827) );
  XNOR U2207 ( .A(n1828), .B(n1827), .Z(c[1361]) );
  NAND U2208 ( .A(b[0]), .B(a[339]), .Z(n1831) );
  XNOR U2209 ( .A(sreg[1362]), .B(n1831), .Z(n1833) );
  NANDN U2210 ( .A(sreg[1361]), .B(n1826), .Z(n1830) );
  NAND U2211 ( .A(n1828), .B(n1827), .Z(n1829) );
  AND U2212 ( .A(n1830), .B(n1829), .Z(n1832) );
  XOR U2213 ( .A(n1833), .B(n1832), .Z(c[1362]) );
  NANDN U2214 ( .A(n1831), .B(sreg[1362]), .Z(n1835) );
  NAND U2215 ( .A(n1833), .B(n1832), .Z(n1834) );
  AND U2216 ( .A(n1835), .B(n1834), .Z(n1838) );
  NAND U2217 ( .A(b[0]), .B(a[340]), .Z(n1836) );
  XNOR U2218 ( .A(sreg[1363]), .B(n1836), .Z(n1837) );
  XNOR U2219 ( .A(n1838), .B(n1837), .Z(c[1363]) );
  NAND U2220 ( .A(b[0]), .B(a[341]), .Z(n1841) );
  XNOR U2221 ( .A(sreg[1364]), .B(n1841), .Z(n1843) );
  NANDN U2222 ( .A(sreg[1363]), .B(n1836), .Z(n1840) );
  NAND U2223 ( .A(n1838), .B(n1837), .Z(n1839) );
  NAND U2224 ( .A(n1840), .B(n1839), .Z(n1842) );
  XNOR U2225 ( .A(n1843), .B(n1842), .Z(c[1364]) );
  NAND U2226 ( .A(b[0]), .B(a[342]), .Z(n1846) );
  XNOR U2227 ( .A(sreg[1365]), .B(n1846), .Z(n1848) );
  NANDN U2228 ( .A(sreg[1364]), .B(n1841), .Z(n1845) );
  NAND U2229 ( .A(n1843), .B(n1842), .Z(n1844) );
  AND U2230 ( .A(n1845), .B(n1844), .Z(n1847) );
  XOR U2231 ( .A(n1848), .B(n1847), .Z(c[1365]) );
  NAND U2232 ( .A(b[0]), .B(a[343]), .Z(n1851) );
  XNOR U2233 ( .A(sreg[1366]), .B(n1851), .Z(n1853) );
  NANDN U2234 ( .A(n1846), .B(sreg[1365]), .Z(n1850) );
  NAND U2235 ( .A(n1848), .B(n1847), .Z(n1849) );
  AND U2236 ( .A(n1850), .B(n1849), .Z(n1852) );
  XNOR U2237 ( .A(n1853), .B(n1852), .Z(c[1366]) );
  NAND U2238 ( .A(b[0]), .B(a[344]), .Z(n1856) );
  XNOR U2239 ( .A(sreg[1367]), .B(n1856), .Z(n1858) );
  NANDN U2240 ( .A(sreg[1366]), .B(n1851), .Z(n1855) );
  NAND U2241 ( .A(n1853), .B(n1852), .Z(n1854) );
  NAND U2242 ( .A(n1855), .B(n1854), .Z(n1857) );
  XNOR U2243 ( .A(n1858), .B(n1857), .Z(c[1367]) );
  NAND U2244 ( .A(b[0]), .B(a[345]), .Z(n1861) );
  XNOR U2245 ( .A(sreg[1368]), .B(n1861), .Z(n1863) );
  NANDN U2246 ( .A(sreg[1367]), .B(n1856), .Z(n1860) );
  NAND U2247 ( .A(n1858), .B(n1857), .Z(n1859) );
  AND U2248 ( .A(n1860), .B(n1859), .Z(n1862) );
  XOR U2249 ( .A(n1863), .B(n1862), .Z(c[1368]) );
  NAND U2250 ( .A(b[0]), .B(a[346]), .Z(n1866) );
  XNOR U2251 ( .A(sreg[1369]), .B(n1866), .Z(n1868) );
  NANDN U2252 ( .A(n1861), .B(sreg[1368]), .Z(n1865) );
  NAND U2253 ( .A(n1863), .B(n1862), .Z(n1864) );
  NAND U2254 ( .A(n1865), .B(n1864), .Z(n1867) );
  XOR U2255 ( .A(n1868), .B(n1867), .Z(c[1369]) );
  NAND U2256 ( .A(b[0]), .B(a[347]), .Z(n1871) );
  XNOR U2257 ( .A(sreg[1370]), .B(n1871), .Z(n1873) );
  NANDN U2258 ( .A(n1866), .B(sreg[1369]), .Z(n1870) );
  NAND U2259 ( .A(n1868), .B(n1867), .Z(n1869) );
  NAND U2260 ( .A(n1870), .B(n1869), .Z(n1872) );
  XOR U2261 ( .A(n1873), .B(n1872), .Z(c[1370]) );
  NANDN U2262 ( .A(n1871), .B(sreg[1370]), .Z(n1875) );
  NAND U2263 ( .A(n1873), .B(n1872), .Z(n1874) );
  AND U2264 ( .A(n1875), .B(n1874), .Z(n1878) );
  NAND U2265 ( .A(b[0]), .B(a[348]), .Z(n1876) );
  XNOR U2266 ( .A(sreg[1371]), .B(n1876), .Z(n1877) );
  XNOR U2267 ( .A(n1878), .B(n1877), .Z(c[1371]) );
  NAND U2268 ( .A(b[0]), .B(a[349]), .Z(n1881) );
  XNOR U2269 ( .A(sreg[1372]), .B(n1881), .Z(n1883) );
  NANDN U2270 ( .A(sreg[1371]), .B(n1876), .Z(n1880) );
  NAND U2271 ( .A(n1878), .B(n1877), .Z(n1879) );
  AND U2272 ( .A(n1880), .B(n1879), .Z(n1882) );
  XOR U2273 ( .A(n1883), .B(n1882), .Z(c[1372]) );
  NAND U2274 ( .A(b[0]), .B(a[350]), .Z(n1886) );
  XNOR U2275 ( .A(sreg[1373]), .B(n1886), .Z(n1888) );
  NANDN U2276 ( .A(n1881), .B(sreg[1372]), .Z(n1885) );
  NAND U2277 ( .A(n1883), .B(n1882), .Z(n1884) );
  NAND U2278 ( .A(n1885), .B(n1884), .Z(n1887) );
  XOR U2279 ( .A(n1888), .B(n1887), .Z(c[1373]) );
  NAND U2280 ( .A(b[0]), .B(a[351]), .Z(n1891) );
  XNOR U2281 ( .A(sreg[1374]), .B(n1891), .Z(n1893) );
  NANDN U2282 ( .A(n1886), .B(sreg[1373]), .Z(n1890) );
  NAND U2283 ( .A(n1888), .B(n1887), .Z(n1889) );
  AND U2284 ( .A(n1890), .B(n1889), .Z(n1892) );
  XNOR U2285 ( .A(n1893), .B(n1892), .Z(c[1374]) );
  NANDN U2286 ( .A(sreg[1374]), .B(n1891), .Z(n1895) );
  NAND U2287 ( .A(n1893), .B(n1892), .Z(n1894) );
  AND U2288 ( .A(n1895), .B(n1894), .Z(n1898) );
  NAND U2289 ( .A(b[0]), .B(a[352]), .Z(n1896) );
  XNOR U2290 ( .A(sreg[1375]), .B(n1896), .Z(n1897) );
  XOR U2291 ( .A(n1898), .B(n1897), .Z(c[1375]) );
  NAND U2292 ( .A(b[0]), .B(a[353]), .Z(n1901) );
  XNOR U2293 ( .A(sreg[1376]), .B(n1901), .Z(n1903) );
  NANDN U2294 ( .A(n1896), .B(sreg[1375]), .Z(n1900) );
  NAND U2295 ( .A(n1898), .B(n1897), .Z(n1899) );
  NAND U2296 ( .A(n1900), .B(n1899), .Z(n1902) );
  XOR U2297 ( .A(n1903), .B(n1902), .Z(c[1376]) );
  NAND U2298 ( .A(b[0]), .B(a[354]), .Z(n1906) );
  XNOR U2299 ( .A(sreg[1377]), .B(n1906), .Z(n1908) );
  NANDN U2300 ( .A(n1901), .B(sreg[1376]), .Z(n1905) );
  NAND U2301 ( .A(n1903), .B(n1902), .Z(n1904) );
  AND U2302 ( .A(n1905), .B(n1904), .Z(n1907) );
  XNOR U2303 ( .A(n1908), .B(n1907), .Z(c[1377]) );
  NANDN U2304 ( .A(sreg[1377]), .B(n1906), .Z(n1910) );
  NAND U2305 ( .A(n1908), .B(n1907), .Z(n1909) );
  AND U2306 ( .A(n1910), .B(n1909), .Z(n1913) );
  NAND U2307 ( .A(b[0]), .B(a[355]), .Z(n1911) );
  XNOR U2308 ( .A(sreg[1378]), .B(n1911), .Z(n1912) );
  XOR U2309 ( .A(n1913), .B(n1912), .Z(c[1378]) );
  NAND U2310 ( .A(b[0]), .B(a[356]), .Z(n1916) );
  XNOR U2311 ( .A(sreg[1379]), .B(n1916), .Z(n1918) );
  NANDN U2312 ( .A(n1911), .B(sreg[1378]), .Z(n1915) );
  NAND U2313 ( .A(n1913), .B(n1912), .Z(n1914) );
  NAND U2314 ( .A(n1915), .B(n1914), .Z(n1917) );
  XOR U2315 ( .A(n1918), .B(n1917), .Z(c[1379]) );
  NAND U2316 ( .A(b[0]), .B(a[357]), .Z(n1921) );
  XNOR U2317 ( .A(sreg[1380]), .B(n1921), .Z(n1923) );
  NANDN U2318 ( .A(n1916), .B(sreg[1379]), .Z(n1920) );
  NAND U2319 ( .A(n1918), .B(n1917), .Z(n1919) );
  AND U2320 ( .A(n1920), .B(n1919), .Z(n1922) );
  XNOR U2321 ( .A(n1923), .B(n1922), .Z(c[1380]) );
  NANDN U2322 ( .A(sreg[1380]), .B(n1921), .Z(n1925) );
  NAND U2323 ( .A(n1923), .B(n1922), .Z(n1924) );
  AND U2324 ( .A(n1925), .B(n1924), .Z(n1928) );
  NAND U2325 ( .A(b[0]), .B(a[358]), .Z(n1926) );
  XNOR U2326 ( .A(sreg[1381]), .B(n1926), .Z(n1927) );
  XOR U2327 ( .A(n1928), .B(n1927), .Z(c[1381]) );
  NAND U2328 ( .A(b[0]), .B(a[359]), .Z(n1931) );
  XNOR U2329 ( .A(sreg[1382]), .B(n1931), .Z(n1933) );
  NANDN U2330 ( .A(n1926), .B(sreg[1381]), .Z(n1930) );
  NAND U2331 ( .A(n1928), .B(n1927), .Z(n1929) );
  NAND U2332 ( .A(n1930), .B(n1929), .Z(n1932) );
  XOR U2333 ( .A(n1933), .B(n1932), .Z(c[1382]) );
  NANDN U2334 ( .A(n1931), .B(sreg[1382]), .Z(n1935) );
  NAND U2335 ( .A(n1933), .B(n1932), .Z(n1934) );
  AND U2336 ( .A(n1935), .B(n1934), .Z(n1938) );
  NAND U2337 ( .A(b[0]), .B(a[360]), .Z(n1936) );
  XNOR U2338 ( .A(sreg[1383]), .B(n1936), .Z(n1937) );
  XNOR U2339 ( .A(n1938), .B(n1937), .Z(c[1383]) );
  NAND U2340 ( .A(b[0]), .B(a[361]), .Z(n1941) );
  XNOR U2341 ( .A(sreg[1384]), .B(n1941), .Z(n1943) );
  NANDN U2342 ( .A(sreg[1383]), .B(n1936), .Z(n1940) );
  NAND U2343 ( .A(n1938), .B(n1937), .Z(n1939) );
  NAND U2344 ( .A(n1940), .B(n1939), .Z(n1942) );
  XNOR U2345 ( .A(n1943), .B(n1942), .Z(c[1384]) );
  NAND U2346 ( .A(b[0]), .B(a[362]), .Z(n1946) );
  XNOR U2347 ( .A(sreg[1385]), .B(n1946), .Z(n1948) );
  NANDN U2348 ( .A(sreg[1384]), .B(n1941), .Z(n1945) );
  NAND U2349 ( .A(n1943), .B(n1942), .Z(n1944) );
  NAND U2350 ( .A(n1945), .B(n1944), .Z(n1947) );
  XNOR U2351 ( .A(n1948), .B(n1947), .Z(c[1385]) );
  NAND U2352 ( .A(b[0]), .B(a[363]), .Z(n1951) );
  XNOR U2353 ( .A(sreg[1386]), .B(n1951), .Z(n1953) );
  NANDN U2354 ( .A(sreg[1385]), .B(n1946), .Z(n1950) );
  NAND U2355 ( .A(n1948), .B(n1947), .Z(n1949) );
  NAND U2356 ( .A(n1950), .B(n1949), .Z(n1952) );
  XNOR U2357 ( .A(n1953), .B(n1952), .Z(c[1386]) );
  NAND U2358 ( .A(b[0]), .B(a[364]), .Z(n1956) );
  XNOR U2359 ( .A(sreg[1387]), .B(n1956), .Z(n1958) );
  NANDN U2360 ( .A(sreg[1386]), .B(n1951), .Z(n1955) );
  NAND U2361 ( .A(n1953), .B(n1952), .Z(n1954) );
  NAND U2362 ( .A(n1955), .B(n1954), .Z(n1957) );
  XNOR U2363 ( .A(n1958), .B(n1957), .Z(c[1387]) );
  NAND U2364 ( .A(b[0]), .B(a[365]), .Z(n1961) );
  XNOR U2365 ( .A(sreg[1388]), .B(n1961), .Z(n1963) );
  NANDN U2366 ( .A(sreg[1387]), .B(n1956), .Z(n1960) );
  NAND U2367 ( .A(n1958), .B(n1957), .Z(n1959) );
  NAND U2368 ( .A(n1960), .B(n1959), .Z(n1962) );
  XNOR U2369 ( .A(n1963), .B(n1962), .Z(c[1388]) );
  NAND U2370 ( .A(b[0]), .B(a[366]), .Z(n1966) );
  XNOR U2371 ( .A(sreg[1389]), .B(n1966), .Z(n1968) );
  NANDN U2372 ( .A(sreg[1388]), .B(n1961), .Z(n1965) );
  NAND U2373 ( .A(n1963), .B(n1962), .Z(n1964) );
  NAND U2374 ( .A(n1965), .B(n1964), .Z(n1967) );
  XNOR U2375 ( .A(n1968), .B(n1967), .Z(c[1389]) );
  NAND U2376 ( .A(b[0]), .B(a[367]), .Z(n1971) );
  XNOR U2377 ( .A(sreg[1390]), .B(n1971), .Z(n1973) );
  NANDN U2378 ( .A(sreg[1389]), .B(n1966), .Z(n1970) );
  NAND U2379 ( .A(n1968), .B(n1967), .Z(n1969) );
  NAND U2380 ( .A(n1970), .B(n1969), .Z(n1972) );
  XNOR U2381 ( .A(n1973), .B(n1972), .Z(c[1390]) );
  AND U2382 ( .A(b[0]), .B(a[368]), .Z(n1978) );
  NANDN U2383 ( .A(sreg[1390]), .B(n1971), .Z(n1975) );
  NAND U2384 ( .A(n1973), .B(n1972), .Z(n1974) );
  NAND U2385 ( .A(n1975), .B(n1974), .Z(n1977) );
  XOR U2386 ( .A(n1977), .B(sreg[1391]), .Z(n1976) );
  XNOR U2387 ( .A(n1978), .B(n1976), .Z(c[1391]) );
  NAND U2388 ( .A(b[0]), .B(a[369]), .Z(n1979) );
  XNOR U2389 ( .A(sreg[1392]), .B(n1979), .Z(n1981) );
  XOR U2390 ( .A(n1981), .B(n1980), .Z(c[1392]) );
  NAND U2391 ( .A(b[0]), .B(a[370]), .Z(n1984) );
  XNOR U2392 ( .A(sreg[1393]), .B(n1984), .Z(n1986) );
  NANDN U2393 ( .A(n1979), .B(sreg[1392]), .Z(n1983) );
  NAND U2394 ( .A(n1981), .B(n1980), .Z(n1982) );
  NAND U2395 ( .A(n1983), .B(n1982), .Z(n1985) );
  XOR U2396 ( .A(n1986), .B(n1985), .Z(c[1393]) );
  NAND U2397 ( .A(b[0]), .B(a[371]), .Z(n1989) );
  XNOR U2398 ( .A(sreg[1394]), .B(n1989), .Z(n1991) );
  NANDN U2399 ( .A(n1984), .B(sreg[1393]), .Z(n1988) );
  NAND U2400 ( .A(n1986), .B(n1985), .Z(n1987) );
  AND U2401 ( .A(n1988), .B(n1987), .Z(n1990) );
  XNOR U2402 ( .A(n1991), .B(n1990), .Z(c[1394]) );
  NANDN U2403 ( .A(sreg[1394]), .B(n1989), .Z(n1993) );
  NAND U2404 ( .A(n1991), .B(n1990), .Z(n1992) );
  AND U2405 ( .A(n1993), .B(n1992), .Z(n1996) );
  NAND U2406 ( .A(b[0]), .B(a[372]), .Z(n1994) );
  XNOR U2407 ( .A(sreg[1395]), .B(n1994), .Z(n1995) );
  XOR U2408 ( .A(n1996), .B(n1995), .Z(c[1395]) );
  NAND U2409 ( .A(b[0]), .B(a[373]), .Z(n1999) );
  XNOR U2410 ( .A(sreg[1396]), .B(n1999), .Z(n2001) );
  NANDN U2411 ( .A(n1994), .B(sreg[1395]), .Z(n1998) );
  NAND U2412 ( .A(n1996), .B(n1995), .Z(n1997) );
  NAND U2413 ( .A(n1998), .B(n1997), .Z(n2000) );
  XOR U2414 ( .A(n2001), .B(n2000), .Z(c[1396]) );
  NAND U2415 ( .A(b[0]), .B(a[374]), .Z(n2004) );
  XNOR U2416 ( .A(sreg[1397]), .B(n2004), .Z(n2006) );
  NANDN U2417 ( .A(n1999), .B(sreg[1396]), .Z(n2003) );
  NAND U2418 ( .A(n2001), .B(n2000), .Z(n2002) );
  AND U2419 ( .A(n2003), .B(n2002), .Z(n2005) );
  XNOR U2420 ( .A(n2006), .B(n2005), .Z(c[1397]) );
  NAND U2421 ( .A(b[0]), .B(a[375]), .Z(n2009) );
  XNOR U2422 ( .A(sreg[1398]), .B(n2009), .Z(n2011) );
  NANDN U2423 ( .A(sreg[1397]), .B(n2004), .Z(n2008) );
  NAND U2424 ( .A(n2006), .B(n2005), .Z(n2007) );
  NAND U2425 ( .A(n2008), .B(n2007), .Z(n2010) );
  XNOR U2426 ( .A(n2011), .B(n2010), .Z(c[1398]) );
  NAND U2427 ( .A(b[0]), .B(a[376]), .Z(n2014) );
  XNOR U2428 ( .A(sreg[1399]), .B(n2014), .Z(n2016) );
  NANDN U2429 ( .A(sreg[1398]), .B(n2009), .Z(n2013) );
  NAND U2430 ( .A(n2011), .B(n2010), .Z(n2012) );
  AND U2431 ( .A(n2013), .B(n2012), .Z(n2015) );
  XOR U2432 ( .A(n2016), .B(n2015), .Z(c[1399]) );
  NANDN U2433 ( .A(n2014), .B(sreg[1399]), .Z(n2018) );
  NAND U2434 ( .A(n2016), .B(n2015), .Z(n2017) );
  AND U2435 ( .A(n2018), .B(n2017), .Z(n2021) );
  NAND U2436 ( .A(b[0]), .B(a[377]), .Z(n2019) );
  XNOR U2437 ( .A(sreg[1400]), .B(n2019), .Z(n2020) );
  XNOR U2438 ( .A(n2021), .B(n2020), .Z(c[1400]) );
  NAND U2439 ( .A(b[0]), .B(a[378]), .Z(n2024) );
  XNOR U2440 ( .A(sreg[1401]), .B(n2024), .Z(n2026) );
  NANDN U2441 ( .A(sreg[1400]), .B(n2019), .Z(n2023) );
  NAND U2442 ( .A(n2021), .B(n2020), .Z(n2022) );
  NAND U2443 ( .A(n2023), .B(n2022), .Z(n2025) );
  XNOR U2444 ( .A(n2026), .B(n2025), .Z(c[1401]) );
  NAND U2445 ( .A(b[0]), .B(a[379]), .Z(n2029) );
  XNOR U2446 ( .A(sreg[1402]), .B(n2029), .Z(n2031) );
  NANDN U2447 ( .A(sreg[1401]), .B(n2024), .Z(n2028) );
  NAND U2448 ( .A(n2026), .B(n2025), .Z(n2027) );
  NAND U2449 ( .A(n2028), .B(n2027), .Z(n2030) );
  XNOR U2450 ( .A(n2031), .B(n2030), .Z(c[1402]) );
  NAND U2451 ( .A(b[0]), .B(a[380]), .Z(n2034) );
  XNOR U2452 ( .A(sreg[1403]), .B(n2034), .Z(n2036) );
  NANDN U2453 ( .A(sreg[1402]), .B(n2029), .Z(n2033) );
  NAND U2454 ( .A(n2031), .B(n2030), .Z(n2032) );
  NAND U2455 ( .A(n2033), .B(n2032), .Z(n2035) );
  XNOR U2456 ( .A(n2036), .B(n2035), .Z(c[1403]) );
  NAND U2457 ( .A(b[0]), .B(a[381]), .Z(n2039) );
  XNOR U2458 ( .A(sreg[1404]), .B(n2039), .Z(n2041) );
  NANDN U2459 ( .A(sreg[1403]), .B(n2034), .Z(n2038) );
  NAND U2460 ( .A(n2036), .B(n2035), .Z(n2037) );
  NAND U2461 ( .A(n2038), .B(n2037), .Z(n2040) );
  XNOR U2462 ( .A(n2041), .B(n2040), .Z(c[1404]) );
  NAND U2463 ( .A(b[0]), .B(a[382]), .Z(n2044) );
  XNOR U2464 ( .A(sreg[1405]), .B(n2044), .Z(n2046) );
  NANDN U2465 ( .A(sreg[1404]), .B(n2039), .Z(n2043) );
  NAND U2466 ( .A(n2041), .B(n2040), .Z(n2042) );
  NAND U2467 ( .A(n2043), .B(n2042), .Z(n2045) );
  XNOR U2468 ( .A(n2046), .B(n2045), .Z(c[1405]) );
  NAND U2469 ( .A(b[0]), .B(a[383]), .Z(n2049) );
  XNOR U2470 ( .A(sreg[1406]), .B(n2049), .Z(n2051) );
  NANDN U2471 ( .A(sreg[1405]), .B(n2044), .Z(n2048) );
  NAND U2472 ( .A(n2046), .B(n2045), .Z(n2047) );
  NAND U2473 ( .A(n2048), .B(n2047), .Z(n2050) );
  XNOR U2474 ( .A(n2051), .B(n2050), .Z(c[1406]) );
  NAND U2475 ( .A(b[0]), .B(a[384]), .Z(n2054) );
  XNOR U2476 ( .A(sreg[1407]), .B(n2054), .Z(n2056) );
  NANDN U2477 ( .A(sreg[1406]), .B(n2049), .Z(n2053) );
  NAND U2478 ( .A(n2051), .B(n2050), .Z(n2052) );
  NAND U2479 ( .A(n2053), .B(n2052), .Z(n2055) );
  XNOR U2480 ( .A(n2056), .B(n2055), .Z(c[1407]) );
  NAND U2481 ( .A(b[0]), .B(a[385]), .Z(n2059) );
  XNOR U2482 ( .A(sreg[1408]), .B(n2059), .Z(n2061) );
  NANDN U2483 ( .A(sreg[1407]), .B(n2054), .Z(n2058) );
  NAND U2484 ( .A(n2056), .B(n2055), .Z(n2057) );
  NAND U2485 ( .A(n2058), .B(n2057), .Z(n2060) );
  XNOR U2486 ( .A(n2061), .B(n2060), .Z(c[1408]) );
  NAND U2487 ( .A(b[0]), .B(a[386]), .Z(n2064) );
  XNOR U2488 ( .A(sreg[1409]), .B(n2064), .Z(n2066) );
  NANDN U2489 ( .A(sreg[1408]), .B(n2059), .Z(n2063) );
  NAND U2490 ( .A(n2061), .B(n2060), .Z(n2062) );
  NAND U2491 ( .A(n2063), .B(n2062), .Z(n2065) );
  XNOR U2492 ( .A(n2066), .B(n2065), .Z(c[1409]) );
  NAND U2493 ( .A(b[0]), .B(a[387]), .Z(n2069) );
  XNOR U2494 ( .A(sreg[1410]), .B(n2069), .Z(n2071) );
  NANDN U2495 ( .A(sreg[1409]), .B(n2064), .Z(n2068) );
  NAND U2496 ( .A(n2066), .B(n2065), .Z(n2067) );
  NAND U2497 ( .A(n2068), .B(n2067), .Z(n2070) );
  XNOR U2498 ( .A(n2071), .B(n2070), .Z(c[1410]) );
  NAND U2499 ( .A(b[0]), .B(a[388]), .Z(n2074) );
  XNOR U2500 ( .A(sreg[1411]), .B(n2074), .Z(n2076) );
  NANDN U2501 ( .A(sreg[1410]), .B(n2069), .Z(n2073) );
  NAND U2502 ( .A(n2071), .B(n2070), .Z(n2072) );
  AND U2503 ( .A(n2073), .B(n2072), .Z(n2075) );
  XOR U2504 ( .A(n2076), .B(n2075), .Z(c[1411]) );
  NANDN U2505 ( .A(n2074), .B(sreg[1411]), .Z(n2078) );
  NAND U2506 ( .A(n2076), .B(n2075), .Z(n2077) );
  AND U2507 ( .A(n2078), .B(n2077), .Z(n2081) );
  NAND U2508 ( .A(b[0]), .B(a[389]), .Z(n2079) );
  XNOR U2509 ( .A(sreg[1412]), .B(n2079), .Z(n2080) );
  XNOR U2510 ( .A(n2081), .B(n2080), .Z(c[1412]) );
  NAND U2511 ( .A(b[0]), .B(a[390]), .Z(n2084) );
  XNOR U2512 ( .A(sreg[1413]), .B(n2084), .Z(n2086) );
  NANDN U2513 ( .A(sreg[1412]), .B(n2079), .Z(n2083) );
  NAND U2514 ( .A(n2081), .B(n2080), .Z(n2082) );
  NAND U2515 ( .A(n2083), .B(n2082), .Z(n2085) );
  XNOR U2516 ( .A(n2086), .B(n2085), .Z(c[1413]) );
  NAND U2517 ( .A(b[0]), .B(a[391]), .Z(n2089) );
  XNOR U2518 ( .A(sreg[1414]), .B(n2089), .Z(n2091) );
  NANDN U2519 ( .A(sreg[1413]), .B(n2084), .Z(n2088) );
  NAND U2520 ( .A(n2086), .B(n2085), .Z(n2087) );
  NAND U2521 ( .A(n2088), .B(n2087), .Z(n2090) );
  XNOR U2522 ( .A(n2091), .B(n2090), .Z(c[1414]) );
  NAND U2523 ( .A(b[0]), .B(a[392]), .Z(n2094) );
  XNOR U2524 ( .A(sreg[1415]), .B(n2094), .Z(n2096) );
  NANDN U2525 ( .A(sreg[1414]), .B(n2089), .Z(n2093) );
  NAND U2526 ( .A(n2091), .B(n2090), .Z(n2092) );
  NAND U2527 ( .A(n2093), .B(n2092), .Z(n2095) );
  XNOR U2528 ( .A(n2096), .B(n2095), .Z(c[1415]) );
  NAND U2529 ( .A(b[0]), .B(a[393]), .Z(n2099) );
  XNOR U2530 ( .A(sreg[1416]), .B(n2099), .Z(n2101) );
  NANDN U2531 ( .A(sreg[1415]), .B(n2094), .Z(n2098) );
  NAND U2532 ( .A(n2096), .B(n2095), .Z(n2097) );
  NAND U2533 ( .A(n2098), .B(n2097), .Z(n2100) );
  XNOR U2534 ( .A(n2101), .B(n2100), .Z(c[1416]) );
  NAND U2535 ( .A(b[0]), .B(a[394]), .Z(n2104) );
  XNOR U2536 ( .A(sreg[1417]), .B(n2104), .Z(n2106) );
  NANDN U2537 ( .A(sreg[1416]), .B(n2099), .Z(n2103) );
  NAND U2538 ( .A(n2101), .B(n2100), .Z(n2102) );
  NAND U2539 ( .A(n2103), .B(n2102), .Z(n2105) );
  XNOR U2540 ( .A(n2106), .B(n2105), .Z(c[1417]) );
  NAND U2541 ( .A(b[0]), .B(a[395]), .Z(n2109) );
  XNOR U2542 ( .A(sreg[1418]), .B(n2109), .Z(n2111) );
  NANDN U2543 ( .A(sreg[1417]), .B(n2104), .Z(n2108) );
  NAND U2544 ( .A(n2106), .B(n2105), .Z(n2107) );
  NAND U2545 ( .A(n2108), .B(n2107), .Z(n2110) );
  XNOR U2546 ( .A(n2111), .B(n2110), .Z(c[1418]) );
  NANDN U2547 ( .A(sreg[1418]), .B(n2109), .Z(n2113) );
  NAND U2548 ( .A(n2111), .B(n2110), .Z(n2112) );
  AND U2549 ( .A(n2113), .B(n2112), .Z(n2116) );
  NAND U2550 ( .A(b[0]), .B(a[396]), .Z(n2114) );
  XNOR U2551 ( .A(sreg[1419]), .B(n2114), .Z(n2115) );
  XOR U2552 ( .A(n2116), .B(n2115), .Z(c[1419]) );
  NAND U2553 ( .A(b[0]), .B(a[397]), .Z(n2119) );
  XNOR U2554 ( .A(sreg[1420]), .B(n2119), .Z(n2121) );
  NANDN U2555 ( .A(n2114), .B(sreg[1419]), .Z(n2118) );
  NAND U2556 ( .A(n2116), .B(n2115), .Z(n2117) );
  NAND U2557 ( .A(n2118), .B(n2117), .Z(n2120) );
  XOR U2558 ( .A(n2121), .B(n2120), .Z(c[1420]) );
  NANDN U2559 ( .A(n2119), .B(sreg[1420]), .Z(n2123) );
  NAND U2560 ( .A(n2121), .B(n2120), .Z(n2122) );
  AND U2561 ( .A(n2123), .B(n2122), .Z(n2125) );
  AND U2562 ( .A(b[0]), .B(a[398]), .Z(n2126) );
  XNOR U2563 ( .A(sreg[1421]), .B(n2126), .Z(n2124) );
  XOR U2564 ( .A(n2125), .B(n2124), .Z(c[1421]) );
  NAND U2565 ( .A(b[0]), .B(a[399]), .Z(n2127) );
  XNOR U2566 ( .A(sreg[1422]), .B(n2127), .Z(n2129) );
  XOR U2567 ( .A(n2129), .B(n2128), .Z(c[1422]) );
  NAND U2568 ( .A(b[0]), .B(a[400]), .Z(n2134) );
  NANDN U2569 ( .A(n2127), .B(sreg[1422]), .Z(n2131) );
  NAND U2570 ( .A(n2129), .B(n2128), .Z(n2130) );
  NAND U2571 ( .A(n2131), .B(n2130), .Z(n2133) );
  XOR U2572 ( .A(n2133), .B(sreg[1423]), .Z(n2132) );
  XNOR U2573 ( .A(n2134), .B(n2132), .Z(c[1423]) );
  NAND U2574 ( .A(b[0]), .B(a[401]), .Z(n2135) );
  XNOR U2575 ( .A(sreg[1424]), .B(n2135), .Z(n2136) );
  XNOR U2576 ( .A(n2137), .B(n2136), .Z(c[1424]) );
  NAND U2577 ( .A(b[0]), .B(a[402]), .Z(n2140) );
  XNOR U2578 ( .A(sreg[1425]), .B(n2140), .Z(n2142) );
  NANDN U2579 ( .A(n2135), .B(sreg[1424]), .Z(n2139) );
  NANDN U2580 ( .A(n2137), .B(n2136), .Z(n2138) );
  NAND U2581 ( .A(n2139), .B(n2138), .Z(n2141) );
  XOR U2582 ( .A(n2142), .B(n2141), .Z(c[1425]) );
  NANDN U2583 ( .A(n2140), .B(sreg[1425]), .Z(n2144) );
  NAND U2584 ( .A(n2142), .B(n2141), .Z(n2143) );
  AND U2585 ( .A(n2144), .B(n2143), .Z(n2147) );
  NAND U2586 ( .A(b[0]), .B(a[403]), .Z(n2145) );
  XNOR U2587 ( .A(sreg[1426]), .B(n2145), .Z(n2146) );
  XNOR U2588 ( .A(n2147), .B(n2146), .Z(c[1426]) );
  NAND U2589 ( .A(b[0]), .B(a[404]), .Z(n2150) );
  XNOR U2590 ( .A(sreg[1427]), .B(n2150), .Z(n2152) );
  NANDN U2591 ( .A(sreg[1426]), .B(n2145), .Z(n2149) );
  NAND U2592 ( .A(n2147), .B(n2146), .Z(n2148) );
  AND U2593 ( .A(n2149), .B(n2148), .Z(n2151) );
  XOR U2594 ( .A(n2152), .B(n2151), .Z(c[1427]) );
  NANDN U2595 ( .A(n2150), .B(sreg[1427]), .Z(n2154) );
  NAND U2596 ( .A(n2152), .B(n2151), .Z(n2153) );
  AND U2597 ( .A(n2154), .B(n2153), .Z(n2157) );
  NAND U2598 ( .A(b[0]), .B(a[405]), .Z(n2155) );
  XNOR U2599 ( .A(sreg[1428]), .B(n2155), .Z(n2156) );
  XNOR U2600 ( .A(n2157), .B(n2156), .Z(c[1428]) );
  NAND U2601 ( .A(b[0]), .B(a[406]), .Z(n2160) );
  XNOR U2602 ( .A(sreg[1429]), .B(n2160), .Z(n2162) );
  NANDN U2603 ( .A(sreg[1428]), .B(n2155), .Z(n2159) );
  NAND U2604 ( .A(n2157), .B(n2156), .Z(n2158) );
  NAND U2605 ( .A(n2159), .B(n2158), .Z(n2161) );
  XNOR U2606 ( .A(n2162), .B(n2161), .Z(c[1429]) );
  NAND U2607 ( .A(b[0]), .B(a[407]), .Z(n2165) );
  XNOR U2608 ( .A(sreg[1430]), .B(n2165), .Z(n2167) );
  NANDN U2609 ( .A(sreg[1429]), .B(n2160), .Z(n2164) );
  NAND U2610 ( .A(n2162), .B(n2161), .Z(n2163) );
  AND U2611 ( .A(n2164), .B(n2163), .Z(n2166) );
  XOR U2612 ( .A(n2167), .B(n2166), .Z(c[1430]) );
  NANDN U2613 ( .A(n2165), .B(sreg[1430]), .Z(n2169) );
  NAND U2614 ( .A(n2167), .B(n2166), .Z(n2168) );
  AND U2615 ( .A(n2169), .B(n2168), .Z(n2172) );
  NAND U2616 ( .A(b[0]), .B(a[408]), .Z(n2170) );
  XNOR U2617 ( .A(sreg[1431]), .B(n2170), .Z(n2171) );
  XNOR U2618 ( .A(n2172), .B(n2171), .Z(c[1431]) );
  NAND U2619 ( .A(b[0]), .B(a[409]), .Z(n2175) );
  XNOR U2620 ( .A(sreg[1432]), .B(n2175), .Z(n2177) );
  NANDN U2621 ( .A(sreg[1431]), .B(n2170), .Z(n2174) );
  NAND U2622 ( .A(n2172), .B(n2171), .Z(n2173) );
  NAND U2623 ( .A(n2174), .B(n2173), .Z(n2176) );
  XNOR U2624 ( .A(n2177), .B(n2176), .Z(c[1432]) );
  NAND U2625 ( .A(b[0]), .B(a[410]), .Z(n2180) );
  XNOR U2626 ( .A(sreg[1433]), .B(n2180), .Z(n2182) );
  NANDN U2627 ( .A(sreg[1432]), .B(n2175), .Z(n2179) );
  NAND U2628 ( .A(n2177), .B(n2176), .Z(n2178) );
  AND U2629 ( .A(n2179), .B(n2178), .Z(n2181) );
  XOR U2630 ( .A(n2182), .B(n2181), .Z(c[1433]) );
  NAND U2631 ( .A(b[0]), .B(a[411]), .Z(n2185) );
  XNOR U2632 ( .A(sreg[1434]), .B(n2185), .Z(n2187) );
  NANDN U2633 ( .A(n2180), .B(sreg[1433]), .Z(n2184) );
  NAND U2634 ( .A(n2182), .B(n2181), .Z(n2183) );
  NAND U2635 ( .A(n2184), .B(n2183), .Z(n2186) );
  XOR U2636 ( .A(n2187), .B(n2186), .Z(c[1434]) );
  NAND U2637 ( .A(b[0]), .B(a[412]), .Z(n2190) );
  XNOR U2638 ( .A(sreg[1435]), .B(n2190), .Z(n2192) );
  NANDN U2639 ( .A(n2185), .B(sreg[1434]), .Z(n2189) );
  NAND U2640 ( .A(n2187), .B(n2186), .Z(n2188) );
  NAND U2641 ( .A(n2189), .B(n2188), .Z(n2191) );
  XOR U2642 ( .A(n2192), .B(n2191), .Z(c[1435]) );
  NAND U2643 ( .A(b[0]), .B(a[413]), .Z(n2195) );
  XNOR U2644 ( .A(sreg[1436]), .B(n2195), .Z(n2197) );
  NANDN U2645 ( .A(n2190), .B(sreg[1435]), .Z(n2194) );
  NAND U2646 ( .A(n2192), .B(n2191), .Z(n2193) );
  NAND U2647 ( .A(n2194), .B(n2193), .Z(n2196) );
  XOR U2648 ( .A(n2197), .B(n2196), .Z(c[1436]) );
  NAND U2649 ( .A(b[0]), .B(a[414]), .Z(n2200) );
  XNOR U2650 ( .A(sreg[1437]), .B(n2200), .Z(n2202) );
  NANDN U2651 ( .A(n2195), .B(sreg[1436]), .Z(n2199) );
  NAND U2652 ( .A(n2197), .B(n2196), .Z(n2198) );
  NAND U2653 ( .A(n2199), .B(n2198), .Z(n2201) );
  XOR U2654 ( .A(n2202), .B(n2201), .Z(c[1437]) );
  NAND U2655 ( .A(b[0]), .B(a[415]), .Z(n2205) );
  XNOR U2656 ( .A(sreg[1438]), .B(n2205), .Z(n2207) );
  NANDN U2657 ( .A(n2200), .B(sreg[1437]), .Z(n2204) );
  NAND U2658 ( .A(n2202), .B(n2201), .Z(n2203) );
  NAND U2659 ( .A(n2204), .B(n2203), .Z(n2206) );
  XOR U2660 ( .A(n2207), .B(n2206), .Z(c[1438]) );
  NAND U2661 ( .A(b[0]), .B(a[416]), .Z(n2210) );
  XNOR U2662 ( .A(sreg[1439]), .B(n2210), .Z(n2212) );
  NANDN U2663 ( .A(n2205), .B(sreg[1438]), .Z(n2209) );
  NAND U2664 ( .A(n2207), .B(n2206), .Z(n2208) );
  NAND U2665 ( .A(n2209), .B(n2208), .Z(n2211) );
  XOR U2666 ( .A(n2212), .B(n2211), .Z(c[1439]) );
  NAND U2667 ( .A(b[0]), .B(a[417]), .Z(n2215) );
  XNOR U2668 ( .A(sreg[1440]), .B(n2215), .Z(n2217) );
  NANDN U2669 ( .A(n2210), .B(sreg[1439]), .Z(n2214) );
  NAND U2670 ( .A(n2212), .B(n2211), .Z(n2213) );
  NAND U2671 ( .A(n2214), .B(n2213), .Z(n2216) );
  XOR U2672 ( .A(n2217), .B(n2216), .Z(c[1440]) );
  NAND U2673 ( .A(b[0]), .B(a[418]), .Z(n2220) );
  XNOR U2674 ( .A(sreg[1441]), .B(n2220), .Z(n2222) );
  NANDN U2675 ( .A(n2215), .B(sreg[1440]), .Z(n2219) );
  NAND U2676 ( .A(n2217), .B(n2216), .Z(n2218) );
  NAND U2677 ( .A(n2219), .B(n2218), .Z(n2221) );
  XOR U2678 ( .A(n2222), .B(n2221), .Z(c[1441]) );
  NAND U2679 ( .A(b[0]), .B(a[419]), .Z(n2225) );
  XNOR U2680 ( .A(sreg[1442]), .B(n2225), .Z(n2227) );
  NANDN U2681 ( .A(n2220), .B(sreg[1441]), .Z(n2224) );
  NAND U2682 ( .A(n2222), .B(n2221), .Z(n2223) );
  NAND U2683 ( .A(n2224), .B(n2223), .Z(n2226) );
  XOR U2684 ( .A(n2227), .B(n2226), .Z(c[1442]) );
  NAND U2685 ( .A(b[0]), .B(a[420]), .Z(n2230) );
  XNOR U2686 ( .A(sreg[1443]), .B(n2230), .Z(n2232) );
  NANDN U2687 ( .A(n2225), .B(sreg[1442]), .Z(n2229) );
  NAND U2688 ( .A(n2227), .B(n2226), .Z(n2228) );
  NAND U2689 ( .A(n2229), .B(n2228), .Z(n2231) );
  XOR U2690 ( .A(n2232), .B(n2231), .Z(c[1443]) );
  NAND U2691 ( .A(b[0]), .B(a[421]), .Z(n2235) );
  XNOR U2692 ( .A(sreg[1444]), .B(n2235), .Z(n2237) );
  NANDN U2693 ( .A(n2230), .B(sreg[1443]), .Z(n2234) );
  NAND U2694 ( .A(n2232), .B(n2231), .Z(n2233) );
  NAND U2695 ( .A(n2234), .B(n2233), .Z(n2236) );
  XOR U2696 ( .A(n2237), .B(n2236), .Z(c[1444]) );
  NAND U2697 ( .A(b[0]), .B(a[422]), .Z(n2240) );
  XNOR U2698 ( .A(sreg[1445]), .B(n2240), .Z(n2242) );
  NANDN U2699 ( .A(n2235), .B(sreg[1444]), .Z(n2239) );
  NAND U2700 ( .A(n2237), .B(n2236), .Z(n2238) );
  NAND U2701 ( .A(n2239), .B(n2238), .Z(n2241) );
  XOR U2702 ( .A(n2242), .B(n2241), .Z(c[1445]) );
  NAND U2703 ( .A(b[0]), .B(a[423]), .Z(n2245) );
  XNOR U2704 ( .A(sreg[1446]), .B(n2245), .Z(n2247) );
  NANDN U2705 ( .A(n2240), .B(sreg[1445]), .Z(n2244) );
  NAND U2706 ( .A(n2242), .B(n2241), .Z(n2243) );
  NAND U2707 ( .A(n2244), .B(n2243), .Z(n2246) );
  XOR U2708 ( .A(n2247), .B(n2246), .Z(c[1446]) );
  NAND U2709 ( .A(b[0]), .B(a[424]), .Z(n2250) );
  XNOR U2710 ( .A(sreg[1447]), .B(n2250), .Z(n2252) );
  NANDN U2711 ( .A(n2245), .B(sreg[1446]), .Z(n2249) );
  NAND U2712 ( .A(n2247), .B(n2246), .Z(n2248) );
  NAND U2713 ( .A(n2249), .B(n2248), .Z(n2251) );
  XOR U2714 ( .A(n2252), .B(n2251), .Z(c[1447]) );
  NAND U2715 ( .A(b[0]), .B(a[425]), .Z(n2255) );
  XNOR U2716 ( .A(sreg[1448]), .B(n2255), .Z(n2257) );
  NANDN U2717 ( .A(n2250), .B(sreg[1447]), .Z(n2254) );
  NAND U2718 ( .A(n2252), .B(n2251), .Z(n2253) );
  NAND U2719 ( .A(n2254), .B(n2253), .Z(n2256) );
  XOR U2720 ( .A(n2257), .B(n2256), .Z(c[1448]) );
  NAND U2721 ( .A(b[0]), .B(a[426]), .Z(n2260) );
  XNOR U2722 ( .A(sreg[1449]), .B(n2260), .Z(n2262) );
  NANDN U2723 ( .A(n2255), .B(sreg[1448]), .Z(n2259) );
  NAND U2724 ( .A(n2257), .B(n2256), .Z(n2258) );
  NAND U2725 ( .A(n2259), .B(n2258), .Z(n2261) );
  XOR U2726 ( .A(n2262), .B(n2261), .Z(c[1449]) );
  NANDN U2727 ( .A(n2260), .B(sreg[1449]), .Z(n2264) );
  NAND U2728 ( .A(n2262), .B(n2261), .Z(n2263) );
  AND U2729 ( .A(n2264), .B(n2263), .Z(n2267) );
  NAND U2730 ( .A(b[0]), .B(a[427]), .Z(n2265) );
  XNOR U2731 ( .A(sreg[1450]), .B(n2265), .Z(n2266) );
  XNOR U2732 ( .A(n2267), .B(n2266), .Z(c[1450]) );
  NANDN U2733 ( .A(sreg[1450]), .B(n2265), .Z(n2269) );
  NAND U2734 ( .A(n2267), .B(n2266), .Z(n2268) );
  AND U2735 ( .A(n2269), .B(n2268), .Z(n2272) );
  NAND U2736 ( .A(b[0]), .B(a[428]), .Z(n2270) );
  XNOR U2737 ( .A(sreg[1451]), .B(n2270), .Z(n2271) );
  XOR U2738 ( .A(n2272), .B(n2271), .Z(c[1451]) );
  NAND U2739 ( .A(b[0]), .B(a[429]), .Z(n2275) );
  XNOR U2740 ( .A(sreg[1452]), .B(n2275), .Z(n2277) );
  NANDN U2741 ( .A(n2270), .B(sreg[1451]), .Z(n2274) );
  NAND U2742 ( .A(n2272), .B(n2271), .Z(n2273) );
  NAND U2743 ( .A(n2274), .B(n2273), .Z(n2276) );
  XOR U2744 ( .A(n2277), .B(n2276), .Z(c[1452]) );
  NANDN U2745 ( .A(n2275), .B(sreg[1452]), .Z(n2279) );
  NAND U2746 ( .A(n2277), .B(n2276), .Z(n2278) );
  AND U2747 ( .A(n2279), .B(n2278), .Z(n2282) );
  NAND U2748 ( .A(b[0]), .B(a[430]), .Z(n2280) );
  XNOR U2749 ( .A(sreg[1453]), .B(n2280), .Z(n2281) );
  XNOR U2750 ( .A(n2282), .B(n2281), .Z(c[1453]) );
  NAND U2751 ( .A(b[0]), .B(a[431]), .Z(n2285) );
  XNOR U2752 ( .A(sreg[1454]), .B(n2285), .Z(n2287) );
  NANDN U2753 ( .A(sreg[1453]), .B(n2280), .Z(n2284) );
  NAND U2754 ( .A(n2282), .B(n2281), .Z(n2283) );
  AND U2755 ( .A(n2284), .B(n2283), .Z(n2286) );
  XOR U2756 ( .A(n2287), .B(n2286), .Z(c[1454]) );
  NANDN U2757 ( .A(n2285), .B(sreg[1454]), .Z(n2289) );
  NAND U2758 ( .A(n2287), .B(n2286), .Z(n2288) );
  AND U2759 ( .A(n2289), .B(n2288), .Z(n2291) );
  AND U2760 ( .A(b[0]), .B(a[432]), .Z(n2292) );
  XNOR U2761 ( .A(sreg[1455]), .B(n2292), .Z(n2290) );
  XOR U2762 ( .A(n2291), .B(n2290), .Z(c[1455]) );
  NAND U2763 ( .A(b[0]), .B(a[433]), .Z(n2293) );
  XNOR U2764 ( .A(sreg[1456]), .B(n2293), .Z(n2295) );
  XOR U2765 ( .A(n2295), .B(n2294), .Z(c[1456]) );
  NAND U2766 ( .A(b[0]), .B(a[434]), .Z(n2298) );
  XNOR U2767 ( .A(sreg[1457]), .B(n2298), .Z(n2300) );
  NANDN U2768 ( .A(n2293), .B(sreg[1456]), .Z(n2297) );
  NAND U2769 ( .A(n2295), .B(n2294), .Z(n2296) );
  NAND U2770 ( .A(n2297), .B(n2296), .Z(n2299) );
  XOR U2771 ( .A(n2300), .B(n2299), .Z(c[1457]) );
  NAND U2772 ( .A(b[0]), .B(a[435]), .Z(n2303) );
  XNOR U2773 ( .A(sreg[1458]), .B(n2303), .Z(n2305) );
  NANDN U2774 ( .A(n2298), .B(sreg[1457]), .Z(n2302) );
  NAND U2775 ( .A(n2300), .B(n2299), .Z(n2301) );
  AND U2776 ( .A(n2302), .B(n2301), .Z(n2304) );
  XNOR U2777 ( .A(n2305), .B(n2304), .Z(c[1458]) );
  NANDN U2778 ( .A(sreg[1458]), .B(n2303), .Z(n2307) );
  NAND U2779 ( .A(n2305), .B(n2304), .Z(n2306) );
  AND U2780 ( .A(n2307), .B(n2306), .Z(n2310) );
  NAND U2781 ( .A(b[0]), .B(a[436]), .Z(n2308) );
  XNOR U2782 ( .A(sreg[1459]), .B(n2308), .Z(n2309) );
  XOR U2783 ( .A(n2310), .B(n2309), .Z(c[1459]) );
  NAND U2784 ( .A(b[0]), .B(a[437]), .Z(n2313) );
  XNOR U2785 ( .A(sreg[1460]), .B(n2313), .Z(n2315) );
  NANDN U2786 ( .A(n2308), .B(sreg[1459]), .Z(n2312) );
  NAND U2787 ( .A(n2310), .B(n2309), .Z(n2311) );
  NAND U2788 ( .A(n2312), .B(n2311), .Z(n2314) );
  XOR U2789 ( .A(n2315), .B(n2314), .Z(c[1460]) );
  NAND U2790 ( .A(b[0]), .B(a[438]), .Z(n2318) );
  XNOR U2791 ( .A(sreg[1461]), .B(n2318), .Z(n2320) );
  NANDN U2792 ( .A(n2313), .B(sreg[1460]), .Z(n2317) );
  NAND U2793 ( .A(n2315), .B(n2314), .Z(n2316) );
  NAND U2794 ( .A(n2317), .B(n2316), .Z(n2319) );
  XOR U2795 ( .A(n2320), .B(n2319), .Z(c[1461]) );
  NAND U2796 ( .A(b[0]), .B(a[439]), .Z(n2323) );
  XNOR U2797 ( .A(sreg[1462]), .B(n2323), .Z(n2325) );
  NANDN U2798 ( .A(n2318), .B(sreg[1461]), .Z(n2322) );
  NAND U2799 ( .A(n2320), .B(n2319), .Z(n2321) );
  NAND U2800 ( .A(n2322), .B(n2321), .Z(n2324) );
  XOR U2801 ( .A(n2325), .B(n2324), .Z(c[1462]) );
  NAND U2802 ( .A(b[0]), .B(a[440]), .Z(n2328) );
  XNOR U2803 ( .A(sreg[1463]), .B(n2328), .Z(n2330) );
  NANDN U2804 ( .A(n2323), .B(sreg[1462]), .Z(n2327) );
  NAND U2805 ( .A(n2325), .B(n2324), .Z(n2326) );
  NAND U2806 ( .A(n2327), .B(n2326), .Z(n2329) );
  XOR U2807 ( .A(n2330), .B(n2329), .Z(c[1463]) );
  NAND U2808 ( .A(b[0]), .B(a[441]), .Z(n2333) );
  XNOR U2809 ( .A(sreg[1464]), .B(n2333), .Z(n2335) );
  NANDN U2810 ( .A(n2328), .B(sreg[1463]), .Z(n2332) );
  NAND U2811 ( .A(n2330), .B(n2329), .Z(n2331) );
  NAND U2812 ( .A(n2332), .B(n2331), .Z(n2334) );
  XOR U2813 ( .A(n2335), .B(n2334), .Z(c[1464]) );
  NAND U2814 ( .A(b[0]), .B(a[442]), .Z(n2338) );
  XNOR U2815 ( .A(sreg[1465]), .B(n2338), .Z(n2340) );
  NANDN U2816 ( .A(n2333), .B(sreg[1464]), .Z(n2337) );
  NAND U2817 ( .A(n2335), .B(n2334), .Z(n2336) );
  NAND U2818 ( .A(n2337), .B(n2336), .Z(n2339) );
  XOR U2819 ( .A(n2340), .B(n2339), .Z(c[1465]) );
  NAND U2820 ( .A(b[0]), .B(a[443]), .Z(n2343) );
  XNOR U2821 ( .A(sreg[1466]), .B(n2343), .Z(n2345) );
  NANDN U2822 ( .A(n2338), .B(sreg[1465]), .Z(n2342) );
  NAND U2823 ( .A(n2340), .B(n2339), .Z(n2341) );
  NAND U2824 ( .A(n2342), .B(n2341), .Z(n2344) );
  XOR U2825 ( .A(n2345), .B(n2344), .Z(c[1466]) );
  NANDN U2826 ( .A(n2343), .B(sreg[1466]), .Z(n2347) );
  NAND U2827 ( .A(n2345), .B(n2344), .Z(n2346) );
  AND U2828 ( .A(n2347), .B(n2346), .Z(n2350) );
  NAND U2829 ( .A(b[0]), .B(a[444]), .Z(n2348) );
  XNOR U2830 ( .A(sreg[1467]), .B(n2348), .Z(n2349) );
  XNOR U2831 ( .A(n2350), .B(n2349), .Z(c[1467]) );
  NANDN U2832 ( .A(sreg[1467]), .B(n2348), .Z(n2352) );
  NAND U2833 ( .A(n2350), .B(n2349), .Z(n2351) );
  AND U2834 ( .A(n2352), .B(n2351), .Z(n2355) );
  NAND U2835 ( .A(b[0]), .B(a[445]), .Z(n2353) );
  XNOR U2836 ( .A(sreg[1468]), .B(n2353), .Z(n2354) );
  XOR U2837 ( .A(n2355), .B(n2354), .Z(c[1468]) );
  NANDN U2838 ( .A(n2353), .B(sreg[1468]), .Z(n2357) );
  NAND U2839 ( .A(n2355), .B(n2354), .Z(n2356) );
  AND U2840 ( .A(n2357), .B(n2356), .Z(n2360) );
  NAND U2841 ( .A(b[0]), .B(a[446]), .Z(n2358) );
  XNOR U2842 ( .A(sreg[1469]), .B(n2358), .Z(n2359) );
  XNOR U2843 ( .A(n2360), .B(n2359), .Z(c[1469]) );
  NAND U2844 ( .A(b[0]), .B(a[447]), .Z(n2363) );
  XNOR U2845 ( .A(sreg[1470]), .B(n2363), .Z(n2365) );
  NANDN U2846 ( .A(sreg[1469]), .B(n2358), .Z(n2362) );
  NAND U2847 ( .A(n2360), .B(n2359), .Z(n2361) );
  NAND U2848 ( .A(n2362), .B(n2361), .Z(n2364) );
  XNOR U2849 ( .A(n2365), .B(n2364), .Z(c[1470]) );
  NAND U2850 ( .A(b[0]), .B(a[448]), .Z(n2368) );
  XNOR U2851 ( .A(sreg[1471]), .B(n2368), .Z(n2370) );
  NANDN U2852 ( .A(sreg[1470]), .B(n2363), .Z(n2367) );
  NAND U2853 ( .A(n2365), .B(n2364), .Z(n2366) );
  NAND U2854 ( .A(n2367), .B(n2366), .Z(n2369) );
  XNOR U2855 ( .A(n2370), .B(n2369), .Z(c[1471]) );
  NANDN U2856 ( .A(sreg[1471]), .B(n2368), .Z(n2372) );
  NAND U2857 ( .A(n2370), .B(n2369), .Z(n2371) );
  AND U2858 ( .A(n2372), .B(n2371), .Z(n2375) );
  NAND U2859 ( .A(b[0]), .B(a[449]), .Z(n2373) );
  XNOR U2860 ( .A(sreg[1472]), .B(n2373), .Z(n2374) );
  XOR U2861 ( .A(n2375), .B(n2374), .Z(c[1472]) );
  NAND U2862 ( .A(b[0]), .B(a[450]), .Z(n2378) );
  XNOR U2863 ( .A(sreg[1473]), .B(n2378), .Z(n2380) );
  NANDN U2864 ( .A(n2373), .B(sreg[1472]), .Z(n2377) );
  NAND U2865 ( .A(n2375), .B(n2374), .Z(n2376) );
  NAND U2866 ( .A(n2377), .B(n2376), .Z(n2379) );
  XOR U2867 ( .A(n2380), .B(n2379), .Z(c[1473]) );
  NAND U2868 ( .A(b[0]), .B(a[451]), .Z(n2383) );
  XNOR U2869 ( .A(sreg[1474]), .B(n2383), .Z(n2385) );
  NANDN U2870 ( .A(n2378), .B(sreg[1473]), .Z(n2382) );
  NAND U2871 ( .A(n2380), .B(n2379), .Z(n2381) );
  AND U2872 ( .A(n2382), .B(n2381), .Z(n2384) );
  XNOR U2873 ( .A(n2385), .B(n2384), .Z(c[1474]) );
  NAND U2874 ( .A(b[0]), .B(a[452]), .Z(n2388) );
  XNOR U2875 ( .A(sreg[1475]), .B(n2388), .Z(n2390) );
  NANDN U2876 ( .A(sreg[1474]), .B(n2383), .Z(n2387) );
  NAND U2877 ( .A(n2385), .B(n2384), .Z(n2386) );
  AND U2878 ( .A(n2387), .B(n2386), .Z(n2389) );
  XOR U2879 ( .A(n2390), .B(n2389), .Z(c[1475]) );
  NAND U2880 ( .A(b[0]), .B(a[453]), .Z(n2393) );
  XNOR U2881 ( .A(sreg[1476]), .B(n2393), .Z(n2395) );
  NANDN U2882 ( .A(n2388), .B(sreg[1475]), .Z(n2392) );
  NAND U2883 ( .A(n2390), .B(n2389), .Z(n2391) );
  NAND U2884 ( .A(n2392), .B(n2391), .Z(n2394) );
  XOR U2885 ( .A(n2395), .B(n2394), .Z(c[1476]) );
  NAND U2886 ( .A(b[0]), .B(a[454]), .Z(n2398) );
  XNOR U2887 ( .A(sreg[1477]), .B(n2398), .Z(n2400) );
  NANDN U2888 ( .A(n2393), .B(sreg[1476]), .Z(n2397) );
  NAND U2889 ( .A(n2395), .B(n2394), .Z(n2396) );
  AND U2890 ( .A(n2397), .B(n2396), .Z(n2399) );
  XNOR U2891 ( .A(n2400), .B(n2399), .Z(c[1477]) );
  NAND U2892 ( .A(b[0]), .B(a[455]), .Z(n2403) );
  XNOR U2893 ( .A(sreg[1478]), .B(n2403), .Z(n2405) );
  NANDN U2894 ( .A(sreg[1477]), .B(n2398), .Z(n2402) );
  NAND U2895 ( .A(n2400), .B(n2399), .Z(n2401) );
  NAND U2896 ( .A(n2402), .B(n2401), .Z(n2404) );
  XNOR U2897 ( .A(n2405), .B(n2404), .Z(c[1478]) );
  NAND U2898 ( .A(b[0]), .B(a[456]), .Z(n2408) );
  XNOR U2899 ( .A(sreg[1479]), .B(n2408), .Z(n2410) );
  NANDN U2900 ( .A(sreg[1478]), .B(n2403), .Z(n2407) );
  NAND U2901 ( .A(n2405), .B(n2404), .Z(n2406) );
  AND U2902 ( .A(n2407), .B(n2406), .Z(n2409) );
  XOR U2903 ( .A(n2410), .B(n2409), .Z(c[1479]) );
  NAND U2904 ( .A(b[0]), .B(a[457]), .Z(n2413) );
  XNOR U2905 ( .A(sreg[1480]), .B(n2413), .Z(n2415) );
  NANDN U2906 ( .A(n2408), .B(sreg[1479]), .Z(n2412) );
  NAND U2907 ( .A(n2410), .B(n2409), .Z(n2411) );
  AND U2908 ( .A(n2412), .B(n2411), .Z(n2414) );
  XNOR U2909 ( .A(n2415), .B(n2414), .Z(c[1480]) );
  NAND U2910 ( .A(b[0]), .B(a[458]), .Z(n2420) );
  NANDN U2911 ( .A(sreg[1480]), .B(n2413), .Z(n2417) );
  NAND U2912 ( .A(n2415), .B(n2414), .Z(n2416) );
  AND U2913 ( .A(n2417), .B(n2416), .Z(n2419) );
  XOR U2914 ( .A(sreg[1481]), .B(n2419), .Z(n2418) );
  XNOR U2915 ( .A(n2420), .B(n2418), .Z(c[1481]) );
  NAND U2916 ( .A(b[0]), .B(a[459]), .Z(n2421) );
  XNOR U2917 ( .A(sreg[1482]), .B(n2421), .Z(n2422) );
  XOR U2918 ( .A(n2423), .B(n2422), .Z(c[1482]) );
  NAND U2919 ( .A(b[0]), .B(a[460]), .Z(n2426) );
  XNOR U2920 ( .A(sreg[1483]), .B(n2426), .Z(n2428) );
  NANDN U2921 ( .A(n2421), .B(sreg[1482]), .Z(n2425) );
  NAND U2922 ( .A(n2423), .B(n2422), .Z(n2424) );
  NAND U2923 ( .A(n2425), .B(n2424), .Z(n2427) );
  XOR U2924 ( .A(n2428), .B(n2427), .Z(c[1483]) );
  NANDN U2925 ( .A(n2426), .B(sreg[1483]), .Z(n2430) );
  NAND U2926 ( .A(n2428), .B(n2427), .Z(n2429) );
  AND U2927 ( .A(n2430), .B(n2429), .Z(n2433) );
  NAND U2928 ( .A(b[0]), .B(a[461]), .Z(n2431) );
  XNOR U2929 ( .A(sreg[1484]), .B(n2431), .Z(n2432) );
  XNOR U2930 ( .A(n2433), .B(n2432), .Z(c[1484]) );
  NAND U2931 ( .A(b[0]), .B(a[462]), .Z(n2436) );
  XNOR U2932 ( .A(sreg[1485]), .B(n2436), .Z(n2438) );
  NANDN U2933 ( .A(sreg[1484]), .B(n2431), .Z(n2435) );
  NAND U2934 ( .A(n2433), .B(n2432), .Z(n2434) );
  AND U2935 ( .A(n2435), .B(n2434), .Z(n2437) );
  XOR U2936 ( .A(n2438), .B(n2437), .Z(c[1485]) );
  NAND U2937 ( .A(b[0]), .B(a[463]), .Z(n2441) );
  XNOR U2938 ( .A(sreg[1486]), .B(n2441), .Z(n2443) );
  NANDN U2939 ( .A(n2436), .B(sreg[1485]), .Z(n2440) );
  NAND U2940 ( .A(n2438), .B(n2437), .Z(n2439) );
  NAND U2941 ( .A(n2440), .B(n2439), .Z(n2442) );
  XOR U2942 ( .A(n2443), .B(n2442), .Z(c[1486]) );
  NAND U2943 ( .A(b[0]), .B(a[464]), .Z(n2446) );
  XNOR U2944 ( .A(sreg[1487]), .B(n2446), .Z(n2448) );
  NANDN U2945 ( .A(n2441), .B(sreg[1486]), .Z(n2445) );
  NAND U2946 ( .A(n2443), .B(n2442), .Z(n2444) );
  NAND U2947 ( .A(n2445), .B(n2444), .Z(n2447) );
  XOR U2948 ( .A(n2448), .B(n2447), .Z(c[1487]) );
  NANDN U2949 ( .A(n2446), .B(sreg[1487]), .Z(n2450) );
  NAND U2950 ( .A(n2448), .B(n2447), .Z(n2449) );
  AND U2951 ( .A(n2450), .B(n2449), .Z(n2453) );
  NAND U2952 ( .A(b[0]), .B(a[465]), .Z(n2451) );
  XNOR U2953 ( .A(sreg[1488]), .B(n2451), .Z(n2452) );
  XNOR U2954 ( .A(n2453), .B(n2452), .Z(c[1488]) );
  NAND U2955 ( .A(b[0]), .B(a[466]), .Z(n2456) );
  XNOR U2956 ( .A(sreg[1489]), .B(n2456), .Z(n2458) );
  NANDN U2957 ( .A(sreg[1488]), .B(n2451), .Z(n2455) );
  NAND U2958 ( .A(n2453), .B(n2452), .Z(n2454) );
  AND U2959 ( .A(n2455), .B(n2454), .Z(n2457) );
  XOR U2960 ( .A(n2458), .B(n2457), .Z(c[1489]) );
  NAND U2961 ( .A(b[0]), .B(a[467]), .Z(n2461) );
  XNOR U2962 ( .A(sreg[1490]), .B(n2461), .Z(n2463) );
  NANDN U2963 ( .A(n2456), .B(sreg[1489]), .Z(n2460) );
  NAND U2964 ( .A(n2458), .B(n2457), .Z(n2459) );
  NAND U2965 ( .A(n2460), .B(n2459), .Z(n2462) );
  XOR U2966 ( .A(n2463), .B(n2462), .Z(c[1490]) );
  NAND U2967 ( .A(b[0]), .B(a[468]), .Z(n2466) );
  XNOR U2968 ( .A(sreg[1491]), .B(n2466), .Z(n2468) );
  NANDN U2969 ( .A(n2461), .B(sreg[1490]), .Z(n2465) );
  NAND U2970 ( .A(n2463), .B(n2462), .Z(n2464) );
  AND U2971 ( .A(n2465), .B(n2464), .Z(n2467) );
  XNOR U2972 ( .A(n2468), .B(n2467), .Z(c[1491]) );
  NAND U2973 ( .A(b[0]), .B(a[469]), .Z(n2471) );
  XNOR U2974 ( .A(sreg[1492]), .B(n2471), .Z(n2473) );
  NANDN U2975 ( .A(sreg[1491]), .B(n2466), .Z(n2470) );
  NAND U2976 ( .A(n2468), .B(n2467), .Z(n2469) );
  NAND U2977 ( .A(n2470), .B(n2469), .Z(n2472) );
  XNOR U2978 ( .A(n2473), .B(n2472), .Z(c[1492]) );
  NAND U2979 ( .A(b[0]), .B(a[470]), .Z(n2476) );
  XNOR U2980 ( .A(sreg[1493]), .B(n2476), .Z(n2478) );
  NANDN U2981 ( .A(sreg[1492]), .B(n2471), .Z(n2475) );
  NAND U2982 ( .A(n2473), .B(n2472), .Z(n2474) );
  AND U2983 ( .A(n2475), .B(n2474), .Z(n2477) );
  XOR U2984 ( .A(n2478), .B(n2477), .Z(c[1493]) );
  NAND U2985 ( .A(b[0]), .B(a[471]), .Z(n2481) );
  XNOR U2986 ( .A(sreg[1494]), .B(n2481), .Z(n2483) );
  NANDN U2987 ( .A(n2476), .B(sreg[1493]), .Z(n2480) );
  NAND U2988 ( .A(n2478), .B(n2477), .Z(n2479) );
  AND U2989 ( .A(n2480), .B(n2479), .Z(n2482) );
  XNOR U2990 ( .A(n2483), .B(n2482), .Z(c[1494]) );
  NAND U2991 ( .A(b[0]), .B(a[472]), .Z(n2486) );
  XNOR U2992 ( .A(sreg[1495]), .B(n2486), .Z(n2488) );
  NANDN U2993 ( .A(sreg[1494]), .B(n2481), .Z(n2485) );
  NAND U2994 ( .A(n2483), .B(n2482), .Z(n2484) );
  NAND U2995 ( .A(n2485), .B(n2484), .Z(n2487) );
  XNOR U2996 ( .A(n2488), .B(n2487), .Z(c[1495]) );
  NAND U2997 ( .A(b[0]), .B(a[473]), .Z(n2491) );
  XNOR U2998 ( .A(sreg[1496]), .B(n2491), .Z(n2493) );
  NANDN U2999 ( .A(sreg[1495]), .B(n2486), .Z(n2490) );
  NAND U3000 ( .A(n2488), .B(n2487), .Z(n2489) );
  AND U3001 ( .A(n2490), .B(n2489), .Z(n2492) );
  XOR U3002 ( .A(n2493), .B(n2492), .Z(c[1496]) );
  NAND U3003 ( .A(b[0]), .B(a[474]), .Z(n2496) );
  XNOR U3004 ( .A(sreg[1497]), .B(n2496), .Z(n2498) );
  NANDN U3005 ( .A(n2491), .B(sreg[1496]), .Z(n2495) );
  NAND U3006 ( .A(n2493), .B(n2492), .Z(n2494) );
  NAND U3007 ( .A(n2495), .B(n2494), .Z(n2497) );
  XOR U3008 ( .A(n2498), .B(n2497), .Z(c[1497]) );
  NANDN U3009 ( .A(n2496), .B(sreg[1497]), .Z(n2500) );
  NAND U3010 ( .A(n2498), .B(n2497), .Z(n2499) );
  AND U3011 ( .A(n2500), .B(n2499), .Z(n2503) );
  NAND U3012 ( .A(b[0]), .B(a[475]), .Z(n2501) );
  XNOR U3013 ( .A(sreg[1498]), .B(n2501), .Z(n2502) );
  XNOR U3014 ( .A(n2503), .B(n2502), .Z(c[1498]) );
  NANDN U3015 ( .A(sreg[1498]), .B(n2501), .Z(n2505) );
  NAND U3016 ( .A(n2503), .B(n2502), .Z(n2504) );
  AND U3017 ( .A(n2505), .B(n2504), .Z(n2508) );
  NAND U3018 ( .A(b[0]), .B(a[476]), .Z(n2506) );
  XNOR U3019 ( .A(sreg[1499]), .B(n2506), .Z(n2507) );
  XOR U3020 ( .A(n2508), .B(n2507), .Z(c[1499]) );
  NAND U3021 ( .A(b[0]), .B(a[477]), .Z(n2511) );
  XNOR U3022 ( .A(sreg[1500]), .B(n2511), .Z(n2513) );
  NANDN U3023 ( .A(n2506), .B(sreg[1499]), .Z(n2510) );
  NAND U3024 ( .A(n2508), .B(n2507), .Z(n2509) );
  AND U3025 ( .A(n2510), .B(n2509), .Z(n2512) );
  XNOR U3026 ( .A(n2513), .B(n2512), .Z(c[1500]) );
  NAND U3027 ( .A(b[0]), .B(a[478]), .Z(n2516) );
  XNOR U3028 ( .A(sreg[1501]), .B(n2516), .Z(n2518) );
  NANDN U3029 ( .A(sreg[1500]), .B(n2511), .Z(n2515) );
  NAND U3030 ( .A(n2513), .B(n2512), .Z(n2514) );
  NAND U3031 ( .A(n2515), .B(n2514), .Z(n2517) );
  XNOR U3032 ( .A(n2518), .B(n2517), .Z(c[1501]) );
  NANDN U3033 ( .A(sreg[1501]), .B(n2516), .Z(n2520) );
  NAND U3034 ( .A(n2518), .B(n2517), .Z(n2519) );
  AND U3035 ( .A(n2520), .B(n2519), .Z(n2523) );
  NAND U3036 ( .A(b[0]), .B(a[479]), .Z(n2521) );
  XNOR U3037 ( .A(sreg[1502]), .B(n2521), .Z(n2522) );
  XOR U3038 ( .A(n2523), .B(n2522), .Z(c[1502]) );
  NAND U3039 ( .A(b[0]), .B(a[480]), .Z(n2526) );
  XNOR U3040 ( .A(sreg[1503]), .B(n2526), .Z(n2528) );
  NANDN U3041 ( .A(n2521), .B(sreg[1502]), .Z(n2525) );
  NAND U3042 ( .A(n2523), .B(n2522), .Z(n2524) );
  AND U3043 ( .A(n2525), .B(n2524), .Z(n2527) );
  XNOR U3044 ( .A(n2528), .B(n2527), .Z(c[1503]) );
  NAND U3045 ( .A(b[0]), .B(a[481]), .Z(n2531) );
  XNOR U3046 ( .A(sreg[1504]), .B(n2531), .Z(n2533) );
  NANDN U3047 ( .A(sreg[1503]), .B(n2526), .Z(n2530) );
  NAND U3048 ( .A(n2528), .B(n2527), .Z(n2529) );
  NAND U3049 ( .A(n2530), .B(n2529), .Z(n2532) );
  XNOR U3050 ( .A(n2533), .B(n2532), .Z(c[1504]) );
  NANDN U3051 ( .A(sreg[1504]), .B(n2531), .Z(n2535) );
  NAND U3052 ( .A(n2533), .B(n2532), .Z(n2534) );
  AND U3053 ( .A(n2535), .B(n2534), .Z(n2538) );
  NAND U3054 ( .A(b[0]), .B(a[482]), .Z(n2536) );
  XNOR U3055 ( .A(sreg[1505]), .B(n2536), .Z(n2537) );
  XOR U3056 ( .A(n2538), .B(n2537), .Z(c[1505]) );
  NAND U3057 ( .A(b[0]), .B(a[483]), .Z(n2541) );
  XNOR U3058 ( .A(sreg[1506]), .B(n2541), .Z(n2543) );
  NANDN U3059 ( .A(n2536), .B(sreg[1505]), .Z(n2540) );
  NAND U3060 ( .A(n2538), .B(n2537), .Z(n2539) );
  AND U3061 ( .A(n2540), .B(n2539), .Z(n2542) );
  XNOR U3062 ( .A(n2543), .B(n2542), .Z(c[1506]) );
  NANDN U3063 ( .A(sreg[1506]), .B(n2541), .Z(n2545) );
  NAND U3064 ( .A(n2543), .B(n2542), .Z(n2544) );
  AND U3065 ( .A(n2545), .B(n2544), .Z(n2548) );
  NAND U3066 ( .A(b[0]), .B(a[484]), .Z(n2546) );
  XNOR U3067 ( .A(sreg[1507]), .B(n2546), .Z(n2547) );
  XOR U3068 ( .A(n2548), .B(n2547), .Z(c[1507]) );
  NAND U3069 ( .A(b[0]), .B(a[485]), .Z(n2551) );
  XNOR U3070 ( .A(sreg[1508]), .B(n2551), .Z(n2553) );
  NANDN U3071 ( .A(n2546), .B(sreg[1507]), .Z(n2550) );
  NAND U3072 ( .A(n2548), .B(n2547), .Z(n2549) );
  NAND U3073 ( .A(n2550), .B(n2549), .Z(n2552) );
  XOR U3074 ( .A(n2553), .B(n2552), .Z(c[1508]) );
  NANDN U3075 ( .A(n2551), .B(sreg[1508]), .Z(n2555) );
  NAND U3076 ( .A(n2553), .B(n2552), .Z(n2554) );
  AND U3077 ( .A(n2555), .B(n2554), .Z(n2558) );
  NAND U3078 ( .A(b[0]), .B(a[486]), .Z(n2556) );
  XNOR U3079 ( .A(sreg[1509]), .B(n2556), .Z(n2557) );
  XNOR U3080 ( .A(n2558), .B(n2557), .Z(c[1509]) );
  NAND U3081 ( .A(b[0]), .B(a[487]), .Z(n2561) );
  XNOR U3082 ( .A(sreg[1510]), .B(n2561), .Z(n2563) );
  NANDN U3083 ( .A(sreg[1509]), .B(n2556), .Z(n2560) );
  NAND U3084 ( .A(n2558), .B(n2557), .Z(n2559) );
  AND U3085 ( .A(n2560), .B(n2559), .Z(n2562) );
  XOR U3086 ( .A(n2563), .B(n2562), .Z(c[1510]) );
  NANDN U3087 ( .A(n2561), .B(sreg[1510]), .Z(n2565) );
  NAND U3088 ( .A(n2563), .B(n2562), .Z(n2564) );
  AND U3089 ( .A(n2565), .B(n2564), .Z(n2567) );
  AND U3090 ( .A(b[0]), .B(a[488]), .Z(n2568) );
  XNOR U3091 ( .A(sreg[1511]), .B(n2568), .Z(n2566) );
  XOR U3092 ( .A(n2567), .B(n2566), .Z(c[1511]) );
  NAND U3093 ( .A(b[0]), .B(a[489]), .Z(n2569) );
  XNOR U3094 ( .A(sreg[1512]), .B(n2569), .Z(n2571) );
  XOR U3095 ( .A(n2571), .B(n2570), .Z(c[1512]) );
  NAND U3096 ( .A(b[0]), .B(a[490]), .Z(n2574) );
  XNOR U3097 ( .A(sreg[1513]), .B(n2574), .Z(n2576) );
  NANDN U3098 ( .A(n2569), .B(sreg[1512]), .Z(n2573) );
  NAND U3099 ( .A(n2571), .B(n2570), .Z(n2572) );
  NAND U3100 ( .A(n2573), .B(n2572), .Z(n2575) );
  XOR U3101 ( .A(n2576), .B(n2575), .Z(c[1513]) );
  NANDN U3102 ( .A(n2574), .B(sreg[1513]), .Z(n2578) );
  NAND U3103 ( .A(n2576), .B(n2575), .Z(n2577) );
  NAND U3104 ( .A(n2578), .B(n2577), .Z(n2581) );
  NAND U3105 ( .A(b[0]), .B(a[491]), .Z(n2580) );
  XOR U3106 ( .A(sreg[1514]), .B(n2580), .Z(n2579) );
  XNOR U3107 ( .A(n2581), .B(n2579), .Z(c[1514]) );
  NAND U3108 ( .A(b[0]), .B(a[492]), .Z(n2582) );
  XNOR U3109 ( .A(sreg[1515]), .B(n2582), .Z(n2583) );
  XOR U3110 ( .A(n2584), .B(n2583), .Z(c[1515]) );
  NANDN U3111 ( .A(n2582), .B(sreg[1515]), .Z(n2586) );
  NAND U3112 ( .A(n2584), .B(n2583), .Z(n2585) );
  AND U3113 ( .A(n2586), .B(n2585), .Z(n2589) );
  NAND U3114 ( .A(b[0]), .B(a[493]), .Z(n2587) );
  XNOR U3115 ( .A(sreg[1516]), .B(n2587), .Z(n2588) );
  XNOR U3116 ( .A(n2589), .B(n2588), .Z(c[1516]) );
  NAND U3117 ( .A(b[0]), .B(a[494]), .Z(n2592) );
  XNOR U3118 ( .A(sreg[1517]), .B(n2592), .Z(n2594) );
  NANDN U3119 ( .A(sreg[1516]), .B(n2587), .Z(n2591) );
  NAND U3120 ( .A(n2589), .B(n2588), .Z(n2590) );
  NAND U3121 ( .A(n2591), .B(n2590), .Z(n2593) );
  XNOR U3122 ( .A(n2594), .B(n2593), .Z(c[1517]) );
  NAND U3123 ( .A(b[0]), .B(a[495]), .Z(n2597) );
  XNOR U3124 ( .A(sreg[1518]), .B(n2597), .Z(n2599) );
  NANDN U3125 ( .A(sreg[1517]), .B(n2592), .Z(n2596) );
  NAND U3126 ( .A(n2594), .B(n2593), .Z(n2595) );
  AND U3127 ( .A(n2596), .B(n2595), .Z(n2598) );
  XOR U3128 ( .A(n2599), .B(n2598), .Z(c[1518]) );
  NANDN U3129 ( .A(n2597), .B(sreg[1518]), .Z(n2601) );
  NAND U3130 ( .A(n2599), .B(n2598), .Z(n2600) );
  AND U3131 ( .A(n2601), .B(n2600), .Z(n2604) );
  NAND U3132 ( .A(b[0]), .B(a[496]), .Z(n2602) );
  XNOR U3133 ( .A(sreg[1519]), .B(n2602), .Z(n2603) );
  XNOR U3134 ( .A(n2604), .B(n2603), .Z(c[1519]) );
  NANDN U3135 ( .A(sreg[1519]), .B(n2602), .Z(n2606) );
  NAND U3136 ( .A(n2604), .B(n2603), .Z(n2605) );
  AND U3137 ( .A(n2606), .B(n2605), .Z(n2609) );
  NAND U3138 ( .A(b[0]), .B(a[497]), .Z(n2607) );
  XNOR U3139 ( .A(sreg[1520]), .B(n2607), .Z(n2608) );
  XOR U3140 ( .A(n2609), .B(n2608), .Z(c[1520]) );
  NAND U3141 ( .A(b[0]), .B(a[498]), .Z(n2612) );
  XNOR U3142 ( .A(sreg[1521]), .B(n2612), .Z(n2614) );
  NANDN U3143 ( .A(n2607), .B(sreg[1520]), .Z(n2611) );
  NAND U3144 ( .A(n2609), .B(n2608), .Z(n2610) );
  AND U3145 ( .A(n2611), .B(n2610), .Z(n2613) );
  XNOR U3146 ( .A(n2614), .B(n2613), .Z(c[1521]) );
  NANDN U3147 ( .A(sreg[1521]), .B(n2612), .Z(n2616) );
  NAND U3148 ( .A(n2614), .B(n2613), .Z(n2615) );
  AND U3149 ( .A(n2616), .B(n2615), .Z(n2619) );
  NAND U3150 ( .A(b[0]), .B(a[499]), .Z(n2617) );
  XNOR U3151 ( .A(sreg[1522]), .B(n2617), .Z(n2618) );
  XOR U3152 ( .A(n2619), .B(n2618), .Z(c[1522]) );
  NAND U3153 ( .A(b[0]), .B(a[500]), .Z(n2622) );
  XNOR U3154 ( .A(sreg[1523]), .B(n2622), .Z(n2624) );
  NANDN U3155 ( .A(n2617), .B(sreg[1522]), .Z(n2621) );
  NAND U3156 ( .A(n2619), .B(n2618), .Z(n2620) );
  NAND U3157 ( .A(n2621), .B(n2620), .Z(n2623) );
  XOR U3158 ( .A(n2624), .B(n2623), .Z(c[1523]) );
  NANDN U3159 ( .A(n2622), .B(sreg[1523]), .Z(n2626) );
  NAND U3160 ( .A(n2624), .B(n2623), .Z(n2625) );
  AND U3161 ( .A(n2626), .B(n2625), .Z(n2629) );
  NAND U3162 ( .A(b[0]), .B(a[501]), .Z(n2627) );
  XNOR U3163 ( .A(sreg[1524]), .B(n2627), .Z(n2628) );
  XNOR U3164 ( .A(n2629), .B(n2628), .Z(c[1524]) );
  NANDN U3165 ( .A(sreg[1524]), .B(n2627), .Z(n2631) );
  NAND U3166 ( .A(n2629), .B(n2628), .Z(n2630) );
  AND U3167 ( .A(n2631), .B(n2630), .Z(n2634) );
  NAND U3168 ( .A(b[0]), .B(a[502]), .Z(n2632) );
  XNOR U3169 ( .A(sreg[1525]), .B(n2632), .Z(n2633) );
  XOR U3170 ( .A(n2634), .B(n2633), .Z(c[1525]) );
  NAND U3171 ( .A(b[0]), .B(a[503]), .Z(n2637) );
  XNOR U3172 ( .A(sreg[1526]), .B(n2637), .Z(n2639) );
  NANDN U3173 ( .A(n2632), .B(sreg[1525]), .Z(n2636) );
  NAND U3174 ( .A(n2634), .B(n2633), .Z(n2635) );
  NAND U3175 ( .A(n2636), .B(n2635), .Z(n2638) );
  XOR U3176 ( .A(n2639), .B(n2638), .Z(c[1526]) );
  NAND U3177 ( .A(b[0]), .B(a[504]), .Z(n2642) );
  XNOR U3178 ( .A(sreg[1527]), .B(n2642), .Z(n2644) );
  NANDN U3179 ( .A(n2637), .B(sreg[1526]), .Z(n2641) );
  NAND U3180 ( .A(n2639), .B(n2638), .Z(n2640) );
  AND U3181 ( .A(n2641), .B(n2640), .Z(n2643) );
  XNOR U3182 ( .A(n2644), .B(n2643), .Z(c[1527]) );
  NAND U3183 ( .A(b[0]), .B(a[505]), .Z(n2647) );
  XNOR U3184 ( .A(sreg[1528]), .B(n2647), .Z(n2649) );
  NANDN U3185 ( .A(sreg[1527]), .B(n2642), .Z(n2646) );
  NAND U3186 ( .A(n2644), .B(n2643), .Z(n2645) );
  AND U3187 ( .A(n2646), .B(n2645), .Z(n2648) );
  XOR U3188 ( .A(n2649), .B(n2648), .Z(c[1528]) );
  NAND U3189 ( .A(b[0]), .B(a[506]), .Z(n2652) );
  XNOR U3190 ( .A(sreg[1529]), .B(n2652), .Z(n2654) );
  NANDN U3191 ( .A(n2647), .B(sreg[1528]), .Z(n2651) );
  NAND U3192 ( .A(n2649), .B(n2648), .Z(n2650) );
  NAND U3193 ( .A(n2651), .B(n2650), .Z(n2653) );
  XOR U3194 ( .A(n2654), .B(n2653), .Z(c[1529]) );
  NAND U3195 ( .A(b[0]), .B(a[507]), .Z(n2657) );
  XNOR U3196 ( .A(sreg[1530]), .B(n2657), .Z(n2659) );
  NANDN U3197 ( .A(n2652), .B(sreg[1529]), .Z(n2656) );
  NAND U3198 ( .A(n2654), .B(n2653), .Z(n2655) );
  NAND U3199 ( .A(n2656), .B(n2655), .Z(n2658) );
  XOR U3200 ( .A(n2659), .B(n2658), .Z(c[1530]) );
  NANDN U3201 ( .A(n2657), .B(sreg[1530]), .Z(n2661) );
  NAND U3202 ( .A(n2659), .B(n2658), .Z(n2660) );
  AND U3203 ( .A(n2661), .B(n2660), .Z(n2664) );
  NAND U3204 ( .A(b[0]), .B(a[508]), .Z(n2662) );
  XNOR U3205 ( .A(sreg[1531]), .B(n2662), .Z(n2663) );
  XNOR U3206 ( .A(n2664), .B(n2663), .Z(c[1531]) );
  NAND U3207 ( .A(b[0]), .B(a[509]), .Z(n2667) );
  XNOR U3208 ( .A(sreg[1532]), .B(n2667), .Z(n2669) );
  NANDN U3209 ( .A(sreg[1531]), .B(n2662), .Z(n2666) );
  NAND U3210 ( .A(n2664), .B(n2663), .Z(n2665) );
  AND U3211 ( .A(n2666), .B(n2665), .Z(n2668) );
  XOR U3212 ( .A(n2669), .B(n2668), .Z(c[1532]) );
  NAND U3213 ( .A(b[0]), .B(a[510]), .Z(n2672) );
  XNOR U3214 ( .A(sreg[1533]), .B(n2672), .Z(n2674) );
  NANDN U3215 ( .A(n2667), .B(sreg[1532]), .Z(n2671) );
  NAND U3216 ( .A(n2669), .B(n2668), .Z(n2670) );
  NAND U3217 ( .A(n2671), .B(n2670), .Z(n2673) );
  XOR U3218 ( .A(n2674), .B(n2673), .Z(c[1533]) );
  NAND U3219 ( .A(b[0]), .B(a[511]), .Z(n2677) );
  XNOR U3220 ( .A(sreg[1534]), .B(n2677), .Z(n2679) );
  NANDN U3221 ( .A(n2672), .B(sreg[1533]), .Z(n2676) );
  NAND U3222 ( .A(n2674), .B(n2673), .Z(n2675) );
  AND U3223 ( .A(n2676), .B(n2675), .Z(n2678) );
  XNOR U3224 ( .A(n2679), .B(n2678), .Z(c[1534]) );
  NANDN U3225 ( .A(sreg[1534]), .B(n2677), .Z(n2681) );
  NAND U3226 ( .A(n2679), .B(n2678), .Z(n2680) );
  AND U3227 ( .A(n2681), .B(n2680), .Z(n2684) );
  NAND U3228 ( .A(b[0]), .B(a[512]), .Z(n2682) );
  XNOR U3229 ( .A(sreg[1535]), .B(n2682), .Z(n2683) );
  XOR U3230 ( .A(n2684), .B(n2683), .Z(c[1535]) );
  NAND U3231 ( .A(b[0]), .B(a[513]), .Z(n2687) );
  XNOR U3232 ( .A(sreg[1536]), .B(n2687), .Z(n2689) );
  NANDN U3233 ( .A(n2682), .B(sreg[1535]), .Z(n2686) );
  NAND U3234 ( .A(n2684), .B(n2683), .Z(n2685) );
  NAND U3235 ( .A(n2686), .B(n2685), .Z(n2688) );
  XOR U3236 ( .A(n2689), .B(n2688), .Z(c[1536]) );
  NANDN U3237 ( .A(n2687), .B(sreg[1536]), .Z(n2691) );
  NAND U3238 ( .A(n2689), .B(n2688), .Z(n2690) );
  AND U3239 ( .A(n2691), .B(n2690), .Z(n2694) );
  NAND U3240 ( .A(b[0]), .B(a[514]), .Z(n2692) );
  XNOR U3241 ( .A(sreg[1537]), .B(n2692), .Z(n2693) );
  XNOR U3242 ( .A(n2694), .B(n2693), .Z(c[1537]) );
  NANDN U3243 ( .A(sreg[1537]), .B(n2692), .Z(n2696) );
  NAND U3244 ( .A(n2694), .B(n2693), .Z(n2695) );
  AND U3245 ( .A(n2696), .B(n2695), .Z(n2699) );
  NAND U3246 ( .A(b[0]), .B(a[515]), .Z(n2697) );
  XNOR U3247 ( .A(sreg[1538]), .B(n2697), .Z(n2698) );
  XOR U3248 ( .A(n2699), .B(n2698), .Z(c[1538]) );
  NAND U3249 ( .A(b[0]), .B(a[516]), .Z(n2702) );
  XNOR U3250 ( .A(sreg[1539]), .B(n2702), .Z(n2704) );
  NANDN U3251 ( .A(n2697), .B(sreg[1538]), .Z(n2701) );
  NAND U3252 ( .A(n2699), .B(n2698), .Z(n2700) );
  AND U3253 ( .A(n2701), .B(n2700), .Z(n2703) );
  XNOR U3254 ( .A(n2704), .B(n2703), .Z(c[1539]) );
  NANDN U3255 ( .A(sreg[1539]), .B(n2702), .Z(n2706) );
  NAND U3256 ( .A(n2704), .B(n2703), .Z(n2705) );
  AND U3257 ( .A(n2706), .B(n2705), .Z(n2709) );
  NAND U3258 ( .A(b[0]), .B(a[517]), .Z(n2707) );
  XNOR U3259 ( .A(sreg[1540]), .B(n2707), .Z(n2708) );
  XOR U3260 ( .A(n2709), .B(n2708), .Z(c[1540]) );
  NAND U3261 ( .A(b[0]), .B(a[518]), .Z(n2712) );
  XNOR U3262 ( .A(sreg[1541]), .B(n2712), .Z(n2714) );
  NANDN U3263 ( .A(n2707), .B(sreg[1540]), .Z(n2711) );
  NAND U3264 ( .A(n2709), .B(n2708), .Z(n2710) );
  NAND U3265 ( .A(n2711), .B(n2710), .Z(n2713) );
  XOR U3266 ( .A(n2714), .B(n2713), .Z(c[1541]) );
  NANDN U3267 ( .A(n2712), .B(sreg[1541]), .Z(n2716) );
  NAND U3268 ( .A(n2714), .B(n2713), .Z(n2715) );
  AND U3269 ( .A(n2716), .B(n2715), .Z(n2719) );
  NAND U3270 ( .A(b[0]), .B(a[519]), .Z(n2717) );
  XNOR U3271 ( .A(sreg[1542]), .B(n2717), .Z(n2718) );
  XNOR U3272 ( .A(n2719), .B(n2718), .Z(c[1542]) );
  NAND U3273 ( .A(b[0]), .B(a[520]), .Z(n2722) );
  XNOR U3274 ( .A(sreg[1543]), .B(n2722), .Z(n2724) );
  NANDN U3275 ( .A(sreg[1542]), .B(n2717), .Z(n2721) );
  NAND U3276 ( .A(n2719), .B(n2718), .Z(n2720) );
  AND U3277 ( .A(n2721), .B(n2720), .Z(n2723) );
  XOR U3278 ( .A(n2724), .B(n2723), .Z(c[1543]) );
  NAND U3279 ( .A(b[0]), .B(a[521]), .Z(n2727) );
  XNOR U3280 ( .A(sreg[1544]), .B(n2727), .Z(n2729) );
  NANDN U3281 ( .A(n2722), .B(sreg[1543]), .Z(n2726) );
  NAND U3282 ( .A(n2724), .B(n2723), .Z(n2725) );
  NAND U3283 ( .A(n2726), .B(n2725), .Z(n2728) );
  XOR U3284 ( .A(n2729), .B(n2728), .Z(c[1544]) );
  NAND U3285 ( .A(b[0]), .B(a[522]), .Z(n2732) );
  XNOR U3286 ( .A(sreg[1545]), .B(n2732), .Z(n2734) );
  NANDN U3287 ( .A(n2727), .B(sreg[1544]), .Z(n2731) );
  NAND U3288 ( .A(n2729), .B(n2728), .Z(n2730) );
  AND U3289 ( .A(n2731), .B(n2730), .Z(n2733) );
  XNOR U3290 ( .A(n2734), .B(n2733), .Z(c[1545]) );
  NAND U3291 ( .A(b[0]), .B(a[523]), .Z(n2737) );
  XNOR U3292 ( .A(sreg[1546]), .B(n2737), .Z(n2739) );
  NANDN U3293 ( .A(sreg[1545]), .B(n2732), .Z(n2736) );
  NAND U3294 ( .A(n2734), .B(n2733), .Z(n2735) );
  NAND U3295 ( .A(n2736), .B(n2735), .Z(n2738) );
  XNOR U3296 ( .A(n2739), .B(n2738), .Z(c[1546]) );
  NANDN U3297 ( .A(sreg[1546]), .B(n2737), .Z(n2741) );
  NAND U3298 ( .A(n2739), .B(n2738), .Z(n2740) );
  AND U3299 ( .A(n2741), .B(n2740), .Z(n2744) );
  NAND U3300 ( .A(b[0]), .B(a[524]), .Z(n2742) );
  XNOR U3301 ( .A(sreg[1547]), .B(n2742), .Z(n2743) );
  XOR U3302 ( .A(n2744), .B(n2743), .Z(c[1547]) );
  NAND U3303 ( .A(b[0]), .B(a[525]), .Z(n2747) );
  XNOR U3304 ( .A(sreg[1548]), .B(n2747), .Z(n2749) );
  NANDN U3305 ( .A(n2742), .B(sreg[1547]), .Z(n2746) );
  NAND U3306 ( .A(n2744), .B(n2743), .Z(n2745) );
  AND U3307 ( .A(n2746), .B(n2745), .Z(n2748) );
  XNOR U3308 ( .A(n2749), .B(n2748), .Z(c[1548]) );
  NAND U3309 ( .A(b[0]), .B(a[526]), .Z(n2752) );
  XNOR U3310 ( .A(sreg[1549]), .B(n2752), .Z(n2754) );
  NANDN U3311 ( .A(sreg[1548]), .B(n2747), .Z(n2751) );
  NAND U3312 ( .A(n2749), .B(n2748), .Z(n2750) );
  NAND U3313 ( .A(n2751), .B(n2750), .Z(n2753) );
  XNOR U3314 ( .A(n2754), .B(n2753), .Z(c[1549]) );
  NANDN U3315 ( .A(sreg[1549]), .B(n2752), .Z(n2756) );
  NAND U3316 ( .A(n2754), .B(n2753), .Z(n2755) );
  AND U3317 ( .A(n2756), .B(n2755), .Z(n2759) );
  NAND U3318 ( .A(b[0]), .B(a[527]), .Z(n2757) );
  XNOR U3319 ( .A(sreg[1550]), .B(n2757), .Z(n2758) );
  XOR U3320 ( .A(n2759), .B(n2758), .Z(c[1550]) );
  NANDN U3321 ( .A(n2757), .B(sreg[1550]), .Z(n2761) );
  NAND U3322 ( .A(n2759), .B(n2758), .Z(n2760) );
  AND U3323 ( .A(n2761), .B(n2760), .Z(n2764) );
  NAND U3324 ( .A(b[0]), .B(a[528]), .Z(n2762) );
  XNOR U3325 ( .A(sreg[1551]), .B(n2762), .Z(n2763) );
  XNOR U3326 ( .A(n2764), .B(n2763), .Z(c[1551]) );
  NAND U3327 ( .A(b[0]), .B(a[529]), .Z(n2767) );
  XNOR U3328 ( .A(sreg[1552]), .B(n2767), .Z(n2769) );
  NANDN U3329 ( .A(sreg[1551]), .B(n2762), .Z(n2766) );
  NAND U3330 ( .A(n2764), .B(n2763), .Z(n2765) );
  NAND U3331 ( .A(n2766), .B(n2765), .Z(n2768) );
  XNOR U3332 ( .A(n2769), .B(n2768), .Z(c[1552]) );
  NANDN U3333 ( .A(sreg[1552]), .B(n2767), .Z(n2771) );
  NAND U3334 ( .A(n2769), .B(n2768), .Z(n2770) );
  AND U3335 ( .A(n2771), .B(n2770), .Z(n2774) );
  NAND U3336 ( .A(b[0]), .B(a[530]), .Z(n2772) );
  XNOR U3337 ( .A(sreg[1553]), .B(n2772), .Z(n2773) );
  XOR U3338 ( .A(n2774), .B(n2773), .Z(c[1553]) );
  NAND U3339 ( .A(b[0]), .B(a[531]), .Z(n2777) );
  XNOR U3340 ( .A(sreg[1554]), .B(n2777), .Z(n2779) );
  NANDN U3341 ( .A(n2772), .B(sreg[1553]), .Z(n2776) );
  NAND U3342 ( .A(n2774), .B(n2773), .Z(n2775) );
  AND U3343 ( .A(n2776), .B(n2775), .Z(n2778) );
  XNOR U3344 ( .A(n2779), .B(n2778), .Z(c[1554]) );
  NAND U3345 ( .A(b[0]), .B(a[532]), .Z(n2782) );
  XNOR U3346 ( .A(sreg[1555]), .B(n2782), .Z(n2784) );
  NANDN U3347 ( .A(sreg[1554]), .B(n2777), .Z(n2781) );
  NAND U3348 ( .A(n2779), .B(n2778), .Z(n2780) );
  NAND U3349 ( .A(n2781), .B(n2780), .Z(n2783) );
  XNOR U3350 ( .A(n2784), .B(n2783), .Z(c[1555]) );
  NAND U3351 ( .A(b[0]), .B(a[533]), .Z(n2787) );
  XNOR U3352 ( .A(sreg[1556]), .B(n2787), .Z(n2789) );
  NANDN U3353 ( .A(sreg[1555]), .B(n2782), .Z(n2786) );
  NAND U3354 ( .A(n2784), .B(n2783), .Z(n2785) );
  AND U3355 ( .A(n2786), .B(n2785), .Z(n2788) );
  XOR U3356 ( .A(n2789), .B(n2788), .Z(c[1556]) );
  NAND U3357 ( .A(b[0]), .B(a[534]), .Z(n2792) );
  XNOR U3358 ( .A(sreg[1557]), .B(n2792), .Z(n2794) );
  NANDN U3359 ( .A(n2787), .B(sreg[1556]), .Z(n2791) );
  NAND U3360 ( .A(n2789), .B(n2788), .Z(n2790) );
  NAND U3361 ( .A(n2791), .B(n2790), .Z(n2793) );
  XOR U3362 ( .A(n2794), .B(n2793), .Z(c[1557]) );
  NAND U3363 ( .A(b[0]), .B(a[535]), .Z(n2797) );
  XNOR U3364 ( .A(sreg[1558]), .B(n2797), .Z(n2799) );
  NANDN U3365 ( .A(n2792), .B(sreg[1557]), .Z(n2796) );
  NAND U3366 ( .A(n2794), .B(n2793), .Z(n2795) );
  NAND U3367 ( .A(n2796), .B(n2795), .Z(n2798) );
  XOR U3368 ( .A(n2799), .B(n2798), .Z(c[1558]) );
  NAND U3369 ( .A(b[0]), .B(a[536]), .Z(n2802) );
  XNOR U3370 ( .A(sreg[1559]), .B(n2802), .Z(n2804) );
  NANDN U3371 ( .A(n2797), .B(sreg[1558]), .Z(n2801) );
  NAND U3372 ( .A(n2799), .B(n2798), .Z(n2800) );
  NAND U3373 ( .A(n2801), .B(n2800), .Z(n2803) );
  XOR U3374 ( .A(n2804), .B(n2803), .Z(c[1559]) );
  NAND U3375 ( .A(b[0]), .B(a[537]), .Z(n2807) );
  XNOR U3376 ( .A(sreg[1560]), .B(n2807), .Z(n2809) );
  NANDN U3377 ( .A(n2802), .B(sreg[1559]), .Z(n2806) );
  NAND U3378 ( .A(n2804), .B(n2803), .Z(n2805) );
  NAND U3379 ( .A(n2806), .B(n2805), .Z(n2808) );
  XOR U3380 ( .A(n2809), .B(n2808), .Z(c[1560]) );
  NAND U3381 ( .A(b[0]), .B(a[538]), .Z(n2812) );
  XNOR U3382 ( .A(sreg[1561]), .B(n2812), .Z(n2814) );
  NANDN U3383 ( .A(n2807), .B(sreg[1560]), .Z(n2811) );
  NAND U3384 ( .A(n2809), .B(n2808), .Z(n2810) );
  NAND U3385 ( .A(n2811), .B(n2810), .Z(n2813) );
  XOR U3386 ( .A(n2814), .B(n2813), .Z(c[1561]) );
  NANDN U3387 ( .A(n2812), .B(sreg[1561]), .Z(n2816) );
  NAND U3388 ( .A(n2814), .B(n2813), .Z(n2815) );
  NAND U3389 ( .A(n2816), .B(n2815), .Z(n2818) );
  AND U3390 ( .A(b[0]), .B(a[539]), .Z(n2819) );
  XNOR U3391 ( .A(n2819), .B(sreg[1562]), .Z(n2817) );
  XNOR U3392 ( .A(n2818), .B(n2817), .Z(c[1562]) );
  NAND U3393 ( .A(b[0]), .B(a[540]), .Z(n2820) );
  XNOR U3394 ( .A(sreg[1563]), .B(n2820), .Z(n2821) );
  XOR U3395 ( .A(n2822), .B(n2821), .Z(c[1563]) );
  NAND U3396 ( .A(b[0]), .B(a[541]), .Z(n2825) );
  XNOR U3397 ( .A(sreg[1564]), .B(n2825), .Z(n2827) );
  NANDN U3398 ( .A(n2820), .B(sreg[1563]), .Z(n2824) );
  NAND U3399 ( .A(n2822), .B(n2821), .Z(n2823) );
  NAND U3400 ( .A(n2824), .B(n2823), .Z(n2826) );
  XOR U3401 ( .A(n2827), .B(n2826), .Z(c[1564]) );
  NAND U3402 ( .A(b[0]), .B(a[542]), .Z(n2830) );
  XNOR U3403 ( .A(sreg[1565]), .B(n2830), .Z(n2832) );
  NANDN U3404 ( .A(n2825), .B(sreg[1564]), .Z(n2829) );
  NAND U3405 ( .A(n2827), .B(n2826), .Z(n2828) );
  AND U3406 ( .A(n2829), .B(n2828), .Z(n2831) );
  XNOR U3407 ( .A(n2832), .B(n2831), .Z(c[1565]) );
  NANDN U3408 ( .A(sreg[1565]), .B(n2830), .Z(n2834) );
  NAND U3409 ( .A(n2832), .B(n2831), .Z(n2833) );
  AND U3410 ( .A(n2834), .B(n2833), .Z(n2837) );
  NAND U3411 ( .A(b[0]), .B(a[543]), .Z(n2835) );
  XNOR U3412 ( .A(sreg[1566]), .B(n2835), .Z(n2836) );
  XOR U3413 ( .A(n2837), .B(n2836), .Z(c[1566]) );
  NAND U3414 ( .A(b[0]), .B(a[544]), .Z(n2840) );
  XNOR U3415 ( .A(sreg[1567]), .B(n2840), .Z(n2842) );
  NANDN U3416 ( .A(n2835), .B(sreg[1566]), .Z(n2839) );
  NAND U3417 ( .A(n2837), .B(n2836), .Z(n2838) );
  NAND U3418 ( .A(n2839), .B(n2838), .Z(n2841) );
  XOR U3419 ( .A(n2842), .B(n2841), .Z(c[1567]) );
  NAND U3420 ( .A(b[0]), .B(a[545]), .Z(n2845) );
  XNOR U3421 ( .A(sreg[1568]), .B(n2845), .Z(n2847) );
  NANDN U3422 ( .A(n2840), .B(sreg[1567]), .Z(n2844) );
  NAND U3423 ( .A(n2842), .B(n2841), .Z(n2843) );
  NAND U3424 ( .A(n2844), .B(n2843), .Z(n2846) );
  XOR U3425 ( .A(n2847), .B(n2846), .Z(c[1568]) );
  NAND U3426 ( .A(b[0]), .B(a[546]), .Z(n2850) );
  XNOR U3427 ( .A(sreg[1569]), .B(n2850), .Z(n2852) );
  NANDN U3428 ( .A(n2845), .B(sreg[1568]), .Z(n2849) );
  NAND U3429 ( .A(n2847), .B(n2846), .Z(n2848) );
  NAND U3430 ( .A(n2849), .B(n2848), .Z(n2851) );
  XOR U3431 ( .A(n2852), .B(n2851), .Z(c[1569]) );
  NAND U3432 ( .A(b[0]), .B(a[547]), .Z(n2855) );
  XNOR U3433 ( .A(sreg[1570]), .B(n2855), .Z(n2857) );
  NANDN U3434 ( .A(n2850), .B(sreg[1569]), .Z(n2854) );
  NAND U3435 ( .A(n2852), .B(n2851), .Z(n2853) );
  NAND U3436 ( .A(n2854), .B(n2853), .Z(n2856) );
  XOR U3437 ( .A(n2857), .B(n2856), .Z(c[1570]) );
  NAND U3438 ( .A(b[0]), .B(a[548]), .Z(n2860) );
  XNOR U3439 ( .A(sreg[1571]), .B(n2860), .Z(n2862) );
  NANDN U3440 ( .A(n2855), .B(sreg[1570]), .Z(n2859) );
  NAND U3441 ( .A(n2857), .B(n2856), .Z(n2858) );
  NAND U3442 ( .A(n2859), .B(n2858), .Z(n2861) );
  XOR U3443 ( .A(n2862), .B(n2861), .Z(c[1571]) );
  NAND U3444 ( .A(b[0]), .B(a[549]), .Z(n2865) );
  XNOR U3445 ( .A(sreg[1572]), .B(n2865), .Z(n2867) );
  NANDN U3446 ( .A(n2860), .B(sreg[1571]), .Z(n2864) );
  NAND U3447 ( .A(n2862), .B(n2861), .Z(n2863) );
  NAND U3448 ( .A(n2864), .B(n2863), .Z(n2866) );
  XOR U3449 ( .A(n2867), .B(n2866), .Z(c[1572]) );
  NAND U3450 ( .A(b[0]), .B(a[550]), .Z(n2870) );
  XNOR U3451 ( .A(sreg[1573]), .B(n2870), .Z(n2872) );
  NANDN U3452 ( .A(n2865), .B(sreg[1572]), .Z(n2869) );
  NAND U3453 ( .A(n2867), .B(n2866), .Z(n2868) );
  NAND U3454 ( .A(n2869), .B(n2868), .Z(n2871) );
  XOR U3455 ( .A(n2872), .B(n2871), .Z(c[1573]) );
  NAND U3456 ( .A(b[0]), .B(a[551]), .Z(n2875) );
  XNOR U3457 ( .A(sreg[1574]), .B(n2875), .Z(n2877) );
  NANDN U3458 ( .A(n2870), .B(sreg[1573]), .Z(n2874) );
  NAND U3459 ( .A(n2872), .B(n2871), .Z(n2873) );
  NAND U3460 ( .A(n2874), .B(n2873), .Z(n2876) );
  XOR U3461 ( .A(n2877), .B(n2876), .Z(c[1574]) );
  NAND U3462 ( .A(b[0]), .B(a[552]), .Z(n2880) );
  XNOR U3463 ( .A(sreg[1575]), .B(n2880), .Z(n2882) );
  NANDN U3464 ( .A(n2875), .B(sreg[1574]), .Z(n2879) );
  NAND U3465 ( .A(n2877), .B(n2876), .Z(n2878) );
  NAND U3466 ( .A(n2879), .B(n2878), .Z(n2881) );
  XOR U3467 ( .A(n2882), .B(n2881), .Z(c[1575]) );
  NAND U3468 ( .A(b[0]), .B(a[553]), .Z(n2885) );
  XNOR U3469 ( .A(sreg[1576]), .B(n2885), .Z(n2887) );
  NANDN U3470 ( .A(n2880), .B(sreg[1575]), .Z(n2884) );
  NAND U3471 ( .A(n2882), .B(n2881), .Z(n2883) );
  NAND U3472 ( .A(n2884), .B(n2883), .Z(n2886) );
  XOR U3473 ( .A(n2887), .B(n2886), .Z(c[1576]) );
  NAND U3474 ( .A(b[0]), .B(a[554]), .Z(n2890) );
  XNOR U3475 ( .A(sreg[1577]), .B(n2890), .Z(n2892) );
  NANDN U3476 ( .A(n2885), .B(sreg[1576]), .Z(n2889) );
  NAND U3477 ( .A(n2887), .B(n2886), .Z(n2888) );
  NAND U3478 ( .A(n2889), .B(n2888), .Z(n2891) );
  XOR U3479 ( .A(n2892), .B(n2891), .Z(c[1577]) );
  NAND U3480 ( .A(b[0]), .B(a[555]), .Z(n2895) );
  XNOR U3481 ( .A(sreg[1578]), .B(n2895), .Z(n2897) );
  NANDN U3482 ( .A(n2890), .B(sreg[1577]), .Z(n2894) );
  NAND U3483 ( .A(n2892), .B(n2891), .Z(n2893) );
  NAND U3484 ( .A(n2894), .B(n2893), .Z(n2896) );
  XOR U3485 ( .A(n2897), .B(n2896), .Z(c[1578]) );
  NAND U3486 ( .A(b[0]), .B(a[556]), .Z(n2900) );
  XNOR U3487 ( .A(sreg[1579]), .B(n2900), .Z(n2902) );
  NANDN U3488 ( .A(n2895), .B(sreg[1578]), .Z(n2899) );
  NAND U3489 ( .A(n2897), .B(n2896), .Z(n2898) );
  NAND U3490 ( .A(n2899), .B(n2898), .Z(n2901) );
  XOR U3491 ( .A(n2902), .B(n2901), .Z(c[1579]) );
  NAND U3492 ( .A(b[0]), .B(a[557]), .Z(n2905) );
  XNOR U3493 ( .A(sreg[1580]), .B(n2905), .Z(n2907) );
  NANDN U3494 ( .A(n2900), .B(sreg[1579]), .Z(n2904) );
  NAND U3495 ( .A(n2902), .B(n2901), .Z(n2903) );
  NAND U3496 ( .A(n2904), .B(n2903), .Z(n2906) );
  XOR U3497 ( .A(n2907), .B(n2906), .Z(c[1580]) );
  NAND U3498 ( .A(b[0]), .B(a[558]), .Z(n2910) );
  XNOR U3499 ( .A(sreg[1581]), .B(n2910), .Z(n2912) );
  NANDN U3500 ( .A(n2905), .B(sreg[1580]), .Z(n2909) );
  NAND U3501 ( .A(n2907), .B(n2906), .Z(n2908) );
  NAND U3502 ( .A(n2909), .B(n2908), .Z(n2911) );
  XOR U3503 ( .A(n2912), .B(n2911), .Z(c[1581]) );
  NAND U3504 ( .A(b[0]), .B(a[559]), .Z(n2915) );
  XNOR U3505 ( .A(sreg[1582]), .B(n2915), .Z(n2917) );
  NANDN U3506 ( .A(n2910), .B(sreg[1581]), .Z(n2914) );
  NAND U3507 ( .A(n2912), .B(n2911), .Z(n2913) );
  NAND U3508 ( .A(n2914), .B(n2913), .Z(n2916) );
  XOR U3509 ( .A(n2917), .B(n2916), .Z(c[1582]) );
  NAND U3510 ( .A(b[0]), .B(a[560]), .Z(n2920) );
  XNOR U3511 ( .A(sreg[1583]), .B(n2920), .Z(n2922) );
  NANDN U3512 ( .A(n2915), .B(sreg[1582]), .Z(n2919) );
  NAND U3513 ( .A(n2917), .B(n2916), .Z(n2918) );
  NAND U3514 ( .A(n2919), .B(n2918), .Z(n2921) );
  XOR U3515 ( .A(n2922), .B(n2921), .Z(c[1583]) );
  NAND U3516 ( .A(b[0]), .B(a[561]), .Z(n2925) );
  XNOR U3517 ( .A(sreg[1584]), .B(n2925), .Z(n2927) );
  NANDN U3518 ( .A(n2920), .B(sreg[1583]), .Z(n2924) );
  NAND U3519 ( .A(n2922), .B(n2921), .Z(n2923) );
  NAND U3520 ( .A(n2924), .B(n2923), .Z(n2926) );
  XOR U3521 ( .A(n2927), .B(n2926), .Z(c[1584]) );
  NAND U3522 ( .A(b[0]), .B(a[562]), .Z(n2930) );
  XNOR U3523 ( .A(sreg[1585]), .B(n2930), .Z(n2932) );
  NANDN U3524 ( .A(n2925), .B(sreg[1584]), .Z(n2929) );
  NAND U3525 ( .A(n2927), .B(n2926), .Z(n2928) );
  NAND U3526 ( .A(n2929), .B(n2928), .Z(n2931) );
  XOR U3527 ( .A(n2932), .B(n2931), .Z(c[1585]) );
  NAND U3528 ( .A(b[0]), .B(a[563]), .Z(n2935) );
  XNOR U3529 ( .A(sreg[1586]), .B(n2935), .Z(n2937) );
  NANDN U3530 ( .A(n2930), .B(sreg[1585]), .Z(n2934) );
  NAND U3531 ( .A(n2932), .B(n2931), .Z(n2933) );
  NAND U3532 ( .A(n2934), .B(n2933), .Z(n2936) );
  XOR U3533 ( .A(n2937), .B(n2936), .Z(c[1586]) );
  NAND U3534 ( .A(b[0]), .B(a[564]), .Z(n2940) );
  XNOR U3535 ( .A(sreg[1587]), .B(n2940), .Z(n2942) );
  NANDN U3536 ( .A(n2935), .B(sreg[1586]), .Z(n2939) );
  NAND U3537 ( .A(n2937), .B(n2936), .Z(n2938) );
  NAND U3538 ( .A(n2939), .B(n2938), .Z(n2941) );
  XOR U3539 ( .A(n2942), .B(n2941), .Z(c[1587]) );
  NAND U3540 ( .A(b[0]), .B(a[565]), .Z(n2945) );
  XNOR U3541 ( .A(sreg[1588]), .B(n2945), .Z(n2947) );
  NANDN U3542 ( .A(n2940), .B(sreg[1587]), .Z(n2944) );
  NAND U3543 ( .A(n2942), .B(n2941), .Z(n2943) );
  NAND U3544 ( .A(n2944), .B(n2943), .Z(n2946) );
  XOR U3545 ( .A(n2947), .B(n2946), .Z(c[1588]) );
  NAND U3546 ( .A(b[0]), .B(a[566]), .Z(n2950) );
  XNOR U3547 ( .A(sreg[1589]), .B(n2950), .Z(n2952) );
  NANDN U3548 ( .A(n2945), .B(sreg[1588]), .Z(n2949) );
  NAND U3549 ( .A(n2947), .B(n2946), .Z(n2948) );
  NAND U3550 ( .A(n2949), .B(n2948), .Z(n2951) );
  XOR U3551 ( .A(n2952), .B(n2951), .Z(c[1589]) );
  NAND U3552 ( .A(b[0]), .B(a[567]), .Z(n2955) );
  XNOR U3553 ( .A(sreg[1590]), .B(n2955), .Z(n2957) );
  NANDN U3554 ( .A(n2950), .B(sreg[1589]), .Z(n2954) );
  NAND U3555 ( .A(n2952), .B(n2951), .Z(n2953) );
  NAND U3556 ( .A(n2954), .B(n2953), .Z(n2956) );
  XOR U3557 ( .A(n2957), .B(n2956), .Z(c[1590]) );
  NAND U3558 ( .A(b[0]), .B(a[568]), .Z(n2960) );
  XNOR U3559 ( .A(sreg[1591]), .B(n2960), .Z(n2962) );
  NANDN U3560 ( .A(n2955), .B(sreg[1590]), .Z(n2959) );
  NAND U3561 ( .A(n2957), .B(n2956), .Z(n2958) );
  NAND U3562 ( .A(n2959), .B(n2958), .Z(n2961) );
  XOR U3563 ( .A(n2962), .B(n2961), .Z(c[1591]) );
  NAND U3564 ( .A(b[0]), .B(a[569]), .Z(n2965) );
  XNOR U3565 ( .A(sreg[1592]), .B(n2965), .Z(n2967) );
  NANDN U3566 ( .A(n2960), .B(sreg[1591]), .Z(n2964) );
  NAND U3567 ( .A(n2962), .B(n2961), .Z(n2963) );
  NAND U3568 ( .A(n2964), .B(n2963), .Z(n2966) );
  XOR U3569 ( .A(n2967), .B(n2966), .Z(c[1592]) );
  NAND U3570 ( .A(b[0]), .B(a[570]), .Z(n2970) );
  XNOR U3571 ( .A(sreg[1593]), .B(n2970), .Z(n2972) );
  NANDN U3572 ( .A(n2965), .B(sreg[1592]), .Z(n2969) );
  NAND U3573 ( .A(n2967), .B(n2966), .Z(n2968) );
  NAND U3574 ( .A(n2969), .B(n2968), .Z(n2971) );
  XOR U3575 ( .A(n2972), .B(n2971), .Z(c[1593]) );
  NAND U3576 ( .A(b[0]), .B(a[571]), .Z(n2975) );
  XNOR U3577 ( .A(sreg[1594]), .B(n2975), .Z(n2977) );
  NANDN U3578 ( .A(n2970), .B(sreg[1593]), .Z(n2974) );
  NAND U3579 ( .A(n2972), .B(n2971), .Z(n2973) );
  NAND U3580 ( .A(n2974), .B(n2973), .Z(n2976) );
  XOR U3581 ( .A(n2977), .B(n2976), .Z(c[1594]) );
  NANDN U3582 ( .A(n2975), .B(sreg[1594]), .Z(n2979) );
  NAND U3583 ( .A(n2977), .B(n2976), .Z(n2978) );
  AND U3584 ( .A(n2979), .B(n2978), .Z(n2982) );
  NAND U3585 ( .A(b[0]), .B(a[572]), .Z(n2980) );
  XNOR U3586 ( .A(sreg[1595]), .B(n2980), .Z(n2981) );
  XNOR U3587 ( .A(n2982), .B(n2981), .Z(c[1595]) );
  NAND U3588 ( .A(b[0]), .B(a[573]), .Z(n2985) );
  XNOR U3589 ( .A(sreg[1596]), .B(n2985), .Z(n2987) );
  NANDN U3590 ( .A(sreg[1595]), .B(n2980), .Z(n2984) );
  NAND U3591 ( .A(n2982), .B(n2981), .Z(n2983) );
  AND U3592 ( .A(n2984), .B(n2983), .Z(n2986) );
  XOR U3593 ( .A(n2987), .B(n2986), .Z(c[1596]) );
  NANDN U3594 ( .A(n2985), .B(sreg[1596]), .Z(n2989) );
  NAND U3595 ( .A(n2987), .B(n2986), .Z(n2988) );
  AND U3596 ( .A(n2989), .B(n2988), .Z(n2992) );
  NAND U3597 ( .A(b[0]), .B(a[574]), .Z(n2990) );
  XNOR U3598 ( .A(sreg[1597]), .B(n2990), .Z(n2991) );
  XNOR U3599 ( .A(n2992), .B(n2991), .Z(c[1597]) );
  NAND U3600 ( .A(b[0]), .B(a[575]), .Z(n2995) );
  XNOR U3601 ( .A(sreg[1598]), .B(n2995), .Z(n2997) );
  NANDN U3602 ( .A(sreg[1597]), .B(n2990), .Z(n2994) );
  NAND U3603 ( .A(n2992), .B(n2991), .Z(n2993) );
  NAND U3604 ( .A(n2994), .B(n2993), .Z(n2996) );
  XNOR U3605 ( .A(n2997), .B(n2996), .Z(c[1598]) );
  NAND U3606 ( .A(b[0]), .B(a[576]), .Z(n3000) );
  XNOR U3607 ( .A(sreg[1599]), .B(n3000), .Z(n3002) );
  NANDN U3608 ( .A(sreg[1598]), .B(n2995), .Z(n2999) );
  NAND U3609 ( .A(n2997), .B(n2996), .Z(n2998) );
  AND U3610 ( .A(n2999), .B(n2998), .Z(n3001) );
  XOR U3611 ( .A(n3002), .B(n3001), .Z(c[1599]) );
  NANDN U3612 ( .A(n3000), .B(sreg[1599]), .Z(n3004) );
  NAND U3613 ( .A(n3002), .B(n3001), .Z(n3003) );
  AND U3614 ( .A(n3004), .B(n3003), .Z(n3007) );
  NAND U3615 ( .A(b[0]), .B(a[577]), .Z(n3005) );
  XNOR U3616 ( .A(sreg[1600]), .B(n3005), .Z(n3006) );
  XNOR U3617 ( .A(n3007), .B(n3006), .Z(c[1600]) );
  NAND U3618 ( .A(b[0]), .B(a[578]), .Z(n3010) );
  XNOR U3619 ( .A(sreg[1601]), .B(n3010), .Z(n3012) );
  NANDN U3620 ( .A(sreg[1600]), .B(n3005), .Z(n3009) );
  NAND U3621 ( .A(n3007), .B(n3006), .Z(n3008) );
  NAND U3622 ( .A(n3009), .B(n3008), .Z(n3011) );
  XNOR U3623 ( .A(n3012), .B(n3011), .Z(c[1601]) );
  NAND U3624 ( .A(b[0]), .B(a[579]), .Z(n3015) );
  XNOR U3625 ( .A(sreg[1602]), .B(n3015), .Z(n3017) );
  NANDN U3626 ( .A(sreg[1601]), .B(n3010), .Z(n3014) );
  NAND U3627 ( .A(n3012), .B(n3011), .Z(n3013) );
  NAND U3628 ( .A(n3014), .B(n3013), .Z(n3016) );
  XNOR U3629 ( .A(n3017), .B(n3016), .Z(c[1602]) );
  NAND U3630 ( .A(b[0]), .B(a[580]), .Z(n3020) );
  XNOR U3631 ( .A(sreg[1603]), .B(n3020), .Z(n3022) );
  NANDN U3632 ( .A(sreg[1602]), .B(n3015), .Z(n3019) );
  NAND U3633 ( .A(n3017), .B(n3016), .Z(n3018) );
  NAND U3634 ( .A(n3019), .B(n3018), .Z(n3021) );
  XNOR U3635 ( .A(n3022), .B(n3021), .Z(c[1603]) );
  NAND U3636 ( .A(b[0]), .B(a[581]), .Z(n3025) );
  XNOR U3637 ( .A(sreg[1604]), .B(n3025), .Z(n3027) );
  NANDN U3638 ( .A(sreg[1603]), .B(n3020), .Z(n3024) );
  NAND U3639 ( .A(n3022), .B(n3021), .Z(n3023) );
  NAND U3640 ( .A(n3024), .B(n3023), .Z(n3026) );
  XNOR U3641 ( .A(n3027), .B(n3026), .Z(c[1604]) );
  NAND U3642 ( .A(b[0]), .B(a[582]), .Z(n3030) );
  XNOR U3643 ( .A(sreg[1605]), .B(n3030), .Z(n3032) );
  NANDN U3644 ( .A(sreg[1604]), .B(n3025), .Z(n3029) );
  NAND U3645 ( .A(n3027), .B(n3026), .Z(n3028) );
  NAND U3646 ( .A(n3029), .B(n3028), .Z(n3031) );
  XNOR U3647 ( .A(n3032), .B(n3031), .Z(c[1605]) );
  NAND U3648 ( .A(b[0]), .B(a[583]), .Z(n3035) );
  XNOR U3649 ( .A(sreg[1606]), .B(n3035), .Z(n3037) );
  NANDN U3650 ( .A(sreg[1605]), .B(n3030), .Z(n3034) );
  NAND U3651 ( .A(n3032), .B(n3031), .Z(n3033) );
  NAND U3652 ( .A(n3034), .B(n3033), .Z(n3036) );
  XNOR U3653 ( .A(n3037), .B(n3036), .Z(c[1606]) );
  NAND U3654 ( .A(b[0]), .B(a[584]), .Z(n3040) );
  XNOR U3655 ( .A(sreg[1607]), .B(n3040), .Z(n3042) );
  NANDN U3656 ( .A(sreg[1606]), .B(n3035), .Z(n3039) );
  NAND U3657 ( .A(n3037), .B(n3036), .Z(n3038) );
  NAND U3658 ( .A(n3039), .B(n3038), .Z(n3041) );
  XNOR U3659 ( .A(n3042), .B(n3041), .Z(c[1607]) );
  NAND U3660 ( .A(b[0]), .B(a[585]), .Z(n3045) );
  XNOR U3661 ( .A(sreg[1608]), .B(n3045), .Z(n3047) );
  NANDN U3662 ( .A(sreg[1607]), .B(n3040), .Z(n3044) );
  NAND U3663 ( .A(n3042), .B(n3041), .Z(n3043) );
  NAND U3664 ( .A(n3044), .B(n3043), .Z(n3046) );
  XNOR U3665 ( .A(n3047), .B(n3046), .Z(c[1608]) );
  NAND U3666 ( .A(b[0]), .B(a[586]), .Z(n3050) );
  XNOR U3667 ( .A(sreg[1609]), .B(n3050), .Z(n3052) );
  NANDN U3668 ( .A(sreg[1608]), .B(n3045), .Z(n3049) );
  NAND U3669 ( .A(n3047), .B(n3046), .Z(n3048) );
  NAND U3670 ( .A(n3049), .B(n3048), .Z(n3051) );
  XNOR U3671 ( .A(n3052), .B(n3051), .Z(c[1609]) );
  NAND U3672 ( .A(b[0]), .B(a[587]), .Z(n3055) );
  XNOR U3673 ( .A(sreg[1610]), .B(n3055), .Z(n3057) );
  NANDN U3674 ( .A(sreg[1609]), .B(n3050), .Z(n3054) );
  NAND U3675 ( .A(n3052), .B(n3051), .Z(n3053) );
  NAND U3676 ( .A(n3054), .B(n3053), .Z(n3056) );
  XNOR U3677 ( .A(n3057), .B(n3056), .Z(c[1610]) );
  NAND U3678 ( .A(b[0]), .B(a[588]), .Z(n3060) );
  XNOR U3679 ( .A(sreg[1611]), .B(n3060), .Z(n3062) );
  NANDN U3680 ( .A(sreg[1610]), .B(n3055), .Z(n3059) );
  NAND U3681 ( .A(n3057), .B(n3056), .Z(n3058) );
  NAND U3682 ( .A(n3059), .B(n3058), .Z(n3061) );
  XNOR U3683 ( .A(n3062), .B(n3061), .Z(c[1611]) );
  NAND U3684 ( .A(b[0]), .B(a[589]), .Z(n3065) );
  XNOR U3685 ( .A(sreg[1612]), .B(n3065), .Z(n3067) );
  NANDN U3686 ( .A(sreg[1611]), .B(n3060), .Z(n3064) );
  NAND U3687 ( .A(n3062), .B(n3061), .Z(n3063) );
  NAND U3688 ( .A(n3064), .B(n3063), .Z(n3066) );
  XNOR U3689 ( .A(n3067), .B(n3066), .Z(c[1612]) );
  NAND U3690 ( .A(b[0]), .B(a[590]), .Z(n3070) );
  XNOR U3691 ( .A(sreg[1613]), .B(n3070), .Z(n3072) );
  NANDN U3692 ( .A(sreg[1612]), .B(n3065), .Z(n3069) );
  NAND U3693 ( .A(n3067), .B(n3066), .Z(n3068) );
  NAND U3694 ( .A(n3069), .B(n3068), .Z(n3071) );
  XNOR U3695 ( .A(n3072), .B(n3071), .Z(c[1613]) );
  NAND U3696 ( .A(b[0]), .B(a[591]), .Z(n3075) );
  XNOR U3697 ( .A(sreg[1614]), .B(n3075), .Z(n3077) );
  NANDN U3698 ( .A(sreg[1613]), .B(n3070), .Z(n3074) );
  NAND U3699 ( .A(n3072), .B(n3071), .Z(n3073) );
  AND U3700 ( .A(n3074), .B(n3073), .Z(n3076) );
  XOR U3701 ( .A(n3077), .B(n3076), .Z(c[1614]) );
  NAND U3702 ( .A(b[0]), .B(a[592]), .Z(n3082) );
  NANDN U3703 ( .A(n3075), .B(sreg[1614]), .Z(n3079) );
  NAND U3704 ( .A(n3077), .B(n3076), .Z(n3078) );
  NAND U3705 ( .A(n3079), .B(n3078), .Z(n3081) );
  XOR U3706 ( .A(sreg[1615]), .B(n3081), .Z(n3080) );
  XNOR U3707 ( .A(n3082), .B(n3080), .Z(c[1615]) );
  NAND U3708 ( .A(b[0]), .B(a[593]), .Z(n3083) );
  XNOR U3709 ( .A(sreg[1616]), .B(n3083), .Z(n3084) );
  XOR U3710 ( .A(n3085), .B(n3084), .Z(c[1616]) );
  NAND U3711 ( .A(b[0]), .B(a[594]), .Z(n3088) );
  XNOR U3712 ( .A(sreg[1617]), .B(n3088), .Z(n3090) );
  NANDN U3713 ( .A(n3083), .B(sreg[1616]), .Z(n3087) );
  NAND U3714 ( .A(n3085), .B(n3084), .Z(n3086) );
  NAND U3715 ( .A(n3087), .B(n3086), .Z(n3089) );
  XOR U3716 ( .A(n3090), .B(n3089), .Z(c[1617]) );
  NAND U3717 ( .A(b[0]), .B(a[595]), .Z(n3093) );
  XNOR U3718 ( .A(sreg[1618]), .B(n3093), .Z(n3095) );
  NANDN U3719 ( .A(n3088), .B(sreg[1617]), .Z(n3092) );
  NAND U3720 ( .A(n3090), .B(n3089), .Z(n3091) );
  NAND U3721 ( .A(n3092), .B(n3091), .Z(n3094) );
  XOR U3722 ( .A(n3095), .B(n3094), .Z(c[1618]) );
  NAND U3723 ( .A(b[0]), .B(a[596]), .Z(n3098) );
  XNOR U3724 ( .A(sreg[1619]), .B(n3098), .Z(n3100) );
  NANDN U3725 ( .A(n3093), .B(sreg[1618]), .Z(n3097) );
  NAND U3726 ( .A(n3095), .B(n3094), .Z(n3096) );
  NAND U3727 ( .A(n3097), .B(n3096), .Z(n3099) );
  XOR U3728 ( .A(n3100), .B(n3099), .Z(c[1619]) );
  NAND U3729 ( .A(b[0]), .B(a[597]), .Z(n3103) );
  XNOR U3730 ( .A(sreg[1620]), .B(n3103), .Z(n3105) );
  NANDN U3731 ( .A(n3098), .B(sreg[1619]), .Z(n3102) );
  NAND U3732 ( .A(n3100), .B(n3099), .Z(n3101) );
  NAND U3733 ( .A(n3102), .B(n3101), .Z(n3104) );
  XOR U3734 ( .A(n3105), .B(n3104), .Z(c[1620]) );
  NAND U3735 ( .A(b[0]), .B(a[598]), .Z(n3108) );
  XNOR U3736 ( .A(sreg[1621]), .B(n3108), .Z(n3110) );
  NANDN U3737 ( .A(n3103), .B(sreg[1620]), .Z(n3107) );
  NAND U3738 ( .A(n3105), .B(n3104), .Z(n3106) );
  NAND U3739 ( .A(n3107), .B(n3106), .Z(n3109) );
  XOR U3740 ( .A(n3110), .B(n3109), .Z(c[1621]) );
  NAND U3741 ( .A(b[0]), .B(a[599]), .Z(n3113) );
  XNOR U3742 ( .A(sreg[1622]), .B(n3113), .Z(n3115) );
  NANDN U3743 ( .A(n3108), .B(sreg[1621]), .Z(n3112) );
  NAND U3744 ( .A(n3110), .B(n3109), .Z(n3111) );
  NAND U3745 ( .A(n3112), .B(n3111), .Z(n3114) );
  XOR U3746 ( .A(n3115), .B(n3114), .Z(c[1622]) );
  NAND U3747 ( .A(b[0]), .B(a[600]), .Z(n3118) );
  XNOR U3748 ( .A(sreg[1623]), .B(n3118), .Z(n3120) );
  NANDN U3749 ( .A(n3113), .B(sreg[1622]), .Z(n3117) );
  NAND U3750 ( .A(n3115), .B(n3114), .Z(n3116) );
  NAND U3751 ( .A(n3117), .B(n3116), .Z(n3119) );
  XOR U3752 ( .A(n3120), .B(n3119), .Z(c[1623]) );
  NAND U3753 ( .A(b[0]), .B(a[601]), .Z(n3123) );
  XNOR U3754 ( .A(sreg[1624]), .B(n3123), .Z(n3125) );
  NANDN U3755 ( .A(n3118), .B(sreg[1623]), .Z(n3122) );
  NAND U3756 ( .A(n3120), .B(n3119), .Z(n3121) );
  AND U3757 ( .A(n3122), .B(n3121), .Z(n3124) );
  XNOR U3758 ( .A(n3125), .B(n3124), .Z(c[1624]) );
  NAND U3759 ( .A(b[0]), .B(a[602]), .Z(n3128) );
  XNOR U3760 ( .A(sreg[1625]), .B(n3128), .Z(n3130) );
  NANDN U3761 ( .A(sreg[1624]), .B(n3123), .Z(n3127) );
  NAND U3762 ( .A(n3125), .B(n3124), .Z(n3126) );
  AND U3763 ( .A(n3127), .B(n3126), .Z(n3129) );
  XOR U3764 ( .A(n3130), .B(n3129), .Z(c[1625]) );
  NAND U3765 ( .A(b[0]), .B(a[603]), .Z(n3133) );
  XNOR U3766 ( .A(sreg[1626]), .B(n3133), .Z(n3135) );
  NANDN U3767 ( .A(n3128), .B(sreg[1625]), .Z(n3132) );
  NAND U3768 ( .A(n3130), .B(n3129), .Z(n3131) );
  NAND U3769 ( .A(n3132), .B(n3131), .Z(n3134) );
  XOR U3770 ( .A(n3135), .B(n3134), .Z(c[1626]) );
  NANDN U3771 ( .A(n3133), .B(sreg[1626]), .Z(n3137) );
  NAND U3772 ( .A(n3135), .B(n3134), .Z(n3136) );
  AND U3773 ( .A(n3137), .B(n3136), .Z(n3140) );
  NAND U3774 ( .A(b[0]), .B(a[604]), .Z(n3138) );
  XNOR U3775 ( .A(sreg[1627]), .B(n3138), .Z(n3139) );
  XNOR U3776 ( .A(n3140), .B(n3139), .Z(c[1627]) );
  NAND U3777 ( .A(b[0]), .B(a[605]), .Z(n3143) );
  XNOR U3778 ( .A(sreg[1628]), .B(n3143), .Z(n3145) );
  NANDN U3779 ( .A(sreg[1627]), .B(n3138), .Z(n3142) );
  NAND U3780 ( .A(n3140), .B(n3139), .Z(n3141) );
  AND U3781 ( .A(n3142), .B(n3141), .Z(n3144) );
  XOR U3782 ( .A(n3145), .B(n3144), .Z(c[1628]) );
  NAND U3783 ( .A(b[0]), .B(a[606]), .Z(n3148) );
  XNOR U3784 ( .A(sreg[1629]), .B(n3148), .Z(n3150) );
  NANDN U3785 ( .A(n3143), .B(sreg[1628]), .Z(n3147) );
  NAND U3786 ( .A(n3145), .B(n3144), .Z(n3146) );
  NAND U3787 ( .A(n3147), .B(n3146), .Z(n3149) );
  XOR U3788 ( .A(n3150), .B(n3149), .Z(c[1629]) );
  NAND U3789 ( .A(b[0]), .B(a[607]), .Z(n3153) );
  XNOR U3790 ( .A(sreg[1630]), .B(n3153), .Z(n3155) );
  NANDN U3791 ( .A(n3148), .B(sreg[1629]), .Z(n3152) );
  NAND U3792 ( .A(n3150), .B(n3149), .Z(n3151) );
  NAND U3793 ( .A(n3152), .B(n3151), .Z(n3154) );
  XOR U3794 ( .A(n3155), .B(n3154), .Z(c[1630]) );
  NAND U3795 ( .A(b[0]), .B(a[608]), .Z(n3158) );
  XNOR U3796 ( .A(sreg[1631]), .B(n3158), .Z(n3160) );
  NANDN U3797 ( .A(n3153), .B(sreg[1630]), .Z(n3157) );
  NAND U3798 ( .A(n3155), .B(n3154), .Z(n3156) );
  NAND U3799 ( .A(n3157), .B(n3156), .Z(n3159) );
  XOR U3800 ( .A(n3160), .B(n3159), .Z(c[1631]) );
  NAND U3801 ( .A(b[0]), .B(a[609]), .Z(n3163) );
  XNOR U3802 ( .A(sreg[1632]), .B(n3163), .Z(n3165) );
  NANDN U3803 ( .A(n3158), .B(sreg[1631]), .Z(n3162) );
  NAND U3804 ( .A(n3160), .B(n3159), .Z(n3161) );
  NAND U3805 ( .A(n3162), .B(n3161), .Z(n3164) );
  XOR U3806 ( .A(n3165), .B(n3164), .Z(c[1632]) );
  NAND U3807 ( .A(b[0]), .B(a[610]), .Z(n3168) );
  XNOR U3808 ( .A(sreg[1633]), .B(n3168), .Z(n3170) );
  NANDN U3809 ( .A(n3163), .B(sreg[1632]), .Z(n3167) );
  NAND U3810 ( .A(n3165), .B(n3164), .Z(n3166) );
  NAND U3811 ( .A(n3167), .B(n3166), .Z(n3169) );
  XOR U3812 ( .A(n3170), .B(n3169), .Z(c[1633]) );
  NAND U3813 ( .A(b[0]), .B(a[611]), .Z(n3173) );
  XNOR U3814 ( .A(sreg[1634]), .B(n3173), .Z(n3175) );
  NANDN U3815 ( .A(n3168), .B(sreg[1633]), .Z(n3172) );
  NAND U3816 ( .A(n3170), .B(n3169), .Z(n3171) );
  NAND U3817 ( .A(n3172), .B(n3171), .Z(n3174) );
  XOR U3818 ( .A(n3175), .B(n3174), .Z(c[1634]) );
  NAND U3819 ( .A(b[0]), .B(a[612]), .Z(n3178) );
  XNOR U3820 ( .A(sreg[1635]), .B(n3178), .Z(n3180) );
  NANDN U3821 ( .A(n3173), .B(sreg[1634]), .Z(n3177) );
  NAND U3822 ( .A(n3175), .B(n3174), .Z(n3176) );
  NAND U3823 ( .A(n3177), .B(n3176), .Z(n3179) );
  XOR U3824 ( .A(n3180), .B(n3179), .Z(c[1635]) );
  NAND U3825 ( .A(b[0]), .B(a[613]), .Z(n3183) );
  XNOR U3826 ( .A(sreg[1636]), .B(n3183), .Z(n3185) );
  NANDN U3827 ( .A(n3178), .B(sreg[1635]), .Z(n3182) );
  NAND U3828 ( .A(n3180), .B(n3179), .Z(n3181) );
  NAND U3829 ( .A(n3182), .B(n3181), .Z(n3184) );
  XOR U3830 ( .A(n3185), .B(n3184), .Z(c[1636]) );
  NAND U3831 ( .A(b[0]), .B(a[614]), .Z(n3188) );
  XNOR U3832 ( .A(sreg[1637]), .B(n3188), .Z(n3190) );
  NANDN U3833 ( .A(n3183), .B(sreg[1636]), .Z(n3187) );
  NAND U3834 ( .A(n3185), .B(n3184), .Z(n3186) );
  NAND U3835 ( .A(n3187), .B(n3186), .Z(n3189) );
  XOR U3836 ( .A(n3190), .B(n3189), .Z(c[1637]) );
  NAND U3837 ( .A(b[0]), .B(a[615]), .Z(n3193) );
  XNOR U3838 ( .A(sreg[1638]), .B(n3193), .Z(n3195) );
  NANDN U3839 ( .A(n3188), .B(sreg[1637]), .Z(n3192) );
  NAND U3840 ( .A(n3190), .B(n3189), .Z(n3191) );
  NAND U3841 ( .A(n3192), .B(n3191), .Z(n3194) );
  XOR U3842 ( .A(n3195), .B(n3194), .Z(c[1638]) );
  NAND U3843 ( .A(b[0]), .B(a[616]), .Z(n3198) );
  XNOR U3844 ( .A(sreg[1639]), .B(n3198), .Z(n3200) );
  NANDN U3845 ( .A(n3193), .B(sreg[1638]), .Z(n3197) );
  NAND U3846 ( .A(n3195), .B(n3194), .Z(n3196) );
  NAND U3847 ( .A(n3197), .B(n3196), .Z(n3199) );
  XOR U3848 ( .A(n3200), .B(n3199), .Z(c[1639]) );
  NAND U3849 ( .A(b[0]), .B(a[617]), .Z(n3203) );
  XNOR U3850 ( .A(sreg[1640]), .B(n3203), .Z(n3205) );
  NANDN U3851 ( .A(n3198), .B(sreg[1639]), .Z(n3202) );
  NAND U3852 ( .A(n3200), .B(n3199), .Z(n3201) );
  NAND U3853 ( .A(n3202), .B(n3201), .Z(n3204) );
  XOR U3854 ( .A(n3205), .B(n3204), .Z(c[1640]) );
  NAND U3855 ( .A(b[0]), .B(a[618]), .Z(n3208) );
  XNOR U3856 ( .A(sreg[1641]), .B(n3208), .Z(n3210) );
  NANDN U3857 ( .A(n3203), .B(sreg[1640]), .Z(n3207) );
  NAND U3858 ( .A(n3205), .B(n3204), .Z(n3206) );
  NAND U3859 ( .A(n3207), .B(n3206), .Z(n3209) );
  XOR U3860 ( .A(n3210), .B(n3209), .Z(c[1641]) );
  NAND U3861 ( .A(b[0]), .B(a[619]), .Z(n3213) );
  XNOR U3862 ( .A(sreg[1642]), .B(n3213), .Z(n3215) );
  NANDN U3863 ( .A(n3208), .B(sreg[1641]), .Z(n3212) );
  NAND U3864 ( .A(n3210), .B(n3209), .Z(n3211) );
  NAND U3865 ( .A(n3212), .B(n3211), .Z(n3214) );
  XOR U3866 ( .A(n3215), .B(n3214), .Z(c[1642]) );
  NAND U3867 ( .A(b[0]), .B(a[620]), .Z(n3218) );
  XNOR U3868 ( .A(sreg[1643]), .B(n3218), .Z(n3220) );
  NANDN U3869 ( .A(n3213), .B(sreg[1642]), .Z(n3217) );
  NAND U3870 ( .A(n3215), .B(n3214), .Z(n3216) );
  NAND U3871 ( .A(n3217), .B(n3216), .Z(n3219) );
  XOR U3872 ( .A(n3220), .B(n3219), .Z(c[1643]) );
  NAND U3873 ( .A(b[0]), .B(a[621]), .Z(n3223) );
  XNOR U3874 ( .A(sreg[1644]), .B(n3223), .Z(n3225) );
  NANDN U3875 ( .A(n3218), .B(sreg[1643]), .Z(n3222) );
  NAND U3876 ( .A(n3220), .B(n3219), .Z(n3221) );
  NAND U3877 ( .A(n3222), .B(n3221), .Z(n3224) );
  XOR U3878 ( .A(n3225), .B(n3224), .Z(c[1644]) );
  NANDN U3879 ( .A(n3223), .B(sreg[1644]), .Z(n3227) );
  NAND U3880 ( .A(n3225), .B(n3224), .Z(n3226) );
  AND U3881 ( .A(n3227), .B(n3226), .Z(n3230) );
  NAND U3882 ( .A(b[0]), .B(a[622]), .Z(n3228) );
  XNOR U3883 ( .A(sreg[1645]), .B(n3228), .Z(n3229) );
  XNOR U3884 ( .A(n3230), .B(n3229), .Z(c[1645]) );
  NAND U3885 ( .A(b[0]), .B(a[623]), .Z(n3233) );
  XNOR U3886 ( .A(sreg[1646]), .B(n3233), .Z(n3235) );
  NANDN U3887 ( .A(sreg[1645]), .B(n3228), .Z(n3232) );
  NAND U3888 ( .A(n3230), .B(n3229), .Z(n3231) );
  NAND U3889 ( .A(n3232), .B(n3231), .Z(n3234) );
  XNOR U3890 ( .A(n3235), .B(n3234), .Z(c[1646]) );
  NAND U3891 ( .A(b[0]), .B(a[624]), .Z(n3238) );
  XNOR U3892 ( .A(sreg[1647]), .B(n3238), .Z(n3240) );
  NANDN U3893 ( .A(sreg[1646]), .B(n3233), .Z(n3237) );
  NAND U3894 ( .A(n3235), .B(n3234), .Z(n3236) );
  NAND U3895 ( .A(n3237), .B(n3236), .Z(n3239) );
  XNOR U3896 ( .A(n3240), .B(n3239), .Z(c[1647]) );
  NAND U3897 ( .A(b[0]), .B(a[625]), .Z(n3243) );
  XNOR U3898 ( .A(sreg[1648]), .B(n3243), .Z(n3245) );
  NANDN U3899 ( .A(sreg[1647]), .B(n3238), .Z(n3242) );
  NAND U3900 ( .A(n3240), .B(n3239), .Z(n3241) );
  NAND U3901 ( .A(n3242), .B(n3241), .Z(n3244) );
  XNOR U3902 ( .A(n3245), .B(n3244), .Z(c[1648]) );
  NAND U3903 ( .A(b[0]), .B(a[626]), .Z(n3248) );
  XNOR U3904 ( .A(sreg[1649]), .B(n3248), .Z(n3250) );
  NANDN U3905 ( .A(sreg[1648]), .B(n3243), .Z(n3247) );
  NAND U3906 ( .A(n3245), .B(n3244), .Z(n3246) );
  NAND U3907 ( .A(n3247), .B(n3246), .Z(n3249) );
  XNOR U3908 ( .A(n3250), .B(n3249), .Z(c[1649]) );
  NAND U3909 ( .A(b[0]), .B(a[627]), .Z(n3253) );
  XNOR U3910 ( .A(sreg[1650]), .B(n3253), .Z(n3255) );
  NANDN U3911 ( .A(sreg[1649]), .B(n3248), .Z(n3252) );
  NAND U3912 ( .A(n3250), .B(n3249), .Z(n3251) );
  NAND U3913 ( .A(n3252), .B(n3251), .Z(n3254) );
  XNOR U3914 ( .A(n3255), .B(n3254), .Z(c[1650]) );
  NANDN U3915 ( .A(sreg[1650]), .B(n3253), .Z(n3257) );
  NAND U3916 ( .A(n3255), .B(n3254), .Z(n3256) );
  AND U3917 ( .A(n3257), .B(n3256), .Z(n3260) );
  NAND U3918 ( .A(b[0]), .B(a[628]), .Z(n3258) );
  XNOR U3919 ( .A(sreg[1651]), .B(n3258), .Z(n3259) );
  XOR U3920 ( .A(n3260), .B(n3259), .Z(c[1651]) );
  NAND U3921 ( .A(b[0]), .B(a[629]), .Z(n3263) );
  XNOR U3922 ( .A(sreg[1652]), .B(n3263), .Z(n3265) );
  NANDN U3923 ( .A(n3258), .B(sreg[1651]), .Z(n3262) );
  NAND U3924 ( .A(n3260), .B(n3259), .Z(n3261) );
  AND U3925 ( .A(n3262), .B(n3261), .Z(n3264) );
  XNOR U3926 ( .A(n3265), .B(n3264), .Z(c[1652]) );
  NANDN U3927 ( .A(sreg[1652]), .B(n3263), .Z(n3267) );
  NAND U3928 ( .A(n3265), .B(n3264), .Z(n3266) );
  AND U3929 ( .A(n3267), .B(n3266), .Z(n3270) );
  NAND U3930 ( .A(b[0]), .B(a[630]), .Z(n3268) );
  XNOR U3931 ( .A(sreg[1653]), .B(n3268), .Z(n3269) );
  XOR U3932 ( .A(n3270), .B(n3269), .Z(c[1653]) );
  NAND U3933 ( .A(b[0]), .B(a[631]), .Z(n3273) );
  XNOR U3934 ( .A(sreg[1654]), .B(n3273), .Z(n3275) );
  NANDN U3935 ( .A(n3268), .B(sreg[1653]), .Z(n3272) );
  NAND U3936 ( .A(n3270), .B(n3269), .Z(n3271) );
  NAND U3937 ( .A(n3272), .B(n3271), .Z(n3274) );
  XOR U3938 ( .A(n3275), .B(n3274), .Z(c[1654]) );
  NAND U3939 ( .A(b[0]), .B(a[632]), .Z(n3278) );
  XNOR U3940 ( .A(sreg[1655]), .B(n3278), .Z(n3280) );
  NANDN U3941 ( .A(n3273), .B(sreg[1654]), .Z(n3277) );
  NAND U3942 ( .A(n3275), .B(n3274), .Z(n3276) );
  AND U3943 ( .A(n3277), .B(n3276), .Z(n3279) );
  XNOR U3944 ( .A(n3280), .B(n3279), .Z(c[1655]) );
  NANDN U3945 ( .A(sreg[1655]), .B(n3278), .Z(n3282) );
  NAND U3946 ( .A(n3280), .B(n3279), .Z(n3281) );
  AND U3947 ( .A(n3282), .B(n3281), .Z(n3285) );
  NAND U3948 ( .A(b[0]), .B(a[633]), .Z(n3283) );
  XNOR U3949 ( .A(sreg[1656]), .B(n3283), .Z(n3284) );
  XOR U3950 ( .A(n3285), .B(n3284), .Z(c[1656]) );
  NAND U3951 ( .A(b[0]), .B(a[634]), .Z(n3288) );
  XNOR U3952 ( .A(sreg[1657]), .B(n3288), .Z(n3290) );
  NANDN U3953 ( .A(n3283), .B(sreg[1656]), .Z(n3287) );
  NAND U3954 ( .A(n3285), .B(n3284), .Z(n3286) );
  NAND U3955 ( .A(n3287), .B(n3286), .Z(n3289) );
  XOR U3956 ( .A(n3290), .B(n3289), .Z(c[1657]) );
  NAND U3957 ( .A(b[0]), .B(a[635]), .Z(n3295) );
  NANDN U3958 ( .A(n3288), .B(sreg[1657]), .Z(n3292) );
  NAND U3959 ( .A(n3290), .B(n3289), .Z(n3291) );
  NAND U3960 ( .A(n3292), .B(n3291), .Z(n3294) );
  XOR U3961 ( .A(sreg[1658]), .B(n3294), .Z(n3293) );
  XNOR U3962 ( .A(n3295), .B(n3293), .Z(c[1658]) );
  NAND U3963 ( .A(b[0]), .B(a[636]), .Z(n3296) );
  XNOR U3964 ( .A(sreg[1659]), .B(n3296), .Z(n3297) );
  XOR U3965 ( .A(n3298), .B(n3297), .Z(c[1659]) );
  NAND U3966 ( .A(b[0]), .B(a[637]), .Z(n3301) );
  XNOR U3967 ( .A(sreg[1660]), .B(n3301), .Z(n3303) );
  NANDN U3968 ( .A(n3296), .B(sreg[1659]), .Z(n3300) );
  NAND U3969 ( .A(n3298), .B(n3297), .Z(n3299) );
  NAND U3970 ( .A(n3300), .B(n3299), .Z(n3302) );
  XOR U3971 ( .A(n3303), .B(n3302), .Z(c[1660]) );
  NANDN U3972 ( .A(n3301), .B(sreg[1660]), .Z(n3305) );
  NAND U3973 ( .A(n3303), .B(n3302), .Z(n3304) );
  AND U3974 ( .A(n3305), .B(n3304), .Z(n3308) );
  NAND U3975 ( .A(b[0]), .B(a[638]), .Z(n3306) );
  XNOR U3976 ( .A(sreg[1661]), .B(n3306), .Z(n3307) );
  XNOR U3977 ( .A(n3308), .B(n3307), .Z(c[1661]) );
  NAND U3978 ( .A(b[0]), .B(a[639]), .Z(n3311) );
  XNOR U3979 ( .A(sreg[1662]), .B(n3311), .Z(n3313) );
  NANDN U3980 ( .A(sreg[1661]), .B(n3306), .Z(n3310) );
  NAND U3981 ( .A(n3308), .B(n3307), .Z(n3309) );
  AND U3982 ( .A(n3310), .B(n3309), .Z(n3312) );
  XOR U3983 ( .A(n3313), .B(n3312), .Z(c[1662]) );
  NAND U3984 ( .A(b[0]), .B(a[640]), .Z(n3316) );
  XNOR U3985 ( .A(sreg[1663]), .B(n3316), .Z(n3318) );
  NANDN U3986 ( .A(n3311), .B(sreg[1662]), .Z(n3315) );
  NAND U3987 ( .A(n3313), .B(n3312), .Z(n3314) );
  NAND U3988 ( .A(n3315), .B(n3314), .Z(n3317) );
  XOR U3989 ( .A(n3318), .B(n3317), .Z(c[1663]) );
  NANDN U3990 ( .A(n3316), .B(sreg[1663]), .Z(n3320) );
  NAND U3991 ( .A(n3318), .B(n3317), .Z(n3319) );
  AND U3992 ( .A(n3320), .B(n3319), .Z(n3323) );
  NAND U3993 ( .A(b[0]), .B(a[641]), .Z(n3321) );
  XNOR U3994 ( .A(sreg[1664]), .B(n3321), .Z(n3322) );
  XNOR U3995 ( .A(n3323), .B(n3322), .Z(c[1664]) );
  NANDN U3996 ( .A(sreg[1664]), .B(n3321), .Z(n3325) );
  NAND U3997 ( .A(n3323), .B(n3322), .Z(n3324) );
  AND U3998 ( .A(n3325), .B(n3324), .Z(n3328) );
  NAND U3999 ( .A(b[0]), .B(a[642]), .Z(n3326) );
  XNOR U4000 ( .A(sreg[1665]), .B(n3326), .Z(n3327) );
  XOR U4001 ( .A(n3328), .B(n3327), .Z(c[1665]) );
  NAND U4002 ( .A(b[0]), .B(a[643]), .Z(n3331) );
  XNOR U4003 ( .A(sreg[1666]), .B(n3331), .Z(n3333) );
  NANDN U4004 ( .A(n3326), .B(sreg[1665]), .Z(n3330) );
  NAND U4005 ( .A(n3328), .B(n3327), .Z(n3329) );
  NAND U4006 ( .A(n3330), .B(n3329), .Z(n3332) );
  XOR U4007 ( .A(n3333), .B(n3332), .Z(c[1666]) );
  NANDN U4008 ( .A(n3331), .B(sreg[1666]), .Z(n3335) );
  NAND U4009 ( .A(n3333), .B(n3332), .Z(n3334) );
  AND U4010 ( .A(n3335), .B(n3334), .Z(n3338) );
  NAND U4011 ( .A(b[0]), .B(a[644]), .Z(n3336) );
  XNOR U4012 ( .A(sreg[1667]), .B(n3336), .Z(n3337) );
  XNOR U4013 ( .A(n3338), .B(n3337), .Z(c[1667]) );
  NANDN U4014 ( .A(sreg[1667]), .B(n3336), .Z(n3340) );
  NAND U4015 ( .A(n3338), .B(n3337), .Z(n3339) );
  AND U4016 ( .A(n3340), .B(n3339), .Z(n3343) );
  NAND U4017 ( .A(b[0]), .B(a[645]), .Z(n3341) );
  XNOR U4018 ( .A(sreg[1668]), .B(n3341), .Z(n3342) );
  XOR U4019 ( .A(n3343), .B(n3342), .Z(c[1668]) );
  NANDN U4020 ( .A(n3341), .B(sreg[1668]), .Z(n3345) );
  NAND U4021 ( .A(n3343), .B(n3342), .Z(n3344) );
  AND U4022 ( .A(n3345), .B(n3344), .Z(n3348) );
  NAND U4023 ( .A(b[0]), .B(a[646]), .Z(n3346) );
  XNOR U4024 ( .A(sreg[1669]), .B(n3346), .Z(n3347) );
  XNOR U4025 ( .A(n3348), .B(n3347), .Z(c[1669]) );
  NANDN U4026 ( .A(sreg[1669]), .B(n3346), .Z(n3350) );
  NAND U4027 ( .A(n3348), .B(n3347), .Z(n3349) );
  AND U4028 ( .A(n3350), .B(n3349), .Z(n3353) );
  NAND U4029 ( .A(b[0]), .B(a[647]), .Z(n3351) );
  XNOR U4030 ( .A(sreg[1670]), .B(n3351), .Z(n3352) );
  XOR U4031 ( .A(n3353), .B(n3352), .Z(c[1670]) );
  NAND U4032 ( .A(b[0]), .B(a[648]), .Z(n3356) );
  XNOR U4033 ( .A(sreg[1671]), .B(n3356), .Z(n3358) );
  NANDN U4034 ( .A(n3351), .B(sreg[1670]), .Z(n3355) );
  NAND U4035 ( .A(n3353), .B(n3352), .Z(n3354) );
  AND U4036 ( .A(n3355), .B(n3354), .Z(n3357) );
  XNOR U4037 ( .A(n3358), .B(n3357), .Z(c[1671]) );
  NAND U4038 ( .A(b[0]), .B(a[649]), .Z(n3361) );
  XNOR U4039 ( .A(sreg[1672]), .B(n3361), .Z(n3363) );
  NANDN U4040 ( .A(sreg[1671]), .B(n3356), .Z(n3360) );
  NAND U4041 ( .A(n3358), .B(n3357), .Z(n3359) );
  NAND U4042 ( .A(n3360), .B(n3359), .Z(n3362) );
  XNOR U4043 ( .A(n3363), .B(n3362), .Z(c[1672]) );
  NAND U4044 ( .A(b[0]), .B(a[650]), .Z(n3366) );
  XNOR U4045 ( .A(sreg[1673]), .B(n3366), .Z(n3368) );
  NANDN U4046 ( .A(sreg[1672]), .B(n3361), .Z(n3365) );
  NAND U4047 ( .A(n3363), .B(n3362), .Z(n3364) );
  AND U4048 ( .A(n3365), .B(n3364), .Z(n3367) );
  XOR U4049 ( .A(n3368), .B(n3367), .Z(c[1673]) );
  NAND U4050 ( .A(b[0]), .B(a[651]), .Z(n3371) );
  XNOR U4051 ( .A(sreg[1674]), .B(n3371), .Z(n3373) );
  NANDN U4052 ( .A(n3366), .B(sreg[1673]), .Z(n3370) );
  NAND U4053 ( .A(n3368), .B(n3367), .Z(n3369) );
  AND U4054 ( .A(n3370), .B(n3369), .Z(n3372) );
  XNOR U4055 ( .A(n3373), .B(n3372), .Z(c[1674]) );
  NAND U4056 ( .A(b[0]), .B(a[652]), .Z(n3376) );
  XNOR U4057 ( .A(sreg[1675]), .B(n3376), .Z(n3378) );
  NANDN U4058 ( .A(sreg[1674]), .B(n3371), .Z(n3375) );
  NAND U4059 ( .A(n3373), .B(n3372), .Z(n3374) );
  NAND U4060 ( .A(n3375), .B(n3374), .Z(n3377) );
  XNOR U4061 ( .A(n3378), .B(n3377), .Z(c[1675]) );
  NAND U4062 ( .A(b[0]), .B(a[653]), .Z(n3381) );
  XNOR U4063 ( .A(sreg[1676]), .B(n3381), .Z(n3383) );
  NANDN U4064 ( .A(sreg[1675]), .B(n3376), .Z(n3380) );
  NAND U4065 ( .A(n3378), .B(n3377), .Z(n3379) );
  AND U4066 ( .A(n3380), .B(n3379), .Z(n3382) );
  XOR U4067 ( .A(n3383), .B(n3382), .Z(c[1676]) );
  NANDN U4068 ( .A(n3381), .B(sreg[1676]), .Z(n3385) );
  NAND U4069 ( .A(n3383), .B(n3382), .Z(n3384) );
  AND U4070 ( .A(n3385), .B(n3384), .Z(n3388) );
  NAND U4071 ( .A(b[0]), .B(a[654]), .Z(n3386) );
  XNOR U4072 ( .A(sreg[1677]), .B(n3386), .Z(n3387) );
  XNOR U4073 ( .A(n3388), .B(n3387), .Z(c[1677]) );
  NAND U4074 ( .A(b[0]), .B(a[655]), .Z(n3391) );
  XNOR U4075 ( .A(sreg[1678]), .B(n3391), .Z(n3393) );
  NANDN U4076 ( .A(sreg[1677]), .B(n3386), .Z(n3390) );
  NAND U4077 ( .A(n3388), .B(n3387), .Z(n3389) );
  NAND U4078 ( .A(n3390), .B(n3389), .Z(n3392) );
  XNOR U4079 ( .A(n3393), .B(n3392), .Z(c[1678]) );
  NANDN U4080 ( .A(sreg[1678]), .B(n3391), .Z(n3395) );
  NAND U4081 ( .A(n3393), .B(n3392), .Z(n3394) );
  AND U4082 ( .A(n3395), .B(n3394), .Z(n3398) );
  NAND U4083 ( .A(b[0]), .B(a[656]), .Z(n3397) );
  XOR U4084 ( .A(sreg[1679]), .B(n3397), .Z(n3396) );
  XNOR U4085 ( .A(n3398), .B(n3396), .Z(c[1679]) );
  AND U4086 ( .A(b[0]), .B(a[657]), .Z(n3401) );
  IV U4087 ( .A(n3401), .Z(n3400) );
  XOR U4088 ( .A(n3400), .B(sreg[1680]), .Z(n3399) );
  XNOR U4089 ( .A(n3402), .B(n3399), .Z(c[1680]) );
  NANDN U4090 ( .A(n3400), .B(sreg[1680]), .Z(n3405) );
  NOR U4091 ( .A(n3401), .B(sreg[1680]), .Z(n3403) );
  NANDN U4092 ( .A(n3403), .B(n3402), .Z(n3404) );
  AND U4093 ( .A(n3405), .B(n3404), .Z(n3408) );
  NAND U4094 ( .A(b[0]), .B(a[658]), .Z(n3406) );
  XNOR U4095 ( .A(sreg[1681]), .B(n3406), .Z(n3407) );
  XNOR U4096 ( .A(n3408), .B(n3407), .Z(c[1681]) );
  NAND U4097 ( .A(b[0]), .B(a[659]), .Z(n3411) );
  XNOR U4098 ( .A(sreg[1682]), .B(n3411), .Z(n3413) );
  NANDN U4099 ( .A(n3406), .B(sreg[1681]), .Z(n3410) );
  NANDN U4100 ( .A(n3408), .B(n3407), .Z(n3409) );
  AND U4101 ( .A(n3410), .B(n3409), .Z(n3412) );
  XNOR U4102 ( .A(n3413), .B(n3412), .Z(c[1682]) );
  NANDN U4103 ( .A(sreg[1682]), .B(n3411), .Z(n3415) );
  NAND U4104 ( .A(n3413), .B(n3412), .Z(n3414) );
  AND U4105 ( .A(n3415), .B(n3414), .Z(n3418) );
  NAND U4106 ( .A(b[0]), .B(a[660]), .Z(n3416) );
  XNOR U4107 ( .A(sreg[1683]), .B(n3416), .Z(n3417) );
  XOR U4108 ( .A(n3418), .B(n3417), .Z(c[1683]) );
  NAND U4109 ( .A(b[0]), .B(a[661]), .Z(n3421) );
  XNOR U4110 ( .A(sreg[1684]), .B(n3421), .Z(n3423) );
  NANDN U4111 ( .A(n3416), .B(sreg[1683]), .Z(n3420) );
  NAND U4112 ( .A(n3418), .B(n3417), .Z(n3419) );
  NAND U4113 ( .A(n3420), .B(n3419), .Z(n3422) );
  XOR U4114 ( .A(n3423), .B(n3422), .Z(c[1684]) );
  NAND U4115 ( .A(b[0]), .B(a[662]), .Z(n3426) );
  XNOR U4116 ( .A(sreg[1685]), .B(n3426), .Z(n3428) );
  NANDN U4117 ( .A(n3421), .B(sreg[1684]), .Z(n3425) );
  NAND U4118 ( .A(n3423), .B(n3422), .Z(n3424) );
  AND U4119 ( .A(n3425), .B(n3424), .Z(n3427) );
  XNOR U4120 ( .A(n3428), .B(n3427), .Z(c[1685]) );
  NANDN U4121 ( .A(sreg[1685]), .B(n3426), .Z(n3430) );
  NAND U4122 ( .A(n3428), .B(n3427), .Z(n3429) );
  AND U4123 ( .A(n3430), .B(n3429), .Z(n3433) );
  NAND U4124 ( .A(b[0]), .B(a[663]), .Z(n3431) );
  XNOR U4125 ( .A(sreg[1686]), .B(n3431), .Z(n3432) );
  XOR U4126 ( .A(n3433), .B(n3432), .Z(c[1686]) );
  NAND U4127 ( .A(b[0]), .B(a[664]), .Z(n3436) );
  XNOR U4128 ( .A(sreg[1687]), .B(n3436), .Z(n3438) );
  NANDN U4129 ( .A(n3431), .B(sreg[1686]), .Z(n3435) );
  NAND U4130 ( .A(n3433), .B(n3432), .Z(n3434) );
  NAND U4131 ( .A(n3435), .B(n3434), .Z(n3437) );
  XOR U4132 ( .A(n3438), .B(n3437), .Z(c[1687]) );
  NAND U4133 ( .A(b[0]), .B(a[665]), .Z(n3441) );
  XNOR U4134 ( .A(sreg[1688]), .B(n3441), .Z(n3443) );
  NANDN U4135 ( .A(n3436), .B(sreg[1687]), .Z(n3440) );
  NAND U4136 ( .A(n3438), .B(n3437), .Z(n3439) );
  AND U4137 ( .A(n3440), .B(n3439), .Z(n3442) );
  XNOR U4138 ( .A(n3443), .B(n3442), .Z(c[1688]) );
  NANDN U4139 ( .A(sreg[1688]), .B(n3441), .Z(n3445) );
  NAND U4140 ( .A(n3443), .B(n3442), .Z(n3444) );
  AND U4141 ( .A(n3445), .B(n3444), .Z(n3448) );
  NAND U4142 ( .A(b[0]), .B(a[666]), .Z(n3446) );
  XNOR U4143 ( .A(sreg[1689]), .B(n3446), .Z(n3447) );
  XOR U4144 ( .A(n3448), .B(n3447), .Z(c[1689]) );
  NAND U4145 ( .A(b[0]), .B(a[667]), .Z(n3451) );
  XNOR U4146 ( .A(sreg[1690]), .B(n3451), .Z(n3453) );
  NANDN U4147 ( .A(n3446), .B(sreg[1689]), .Z(n3450) );
  NAND U4148 ( .A(n3448), .B(n3447), .Z(n3449) );
  NAND U4149 ( .A(n3450), .B(n3449), .Z(n3452) );
  XOR U4150 ( .A(n3453), .B(n3452), .Z(c[1690]) );
  NAND U4151 ( .A(b[0]), .B(a[668]), .Z(n3456) );
  XNOR U4152 ( .A(sreg[1691]), .B(n3456), .Z(n3458) );
  NANDN U4153 ( .A(n3451), .B(sreg[1690]), .Z(n3455) );
  NAND U4154 ( .A(n3453), .B(n3452), .Z(n3454) );
  AND U4155 ( .A(n3455), .B(n3454), .Z(n3457) );
  XNOR U4156 ( .A(n3458), .B(n3457), .Z(c[1691]) );
  NAND U4157 ( .A(b[0]), .B(a[669]), .Z(n3461) );
  XNOR U4158 ( .A(sreg[1692]), .B(n3461), .Z(n3463) );
  NANDN U4159 ( .A(sreg[1691]), .B(n3456), .Z(n3460) );
  NAND U4160 ( .A(n3458), .B(n3457), .Z(n3459) );
  NAND U4161 ( .A(n3460), .B(n3459), .Z(n3462) );
  XNOR U4162 ( .A(n3463), .B(n3462), .Z(c[1692]) );
  NAND U4163 ( .A(b[0]), .B(a[670]), .Z(n3466) );
  XNOR U4164 ( .A(sreg[1693]), .B(n3466), .Z(n3468) );
  NANDN U4165 ( .A(sreg[1692]), .B(n3461), .Z(n3465) );
  NAND U4166 ( .A(n3463), .B(n3462), .Z(n3464) );
  NAND U4167 ( .A(n3465), .B(n3464), .Z(n3467) );
  XNOR U4168 ( .A(n3468), .B(n3467), .Z(c[1693]) );
  NAND U4169 ( .A(b[0]), .B(a[671]), .Z(n3471) );
  XNOR U4170 ( .A(sreg[1694]), .B(n3471), .Z(n3473) );
  NANDN U4171 ( .A(sreg[1693]), .B(n3466), .Z(n3470) );
  NAND U4172 ( .A(n3468), .B(n3467), .Z(n3469) );
  NAND U4173 ( .A(n3470), .B(n3469), .Z(n3472) );
  XNOR U4174 ( .A(n3473), .B(n3472), .Z(c[1694]) );
  NAND U4175 ( .A(b[0]), .B(a[672]), .Z(n3476) );
  XNOR U4176 ( .A(sreg[1695]), .B(n3476), .Z(n3478) );
  NANDN U4177 ( .A(sreg[1694]), .B(n3471), .Z(n3475) );
  NAND U4178 ( .A(n3473), .B(n3472), .Z(n3474) );
  NAND U4179 ( .A(n3475), .B(n3474), .Z(n3477) );
  XNOR U4180 ( .A(n3478), .B(n3477), .Z(c[1695]) );
  NAND U4181 ( .A(b[0]), .B(a[673]), .Z(n3481) );
  XNOR U4182 ( .A(sreg[1696]), .B(n3481), .Z(n3483) );
  NANDN U4183 ( .A(sreg[1695]), .B(n3476), .Z(n3480) );
  NAND U4184 ( .A(n3478), .B(n3477), .Z(n3479) );
  NAND U4185 ( .A(n3480), .B(n3479), .Z(n3482) );
  XNOR U4186 ( .A(n3483), .B(n3482), .Z(c[1696]) );
  NAND U4187 ( .A(b[0]), .B(a[674]), .Z(n3486) );
  XNOR U4188 ( .A(sreg[1697]), .B(n3486), .Z(n3488) );
  NANDN U4189 ( .A(sreg[1696]), .B(n3481), .Z(n3485) );
  NAND U4190 ( .A(n3483), .B(n3482), .Z(n3484) );
  NAND U4191 ( .A(n3485), .B(n3484), .Z(n3487) );
  XNOR U4192 ( .A(n3488), .B(n3487), .Z(c[1697]) );
  NAND U4193 ( .A(b[0]), .B(a[675]), .Z(n3491) );
  XNOR U4194 ( .A(sreg[1698]), .B(n3491), .Z(n3493) );
  NANDN U4195 ( .A(sreg[1697]), .B(n3486), .Z(n3490) );
  NAND U4196 ( .A(n3488), .B(n3487), .Z(n3489) );
  AND U4197 ( .A(n3490), .B(n3489), .Z(n3492) );
  XOR U4198 ( .A(n3493), .B(n3492), .Z(c[1698]) );
  NANDN U4199 ( .A(n3491), .B(sreg[1698]), .Z(n3495) );
  NAND U4200 ( .A(n3493), .B(n3492), .Z(n3494) );
  AND U4201 ( .A(n3495), .B(n3494), .Z(n3498) );
  NAND U4202 ( .A(b[0]), .B(a[676]), .Z(n3496) );
  XNOR U4203 ( .A(sreg[1699]), .B(n3496), .Z(n3497) );
  XNOR U4204 ( .A(n3498), .B(n3497), .Z(c[1699]) );
  NAND U4205 ( .A(b[0]), .B(a[677]), .Z(n3501) );
  XNOR U4206 ( .A(sreg[1700]), .B(n3501), .Z(n3503) );
  NANDN U4207 ( .A(sreg[1699]), .B(n3496), .Z(n3500) );
  NAND U4208 ( .A(n3498), .B(n3497), .Z(n3499) );
  NAND U4209 ( .A(n3500), .B(n3499), .Z(n3502) );
  XNOR U4210 ( .A(n3503), .B(n3502), .Z(c[1700]) );
  NAND U4211 ( .A(b[0]), .B(a[678]), .Z(n3506) );
  XNOR U4212 ( .A(sreg[1701]), .B(n3506), .Z(n3508) );
  NANDN U4213 ( .A(sreg[1700]), .B(n3501), .Z(n3505) );
  NAND U4214 ( .A(n3503), .B(n3502), .Z(n3504) );
  NAND U4215 ( .A(n3505), .B(n3504), .Z(n3507) );
  XNOR U4216 ( .A(n3508), .B(n3507), .Z(c[1701]) );
  NAND U4217 ( .A(b[0]), .B(a[679]), .Z(n3511) );
  XNOR U4218 ( .A(sreg[1702]), .B(n3511), .Z(n3513) );
  NANDN U4219 ( .A(sreg[1701]), .B(n3506), .Z(n3510) );
  NAND U4220 ( .A(n3508), .B(n3507), .Z(n3509) );
  NAND U4221 ( .A(n3510), .B(n3509), .Z(n3512) );
  XNOR U4222 ( .A(n3513), .B(n3512), .Z(c[1702]) );
  NAND U4223 ( .A(b[0]), .B(a[680]), .Z(n3516) );
  XNOR U4224 ( .A(sreg[1703]), .B(n3516), .Z(n3518) );
  NANDN U4225 ( .A(sreg[1702]), .B(n3511), .Z(n3515) );
  NAND U4226 ( .A(n3513), .B(n3512), .Z(n3514) );
  NAND U4227 ( .A(n3515), .B(n3514), .Z(n3517) );
  XNOR U4228 ( .A(n3518), .B(n3517), .Z(c[1703]) );
  NAND U4229 ( .A(b[0]), .B(a[681]), .Z(n3521) );
  XNOR U4230 ( .A(sreg[1704]), .B(n3521), .Z(n3523) );
  NANDN U4231 ( .A(sreg[1703]), .B(n3516), .Z(n3520) );
  NAND U4232 ( .A(n3518), .B(n3517), .Z(n3519) );
  NAND U4233 ( .A(n3520), .B(n3519), .Z(n3522) );
  XNOR U4234 ( .A(n3523), .B(n3522), .Z(c[1704]) );
  NAND U4235 ( .A(b[0]), .B(a[682]), .Z(n3526) );
  XNOR U4236 ( .A(sreg[1705]), .B(n3526), .Z(n3528) );
  NANDN U4237 ( .A(sreg[1704]), .B(n3521), .Z(n3525) );
  NAND U4238 ( .A(n3523), .B(n3522), .Z(n3524) );
  NAND U4239 ( .A(n3525), .B(n3524), .Z(n3527) );
  XNOR U4240 ( .A(n3528), .B(n3527), .Z(c[1705]) );
  NAND U4241 ( .A(b[0]), .B(a[683]), .Z(n3531) );
  XNOR U4242 ( .A(sreg[1706]), .B(n3531), .Z(n3533) );
  NANDN U4243 ( .A(sreg[1705]), .B(n3526), .Z(n3530) );
  NAND U4244 ( .A(n3528), .B(n3527), .Z(n3529) );
  NAND U4245 ( .A(n3530), .B(n3529), .Z(n3532) );
  XNOR U4246 ( .A(n3533), .B(n3532), .Z(c[1706]) );
  NAND U4247 ( .A(b[0]), .B(a[684]), .Z(n3536) );
  XNOR U4248 ( .A(sreg[1707]), .B(n3536), .Z(n3538) );
  NANDN U4249 ( .A(sreg[1706]), .B(n3531), .Z(n3535) );
  NAND U4250 ( .A(n3533), .B(n3532), .Z(n3534) );
  NAND U4251 ( .A(n3535), .B(n3534), .Z(n3537) );
  XNOR U4252 ( .A(n3538), .B(n3537), .Z(c[1707]) );
  NANDN U4253 ( .A(sreg[1707]), .B(n3536), .Z(n3540) );
  NAND U4254 ( .A(n3538), .B(n3537), .Z(n3539) );
  AND U4255 ( .A(n3540), .B(n3539), .Z(n3543) );
  NAND U4256 ( .A(b[0]), .B(a[685]), .Z(n3541) );
  XNOR U4257 ( .A(sreg[1708]), .B(n3541), .Z(n3542) );
  XOR U4258 ( .A(n3543), .B(n3542), .Z(c[1708]) );
  NANDN U4259 ( .A(n3541), .B(sreg[1708]), .Z(n3545) );
  NAND U4260 ( .A(n3543), .B(n3542), .Z(n3544) );
  AND U4261 ( .A(n3545), .B(n3544), .Z(n3547) );
  AND U4262 ( .A(b[0]), .B(a[686]), .Z(n3548) );
  XNOR U4263 ( .A(sreg[1709]), .B(n3548), .Z(n3546) );
  XOR U4264 ( .A(n3547), .B(n3546), .Z(c[1709]) );
  NAND U4265 ( .A(b[0]), .B(a[687]), .Z(n3549) );
  XNOR U4266 ( .A(sreg[1710]), .B(n3549), .Z(n3551) );
  XOR U4267 ( .A(n3551), .B(n3550), .Z(c[1710]) );
  NAND U4268 ( .A(b[0]), .B(a[688]), .Z(n3554) );
  XNOR U4269 ( .A(sreg[1711]), .B(n3554), .Z(n3556) );
  NANDN U4270 ( .A(n3549), .B(sreg[1710]), .Z(n3553) );
  NAND U4271 ( .A(n3551), .B(n3550), .Z(n3552) );
  NAND U4272 ( .A(n3553), .B(n3552), .Z(n3555) );
  XOR U4273 ( .A(n3556), .B(n3555), .Z(c[1711]) );
  NANDN U4274 ( .A(n3554), .B(sreg[1711]), .Z(n3558) );
  NAND U4275 ( .A(n3556), .B(n3555), .Z(n3557) );
  NAND U4276 ( .A(n3558), .B(n3557), .Z(n3561) );
  NAND U4277 ( .A(b[0]), .B(a[689]), .Z(n3560) );
  XOR U4278 ( .A(sreg[1712]), .B(n3560), .Z(n3559) );
  XNOR U4279 ( .A(n3561), .B(n3559), .Z(c[1712]) );
  NAND U4280 ( .A(b[0]), .B(a[690]), .Z(n3562) );
  XNOR U4281 ( .A(sreg[1713]), .B(n3562), .Z(n3563) );
  XOR U4282 ( .A(n3564), .B(n3563), .Z(c[1713]) );
  NANDN U4283 ( .A(n3562), .B(sreg[1713]), .Z(n3566) );
  NAND U4284 ( .A(n3564), .B(n3563), .Z(n3565) );
  AND U4285 ( .A(n3566), .B(n3565), .Z(n3569) );
  NAND U4286 ( .A(b[0]), .B(a[691]), .Z(n3567) );
  XNOR U4287 ( .A(sreg[1714]), .B(n3567), .Z(n3568) );
  XNOR U4288 ( .A(n3569), .B(n3568), .Z(c[1714]) );
  NAND U4289 ( .A(b[0]), .B(a[692]), .Z(n3572) );
  XNOR U4290 ( .A(sreg[1715]), .B(n3572), .Z(n3574) );
  NANDN U4291 ( .A(sreg[1714]), .B(n3567), .Z(n3571) );
  NAND U4292 ( .A(n3569), .B(n3568), .Z(n3570) );
  NAND U4293 ( .A(n3571), .B(n3570), .Z(n3573) );
  XNOR U4294 ( .A(n3574), .B(n3573), .Z(c[1715]) );
  NAND U4295 ( .A(b[0]), .B(a[693]), .Z(n3577) );
  XNOR U4296 ( .A(sreg[1716]), .B(n3577), .Z(n3579) );
  NANDN U4297 ( .A(sreg[1715]), .B(n3572), .Z(n3576) );
  NAND U4298 ( .A(n3574), .B(n3573), .Z(n3575) );
  NAND U4299 ( .A(n3576), .B(n3575), .Z(n3578) );
  XNOR U4300 ( .A(n3579), .B(n3578), .Z(c[1716]) );
  NAND U4301 ( .A(b[0]), .B(a[694]), .Z(n3582) );
  XNOR U4302 ( .A(sreg[1717]), .B(n3582), .Z(n3584) );
  NANDN U4303 ( .A(sreg[1716]), .B(n3577), .Z(n3581) );
  NAND U4304 ( .A(n3579), .B(n3578), .Z(n3580) );
  NAND U4305 ( .A(n3581), .B(n3580), .Z(n3583) );
  XNOR U4306 ( .A(n3584), .B(n3583), .Z(c[1717]) );
  NAND U4307 ( .A(b[0]), .B(a[695]), .Z(n3587) );
  XNOR U4308 ( .A(sreg[1718]), .B(n3587), .Z(n3589) );
  NANDN U4309 ( .A(sreg[1717]), .B(n3582), .Z(n3586) );
  NAND U4310 ( .A(n3584), .B(n3583), .Z(n3585) );
  NAND U4311 ( .A(n3586), .B(n3585), .Z(n3588) );
  XNOR U4312 ( .A(n3589), .B(n3588), .Z(c[1718]) );
  NAND U4313 ( .A(b[0]), .B(a[696]), .Z(n3592) );
  XNOR U4314 ( .A(sreg[1719]), .B(n3592), .Z(n3594) );
  NANDN U4315 ( .A(sreg[1718]), .B(n3587), .Z(n3591) );
  NAND U4316 ( .A(n3589), .B(n3588), .Z(n3590) );
  NAND U4317 ( .A(n3591), .B(n3590), .Z(n3593) );
  XNOR U4318 ( .A(n3594), .B(n3593), .Z(c[1719]) );
  NAND U4319 ( .A(b[0]), .B(a[697]), .Z(n3597) );
  XNOR U4320 ( .A(sreg[1720]), .B(n3597), .Z(n3599) );
  NANDN U4321 ( .A(sreg[1719]), .B(n3592), .Z(n3596) );
  NAND U4322 ( .A(n3594), .B(n3593), .Z(n3595) );
  NAND U4323 ( .A(n3596), .B(n3595), .Z(n3598) );
  XNOR U4324 ( .A(n3599), .B(n3598), .Z(c[1720]) );
  NANDN U4325 ( .A(sreg[1720]), .B(n3597), .Z(n3601) );
  NAND U4326 ( .A(n3599), .B(n3598), .Z(n3600) );
  AND U4327 ( .A(n3601), .B(n3600), .Z(n3604) );
  NAND U4328 ( .A(b[0]), .B(a[698]), .Z(n3602) );
  XNOR U4329 ( .A(sreg[1721]), .B(n3602), .Z(n3603) );
  XOR U4330 ( .A(n3604), .B(n3603), .Z(c[1721]) );
  NAND U4331 ( .A(b[0]), .B(a[699]), .Z(n3607) );
  XNOR U4332 ( .A(sreg[1722]), .B(n3607), .Z(n3609) );
  NANDN U4333 ( .A(n3602), .B(sreg[1721]), .Z(n3606) );
  NAND U4334 ( .A(n3604), .B(n3603), .Z(n3605) );
  AND U4335 ( .A(n3606), .B(n3605), .Z(n3608) );
  XNOR U4336 ( .A(n3609), .B(n3608), .Z(c[1722]) );
  NAND U4337 ( .A(b[0]), .B(a[700]), .Z(n3612) );
  XNOR U4338 ( .A(sreg[1723]), .B(n3612), .Z(n3614) );
  NANDN U4339 ( .A(sreg[1722]), .B(n3607), .Z(n3611) );
  NAND U4340 ( .A(n3609), .B(n3608), .Z(n3610) );
  NAND U4341 ( .A(n3611), .B(n3610), .Z(n3613) );
  XNOR U4342 ( .A(n3614), .B(n3613), .Z(c[1723]) );
  NAND U4343 ( .A(b[0]), .B(a[701]), .Z(n3617) );
  XNOR U4344 ( .A(sreg[1724]), .B(n3617), .Z(n3619) );
  NANDN U4345 ( .A(sreg[1723]), .B(n3612), .Z(n3616) );
  NAND U4346 ( .A(n3614), .B(n3613), .Z(n3615) );
  AND U4347 ( .A(n3616), .B(n3615), .Z(n3618) );
  XOR U4348 ( .A(n3619), .B(n3618), .Z(c[1724]) );
  NAND U4349 ( .A(b[0]), .B(a[702]), .Z(n3622) );
  XNOR U4350 ( .A(sreg[1725]), .B(n3622), .Z(n3624) );
  NANDN U4351 ( .A(n3617), .B(sreg[1724]), .Z(n3621) );
  NAND U4352 ( .A(n3619), .B(n3618), .Z(n3620) );
  NAND U4353 ( .A(n3621), .B(n3620), .Z(n3623) );
  XOR U4354 ( .A(n3624), .B(n3623), .Z(c[1725]) );
  NAND U4355 ( .A(b[0]), .B(a[703]), .Z(n3627) );
  XNOR U4356 ( .A(sreg[1726]), .B(n3627), .Z(n3629) );
  NANDN U4357 ( .A(n3622), .B(sreg[1725]), .Z(n3626) );
  NAND U4358 ( .A(n3624), .B(n3623), .Z(n3625) );
  AND U4359 ( .A(n3626), .B(n3625), .Z(n3628) );
  XNOR U4360 ( .A(n3629), .B(n3628), .Z(c[1726]) );
  NAND U4361 ( .A(b[0]), .B(a[704]), .Z(n3632) );
  XNOR U4362 ( .A(sreg[1727]), .B(n3632), .Z(n3634) );
  NANDN U4363 ( .A(sreg[1726]), .B(n3627), .Z(n3631) );
  NAND U4364 ( .A(n3629), .B(n3628), .Z(n3630) );
  NAND U4365 ( .A(n3631), .B(n3630), .Z(n3633) );
  XNOR U4366 ( .A(n3634), .B(n3633), .Z(c[1727]) );
  NAND U4367 ( .A(b[0]), .B(a[705]), .Z(n3637) );
  XNOR U4368 ( .A(sreg[1728]), .B(n3637), .Z(n3639) );
  NANDN U4369 ( .A(sreg[1727]), .B(n3632), .Z(n3636) );
  NAND U4370 ( .A(n3634), .B(n3633), .Z(n3635) );
  AND U4371 ( .A(n3636), .B(n3635), .Z(n3638) );
  XOR U4372 ( .A(n3639), .B(n3638), .Z(c[1728]) );
  NAND U4373 ( .A(b[0]), .B(a[706]), .Z(n3642) );
  XNOR U4374 ( .A(sreg[1729]), .B(n3642), .Z(n3644) );
  NANDN U4375 ( .A(n3637), .B(sreg[1728]), .Z(n3641) );
  NAND U4376 ( .A(n3639), .B(n3638), .Z(n3640) );
  NAND U4377 ( .A(n3641), .B(n3640), .Z(n3643) );
  XOR U4378 ( .A(n3644), .B(n3643), .Z(c[1729]) );
  NAND U4379 ( .A(b[0]), .B(a[707]), .Z(n3647) );
  XNOR U4380 ( .A(sreg[1730]), .B(n3647), .Z(n3649) );
  NANDN U4381 ( .A(n3642), .B(sreg[1729]), .Z(n3646) );
  NAND U4382 ( .A(n3644), .B(n3643), .Z(n3645) );
  AND U4383 ( .A(n3646), .B(n3645), .Z(n3648) );
  XNOR U4384 ( .A(n3649), .B(n3648), .Z(c[1730]) );
  NAND U4385 ( .A(b[0]), .B(a[708]), .Z(n3652) );
  XNOR U4386 ( .A(sreg[1731]), .B(n3652), .Z(n3654) );
  NANDN U4387 ( .A(sreg[1730]), .B(n3647), .Z(n3651) );
  NAND U4388 ( .A(n3649), .B(n3648), .Z(n3650) );
  AND U4389 ( .A(n3651), .B(n3650), .Z(n3653) );
  XOR U4390 ( .A(n3654), .B(n3653), .Z(c[1731]) );
  NAND U4391 ( .A(b[0]), .B(a[709]), .Z(n3657) );
  XNOR U4392 ( .A(sreg[1732]), .B(n3657), .Z(n3659) );
  NANDN U4393 ( .A(n3652), .B(sreg[1731]), .Z(n3656) );
  NAND U4394 ( .A(n3654), .B(n3653), .Z(n3655) );
  NAND U4395 ( .A(n3656), .B(n3655), .Z(n3658) );
  XOR U4396 ( .A(n3659), .B(n3658), .Z(c[1732]) );
  NAND U4397 ( .A(b[0]), .B(a[710]), .Z(n3662) );
  XNOR U4398 ( .A(sreg[1733]), .B(n3662), .Z(n3664) );
  NANDN U4399 ( .A(n3657), .B(sreg[1732]), .Z(n3661) );
  NAND U4400 ( .A(n3659), .B(n3658), .Z(n3660) );
  AND U4401 ( .A(n3661), .B(n3660), .Z(n3663) );
  XNOR U4402 ( .A(n3664), .B(n3663), .Z(c[1733]) );
  NAND U4403 ( .A(b[0]), .B(a[711]), .Z(n3667) );
  XNOR U4404 ( .A(sreg[1734]), .B(n3667), .Z(n3669) );
  NANDN U4405 ( .A(sreg[1733]), .B(n3662), .Z(n3666) );
  NAND U4406 ( .A(n3664), .B(n3663), .Z(n3665) );
  NAND U4407 ( .A(n3666), .B(n3665), .Z(n3668) );
  XNOR U4408 ( .A(n3669), .B(n3668), .Z(c[1734]) );
  NAND U4409 ( .A(b[0]), .B(a[712]), .Z(n3672) );
  XNOR U4410 ( .A(sreg[1735]), .B(n3672), .Z(n3674) );
  NANDN U4411 ( .A(sreg[1734]), .B(n3667), .Z(n3671) );
  NAND U4412 ( .A(n3669), .B(n3668), .Z(n3670) );
  NAND U4413 ( .A(n3671), .B(n3670), .Z(n3673) );
  XNOR U4414 ( .A(n3674), .B(n3673), .Z(c[1735]) );
  NAND U4415 ( .A(b[0]), .B(a[713]), .Z(n3677) );
  XNOR U4416 ( .A(sreg[1736]), .B(n3677), .Z(n3679) );
  NANDN U4417 ( .A(sreg[1735]), .B(n3672), .Z(n3676) );
  NAND U4418 ( .A(n3674), .B(n3673), .Z(n3675) );
  NAND U4419 ( .A(n3676), .B(n3675), .Z(n3678) );
  XNOR U4420 ( .A(n3679), .B(n3678), .Z(c[1736]) );
  NAND U4421 ( .A(b[0]), .B(a[714]), .Z(n3682) );
  XNOR U4422 ( .A(sreg[1737]), .B(n3682), .Z(n3684) );
  NANDN U4423 ( .A(sreg[1736]), .B(n3677), .Z(n3681) );
  NAND U4424 ( .A(n3679), .B(n3678), .Z(n3680) );
  NAND U4425 ( .A(n3681), .B(n3680), .Z(n3683) );
  XNOR U4426 ( .A(n3684), .B(n3683), .Z(c[1737]) );
  NAND U4427 ( .A(b[0]), .B(a[715]), .Z(n3687) );
  XNOR U4428 ( .A(sreg[1738]), .B(n3687), .Z(n3689) );
  NANDN U4429 ( .A(sreg[1737]), .B(n3682), .Z(n3686) );
  NAND U4430 ( .A(n3684), .B(n3683), .Z(n3685) );
  NAND U4431 ( .A(n3686), .B(n3685), .Z(n3688) );
  XNOR U4432 ( .A(n3689), .B(n3688), .Z(c[1738]) );
  NAND U4433 ( .A(b[0]), .B(a[716]), .Z(n3692) );
  XNOR U4434 ( .A(sreg[1739]), .B(n3692), .Z(n3694) );
  NANDN U4435 ( .A(sreg[1738]), .B(n3687), .Z(n3691) );
  NAND U4436 ( .A(n3689), .B(n3688), .Z(n3690) );
  NAND U4437 ( .A(n3691), .B(n3690), .Z(n3693) );
  XNOR U4438 ( .A(n3694), .B(n3693), .Z(c[1739]) );
  NAND U4439 ( .A(b[0]), .B(a[717]), .Z(n3697) );
  XNOR U4440 ( .A(sreg[1740]), .B(n3697), .Z(n3699) );
  NANDN U4441 ( .A(sreg[1739]), .B(n3692), .Z(n3696) );
  NAND U4442 ( .A(n3694), .B(n3693), .Z(n3695) );
  NAND U4443 ( .A(n3696), .B(n3695), .Z(n3698) );
  XNOR U4444 ( .A(n3699), .B(n3698), .Z(c[1740]) );
  NANDN U4445 ( .A(sreg[1740]), .B(n3697), .Z(n3701) );
  NAND U4446 ( .A(n3699), .B(n3698), .Z(n3700) );
  AND U4447 ( .A(n3701), .B(n3700), .Z(n3704) );
  NAND U4448 ( .A(b[0]), .B(a[718]), .Z(n3702) );
  XNOR U4449 ( .A(sreg[1741]), .B(n3702), .Z(n3703) );
  XOR U4450 ( .A(n3704), .B(n3703), .Z(c[1741]) );
  NAND U4451 ( .A(b[0]), .B(a[719]), .Z(n3707) );
  XNOR U4452 ( .A(sreg[1742]), .B(n3707), .Z(n3709) );
  NANDN U4453 ( .A(n3702), .B(sreg[1741]), .Z(n3706) );
  NAND U4454 ( .A(n3704), .B(n3703), .Z(n3705) );
  NAND U4455 ( .A(n3706), .B(n3705), .Z(n3708) );
  XOR U4456 ( .A(n3709), .B(n3708), .Z(c[1742]) );
  NAND U4457 ( .A(b[0]), .B(a[720]), .Z(n3712) );
  XNOR U4458 ( .A(sreg[1743]), .B(n3712), .Z(n3714) );
  NANDN U4459 ( .A(n3707), .B(sreg[1742]), .Z(n3711) );
  NAND U4460 ( .A(n3709), .B(n3708), .Z(n3710) );
  AND U4461 ( .A(n3711), .B(n3710), .Z(n3713) );
  XNOR U4462 ( .A(n3714), .B(n3713), .Z(c[1743]) );
  NAND U4463 ( .A(b[0]), .B(a[721]), .Z(n3717) );
  XNOR U4464 ( .A(sreg[1744]), .B(n3717), .Z(n3719) );
  NANDN U4465 ( .A(sreg[1743]), .B(n3712), .Z(n3716) );
  NAND U4466 ( .A(n3714), .B(n3713), .Z(n3715) );
  AND U4467 ( .A(n3716), .B(n3715), .Z(n3718) );
  XOR U4468 ( .A(n3719), .B(n3718), .Z(c[1744]) );
  NAND U4469 ( .A(b[0]), .B(a[722]), .Z(n3722) );
  XNOR U4470 ( .A(sreg[1745]), .B(n3722), .Z(n3724) );
  NANDN U4471 ( .A(n3717), .B(sreg[1744]), .Z(n3721) );
  NAND U4472 ( .A(n3719), .B(n3718), .Z(n3720) );
  NAND U4473 ( .A(n3721), .B(n3720), .Z(n3723) );
  XOR U4474 ( .A(n3724), .B(n3723), .Z(c[1745]) );
  NAND U4475 ( .A(b[0]), .B(a[723]), .Z(n3727) );
  XNOR U4476 ( .A(sreg[1746]), .B(n3727), .Z(n3729) );
  NANDN U4477 ( .A(n3722), .B(sreg[1745]), .Z(n3726) );
  NAND U4478 ( .A(n3724), .B(n3723), .Z(n3725) );
  AND U4479 ( .A(n3726), .B(n3725), .Z(n3728) );
  XNOR U4480 ( .A(n3729), .B(n3728), .Z(c[1746]) );
  NANDN U4481 ( .A(sreg[1746]), .B(n3727), .Z(n3731) );
  NAND U4482 ( .A(n3729), .B(n3728), .Z(n3730) );
  AND U4483 ( .A(n3731), .B(n3730), .Z(n3734) );
  NAND U4484 ( .A(b[0]), .B(a[724]), .Z(n3732) );
  XNOR U4485 ( .A(sreg[1747]), .B(n3732), .Z(n3733) );
  XOR U4486 ( .A(n3734), .B(n3733), .Z(c[1747]) );
  NAND U4487 ( .A(b[0]), .B(a[725]), .Z(n3737) );
  XNOR U4488 ( .A(sreg[1748]), .B(n3737), .Z(n3739) );
  NANDN U4489 ( .A(n3732), .B(sreg[1747]), .Z(n3736) );
  NAND U4490 ( .A(n3734), .B(n3733), .Z(n3735) );
  NAND U4491 ( .A(n3736), .B(n3735), .Z(n3738) );
  XOR U4492 ( .A(n3739), .B(n3738), .Z(c[1748]) );
  NAND U4493 ( .A(b[0]), .B(a[726]), .Z(n3742) );
  XNOR U4494 ( .A(sreg[1749]), .B(n3742), .Z(n3744) );
  NANDN U4495 ( .A(n3737), .B(sreg[1748]), .Z(n3741) );
  NAND U4496 ( .A(n3739), .B(n3738), .Z(n3740) );
  NAND U4497 ( .A(n3741), .B(n3740), .Z(n3743) );
  XOR U4498 ( .A(n3744), .B(n3743), .Z(c[1749]) );
  NAND U4499 ( .A(b[0]), .B(a[727]), .Z(n3747) );
  XNOR U4500 ( .A(sreg[1750]), .B(n3747), .Z(n3749) );
  NANDN U4501 ( .A(n3742), .B(sreg[1749]), .Z(n3746) );
  NAND U4502 ( .A(n3744), .B(n3743), .Z(n3745) );
  NAND U4503 ( .A(n3746), .B(n3745), .Z(n3748) );
  XOR U4504 ( .A(n3749), .B(n3748), .Z(c[1750]) );
  NANDN U4505 ( .A(n3747), .B(sreg[1750]), .Z(n3751) );
  NAND U4506 ( .A(n3749), .B(n3748), .Z(n3750) );
  AND U4507 ( .A(n3751), .B(n3750), .Z(n3754) );
  NAND U4508 ( .A(b[0]), .B(a[728]), .Z(n3752) );
  XNOR U4509 ( .A(sreg[1751]), .B(n3752), .Z(n3753) );
  XNOR U4510 ( .A(n3754), .B(n3753), .Z(c[1751]) );
  NAND U4511 ( .A(b[0]), .B(a[729]), .Z(n3757) );
  XNOR U4512 ( .A(sreg[1752]), .B(n3757), .Z(n3759) );
  NANDN U4513 ( .A(sreg[1751]), .B(n3752), .Z(n3756) );
  NAND U4514 ( .A(n3754), .B(n3753), .Z(n3755) );
  NAND U4515 ( .A(n3756), .B(n3755), .Z(n3758) );
  XNOR U4516 ( .A(n3759), .B(n3758), .Z(c[1752]) );
  NANDN U4517 ( .A(sreg[1752]), .B(n3757), .Z(n3761) );
  NAND U4518 ( .A(n3759), .B(n3758), .Z(n3760) );
  AND U4519 ( .A(n3761), .B(n3760), .Z(n3764) );
  NAND U4520 ( .A(b[0]), .B(a[730]), .Z(n3762) );
  XNOR U4521 ( .A(sreg[1753]), .B(n3762), .Z(n3763) );
  XOR U4522 ( .A(n3764), .B(n3763), .Z(c[1753]) );
  NAND U4523 ( .A(b[0]), .B(a[731]), .Z(n3767) );
  XNOR U4524 ( .A(sreg[1754]), .B(n3767), .Z(n3769) );
  NANDN U4525 ( .A(n3762), .B(sreg[1753]), .Z(n3766) );
  NAND U4526 ( .A(n3764), .B(n3763), .Z(n3765) );
  AND U4527 ( .A(n3766), .B(n3765), .Z(n3768) );
  XNOR U4528 ( .A(n3769), .B(n3768), .Z(c[1754]) );
  NAND U4529 ( .A(b[0]), .B(a[732]), .Z(n3772) );
  XNOR U4530 ( .A(sreg[1755]), .B(n3772), .Z(n3774) );
  NANDN U4531 ( .A(sreg[1754]), .B(n3767), .Z(n3771) );
  NAND U4532 ( .A(n3769), .B(n3768), .Z(n3770) );
  NAND U4533 ( .A(n3771), .B(n3770), .Z(n3773) );
  XNOR U4534 ( .A(n3774), .B(n3773), .Z(c[1755]) );
  NANDN U4535 ( .A(sreg[1755]), .B(n3772), .Z(n3776) );
  NAND U4536 ( .A(n3774), .B(n3773), .Z(n3775) );
  AND U4537 ( .A(n3776), .B(n3775), .Z(n3779) );
  NAND U4538 ( .A(b[0]), .B(a[733]), .Z(n3777) );
  XNOR U4539 ( .A(sreg[1756]), .B(n3777), .Z(n3778) );
  XOR U4540 ( .A(n3779), .B(n3778), .Z(c[1756]) );
  NAND U4541 ( .A(b[0]), .B(a[734]), .Z(n3782) );
  XNOR U4542 ( .A(sreg[1757]), .B(n3782), .Z(n3784) );
  NANDN U4543 ( .A(n3777), .B(sreg[1756]), .Z(n3781) );
  NAND U4544 ( .A(n3779), .B(n3778), .Z(n3780) );
  AND U4545 ( .A(n3781), .B(n3780), .Z(n3783) );
  XNOR U4546 ( .A(n3784), .B(n3783), .Z(c[1757]) );
  NAND U4547 ( .A(b[0]), .B(a[735]), .Z(n3787) );
  XNOR U4548 ( .A(sreg[1758]), .B(n3787), .Z(n3789) );
  NANDN U4549 ( .A(sreg[1757]), .B(n3782), .Z(n3786) );
  NAND U4550 ( .A(n3784), .B(n3783), .Z(n3785) );
  NAND U4551 ( .A(n3786), .B(n3785), .Z(n3788) );
  XNOR U4552 ( .A(n3789), .B(n3788), .Z(c[1758]) );
  NANDN U4553 ( .A(sreg[1758]), .B(n3787), .Z(n3791) );
  NAND U4554 ( .A(n3789), .B(n3788), .Z(n3790) );
  AND U4555 ( .A(n3791), .B(n3790), .Z(n3794) );
  NAND U4556 ( .A(b[0]), .B(a[736]), .Z(n3792) );
  XNOR U4557 ( .A(sreg[1759]), .B(n3792), .Z(n3793) );
  XOR U4558 ( .A(n3794), .B(n3793), .Z(c[1759]) );
  NAND U4559 ( .A(b[0]), .B(a[737]), .Z(n3797) );
  XNOR U4560 ( .A(sreg[1760]), .B(n3797), .Z(n3799) );
  NANDN U4561 ( .A(n3792), .B(sreg[1759]), .Z(n3796) );
  NAND U4562 ( .A(n3794), .B(n3793), .Z(n3795) );
  AND U4563 ( .A(n3796), .B(n3795), .Z(n3798) );
  XNOR U4564 ( .A(n3799), .B(n3798), .Z(c[1760]) );
  NANDN U4565 ( .A(sreg[1760]), .B(n3797), .Z(n3801) );
  NAND U4566 ( .A(n3799), .B(n3798), .Z(n3800) );
  AND U4567 ( .A(n3801), .B(n3800), .Z(n3804) );
  NAND U4568 ( .A(b[0]), .B(a[738]), .Z(n3802) );
  XNOR U4569 ( .A(sreg[1761]), .B(n3802), .Z(n3803) );
  XOR U4570 ( .A(n3804), .B(n3803), .Z(c[1761]) );
  NAND U4571 ( .A(b[0]), .B(a[739]), .Z(n3807) );
  XNOR U4572 ( .A(sreg[1762]), .B(n3807), .Z(n3809) );
  NANDN U4573 ( .A(n3802), .B(sreg[1761]), .Z(n3806) );
  NAND U4574 ( .A(n3804), .B(n3803), .Z(n3805) );
  NAND U4575 ( .A(n3806), .B(n3805), .Z(n3808) );
  XOR U4576 ( .A(n3809), .B(n3808), .Z(c[1762]) );
  NAND U4577 ( .A(b[0]), .B(a[740]), .Z(n3812) );
  XNOR U4578 ( .A(sreg[1763]), .B(n3812), .Z(n3814) );
  NANDN U4579 ( .A(n3807), .B(sreg[1762]), .Z(n3811) );
  NAND U4580 ( .A(n3809), .B(n3808), .Z(n3810) );
  AND U4581 ( .A(n3811), .B(n3810), .Z(n3813) );
  XNOR U4582 ( .A(n3814), .B(n3813), .Z(c[1763]) );
  NANDN U4583 ( .A(sreg[1763]), .B(n3812), .Z(n3816) );
  NAND U4584 ( .A(n3814), .B(n3813), .Z(n3815) );
  AND U4585 ( .A(n3816), .B(n3815), .Z(n3819) );
  NAND U4586 ( .A(b[0]), .B(a[741]), .Z(n3817) );
  XNOR U4587 ( .A(sreg[1764]), .B(n3817), .Z(n3818) );
  XOR U4588 ( .A(n3819), .B(n3818), .Z(c[1764]) );
  NAND U4589 ( .A(b[0]), .B(a[742]), .Z(n3822) );
  XNOR U4590 ( .A(sreg[1765]), .B(n3822), .Z(n3824) );
  NANDN U4591 ( .A(n3817), .B(sreg[1764]), .Z(n3821) );
  NAND U4592 ( .A(n3819), .B(n3818), .Z(n3820) );
  NAND U4593 ( .A(n3821), .B(n3820), .Z(n3823) );
  XOR U4594 ( .A(n3824), .B(n3823), .Z(c[1765]) );
  AND U4595 ( .A(b[0]), .B(a[743]), .Z(n3828) );
  NANDN U4596 ( .A(n3822), .B(sreg[1765]), .Z(n3826) );
  NAND U4597 ( .A(n3824), .B(n3823), .Z(n3825) );
  AND U4598 ( .A(n3826), .B(n3825), .Z(n3829) );
  XNOR U4599 ( .A(sreg[1766]), .B(n3829), .Z(n3827) );
  XOR U4600 ( .A(n3828), .B(n3827), .Z(c[1766]) );
  NAND U4601 ( .A(b[0]), .B(a[744]), .Z(n3830) );
  XNOR U4602 ( .A(sreg[1767]), .B(n3830), .Z(n3831) );
  XNOR U4603 ( .A(n3832), .B(n3831), .Z(c[1767]) );
  NAND U4604 ( .A(b[0]), .B(a[745]), .Z(n3835) );
  XNOR U4605 ( .A(sreg[1768]), .B(n3835), .Z(n3837) );
  NANDN U4606 ( .A(n3830), .B(sreg[1767]), .Z(n3834) );
  NANDN U4607 ( .A(n3832), .B(n3831), .Z(n3833) );
  NAND U4608 ( .A(n3834), .B(n3833), .Z(n3836) );
  XOR U4609 ( .A(n3837), .B(n3836), .Z(c[1768]) );
  NANDN U4610 ( .A(n3835), .B(sreg[1768]), .Z(n3839) );
  NAND U4611 ( .A(n3837), .B(n3836), .Z(n3838) );
  NAND U4612 ( .A(n3839), .B(n3838), .Z(n3842) );
  NAND U4613 ( .A(b[0]), .B(a[746]), .Z(n3841) );
  XOR U4614 ( .A(sreg[1769]), .B(n3841), .Z(n3840) );
  XNOR U4615 ( .A(n3842), .B(n3840), .Z(c[1769]) );
  NAND U4616 ( .A(b[0]), .B(a[747]), .Z(n3843) );
  XNOR U4617 ( .A(sreg[1770]), .B(n3843), .Z(n3844) );
  XOR U4618 ( .A(n3845), .B(n3844), .Z(c[1770]) );
  NAND U4619 ( .A(b[0]), .B(a[748]), .Z(n3848) );
  XNOR U4620 ( .A(sreg[1771]), .B(n3848), .Z(n3850) );
  NANDN U4621 ( .A(n3843), .B(sreg[1770]), .Z(n3847) );
  NAND U4622 ( .A(n3845), .B(n3844), .Z(n3846) );
  NAND U4623 ( .A(n3847), .B(n3846), .Z(n3849) );
  XOR U4624 ( .A(n3850), .B(n3849), .Z(c[1771]) );
  AND U4625 ( .A(b[0]), .B(a[749]), .Z(n3854) );
  NANDN U4626 ( .A(n3848), .B(sreg[1771]), .Z(n3852) );
  NAND U4627 ( .A(n3850), .B(n3849), .Z(n3851) );
  AND U4628 ( .A(n3852), .B(n3851), .Z(n3855) );
  XNOR U4629 ( .A(sreg[1772]), .B(n3855), .Z(n3853) );
  XOR U4630 ( .A(n3854), .B(n3853), .Z(c[1772]) );
  NAND U4631 ( .A(b[0]), .B(a[750]), .Z(n3856) );
  XNOR U4632 ( .A(sreg[1773]), .B(n3856), .Z(n3857) );
  XNOR U4633 ( .A(n3858), .B(n3857), .Z(c[1773]) );
  NAND U4634 ( .A(b[0]), .B(a[751]), .Z(n3861) );
  XNOR U4635 ( .A(sreg[1774]), .B(n3861), .Z(n3863) );
  NANDN U4636 ( .A(n3856), .B(sreg[1773]), .Z(n3860) );
  NANDN U4637 ( .A(n3858), .B(n3857), .Z(n3859) );
  NAND U4638 ( .A(n3860), .B(n3859), .Z(n3862) );
  XOR U4639 ( .A(n3863), .B(n3862), .Z(c[1774]) );
  NAND U4640 ( .A(b[0]), .B(a[752]), .Z(n3868) );
  NANDN U4641 ( .A(n3861), .B(sreg[1774]), .Z(n3865) );
  NAND U4642 ( .A(n3863), .B(n3862), .Z(n3864) );
  NAND U4643 ( .A(n3865), .B(n3864), .Z(n3867) );
  XOR U4644 ( .A(n3867), .B(sreg[1775]), .Z(n3866) );
  XNOR U4645 ( .A(n3868), .B(n3866), .Z(c[1775]) );
  NAND U4646 ( .A(b[0]), .B(a[753]), .Z(n3869) );
  XNOR U4647 ( .A(sreg[1776]), .B(n3869), .Z(n3870) );
  XNOR U4648 ( .A(n3871), .B(n3870), .Z(c[1776]) );
  NAND U4649 ( .A(b[0]), .B(a[754]), .Z(n3874) );
  XNOR U4650 ( .A(sreg[1777]), .B(n3874), .Z(n3876) );
  NANDN U4651 ( .A(n3869), .B(sreg[1776]), .Z(n3873) );
  NANDN U4652 ( .A(n3871), .B(n3870), .Z(n3872) );
  NAND U4653 ( .A(n3873), .B(n3872), .Z(n3875) );
  XOR U4654 ( .A(n3876), .B(n3875), .Z(c[1777]) );
  NAND U4655 ( .A(b[0]), .B(a[755]), .Z(n3879) );
  XNOR U4656 ( .A(sreg[1778]), .B(n3879), .Z(n3881) );
  NANDN U4657 ( .A(n3874), .B(sreg[1777]), .Z(n3878) );
  NAND U4658 ( .A(n3876), .B(n3875), .Z(n3877) );
  NAND U4659 ( .A(n3878), .B(n3877), .Z(n3880) );
  XOR U4660 ( .A(n3881), .B(n3880), .Z(c[1778]) );
  NAND U4661 ( .A(b[0]), .B(a[756]), .Z(n3884) );
  XNOR U4662 ( .A(sreg[1779]), .B(n3884), .Z(n3886) );
  NANDN U4663 ( .A(n3879), .B(sreg[1778]), .Z(n3883) );
  NAND U4664 ( .A(n3881), .B(n3880), .Z(n3882) );
  NAND U4665 ( .A(n3883), .B(n3882), .Z(n3885) );
  XOR U4666 ( .A(n3886), .B(n3885), .Z(c[1779]) );
  NAND U4667 ( .A(b[0]), .B(a[757]), .Z(n3889) );
  XNOR U4668 ( .A(sreg[1780]), .B(n3889), .Z(n3891) );
  NANDN U4669 ( .A(n3884), .B(sreg[1779]), .Z(n3888) );
  NAND U4670 ( .A(n3886), .B(n3885), .Z(n3887) );
  NAND U4671 ( .A(n3888), .B(n3887), .Z(n3890) );
  XOR U4672 ( .A(n3891), .B(n3890), .Z(c[1780]) );
  NAND U4673 ( .A(b[0]), .B(a[758]), .Z(n3894) );
  XNOR U4674 ( .A(sreg[1781]), .B(n3894), .Z(n3896) );
  NANDN U4675 ( .A(n3889), .B(sreg[1780]), .Z(n3893) );
  NAND U4676 ( .A(n3891), .B(n3890), .Z(n3892) );
  NAND U4677 ( .A(n3893), .B(n3892), .Z(n3895) );
  XOR U4678 ( .A(n3896), .B(n3895), .Z(c[1781]) );
  NANDN U4679 ( .A(n3894), .B(sreg[1781]), .Z(n3898) );
  NAND U4680 ( .A(n3896), .B(n3895), .Z(n3897) );
  AND U4681 ( .A(n3898), .B(n3897), .Z(n3901) );
  NAND U4682 ( .A(b[0]), .B(a[759]), .Z(n3899) );
  XNOR U4683 ( .A(sreg[1782]), .B(n3899), .Z(n3900) );
  XNOR U4684 ( .A(n3901), .B(n3900), .Z(c[1782]) );
  NAND U4685 ( .A(b[0]), .B(a[760]), .Z(n3904) );
  XNOR U4686 ( .A(sreg[1783]), .B(n3904), .Z(n3906) );
  NANDN U4687 ( .A(sreg[1782]), .B(n3899), .Z(n3903) );
  NAND U4688 ( .A(n3901), .B(n3900), .Z(n3902) );
  NAND U4689 ( .A(n3903), .B(n3902), .Z(n3905) );
  XNOR U4690 ( .A(n3906), .B(n3905), .Z(c[1783]) );
  NAND U4691 ( .A(b[0]), .B(a[761]), .Z(n3909) );
  XNOR U4692 ( .A(sreg[1784]), .B(n3909), .Z(n3911) );
  NANDN U4693 ( .A(sreg[1783]), .B(n3904), .Z(n3908) );
  NAND U4694 ( .A(n3906), .B(n3905), .Z(n3907) );
  NAND U4695 ( .A(n3908), .B(n3907), .Z(n3910) );
  XNOR U4696 ( .A(n3911), .B(n3910), .Z(c[1784]) );
  NAND U4697 ( .A(b[0]), .B(a[762]), .Z(n3914) );
  XNOR U4698 ( .A(sreg[1785]), .B(n3914), .Z(n3916) );
  NANDN U4699 ( .A(sreg[1784]), .B(n3909), .Z(n3913) );
  NAND U4700 ( .A(n3911), .B(n3910), .Z(n3912) );
  NAND U4701 ( .A(n3913), .B(n3912), .Z(n3915) );
  XNOR U4702 ( .A(n3916), .B(n3915), .Z(c[1785]) );
  NAND U4703 ( .A(b[0]), .B(a[763]), .Z(n3919) );
  XNOR U4704 ( .A(sreg[1786]), .B(n3919), .Z(n3921) );
  NANDN U4705 ( .A(sreg[1785]), .B(n3914), .Z(n3918) );
  NAND U4706 ( .A(n3916), .B(n3915), .Z(n3917) );
  NAND U4707 ( .A(n3918), .B(n3917), .Z(n3920) );
  XNOR U4708 ( .A(n3921), .B(n3920), .Z(c[1786]) );
  NAND U4709 ( .A(b[0]), .B(a[764]), .Z(n3924) );
  XNOR U4710 ( .A(sreg[1787]), .B(n3924), .Z(n3926) );
  NANDN U4711 ( .A(sreg[1786]), .B(n3919), .Z(n3923) );
  NAND U4712 ( .A(n3921), .B(n3920), .Z(n3922) );
  NAND U4713 ( .A(n3923), .B(n3922), .Z(n3925) );
  XNOR U4714 ( .A(n3926), .B(n3925), .Z(c[1787]) );
  NAND U4715 ( .A(b[0]), .B(a[765]), .Z(n3929) );
  XNOR U4716 ( .A(sreg[1788]), .B(n3929), .Z(n3931) );
  NANDN U4717 ( .A(sreg[1787]), .B(n3924), .Z(n3928) );
  NAND U4718 ( .A(n3926), .B(n3925), .Z(n3927) );
  NAND U4719 ( .A(n3928), .B(n3927), .Z(n3930) );
  XNOR U4720 ( .A(n3931), .B(n3930), .Z(c[1788]) );
  NAND U4721 ( .A(b[0]), .B(a[766]), .Z(n3934) );
  XNOR U4722 ( .A(sreg[1789]), .B(n3934), .Z(n3936) );
  NANDN U4723 ( .A(sreg[1788]), .B(n3929), .Z(n3933) );
  NAND U4724 ( .A(n3931), .B(n3930), .Z(n3932) );
  NAND U4725 ( .A(n3933), .B(n3932), .Z(n3935) );
  XNOR U4726 ( .A(n3936), .B(n3935), .Z(c[1789]) );
  NAND U4727 ( .A(b[0]), .B(a[767]), .Z(n3939) );
  XNOR U4728 ( .A(sreg[1790]), .B(n3939), .Z(n3941) );
  NANDN U4729 ( .A(sreg[1789]), .B(n3934), .Z(n3938) );
  NAND U4730 ( .A(n3936), .B(n3935), .Z(n3937) );
  NAND U4731 ( .A(n3938), .B(n3937), .Z(n3940) );
  XNOR U4732 ( .A(n3941), .B(n3940), .Z(c[1790]) );
  NAND U4733 ( .A(b[0]), .B(a[768]), .Z(n3944) );
  XNOR U4734 ( .A(sreg[1791]), .B(n3944), .Z(n3946) );
  NANDN U4735 ( .A(sreg[1790]), .B(n3939), .Z(n3943) );
  NAND U4736 ( .A(n3941), .B(n3940), .Z(n3942) );
  NAND U4737 ( .A(n3943), .B(n3942), .Z(n3945) );
  XNOR U4738 ( .A(n3946), .B(n3945), .Z(c[1791]) );
  NAND U4739 ( .A(b[0]), .B(a[769]), .Z(n3949) );
  XNOR U4740 ( .A(sreg[1792]), .B(n3949), .Z(n3951) );
  NANDN U4741 ( .A(sreg[1791]), .B(n3944), .Z(n3948) );
  NAND U4742 ( .A(n3946), .B(n3945), .Z(n3947) );
  NAND U4743 ( .A(n3948), .B(n3947), .Z(n3950) );
  XNOR U4744 ( .A(n3951), .B(n3950), .Z(c[1792]) );
  NAND U4745 ( .A(b[0]), .B(a[770]), .Z(n3954) );
  XNOR U4746 ( .A(sreg[1793]), .B(n3954), .Z(n3956) );
  NANDN U4747 ( .A(sreg[1792]), .B(n3949), .Z(n3953) );
  NAND U4748 ( .A(n3951), .B(n3950), .Z(n3952) );
  NAND U4749 ( .A(n3953), .B(n3952), .Z(n3955) );
  XNOR U4750 ( .A(n3956), .B(n3955), .Z(c[1793]) );
  NANDN U4751 ( .A(sreg[1793]), .B(n3954), .Z(n3958) );
  NAND U4752 ( .A(n3956), .B(n3955), .Z(n3957) );
  AND U4753 ( .A(n3958), .B(n3957), .Z(n3961) );
  NAND U4754 ( .A(b[0]), .B(a[771]), .Z(n3959) );
  XNOR U4755 ( .A(sreg[1794]), .B(n3959), .Z(n3960) );
  XOR U4756 ( .A(n3961), .B(n3960), .Z(c[1794]) );
  NAND U4757 ( .A(b[0]), .B(a[772]), .Z(n3964) );
  XNOR U4758 ( .A(sreg[1795]), .B(n3964), .Z(n3966) );
  NANDN U4759 ( .A(n3959), .B(sreg[1794]), .Z(n3963) );
  NAND U4760 ( .A(n3961), .B(n3960), .Z(n3962) );
  NAND U4761 ( .A(n3963), .B(n3962), .Z(n3965) );
  XOR U4762 ( .A(n3966), .B(n3965), .Z(c[1795]) );
  NANDN U4763 ( .A(n3964), .B(sreg[1795]), .Z(n3968) );
  NAND U4764 ( .A(n3966), .B(n3965), .Z(n3967) );
  AND U4765 ( .A(n3968), .B(n3967), .Z(n3971) );
  NAND U4766 ( .A(b[0]), .B(a[773]), .Z(n3969) );
  XNOR U4767 ( .A(sreg[1796]), .B(n3969), .Z(n3970) );
  XNOR U4768 ( .A(n3971), .B(n3970), .Z(c[1796]) );
  NAND U4769 ( .A(b[0]), .B(a[774]), .Z(n3974) );
  XNOR U4770 ( .A(sreg[1797]), .B(n3974), .Z(n3976) );
  NANDN U4771 ( .A(sreg[1796]), .B(n3969), .Z(n3973) );
  NAND U4772 ( .A(n3971), .B(n3970), .Z(n3972) );
  AND U4773 ( .A(n3973), .B(n3972), .Z(n3975) );
  XOR U4774 ( .A(n3976), .B(n3975), .Z(c[1797]) );
  NAND U4775 ( .A(b[0]), .B(a[775]), .Z(n3979) );
  XNOR U4776 ( .A(sreg[1798]), .B(n3979), .Z(n3981) );
  NANDN U4777 ( .A(n3974), .B(sreg[1797]), .Z(n3978) );
  NAND U4778 ( .A(n3976), .B(n3975), .Z(n3977) );
  NAND U4779 ( .A(n3978), .B(n3977), .Z(n3980) );
  XOR U4780 ( .A(n3981), .B(n3980), .Z(c[1798]) );
  NANDN U4781 ( .A(n3979), .B(sreg[1798]), .Z(n3983) );
  NAND U4782 ( .A(n3981), .B(n3980), .Z(n3982) );
  AND U4783 ( .A(n3983), .B(n3982), .Z(n3986) );
  NAND U4784 ( .A(b[0]), .B(a[776]), .Z(n3984) );
  XNOR U4785 ( .A(sreg[1799]), .B(n3984), .Z(n3985) );
  XNOR U4786 ( .A(n3986), .B(n3985), .Z(c[1799]) );
  NAND U4787 ( .A(b[0]), .B(a[777]), .Z(n3989) );
  XNOR U4788 ( .A(sreg[1800]), .B(n3989), .Z(n3991) );
  NANDN U4789 ( .A(sreg[1799]), .B(n3984), .Z(n3988) );
  NAND U4790 ( .A(n3986), .B(n3985), .Z(n3987) );
  NAND U4791 ( .A(n3988), .B(n3987), .Z(n3990) );
  XNOR U4792 ( .A(n3991), .B(n3990), .Z(c[1800]) );
  NANDN U4793 ( .A(sreg[1800]), .B(n3989), .Z(n3993) );
  NAND U4794 ( .A(n3991), .B(n3990), .Z(n3992) );
  AND U4795 ( .A(n3993), .B(n3992), .Z(n3996) );
  NAND U4796 ( .A(b[0]), .B(a[778]), .Z(n3994) );
  XNOR U4797 ( .A(sreg[1801]), .B(n3994), .Z(n3995) );
  XOR U4798 ( .A(n3996), .B(n3995), .Z(c[1801]) );
  NAND U4799 ( .A(b[0]), .B(a[779]), .Z(n3999) );
  XNOR U4800 ( .A(sreg[1802]), .B(n3999), .Z(n4001) );
  NANDN U4801 ( .A(n3994), .B(sreg[1801]), .Z(n3998) );
  NAND U4802 ( .A(n3996), .B(n3995), .Z(n3997) );
  AND U4803 ( .A(n3998), .B(n3997), .Z(n4000) );
  XNOR U4804 ( .A(n4001), .B(n4000), .Z(c[1802]) );
  NAND U4805 ( .A(b[0]), .B(a[780]), .Z(n4004) );
  XNOR U4806 ( .A(sreg[1803]), .B(n4004), .Z(n4006) );
  NANDN U4807 ( .A(sreg[1802]), .B(n3999), .Z(n4003) );
  NAND U4808 ( .A(n4001), .B(n4000), .Z(n4002) );
  NAND U4809 ( .A(n4003), .B(n4002), .Z(n4005) );
  XNOR U4810 ( .A(n4006), .B(n4005), .Z(c[1803]) );
  NANDN U4811 ( .A(sreg[1803]), .B(n4004), .Z(n4008) );
  NAND U4812 ( .A(n4006), .B(n4005), .Z(n4007) );
  AND U4813 ( .A(n4008), .B(n4007), .Z(n4011) );
  NAND U4814 ( .A(b[0]), .B(a[781]), .Z(n4009) );
  XNOR U4815 ( .A(sreg[1804]), .B(n4009), .Z(n4010) );
  XOR U4816 ( .A(n4011), .B(n4010), .Z(c[1804]) );
  NAND U4817 ( .A(b[0]), .B(a[782]), .Z(n4014) );
  XNOR U4818 ( .A(sreg[1805]), .B(n4014), .Z(n4016) );
  NANDN U4819 ( .A(n4009), .B(sreg[1804]), .Z(n4013) );
  NAND U4820 ( .A(n4011), .B(n4010), .Z(n4012) );
  NAND U4821 ( .A(n4013), .B(n4012), .Z(n4015) );
  XOR U4822 ( .A(n4016), .B(n4015), .Z(c[1805]) );
  NAND U4823 ( .A(b[0]), .B(a[783]), .Z(n4019) );
  XNOR U4824 ( .A(sreg[1806]), .B(n4019), .Z(n4021) );
  NANDN U4825 ( .A(n4014), .B(sreg[1805]), .Z(n4018) );
  NAND U4826 ( .A(n4016), .B(n4015), .Z(n4017) );
  NAND U4827 ( .A(n4018), .B(n4017), .Z(n4020) );
  XOR U4828 ( .A(n4021), .B(n4020), .Z(c[1806]) );
  NAND U4829 ( .A(b[0]), .B(a[784]), .Z(n4024) );
  XNOR U4830 ( .A(sreg[1807]), .B(n4024), .Z(n4026) );
  NANDN U4831 ( .A(n4019), .B(sreg[1806]), .Z(n4023) );
  NAND U4832 ( .A(n4021), .B(n4020), .Z(n4022) );
  NAND U4833 ( .A(n4023), .B(n4022), .Z(n4025) );
  XOR U4834 ( .A(n4026), .B(n4025), .Z(c[1807]) );
  NAND U4835 ( .A(b[0]), .B(a[785]), .Z(n4029) );
  XNOR U4836 ( .A(sreg[1808]), .B(n4029), .Z(n4031) );
  NANDN U4837 ( .A(n4024), .B(sreg[1807]), .Z(n4028) );
  NAND U4838 ( .A(n4026), .B(n4025), .Z(n4027) );
  NAND U4839 ( .A(n4028), .B(n4027), .Z(n4030) );
  XOR U4840 ( .A(n4031), .B(n4030), .Z(c[1808]) );
  NAND U4841 ( .A(b[0]), .B(a[786]), .Z(n4034) );
  XNOR U4842 ( .A(sreg[1809]), .B(n4034), .Z(n4036) );
  NANDN U4843 ( .A(n4029), .B(sreg[1808]), .Z(n4033) );
  NAND U4844 ( .A(n4031), .B(n4030), .Z(n4032) );
  NAND U4845 ( .A(n4033), .B(n4032), .Z(n4035) );
  XOR U4846 ( .A(n4036), .B(n4035), .Z(c[1809]) );
  NAND U4847 ( .A(b[0]), .B(a[787]), .Z(n4039) );
  XNOR U4848 ( .A(sreg[1810]), .B(n4039), .Z(n4041) );
  NANDN U4849 ( .A(n4034), .B(sreg[1809]), .Z(n4038) );
  NAND U4850 ( .A(n4036), .B(n4035), .Z(n4037) );
  NAND U4851 ( .A(n4038), .B(n4037), .Z(n4040) );
  XOR U4852 ( .A(n4041), .B(n4040), .Z(c[1810]) );
  NAND U4853 ( .A(b[0]), .B(a[788]), .Z(n4044) );
  XNOR U4854 ( .A(sreg[1811]), .B(n4044), .Z(n4046) );
  NANDN U4855 ( .A(n4039), .B(sreg[1810]), .Z(n4043) );
  NAND U4856 ( .A(n4041), .B(n4040), .Z(n4042) );
  NAND U4857 ( .A(n4043), .B(n4042), .Z(n4045) );
  XOR U4858 ( .A(n4046), .B(n4045), .Z(c[1811]) );
  NAND U4859 ( .A(b[0]), .B(a[789]), .Z(n4049) );
  XNOR U4860 ( .A(sreg[1812]), .B(n4049), .Z(n4051) );
  NANDN U4861 ( .A(n4044), .B(sreg[1811]), .Z(n4048) );
  NAND U4862 ( .A(n4046), .B(n4045), .Z(n4047) );
  NAND U4863 ( .A(n4048), .B(n4047), .Z(n4050) );
  XOR U4864 ( .A(n4051), .B(n4050), .Z(c[1812]) );
  NAND U4865 ( .A(b[0]), .B(a[790]), .Z(n4054) );
  XNOR U4866 ( .A(sreg[1813]), .B(n4054), .Z(n4056) );
  NANDN U4867 ( .A(n4049), .B(sreg[1812]), .Z(n4053) );
  NAND U4868 ( .A(n4051), .B(n4050), .Z(n4052) );
  NAND U4869 ( .A(n4053), .B(n4052), .Z(n4055) );
  XOR U4870 ( .A(n4056), .B(n4055), .Z(c[1813]) );
  NAND U4871 ( .A(b[0]), .B(a[791]), .Z(n4059) );
  XNOR U4872 ( .A(sreg[1814]), .B(n4059), .Z(n4061) );
  NANDN U4873 ( .A(n4054), .B(sreg[1813]), .Z(n4058) );
  NAND U4874 ( .A(n4056), .B(n4055), .Z(n4057) );
  NAND U4875 ( .A(n4058), .B(n4057), .Z(n4060) );
  XOR U4876 ( .A(n4061), .B(n4060), .Z(c[1814]) );
  NANDN U4877 ( .A(n4059), .B(sreg[1814]), .Z(n4063) );
  NAND U4878 ( .A(n4061), .B(n4060), .Z(n4062) );
  AND U4879 ( .A(n4063), .B(n4062), .Z(n4066) );
  NAND U4880 ( .A(b[0]), .B(a[792]), .Z(n4064) );
  XNOR U4881 ( .A(sreg[1815]), .B(n4064), .Z(n4065) );
  XNOR U4882 ( .A(n4066), .B(n4065), .Z(c[1815]) );
  NANDN U4883 ( .A(sreg[1815]), .B(n4064), .Z(n4068) );
  NAND U4884 ( .A(n4066), .B(n4065), .Z(n4067) );
  AND U4885 ( .A(n4068), .B(n4067), .Z(n4071) );
  NAND U4886 ( .A(b[0]), .B(a[793]), .Z(n4069) );
  XNOR U4887 ( .A(sreg[1816]), .B(n4069), .Z(n4070) );
  XOR U4888 ( .A(n4071), .B(n4070), .Z(c[1816]) );
  NAND U4889 ( .A(b[0]), .B(a[794]), .Z(n4074) );
  XNOR U4890 ( .A(sreg[1817]), .B(n4074), .Z(n4076) );
  NANDN U4891 ( .A(n4069), .B(sreg[1816]), .Z(n4073) );
  NAND U4892 ( .A(n4071), .B(n4070), .Z(n4072) );
  NAND U4893 ( .A(n4073), .B(n4072), .Z(n4075) );
  XOR U4894 ( .A(n4076), .B(n4075), .Z(c[1817]) );
  NAND U4895 ( .A(b[0]), .B(a[795]), .Z(n4079) );
  XNOR U4896 ( .A(sreg[1818]), .B(n4079), .Z(n4081) );
  NANDN U4897 ( .A(n4074), .B(sreg[1817]), .Z(n4078) );
  NAND U4898 ( .A(n4076), .B(n4075), .Z(n4077) );
  NAND U4899 ( .A(n4078), .B(n4077), .Z(n4080) );
  XOR U4900 ( .A(n4081), .B(n4080), .Z(c[1818]) );
  NAND U4901 ( .A(b[0]), .B(a[796]), .Z(n4084) );
  XNOR U4902 ( .A(sreg[1819]), .B(n4084), .Z(n4086) );
  NANDN U4903 ( .A(n4079), .B(sreg[1818]), .Z(n4083) );
  NAND U4904 ( .A(n4081), .B(n4080), .Z(n4082) );
  NAND U4905 ( .A(n4083), .B(n4082), .Z(n4085) );
  XOR U4906 ( .A(n4086), .B(n4085), .Z(c[1819]) );
  NAND U4907 ( .A(b[0]), .B(a[797]), .Z(n4089) );
  XNOR U4908 ( .A(sreg[1820]), .B(n4089), .Z(n4091) );
  NANDN U4909 ( .A(n4084), .B(sreg[1819]), .Z(n4088) );
  NAND U4910 ( .A(n4086), .B(n4085), .Z(n4087) );
  NAND U4911 ( .A(n4088), .B(n4087), .Z(n4090) );
  XOR U4912 ( .A(n4091), .B(n4090), .Z(c[1820]) );
  NAND U4913 ( .A(b[0]), .B(a[798]), .Z(n4094) );
  XNOR U4914 ( .A(sreg[1821]), .B(n4094), .Z(n4096) );
  NANDN U4915 ( .A(n4089), .B(sreg[1820]), .Z(n4093) );
  NAND U4916 ( .A(n4091), .B(n4090), .Z(n4092) );
  NAND U4917 ( .A(n4093), .B(n4092), .Z(n4095) );
  XOR U4918 ( .A(n4096), .B(n4095), .Z(c[1821]) );
  NAND U4919 ( .A(b[0]), .B(a[799]), .Z(n4099) );
  XNOR U4920 ( .A(sreg[1822]), .B(n4099), .Z(n4101) );
  NANDN U4921 ( .A(n4094), .B(sreg[1821]), .Z(n4098) );
  NAND U4922 ( .A(n4096), .B(n4095), .Z(n4097) );
  NAND U4923 ( .A(n4098), .B(n4097), .Z(n4100) );
  XOR U4924 ( .A(n4101), .B(n4100), .Z(c[1822]) );
  NAND U4925 ( .A(b[0]), .B(a[800]), .Z(n4104) );
  XNOR U4926 ( .A(sreg[1823]), .B(n4104), .Z(n4106) );
  NANDN U4927 ( .A(n4099), .B(sreg[1822]), .Z(n4103) );
  NAND U4928 ( .A(n4101), .B(n4100), .Z(n4102) );
  NAND U4929 ( .A(n4103), .B(n4102), .Z(n4105) );
  XOR U4930 ( .A(n4106), .B(n4105), .Z(c[1823]) );
  NAND U4931 ( .A(b[0]), .B(a[801]), .Z(n4109) );
  XNOR U4932 ( .A(sreg[1824]), .B(n4109), .Z(n4111) );
  NANDN U4933 ( .A(n4104), .B(sreg[1823]), .Z(n4108) );
  NAND U4934 ( .A(n4106), .B(n4105), .Z(n4107) );
  NAND U4935 ( .A(n4108), .B(n4107), .Z(n4110) );
  XOR U4936 ( .A(n4111), .B(n4110), .Z(c[1824]) );
  NAND U4937 ( .A(b[0]), .B(a[802]), .Z(n4114) );
  XNOR U4938 ( .A(sreg[1825]), .B(n4114), .Z(n4116) );
  NANDN U4939 ( .A(n4109), .B(sreg[1824]), .Z(n4113) );
  NAND U4940 ( .A(n4111), .B(n4110), .Z(n4112) );
  NAND U4941 ( .A(n4113), .B(n4112), .Z(n4115) );
  XOR U4942 ( .A(n4116), .B(n4115), .Z(c[1825]) );
  NAND U4943 ( .A(b[0]), .B(a[803]), .Z(n4119) );
  XNOR U4944 ( .A(sreg[1826]), .B(n4119), .Z(n4121) );
  NANDN U4945 ( .A(n4114), .B(sreg[1825]), .Z(n4118) );
  NAND U4946 ( .A(n4116), .B(n4115), .Z(n4117) );
  NAND U4947 ( .A(n4118), .B(n4117), .Z(n4120) );
  XOR U4948 ( .A(n4121), .B(n4120), .Z(c[1826]) );
  NANDN U4949 ( .A(n4119), .B(sreg[1826]), .Z(n4123) );
  NAND U4950 ( .A(n4121), .B(n4120), .Z(n4122) );
  AND U4951 ( .A(n4123), .B(n4122), .Z(n4126) );
  NAND U4952 ( .A(b[0]), .B(a[804]), .Z(n4124) );
  XNOR U4953 ( .A(sreg[1827]), .B(n4124), .Z(n4125) );
  XNOR U4954 ( .A(n4126), .B(n4125), .Z(c[1827]) );
  NAND U4955 ( .A(b[0]), .B(a[805]), .Z(n4129) );
  XNOR U4956 ( .A(sreg[1828]), .B(n4129), .Z(n4131) );
  NANDN U4957 ( .A(sreg[1827]), .B(n4124), .Z(n4128) );
  NAND U4958 ( .A(n4126), .B(n4125), .Z(n4127) );
  AND U4959 ( .A(n4128), .B(n4127), .Z(n4130) );
  XOR U4960 ( .A(n4131), .B(n4130), .Z(c[1828]) );
  NAND U4961 ( .A(b[0]), .B(a[806]), .Z(n4134) );
  XNOR U4962 ( .A(sreg[1829]), .B(n4134), .Z(n4136) );
  NANDN U4963 ( .A(n4129), .B(sreg[1828]), .Z(n4133) );
  NAND U4964 ( .A(n4131), .B(n4130), .Z(n4132) );
  NAND U4965 ( .A(n4133), .B(n4132), .Z(n4135) );
  XOR U4966 ( .A(n4136), .B(n4135), .Z(c[1829]) );
  NAND U4967 ( .A(b[0]), .B(a[807]), .Z(n4139) );
  XNOR U4968 ( .A(sreg[1830]), .B(n4139), .Z(n4141) );
  NANDN U4969 ( .A(n4134), .B(sreg[1829]), .Z(n4138) );
  NAND U4970 ( .A(n4136), .B(n4135), .Z(n4137) );
  AND U4971 ( .A(n4138), .B(n4137), .Z(n4140) );
  XNOR U4972 ( .A(n4141), .B(n4140), .Z(c[1830]) );
  NAND U4973 ( .A(b[0]), .B(a[808]), .Z(n4144) );
  XNOR U4974 ( .A(sreg[1831]), .B(n4144), .Z(n4146) );
  NANDN U4975 ( .A(sreg[1830]), .B(n4139), .Z(n4143) );
  NAND U4976 ( .A(n4141), .B(n4140), .Z(n4142) );
  NAND U4977 ( .A(n4143), .B(n4142), .Z(n4145) );
  XNOR U4978 ( .A(n4146), .B(n4145), .Z(c[1831]) );
  NAND U4979 ( .A(b[0]), .B(a[809]), .Z(n4149) );
  XNOR U4980 ( .A(sreg[1832]), .B(n4149), .Z(n4151) );
  NANDN U4981 ( .A(sreg[1831]), .B(n4144), .Z(n4148) );
  NAND U4982 ( .A(n4146), .B(n4145), .Z(n4147) );
  AND U4983 ( .A(n4148), .B(n4147), .Z(n4150) );
  XOR U4984 ( .A(n4151), .B(n4150), .Z(c[1832]) );
  NANDN U4985 ( .A(n4149), .B(sreg[1832]), .Z(n4153) );
  NAND U4986 ( .A(n4151), .B(n4150), .Z(n4152) );
  AND U4987 ( .A(n4153), .B(n4152), .Z(n4156) );
  NAND U4988 ( .A(b[0]), .B(a[810]), .Z(n4154) );
  XNOR U4989 ( .A(sreg[1833]), .B(n4154), .Z(n4155) );
  XNOR U4990 ( .A(n4156), .B(n4155), .Z(c[1833]) );
  NAND U4991 ( .A(b[0]), .B(a[811]), .Z(n4159) );
  XNOR U4992 ( .A(sreg[1834]), .B(n4159), .Z(n4161) );
  NANDN U4993 ( .A(sreg[1833]), .B(n4154), .Z(n4158) );
  NAND U4994 ( .A(n4156), .B(n4155), .Z(n4157) );
  NAND U4995 ( .A(n4158), .B(n4157), .Z(n4160) );
  XNOR U4996 ( .A(n4161), .B(n4160), .Z(c[1834]) );
  NANDN U4997 ( .A(sreg[1834]), .B(n4159), .Z(n4163) );
  NAND U4998 ( .A(n4161), .B(n4160), .Z(n4162) );
  AND U4999 ( .A(n4163), .B(n4162), .Z(n4166) );
  NAND U5000 ( .A(b[0]), .B(a[812]), .Z(n4164) );
  XNOR U5001 ( .A(sreg[1835]), .B(n4164), .Z(n4165) );
  XOR U5002 ( .A(n4166), .B(n4165), .Z(c[1835]) );
  NAND U5003 ( .A(b[0]), .B(a[813]), .Z(n4169) );
  XNOR U5004 ( .A(sreg[1836]), .B(n4169), .Z(n4171) );
  NANDN U5005 ( .A(n4164), .B(sreg[1835]), .Z(n4168) );
  NAND U5006 ( .A(n4166), .B(n4165), .Z(n4167) );
  NAND U5007 ( .A(n4168), .B(n4167), .Z(n4170) );
  XOR U5008 ( .A(n4171), .B(n4170), .Z(c[1836]) );
  NANDN U5009 ( .A(n4169), .B(sreg[1836]), .Z(n4173) );
  NAND U5010 ( .A(n4171), .B(n4170), .Z(n4172) );
  AND U5011 ( .A(n4173), .B(n4172), .Z(n4176) );
  NAND U5012 ( .A(b[0]), .B(a[814]), .Z(n4174) );
  XNOR U5013 ( .A(sreg[1837]), .B(n4174), .Z(n4175) );
  XNOR U5014 ( .A(n4176), .B(n4175), .Z(c[1837]) );
  NAND U5015 ( .A(b[0]), .B(a[815]), .Z(n4179) );
  XNOR U5016 ( .A(sreg[1838]), .B(n4179), .Z(n4181) );
  NANDN U5017 ( .A(sreg[1837]), .B(n4174), .Z(n4178) );
  NAND U5018 ( .A(n4176), .B(n4175), .Z(n4177) );
  AND U5019 ( .A(n4178), .B(n4177), .Z(n4180) );
  XOR U5020 ( .A(n4181), .B(n4180), .Z(c[1838]) );
  NAND U5021 ( .A(b[0]), .B(a[816]), .Z(n4184) );
  XNOR U5022 ( .A(sreg[1839]), .B(n4184), .Z(n4186) );
  NANDN U5023 ( .A(n4179), .B(sreg[1838]), .Z(n4183) );
  NAND U5024 ( .A(n4181), .B(n4180), .Z(n4182) );
  NAND U5025 ( .A(n4183), .B(n4182), .Z(n4185) );
  XOR U5026 ( .A(n4186), .B(n4185), .Z(c[1839]) );
  NANDN U5027 ( .A(n4184), .B(sreg[1839]), .Z(n4188) );
  NAND U5028 ( .A(n4186), .B(n4185), .Z(n4187) );
  AND U5029 ( .A(n4188), .B(n4187), .Z(n4191) );
  NAND U5030 ( .A(b[0]), .B(a[817]), .Z(n4189) );
  XNOR U5031 ( .A(sreg[1840]), .B(n4189), .Z(n4190) );
  XNOR U5032 ( .A(n4191), .B(n4190), .Z(c[1840]) );
  NAND U5033 ( .A(b[0]), .B(a[818]), .Z(n4194) );
  XNOR U5034 ( .A(sreg[1841]), .B(n4194), .Z(n4196) );
  NANDN U5035 ( .A(sreg[1840]), .B(n4189), .Z(n4193) );
  NAND U5036 ( .A(n4191), .B(n4190), .Z(n4192) );
  AND U5037 ( .A(n4193), .B(n4192), .Z(n4195) );
  XOR U5038 ( .A(n4196), .B(n4195), .Z(c[1841]) );
  NAND U5039 ( .A(b[0]), .B(a[819]), .Z(n4199) );
  XNOR U5040 ( .A(sreg[1842]), .B(n4199), .Z(n4201) );
  NANDN U5041 ( .A(n4194), .B(sreg[1841]), .Z(n4198) );
  NAND U5042 ( .A(n4196), .B(n4195), .Z(n4197) );
  NAND U5043 ( .A(n4198), .B(n4197), .Z(n4200) );
  XOR U5044 ( .A(n4201), .B(n4200), .Z(c[1842]) );
  NAND U5045 ( .A(b[0]), .B(a[820]), .Z(n4204) );
  XNOR U5046 ( .A(sreg[1843]), .B(n4204), .Z(n4206) );
  NANDN U5047 ( .A(n4199), .B(sreg[1842]), .Z(n4203) );
  NAND U5048 ( .A(n4201), .B(n4200), .Z(n4202) );
  AND U5049 ( .A(n4203), .B(n4202), .Z(n4205) );
  XNOR U5050 ( .A(n4206), .B(n4205), .Z(c[1843]) );
  NANDN U5051 ( .A(sreg[1843]), .B(n4204), .Z(n4208) );
  NAND U5052 ( .A(n4206), .B(n4205), .Z(n4207) );
  AND U5053 ( .A(n4208), .B(n4207), .Z(n4211) );
  NAND U5054 ( .A(b[0]), .B(a[821]), .Z(n4209) );
  XNOR U5055 ( .A(sreg[1844]), .B(n4209), .Z(n4210) );
  XOR U5056 ( .A(n4211), .B(n4210), .Z(c[1844]) );
  NAND U5057 ( .A(b[0]), .B(a[822]), .Z(n4214) );
  XNOR U5058 ( .A(sreg[1845]), .B(n4214), .Z(n4216) );
  NANDN U5059 ( .A(n4209), .B(sreg[1844]), .Z(n4213) );
  NAND U5060 ( .A(n4211), .B(n4210), .Z(n4212) );
  NAND U5061 ( .A(n4213), .B(n4212), .Z(n4215) );
  XOR U5062 ( .A(n4216), .B(n4215), .Z(c[1845]) );
  NAND U5063 ( .A(b[0]), .B(a[823]), .Z(n4219) );
  XNOR U5064 ( .A(sreg[1846]), .B(n4219), .Z(n4221) );
  NANDN U5065 ( .A(n4214), .B(sreg[1845]), .Z(n4218) );
  NAND U5066 ( .A(n4216), .B(n4215), .Z(n4217) );
  AND U5067 ( .A(n4218), .B(n4217), .Z(n4220) );
  XNOR U5068 ( .A(n4221), .B(n4220), .Z(c[1846]) );
  NAND U5069 ( .A(b[0]), .B(a[824]), .Z(n4224) );
  XNOR U5070 ( .A(sreg[1847]), .B(n4224), .Z(n4226) );
  NANDN U5071 ( .A(sreg[1846]), .B(n4219), .Z(n4223) );
  NAND U5072 ( .A(n4221), .B(n4220), .Z(n4222) );
  AND U5073 ( .A(n4223), .B(n4222), .Z(n4225) );
  XOR U5074 ( .A(n4226), .B(n4225), .Z(c[1847]) );
  NAND U5075 ( .A(b[0]), .B(a[825]), .Z(n4229) );
  XNOR U5076 ( .A(sreg[1848]), .B(n4229), .Z(n4231) );
  NANDN U5077 ( .A(n4224), .B(sreg[1847]), .Z(n4228) );
  NAND U5078 ( .A(n4226), .B(n4225), .Z(n4227) );
  NAND U5079 ( .A(n4228), .B(n4227), .Z(n4230) );
  XOR U5080 ( .A(n4231), .B(n4230), .Z(c[1848]) );
  NAND U5081 ( .A(b[0]), .B(a[826]), .Z(n4234) );
  XNOR U5082 ( .A(sreg[1849]), .B(n4234), .Z(n4236) );
  NANDN U5083 ( .A(n4229), .B(sreg[1848]), .Z(n4233) );
  NAND U5084 ( .A(n4231), .B(n4230), .Z(n4232) );
  NAND U5085 ( .A(n4233), .B(n4232), .Z(n4235) );
  XOR U5086 ( .A(n4236), .B(n4235), .Z(c[1849]) );
  NAND U5087 ( .A(b[0]), .B(a[827]), .Z(n4240) );
  NANDN U5088 ( .A(n4234), .B(sreg[1849]), .Z(n4238) );
  NAND U5089 ( .A(n4236), .B(n4235), .Z(n4237) );
  AND U5090 ( .A(n4238), .B(n4237), .Z(n4241) );
  XNOR U5091 ( .A(n4241), .B(sreg[1850]), .Z(n4239) );
  XNOR U5092 ( .A(n4240), .B(n4239), .Z(c[1850]) );
  NAND U5093 ( .A(b[0]), .B(a[828]), .Z(n4242) );
  XNOR U5094 ( .A(sreg[1851]), .B(n4242), .Z(n4244) );
  XOR U5095 ( .A(n4244), .B(n4243), .Z(c[1851]) );
  NAND U5096 ( .A(b[0]), .B(a[829]), .Z(n4247) );
  XNOR U5097 ( .A(sreg[1852]), .B(n4247), .Z(n4249) );
  NANDN U5098 ( .A(n4242), .B(sreg[1851]), .Z(n4246) );
  NAND U5099 ( .A(n4244), .B(n4243), .Z(n4245) );
  NAND U5100 ( .A(n4246), .B(n4245), .Z(n4248) );
  XOR U5101 ( .A(n4249), .B(n4248), .Z(c[1852]) );
  NAND U5102 ( .A(b[0]), .B(a[830]), .Z(n4252) );
  XNOR U5103 ( .A(sreg[1853]), .B(n4252), .Z(n4254) );
  NANDN U5104 ( .A(n4247), .B(sreg[1852]), .Z(n4251) );
  NAND U5105 ( .A(n4249), .B(n4248), .Z(n4250) );
  NAND U5106 ( .A(n4251), .B(n4250), .Z(n4253) );
  XOR U5107 ( .A(n4254), .B(n4253), .Z(c[1853]) );
  NAND U5108 ( .A(b[0]), .B(a[831]), .Z(n4257) );
  XNOR U5109 ( .A(sreg[1854]), .B(n4257), .Z(n4259) );
  NANDN U5110 ( .A(n4252), .B(sreg[1853]), .Z(n4256) );
  NAND U5111 ( .A(n4254), .B(n4253), .Z(n4255) );
  NAND U5112 ( .A(n4256), .B(n4255), .Z(n4258) );
  XOR U5113 ( .A(n4259), .B(n4258), .Z(c[1854]) );
  NANDN U5114 ( .A(n4257), .B(sreg[1854]), .Z(n4261) );
  NAND U5115 ( .A(n4259), .B(n4258), .Z(n4260) );
  AND U5116 ( .A(n4261), .B(n4260), .Z(n4264) );
  NAND U5117 ( .A(b[0]), .B(a[832]), .Z(n4262) );
  XNOR U5118 ( .A(sreg[1855]), .B(n4262), .Z(n4263) );
  XNOR U5119 ( .A(n4264), .B(n4263), .Z(c[1855]) );
  NAND U5120 ( .A(b[0]), .B(a[833]), .Z(n4267) );
  XNOR U5121 ( .A(sreg[1856]), .B(n4267), .Z(n4269) );
  NANDN U5122 ( .A(sreg[1855]), .B(n4262), .Z(n4266) );
  NAND U5123 ( .A(n4264), .B(n4263), .Z(n4265) );
  NAND U5124 ( .A(n4266), .B(n4265), .Z(n4268) );
  XNOR U5125 ( .A(n4269), .B(n4268), .Z(c[1856]) );
  NAND U5126 ( .A(b[0]), .B(a[834]), .Z(n4272) );
  XNOR U5127 ( .A(sreg[1857]), .B(n4272), .Z(n4274) );
  NANDN U5128 ( .A(sreg[1856]), .B(n4267), .Z(n4271) );
  NAND U5129 ( .A(n4269), .B(n4268), .Z(n4270) );
  NAND U5130 ( .A(n4271), .B(n4270), .Z(n4273) );
  XNOR U5131 ( .A(n4274), .B(n4273), .Z(c[1857]) );
  NAND U5132 ( .A(b[0]), .B(a[835]), .Z(n4277) );
  XNOR U5133 ( .A(sreg[1858]), .B(n4277), .Z(n4279) );
  NANDN U5134 ( .A(sreg[1857]), .B(n4272), .Z(n4276) );
  NAND U5135 ( .A(n4274), .B(n4273), .Z(n4275) );
  NAND U5136 ( .A(n4276), .B(n4275), .Z(n4278) );
  XNOR U5137 ( .A(n4279), .B(n4278), .Z(c[1858]) );
  NAND U5138 ( .A(b[0]), .B(a[836]), .Z(n4282) );
  XNOR U5139 ( .A(sreg[1859]), .B(n4282), .Z(n4284) );
  NANDN U5140 ( .A(sreg[1858]), .B(n4277), .Z(n4281) );
  NAND U5141 ( .A(n4279), .B(n4278), .Z(n4280) );
  NAND U5142 ( .A(n4281), .B(n4280), .Z(n4283) );
  XNOR U5143 ( .A(n4284), .B(n4283), .Z(c[1859]) );
  NAND U5144 ( .A(b[0]), .B(a[837]), .Z(n4287) );
  XNOR U5145 ( .A(sreg[1860]), .B(n4287), .Z(n4289) );
  NANDN U5146 ( .A(sreg[1859]), .B(n4282), .Z(n4286) );
  NAND U5147 ( .A(n4284), .B(n4283), .Z(n4285) );
  NAND U5148 ( .A(n4286), .B(n4285), .Z(n4288) );
  XNOR U5149 ( .A(n4289), .B(n4288), .Z(c[1860]) );
  NAND U5150 ( .A(b[0]), .B(a[838]), .Z(n4292) );
  XNOR U5151 ( .A(sreg[1861]), .B(n4292), .Z(n4294) );
  NANDN U5152 ( .A(sreg[1860]), .B(n4287), .Z(n4291) );
  NAND U5153 ( .A(n4289), .B(n4288), .Z(n4290) );
  NAND U5154 ( .A(n4291), .B(n4290), .Z(n4293) );
  XNOR U5155 ( .A(n4294), .B(n4293), .Z(c[1861]) );
  NAND U5156 ( .A(b[0]), .B(a[839]), .Z(n4297) );
  XNOR U5157 ( .A(sreg[1862]), .B(n4297), .Z(n4299) );
  NANDN U5158 ( .A(sreg[1861]), .B(n4292), .Z(n4296) );
  NAND U5159 ( .A(n4294), .B(n4293), .Z(n4295) );
  NAND U5160 ( .A(n4296), .B(n4295), .Z(n4298) );
  XNOR U5161 ( .A(n4299), .B(n4298), .Z(c[1862]) );
  NAND U5162 ( .A(b[0]), .B(a[840]), .Z(n4302) );
  XNOR U5163 ( .A(sreg[1863]), .B(n4302), .Z(n4304) );
  NANDN U5164 ( .A(sreg[1862]), .B(n4297), .Z(n4301) );
  NAND U5165 ( .A(n4299), .B(n4298), .Z(n4300) );
  NAND U5166 ( .A(n4301), .B(n4300), .Z(n4303) );
  XNOR U5167 ( .A(n4304), .B(n4303), .Z(c[1863]) );
  NAND U5168 ( .A(b[0]), .B(a[841]), .Z(n4307) );
  XNOR U5169 ( .A(sreg[1864]), .B(n4307), .Z(n4309) );
  NANDN U5170 ( .A(sreg[1863]), .B(n4302), .Z(n4306) );
  NAND U5171 ( .A(n4304), .B(n4303), .Z(n4305) );
  NAND U5172 ( .A(n4306), .B(n4305), .Z(n4308) );
  XNOR U5173 ( .A(n4309), .B(n4308), .Z(c[1864]) );
  NAND U5174 ( .A(b[0]), .B(a[842]), .Z(n4312) );
  XNOR U5175 ( .A(sreg[1865]), .B(n4312), .Z(n4314) );
  NANDN U5176 ( .A(sreg[1864]), .B(n4307), .Z(n4311) );
  NAND U5177 ( .A(n4309), .B(n4308), .Z(n4310) );
  NAND U5178 ( .A(n4311), .B(n4310), .Z(n4313) );
  XNOR U5179 ( .A(n4314), .B(n4313), .Z(c[1865]) );
  NAND U5180 ( .A(b[0]), .B(a[843]), .Z(n4317) );
  XNOR U5181 ( .A(sreg[1866]), .B(n4317), .Z(n4319) );
  NANDN U5182 ( .A(sreg[1865]), .B(n4312), .Z(n4316) );
  NAND U5183 ( .A(n4314), .B(n4313), .Z(n4315) );
  NAND U5184 ( .A(n4316), .B(n4315), .Z(n4318) );
  XNOR U5185 ( .A(n4319), .B(n4318), .Z(c[1866]) );
  NAND U5186 ( .A(b[0]), .B(a[844]), .Z(n4322) );
  XNOR U5187 ( .A(sreg[1867]), .B(n4322), .Z(n4324) );
  NANDN U5188 ( .A(sreg[1866]), .B(n4317), .Z(n4321) );
  NAND U5189 ( .A(n4319), .B(n4318), .Z(n4320) );
  NAND U5190 ( .A(n4321), .B(n4320), .Z(n4323) );
  XNOR U5191 ( .A(n4324), .B(n4323), .Z(c[1867]) );
  NAND U5192 ( .A(b[0]), .B(a[845]), .Z(n4327) );
  XNOR U5193 ( .A(sreg[1868]), .B(n4327), .Z(n4329) );
  NANDN U5194 ( .A(sreg[1867]), .B(n4322), .Z(n4326) );
  NAND U5195 ( .A(n4324), .B(n4323), .Z(n4325) );
  NAND U5196 ( .A(n4326), .B(n4325), .Z(n4328) );
  XNOR U5197 ( .A(n4329), .B(n4328), .Z(c[1868]) );
  NAND U5198 ( .A(b[0]), .B(a[846]), .Z(n4332) );
  XNOR U5199 ( .A(sreg[1869]), .B(n4332), .Z(n4334) );
  NANDN U5200 ( .A(sreg[1868]), .B(n4327), .Z(n4331) );
  NAND U5201 ( .A(n4329), .B(n4328), .Z(n4330) );
  NAND U5202 ( .A(n4331), .B(n4330), .Z(n4333) );
  XNOR U5203 ( .A(n4334), .B(n4333), .Z(c[1869]) );
  NAND U5204 ( .A(b[0]), .B(a[847]), .Z(n4337) );
  XNOR U5205 ( .A(sreg[1870]), .B(n4337), .Z(n4339) );
  NANDN U5206 ( .A(sreg[1869]), .B(n4332), .Z(n4336) );
  NAND U5207 ( .A(n4334), .B(n4333), .Z(n4335) );
  NAND U5208 ( .A(n4336), .B(n4335), .Z(n4338) );
  XNOR U5209 ( .A(n4339), .B(n4338), .Z(c[1870]) );
  NAND U5210 ( .A(b[0]), .B(a[848]), .Z(n4344) );
  NANDN U5211 ( .A(sreg[1870]), .B(n4337), .Z(n4341) );
  NAND U5212 ( .A(n4339), .B(n4338), .Z(n4340) );
  AND U5213 ( .A(n4341), .B(n4340), .Z(n4343) );
  XOR U5214 ( .A(sreg[1871]), .B(n4343), .Z(n4342) );
  XNOR U5215 ( .A(n4344), .B(n4342), .Z(c[1871]) );
  NAND U5216 ( .A(b[0]), .B(a[849]), .Z(n4345) );
  XNOR U5217 ( .A(sreg[1872]), .B(n4345), .Z(n4346) );
  XOR U5218 ( .A(n4347), .B(n4346), .Z(c[1872]) );
  NAND U5219 ( .A(b[0]), .B(a[850]), .Z(n4350) );
  XNOR U5220 ( .A(sreg[1873]), .B(n4350), .Z(n4352) );
  NANDN U5221 ( .A(n4345), .B(sreg[1872]), .Z(n4349) );
  NAND U5222 ( .A(n4347), .B(n4346), .Z(n4348) );
  NAND U5223 ( .A(n4349), .B(n4348), .Z(n4351) );
  XOR U5224 ( .A(n4352), .B(n4351), .Z(c[1873]) );
  NAND U5225 ( .A(b[0]), .B(a[851]), .Z(n4355) );
  XNOR U5226 ( .A(sreg[1874]), .B(n4355), .Z(n4357) );
  NANDN U5227 ( .A(n4350), .B(sreg[1873]), .Z(n4354) );
  NAND U5228 ( .A(n4352), .B(n4351), .Z(n4353) );
  NAND U5229 ( .A(n4354), .B(n4353), .Z(n4356) );
  XOR U5230 ( .A(n4357), .B(n4356), .Z(c[1874]) );
  NAND U5231 ( .A(b[0]), .B(a[852]), .Z(n4360) );
  XNOR U5232 ( .A(sreg[1875]), .B(n4360), .Z(n4362) );
  NANDN U5233 ( .A(n4355), .B(sreg[1874]), .Z(n4359) );
  NAND U5234 ( .A(n4357), .B(n4356), .Z(n4358) );
  NAND U5235 ( .A(n4359), .B(n4358), .Z(n4361) );
  XOR U5236 ( .A(n4362), .B(n4361), .Z(c[1875]) );
  NAND U5237 ( .A(b[0]), .B(a[853]), .Z(n4365) );
  XNOR U5238 ( .A(sreg[1876]), .B(n4365), .Z(n4367) );
  NANDN U5239 ( .A(n4360), .B(sreg[1875]), .Z(n4364) );
  NAND U5240 ( .A(n4362), .B(n4361), .Z(n4363) );
  NAND U5241 ( .A(n4364), .B(n4363), .Z(n4366) );
  XOR U5242 ( .A(n4367), .B(n4366), .Z(c[1876]) );
  NANDN U5243 ( .A(n4365), .B(sreg[1876]), .Z(n4369) );
  NAND U5244 ( .A(n4367), .B(n4366), .Z(n4368) );
  AND U5245 ( .A(n4369), .B(n4368), .Z(n4372) );
  NAND U5246 ( .A(b[0]), .B(a[854]), .Z(n4370) );
  XNOR U5247 ( .A(sreg[1877]), .B(n4370), .Z(n4371) );
  XNOR U5248 ( .A(n4372), .B(n4371), .Z(c[1877]) );
  NAND U5249 ( .A(b[0]), .B(a[855]), .Z(n4375) );
  XNOR U5250 ( .A(sreg[1878]), .B(n4375), .Z(n4377) );
  NANDN U5251 ( .A(sreg[1877]), .B(n4370), .Z(n4374) );
  NAND U5252 ( .A(n4372), .B(n4371), .Z(n4373) );
  AND U5253 ( .A(n4374), .B(n4373), .Z(n4376) );
  XOR U5254 ( .A(n4377), .B(n4376), .Z(c[1878]) );
  NAND U5255 ( .A(b[0]), .B(a[856]), .Z(n4380) );
  XNOR U5256 ( .A(sreg[1879]), .B(n4380), .Z(n4382) );
  NANDN U5257 ( .A(n4375), .B(sreg[1878]), .Z(n4379) );
  NAND U5258 ( .A(n4377), .B(n4376), .Z(n4378) );
  NAND U5259 ( .A(n4379), .B(n4378), .Z(n4381) );
  XOR U5260 ( .A(n4382), .B(n4381), .Z(c[1879]) );
  NAND U5261 ( .A(b[0]), .B(a[857]), .Z(n4385) );
  XNOR U5262 ( .A(sreg[1880]), .B(n4385), .Z(n4387) );
  NANDN U5263 ( .A(n4380), .B(sreg[1879]), .Z(n4384) );
  NAND U5264 ( .A(n4382), .B(n4381), .Z(n4383) );
  AND U5265 ( .A(n4384), .B(n4383), .Z(n4386) );
  XNOR U5266 ( .A(n4387), .B(n4386), .Z(c[1880]) );
  NANDN U5267 ( .A(sreg[1880]), .B(n4385), .Z(n4389) );
  NAND U5268 ( .A(n4387), .B(n4386), .Z(n4388) );
  AND U5269 ( .A(n4389), .B(n4388), .Z(n4392) );
  NAND U5270 ( .A(b[0]), .B(a[858]), .Z(n4390) );
  XNOR U5271 ( .A(sreg[1881]), .B(n4390), .Z(n4391) );
  XOR U5272 ( .A(n4392), .B(n4391), .Z(c[1881]) );
  NAND U5273 ( .A(b[0]), .B(a[859]), .Z(n4395) );
  XNOR U5274 ( .A(sreg[1882]), .B(n4395), .Z(n4397) );
  NANDN U5275 ( .A(n4390), .B(sreg[1881]), .Z(n4394) );
  NAND U5276 ( .A(n4392), .B(n4391), .Z(n4393) );
  NAND U5277 ( .A(n4394), .B(n4393), .Z(n4396) );
  XOR U5278 ( .A(n4397), .B(n4396), .Z(c[1882]) );
  NANDN U5279 ( .A(n4395), .B(sreg[1882]), .Z(n4399) );
  NAND U5280 ( .A(n4397), .B(n4396), .Z(n4398) );
  AND U5281 ( .A(n4399), .B(n4398), .Z(n4402) );
  NAND U5282 ( .A(b[0]), .B(a[860]), .Z(n4400) );
  XNOR U5283 ( .A(sreg[1883]), .B(n4400), .Z(n4401) );
  XNOR U5284 ( .A(n4402), .B(n4401), .Z(c[1883]) );
  NAND U5285 ( .A(b[0]), .B(a[861]), .Z(n4405) );
  XNOR U5286 ( .A(sreg[1884]), .B(n4405), .Z(n4407) );
  NANDN U5287 ( .A(sreg[1883]), .B(n4400), .Z(n4404) );
  NAND U5288 ( .A(n4402), .B(n4401), .Z(n4403) );
  AND U5289 ( .A(n4404), .B(n4403), .Z(n4406) );
  XOR U5290 ( .A(n4407), .B(n4406), .Z(c[1884]) );
  NAND U5291 ( .A(b[0]), .B(a[862]), .Z(n4410) );
  XNOR U5292 ( .A(sreg[1885]), .B(n4410), .Z(n4412) );
  NANDN U5293 ( .A(n4405), .B(sreg[1884]), .Z(n4409) );
  NAND U5294 ( .A(n4407), .B(n4406), .Z(n4408) );
  NAND U5295 ( .A(n4409), .B(n4408), .Z(n4411) );
  XOR U5296 ( .A(n4412), .B(n4411), .Z(c[1885]) );
  NANDN U5297 ( .A(n4410), .B(sreg[1885]), .Z(n4414) );
  NAND U5298 ( .A(n4412), .B(n4411), .Z(n4413) );
  AND U5299 ( .A(n4414), .B(n4413), .Z(n4417) );
  NAND U5300 ( .A(b[0]), .B(a[863]), .Z(n4415) );
  XNOR U5301 ( .A(sreg[1886]), .B(n4415), .Z(n4416) );
  XNOR U5302 ( .A(n4417), .B(n4416), .Z(c[1886]) );
  NAND U5303 ( .A(b[0]), .B(a[864]), .Z(n4420) );
  XNOR U5304 ( .A(sreg[1887]), .B(n4420), .Z(n4422) );
  NANDN U5305 ( .A(sreg[1886]), .B(n4415), .Z(n4419) );
  NAND U5306 ( .A(n4417), .B(n4416), .Z(n4418) );
  AND U5307 ( .A(n4419), .B(n4418), .Z(n4421) );
  XOR U5308 ( .A(n4422), .B(n4421), .Z(c[1887]) );
  NAND U5309 ( .A(b[0]), .B(a[865]), .Z(n4425) );
  XNOR U5310 ( .A(sreg[1888]), .B(n4425), .Z(n4427) );
  NANDN U5311 ( .A(n4420), .B(sreg[1887]), .Z(n4424) );
  NAND U5312 ( .A(n4422), .B(n4421), .Z(n4423) );
  NAND U5313 ( .A(n4424), .B(n4423), .Z(n4426) );
  XOR U5314 ( .A(n4427), .B(n4426), .Z(c[1888]) );
  NANDN U5315 ( .A(n4425), .B(sreg[1888]), .Z(n4429) );
  NAND U5316 ( .A(n4427), .B(n4426), .Z(n4428) );
  AND U5317 ( .A(n4429), .B(n4428), .Z(n4432) );
  NAND U5318 ( .A(b[0]), .B(a[866]), .Z(n4430) );
  XNOR U5319 ( .A(sreg[1889]), .B(n4430), .Z(n4431) );
  XNOR U5320 ( .A(n4432), .B(n4431), .Z(c[1889]) );
  NAND U5321 ( .A(b[0]), .B(a[867]), .Z(n4435) );
  XNOR U5322 ( .A(sreg[1890]), .B(n4435), .Z(n4437) );
  NANDN U5323 ( .A(sreg[1889]), .B(n4430), .Z(n4434) );
  NAND U5324 ( .A(n4432), .B(n4431), .Z(n4433) );
  NAND U5325 ( .A(n4434), .B(n4433), .Z(n4436) );
  XNOR U5326 ( .A(n4437), .B(n4436), .Z(c[1890]) );
  NANDN U5327 ( .A(sreg[1890]), .B(n4435), .Z(n4439) );
  NAND U5328 ( .A(n4437), .B(n4436), .Z(n4438) );
  AND U5329 ( .A(n4439), .B(n4438), .Z(n4442) );
  NAND U5330 ( .A(b[0]), .B(a[868]), .Z(n4440) );
  XNOR U5331 ( .A(sreg[1891]), .B(n4440), .Z(n4441) );
  XOR U5332 ( .A(n4442), .B(n4441), .Z(c[1891]) );
  NAND U5333 ( .A(b[0]), .B(a[869]), .Z(n4445) );
  XNOR U5334 ( .A(sreg[1892]), .B(n4445), .Z(n4447) );
  NANDN U5335 ( .A(n4440), .B(sreg[1891]), .Z(n4444) );
  NAND U5336 ( .A(n4442), .B(n4441), .Z(n4443) );
  AND U5337 ( .A(n4444), .B(n4443), .Z(n4446) );
  XNOR U5338 ( .A(n4447), .B(n4446), .Z(c[1892]) );
  NAND U5339 ( .A(b[0]), .B(a[870]), .Z(n4450) );
  XNOR U5340 ( .A(sreg[1893]), .B(n4450), .Z(n4452) );
  NANDN U5341 ( .A(sreg[1892]), .B(n4445), .Z(n4449) );
  NAND U5342 ( .A(n4447), .B(n4446), .Z(n4448) );
  NAND U5343 ( .A(n4449), .B(n4448), .Z(n4451) );
  XNOR U5344 ( .A(n4452), .B(n4451), .Z(c[1893]) );
  NAND U5345 ( .A(b[0]), .B(a[871]), .Z(n4455) );
  XNOR U5346 ( .A(sreg[1894]), .B(n4455), .Z(n4457) );
  NANDN U5347 ( .A(sreg[1893]), .B(n4450), .Z(n4454) );
  NAND U5348 ( .A(n4452), .B(n4451), .Z(n4453) );
  AND U5349 ( .A(n4454), .B(n4453), .Z(n4456) );
  XOR U5350 ( .A(n4457), .B(n4456), .Z(c[1894]) );
  NAND U5351 ( .A(b[0]), .B(a[872]), .Z(n4460) );
  XNOR U5352 ( .A(sreg[1895]), .B(n4460), .Z(n4462) );
  NANDN U5353 ( .A(n4455), .B(sreg[1894]), .Z(n4459) );
  NAND U5354 ( .A(n4457), .B(n4456), .Z(n4458) );
  AND U5355 ( .A(n4459), .B(n4458), .Z(n4461) );
  XNOR U5356 ( .A(n4462), .B(n4461), .Z(c[1895]) );
  NAND U5357 ( .A(b[0]), .B(a[873]), .Z(n4465) );
  XNOR U5358 ( .A(sreg[1896]), .B(n4465), .Z(n4467) );
  NANDN U5359 ( .A(sreg[1895]), .B(n4460), .Z(n4464) );
  NAND U5360 ( .A(n4462), .B(n4461), .Z(n4463) );
  NAND U5361 ( .A(n4464), .B(n4463), .Z(n4466) );
  XNOR U5362 ( .A(n4467), .B(n4466), .Z(c[1896]) );
  NAND U5363 ( .A(b[0]), .B(a[874]), .Z(n4470) );
  XNOR U5364 ( .A(sreg[1897]), .B(n4470), .Z(n4472) );
  NANDN U5365 ( .A(sreg[1896]), .B(n4465), .Z(n4469) );
  NAND U5366 ( .A(n4467), .B(n4466), .Z(n4468) );
  AND U5367 ( .A(n4469), .B(n4468), .Z(n4471) );
  XOR U5368 ( .A(n4472), .B(n4471), .Z(c[1897]) );
  NAND U5369 ( .A(b[0]), .B(a[875]), .Z(n4475) );
  XNOR U5370 ( .A(sreg[1898]), .B(n4475), .Z(n4477) );
  NANDN U5371 ( .A(n4470), .B(sreg[1897]), .Z(n4474) );
  NAND U5372 ( .A(n4472), .B(n4471), .Z(n4473) );
  NAND U5373 ( .A(n4474), .B(n4473), .Z(n4476) );
  XOR U5374 ( .A(n4477), .B(n4476), .Z(c[1898]) );
  NANDN U5375 ( .A(n4475), .B(sreg[1898]), .Z(n4479) );
  NAND U5376 ( .A(n4477), .B(n4476), .Z(n4478) );
  AND U5377 ( .A(n4479), .B(n4478), .Z(n4482) );
  NAND U5378 ( .A(b[0]), .B(a[876]), .Z(n4480) );
  XNOR U5379 ( .A(sreg[1899]), .B(n4480), .Z(n4481) );
  XNOR U5380 ( .A(n4482), .B(n4481), .Z(c[1899]) );
  NANDN U5381 ( .A(sreg[1899]), .B(n4480), .Z(n4484) );
  NAND U5382 ( .A(n4482), .B(n4481), .Z(n4483) );
  AND U5383 ( .A(n4484), .B(n4483), .Z(n4487) );
  NAND U5384 ( .A(b[0]), .B(a[877]), .Z(n4485) );
  XNOR U5385 ( .A(sreg[1900]), .B(n4485), .Z(n4486) );
  XOR U5386 ( .A(n4487), .B(n4486), .Z(c[1900]) );
  NANDN U5387 ( .A(n4485), .B(sreg[1900]), .Z(n4489) );
  NAND U5388 ( .A(n4487), .B(n4486), .Z(n4488) );
  AND U5389 ( .A(n4489), .B(n4488), .Z(n4491) );
  AND U5390 ( .A(b[0]), .B(a[878]), .Z(n4492) );
  XNOR U5391 ( .A(sreg[1901]), .B(n4492), .Z(n4490) );
  XOR U5392 ( .A(n4491), .B(n4490), .Z(c[1901]) );
  NAND U5393 ( .A(b[0]), .B(a[879]), .Z(n4493) );
  XNOR U5394 ( .A(sreg[1902]), .B(n4493), .Z(n4495) );
  XOR U5395 ( .A(n4495), .B(n4494), .Z(c[1902]) );
  NAND U5396 ( .A(b[0]), .B(a[880]), .Z(n4500) );
  NANDN U5397 ( .A(n4493), .B(sreg[1902]), .Z(n4497) );
  NAND U5398 ( .A(n4495), .B(n4494), .Z(n4496) );
  NAND U5399 ( .A(n4497), .B(n4496), .Z(n4499) );
  XOR U5400 ( .A(n4499), .B(sreg[1903]), .Z(n4498) );
  XNOR U5401 ( .A(n4500), .B(n4498), .Z(c[1903]) );
  NAND U5402 ( .A(b[0]), .B(a[881]), .Z(n4501) );
  XNOR U5403 ( .A(sreg[1904]), .B(n4501), .Z(n4502) );
  XNOR U5404 ( .A(n4503), .B(n4502), .Z(c[1904]) );
  NAND U5405 ( .A(b[0]), .B(a[882]), .Z(n4506) );
  XNOR U5406 ( .A(sreg[1905]), .B(n4506), .Z(n4508) );
  NANDN U5407 ( .A(n4501), .B(sreg[1904]), .Z(n4505) );
  NANDN U5408 ( .A(n4503), .B(n4502), .Z(n4504) );
  NAND U5409 ( .A(n4505), .B(n4504), .Z(n4507) );
  XOR U5410 ( .A(n4508), .B(n4507), .Z(c[1905]) );
  NAND U5411 ( .A(b[0]), .B(a[883]), .Z(n4511) );
  XNOR U5412 ( .A(sreg[1906]), .B(n4511), .Z(n4513) );
  NANDN U5413 ( .A(n4506), .B(sreg[1905]), .Z(n4510) );
  NAND U5414 ( .A(n4508), .B(n4507), .Z(n4509) );
  AND U5415 ( .A(n4510), .B(n4509), .Z(n4512) );
  XNOR U5416 ( .A(n4513), .B(n4512), .Z(c[1906]) );
  NANDN U5417 ( .A(sreg[1906]), .B(n4511), .Z(n4515) );
  NAND U5418 ( .A(n4513), .B(n4512), .Z(n4514) );
  AND U5419 ( .A(n4515), .B(n4514), .Z(n4518) );
  NAND U5420 ( .A(b[0]), .B(a[884]), .Z(n4516) );
  XNOR U5421 ( .A(sreg[1907]), .B(n4516), .Z(n4517) );
  XOR U5422 ( .A(n4518), .B(n4517), .Z(c[1907]) );
  NAND U5423 ( .A(b[0]), .B(a[885]), .Z(n4521) );
  XNOR U5424 ( .A(sreg[1908]), .B(n4521), .Z(n4523) );
  NANDN U5425 ( .A(n4516), .B(sreg[1907]), .Z(n4520) );
  NAND U5426 ( .A(n4518), .B(n4517), .Z(n4519) );
  NAND U5427 ( .A(n4520), .B(n4519), .Z(n4522) );
  XOR U5428 ( .A(n4523), .B(n4522), .Z(c[1908]) );
  NAND U5429 ( .A(b[0]), .B(a[886]), .Z(n4526) );
  XNOR U5430 ( .A(sreg[1909]), .B(n4526), .Z(n4528) );
  NANDN U5431 ( .A(n4521), .B(sreg[1908]), .Z(n4525) );
  NAND U5432 ( .A(n4523), .B(n4522), .Z(n4524) );
  NAND U5433 ( .A(n4525), .B(n4524), .Z(n4527) );
  XOR U5434 ( .A(n4528), .B(n4527), .Z(c[1909]) );
  NAND U5435 ( .A(b[0]), .B(a[887]), .Z(n4531) );
  XNOR U5436 ( .A(sreg[1910]), .B(n4531), .Z(n4533) );
  NANDN U5437 ( .A(n4526), .B(sreg[1909]), .Z(n4530) );
  NAND U5438 ( .A(n4528), .B(n4527), .Z(n4529) );
  NAND U5439 ( .A(n4530), .B(n4529), .Z(n4532) );
  XOR U5440 ( .A(n4533), .B(n4532), .Z(c[1910]) );
  NAND U5441 ( .A(b[0]), .B(a[888]), .Z(n4536) );
  XNOR U5442 ( .A(sreg[1911]), .B(n4536), .Z(n4538) );
  NANDN U5443 ( .A(n4531), .B(sreg[1910]), .Z(n4535) );
  NAND U5444 ( .A(n4533), .B(n4532), .Z(n4534) );
  NAND U5445 ( .A(n4535), .B(n4534), .Z(n4537) );
  XOR U5446 ( .A(n4538), .B(n4537), .Z(c[1911]) );
  NAND U5447 ( .A(b[0]), .B(a[889]), .Z(n4541) );
  XNOR U5448 ( .A(sreg[1912]), .B(n4541), .Z(n4543) );
  NANDN U5449 ( .A(n4536), .B(sreg[1911]), .Z(n4540) );
  NAND U5450 ( .A(n4538), .B(n4537), .Z(n4539) );
  NAND U5451 ( .A(n4540), .B(n4539), .Z(n4542) );
  XOR U5452 ( .A(n4543), .B(n4542), .Z(c[1912]) );
  NANDN U5453 ( .A(n4541), .B(sreg[1912]), .Z(n4545) );
  NAND U5454 ( .A(n4543), .B(n4542), .Z(n4544) );
  AND U5455 ( .A(n4545), .B(n4544), .Z(n4547) );
  AND U5456 ( .A(b[0]), .B(a[890]), .Z(n4548) );
  XNOR U5457 ( .A(sreg[1913]), .B(n4548), .Z(n4546) );
  XOR U5458 ( .A(n4547), .B(n4546), .Z(c[1913]) );
  AND U5459 ( .A(b[0]), .B(a[891]), .Z(n4551) );
  XNOR U5460 ( .A(sreg[1914]), .B(n4550), .Z(n4549) );
  XNOR U5461 ( .A(n4551), .B(n4549), .Z(c[1914]) );
  NAND U5462 ( .A(b[0]), .B(a[892]), .Z(n4552) );
  XNOR U5463 ( .A(sreg[1915]), .B(n4552), .Z(n4553) );
  XOR U5464 ( .A(n4554), .B(n4553), .Z(c[1915]) );
  NAND U5465 ( .A(b[0]), .B(a[893]), .Z(n4557) );
  XNOR U5466 ( .A(sreg[1916]), .B(n4557), .Z(n4559) );
  NANDN U5467 ( .A(n4552), .B(sreg[1915]), .Z(n4556) );
  NAND U5468 ( .A(n4554), .B(n4553), .Z(n4555) );
  NAND U5469 ( .A(n4556), .B(n4555), .Z(n4558) );
  XOR U5470 ( .A(n4559), .B(n4558), .Z(c[1916]) );
  NAND U5471 ( .A(b[0]), .B(a[894]), .Z(n4562) );
  XNOR U5472 ( .A(sreg[1917]), .B(n4562), .Z(n4564) );
  NANDN U5473 ( .A(n4557), .B(sreg[1916]), .Z(n4561) );
  NAND U5474 ( .A(n4559), .B(n4558), .Z(n4560) );
  NAND U5475 ( .A(n4561), .B(n4560), .Z(n4563) );
  XOR U5476 ( .A(n4564), .B(n4563), .Z(c[1917]) );
  NAND U5477 ( .A(b[0]), .B(a[895]), .Z(n4567) );
  XNOR U5478 ( .A(sreg[1918]), .B(n4567), .Z(n4569) );
  NANDN U5479 ( .A(n4562), .B(sreg[1917]), .Z(n4566) );
  NAND U5480 ( .A(n4564), .B(n4563), .Z(n4565) );
  NAND U5481 ( .A(n4566), .B(n4565), .Z(n4568) );
  XOR U5482 ( .A(n4569), .B(n4568), .Z(c[1918]) );
  NAND U5483 ( .A(b[0]), .B(a[896]), .Z(n4572) );
  XNOR U5484 ( .A(sreg[1919]), .B(n4572), .Z(n4574) );
  NANDN U5485 ( .A(n4567), .B(sreg[1918]), .Z(n4571) );
  NAND U5486 ( .A(n4569), .B(n4568), .Z(n4570) );
  NAND U5487 ( .A(n4571), .B(n4570), .Z(n4573) );
  XOR U5488 ( .A(n4574), .B(n4573), .Z(c[1919]) );
  NAND U5489 ( .A(b[0]), .B(a[897]), .Z(n4577) );
  XNOR U5490 ( .A(sreg[1920]), .B(n4577), .Z(n4579) );
  NANDN U5491 ( .A(n4572), .B(sreg[1919]), .Z(n4576) );
  NAND U5492 ( .A(n4574), .B(n4573), .Z(n4575) );
  NAND U5493 ( .A(n4576), .B(n4575), .Z(n4578) );
  XOR U5494 ( .A(n4579), .B(n4578), .Z(c[1920]) );
  NAND U5495 ( .A(b[0]), .B(a[898]), .Z(n4582) );
  XNOR U5496 ( .A(sreg[1921]), .B(n4582), .Z(n4584) );
  NANDN U5497 ( .A(n4577), .B(sreg[1920]), .Z(n4581) );
  NAND U5498 ( .A(n4579), .B(n4578), .Z(n4580) );
  NAND U5499 ( .A(n4581), .B(n4580), .Z(n4583) );
  XOR U5500 ( .A(n4584), .B(n4583), .Z(c[1921]) );
  NAND U5501 ( .A(b[0]), .B(a[899]), .Z(n4587) );
  XNOR U5502 ( .A(sreg[1922]), .B(n4587), .Z(n4589) );
  NANDN U5503 ( .A(n4582), .B(sreg[1921]), .Z(n4586) );
  NAND U5504 ( .A(n4584), .B(n4583), .Z(n4585) );
  NAND U5505 ( .A(n4586), .B(n4585), .Z(n4588) );
  XOR U5506 ( .A(n4589), .B(n4588), .Z(c[1922]) );
  NAND U5507 ( .A(b[0]), .B(a[900]), .Z(n4592) );
  XNOR U5508 ( .A(sreg[1923]), .B(n4592), .Z(n4594) );
  NANDN U5509 ( .A(n4587), .B(sreg[1922]), .Z(n4591) );
  NAND U5510 ( .A(n4589), .B(n4588), .Z(n4590) );
  NAND U5511 ( .A(n4591), .B(n4590), .Z(n4593) );
  XOR U5512 ( .A(n4594), .B(n4593), .Z(c[1923]) );
  NAND U5513 ( .A(b[0]), .B(a[901]), .Z(n4597) );
  XNOR U5514 ( .A(sreg[1924]), .B(n4597), .Z(n4599) );
  NANDN U5515 ( .A(n4592), .B(sreg[1923]), .Z(n4596) );
  NAND U5516 ( .A(n4594), .B(n4593), .Z(n4595) );
  NAND U5517 ( .A(n4596), .B(n4595), .Z(n4598) );
  XOR U5518 ( .A(n4599), .B(n4598), .Z(c[1924]) );
  NAND U5519 ( .A(b[0]), .B(a[902]), .Z(n4602) );
  XNOR U5520 ( .A(sreg[1925]), .B(n4602), .Z(n4604) );
  NANDN U5521 ( .A(n4597), .B(sreg[1924]), .Z(n4601) );
  NAND U5522 ( .A(n4599), .B(n4598), .Z(n4600) );
  NAND U5523 ( .A(n4601), .B(n4600), .Z(n4603) );
  XOR U5524 ( .A(n4604), .B(n4603), .Z(c[1925]) );
  NAND U5525 ( .A(b[0]), .B(a[903]), .Z(n4607) );
  XNOR U5526 ( .A(sreg[1926]), .B(n4607), .Z(n4609) );
  NANDN U5527 ( .A(n4602), .B(sreg[1925]), .Z(n4606) );
  NAND U5528 ( .A(n4604), .B(n4603), .Z(n4605) );
  NAND U5529 ( .A(n4606), .B(n4605), .Z(n4608) );
  XOR U5530 ( .A(n4609), .B(n4608), .Z(c[1926]) );
  NAND U5531 ( .A(b[0]), .B(a[904]), .Z(n4612) );
  XNOR U5532 ( .A(sreg[1927]), .B(n4612), .Z(n4614) );
  NANDN U5533 ( .A(n4607), .B(sreg[1926]), .Z(n4611) );
  NAND U5534 ( .A(n4609), .B(n4608), .Z(n4610) );
  NAND U5535 ( .A(n4611), .B(n4610), .Z(n4613) );
  XOR U5536 ( .A(n4614), .B(n4613), .Z(c[1927]) );
  NAND U5537 ( .A(b[0]), .B(a[905]), .Z(n4617) );
  XNOR U5538 ( .A(sreg[1928]), .B(n4617), .Z(n4619) );
  NANDN U5539 ( .A(n4612), .B(sreg[1927]), .Z(n4616) );
  NAND U5540 ( .A(n4614), .B(n4613), .Z(n4615) );
  NAND U5541 ( .A(n4616), .B(n4615), .Z(n4618) );
  XOR U5542 ( .A(n4619), .B(n4618), .Z(c[1928]) );
  NANDN U5543 ( .A(n4617), .B(sreg[1928]), .Z(n4621) );
  NAND U5544 ( .A(n4619), .B(n4618), .Z(n4620) );
  AND U5545 ( .A(n4621), .B(n4620), .Z(n4624) );
  NAND U5546 ( .A(b[0]), .B(a[906]), .Z(n4622) );
  XNOR U5547 ( .A(sreg[1929]), .B(n4622), .Z(n4623) );
  XNOR U5548 ( .A(n4624), .B(n4623), .Z(c[1929]) );
  NAND U5549 ( .A(b[0]), .B(a[907]), .Z(n4627) );
  XNOR U5550 ( .A(sreg[1930]), .B(n4627), .Z(n4629) );
  NANDN U5551 ( .A(sreg[1929]), .B(n4622), .Z(n4626) );
  NAND U5552 ( .A(n4624), .B(n4623), .Z(n4625) );
  NAND U5553 ( .A(n4626), .B(n4625), .Z(n4628) );
  XNOR U5554 ( .A(n4629), .B(n4628), .Z(c[1930]) );
  NAND U5555 ( .A(b[0]), .B(a[908]), .Z(n4632) );
  XNOR U5556 ( .A(sreg[1931]), .B(n4632), .Z(n4634) );
  NANDN U5557 ( .A(sreg[1930]), .B(n4627), .Z(n4631) );
  NAND U5558 ( .A(n4629), .B(n4628), .Z(n4630) );
  AND U5559 ( .A(n4631), .B(n4630), .Z(n4633) );
  XOR U5560 ( .A(n4634), .B(n4633), .Z(c[1931]) );
  NAND U5561 ( .A(b[0]), .B(a[909]), .Z(n4637) );
  XNOR U5562 ( .A(sreg[1932]), .B(n4637), .Z(n4639) );
  NANDN U5563 ( .A(n4632), .B(sreg[1931]), .Z(n4636) );
  NAND U5564 ( .A(n4634), .B(n4633), .Z(n4635) );
  AND U5565 ( .A(n4636), .B(n4635), .Z(n4638) );
  XNOR U5566 ( .A(n4639), .B(n4638), .Z(c[1932]) );
  NAND U5567 ( .A(b[0]), .B(a[910]), .Z(n4642) );
  XNOR U5568 ( .A(sreg[1933]), .B(n4642), .Z(n4644) );
  NANDN U5569 ( .A(sreg[1932]), .B(n4637), .Z(n4641) );
  NAND U5570 ( .A(n4639), .B(n4638), .Z(n4640) );
  NAND U5571 ( .A(n4641), .B(n4640), .Z(n4643) );
  XNOR U5572 ( .A(n4644), .B(n4643), .Z(c[1933]) );
  NAND U5573 ( .A(b[0]), .B(a[911]), .Z(n4647) );
  XNOR U5574 ( .A(sreg[1934]), .B(n4647), .Z(n4649) );
  NANDN U5575 ( .A(sreg[1933]), .B(n4642), .Z(n4646) );
  NAND U5576 ( .A(n4644), .B(n4643), .Z(n4645) );
  AND U5577 ( .A(n4646), .B(n4645), .Z(n4648) );
  XOR U5578 ( .A(n4649), .B(n4648), .Z(c[1934]) );
  NANDN U5579 ( .A(n4647), .B(sreg[1934]), .Z(n4651) );
  NAND U5580 ( .A(n4649), .B(n4648), .Z(n4650) );
  AND U5581 ( .A(n4651), .B(n4650), .Z(n4653) );
  AND U5582 ( .A(b[0]), .B(a[912]), .Z(n4654) );
  XNOR U5583 ( .A(sreg[1935]), .B(n4654), .Z(n4652) );
  XOR U5584 ( .A(n4653), .B(n4652), .Z(c[1935]) );
  NAND U5585 ( .A(b[0]), .B(a[913]), .Z(n4655) );
  XNOR U5586 ( .A(sreg[1936]), .B(n4655), .Z(n4657) );
  XOR U5587 ( .A(n4657), .B(n4656), .Z(c[1936]) );
  NAND U5588 ( .A(b[0]), .B(a[914]), .Z(n4660) );
  XNOR U5589 ( .A(sreg[1937]), .B(n4660), .Z(n4662) );
  NANDN U5590 ( .A(n4655), .B(sreg[1936]), .Z(n4659) );
  NAND U5591 ( .A(n4657), .B(n4656), .Z(n4658) );
  NAND U5592 ( .A(n4659), .B(n4658), .Z(n4661) );
  XOR U5593 ( .A(n4662), .B(n4661), .Z(c[1937]) );
  NAND U5594 ( .A(b[0]), .B(a[915]), .Z(n4665) );
  XNOR U5595 ( .A(sreg[1938]), .B(n4665), .Z(n4667) );
  NANDN U5596 ( .A(n4660), .B(sreg[1937]), .Z(n4664) );
  NAND U5597 ( .A(n4662), .B(n4661), .Z(n4663) );
  NAND U5598 ( .A(n4664), .B(n4663), .Z(n4666) );
  XOR U5599 ( .A(n4667), .B(n4666), .Z(c[1938]) );
  NAND U5600 ( .A(b[0]), .B(a[916]), .Z(n4670) );
  XNOR U5601 ( .A(sreg[1939]), .B(n4670), .Z(n4672) );
  NANDN U5602 ( .A(n4665), .B(sreg[1938]), .Z(n4669) );
  NAND U5603 ( .A(n4667), .B(n4666), .Z(n4668) );
  NAND U5604 ( .A(n4669), .B(n4668), .Z(n4671) );
  XOR U5605 ( .A(n4672), .B(n4671), .Z(c[1939]) );
  NANDN U5606 ( .A(n4670), .B(sreg[1939]), .Z(n4674) );
  NAND U5607 ( .A(n4672), .B(n4671), .Z(n4673) );
  AND U5608 ( .A(n4674), .B(n4673), .Z(n4677) );
  NAND U5609 ( .A(b[0]), .B(a[917]), .Z(n4675) );
  XNOR U5610 ( .A(sreg[1940]), .B(n4675), .Z(n4676) );
  XNOR U5611 ( .A(n4677), .B(n4676), .Z(c[1940]) );
  NAND U5612 ( .A(b[0]), .B(a[918]), .Z(n4680) );
  XNOR U5613 ( .A(sreg[1941]), .B(n4680), .Z(n4682) );
  NANDN U5614 ( .A(sreg[1940]), .B(n4675), .Z(n4679) );
  NAND U5615 ( .A(n4677), .B(n4676), .Z(n4678) );
  NAND U5616 ( .A(n4679), .B(n4678), .Z(n4681) );
  XNOR U5617 ( .A(n4682), .B(n4681), .Z(c[1941]) );
  NAND U5618 ( .A(b[0]), .B(a[919]), .Z(n4685) );
  XNOR U5619 ( .A(sreg[1942]), .B(n4685), .Z(n4687) );
  NANDN U5620 ( .A(sreg[1941]), .B(n4680), .Z(n4684) );
  NAND U5621 ( .A(n4682), .B(n4681), .Z(n4683) );
  AND U5622 ( .A(n4684), .B(n4683), .Z(n4686) );
  XOR U5623 ( .A(n4687), .B(n4686), .Z(c[1942]) );
  NAND U5624 ( .A(b[0]), .B(a[920]), .Z(n4690) );
  XNOR U5625 ( .A(sreg[1943]), .B(n4690), .Z(n4692) );
  NANDN U5626 ( .A(n4685), .B(sreg[1942]), .Z(n4689) );
  NAND U5627 ( .A(n4687), .B(n4686), .Z(n4688) );
  AND U5628 ( .A(n4689), .B(n4688), .Z(n4691) );
  XNOR U5629 ( .A(n4692), .B(n4691), .Z(c[1943]) );
  NAND U5630 ( .A(b[0]), .B(a[921]), .Z(n4695) );
  XNOR U5631 ( .A(sreg[1944]), .B(n4695), .Z(n4697) );
  NANDN U5632 ( .A(sreg[1943]), .B(n4690), .Z(n4694) );
  NAND U5633 ( .A(n4692), .B(n4691), .Z(n4693) );
  NAND U5634 ( .A(n4694), .B(n4693), .Z(n4696) );
  XNOR U5635 ( .A(n4697), .B(n4696), .Z(c[1944]) );
  NANDN U5636 ( .A(sreg[1944]), .B(n4695), .Z(n4699) );
  NAND U5637 ( .A(n4697), .B(n4696), .Z(n4698) );
  AND U5638 ( .A(n4699), .B(n4698), .Z(n4702) );
  NAND U5639 ( .A(b[0]), .B(a[922]), .Z(n4700) );
  XNOR U5640 ( .A(sreg[1945]), .B(n4700), .Z(n4701) );
  XOR U5641 ( .A(n4702), .B(n4701), .Z(c[1945]) );
  NAND U5642 ( .A(b[0]), .B(a[923]), .Z(n4705) );
  XNOR U5643 ( .A(sreg[1946]), .B(n4705), .Z(n4707) );
  NANDN U5644 ( .A(n4700), .B(sreg[1945]), .Z(n4704) );
  NAND U5645 ( .A(n4702), .B(n4701), .Z(n4703) );
  NAND U5646 ( .A(n4704), .B(n4703), .Z(n4706) );
  XOR U5647 ( .A(n4707), .B(n4706), .Z(c[1946]) );
  NANDN U5648 ( .A(n4705), .B(sreg[1946]), .Z(n4709) );
  NAND U5649 ( .A(n4707), .B(n4706), .Z(n4708) );
  AND U5650 ( .A(n4709), .B(n4708), .Z(n4712) );
  NAND U5651 ( .A(b[0]), .B(a[924]), .Z(n4710) );
  XNOR U5652 ( .A(sreg[1947]), .B(n4710), .Z(n4711) );
  XNOR U5653 ( .A(n4712), .B(n4711), .Z(c[1947]) );
  NAND U5654 ( .A(b[0]), .B(a[925]), .Z(n4715) );
  XNOR U5655 ( .A(sreg[1948]), .B(n4715), .Z(n4717) );
  NANDN U5656 ( .A(sreg[1947]), .B(n4710), .Z(n4714) );
  NAND U5657 ( .A(n4712), .B(n4711), .Z(n4713) );
  AND U5658 ( .A(n4714), .B(n4713), .Z(n4716) );
  XOR U5659 ( .A(n4717), .B(n4716), .Z(c[1948]) );
  NAND U5660 ( .A(b[0]), .B(a[926]), .Z(n4720) );
  XNOR U5661 ( .A(sreg[1949]), .B(n4720), .Z(n4722) );
  NANDN U5662 ( .A(n4715), .B(sreg[1948]), .Z(n4719) );
  NAND U5663 ( .A(n4717), .B(n4716), .Z(n4718) );
  NAND U5664 ( .A(n4719), .B(n4718), .Z(n4721) );
  XOR U5665 ( .A(n4722), .B(n4721), .Z(c[1949]) );
  NAND U5666 ( .A(b[0]), .B(a[927]), .Z(n4725) );
  XNOR U5667 ( .A(sreg[1950]), .B(n4725), .Z(n4727) );
  NANDN U5668 ( .A(n4720), .B(sreg[1949]), .Z(n4724) );
  NAND U5669 ( .A(n4722), .B(n4721), .Z(n4723) );
  AND U5670 ( .A(n4724), .B(n4723), .Z(n4726) );
  XNOR U5671 ( .A(n4727), .B(n4726), .Z(c[1950]) );
  NAND U5672 ( .A(b[0]), .B(a[928]), .Z(n4730) );
  XNOR U5673 ( .A(sreg[1951]), .B(n4730), .Z(n4732) );
  NANDN U5674 ( .A(sreg[1950]), .B(n4725), .Z(n4729) );
  NAND U5675 ( .A(n4727), .B(n4726), .Z(n4728) );
  AND U5676 ( .A(n4729), .B(n4728), .Z(n4731) );
  XOR U5677 ( .A(n4732), .B(n4731), .Z(c[1951]) );
  NAND U5678 ( .A(b[0]), .B(a[929]), .Z(n4735) );
  XNOR U5679 ( .A(sreg[1952]), .B(n4735), .Z(n4737) );
  NANDN U5680 ( .A(n4730), .B(sreg[1951]), .Z(n4734) );
  NAND U5681 ( .A(n4732), .B(n4731), .Z(n4733) );
  NAND U5682 ( .A(n4734), .B(n4733), .Z(n4736) );
  XOR U5683 ( .A(n4737), .B(n4736), .Z(c[1952]) );
  NANDN U5684 ( .A(n4735), .B(sreg[1952]), .Z(n4739) );
  NAND U5685 ( .A(n4737), .B(n4736), .Z(n4738) );
  AND U5686 ( .A(n4739), .B(n4738), .Z(n4742) );
  NAND U5687 ( .A(b[0]), .B(a[930]), .Z(n4740) );
  XNOR U5688 ( .A(sreg[1953]), .B(n4740), .Z(n4741) );
  XNOR U5689 ( .A(n4742), .B(n4741), .Z(c[1953]) );
  NANDN U5690 ( .A(sreg[1953]), .B(n4740), .Z(n4744) );
  NAND U5691 ( .A(n4742), .B(n4741), .Z(n4743) );
  AND U5692 ( .A(n4744), .B(n4743), .Z(n4747) );
  NAND U5693 ( .A(b[0]), .B(a[931]), .Z(n4745) );
  XNOR U5694 ( .A(sreg[1954]), .B(n4745), .Z(n4746) );
  XOR U5695 ( .A(n4747), .B(n4746), .Z(c[1954]) );
  NAND U5696 ( .A(b[0]), .B(a[932]), .Z(n4750) );
  XNOR U5697 ( .A(sreg[1955]), .B(n4750), .Z(n4752) );
  NANDN U5698 ( .A(n4745), .B(sreg[1954]), .Z(n4749) );
  NAND U5699 ( .A(n4747), .B(n4746), .Z(n4748) );
  NAND U5700 ( .A(n4749), .B(n4748), .Z(n4751) );
  XOR U5701 ( .A(n4752), .B(n4751), .Z(c[1955]) );
  NAND U5702 ( .A(b[0]), .B(a[933]), .Z(n4755) );
  XNOR U5703 ( .A(sreg[1956]), .B(n4755), .Z(n4757) );
  NANDN U5704 ( .A(n4750), .B(sreg[1955]), .Z(n4754) );
  NAND U5705 ( .A(n4752), .B(n4751), .Z(n4753) );
  NAND U5706 ( .A(n4754), .B(n4753), .Z(n4756) );
  XOR U5707 ( .A(n4757), .B(n4756), .Z(c[1956]) );
  NAND U5708 ( .A(b[0]), .B(a[934]), .Z(n4760) );
  XNOR U5709 ( .A(sreg[1957]), .B(n4760), .Z(n4762) );
  NANDN U5710 ( .A(n4755), .B(sreg[1956]), .Z(n4759) );
  NAND U5711 ( .A(n4757), .B(n4756), .Z(n4758) );
  NAND U5712 ( .A(n4759), .B(n4758), .Z(n4761) );
  XOR U5713 ( .A(n4762), .B(n4761), .Z(c[1957]) );
  NAND U5714 ( .A(b[0]), .B(a[935]), .Z(n4765) );
  XNOR U5715 ( .A(sreg[1958]), .B(n4765), .Z(n4767) );
  NANDN U5716 ( .A(n4760), .B(sreg[1957]), .Z(n4764) );
  NAND U5717 ( .A(n4762), .B(n4761), .Z(n4763) );
  NAND U5718 ( .A(n4764), .B(n4763), .Z(n4766) );
  XOR U5719 ( .A(n4767), .B(n4766), .Z(c[1958]) );
  NAND U5720 ( .A(b[0]), .B(a[936]), .Z(n4772) );
  NANDN U5721 ( .A(n4765), .B(sreg[1958]), .Z(n4769) );
  NAND U5722 ( .A(n4767), .B(n4766), .Z(n4768) );
  NAND U5723 ( .A(n4769), .B(n4768), .Z(n4771) );
  XOR U5724 ( .A(sreg[1959]), .B(n4771), .Z(n4770) );
  XNOR U5725 ( .A(n4772), .B(n4770), .Z(c[1959]) );
  NAND U5726 ( .A(b[0]), .B(a[937]), .Z(n4773) );
  XNOR U5727 ( .A(sreg[1960]), .B(n4773), .Z(n4774) );
  XOR U5728 ( .A(n4775), .B(n4774), .Z(c[1960]) );
  NANDN U5729 ( .A(n4773), .B(sreg[1960]), .Z(n4777) );
  NAND U5730 ( .A(n4775), .B(n4774), .Z(n4776) );
  AND U5731 ( .A(n4777), .B(n4776), .Z(n4779) );
  AND U5732 ( .A(b[0]), .B(a[938]), .Z(n4780) );
  XNOR U5733 ( .A(sreg[1961]), .B(n4780), .Z(n4778) );
  XOR U5734 ( .A(n4779), .B(n4778), .Z(c[1961]) );
  NAND U5735 ( .A(b[0]), .B(a[939]), .Z(n4781) );
  XNOR U5736 ( .A(sreg[1962]), .B(n4781), .Z(n4782) );
  XOR U5737 ( .A(n4783), .B(n4782), .Z(c[1962]) );
  NAND U5738 ( .A(b[0]), .B(a[940]), .Z(n4786) );
  XNOR U5739 ( .A(sreg[1963]), .B(n4786), .Z(n4788) );
  NANDN U5740 ( .A(n4781), .B(sreg[1962]), .Z(n4785) );
  NAND U5741 ( .A(n4783), .B(n4782), .Z(n4784) );
  NAND U5742 ( .A(n4785), .B(n4784), .Z(n4787) );
  XOR U5743 ( .A(n4788), .B(n4787), .Z(c[1963]) );
  NAND U5744 ( .A(b[0]), .B(a[941]), .Z(n4791) );
  XNOR U5745 ( .A(sreg[1964]), .B(n4791), .Z(n4793) );
  NANDN U5746 ( .A(n4786), .B(sreg[1963]), .Z(n4790) );
  NAND U5747 ( .A(n4788), .B(n4787), .Z(n4789) );
  AND U5748 ( .A(n4790), .B(n4789), .Z(n4792) );
  XNOR U5749 ( .A(n4793), .B(n4792), .Z(c[1964]) );
  NANDN U5750 ( .A(sreg[1964]), .B(n4791), .Z(n4795) );
  NAND U5751 ( .A(n4793), .B(n4792), .Z(n4794) );
  AND U5752 ( .A(n4795), .B(n4794), .Z(n4798) );
  NAND U5753 ( .A(b[0]), .B(a[942]), .Z(n4796) );
  XNOR U5754 ( .A(sreg[1965]), .B(n4796), .Z(n4797) );
  XOR U5755 ( .A(n4798), .B(n4797), .Z(c[1965]) );
  NAND U5756 ( .A(b[0]), .B(a[943]), .Z(n4801) );
  XNOR U5757 ( .A(sreg[1966]), .B(n4801), .Z(n4803) );
  NANDN U5758 ( .A(n4796), .B(sreg[1965]), .Z(n4800) );
  NAND U5759 ( .A(n4798), .B(n4797), .Z(n4799) );
  NAND U5760 ( .A(n4800), .B(n4799), .Z(n4802) );
  XOR U5761 ( .A(n4803), .B(n4802), .Z(c[1966]) );
  AND U5762 ( .A(b[0]), .B(a[944]), .Z(n4807) );
  NANDN U5763 ( .A(n4801), .B(sreg[1966]), .Z(n4805) );
  NAND U5764 ( .A(n4803), .B(n4802), .Z(n4804) );
  AND U5765 ( .A(n4805), .B(n4804), .Z(n4808) );
  XNOR U5766 ( .A(sreg[1967]), .B(n4808), .Z(n4806) );
  XOR U5767 ( .A(n4807), .B(n4806), .Z(c[1967]) );
  NAND U5768 ( .A(b[0]), .B(a[945]), .Z(n4809) );
  XNOR U5769 ( .A(sreg[1968]), .B(n4809), .Z(n4810) );
  XNOR U5770 ( .A(n4811), .B(n4810), .Z(c[1968]) );
  NAND U5771 ( .A(b[0]), .B(a[946]), .Z(n4814) );
  XNOR U5772 ( .A(sreg[1969]), .B(n4814), .Z(n4816) );
  NANDN U5773 ( .A(n4809), .B(sreg[1968]), .Z(n4813) );
  NANDN U5774 ( .A(n4811), .B(n4810), .Z(n4812) );
  NAND U5775 ( .A(n4813), .B(n4812), .Z(n4815) );
  XOR U5776 ( .A(n4816), .B(n4815), .Z(c[1969]) );
  NANDN U5777 ( .A(n4814), .B(sreg[1969]), .Z(n4818) );
  NAND U5778 ( .A(n4816), .B(n4815), .Z(n4817) );
  NAND U5779 ( .A(n4818), .B(n4817), .Z(n4821) );
  NAND U5780 ( .A(b[0]), .B(a[947]), .Z(n4820) );
  XOR U5781 ( .A(sreg[1970]), .B(n4820), .Z(n4819) );
  XNOR U5782 ( .A(n4821), .B(n4819), .Z(c[1970]) );
  NAND U5783 ( .A(b[0]), .B(a[948]), .Z(n4822) );
  XNOR U5784 ( .A(sreg[1971]), .B(n4822), .Z(n4823) );
  XOR U5785 ( .A(n4824), .B(n4823), .Z(c[1971]) );
  NANDN U5786 ( .A(n4822), .B(sreg[1971]), .Z(n4826) );
  NAND U5787 ( .A(n4824), .B(n4823), .Z(n4825) );
  AND U5788 ( .A(n4826), .B(n4825), .Z(n4829) );
  NAND U5789 ( .A(b[0]), .B(a[949]), .Z(n4827) );
  XNOR U5790 ( .A(sreg[1972]), .B(n4827), .Z(n4828) );
  XNOR U5791 ( .A(n4829), .B(n4828), .Z(c[1972]) );
  NAND U5792 ( .A(b[0]), .B(a[950]), .Z(n4832) );
  XNOR U5793 ( .A(sreg[1973]), .B(n4832), .Z(n4834) );
  NANDN U5794 ( .A(sreg[1972]), .B(n4827), .Z(n4831) );
  NAND U5795 ( .A(n4829), .B(n4828), .Z(n4830) );
  AND U5796 ( .A(n4831), .B(n4830), .Z(n4833) );
  XOR U5797 ( .A(n4834), .B(n4833), .Z(c[1973]) );
  NAND U5798 ( .A(b[0]), .B(a[951]), .Z(n4837) );
  XNOR U5799 ( .A(sreg[1974]), .B(n4837), .Z(n4839) );
  NANDN U5800 ( .A(n4832), .B(sreg[1973]), .Z(n4836) );
  NAND U5801 ( .A(n4834), .B(n4833), .Z(n4835) );
  NAND U5802 ( .A(n4836), .B(n4835), .Z(n4838) );
  XOR U5803 ( .A(n4839), .B(n4838), .Z(c[1974]) );
  NANDN U5804 ( .A(n4837), .B(sreg[1974]), .Z(n4841) );
  NAND U5805 ( .A(n4839), .B(n4838), .Z(n4840) );
  AND U5806 ( .A(n4841), .B(n4840), .Z(n4844) );
  NAND U5807 ( .A(b[0]), .B(a[952]), .Z(n4842) );
  XNOR U5808 ( .A(sreg[1975]), .B(n4842), .Z(n4843) );
  XNOR U5809 ( .A(n4844), .B(n4843), .Z(c[1975]) );
  NANDN U5810 ( .A(sreg[1975]), .B(n4842), .Z(n4846) );
  NAND U5811 ( .A(n4844), .B(n4843), .Z(n4845) );
  AND U5812 ( .A(n4846), .B(n4845), .Z(n4849) );
  NAND U5813 ( .A(b[0]), .B(a[953]), .Z(n4847) );
  XNOR U5814 ( .A(sreg[1976]), .B(n4847), .Z(n4848) );
  XOR U5815 ( .A(n4849), .B(n4848), .Z(c[1976]) );
  NAND U5816 ( .A(b[0]), .B(a[954]), .Z(n4852) );
  XNOR U5817 ( .A(sreg[1977]), .B(n4852), .Z(n4854) );
  NANDN U5818 ( .A(n4847), .B(sreg[1976]), .Z(n4851) );
  NAND U5819 ( .A(n4849), .B(n4848), .Z(n4850) );
  NAND U5820 ( .A(n4851), .B(n4850), .Z(n4853) );
  XOR U5821 ( .A(n4854), .B(n4853), .Z(c[1977]) );
  NAND U5822 ( .A(b[0]), .B(a[955]), .Z(n4857) );
  XNOR U5823 ( .A(sreg[1978]), .B(n4857), .Z(n4859) );
  NANDN U5824 ( .A(n4852), .B(sreg[1977]), .Z(n4856) );
  NAND U5825 ( .A(n4854), .B(n4853), .Z(n4855) );
  AND U5826 ( .A(n4856), .B(n4855), .Z(n4858) );
  XNOR U5827 ( .A(n4859), .B(n4858), .Z(c[1978]) );
  NAND U5828 ( .A(b[0]), .B(a[956]), .Z(n4862) );
  XNOR U5829 ( .A(sreg[1979]), .B(n4862), .Z(n4864) );
  NANDN U5830 ( .A(sreg[1978]), .B(n4857), .Z(n4861) );
  NAND U5831 ( .A(n4859), .B(n4858), .Z(n4860) );
  AND U5832 ( .A(n4861), .B(n4860), .Z(n4863) );
  XOR U5833 ( .A(n4864), .B(n4863), .Z(c[1979]) );
  NAND U5834 ( .A(b[0]), .B(a[957]), .Z(n4867) );
  XNOR U5835 ( .A(sreg[1980]), .B(n4867), .Z(n4869) );
  NANDN U5836 ( .A(n4862), .B(sreg[1979]), .Z(n4866) );
  NAND U5837 ( .A(n4864), .B(n4863), .Z(n4865) );
  NAND U5838 ( .A(n4866), .B(n4865), .Z(n4868) );
  XOR U5839 ( .A(n4869), .B(n4868), .Z(c[1980]) );
  NANDN U5840 ( .A(n4867), .B(sreg[1980]), .Z(n4871) );
  NAND U5841 ( .A(n4869), .B(n4868), .Z(n4870) );
  AND U5842 ( .A(n4871), .B(n4870), .Z(n4874) );
  NAND U5843 ( .A(b[0]), .B(a[958]), .Z(n4872) );
  XNOR U5844 ( .A(sreg[1981]), .B(n4872), .Z(n4873) );
  XNOR U5845 ( .A(n4874), .B(n4873), .Z(c[1981]) );
  NAND U5846 ( .A(b[0]), .B(a[959]), .Z(n4877) );
  XNOR U5847 ( .A(sreg[1982]), .B(n4877), .Z(n4879) );
  NANDN U5848 ( .A(sreg[1981]), .B(n4872), .Z(n4876) );
  NAND U5849 ( .A(n4874), .B(n4873), .Z(n4875) );
  NAND U5850 ( .A(n4876), .B(n4875), .Z(n4878) );
  XNOR U5851 ( .A(n4879), .B(n4878), .Z(c[1982]) );
  NAND U5852 ( .A(b[0]), .B(a[960]), .Z(n4882) );
  XNOR U5853 ( .A(sreg[1983]), .B(n4882), .Z(n4884) );
  NANDN U5854 ( .A(sreg[1982]), .B(n4877), .Z(n4881) );
  NAND U5855 ( .A(n4879), .B(n4878), .Z(n4880) );
  AND U5856 ( .A(n4881), .B(n4880), .Z(n4883) );
  XOR U5857 ( .A(n4884), .B(n4883), .Z(c[1983]) );
  NANDN U5858 ( .A(n4882), .B(sreg[1983]), .Z(n4886) );
  NAND U5859 ( .A(n4884), .B(n4883), .Z(n4885) );
  AND U5860 ( .A(n4886), .B(n4885), .Z(n4889) );
  NAND U5861 ( .A(b[0]), .B(a[961]), .Z(n4887) );
  XNOR U5862 ( .A(sreg[1984]), .B(n4887), .Z(n4888) );
  XNOR U5863 ( .A(n4889), .B(n4888), .Z(c[1984]) );
  NAND U5864 ( .A(b[0]), .B(a[962]), .Z(n4892) );
  XNOR U5865 ( .A(sreg[1985]), .B(n4892), .Z(n4894) );
  NANDN U5866 ( .A(sreg[1984]), .B(n4887), .Z(n4891) );
  NAND U5867 ( .A(n4889), .B(n4888), .Z(n4890) );
  NAND U5868 ( .A(n4891), .B(n4890), .Z(n4893) );
  XNOR U5869 ( .A(n4894), .B(n4893), .Z(c[1985]) );
  NANDN U5870 ( .A(sreg[1985]), .B(n4892), .Z(n4896) );
  NAND U5871 ( .A(n4894), .B(n4893), .Z(n4895) );
  AND U5872 ( .A(n4896), .B(n4895), .Z(n4899) );
  NAND U5873 ( .A(b[0]), .B(a[963]), .Z(n4897) );
  XNOR U5874 ( .A(sreg[1986]), .B(n4897), .Z(n4898) );
  XOR U5875 ( .A(n4899), .B(n4898), .Z(c[1986]) );
  NAND U5876 ( .A(b[0]), .B(a[964]), .Z(n4902) );
  XNOR U5877 ( .A(sreg[1987]), .B(n4902), .Z(n4904) );
  NANDN U5878 ( .A(n4897), .B(sreg[1986]), .Z(n4901) );
  NAND U5879 ( .A(n4899), .B(n4898), .Z(n4900) );
  NAND U5880 ( .A(n4901), .B(n4900), .Z(n4903) );
  XOR U5881 ( .A(n4904), .B(n4903), .Z(c[1987]) );
  NAND U5882 ( .A(b[0]), .B(a[965]), .Z(n4907) );
  XNOR U5883 ( .A(sreg[1988]), .B(n4907), .Z(n4909) );
  NANDN U5884 ( .A(n4902), .B(sreg[1987]), .Z(n4906) );
  NAND U5885 ( .A(n4904), .B(n4903), .Z(n4905) );
  AND U5886 ( .A(n4906), .B(n4905), .Z(n4908) );
  XNOR U5887 ( .A(n4909), .B(n4908), .Z(c[1988]) );
  NANDN U5888 ( .A(sreg[1988]), .B(n4907), .Z(n4911) );
  NAND U5889 ( .A(n4909), .B(n4908), .Z(n4910) );
  AND U5890 ( .A(n4911), .B(n4910), .Z(n4914) );
  NAND U5891 ( .A(b[0]), .B(a[966]), .Z(n4912) );
  XNOR U5892 ( .A(sreg[1989]), .B(n4912), .Z(n4913) );
  XOR U5893 ( .A(n4914), .B(n4913), .Z(c[1989]) );
  NAND U5894 ( .A(b[0]), .B(a[967]), .Z(n4917) );
  XNOR U5895 ( .A(sreg[1990]), .B(n4917), .Z(n4919) );
  NANDN U5896 ( .A(n4912), .B(sreg[1989]), .Z(n4916) );
  NAND U5897 ( .A(n4914), .B(n4913), .Z(n4915) );
  NAND U5898 ( .A(n4916), .B(n4915), .Z(n4918) );
  XOR U5899 ( .A(n4919), .B(n4918), .Z(c[1990]) );
  NAND U5900 ( .A(b[0]), .B(a[968]), .Z(n4922) );
  XNOR U5901 ( .A(sreg[1991]), .B(n4922), .Z(n4924) );
  NANDN U5902 ( .A(n4917), .B(sreg[1990]), .Z(n4921) );
  NAND U5903 ( .A(n4919), .B(n4918), .Z(n4920) );
  NAND U5904 ( .A(n4921), .B(n4920), .Z(n4923) );
  XOR U5905 ( .A(n4924), .B(n4923), .Z(c[1991]) );
  NAND U5906 ( .A(b[0]), .B(a[969]), .Z(n4927) );
  XNOR U5907 ( .A(sreg[1992]), .B(n4927), .Z(n4929) );
  NANDN U5908 ( .A(n4922), .B(sreg[1991]), .Z(n4926) );
  NAND U5909 ( .A(n4924), .B(n4923), .Z(n4925) );
  NAND U5910 ( .A(n4926), .B(n4925), .Z(n4928) );
  XOR U5911 ( .A(n4929), .B(n4928), .Z(c[1992]) );
  NAND U5912 ( .A(b[0]), .B(a[970]), .Z(n4932) );
  XNOR U5913 ( .A(sreg[1993]), .B(n4932), .Z(n4934) );
  NANDN U5914 ( .A(n4927), .B(sreg[1992]), .Z(n4931) );
  NAND U5915 ( .A(n4929), .B(n4928), .Z(n4930) );
  AND U5916 ( .A(n4931), .B(n4930), .Z(n4933) );
  XNOR U5917 ( .A(n4934), .B(n4933), .Z(c[1993]) );
  NAND U5918 ( .A(b[0]), .B(a[971]), .Z(n4937) );
  XNOR U5919 ( .A(sreg[1994]), .B(n4937), .Z(n4939) );
  NANDN U5920 ( .A(sreg[1993]), .B(n4932), .Z(n4936) );
  NAND U5921 ( .A(n4934), .B(n4933), .Z(n4935) );
  AND U5922 ( .A(n4936), .B(n4935), .Z(n4938) );
  XOR U5923 ( .A(n4939), .B(n4938), .Z(c[1994]) );
  NAND U5924 ( .A(b[0]), .B(a[972]), .Z(n4942) );
  XNOR U5925 ( .A(sreg[1995]), .B(n4942), .Z(n4944) );
  NANDN U5926 ( .A(n4937), .B(sreg[1994]), .Z(n4941) );
  NAND U5927 ( .A(n4939), .B(n4938), .Z(n4940) );
  NAND U5928 ( .A(n4941), .B(n4940), .Z(n4943) );
  XOR U5929 ( .A(n4944), .B(n4943), .Z(c[1995]) );
  NANDN U5930 ( .A(n4942), .B(sreg[1995]), .Z(n4946) );
  NAND U5931 ( .A(n4944), .B(n4943), .Z(n4945) );
  AND U5932 ( .A(n4946), .B(n4945), .Z(n4949) );
  NAND U5933 ( .A(b[0]), .B(a[973]), .Z(n4947) );
  XNOR U5934 ( .A(sreg[1996]), .B(n4947), .Z(n4948) );
  XNOR U5935 ( .A(n4949), .B(n4948), .Z(c[1996]) );
  NANDN U5936 ( .A(sreg[1996]), .B(n4947), .Z(n4951) );
  NAND U5937 ( .A(n4949), .B(n4948), .Z(n4950) );
  AND U5938 ( .A(n4951), .B(n4950), .Z(n4954) );
  NAND U5939 ( .A(b[0]), .B(a[974]), .Z(n4952) );
  XNOR U5940 ( .A(sreg[1997]), .B(n4952), .Z(n4953) );
  XOR U5941 ( .A(n4954), .B(n4953), .Z(c[1997]) );
  NAND U5942 ( .A(b[0]), .B(a[975]), .Z(n4957) );
  XNOR U5943 ( .A(sreg[1998]), .B(n4957), .Z(n4959) );
  NANDN U5944 ( .A(n4952), .B(sreg[1997]), .Z(n4956) );
  NAND U5945 ( .A(n4954), .B(n4953), .Z(n4955) );
  NAND U5946 ( .A(n4956), .B(n4955), .Z(n4958) );
  XOR U5947 ( .A(n4959), .B(n4958), .Z(c[1998]) );
  NANDN U5948 ( .A(n4957), .B(sreg[1998]), .Z(n4961) );
  NAND U5949 ( .A(n4959), .B(n4958), .Z(n4960) );
  AND U5950 ( .A(n4961), .B(n4960), .Z(n4963) );
  AND U5951 ( .A(b[0]), .B(a[976]), .Z(n4964) );
  XNOR U5952 ( .A(sreg[1999]), .B(n4964), .Z(n4962) );
  XOR U5953 ( .A(n4963), .B(n4962), .Z(c[1999]) );
  NAND U5954 ( .A(b[0]), .B(a[977]), .Z(n4965) );
  XNOR U5955 ( .A(sreg[2000]), .B(n4965), .Z(n4967) );
  XOR U5956 ( .A(n4967), .B(n4966), .Z(c[2000]) );
  NAND U5957 ( .A(b[0]), .B(a[978]), .Z(n4970) );
  XNOR U5958 ( .A(sreg[2001]), .B(n4970), .Z(n4972) );
  NANDN U5959 ( .A(n4965), .B(sreg[2000]), .Z(n4969) );
  NAND U5960 ( .A(n4967), .B(n4966), .Z(n4968) );
  NAND U5961 ( .A(n4969), .B(n4968), .Z(n4971) );
  XOR U5962 ( .A(n4972), .B(n4971), .Z(c[2001]) );
  NANDN U5963 ( .A(n4970), .B(sreg[2001]), .Z(n4974) );
  NAND U5964 ( .A(n4972), .B(n4971), .Z(n4973) );
  NAND U5965 ( .A(n4974), .B(n4973), .Z(n4977) );
  NAND U5966 ( .A(b[0]), .B(a[979]), .Z(n4976) );
  XOR U5967 ( .A(sreg[2002]), .B(n4976), .Z(n4975) );
  XNOR U5968 ( .A(n4977), .B(n4975), .Z(c[2002]) );
  NAND U5969 ( .A(b[0]), .B(a[980]), .Z(n4978) );
  XNOR U5970 ( .A(sreg[2003]), .B(n4978), .Z(n4979) );
  XOR U5971 ( .A(n4980), .B(n4979), .Z(c[2003]) );
  NAND U5972 ( .A(b[0]), .B(a[981]), .Z(n4983) );
  XNOR U5973 ( .A(sreg[2004]), .B(n4983), .Z(n4985) );
  NANDN U5974 ( .A(sreg[2003]), .B(n4978), .Z(n4982) );
  NANDN U5975 ( .A(n4980), .B(n4979), .Z(n4981) );
  AND U5976 ( .A(n4982), .B(n4981), .Z(n4984) );
  XOR U5977 ( .A(n4985), .B(n4984), .Z(c[2004]) );
  AND U5978 ( .A(b[0]), .B(a[982]), .Z(n4989) );
  NANDN U5979 ( .A(n4983), .B(sreg[2004]), .Z(n4987) );
  NAND U5980 ( .A(n4985), .B(n4984), .Z(n4986) );
  AND U5981 ( .A(n4987), .B(n4986), .Z(n4990) );
  XNOR U5982 ( .A(sreg[2005]), .B(n4990), .Z(n4988) );
  XOR U5983 ( .A(n4989), .B(n4988), .Z(c[2005]) );
  NAND U5984 ( .A(b[0]), .B(a[983]), .Z(n4991) );
  XNOR U5985 ( .A(sreg[2006]), .B(n4991), .Z(n4992) );
  XNOR U5986 ( .A(n4993), .B(n4992), .Z(c[2006]) );
  NANDN U5987 ( .A(sreg[2006]), .B(n4991), .Z(n4995) );
  NAND U5988 ( .A(n4993), .B(n4992), .Z(n4994) );
  AND U5989 ( .A(n4995), .B(n4994), .Z(n4998) );
  NAND U5990 ( .A(b[0]), .B(a[984]), .Z(n4996) );
  XNOR U5991 ( .A(sreg[2007]), .B(n4996), .Z(n4997) );
  XOR U5992 ( .A(n4998), .B(n4997), .Z(c[2007]) );
  NAND U5993 ( .A(b[0]), .B(a[985]), .Z(n5001) );
  XNOR U5994 ( .A(sreg[2008]), .B(n5001), .Z(n5003) );
  NANDN U5995 ( .A(n4996), .B(sreg[2007]), .Z(n5000) );
  NAND U5996 ( .A(n4998), .B(n4997), .Z(n4999) );
  NAND U5997 ( .A(n5000), .B(n4999), .Z(n5002) );
  XOR U5998 ( .A(n5003), .B(n5002), .Z(c[2008]) );
  NAND U5999 ( .A(b[0]), .B(a[986]), .Z(n5006) );
  XNOR U6000 ( .A(sreg[2009]), .B(n5006), .Z(n5008) );
  NANDN U6001 ( .A(n5001), .B(sreg[2008]), .Z(n5005) );
  NAND U6002 ( .A(n5003), .B(n5002), .Z(n5004) );
  NAND U6003 ( .A(n5005), .B(n5004), .Z(n5007) );
  XOR U6004 ( .A(n5008), .B(n5007), .Z(c[2009]) );
  NAND U6005 ( .A(b[0]), .B(a[987]), .Z(n5013) );
  NANDN U6006 ( .A(n5006), .B(sreg[2009]), .Z(n5010) );
  NAND U6007 ( .A(n5008), .B(n5007), .Z(n5009) );
  NAND U6008 ( .A(n5010), .B(n5009), .Z(n5012) );
  XOR U6009 ( .A(n5012), .B(sreg[2010]), .Z(n5011) );
  XNOR U6010 ( .A(n5013), .B(n5011), .Z(c[2010]) );
  NAND U6011 ( .A(b[0]), .B(a[988]), .Z(n5014) );
  XNOR U6012 ( .A(sreg[2011]), .B(n5014), .Z(n5015) );
  XNOR U6013 ( .A(n5016), .B(n5015), .Z(c[2011]) );
  NAND U6014 ( .A(b[0]), .B(a[989]), .Z(n5019) );
  XNOR U6015 ( .A(sreg[2012]), .B(n5019), .Z(n5021) );
  NANDN U6016 ( .A(n5014), .B(sreg[2011]), .Z(n5018) );
  NANDN U6017 ( .A(n5016), .B(n5015), .Z(n5017) );
  NAND U6018 ( .A(n5018), .B(n5017), .Z(n5020) );
  XOR U6019 ( .A(n5021), .B(n5020), .Z(c[2012]) );
  NANDN U6020 ( .A(n5019), .B(sreg[2012]), .Z(n5023) );
  NAND U6021 ( .A(n5021), .B(n5020), .Z(n5022) );
  NAND U6022 ( .A(n5023), .B(n5022), .Z(n5026) );
  NAND U6023 ( .A(b[0]), .B(a[990]), .Z(n5025) );
  XOR U6024 ( .A(sreg[2013]), .B(n5025), .Z(n5024) );
  XNOR U6025 ( .A(n5026), .B(n5024), .Z(c[2013]) );
  NAND U6026 ( .A(b[0]), .B(a[991]), .Z(n5028) );
  XOR U6027 ( .A(sreg[2014]), .B(n5028), .Z(n5027) );
  XNOR U6028 ( .A(n5029), .B(n5027), .Z(c[2014]) );
  NAND U6029 ( .A(b[0]), .B(a[992]), .Z(n5030) );
  XNOR U6030 ( .A(sreg[2015]), .B(n5030), .Z(n5031) );
  XOR U6031 ( .A(n5032), .B(n5031), .Z(c[2015]) );
  AND U6032 ( .A(b[0]), .B(a[993]), .Z(n5036) );
  NANDN U6033 ( .A(n5030), .B(sreg[2015]), .Z(n5034) );
  NAND U6034 ( .A(n5032), .B(n5031), .Z(n5033) );
  AND U6035 ( .A(n5034), .B(n5033), .Z(n5037) );
  XNOR U6036 ( .A(sreg[2016]), .B(n5037), .Z(n5035) );
  XOR U6037 ( .A(n5036), .B(n5035), .Z(c[2016]) );
  AND U6038 ( .A(b[0]), .B(a[994]), .Z(n5039) );
  XNOR U6039 ( .A(sreg[2017]), .B(n5040), .Z(n5038) );
  XOR U6040 ( .A(n5039), .B(n5038), .Z(c[2017]) );
  NAND U6041 ( .A(b[0]), .B(a[995]), .Z(n5041) );
  XNOR U6042 ( .A(sreg[2018]), .B(n5041), .Z(n5042) );
  XNOR U6043 ( .A(n5043), .B(n5042), .Z(c[2018]) );
  NAND U6044 ( .A(b[0]), .B(a[996]), .Z(n5046) );
  XNOR U6045 ( .A(sreg[2019]), .B(n5046), .Z(n5048) );
  NANDN U6046 ( .A(n5041), .B(sreg[2018]), .Z(n5045) );
  NANDN U6047 ( .A(n5043), .B(n5042), .Z(n5044) );
  NAND U6048 ( .A(n5045), .B(n5044), .Z(n5047) );
  XOR U6049 ( .A(n5048), .B(n5047), .Z(c[2019]) );
  NAND U6050 ( .A(b[0]), .B(a[997]), .Z(n5051) );
  XNOR U6051 ( .A(sreg[2020]), .B(n5051), .Z(n5053) );
  NANDN U6052 ( .A(n5046), .B(sreg[2019]), .Z(n5050) );
  NAND U6053 ( .A(n5048), .B(n5047), .Z(n5049) );
  NAND U6054 ( .A(n5050), .B(n5049), .Z(n5052) );
  XOR U6055 ( .A(n5053), .B(n5052), .Z(c[2020]) );
  NAND U6056 ( .A(b[0]), .B(a[998]), .Z(n5056) );
  XNOR U6057 ( .A(sreg[2021]), .B(n5056), .Z(n5058) );
  NANDN U6058 ( .A(n5051), .B(sreg[2020]), .Z(n5055) );
  NAND U6059 ( .A(n5053), .B(n5052), .Z(n5054) );
  AND U6060 ( .A(n5055), .B(n5054), .Z(n5057) );
  XNOR U6061 ( .A(n5058), .B(n5057), .Z(c[2021]) );
  NANDN U6062 ( .A(sreg[2021]), .B(n5056), .Z(n5060) );
  NAND U6063 ( .A(n5058), .B(n5057), .Z(n5059) );
  AND U6064 ( .A(n5060), .B(n5059), .Z(n5063) );
  NAND U6065 ( .A(b[0]), .B(a[999]), .Z(n5061) );
  XNOR U6066 ( .A(sreg[2022]), .B(n5061), .Z(n5062) );
  XOR U6067 ( .A(n5063), .B(n5062), .Z(c[2022]) );
  NAND U6068 ( .A(b[0]), .B(a[1000]), .Z(n5066) );
  XNOR U6069 ( .A(sreg[2023]), .B(n5066), .Z(n5068) );
  NANDN U6070 ( .A(n5061), .B(sreg[2022]), .Z(n5065) );
  NAND U6071 ( .A(n5063), .B(n5062), .Z(n5064) );
  NAND U6072 ( .A(n5065), .B(n5064), .Z(n5067) );
  XOR U6073 ( .A(n5068), .B(n5067), .Z(c[2023]) );
  NAND U6074 ( .A(b[0]), .B(a[1001]), .Z(n5071) );
  XNOR U6075 ( .A(sreg[2024]), .B(n5071), .Z(n5073) );
  NANDN U6076 ( .A(n5066), .B(sreg[2023]), .Z(n5070) );
  NAND U6077 ( .A(n5068), .B(n5067), .Z(n5069) );
  NAND U6078 ( .A(n5070), .B(n5069), .Z(n5072) );
  XOR U6079 ( .A(n5073), .B(n5072), .Z(c[2024]) );
  NAND U6080 ( .A(b[0]), .B(a[1002]), .Z(n5076) );
  XNOR U6081 ( .A(sreg[2025]), .B(n5076), .Z(n5078) );
  NANDN U6082 ( .A(n5071), .B(sreg[2024]), .Z(n5075) );
  NAND U6083 ( .A(n5073), .B(n5072), .Z(n5074) );
  NAND U6084 ( .A(n5075), .B(n5074), .Z(n5077) );
  XOR U6085 ( .A(n5078), .B(n5077), .Z(c[2025]) );
  NAND U6086 ( .A(b[0]), .B(a[1003]), .Z(n5081) );
  XNOR U6087 ( .A(sreg[2026]), .B(n5081), .Z(n5083) );
  NANDN U6088 ( .A(n5076), .B(sreg[2025]), .Z(n5080) );
  NAND U6089 ( .A(n5078), .B(n5077), .Z(n5079) );
  NAND U6090 ( .A(n5080), .B(n5079), .Z(n5082) );
  XOR U6091 ( .A(n5083), .B(n5082), .Z(c[2026]) );
  NAND U6092 ( .A(b[0]), .B(a[1004]), .Z(n5086) );
  XNOR U6093 ( .A(sreg[2027]), .B(n5086), .Z(n5088) );
  NANDN U6094 ( .A(n5081), .B(sreg[2026]), .Z(n5085) );
  NAND U6095 ( .A(n5083), .B(n5082), .Z(n5084) );
  NAND U6096 ( .A(n5085), .B(n5084), .Z(n5087) );
  XOR U6097 ( .A(n5088), .B(n5087), .Z(c[2027]) );
  NAND U6098 ( .A(b[0]), .B(a[1005]), .Z(n5091) );
  XNOR U6099 ( .A(sreg[2028]), .B(n5091), .Z(n5093) );
  NANDN U6100 ( .A(n5086), .B(sreg[2027]), .Z(n5090) );
  NAND U6101 ( .A(n5088), .B(n5087), .Z(n5089) );
  NAND U6102 ( .A(n5090), .B(n5089), .Z(n5092) );
  XOR U6103 ( .A(n5093), .B(n5092), .Z(c[2028]) );
  NAND U6104 ( .A(b[0]), .B(a[1006]), .Z(n5096) );
  XNOR U6105 ( .A(sreg[2029]), .B(n5096), .Z(n5098) );
  NANDN U6106 ( .A(n5091), .B(sreg[2028]), .Z(n5095) );
  NAND U6107 ( .A(n5093), .B(n5092), .Z(n5094) );
  NAND U6108 ( .A(n5095), .B(n5094), .Z(n5097) );
  XOR U6109 ( .A(n5098), .B(n5097), .Z(c[2029]) );
  NAND U6110 ( .A(b[0]), .B(a[1007]), .Z(n5101) );
  XNOR U6111 ( .A(sreg[2030]), .B(n5101), .Z(n5103) );
  NANDN U6112 ( .A(n5096), .B(sreg[2029]), .Z(n5100) );
  NAND U6113 ( .A(n5098), .B(n5097), .Z(n5099) );
  NAND U6114 ( .A(n5100), .B(n5099), .Z(n5102) );
  XOR U6115 ( .A(n5103), .B(n5102), .Z(c[2030]) );
  NAND U6116 ( .A(b[0]), .B(a[1008]), .Z(n5106) );
  XNOR U6117 ( .A(sreg[2031]), .B(n5106), .Z(n5108) );
  NANDN U6118 ( .A(n5101), .B(sreg[2030]), .Z(n5105) );
  NAND U6119 ( .A(n5103), .B(n5102), .Z(n5104) );
  NAND U6120 ( .A(n5105), .B(n5104), .Z(n5107) );
  XOR U6121 ( .A(n5108), .B(n5107), .Z(c[2031]) );
  NAND U6122 ( .A(b[0]), .B(a[1009]), .Z(n5111) );
  XNOR U6123 ( .A(sreg[2032]), .B(n5111), .Z(n5113) );
  NANDN U6124 ( .A(n5106), .B(sreg[2031]), .Z(n5110) );
  NAND U6125 ( .A(n5108), .B(n5107), .Z(n5109) );
  NAND U6126 ( .A(n5110), .B(n5109), .Z(n5112) );
  XOR U6127 ( .A(n5113), .B(n5112), .Z(c[2032]) );
  NAND U6128 ( .A(b[0]), .B(a[1010]), .Z(n5116) );
  XNOR U6129 ( .A(sreg[2033]), .B(n5116), .Z(n5118) );
  NANDN U6130 ( .A(n5111), .B(sreg[2032]), .Z(n5115) );
  NAND U6131 ( .A(n5113), .B(n5112), .Z(n5114) );
  NAND U6132 ( .A(n5115), .B(n5114), .Z(n5117) );
  XOR U6133 ( .A(n5118), .B(n5117), .Z(c[2033]) );
  NAND U6134 ( .A(b[0]), .B(a[1011]), .Z(n5121) );
  XNOR U6135 ( .A(sreg[2034]), .B(n5121), .Z(n5123) );
  NANDN U6136 ( .A(n5116), .B(sreg[2033]), .Z(n5120) );
  NAND U6137 ( .A(n5118), .B(n5117), .Z(n5119) );
  NAND U6138 ( .A(n5120), .B(n5119), .Z(n5122) );
  XOR U6139 ( .A(n5123), .B(n5122), .Z(c[2034]) );
  NAND U6140 ( .A(b[0]), .B(a[1012]), .Z(n5126) );
  XNOR U6141 ( .A(sreg[2035]), .B(n5126), .Z(n5128) );
  NANDN U6142 ( .A(n5121), .B(sreg[2034]), .Z(n5125) );
  NAND U6143 ( .A(n5123), .B(n5122), .Z(n5124) );
  NAND U6144 ( .A(n5125), .B(n5124), .Z(n5127) );
  XOR U6145 ( .A(n5128), .B(n5127), .Z(c[2035]) );
  NAND U6146 ( .A(b[0]), .B(a[1013]), .Z(n5131) );
  XNOR U6147 ( .A(sreg[2036]), .B(n5131), .Z(n5133) );
  NANDN U6148 ( .A(n5126), .B(sreg[2035]), .Z(n5130) );
  NAND U6149 ( .A(n5128), .B(n5127), .Z(n5129) );
  NAND U6150 ( .A(n5130), .B(n5129), .Z(n5132) );
  XOR U6151 ( .A(n5133), .B(n5132), .Z(c[2036]) );
  NAND U6152 ( .A(b[0]), .B(a[1014]), .Z(n5136) );
  XNOR U6153 ( .A(sreg[2037]), .B(n5136), .Z(n5138) );
  NANDN U6154 ( .A(n5131), .B(sreg[2036]), .Z(n5135) );
  NAND U6155 ( .A(n5133), .B(n5132), .Z(n5134) );
  NAND U6156 ( .A(n5135), .B(n5134), .Z(n5137) );
  XOR U6157 ( .A(n5138), .B(n5137), .Z(c[2037]) );
  NAND U6158 ( .A(b[0]), .B(a[1015]), .Z(n5141) );
  XNOR U6159 ( .A(sreg[2038]), .B(n5141), .Z(n5143) );
  NANDN U6160 ( .A(n5136), .B(sreg[2037]), .Z(n5140) );
  NAND U6161 ( .A(n5138), .B(n5137), .Z(n5139) );
  NAND U6162 ( .A(n5140), .B(n5139), .Z(n5142) );
  XOR U6163 ( .A(n5143), .B(n5142), .Z(c[2038]) );
  NAND U6164 ( .A(b[0]), .B(a[1016]), .Z(n5146) );
  XNOR U6165 ( .A(sreg[2039]), .B(n5146), .Z(n5148) );
  NANDN U6166 ( .A(n5141), .B(sreg[2038]), .Z(n5145) );
  NAND U6167 ( .A(n5143), .B(n5142), .Z(n5144) );
  NAND U6168 ( .A(n5145), .B(n5144), .Z(n5147) );
  XOR U6169 ( .A(n5148), .B(n5147), .Z(c[2039]) );
  NAND U6170 ( .A(b[0]), .B(a[1017]), .Z(n5151) );
  XNOR U6171 ( .A(sreg[2040]), .B(n5151), .Z(n5153) );
  NANDN U6172 ( .A(n5146), .B(sreg[2039]), .Z(n5150) );
  NAND U6173 ( .A(n5148), .B(n5147), .Z(n5149) );
  AND U6174 ( .A(n5150), .B(n5149), .Z(n5152) );
  XNOR U6175 ( .A(n5153), .B(n5152), .Z(c[2040]) );
  NANDN U6176 ( .A(sreg[2040]), .B(n5151), .Z(n5155) );
  NAND U6177 ( .A(n5153), .B(n5152), .Z(n5154) );
  AND U6178 ( .A(n5155), .B(n5154), .Z(n5158) );
  NAND U6179 ( .A(b[0]), .B(a[1018]), .Z(n5156) );
  XNOR U6180 ( .A(sreg[2041]), .B(n5156), .Z(n5157) );
  XOR U6181 ( .A(n5158), .B(n5157), .Z(c[2041]) );
  NANDN U6182 ( .A(n5156), .B(sreg[2041]), .Z(n5160) );
  NAND U6183 ( .A(n5158), .B(n5157), .Z(n5159) );
  AND U6184 ( .A(n5160), .B(n5159), .Z(n5163) );
  NAND U6185 ( .A(b[0]), .B(a[1019]), .Z(n5161) );
  XNOR U6186 ( .A(sreg[2042]), .B(n5161), .Z(n5162) );
  XNOR U6187 ( .A(n5163), .B(n5162), .Z(c[2042]) );
  NAND U6188 ( .A(b[0]), .B(a[1020]), .Z(n5166) );
  XNOR U6189 ( .A(sreg[2043]), .B(n5166), .Z(n5168) );
  NANDN U6190 ( .A(sreg[2042]), .B(n5161), .Z(n5165) );
  NAND U6191 ( .A(n5163), .B(n5162), .Z(n5164) );
  NAND U6192 ( .A(n5165), .B(n5164), .Z(n5167) );
  XNOR U6193 ( .A(n5168), .B(n5167), .Z(c[2043]) );
  NANDN U6194 ( .A(sreg[2043]), .B(n5166), .Z(n5170) );
  NAND U6195 ( .A(n5168), .B(n5167), .Z(n5169) );
  AND U6196 ( .A(n5170), .B(n5169), .Z(n5173) );
  NAND U6197 ( .A(b[0]), .B(a[1021]), .Z(n5171) );
  XNOR U6198 ( .A(sreg[2044]), .B(n5171), .Z(n5172) );
  XOR U6199 ( .A(n5173), .B(n5172), .Z(c[2044]) );
  NANDN U6200 ( .A(n5171), .B(sreg[2044]), .Z(n5175) );
  NAND U6201 ( .A(n5173), .B(n5172), .Z(n5174) );
  AND U6202 ( .A(n5175), .B(n5174), .Z(n5178) );
  NAND U6203 ( .A(b[0]), .B(a[1022]), .Z(n5176) );
  XNOR U6204 ( .A(sreg[2045]), .B(n5176), .Z(n5177) );
  XNOR U6205 ( .A(n5178), .B(n5177), .Z(c[2045]) );
  NANDN U6206 ( .A(sreg[2045]), .B(n5176), .Z(n5180) );
  NAND U6207 ( .A(n5178), .B(n5177), .Z(n5179) );
  AND U6208 ( .A(n5180), .B(n5179), .Z(n5183) );
  NAND U6209 ( .A(b[0]), .B(a[1023]), .Z(n5182) );
  XOR U6210 ( .A(n5182), .B(sreg[2046]), .Z(n5181) );
  XNOR U6211 ( .A(n5183), .B(n5181), .Z(c[2046]) );
endmodule

