
module mult_N128_CC16 ( clk, rst, a, b, c );
  input [127:0] a;
  input [7:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671;
  wire   [127:8] swire;
  wire   [255:128] sreg;

  DFF \sreg_reg[128]  ( .D(swire[8]), .CLK(clk), .RST(rst), .Q(sreg[128]) );
  DFF \sreg_reg[129]  ( .D(swire[9]), .CLK(clk), .RST(rst), .Q(sreg[129]) );
  DFF \sreg_reg[130]  ( .D(swire[10]), .CLK(clk), .RST(rst), .Q(sreg[130]) );
  DFF \sreg_reg[131]  ( .D(swire[11]), .CLK(clk), .RST(rst), .Q(sreg[131]) );
  DFF \sreg_reg[132]  ( .D(swire[12]), .CLK(clk), .RST(rst), .Q(sreg[132]) );
  DFF \sreg_reg[133]  ( .D(swire[13]), .CLK(clk), .RST(rst), .Q(sreg[133]) );
  DFF \sreg_reg[134]  ( .D(swire[14]), .CLK(clk), .RST(rst), .Q(sreg[134]) );
  DFF \sreg_reg[135]  ( .D(swire[15]), .CLK(clk), .RST(rst), .Q(sreg[135]) );
  DFF \sreg_reg[136]  ( .D(swire[16]), .CLK(clk), .RST(rst), .Q(sreg[136]) );
  DFF \sreg_reg[137]  ( .D(swire[17]), .CLK(clk), .RST(rst), .Q(sreg[137]) );
  DFF \sreg_reg[138]  ( .D(swire[18]), .CLK(clk), .RST(rst), .Q(sreg[138]) );
  DFF \sreg_reg[139]  ( .D(swire[19]), .CLK(clk), .RST(rst), .Q(sreg[139]) );
  DFF \sreg_reg[140]  ( .D(swire[20]), .CLK(clk), .RST(rst), .Q(sreg[140]) );
  DFF \sreg_reg[141]  ( .D(swire[21]), .CLK(clk), .RST(rst), .Q(sreg[141]) );
  DFF \sreg_reg[142]  ( .D(swire[22]), .CLK(clk), .RST(rst), .Q(sreg[142]) );
  DFF \sreg_reg[143]  ( .D(swire[23]), .CLK(clk), .RST(rst), .Q(sreg[143]) );
  DFF \sreg_reg[144]  ( .D(swire[24]), .CLK(clk), .RST(rst), .Q(sreg[144]) );
  DFF \sreg_reg[145]  ( .D(swire[25]), .CLK(clk), .RST(rst), .Q(sreg[145]) );
  DFF \sreg_reg[146]  ( .D(swire[26]), .CLK(clk), .RST(rst), .Q(sreg[146]) );
  DFF \sreg_reg[147]  ( .D(swire[27]), .CLK(clk), .RST(rst), .Q(sreg[147]) );
  DFF \sreg_reg[148]  ( .D(swire[28]), .CLK(clk), .RST(rst), .Q(sreg[148]) );
  DFF \sreg_reg[149]  ( .D(swire[29]), .CLK(clk), .RST(rst), .Q(sreg[149]) );
  DFF \sreg_reg[150]  ( .D(swire[30]), .CLK(clk), .RST(rst), .Q(sreg[150]) );
  DFF \sreg_reg[151]  ( .D(swire[31]), .CLK(clk), .RST(rst), .Q(sreg[151]) );
  DFF \sreg_reg[152]  ( .D(swire[32]), .CLK(clk), .RST(rst), .Q(sreg[152]) );
  DFF \sreg_reg[153]  ( .D(swire[33]), .CLK(clk), .RST(rst), .Q(sreg[153]) );
  DFF \sreg_reg[154]  ( .D(swire[34]), .CLK(clk), .RST(rst), .Q(sreg[154]) );
  DFF \sreg_reg[155]  ( .D(swire[35]), .CLK(clk), .RST(rst), .Q(sreg[155]) );
  DFF \sreg_reg[156]  ( .D(swire[36]), .CLK(clk), .RST(rst), .Q(sreg[156]) );
  DFF \sreg_reg[157]  ( .D(swire[37]), .CLK(clk), .RST(rst), .Q(sreg[157]) );
  DFF \sreg_reg[158]  ( .D(swire[38]), .CLK(clk), .RST(rst), .Q(sreg[158]) );
  DFF \sreg_reg[159]  ( .D(swire[39]), .CLK(clk), .RST(rst), .Q(sreg[159]) );
  DFF \sreg_reg[160]  ( .D(swire[40]), .CLK(clk), .RST(rst), .Q(sreg[160]) );
  DFF \sreg_reg[161]  ( .D(swire[41]), .CLK(clk), .RST(rst), .Q(sreg[161]) );
  DFF \sreg_reg[162]  ( .D(swire[42]), .CLK(clk), .RST(rst), .Q(sreg[162]) );
  DFF \sreg_reg[163]  ( .D(swire[43]), .CLK(clk), .RST(rst), .Q(sreg[163]) );
  DFF \sreg_reg[164]  ( .D(swire[44]), .CLK(clk), .RST(rst), .Q(sreg[164]) );
  DFF \sreg_reg[165]  ( .D(swire[45]), .CLK(clk), .RST(rst), .Q(sreg[165]) );
  DFF \sreg_reg[166]  ( .D(swire[46]), .CLK(clk), .RST(rst), .Q(sreg[166]) );
  DFF \sreg_reg[167]  ( .D(swire[47]), .CLK(clk), .RST(rst), .Q(sreg[167]) );
  DFF \sreg_reg[168]  ( .D(swire[48]), .CLK(clk), .RST(rst), .Q(sreg[168]) );
  DFF \sreg_reg[169]  ( .D(swire[49]), .CLK(clk), .RST(rst), .Q(sreg[169]) );
  DFF \sreg_reg[170]  ( .D(swire[50]), .CLK(clk), .RST(rst), .Q(sreg[170]) );
  DFF \sreg_reg[171]  ( .D(swire[51]), .CLK(clk), .RST(rst), .Q(sreg[171]) );
  DFF \sreg_reg[172]  ( .D(swire[52]), .CLK(clk), .RST(rst), .Q(sreg[172]) );
  DFF \sreg_reg[173]  ( .D(swire[53]), .CLK(clk), .RST(rst), .Q(sreg[173]) );
  DFF \sreg_reg[174]  ( .D(swire[54]), .CLK(clk), .RST(rst), .Q(sreg[174]) );
  DFF \sreg_reg[175]  ( .D(swire[55]), .CLK(clk), .RST(rst), .Q(sreg[175]) );
  DFF \sreg_reg[176]  ( .D(swire[56]), .CLK(clk), .RST(rst), .Q(sreg[176]) );
  DFF \sreg_reg[177]  ( .D(swire[57]), .CLK(clk), .RST(rst), .Q(sreg[177]) );
  DFF \sreg_reg[178]  ( .D(swire[58]), .CLK(clk), .RST(rst), .Q(sreg[178]) );
  DFF \sreg_reg[179]  ( .D(swire[59]), .CLK(clk), .RST(rst), .Q(sreg[179]) );
  DFF \sreg_reg[180]  ( .D(swire[60]), .CLK(clk), .RST(rst), .Q(sreg[180]) );
  DFF \sreg_reg[181]  ( .D(swire[61]), .CLK(clk), .RST(rst), .Q(sreg[181]) );
  DFF \sreg_reg[182]  ( .D(swire[62]), .CLK(clk), .RST(rst), .Q(sreg[182]) );
  DFF \sreg_reg[183]  ( .D(swire[63]), .CLK(clk), .RST(rst), .Q(sreg[183]) );
  DFF \sreg_reg[184]  ( .D(swire[64]), .CLK(clk), .RST(rst), .Q(sreg[184]) );
  DFF \sreg_reg[185]  ( .D(swire[65]), .CLK(clk), .RST(rst), .Q(sreg[185]) );
  DFF \sreg_reg[186]  ( .D(swire[66]), .CLK(clk), .RST(rst), .Q(sreg[186]) );
  DFF \sreg_reg[187]  ( .D(swire[67]), .CLK(clk), .RST(rst), .Q(sreg[187]) );
  DFF \sreg_reg[188]  ( .D(swire[68]), .CLK(clk), .RST(rst), .Q(sreg[188]) );
  DFF \sreg_reg[189]  ( .D(swire[69]), .CLK(clk), .RST(rst), .Q(sreg[189]) );
  DFF \sreg_reg[190]  ( .D(swire[70]), .CLK(clk), .RST(rst), .Q(sreg[190]) );
  DFF \sreg_reg[191]  ( .D(swire[71]), .CLK(clk), .RST(rst), .Q(sreg[191]) );
  DFF \sreg_reg[192]  ( .D(swire[72]), .CLK(clk), .RST(rst), .Q(sreg[192]) );
  DFF \sreg_reg[193]  ( .D(swire[73]), .CLK(clk), .RST(rst), .Q(sreg[193]) );
  DFF \sreg_reg[194]  ( .D(swire[74]), .CLK(clk), .RST(rst), .Q(sreg[194]) );
  DFF \sreg_reg[195]  ( .D(swire[75]), .CLK(clk), .RST(rst), .Q(sreg[195]) );
  DFF \sreg_reg[196]  ( .D(swire[76]), .CLK(clk), .RST(rst), .Q(sreg[196]) );
  DFF \sreg_reg[197]  ( .D(swire[77]), .CLK(clk), .RST(rst), .Q(sreg[197]) );
  DFF \sreg_reg[198]  ( .D(swire[78]), .CLK(clk), .RST(rst), .Q(sreg[198]) );
  DFF \sreg_reg[199]  ( .D(swire[79]), .CLK(clk), .RST(rst), .Q(sreg[199]) );
  DFF \sreg_reg[200]  ( .D(swire[80]), .CLK(clk), .RST(rst), .Q(sreg[200]) );
  DFF \sreg_reg[201]  ( .D(swire[81]), .CLK(clk), .RST(rst), .Q(sreg[201]) );
  DFF \sreg_reg[202]  ( .D(swire[82]), .CLK(clk), .RST(rst), .Q(sreg[202]) );
  DFF \sreg_reg[203]  ( .D(swire[83]), .CLK(clk), .RST(rst), .Q(sreg[203]) );
  DFF \sreg_reg[204]  ( .D(swire[84]), .CLK(clk), .RST(rst), .Q(sreg[204]) );
  DFF \sreg_reg[205]  ( .D(swire[85]), .CLK(clk), .RST(rst), .Q(sreg[205]) );
  DFF \sreg_reg[206]  ( .D(swire[86]), .CLK(clk), .RST(rst), .Q(sreg[206]) );
  DFF \sreg_reg[207]  ( .D(swire[87]), .CLK(clk), .RST(rst), .Q(sreg[207]) );
  DFF \sreg_reg[208]  ( .D(swire[88]), .CLK(clk), .RST(rst), .Q(sreg[208]) );
  DFF \sreg_reg[209]  ( .D(swire[89]), .CLK(clk), .RST(rst), .Q(sreg[209]) );
  DFF \sreg_reg[210]  ( .D(swire[90]), .CLK(clk), .RST(rst), .Q(sreg[210]) );
  DFF \sreg_reg[211]  ( .D(swire[91]), .CLK(clk), .RST(rst), .Q(sreg[211]) );
  DFF \sreg_reg[212]  ( .D(swire[92]), .CLK(clk), .RST(rst), .Q(sreg[212]) );
  DFF \sreg_reg[213]  ( .D(swire[93]), .CLK(clk), .RST(rst), .Q(sreg[213]) );
  DFF \sreg_reg[214]  ( .D(swire[94]), .CLK(clk), .RST(rst), .Q(sreg[214]) );
  DFF \sreg_reg[215]  ( .D(swire[95]), .CLK(clk), .RST(rst), .Q(sreg[215]) );
  DFF \sreg_reg[216]  ( .D(swire[96]), .CLK(clk), .RST(rst), .Q(sreg[216]) );
  DFF \sreg_reg[217]  ( .D(swire[97]), .CLK(clk), .RST(rst), .Q(sreg[217]) );
  DFF \sreg_reg[218]  ( .D(swire[98]), .CLK(clk), .RST(rst), .Q(sreg[218]) );
  DFF \sreg_reg[219]  ( .D(swire[99]), .CLK(clk), .RST(rst), .Q(sreg[219]) );
  DFF \sreg_reg[220]  ( .D(swire[100]), .CLK(clk), .RST(rst), .Q(sreg[220]) );
  DFF \sreg_reg[221]  ( .D(swire[101]), .CLK(clk), .RST(rst), .Q(sreg[221]) );
  DFF \sreg_reg[222]  ( .D(swire[102]), .CLK(clk), .RST(rst), .Q(sreg[222]) );
  DFF \sreg_reg[223]  ( .D(swire[103]), .CLK(clk), .RST(rst), .Q(sreg[223]) );
  DFF \sreg_reg[224]  ( .D(swire[104]), .CLK(clk), .RST(rst), .Q(sreg[224]) );
  DFF \sreg_reg[225]  ( .D(swire[105]), .CLK(clk), .RST(rst), .Q(sreg[225]) );
  DFF \sreg_reg[226]  ( .D(swire[106]), .CLK(clk), .RST(rst), .Q(sreg[226]) );
  DFF \sreg_reg[227]  ( .D(swire[107]), .CLK(clk), .RST(rst), .Q(sreg[227]) );
  DFF \sreg_reg[228]  ( .D(swire[108]), .CLK(clk), .RST(rst), .Q(sreg[228]) );
  DFF \sreg_reg[229]  ( .D(swire[109]), .CLK(clk), .RST(rst), .Q(sreg[229]) );
  DFF \sreg_reg[230]  ( .D(swire[110]), .CLK(clk), .RST(rst), .Q(sreg[230]) );
  DFF \sreg_reg[231]  ( .D(swire[111]), .CLK(clk), .RST(rst), .Q(sreg[231]) );
  DFF \sreg_reg[232]  ( .D(swire[112]), .CLK(clk), .RST(rst), .Q(sreg[232]) );
  DFF \sreg_reg[233]  ( .D(swire[113]), .CLK(clk), .RST(rst), .Q(sreg[233]) );
  DFF \sreg_reg[234]  ( .D(swire[114]), .CLK(clk), .RST(rst), .Q(sreg[234]) );
  DFF \sreg_reg[235]  ( .D(swire[115]), .CLK(clk), .RST(rst), .Q(sreg[235]) );
  DFF \sreg_reg[236]  ( .D(swire[116]), .CLK(clk), .RST(rst), .Q(sreg[236]) );
  DFF \sreg_reg[237]  ( .D(swire[117]), .CLK(clk), .RST(rst), .Q(sreg[237]) );
  DFF \sreg_reg[238]  ( .D(swire[118]), .CLK(clk), .RST(rst), .Q(sreg[238]) );
  DFF \sreg_reg[239]  ( .D(swire[119]), .CLK(clk), .RST(rst), .Q(sreg[239]) );
  DFF \sreg_reg[240]  ( .D(swire[120]), .CLK(clk), .RST(rst), .Q(sreg[240]) );
  DFF \sreg_reg[241]  ( .D(swire[121]), .CLK(clk), .RST(rst), .Q(sreg[241]) );
  DFF \sreg_reg[242]  ( .D(swire[122]), .CLK(clk), .RST(rst), .Q(sreg[242]) );
  DFF \sreg_reg[243]  ( .D(swire[123]), .CLK(clk), .RST(rst), .Q(sreg[243]) );
  DFF \sreg_reg[244]  ( .D(swire[124]), .CLK(clk), .RST(rst), .Q(sreg[244]) );
  DFF \sreg_reg[245]  ( .D(swire[125]), .CLK(clk), .RST(rst), .Q(sreg[245]) );
  DFF \sreg_reg[246]  ( .D(swire[126]), .CLK(clk), .RST(rst), .Q(sreg[246]) );
  DFF \sreg_reg[247]  ( .D(swire[127]), .CLK(clk), .RST(rst), .Q(sreg[247]) );
  DFF \sreg_reg[127]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[126]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[125]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[124]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[123]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[122]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[121]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[120]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[119]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[118]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[117]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[116]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[115]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[114]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[113]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[112]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[111]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[110]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[109]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[108]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[107]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[106]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[105]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[104]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[103]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[102]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[101]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[100]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[99]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[98]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[97]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[96]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[95]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[94]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[93]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[92]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[91]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[90]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[89]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[88]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[87]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[86]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[85]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[84]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[83]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[82]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[81]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[80]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[79]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[78]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[77]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[76]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[75]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[74]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[73]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[72]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[71]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[70]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[69]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[68]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[67]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[66]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[65]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[64]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[63]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[62]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[61]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[60]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[59]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[58]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[57]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[56]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[55]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[54]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[53]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[52]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[51]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[50]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[49]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[48]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[47]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[46]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[45]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[44]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[43]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[42]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[41]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[40]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[39]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[38]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[37]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[36]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[35]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[34]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[33]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[32]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[31]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[30]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[29]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[28]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[27]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[26]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[25]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[24]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[23]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[22]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[21]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[20]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[19]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[18]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[17]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[16]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[15]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[14]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[13]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[12]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[11]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[10]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[9]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[8]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[0]) );
  XNOR U11 ( .A(n1731), .B(n1747), .Z(n1727) );
  XOR U12 ( .A(n1631), .B(n1651), .Z(n1636) );
  XOR U13 ( .A(n1663), .B(n1683), .Z(n1668) );
  XOR U14 ( .A(n1758), .B(n1778), .Z(n1764) );
  XOR U15 ( .A(n1868), .B(n1874), .Z(n1847) );
  XOR U16 ( .A(n1900), .B(n1906), .Z(n1879) );
  XOR U17 ( .A(n1980), .B(n2000), .Z(n1986) );
  XOR U18 ( .A(n2090), .B(n2096), .Z(n2069) );
  XOR U19 ( .A(n2122), .B(n2128), .Z(n2101) );
  XOR U20 ( .A(n2202), .B(n2222), .Z(n2208) );
  XOR U21 ( .A(n2312), .B(n2318), .Z(n2291) );
  XOR U22 ( .A(n2344), .B(n2350), .Z(n2323) );
  XOR U23 ( .A(n2424), .B(n2444), .Z(n2430) );
  XOR U24 ( .A(n2534), .B(n2540), .Z(n2513) );
  XOR U25 ( .A(n2566), .B(n2572), .Z(n2545) );
  XOR U26 ( .A(n2646), .B(n2666), .Z(n2652) );
  XOR U27 ( .A(n2756), .B(n2762), .Z(n2735) );
  XOR U28 ( .A(n2788), .B(n2794), .Z(n2767) );
  XOR U29 ( .A(n2868), .B(n2888), .Z(n2874) );
  XOR U30 ( .A(n2978), .B(n2984), .Z(n2957) );
  XOR U31 ( .A(n3010), .B(n3016), .Z(n2989) );
  XOR U32 ( .A(n3090), .B(n3110), .Z(n3096) );
  XOR U33 ( .A(n3200), .B(n3206), .Z(n3179) );
  XOR U34 ( .A(n3232), .B(n3238), .Z(n3211) );
  XOR U35 ( .A(n3312), .B(n3332), .Z(n3318) );
  XOR U36 ( .A(n3422), .B(n3428), .Z(n3401) );
  XOR U37 ( .A(n3454), .B(n3460), .Z(n3433) );
  XOR U38 ( .A(n3534), .B(n3554), .Z(n3540) );
  XOR U39 ( .A(n3644), .B(n3650), .Z(n3623) );
  XOR U40 ( .A(n3676), .B(n3682), .Z(n3655) );
  XOR U41 ( .A(n3756), .B(n3776), .Z(n3762) );
  XOR U42 ( .A(n3866), .B(n3872), .Z(n3845) );
  XOR U43 ( .A(n3898), .B(n3904), .Z(n3877) );
  XOR U44 ( .A(n3978), .B(n3998), .Z(n3984) );
  XOR U45 ( .A(n4088), .B(n4094), .Z(n4067) );
  XOR U46 ( .A(n4120), .B(n4126), .Z(n4099) );
  XOR U47 ( .A(n4200), .B(n4220), .Z(n4206) );
  XOR U48 ( .A(n4310), .B(n4316), .Z(n4289) );
  XOR U49 ( .A(n4342), .B(n4348), .Z(n4321) );
  XOR U50 ( .A(n4453), .B(n4473), .Z(n4459) );
  XNOR U51 ( .A(n4551), .B(n4571), .Z(n4559) );
  XOR U52 ( .A(n1789), .B(n1809), .Z(n1795) );
  XOR U53 ( .A(n2011), .B(n2031), .Z(n2017) );
  XOR U54 ( .A(n2233), .B(n2253), .Z(n2239) );
  XOR U55 ( .A(n2455), .B(n2475), .Z(n2461) );
  XOR U56 ( .A(n2677), .B(n2697), .Z(n2683) );
  XOR U57 ( .A(n2899), .B(n2919), .Z(n2905) );
  XOR U58 ( .A(n3121), .B(n3141), .Z(n3127) );
  XOR U59 ( .A(n3343), .B(n3363), .Z(n3349) );
  XOR U60 ( .A(n3565), .B(n3585), .Z(n3571) );
  XOR U61 ( .A(n3787), .B(n3807), .Z(n3793) );
  XOR U62 ( .A(n4009), .B(n4029), .Z(n4015) );
  XOR U63 ( .A(n4231), .B(n4251), .Z(n4237) );
  XNOR U64 ( .A(n4395), .B(n4411), .Z(n4391) );
  XNOR U65 ( .A(n4586), .B(n4607), .Z(n4595) );
  XNOR U66 ( .A(n4522), .B(n4533), .Z(n4504) );
  XOR U67 ( .A(n1637), .B(n1642), .Z(n1614) );
  XOR U68 ( .A(n1700), .B(n1706), .Z(n1679) );
  XNOR U69 ( .A(n1773), .B(n1763), .Z(n1743) );
  XOR U70 ( .A(n1888), .B(n1878), .Z(n1852) );
  XNOR U71 ( .A(n1995), .B(n1985), .Z(n1965) );
  XOR U72 ( .A(n2110), .B(n2100), .Z(n2074) );
  XNOR U73 ( .A(n2217), .B(n2207), .Z(n2187) );
  XOR U74 ( .A(n2332), .B(n2322), .Z(n2296) );
  XNOR U75 ( .A(n2439), .B(n2429), .Z(n2409) );
  XOR U76 ( .A(n2554), .B(n2544), .Z(n2518) );
  XNOR U77 ( .A(n2661), .B(n2651), .Z(n2631) );
  XOR U78 ( .A(n2776), .B(n2766), .Z(n2740) );
  XNOR U79 ( .A(n2883), .B(n2873), .Z(n2853) );
  XOR U80 ( .A(n2998), .B(n2988), .Z(n2962) );
  XNOR U81 ( .A(n3105), .B(n3095), .Z(n3075) );
  XOR U82 ( .A(n3220), .B(n3210), .Z(n3184) );
  XNOR U83 ( .A(n3327), .B(n3317), .Z(n3297) );
  XOR U84 ( .A(n3442), .B(n3432), .Z(n3406) );
  XNOR U85 ( .A(n3549), .B(n3539), .Z(n3519) );
  XOR U86 ( .A(n3664), .B(n3654), .Z(n3628) );
  XNOR U87 ( .A(n3771), .B(n3761), .Z(n3741) );
  XOR U88 ( .A(n3886), .B(n3876), .Z(n3850) );
  XNOR U89 ( .A(n3993), .B(n3983), .Z(n3963) );
  XOR U90 ( .A(n4108), .B(n4098), .Z(n4072) );
  XNOR U91 ( .A(n4215), .B(n4205), .Z(n4185) );
  XOR U92 ( .A(n4298), .B(n4288), .Z(n4274) );
  XOR U93 ( .A(n4362), .B(n4352), .Z(n4326) );
  XNOR U94 ( .A(n4468), .B(n4458), .Z(n4433) );
  XOR U95 ( .A(n863), .B(n890), .Z(n868) );
  XOR U96 ( .A(n939), .B(n966), .Z(n944) );
  XOR U97 ( .A(n1015), .B(n1042), .Z(n1020) );
  XOR U98 ( .A(n1091), .B(n1578), .Z(n1096) );
  XNOR U99 ( .A(n1953), .B(n1969), .Z(n1949) );
  XNOR U100 ( .A(n2175), .B(n2191), .Z(n2171) );
  XNOR U101 ( .A(n2397), .B(n2413), .Z(n2393) );
  XNOR U102 ( .A(n2619), .B(n2635), .Z(n2615) );
  XNOR U103 ( .A(n2841), .B(n2857), .Z(n2837) );
  XNOR U104 ( .A(n3063), .B(n3079), .Z(n3059) );
  XNOR U105 ( .A(n3285), .B(n3301), .Z(n3281) );
  XNOR U106 ( .A(n3507), .B(n3523), .Z(n3503) );
  XNOR U107 ( .A(n3729), .B(n3745), .Z(n3725) );
  XNOR U108 ( .A(n3951), .B(n3967), .Z(n3947) );
  XNOR U109 ( .A(n4173), .B(n4189), .Z(n4169) );
  XOR U110 ( .A(n1669), .B(n1674), .Z(n1647) );
  XOR U111 ( .A(n1727), .B(n1737), .Z(n1711) );
  XNOR U112 ( .A(n1804), .B(n1794), .Z(n1769) );
  XOR U113 ( .A(n1856), .B(n1846), .Z(n1832) );
  XNOR U114 ( .A(n1909), .B(n1908), .Z(n1885) );
  XNOR U115 ( .A(n1958), .B(n1957), .Z(n1917) );
  XNOR U116 ( .A(n2026), .B(n2016), .Z(n1991) );
  XOR U117 ( .A(n2078), .B(n2068), .Z(n2054) );
  XNOR U118 ( .A(n2131), .B(n2130), .Z(n2107) );
  XNOR U119 ( .A(n2180), .B(n2179), .Z(n2139) );
  XNOR U120 ( .A(n2248), .B(n2238), .Z(n2213) );
  XOR U121 ( .A(n2300), .B(n2290), .Z(n2276) );
  XNOR U122 ( .A(n2353), .B(n2352), .Z(n2329) );
  XNOR U123 ( .A(n2402), .B(n2401), .Z(n2361) );
  XNOR U124 ( .A(n2470), .B(n2460), .Z(n2435) );
  XOR U125 ( .A(n2522), .B(n2512), .Z(n2498) );
  XNOR U126 ( .A(n2575), .B(n2574), .Z(n2551) );
  XNOR U127 ( .A(n2624), .B(n2623), .Z(n2583) );
  XNOR U128 ( .A(n2692), .B(n2682), .Z(n2657) );
  XOR U129 ( .A(n2744), .B(n2734), .Z(n2720) );
  XNOR U130 ( .A(n2797), .B(n2796), .Z(n2773) );
  XNOR U131 ( .A(n2846), .B(n2845), .Z(n2805) );
  XNOR U132 ( .A(n2914), .B(n2904), .Z(n2879) );
  XOR U133 ( .A(n2966), .B(n2956), .Z(n2942) );
  XNOR U134 ( .A(n3019), .B(n3018), .Z(n2995) );
  XNOR U135 ( .A(n3068), .B(n3067), .Z(n3027) );
  XNOR U136 ( .A(n3136), .B(n3126), .Z(n3101) );
  XOR U137 ( .A(n3188), .B(n3178), .Z(n3164) );
  XNOR U138 ( .A(n3241), .B(n3240), .Z(n3217) );
  XNOR U139 ( .A(n3290), .B(n3289), .Z(n3249) );
  XNOR U140 ( .A(n3358), .B(n3348), .Z(n3323) );
  XOR U141 ( .A(n3410), .B(n3400), .Z(n3386) );
  XNOR U142 ( .A(n3463), .B(n3462), .Z(n3439) );
  XNOR U143 ( .A(n3512), .B(n3511), .Z(n3471) );
  XNOR U144 ( .A(n3580), .B(n3570), .Z(n3545) );
  XOR U145 ( .A(n3632), .B(n3622), .Z(n3608) );
  XNOR U146 ( .A(n3685), .B(n3684), .Z(n3661) );
  XNOR U147 ( .A(n3734), .B(n3733), .Z(n3693) );
  XNOR U148 ( .A(n3802), .B(n3792), .Z(n3767) );
  XOR U149 ( .A(n3854), .B(n3844), .Z(n3830) );
  XNOR U150 ( .A(n3907), .B(n3906), .Z(n3883) );
  XNOR U151 ( .A(n3956), .B(n3955), .Z(n3915) );
  XNOR U152 ( .A(n4024), .B(n4014), .Z(n3989) );
  XOR U153 ( .A(n4076), .B(n4066), .Z(n4052) );
  XNOR U154 ( .A(n4129), .B(n4128), .Z(n4105) );
  XNOR U155 ( .A(n4178), .B(n4177), .Z(n4137) );
  XNOR U156 ( .A(n4246), .B(n4236), .Z(n4211) );
  XOR U157 ( .A(n4330), .B(n4320), .Z(n4294) );
  XNOR U158 ( .A(n4400), .B(n4399), .Z(n4359) );
  XNOR U159 ( .A(n4437), .B(n4427), .Z(n4407) );
  XOR U160 ( .A(n4496), .B(n4490), .Z(n4464) );
  XNOR U161 ( .A(n4622), .B(n4630), .Z(n4618) );
  XNOR U162 ( .A(n4559), .B(n4567), .Z(n4555) );
  AND U163 ( .A(n293), .B(n292), .Z(n260) );
  XOR U164 ( .A(n901), .B(n928), .Z(n906) );
  XOR U165 ( .A(n977), .B(n1004), .Z(n982) );
  XOR U166 ( .A(n1053), .B(n1080), .Z(n1058) );
  XOR U167 ( .A(n1595), .B(n1609), .Z(n1600) );
  XNOR U168 ( .A(n1641), .B(n1640), .Z(n1615) );
  XNOR U169 ( .A(n1673), .B(n1672), .Z(n1648) );
  XNOR U170 ( .A(n1705), .B(n1704), .Z(n1680) );
  XOR U171 ( .A(n1836), .B(n1826), .Z(n1800) );
  XNOR U172 ( .A(n1845), .B(n1844), .Z(n1833) );
  XNOR U173 ( .A(n1877), .B(n1876), .Z(n1853) );
  XOR U174 ( .A(n1920), .B(n1910), .Z(n1884) );
  XOR U175 ( .A(n2058), .B(n2048), .Z(n2022) );
  XNOR U176 ( .A(n2067), .B(n2066), .Z(n2055) );
  XNOR U177 ( .A(n2099), .B(n2098), .Z(n2075) );
  XOR U178 ( .A(n2142), .B(n2132), .Z(n2106) );
  XOR U179 ( .A(n2280), .B(n2270), .Z(n2244) );
  XNOR U180 ( .A(n2289), .B(n2288), .Z(n2277) );
  XNOR U181 ( .A(n2321), .B(n2320), .Z(n2297) );
  XOR U182 ( .A(n2364), .B(n2354), .Z(n2328) );
  XOR U183 ( .A(n2502), .B(n2492), .Z(n2466) );
  XNOR U184 ( .A(n2511), .B(n2510), .Z(n2499) );
  XNOR U185 ( .A(n2543), .B(n2542), .Z(n2519) );
  XOR U186 ( .A(n2586), .B(n2576), .Z(n2550) );
  XOR U187 ( .A(n2724), .B(n2714), .Z(n2688) );
  XNOR U188 ( .A(n2733), .B(n2732), .Z(n2721) );
  XNOR U189 ( .A(n2765), .B(n2764), .Z(n2741) );
  XOR U190 ( .A(n2808), .B(n2798), .Z(n2772) );
  XOR U191 ( .A(n2946), .B(n2936), .Z(n2910) );
  XNOR U192 ( .A(n2955), .B(n2954), .Z(n2943) );
  XNOR U193 ( .A(n2987), .B(n2986), .Z(n2963) );
  XOR U194 ( .A(n3030), .B(n3020), .Z(n2994) );
  XOR U195 ( .A(n3168), .B(n3158), .Z(n3132) );
  XNOR U196 ( .A(n3177), .B(n3176), .Z(n3165) );
  XNOR U197 ( .A(n3209), .B(n3208), .Z(n3185) );
  XOR U198 ( .A(n3252), .B(n3242), .Z(n3216) );
  XOR U199 ( .A(n3390), .B(n3380), .Z(n3354) );
  XNOR U200 ( .A(n3399), .B(n3398), .Z(n3387) );
  XNOR U201 ( .A(n3431), .B(n3430), .Z(n3407) );
  XOR U202 ( .A(n3474), .B(n3464), .Z(n3438) );
  XOR U203 ( .A(n3612), .B(n3602), .Z(n3576) );
  XNOR U204 ( .A(n3621), .B(n3620), .Z(n3609) );
  XNOR U205 ( .A(n3653), .B(n3652), .Z(n3629) );
  XOR U206 ( .A(n3696), .B(n3686), .Z(n3660) );
  XOR U207 ( .A(n3834), .B(n3824), .Z(n3798) );
  XNOR U208 ( .A(n3843), .B(n3842), .Z(n3831) );
  XNOR U209 ( .A(n3875), .B(n3874), .Z(n3851) );
  XOR U210 ( .A(n3918), .B(n3908), .Z(n3882) );
  XOR U211 ( .A(n4056), .B(n4046), .Z(n4020) );
  XNOR U212 ( .A(n4065), .B(n4064), .Z(n4053) );
  XNOR U213 ( .A(n4097), .B(n4096), .Z(n4073) );
  XOR U214 ( .A(n4140), .B(n4130), .Z(n4104) );
  XOR U215 ( .A(n4278), .B(n4268), .Z(n4242) );
  XNOR U216 ( .A(n4287), .B(n4286), .Z(n4275) );
  XNOR U217 ( .A(n4319), .B(n4318), .Z(n4295) );
  XNOR U218 ( .A(n4351), .B(n4350), .Z(n4327) );
  XOR U219 ( .A(n4391), .B(n4401), .Z(n4358) );
  AND U220 ( .A(a[1]), .B(n4656), .Z(n4667) );
  XNOR U221 ( .A(n4595), .B(n4603), .Z(n4591) );
  XNOR U222 ( .A(n4504), .B(n4529), .Z(n4495) );
  XNOR U223 ( .A(n1743), .B(n1741), .Z(n1714) );
  XNOR U224 ( .A(n1965), .B(n1963), .Z(n1919) );
  XNOR U225 ( .A(n2187), .B(n2185), .Z(n2141) );
  XNOR U226 ( .A(n2409), .B(n2407), .Z(n2363) );
  XNOR U227 ( .A(n2631), .B(n2629), .Z(n2585) );
  XNOR U228 ( .A(n2853), .B(n2851), .Z(n2807) );
  XNOR U229 ( .A(n3075), .B(n3073), .Z(n3029) );
  XNOR U230 ( .A(n3297), .B(n3295), .Z(n3251) );
  XNOR U231 ( .A(n3519), .B(n3517), .Z(n3473) );
  XNOR U232 ( .A(n3741), .B(n3739), .Z(n3695) );
  XNOR U233 ( .A(n3963), .B(n3961), .Z(n3917) );
  XNOR U234 ( .A(n4185), .B(n4183), .Z(n4139) );
  XNOR U235 ( .A(n4433), .B(n4431), .Z(n4409) );
  AND U236 ( .A(n325), .B(n324), .Z(n292) );
  XOR U237 ( .A(n4516), .B(n4534), .Z(n4521) );
  XOR U238 ( .A(n1589), .B(n1618), .Z(n1594) );
  XNOR U239 ( .A(n1702), .B(n1667), .Z(n1669) );
  XOR U240 ( .A(n1820), .B(n1842), .Z(n1827) );
  XNOR U241 ( .A(n1905), .B(n1904), .Z(n1888) );
  XOR U242 ( .A(n2042), .B(n2064), .Z(n2049) );
  XNOR U243 ( .A(n2127), .B(n2126), .Z(n2110) );
  XOR U244 ( .A(n2264), .B(n2286), .Z(n2271) );
  XNOR U245 ( .A(n2349), .B(n2348), .Z(n2332) );
  XOR U246 ( .A(n2486), .B(n2508), .Z(n2493) );
  XNOR U247 ( .A(n2571), .B(n2570), .Z(n2554) );
  XOR U248 ( .A(n2708), .B(n2730), .Z(n2715) );
  XNOR U249 ( .A(n2793), .B(n2792), .Z(n2776) );
  XOR U250 ( .A(n2930), .B(n2952), .Z(n2937) );
  XNOR U251 ( .A(n3015), .B(n3014), .Z(n2998) );
  XOR U252 ( .A(n3152), .B(n3174), .Z(n3159) );
  XNOR U253 ( .A(n3237), .B(n3236), .Z(n3220) );
  XOR U254 ( .A(n3374), .B(n3396), .Z(n3381) );
  XNOR U255 ( .A(n3459), .B(n3458), .Z(n3442) );
  XOR U256 ( .A(n3596), .B(n3618), .Z(n3603) );
  XNOR U257 ( .A(n3681), .B(n3680), .Z(n3664) );
  XOR U258 ( .A(n3818), .B(n3840), .Z(n3825) );
  XNOR U259 ( .A(n3903), .B(n3902), .Z(n3886) );
  XOR U260 ( .A(n4040), .B(n4062), .Z(n4047) );
  XNOR U261 ( .A(n4125), .B(n4124), .Z(n4108) );
  XOR U262 ( .A(n4262), .B(n4284), .Z(n4269) );
  XNOR U263 ( .A(n4347), .B(n4346), .Z(n4330) );
  XOR U264 ( .A(n249), .B(n268), .Z(n259) );
  XOR U265 ( .A(n313), .B(n333), .Z(n323) );
  XOR U266 ( .A(n378), .B(n398), .Z(n388) );
  XOR U267 ( .A(n451), .B(n472), .Z(n461) );
  XOR U268 ( .A(n519), .B(n540), .Z(n529) );
  XOR U269 ( .A(n587), .B(n608), .Z(n597) );
  XOR U270 ( .A(n655), .B(n676), .Z(n665) );
  XOR U271 ( .A(n723), .B(n744), .Z(n733) );
  XOR U272 ( .A(n793), .B(n814), .Z(n803) );
  XOR U273 ( .A(n869), .B(n889), .Z(n878) );
  XOR U274 ( .A(n945), .B(n965), .Z(n954) );
  XOR U275 ( .A(n1021), .B(n1041), .Z(n1030) );
  XOR U276 ( .A(n1097), .B(n1577), .Z(n1106) );
  XNOR U277 ( .A(n1736), .B(n1735), .Z(n1712) );
  XOR U278 ( .A(n1949), .B(n1959), .Z(n1916) );
  XOR U279 ( .A(n2171), .B(n2181), .Z(n2138) );
  XOR U280 ( .A(n2393), .B(n2403), .Z(n2360) );
  XOR U281 ( .A(n2615), .B(n2625), .Z(n2582) );
  XOR U282 ( .A(n2837), .B(n2847), .Z(n2804) );
  XOR U283 ( .A(n3059), .B(n3069), .Z(n3026) );
  XOR U284 ( .A(n3281), .B(n3291), .Z(n3248) );
  XOR U285 ( .A(n3503), .B(n3513), .Z(n3470) );
  XOR U286 ( .A(n3725), .B(n3735), .Z(n3692) );
  XOR U287 ( .A(n3947), .B(n3957), .Z(n3914) );
  XOR U288 ( .A(n4169), .B(n4179), .Z(n4136) );
  XNOR U289 ( .A(n1615), .B(n1613), .Z(n1603) );
  XNOR U290 ( .A(n1680), .B(n1678), .Z(n1650) );
  XNOR U291 ( .A(n1769), .B(n1767), .Z(n1745) );
  XNOR U292 ( .A(n1833), .B(n1831), .Z(n1803) );
  XNOR U293 ( .A(n1885), .B(n1883), .Z(n1855) );
  XNOR U294 ( .A(n1991), .B(n1989), .Z(n1967) );
  XNOR U295 ( .A(n2055), .B(n2053), .Z(n2025) );
  XNOR U296 ( .A(n2107), .B(n2105), .Z(n2077) );
  XNOR U297 ( .A(n2213), .B(n2211), .Z(n2189) );
  XNOR U298 ( .A(n2277), .B(n2275), .Z(n2247) );
  XNOR U299 ( .A(n2329), .B(n2327), .Z(n2299) );
  XNOR U300 ( .A(n2435), .B(n2433), .Z(n2411) );
  XNOR U301 ( .A(n2499), .B(n2497), .Z(n2469) );
  XNOR U302 ( .A(n2551), .B(n2549), .Z(n2521) );
  XNOR U303 ( .A(n2657), .B(n2655), .Z(n2633) );
  XNOR U304 ( .A(n2721), .B(n2719), .Z(n2691) );
  XNOR U305 ( .A(n2773), .B(n2771), .Z(n2743) );
  XNOR U306 ( .A(n2879), .B(n2877), .Z(n2855) );
  XNOR U307 ( .A(n2943), .B(n2941), .Z(n2913) );
  XNOR U308 ( .A(n2995), .B(n2993), .Z(n2965) );
  XNOR U309 ( .A(n3101), .B(n3099), .Z(n3077) );
  XNOR U310 ( .A(n3165), .B(n3163), .Z(n3135) );
  XNOR U311 ( .A(n3217), .B(n3215), .Z(n3187) );
  XNOR U312 ( .A(n3323), .B(n3321), .Z(n3299) );
  XNOR U313 ( .A(n3387), .B(n3385), .Z(n3357) );
  XNOR U314 ( .A(n3439), .B(n3437), .Z(n3409) );
  XNOR U315 ( .A(n3545), .B(n3543), .Z(n3521) );
  XNOR U316 ( .A(n3609), .B(n3607), .Z(n3579) );
  XNOR U317 ( .A(n3661), .B(n3659), .Z(n3631) );
  XNOR U318 ( .A(n3767), .B(n3765), .Z(n3743) );
  XNOR U319 ( .A(n3831), .B(n3829), .Z(n3801) );
  XNOR U320 ( .A(n3883), .B(n3881), .Z(n3853) );
  XNOR U321 ( .A(n3989), .B(n3987), .Z(n3965) );
  XNOR U322 ( .A(n4053), .B(n4051), .Z(n4023) );
  XNOR U323 ( .A(n4105), .B(n4103), .Z(n4075) );
  XNOR U324 ( .A(n4211), .B(n4209), .Z(n4187) );
  XNOR U325 ( .A(n4275), .B(n4273), .Z(n4245) );
  XNOR U326 ( .A(n4327), .B(n4325), .Z(n4297) );
  XNOR U327 ( .A(n4407), .B(n4405), .Z(n4361) );
  XNOR U328 ( .A(n4465), .B(n4463), .Z(n4436) );
  XNOR U329 ( .A(n4658), .B(n4659), .Z(n4653) );
  XNOR U330 ( .A(n4618), .B(n4617), .Z(n4606) );
  XNOR U331 ( .A(n4555), .B(n4554), .Z(n4532) );
  AND U332 ( .A(n358), .B(n357), .Z(n324) );
  XOR U333 ( .A(n4545), .B(n4572), .Z(n4550) );
  XNOR U334 ( .A(n1670), .B(n1635), .Z(n1637) );
  XNOR U335 ( .A(n1733), .B(n1699), .Z(n1700) );
  XNOR U336 ( .A(n1873), .B(n1872), .Z(n1856) );
  XNOR U337 ( .A(n1955), .B(n1936), .Z(n1920) );
  XNOR U338 ( .A(n2095), .B(n2094), .Z(n2078) );
  XNOR U339 ( .A(n2177), .B(n2158), .Z(n2142) );
  XNOR U340 ( .A(n2317), .B(n2316), .Z(n2300) );
  XNOR U341 ( .A(n2399), .B(n2380), .Z(n2364) );
  XNOR U342 ( .A(n2539), .B(n2538), .Z(n2522) );
  XNOR U343 ( .A(n2621), .B(n2602), .Z(n2586) );
  XNOR U344 ( .A(n2761), .B(n2760), .Z(n2744) );
  XNOR U345 ( .A(n2843), .B(n2824), .Z(n2808) );
  XNOR U346 ( .A(n2983), .B(n2982), .Z(n2966) );
  XNOR U347 ( .A(n3065), .B(n3046), .Z(n3030) );
  XNOR U348 ( .A(n3205), .B(n3204), .Z(n3188) );
  XNOR U349 ( .A(n3287), .B(n3268), .Z(n3252) );
  XNOR U350 ( .A(n3427), .B(n3426), .Z(n3410) );
  XNOR U351 ( .A(n3509), .B(n3490), .Z(n3474) );
  XNOR U352 ( .A(n3649), .B(n3648), .Z(n3632) );
  XNOR U353 ( .A(n3731), .B(n3712), .Z(n3696) );
  XNOR U354 ( .A(n3871), .B(n3870), .Z(n3854) );
  XNOR U355 ( .A(n3953), .B(n3934), .Z(n3918) );
  XNOR U356 ( .A(n4093), .B(n4092), .Z(n4076) );
  XNOR U357 ( .A(n4175), .B(n4156), .Z(n4140) );
  XNOR U358 ( .A(n4315), .B(n4314), .Z(n4298) );
  XNOR U359 ( .A(n4397), .B(n4378), .Z(n4362) );
  XOR U360 ( .A(n4422), .B(n4442), .Z(n4428) );
  XOR U361 ( .A(n4484), .B(n4501), .Z(n4491) );
  XOR U362 ( .A(n281), .B(n300), .Z(n291) );
  XOR U363 ( .A(n346), .B(n365), .Z(n356) );
  XOR U364 ( .A(n411), .B(n438), .Z(n421) );
  XOR U365 ( .A(n485), .B(n506), .Z(n495) );
  XOR U366 ( .A(n553), .B(n574), .Z(n563) );
  XOR U367 ( .A(n621), .B(n642), .Z(n631) );
  XOR U368 ( .A(n689), .B(n710), .Z(n699) );
  XOR U369 ( .A(n757), .B(n780), .Z(n767) );
  XOR U370 ( .A(n827), .B(n848), .Z(n837) );
  XOR U371 ( .A(n907), .B(n927), .Z(n916) );
  XOR U372 ( .A(n983), .B(n1003), .Z(n992) );
  XOR U373 ( .A(n1059), .B(n1079), .Z(n1068) );
  XNOR U374 ( .A(n1601), .B(n1599), .Z(n1576) );
  XNOR U375 ( .A(n1648), .B(n1646), .Z(n1617) );
  XNOR U376 ( .A(n1712), .B(n1710), .Z(n1682) );
  XNOR U377 ( .A(n1801), .B(n1799), .Z(n1772) );
  XNOR U378 ( .A(n1853), .B(n1851), .Z(n1835) );
  XNOR U379 ( .A(n1917), .B(n1915), .Z(n1887) );
  XNOR U380 ( .A(n2023), .B(n2021), .Z(n1994) );
  XNOR U381 ( .A(n2075), .B(n2073), .Z(n2057) );
  XNOR U382 ( .A(n2139), .B(n2137), .Z(n2109) );
  XNOR U383 ( .A(n2245), .B(n2243), .Z(n2216) );
  XNOR U384 ( .A(n2297), .B(n2295), .Z(n2279) );
  XNOR U385 ( .A(n2361), .B(n2359), .Z(n2331) );
  XNOR U386 ( .A(n2467), .B(n2465), .Z(n2438) );
  XNOR U387 ( .A(n2519), .B(n2517), .Z(n2501) );
  XNOR U388 ( .A(n2583), .B(n2581), .Z(n2553) );
  XNOR U389 ( .A(n2689), .B(n2687), .Z(n2660) );
  XNOR U390 ( .A(n2741), .B(n2739), .Z(n2723) );
  XNOR U391 ( .A(n2805), .B(n2803), .Z(n2775) );
  XNOR U392 ( .A(n2911), .B(n2909), .Z(n2882) );
  XNOR U393 ( .A(n2963), .B(n2961), .Z(n2945) );
  XNOR U394 ( .A(n3027), .B(n3025), .Z(n2997) );
  XNOR U395 ( .A(n3133), .B(n3131), .Z(n3104) );
  XNOR U396 ( .A(n3185), .B(n3183), .Z(n3167) );
  XNOR U397 ( .A(n3249), .B(n3247), .Z(n3219) );
  XNOR U398 ( .A(n3355), .B(n3353), .Z(n3326) );
  XNOR U399 ( .A(n3407), .B(n3405), .Z(n3389) );
  XNOR U400 ( .A(n3471), .B(n3469), .Z(n3441) );
  XNOR U401 ( .A(n3577), .B(n3575), .Z(n3548) );
  XNOR U402 ( .A(n3629), .B(n3627), .Z(n3611) );
  XNOR U403 ( .A(n3693), .B(n3691), .Z(n3663) );
  XNOR U404 ( .A(n3799), .B(n3797), .Z(n3770) );
  XNOR U405 ( .A(n3851), .B(n3849), .Z(n3833) );
  XNOR U406 ( .A(n3915), .B(n3913), .Z(n3885) );
  XNOR U407 ( .A(n4021), .B(n4019), .Z(n3992) );
  XNOR U408 ( .A(n4073), .B(n4071), .Z(n4055) );
  XNOR U409 ( .A(n4137), .B(n4135), .Z(n4107) );
  XNOR U410 ( .A(n4243), .B(n4241), .Z(n4214) );
  XNOR U411 ( .A(n4295), .B(n4293), .Z(n4277) );
  XNOR U412 ( .A(n4359), .B(n4357), .Z(n4329) );
  XNOR U413 ( .A(n4639), .B(n4638), .Z(n4633) );
  XNOR U414 ( .A(n4591), .B(n4590), .Z(n4570) );
  XNOR U415 ( .A(n4495), .B(n4494), .Z(n4467) );
  XNOR U416 ( .A(n1745), .B(n1744), .Z(n1140) );
  XNOR U417 ( .A(n1967), .B(n1966), .Z(n1175) );
  XNOR U418 ( .A(n2189), .B(n2188), .Z(n1210) );
  XNOR U419 ( .A(n2411), .B(n2410), .Z(n1245) );
  XNOR U420 ( .A(n2633), .B(n2632), .Z(n1280) );
  XNOR U421 ( .A(n2855), .B(n2854), .Z(n1315) );
  XNOR U422 ( .A(n3077), .B(n3076), .Z(n1350) );
  XNOR U423 ( .A(n3299), .B(n3298), .Z(n1385) );
  XNOR U424 ( .A(n3521), .B(n3520), .Z(n1420) );
  XNOR U425 ( .A(n3743), .B(n3742), .Z(n1455) );
  XNOR U426 ( .A(n3965), .B(n3964), .Z(n1490) );
  XNOR U427 ( .A(n4187), .B(n4186), .Z(n1525) );
  XNOR U428 ( .A(n4409), .B(n4408), .Z(n1560) );
  XOR U429 ( .A(n4653), .B(n4660), .Z(n4648) );
  AND U430 ( .A(n390), .B(n389), .Z(n357) );
  NAND U431 ( .A(n261), .B(n260), .Z(n222) );
  XNOR U432 ( .A(n1), .B(n2), .Z(swire[9]) );
  XNOR U433 ( .A(n3), .B(n4), .Z(swire[99]) );
  XNOR U434 ( .A(n5), .B(n6), .Z(swire[98]) );
  XNOR U435 ( .A(n7), .B(n8), .Z(swire[97]) );
  XNOR U436 ( .A(n9), .B(n10), .Z(swire[96]) );
  XNOR U437 ( .A(n11), .B(n12), .Z(swire[95]) );
  XNOR U438 ( .A(n13), .B(n14), .Z(swire[94]) );
  XNOR U439 ( .A(n15), .B(n16), .Z(swire[93]) );
  XNOR U440 ( .A(n17), .B(n18), .Z(swire[92]) );
  XNOR U441 ( .A(n19), .B(n20), .Z(swire[91]) );
  XNOR U442 ( .A(n21), .B(n22), .Z(swire[90]) );
  XNOR U443 ( .A(n23), .B(n24), .Z(swire[8]) );
  XNOR U444 ( .A(n25), .B(n26), .Z(swire[89]) );
  XNOR U445 ( .A(n27), .B(n28), .Z(swire[88]) );
  XNOR U446 ( .A(n29), .B(n30), .Z(swire[87]) );
  XNOR U447 ( .A(n31), .B(n32), .Z(swire[86]) );
  XNOR U448 ( .A(n33), .B(n34), .Z(swire[85]) );
  XNOR U449 ( .A(n35), .B(n36), .Z(swire[84]) );
  XNOR U450 ( .A(n37), .B(n38), .Z(swire[83]) );
  XNOR U451 ( .A(n39), .B(n40), .Z(swire[82]) );
  XNOR U452 ( .A(n41), .B(n42), .Z(swire[81]) );
  XNOR U453 ( .A(n43), .B(n44), .Z(swire[80]) );
  XNOR U454 ( .A(n45), .B(n46), .Z(swire[79]) );
  XNOR U455 ( .A(n47), .B(n48), .Z(swire[78]) );
  XNOR U456 ( .A(n49), .B(n50), .Z(swire[77]) );
  XNOR U457 ( .A(n51), .B(n52), .Z(swire[76]) );
  XNOR U458 ( .A(n53), .B(n54), .Z(swire[75]) );
  XNOR U459 ( .A(n55), .B(n56), .Z(swire[74]) );
  XNOR U460 ( .A(n57), .B(n58), .Z(swire[73]) );
  XNOR U461 ( .A(n59), .B(n60), .Z(swire[72]) );
  XNOR U462 ( .A(n61), .B(n62), .Z(swire[71]) );
  XNOR U463 ( .A(n63), .B(n64), .Z(swire[70]) );
  XNOR U464 ( .A(n65), .B(n66), .Z(swire[69]) );
  XNOR U465 ( .A(n67), .B(n68), .Z(swire[68]) );
  XNOR U466 ( .A(n69), .B(n70), .Z(swire[67]) );
  XNOR U467 ( .A(n71), .B(n72), .Z(swire[66]) );
  XNOR U468 ( .A(n73), .B(n74), .Z(swire[65]) );
  XNOR U469 ( .A(n75), .B(n76), .Z(swire[64]) );
  XNOR U470 ( .A(n77), .B(n78), .Z(swire[63]) );
  XNOR U471 ( .A(n79), .B(n80), .Z(swire[62]) );
  XNOR U472 ( .A(n81), .B(n82), .Z(swire[61]) );
  XNOR U473 ( .A(n83), .B(n84), .Z(swire[60]) );
  XNOR U474 ( .A(n85), .B(n86), .Z(swire[59]) );
  XNOR U475 ( .A(n87), .B(n88), .Z(swire[58]) );
  XNOR U476 ( .A(n89), .B(n90), .Z(swire[57]) );
  XNOR U477 ( .A(n91), .B(n92), .Z(swire[56]) );
  XNOR U478 ( .A(n93), .B(n94), .Z(swire[55]) );
  XNOR U479 ( .A(n95), .B(n96), .Z(swire[54]) );
  XNOR U480 ( .A(n97), .B(n98), .Z(swire[53]) );
  XNOR U481 ( .A(n99), .B(n100), .Z(swire[52]) );
  XNOR U482 ( .A(n101), .B(n102), .Z(swire[51]) );
  XNOR U483 ( .A(n103), .B(n104), .Z(swire[50]) );
  XNOR U484 ( .A(n105), .B(n106), .Z(swire[49]) );
  XNOR U485 ( .A(n107), .B(n108), .Z(swire[48]) );
  XNOR U486 ( .A(n109), .B(n110), .Z(swire[47]) );
  XNOR U487 ( .A(n111), .B(n112), .Z(swire[46]) );
  XNOR U488 ( .A(n113), .B(n114), .Z(swire[45]) );
  XNOR U489 ( .A(n115), .B(n116), .Z(swire[44]) );
  XNOR U490 ( .A(n117), .B(n118), .Z(swire[43]) );
  XNOR U491 ( .A(n119), .B(n120), .Z(swire[42]) );
  XNOR U492 ( .A(n121), .B(n122), .Z(swire[41]) );
  XNOR U493 ( .A(n123), .B(n124), .Z(swire[40]) );
  XNOR U494 ( .A(n125), .B(n126), .Z(swire[39]) );
  XNOR U495 ( .A(n127), .B(n128), .Z(swire[38]) );
  XNOR U496 ( .A(n129), .B(n130), .Z(swire[37]) );
  XNOR U497 ( .A(n131), .B(n132), .Z(swire[36]) );
  XNOR U498 ( .A(n133), .B(n134), .Z(swire[35]) );
  XNOR U499 ( .A(n135), .B(n136), .Z(swire[34]) );
  XNOR U500 ( .A(n137), .B(n138), .Z(swire[33]) );
  XNOR U501 ( .A(n139), .B(n140), .Z(swire[32]) );
  XNOR U502 ( .A(n141), .B(n142), .Z(swire[31]) );
  XNOR U503 ( .A(n143), .B(n144), .Z(swire[30]) );
  XNOR U504 ( .A(n145), .B(n146), .Z(swire[29]) );
  XNOR U505 ( .A(n147), .B(n148), .Z(swire[28]) );
  XNOR U506 ( .A(n149), .B(n150), .Z(swire[27]) );
  XNOR U507 ( .A(n151), .B(n152), .Z(swire[26]) );
  XNOR U508 ( .A(n153), .B(n154), .Z(swire[25]) );
  XNOR U509 ( .A(n155), .B(n156), .Z(swire[24]) );
  XNOR U510 ( .A(n157), .B(n158), .Z(swire[23]) );
  XNOR U511 ( .A(n159), .B(n160), .Z(swire[22]) );
  XNOR U512 ( .A(n161), .B(n162), .Z(swire[21]) );
  XNOR U513 ( .A(n163), .B(n164), .Z(swire[20]) );
  XNOR U514 ( .A(n165), .B(n166), .Z(swire[19]) );
  XNOR U515 ( .A(n167), .B(n168), .Z(swire[18]) );
  XNOR U516 ( .A(n169), .B(n170), .Z(swire[17]) );
  XNOR U517 ( .A(n171), .B(n172), .Z(swire[16]) );
  XNOR U518 ( .A(n173), .B(n174), .Z(swire[15]) );
  XNOR U519 ( .A(n175), .B(n176), .Z(swire[14]) );
  XNOR U520 ( .A(n177), .B(n178), .Z(swire[13]) );
  XNOR U521 ( .A(n179), .B(n180), .Z(swire[12]) );
  XOR U522 ( .A(n181), .B(n182), .Z(swire[127]) );
  XOR U523 ( .A(n183), .B(n184), .Z(n182) );
  XOR U524 ( .A(n185), .B(n186), .Z(n184) );
  ANDN U525 ( .B(a[127]), .A(n187), .Z(n186) );
  AND U526 ( .A(b[1]), .B(a[126]), .Z(n185) );
  XOR U527 ( .A(n188), .B(n189), .Z(n183) );
  AND U528 ( .A(b[2]), .B(a[125]), .Z(n189) );
  AND U529 ( .A(b[3]), .B(a[124]), .Z(n188) );
  XOR U530 ( .A(n190), .B(n191), .Z(n181) );
  XOR U531 ( .A(n192), .B(n193), .Z(n191) );
  AND U532 ( .A(b[4]), .B(a[123]), .Z(n193) );
  AND U533 ( .A(b[5]), .B(a[122]), .Z(n192) );
  XOR U534 ( .A(n194), .B(n195), .Z(n190) );
  AND U535 ( .A(b[6]), .B(a[121]), .Z(n195) );
  AND U536 ( .A(b[7]), .B(a[120]), .Z(n194) );
  XOR U537 ( .A(n196), .B(n197), .Z(swire[126]) );
  XOR U538 ( .A(n198), .B(n199), .Z(n197) );
  XNOR U539 ( .A(n200), .B(n201), .Z(n199) );
  ANDN U540 ( .B(a[126]), .A(n187), .Z(n200) );
  XOR U541 ( .A(n202), .B(n203), .Z(n198) );
  XNOR U542 ( .A(n201), .B(n204), .Z(n203) );
  XNOR U543 ( .A(n205), .B(n206), .Z(n204) );
  AND U544 ( .A(b[3]), .B(a[123]), .Z(n205) );
  XOR U545 ( .A(n207), .B(n208), .Z(n201) );
  OR U546 ( .A(n209), .B(n210), .Z(n208) );
  XOR U547 ( .A(n211), .B(n212), .Z(n202) );
  XOR U548 ( .A(n213), .B(n214), .Z(n212) );
  AND U549 ( .A(b[4]), .B(a[122]), .Z(n214) );
  AND U550 ( .A(b[5]), .B(a[121]), .Z(n213) );
  XOR U551 ( .A(n215), .B(n216), .Z(n211) );
  AND U552 ( .A(b[6]), .B(a[120]), .Z(n216) );
  AND U553 ( .A(b[7]), .B(a[119]), .Z(n215) );
  XOR U554 ( .A(n217), .B(n218), .Z(n196) );
  XNOR U555 ( .A(n219), .B(n206), .Z(n218) );
  NANDN U556 ( .A(n220), .B(n221), .Z(n206) );
  AND U557 ( .A(b[2]), .B(a[124]), .Z(n219) );
  AND U558 ( .A(b[1]), .B(a[125]), .Z(n217) );
  XNOR U559 ( .A(n222), .B(n223), .Z(swire[125]) );
  XOR U560 ( .A(n221), .B(n224), .Z(n223) );
  XOR U561 ( .A(n220), .B(n222), .Z(n224) );
  NANDN U562 ( .A(n187), .B(a[125]), .Z(n220) );
  XOR U563 ( .A(n209), .B(n210), .Z(n221) );
  XOR U564 ( .A(n207), .B(n225), .Z(n210) );
  NAND U565 ( .A(b[1]), .B(a[124]), .Z(n225) );
  XOR U566 ( .A(n226), .B(n227), .Z(n209) );
  XOR U567 ( .A(n207), .B(n228), .Z(n227) );
  XOR U568 ( .A(n229), .B(n230), .Z(n228) );
  AND U569 ( .A(b[2]), .B(a[123]), .Z(n229) );
  ANDN U570 ( .B(n231), .A(n232), .Z(n207) );
  XOR U571 ( .A(n233), .B(n234), .Z(n226) );
  XNOR U572 ( .A(n230), .B(n235), .Z(n234) );
  XOR U573 ( .A(n236), .B(n237), .Z(n235) );
  XOR U574 ( .A(n238), .B(n239), .Z(n237) );
  XOR U575 ( .A(n240), .B(n241), .Z(n239) );
  XOR U576 ( .A(n242), .B(n243), .Z(n241) );
  AND U577 ( .A(b[5]), .B(a[120]), .Z(n242) );
  XOR U578 ( .A(n244), .B(n245), .Z(n240) );
  AND U579 ( .A(b[6]), .B(a[119]), .Z(n245) );
  AND U580 ( .A(b[7]), .B(a[118]), .Z(n244) );
  XOR U581 ( .A(n246), .B(n243), .Z(n236) );
  XOR U582 ( .A(n247), .B(n248), .Z(n243) );
  NOR U583 ( .A(n249), .B(n250), .Z(n247) );
  AND U584 ( .A(b[4]), .B(a[121]), .Z(n246) );
  XNOR U585 ( .A(n251), .B(n252), .Z(n230) );
  NANDN U586 ( .A(n253), .B(n254), .Z(n252) );
  XOR U587 ( .A(n255), .B(n238), .Z(n233) );
  XNOR U588 ( .A(n256), .B(n257), .Z(n238) );
  AND U589 ( .A(n258), .B(n259), .Z(n256) );
  AND U590 ( .A(b[3]), .B(a[122]), .Z(n255) );
  XNOR U591 ( .A(n260), .B(n261), .Z(swire[124]) );
  XOR U592 ( .A(n231), .B(n262), .Z(n261) );
  XOR U593 ( .A(n232), .B(n260), .Z(n262) );
  NANDN U594 ( .A(n187), .B(a[124]), .Z(n232) );
  XNOR U595 ( .A(n253), .B(n254), .Z(n231) );
  XOR U596 ( .A(n251), .B(n263), .Z(n254) );
  NAND U597 ( .A(b[1]), .B(a[123]), .Z(n263) );
  XOR U598 ( .A(n259), .B(n264), .Z(n253) );
  XOR U599 ( .A(n251), .B(n258), .Z(n264) );
  XNOR U600 ( .A(n265), .B(n257), .Z(n258) );
  AND U601 ( .A(b[2]), .B(a[122]), .Z(n265) );
  NANDN U602 ( .A(n266), .B(n267), .Z(n251) );
  XNOR U603 ( .A(n257), .B(n250), .Z(n268) );
  XOR U604 ( .A(n269), .B(n270), .Z(n250) );
  XOR U605 ( .A(n248), .B(n271), .Z(n270) );
  XOR U606 ( .A(n272), .B(n273), .Z(n271) );
  XNOR U607 ( .A(n274), .B(n275), .Z(n273) );
  AND U608 ( .A(b[5]), .B(a[119]), .Z(n274) );
  XOR U609 ( .A(n276), .B(n277), .Z(n272) );
  AND U610 ( .A(b[6]), .B(a[118]), .Z(n277) );
  AND U611 ( .A(b[7]), .B(a[117]), .Z(n276) );
  XOR U612 ( .A(n278), .B(n275), .Z(n269) );
  XOR U613 ( .A(n279), .B(n280), .Z(n275) );
  NOR U614 ( .A(n281), .B(n282), .Z(n279) );
  AND U615 ( .A(b[4]), .B(a[120]), .Z(n278) );
  XNOR U616 ( .A(n283), .B(n284), .Z(n257) );
  NANDN U617 ( .A(n285), .B(n286), .Z(n284) );
  XNOR U618 ( .A(n287), .B(n248), .Z(n249) );
  XNOR U619 ( .A(n288), .B(n289), .Z(n248) );
  AND U620 ( .A(n290), .B(n291), .Z(n288) );
  AND U621 ( .A(b[3]), .B(a[121]), .Z(n287) );
  XNOR U622 ( .A(n292), .B(n293), .Z(swire[123]) );
  XOR U623 ( .A(n267), .B(n294), .Z(n293) );
  XOR U624 ( .A(n266), .B(n292), .Z(n294) );
  NANDN U625 ( .A(n187), .B(a[123]), .Z(n266) );
  XNOR U626 ( .A(n285), .B(n286), .Z(n267) );
  XOR U627 ( .A(n283), .B(n295), .Z(n286) );
  NAND U628 ( .A(b[1]), .B(a[122]), .Z(n295) );
  XOR U629 ( .A(n291), .B(n296), .Z(n285) );
  XOR U630 ( .A(n283), .B(n290), .Z(n296) );
  XNOR U631 ( .A(n297), .B(n289), .Z(n290) );
  AND U632 ( .A(b[2]), .B(a[121]), .Z(n297) );
  NANDN U633 ( .A(n298), .B(n299), .Z(n283) );
  XNOR U634 ( .A(n289), .B(n282), .Z(n300) );
  XOR U635 ( .A(n301), .B(n302), .Z(n282) );
  XOR U636 ( .A(n280), .B(n303), .Z(n302) );
  XOR U637 ( .A(n304), .B(n305), .Z(n303) );
  XNOR U638 ( .A(n306), .B(n307), .Z(n305) );
  AND U639 ( .A(b[5]), .B(a[118]), .Z(n306) );
  XOR U640 ( .A(n308), .B(n309), .Z(n304) );
  AND U641 ( .A(b[6]), .B(a[117]), .Z(n309) );
  AND U642 ( .A(b[7]), .B(a[116]), .Z(n308) );
  XOR U643 ( .A(n310), .B(n307), .Z(n301) );
  XOR U644 ( .A(n311), .B(n312), .Z(n307) );
  NOR U645 ( .A(n313), .B(n314), .Z(n311) );
  AND U646 ( .A(b[4]), .B(a[119]), .Z(n310) );
  XNOR U647 ( .A(n315), .B(n316), .Z(n289) );
  NANDN U648 ( .A(n317), .B(n318), .Z(n316) );
  XNOR U649 ( .A(n319), .B(n280), .Z(n281) );
  XNOR U650 ( .A(n320), .B(n321), .Z(n280) );
  AND U651 ( .A(n322), .B(n323), .Z(n320) );
  AND U652 ( .A(b[3]), .B(a[120]), .Z(n319) );
  XNOR U653 ( .A(n324), .B(n325), .Z(swire[122]) );
  XOR U654 ( .A(n299), .B(n327), .Z(n325) );
  XNOR U655 ( .A(n298), .B(n326), .Z(n327) );
  IV U656 ( .A(n324), .Z(n326) );
  NANDN U657 ( .A(n187), .B(a[122]), .Z(n298) );
  XNOR U658 ( .A(n317), .B(n318), .Z(n299) );
  XOR U659 ( .A(n315), .B(n328), .Z(n318) );
  NAND U660 ( .A(b[1]), .B(a[121]), .Z(n328) );
  XOR U661 ( .A(n323), .B(n329), .Z(n317) );
  XOR U662 ( .A(n315), .B(n322), .Z(n329) );
  XNOR U663 ( .A(n330), .B(n321), .Z(n322) );
  AND U664 ( .A(b[2]), .B(a[120]), .Z(n330) );
  NANDN U665 ( .A(n331), .B(n332), .Z(n315) );
  XNOR U666 ( .A(n321), .B(n314), .Z(n333) );
  XOR U667 ( .A(n334), .B(n335), .Z(n314) );
  XOR U668 ( .A(n312), .B(n336), .Z(n335) );
  XOR U669 ( .A(n337), .B(n338), .Z(n336) );
  XNOR U670 ( .A(n339), .B(n340), .Z(n338) );
  AND U671 ( .A(b[5]), .B(a[117]), .Z(n339) );
  XOR U672 ( .A(n341), .B(n342), .Z(n337) );
  AND U673 ( .A(b[6]), .B(a[116]), .Z(n342) );
  AND U674 ( .A(b[7]), .B(a[115]), .Z(n341) );
  XOR U675 ( .A(n343), .B(n340), .Z(n334) );
  XOR U676 ( .A(n344), .B(n345), .Z(n340) );
  NOR U677 ( .A(n346), .B(n347), .Z(n344) );
  AND U678 ( .A(b[4]), .B(a[118]), .Z(n343) );
  XNOR U679 ( .A(n348), .B(n349), .Z(n321) );
  NANDN U680 ( .A(n350), .B(n351), .Z(n349) );
  XNOR U681 ( .A(n352), .B(n312), .Z(n313) );
  XNOR U682 ( .A(n353), .B(n354), .Z(n312) );
  AND U683 ( .A(n355), .B(n356), .Z(n353) );
  AND U684 ( .A(b[3]), .B(a[119]), .Z(n352) );
  XNOR U685 ( .A(n357), .B(n358), .Z(swire[121]) );
  XOR U686 ( .A(n332), .B(n359), .Z(n358) );
  XOR U687 ( .A(n331), .B(n357), .Z(n359) );
  NANDN U688 ( .A(n187), .B(a[121]), .Z(n331) );
  XNOR U689 ( .A(n350), .B(n351), .Z(n332) );
  XOR U690 ( .A(n348), .B(n360), .Z(n351) );
  NAND U691 ( .A(b[1]), .B(a[120]), .Z(n360) );
  XOR U692 ( .A(n356), .B(n361), .Z(n350) );
  XOR U693 ( .A(n348), .B(n355), .Z(n361) );
  XNOR U694 ( .A(n362), .B(n354), .Z(n355) );
  AND U695 ( .A(b[2]), .B(a[119]), .Z(n362) );
  NANDN U696 ( .A(n363), .B(n364), .Z(n348) );
  XNOR U697 ( .A(n354), .B(n347), .Z(n365) );
  XOR U698 ( .A(n366), .B(n367), .Z(n347) );
  XOR U699 ( .A(n345), .B(n368), .Z(n367) );
  XOR U700 ( .A(n369), .B(n370), .Z(n368) );
  XNOR U701 ( .A(n371), .B(n372), .Z(n370) );
  AND U702 ( .A(b[5]), .B(a[116]), .Z(n371) );
  XOR U703 ( .A(n373), .B(n374), .Z(n369) );
  AND U704 ( .A(b[6]), .B(a[115]), .Z(n374) );
  AND U705 ( .A(b[7]), .B(a[114]), .Z(n373) );
  XOR U706 ( .A(n375), .B(n372), .Z(n366) );
  XOR U707 ( .A(n376), .B(n377), .Z(n372) );
  NOR U708 ( .A(n378), .B(n379), .Z(n376) );
  AND U709 ( .A(b[4]), .B(a[117]), .Z(n375) );
  XNOR U710 ( .A(n380), .B(n381), .Z(n354) );
  NANDN U711 ( .A(n382), .B(n383), .Z(n381) );
  XNOR U712 ( .A(n384), .B(n345), .Z(n346) );
  XNOR U713 ( .A(n385), .B(n386), .Z(n345) );
  AND U714 ( .A(n387), .B(n388), .Z(n385) );
  AND U715 ( .A(b[3]), .B(a[118]), .Z(n384) );
  XNOR U716 ( .A(n389), .B(n390), .Z(swire[120]) );
  XOR U717 ( .A(n364), .B(n392), .Z(n390) );
  XNOR U718 ( .A(n363), .B(n391), .Z(n392) );
  IV U719 ( .A(n389), .Z(n391) );
  NANDN U720 ( .A(n187), .B(a[120]), .Z(n363) );
  XNOR U721 ( .A(n382), .B(n383), .Z(n364) );
  XOR U722 ( .A(n380), .B(n393), .Z(n383) );
  NAND U723 ( .A(b[1]), .B(a[119]), .Z(n393) );
  XOR U724 ( .A(n388), .B(n394), .Z(n382) );
  XOR U725 ( .A(n380), .B(n387), .Z(n394) );
  XNOR U726 ( .A(n395), .B(n386), .Z(n387) );
  AND U727 ( .A(b[2]), .B(a[118]), .Z(n395) );
  NANDN U728 ( .A(n396), .B(n397), .Z(n380) );
  XNOR U729 ( .A(n386), .B(n379), .Z(n398) );
  XOR U730 ( .A(n399), .B(n400), .Z(n379) );
  XOR U731 ( .A(n377), .B(n401), .Z(n400) );
  XOR U732 ( .A(n402), .B(n403), .Z(n401) );
  XNOR U733 ( .A(n404), .B(n405), .Z(n403) );
  AND U734 ( .A(b[5]), .B(a[115]), .Z(n404) );
  XOR U735 ( .A(n406), .B(n407), .Z(n402) );
  AND U736 ( .A(b[6]), .B(a[114]), .Z(n407) );
  AND U737 ( .A(b[7]), .B(a[113]), .Z(n406) );
  XOR U738 ( .A(n408), .B(n405), .Z(n399) );
  XOR U739 ( .A(n409), .B(n410), .Z(n405) );
  NOR U740 ( .A(n411), .B(n412), .Z(n409) );
  AND U741 ( .A(b[4]), .B(a[116]), .Z(n408) );
  XNOR U742 ( .A(n413), .B(n414), .Z(n386) );
  NANDN U743 ( .A(n415), .B(n416), .Z(n414) );
  XNOR U744 ( .A(n417), .B(n377), .Z(n378) );
  XNOR U745 ( .A(n418), .B(n419), .Z(n377) );
  AND U746 ( .A(n420), .B(n421), .Z(n418) );
  AND U747 ( .A(b[3]), .B(a[117]), .Z(n417) );
  XNOR U748 ( .A(n422), .B(n423), .Z(n389) );
  NOR U749 ( .A(n424), .B(n425), .Z(n422) );
  XNOR U750 ( .A(n426), .B(n427), .Z(swire[11]) );
  XOR U751 ( .A(n425), .B(n424), .Z(swire[119]) );
  XOR U752 ( .A(sreg[247]), .B(n423), .Z(n424) );
  XOR U753 ( .A(n397), .B(n428), .Z(n425) );
  XNOR U754 ( .A(n396), .B(n423), .Z(n428) );
  XOR U755 ( .A(n429), .B(n430), .Z(n423) );
  NOR U756 ( .A(n431), .B(n432), .Z(n429) );
  NANDN U757 ( .A(n187), .B(a[119]), .Z(n396) );
  XNOR U758 ( .A(n415), .B(n416), .Z(n397) );
  XOR U759 ( .A(n413), .B(n433), .Z(n416) );
  NAND U760 ( .A(b[1]), .B(a[118]), .Z(n433) );
  XOR U761 ( .A(n421), .B(n434), .Z(n415) );
  XOR U762 ( .A(n413), .B(n420), .Z(n434) );
  XNOR U763 ( .A(n435), .B(n419), .Z(n420) );
  AND U764 ( .A(b[2]), .B(a[117]), .Z(n435) );
  NANDN U765 ( .A(n436), .B(n437), .Z(n413) );
  XNOR U766 ( .A(n419), .B(n412), .Z(n438) );
  XOR U767 ( .A(n439), .B(n440), .Z(n412) );
  XOR U768 ( .A(n410), .B(n441), .Z(n440) );
  XOR U769 ( .A(n442), .B(n443), .Z(n441) );
  XNOR U770 ( .A(n444), .B(n445), .Z(n443) );
  AND U771 ( .A(b[5]), .B(a[114]), .Z(n444) );
  XOR U772 ( .A(n446), .B(n447), .Z(n442) );
  AND U773 ( .A(b[6]), .B(a[113]), .Z(n447) );
  AND U774 ( .A(b[7]), .B(a[112]), .Z(n446) );
  XOR U775 ( .A(n448), .B(n445), .Z(n439) );
  XOR U776 ( .A(n449), .B(n450), .Z(n445) );
  NOR U777 ( .A(n451), .B(n452), .Z(n449) );
  AND U778 ( .A(b[4]), .B(a[115]), .Z(n448) );
  XNOR U779 ( .A(n453), .B(n454), .Z(n419) );
  NANDN U780 ( .A(n455), .B(n456), .Z(n454) );
  XNOR U781 ( .A(n457), .B(n410), .Z(n411) );
  XNOR U782 ( .A(n458), .B(n459), .Z(n410) );
  AND U783 ( .A(n460), .B(n461), .Z(n458) );
  AND U784 ( .A(b[3]), .B(a[116]), .Z(n457) );
  XOR U785 ( .A(n432), .B(n431), .Z(swire[118]) );
  XOR U786 ( .A(sreg[246]), .B(n430), .Z(n431) );
  XOR U787 ( .A(n437), .B(n462), .Z(n432) );
  XNOR U788 ( .A(n436), .B(n430), .Z(n462) );
  XOR U789 ( .A(n463), .B(n464), .Z(n430) );
  NOR U790 ( .A(n465), .B(n466), .Z(n463) );
  NANDN U791 ( .A(n187), .B(a[118]), .Z(n436) );
  XNOR U792 ( .A(n455), .B(n456), .Z(n437) );
  XOR U793 ( .A(n453), .B(n467), .Z(n456) );
  NAND U794 ( .A(b[1]), .B(a[117]), .Z(n467) );
  XOR U795 ( .A(n461), .B(n468), .Z(n455) );
  XOR U796 ( .A(n453), .B(n460), .Z(n468) );
  XNOR U797 ( .A(n469), .B(n459), .Z(n460) );
  AND U798 ( .A(b[2]), .B(a[116]), .Z(n469) );
  NANDN U799 ( .A(n470), .B(n471), .Z(n453) );
  XNOR U800 ( .A(n459), .B(n452), .Z(n472) );
  XOR U801 ( .A(n473), .B(n474), .Z(n452) );
  XOR U802 ( .A(n450), .B(n475), .Z(n474) );
  XOR U803 ( .A(n476), .B(n477), .Z(n475) );
  XNOR U804 ( .A(n478), .B(n479), .Z(n477) );
  AND U805 ( .A(b[5]), .B(a[113]), .Z(n478) );
  XOR U806 ( .A(n480), .B(n481), .Z(n476) );
  AND U807 ( .A(b[6]), .B(a[112]), .Z(n481) );
  AND U808 ( .A(b[7]), .B(a[111]), .Z(n480) );
  XOR U809 ( .A(n482), .B(n479), .Z(n473) );
  XOR U810 ( .A(n483), .B(n484), .Z(n479) );
  NOR U811 ( .A(n485), .B(n486), .Z(n483) );
  AND U812 ( .A(b[4]), .B(a[114]), .Z(n482) );
  XNOR U813 ( .A(n487), .B(n488), .Z(n459) );
  NANDN U814 ( .A(n489), .B(n490), .Z(n488) );
  XNOR U815 ( .A(n491), .B(n450), .Z(n451) );
  XNOR U816 ( .A(n492), .B(n493), .Z(n450) );
  AND U817 ( .A(n494), .B(n495), .Z(n492) );
  AND U818 ( .A(b[3]), .B(a[115]), .Z(n491) );
  XOR U819 ( .A(n466), .B(n465), .Z(swire[117]) );
  XOR U820 ( .A(sreg[245]), .B(n464), .Z(n465) );
  XOR U821 ( .A(n471), .B(n496), .Z(n466) );
  XNOR U822 ( .A(n470), .B(n464), .Z(n496) );
  XOR U823 ( .A(n497), .B(n498), .Z(n464) );
  NOR U824 ( .A(n499), .B(n500), .Z(n497) );
  NANDN U825 ( .A(n187), .B(a[117]), .Z(n470) );
  XNOR U826 ( .A(n489), .B(n490), .Z(n471) );
  XOR U827 ( .A(n487), .B(n501), .Z(n490) );
  NAND U828 ( .A(b[1]), .B(a[116]), .Z(n501) );
  XOR U829 ( .A(n495), .B(n502), .Z(n489) );
  XOR U830 ( .A(n487), .B(n494), .Z(n502) );
  XNOR U831 ( .A(n503), .B(n493), .Z(n494) );
  AND U832 ( .A(b[2]), .B(a[115]), .Z(n503) );
  NANDN U833 ( .A(n504), .B(n505), .Z(n487) );
  XNOR U834 ( .A(n493), .B(n486), .Z(n506) );
  XOR U835 ( .A(n507), .B(n508), .Z(n486) );
  XOR U836 ( .A(n484), .B(n509), .Z(n508) );
  XOR U837 ( .A(n510), .B(n511), .Z(n509) );
  XNOR U838 ( .A(n512), .B(n513), .Z(n511) );
  AND U839 ( .A(b[5]), .B(a[112]), .Z(n512) );
  XOR U840 ( .A(n514), .B(n515), .Z(n510) );
  AND U841 ( .A(b[6]), .B(a[111]), .Z(n515) );
  AND U842 ( .A(b[7]), .B(a[110]), .Z(n514) );
  XOR U843 ( .A(n516), .B(n513), .Z(n507) );
  XOR U844 ( .A(n517), .B(n518), .Z(n513) );
  NOR U845 ( .A(n519), .B(n520), .Z(n517) );
  AND U846 ( .A(b[4]), .B(a[113]), .Z(n516) );
  XNOR U847 ( .A(n521), .B(n522), .Z(n493) );
  NANDN U848 ( .A(n523), .B(n524), .Z(n522) );
  XNOR U849 ( .A(n525), .B(n484), .Z(n485) );
  XNOR U850 ( .A(n526), .B(n527), .Z(n484) );
  AND U851 ( .A(n528), .B(n529), .Z(n526) );
  AND U852 ( .A(b[3]), .B(a[114]), .Z(n525) );
  XOR U853 ( .A(n500), .B(n499), .Z(swire[116]) );
  XOR U854 ( .A(sreg[244]), .B(n498), .Z(n499) );
  XOR U855 ( .A(n505), .B(n530), .Z(n500) );
  XNOR U856 ( .A(n504), .B(n498), .Z(n530) );
  XOR U857 ( .A(n531), .B(n532), .Z(n498) );
  NOR U858 ( .A(n533), .B(n534), .Z(n531) );
  NANDN U859 ( .A(n187), .B(a[116]), .Z(n504) );
  XNOR U860 ( .A(n523), .B(n524), .Z(n505) );
  XOR U861 ( .A(n521), .B(n535), .Z(n524) );
  NAND U862 ( .A(b[1]), .B(a[115]), .Z(n535) );
  XOR U863 ( .A(n529), .B(n536), .Z(n523) );
  XOR U864 ( .A(n521), .B(n528), .Z(n536) );
  XNOR U865 ( .A(n537), .B(n527), .Z(n528) );
  AND U866 ( .A(b[2]), .B(a[114]), .Z(n537) );
  NANDN U867 ( .A(n538), .B(n539), .Z(n521) );
  XNOR U868 ( .A(n527), .B(n520), .Z(n540) );
  XOR U869 ( .A(n541), .B(n542), .Z(n520) );
  XOR U870 ( .A(n518), .B(n543), .Z(n542) );
  XOR U871 ( .A(n544), .B(n545), .Z(n543) );
  XNOR U872 ( .A(n546), .B(n547), .Z(n545) );
  AND U873 ( .A(b[5]), .B(a[111]), .Z(n546) );
  XOR U874 ( .A(n548), .B(n549), .Z(n544) );
  AND U875 ( .A(b[6]), .B(a[110]), .Z(n549) );
  AND U876 ( .A(b[7]), .B(a[109]), .Z(n548) );
  XOR U877 ( .A(n550), .B(n547), .Z(n541) );
  XOR U878 ( .A(n551), .B(n552), .Z(n547) );
  NOR U879 ( .A(n553), .B(n554), .Z(n551) );
  AND U880 ( .A(b[4]), .B(a[112]), .Z(n550) );
  XNOR U881 ( .A(n555), .B(n556), .Z(n527) );
  NANDN U882 ( .A(n557), .B(n558), .Z(n556) );
  XNOR U883 ( .A(n559), .B(n518), .Z(n519) );
  XNOR U884 ( .A(n560), .B(n561), .Z(n518) );
  AND U885 ( .A(n562), .B(n563), .Z(n560) );
  AND U886 ( .A(b[3]), .B(a[113]), .Z(n559) );
  XOR U887 ( .A(n534), .B(n533), .Z(swire[115]) );
  XOR U888 ( .A(sreg[243]), .B(n532), .Z(n533) );
  XOR U889 ( .A(n539), .B(n564), .Z(n534) );
  XNOR U890 ( .A(n538), .B(n532), .Z(n564) );
  XOR U891 ( .A(n565), .B(n566), .Z(n532) );
  NOR U892 ( .A(n567), .B(n568), .Z(n565) );
  NANDN U893 ( .A(n187), .B(a[115]), .Z(n538) );
  XNOR U894 ( .A(n557), .B(n558), .Z(n539) );
  XOR U895 ( .A(n555), .B(n569), .Z(n558) );
  NAND U896 ( .A(b[1]), .B(a[114]), .Z(n569) );
  XOR U897 ( .A(n563), .B(n570), .Z(n557) );
  XOR U898 ( .A(n555), .B(n562), .Z(n570) );
  XNOR U899 ( .A(n571), .B(n561), .Z(n562) );
  AND U900 ( .A(b[2]), .B(a[113]), .Z(n571) );
  NANDN U901 ( .A(n572), .B(n573), .Z(n555) );
  XNOR U902 ( .A(n561), .B(n554), .Z(n574) );
  XOR U903 ( .A(n575), .B(n576), .Z(n554) );
  XOR U904 ( .A(n552), .B(n577), .Z(n576) );
  XOR U905 ( .A(n578), .B(n579), .Z(n577) );
  XNOR U906 ( .A(n580), .B(n581), .Z(n579) );
  AND U907 ( .A(b[5]), .B(a[110]), .Z(n580) );
  XOR U908 ( .A(n582), .B(n583), .Z(n578) );
  AND U909 ( .A(b[6]), .B(a[109]), .Z(n583) );
  AND U910 ( .A(b[7]), .B(a[108]), .Z(n582) );
  XOR U911 ( .A(n584), .B(n581), .Z(n575) );
  XOR U912 ( .A(n585), .B(n586), .Z(n581) );
  NOR U913 ( .A(n587), .B(n588), .Z(n585) );
  AND U914 ( .A(b[4]), .B(a[111]), .Z(n584) );
  XNOR U915 ( .A(n589), .B(n590), .Z(n561) );
  NANDN U916 ( .A(n591), .B(n592), .Z(n590) );
  XNOR U917 ( .A(n593), .B(n552), .Z(n553) );
  XNOR U918 ( .A(n594), .B(n595), .Z(n552) );
  AND U919 ( .A(n596), .B(n597), .Z(n594) );
  AND U920 ( .A(b[3]), .B(a[112]), .Z(n593) );
  XOR U921 ( .A(n568), .B(n567), .Z(swire[114]) );
  XOR U922 ( .A(sreg[242]), .B(n566), .Z(n567) );
  XOR U923 ( .A(n573), .B(n598), .Z(n568) );
  XNOR U924 ( .A(n572), .B(n566), .Z(n598) );
  XOR U925 ( .A(n599), .B(n600), .Z(n566) );
  NOR U926 ( .A(n601), .B(n602), .Z(n599) );
  NANDN U927 ( .A(n187), .B(a[114]), .Z(n572) );
  XNOR U928 ( .A(n591), .B(n592), .Z(n573) );
  XOR U929 ( .A(n589), .B(n603), .Z(n592) );
  NAND U930 ( .A(b[1]), .B(a[113]), .Z(n603) );
  XOR U931 ( .A(n597), .B(n604), .Z(n591) );
  XOR U932 ( .A(n589), .B(n596), .Z(n604) );
  XNOR U933 ( .A(n605), .B(n595), .Z(n596) );
  AND U934 ( .A(b[2]), .B(a[112]), .Z(n605) );
  NANDN U935 ( .A(n606), .B(n607), .Z(n589) );
  XNOR U936 ( .A(n595), .B(n588), .Z(n608) );
  XOR U937 ( .A(n609), .B(n610), .Z(n588) );
  XOR U938 ( .A(n586), .B(n611), .Z(n610) );
  XOR U939 ( .A(n612), .B(n613), .Z(n611) );
  XNOR U940 ( .A(n614), .B(n615), .Z(n613) );
  AND U941 ( .A(b[5]), .B(a[109]), .Z(n614) );
  XOR U942 ( .A(n616), .B(n617), .Z(n612) );
  AND U943 ( .A(b[6]), .B(a[108]), .Z(n617) );
  AND U944 ( .A(b[7]), .B(a[107]), .Z(n616) );
  XOR U945 ( .A(n618), .B(n615), .Z(n609) );
  XOR U946 ( .A(n619), .B(n620), .Z(n615) );
  NOR U947 ( .A(n621), .B(n622), .Z(n619) );
  AND U948 ( .A(b[4]), .B(a[110]), .Z(n618) );
  XNOR U949 ( .A(n623), .B(n624), .Z(n595) );
  NANDN U950 ( .A(n625), .B(n626), .Z(n624) );
  XNOR U951 ( .A(n627), .B(n586), .Z(n587) );
  XNOR U952 ( .A(n628), .B(n629), .Z(n586) );
  AND U953 ( .A(n630), .B(n631), .Z(n628) );
  AND U954 ( .A(b[3]), .B(a[111]), .Z(n627) );
  XOR U955 ( .A(n602), .B(n601), .Z(swire[113]) );
  XOR U956 ( .A(sreg[241]), .B(n600), .Z(n601) );
  XOR U957 ( .A(n607), .B(n632), .Z(n602) );
  XNOR U958 ( .A(n606), .B(n600), .Z(n632) );
  XOR U959 ( .A(n633), .B(n634), .Z(n600) );
  NOR U960 ( .A(n635), .B(n636), .Z(n633) );
  NANDN U961 ( .A(n187), .B(a[113]), .Z(n606) );
  XNOR U962 ( .A(n625), .B(n626), .Z(n607) );
  XOR U963 ( .A(n623), .B(n637), .Z(n626) );
  NAND U964 ( .A(b[1]), .B(a[112]), .Z(n637) );
  XOR U965 ( .A(n631), .B(n638), .Z(n625) );
  XOR U966 ( .A(n623), .B(n630), .Z(n638) );
  XNOR U967 ( .A(n639), .B(n629), .Z(n630) );
  AND U968 ( .A(b[2]), .B(a[111]), .Z(n639) );
  NANDN U969 ( .A(n640), .B(n641), .Z(n623) );
  XNOR U970 ( .A(n629), .B(n622), .Z(n642) );
  XOR U971 ( .A(n643), .B(n644), .Z(n622) );
  XOR U972 ( .A(n620), .B(n645), .Z(n644) );
  XOR U973 ( .A(n646), .B(n647), .Z(n645) );
  XNOR U974 ( .A(n648), .B(n649), .Z(n647) );
  AND U975 ( .A(b[5]), .B(a[108]), .Z(n648) );
  XOR U976 ( .A(n650), .B(n651), .Z(n646) );
  AND U977 ( .A(b[6]), .B(a[107]), .Z(n651) );
  AND U978 ( .A(b[7]), .B(a[106]), .Z(n650) );
  XOR U979 ( .A(n652), .B(n649), .Z(n643) );
  XOR U980 ( .A(n653), .B(n654), .Z(n649) );
  NOR U981 ( .A(n655), .B(n656), .Z(n653) );
  AND U982 ( .A(b[4]), .B(a[109]), .Z(n652) );
  XNOR U983 ( .A(n657), .B(n658), .Z(n629) );
  NANDN U984 ( .A(n659), .B(n660), .Z(n658) );
  XNOR U985 ( .A(n661), .B(n620), .Z(n621) );
  XNOR U986 ( .A(n662), .B(n663), .Z(n620) );
  AND U987 ( .A(n664), .B(n665), .Z(n662) );
  AND U988 ( .A(b[3]), .B(a[110]), .Z(n661) );
  XOR U989 ( .A(n636), .B(n635), .Z(swire[112]) );
  XOR U990 ( .A(sreg[240]), .B(n634), .Z(n635) );
  XOR U991 ( .A(n641), .B(n666), .Z(n636) );
  XNOR U992 ( .A(n640), .B(n634), .Z(n666) );
  XOR U993 ( .A(n667), .B(n668), .Z(n634) );
  NOR U994 ( .A(n669), .B(n670), .Z(n667) );
  NANDN U995 ( .A(n187), .B(a[112]), .Z(n640) );
  XNOR U996 ( .A(n659), .B(n660), .Z(n641) );
  XOR U997 ( .A(n657), .B(n671), .Z(n660) );
  NAND U998 ( .A(b[1]), .B(a[111]), .Z(n671) );
  XOR U999 ( .A(n665), .B(n672), .Z(n659) );
  XOR U1000 ( .A(n657), .B(n664), .Z(n672) );
  XNOR U1001 ( .A(n673), .B(n663), .Z(n664) );
  AND U1002 ( .A(b[2]), .B(a[110]), .Z(n673) );
  NANDN U1003 ( .A(n674), .B(n675), .Z(n657) );
  XNOR U1004 ( .A(n663), .B(n656), .Z(n676) );
  XOR U1005 ( .A(n677), .B(n678), .Z(n656) );
  XOR U1006 ( .A(n654), .B(n679), .Z(n678) );
  XOR U1007 ( .A(n680), .B(n681), .Z(n679) );
  XNOR U1008 ( .A(n682), .B(n683), .Z(n681) );
  AND U1009 ( .A(b[5]), .B(a[107]), .Z(n682) );
  XOR U1010 ( .A(n684), .B(n685), .Z(n680) );
  AND U1011 ( .A(b[6]), .B(a[106]), .Z(n685) );
  AND U1012 ( .A(b[7]), .B(a[105]), .Z(n684) );
  XOR U1013 ( .A(n686), .B(n683), .Z(n677) );
  XOR U1014 ( .A(n687), .B(n688), .Z(n683) );
  NOR U1015 ( .A(n689), .B(n690), .Z(n687) );
  AND U1016 ( .A(b[4]), .B(a[108]), .Z(n686) );
  XNOR U1017 ( .A(n691), .B(n692), .Z(n663) );
  NANDN U1018 ( .A(n693), .B(n694), .Z(n692) );
  XNOR U1019 ( .A(n695), .B(n654), .Z(n655) );
  XNOR U1020 ( .A(n696), .B(n697), .Z(n654) );
  AND U1021 ( .A(n698), .B(n699), .Z(n696) );
  AND U1022 ( .A(b[3]), .B(a[109]), .Z(n695) );
  XOR U1023 ( .A(n670), .B(n669), .Z(swire[111]) );
  XOR U1024 ( .A(sreg[239]), .B(n668), .Z(n669) );
  XOR U1025 ( .A(n675), .B(n700), .Z(n670) );
  XNOR U1026 ( .A(n674), .B(n668), .Z(n700) );
  XOR U1027 ( .A(n701), .B(n702), .Z(n668) );
  NOR U1028 ( .A(n703), .B(n704), .Z(n701) );
  NANDN U1029 ( .A(n187), .B(a[111]), .Z(n674) );
  XNOR U1030 ( .A(n693), .B(n694), .Z(n675) );
  XOR U1031 ( .A(n691), .B(n705), .Z(n694) );
  NAND U1032 ( .A(b[1]), .B(a[110]), .Z(n705) );
  XOR U1033 ( .A(n699), .B(n706), .Z(n693) );
  XOR U1034 ( .A(n691), .B(n698), .Z(n706) );
  XNOR U1035 ( .A(n707), .B(n697), .Z(n698) );
  AND U1036 ( .A(b[2]), .B(a[109]), .Z(n707) );
  NANDN U1037 ( .A(n708), .B(n709), .Z(n691) );
  XNOR U1038 ( .A(n697), .B(n690), .Z(n710) );
  XOR U1039 ( .A(n711), .B(n712), .Z(n690) );
  XOR U1040 ( .A(n688), .B(n713), .Z(n712) );
  XOR U1041 ( .A(n714), .B(n715), .Z(n713) );
  XNOR U1042 ( .A(n716), .B(n717), .Z(n715) );
  AND U1043 ( .A(b[5]), .B(a[106]), .Z(n716) );
  XOR U1044 ( .A(n718), .B(n719), .Z(n714) );
  AND U1045 ( .A(b[6]), .B(a[105]), .Z(n719) );
  AND U1046 ( .A(b[7]), .B(a[104]), .Z(n718) );
  XOR U1047 ( .A(n720), .B(n717), .Z(n711) );
  XOR U1048 ( .A(n721), .B(n722), .Z(n717) );
  NOR U1049 ( .A(n723), .B(n724), .Z(n721) );
  AND U1050 ( .A(b[4]), .B(a[107]), .Z(n720) );
  XNOR U1051 ( .A(n725), .B(n726), .Z(n697) );
  NANDN U1052 ( .A(n727), .B(n728), .Z(n726) );
  XNOR U1053 ( .A(n729), .B(n688), .Z(n689) );
  XNOR U1054 ( .A(n730), .B(n731), .Z(n688) );
  AND U1055 ( .A(n732), .B(n733), .Z(n730) );
  AND U1056 ( .A(b[3]), .B(a[108]), .Z(n729) );
  XOR U1057 ( .A(n704), .B(n703), .Z(swire[110]) );
  XOR U1058 ( .A(sreg[238]), .B(n702), .Z(n703) );
  XOR U1059 ( .A(n709), .B(n734), .Z(n704) );
  XNOR U1060 ( .A(n708), .B(n702), .Z(n734) );
  XOR U1061 ( .A(n735), .B(n736), .Z(n702) );
  NOR U1062 ( .A(n737), .B(n738), .Z(n735) );
  NANDN U1063 ( .A(n187), .B(a[110]), .Z(n708) );
  XNOR U1064 ( .A(n727), .B(n728), .Z(n709) );
  XOR U1065 ( .A(n725), .B(n739), .Z(n728) );
  NAND U1066 ( .A(b[1]), .B(a[109]), .Z(n739) );
  XOR U1067 ( .A(n733), .B(n740), .Z(n727) );
  XOR U1068 ( .A(n725), .B(n732), .Z(n740) );
  XNOR U1069 ( .A(n741), .B(n731), .Z(n732) );
  AND U1070 ( .A(b[2]), .B(a[108]), .Z(n741) );
  NANDN U1071 ( .A(n742), .B(n743), .Z(n725) );
  XNOR U1072 ( .A(n731), .B(n724), .Z(n744) );
  XOR U1073 ( .A(n745), .B(n746), .Z(n724) );
  XOR U1074 ( .A(n722), .B(n747), .Z(n746) );
  XOR U1075 ( .A(n748), .B(n749), .Z(n747) );
  XNOR U1076 ( .A(n750), .B(n751), .Z(n749) );
  AND U1077 ( .A(b[5]), .B(a[105]), .Z(n750) );
  XOR U1078 ( .A(n752), .B(n753), .Z(n748) );
  AND U1079 ( .A(b[6]), .B(a[104]), .Z(n753) );
  AND U1080 ( .A(b[7]), .B(a[103]), .Z(n752) );
  XOR U1081 ( .A(n754), .B(n751), .Z(n745) );
  XOR U1082 ( .A(n755), .B(n756), .Z(n751) );
  NOR U1083 ( .A(n757), .B(n758), .Z(n755) );
  AND U1084 ( .A(b[4]), .B(a[106]), .Z(n754) );
  XNOR U1085 ( .A(n759), .B(n760), .Z(n731) );
  NANDN U1086 ( .A(n761), .B(n762), .Z(n760) );
  XNOR U1087 ( .A(n763), .B(n722), .Z(n723) );
  XNOR U1088 ( .A(n764), .B(n765), .Z(n722) );
  AND U1089 ( .A(n766), .B(n767), .Z(n764) );
  AND U1090 ( .A(b[3]), .B(a[107]), .Z(n763) );
  XNOR U1091 ( .A(n768), .B(n769), .Z(swire[10]) );
  XOR U1092 ( .A(n738), .B(n737), .Z(swire[109]) );
  XOR U1093 ( .A(sreg[237]), .B(n736), .Z(n737) );
  XOR U1094 ( .A(n743), .B(n770), .Z(n738) );
  XNOR U1095 ( .A(n742), .B(n736), .Z(n770) );
  XOR U1096 ( .A(n771), .B(n772), .Z(n736) );
  NOR U1097 ( .A(n773), .B(n774), .Z(n771) );
  NANDN U1098 ( .A(n187), .B(a[109]), .Z(n742) );
  XNOR U1099 ( .A(n761), .B(n762), .Z(n743) );
  XOR U1100 ( .A(n759), .B(n775), .Z(n762) );
  NAND U1101 ( .A(b[1]), .B(a[108]), .Z(n775) );
  XOR U1102 ( .A(n767), .B(n776), .Z(n761) );
  XOR U1103 ( .A(n759), .B(n766), .Z(n776) );
  XNOR U1104 ( .A(n777), .B(n765), .Z(n766) );
  AND U1105 ( .A(b[2]), .B(a[107]), .Z(n777) );
  NANDN U1106 ( .A(n778), .B(n779), .Z(n759) );
  XNOR U1107 ( .A(n765), .B(n758), .Z(n780) );
  XOR U1108 ( .A(n781), .B(n782), .Z(n758) );
  XOR U1109 ( .A(n756), .B(n783), .Z(n782) );
  XOR U1110 ( .A(n784), .B(n785), .Z(n783) );
  XNOR U1111 ( .A(n786), .B(n787), .Z(n785) );
  AND U1112 ( .A(b[5]), .B(a[104]), .Z(n786) );
  XOR U1113 ( .A(n788), .B(n789), .Z(n784) );
  AND U1114 ( .A(b[6]), .B(a[103]), .Z(n789) );
  AND U1115 ( .A(b[7]), .B(a[102]), .Z(n788) );
  XOR U1116 ( .A(n790), .B(n787), .Z(n781) );
  XOR U1117 ( .A(n791), .B(n792), .Z(n787) );
  NOR U1118 ( .A(n793), .B(n794), .Z(n791) );
  AND U1119 ( .A(b[4]), .B(a[105]), .Z(n790) );
  XNOR U1120 ( .A(n795), .B(n796), .Z(n765) );
  NANDN U1121 ( .A(n797), .B(n798), .Z(n796) );
  XNOR U1122 ( .A(n799), .B(n756), .Z(n757) );
  XNOR U1123 ( .A(n800), .B(n801), .Z(n756) );
  AND U1124 ( .A(n802), .B(n803), .Z(n800) );
  AND U1125 ( .A(b[3]), .B(a[106]), .Z(n799) );
  XOR U1126 ( .A(n774), .B(n773), .Z(swire[108]) );
  XOR U1127 ( .A(sreg[236]), .B(n772), .Z(n773) );
  XOR U1128 ( .A(n779), .B(n804), .Z(n774) );
  XNOR U1129 ( .A(n778), .B(n772), .Z(n804) );
  XOR U1130 ( .A(n805), .B(n806), .Z(n772) );
  NOR U1131 ( .A(n807), .B(n808), .Z(n805) );
  NANDN U1132 ( .A(n187), .B(a[108]), .Z(n778) );
  XNOR U1133 ( .A(n797), .B(n798), .Z(n779) );
  XOR U1134 ( .A(n795), .B(n809), .Z(n798) );
  NAND U1135 ( .A(b[1]), .B(a[107]), .Z(n809) );
  XOR U1136 ( .A(n803), .B(n810), .Z(n797) );
  XOR U1137 ( .A(n795), .B(n802), .Z(n810) );
  XNOR U1138 ( .A(n811), .B(n801), .Z(n802) );
  AND U1139 ( .A(b[2]), .B(a[106]), .Z(n811) );
  NANDN U1140 ( .A(n812), .B(n813), .Z(n795) );
  XNOR U1141 ( .A(n801), .B(n794), .Z(n814) );
  XOR U1142 ( .A(n815), .B(n816), .Z(n794) );
  XOR U1143 ( .A(n792), .B(n817), .Z(n816) );
  XOR U1144 ( .A(n818), .B(n819), .Z(n817) );
  XNOR U1145 ( .A(n820), .B(n821), .Z(n819) );
  AND U1146 ( .A(b[5]), .B(a[103]), .Z(n820) );
  XOR U1147 ( .A(n822), .B(n823), .Z(n818) );
  AND U1148 ( .A(b[6]), .B(a[102]), .Z(n823) );
  AND U1149 ( .A(b[7]), .B(a[101]), .Z(n822) );
  XOR U1150 ( .A(n824), .B(n821), .Z(n815) );
  XOR U1151 ( .A(n825), .B(n826), .Z(n821) );
  NOR U1152 ( .A(n827), .B(n828), .Z(n825) );
  AND U1153 ( .A(b[4]), .B(a[104]), .Z(n824) );
  XNOR U1154 ( .A(n829), .B(n830), .Z(n801) );
  NANDN U1155 ( .A(n831), .B(n832), .Z(n830) );
  XNOR U1156 ( .A(n833), .B(n792), .Z(n793) );
  XNOR U1157 ( .A(n834), .B(n835), .Z(n792) );
  AND U1158 ( .A(n836), .B(n837), .Z(n834) );
  AND U1159 ( .A(b[3]), .B(a[105]), .Z(n833) );
  XOR U1160 ( .A(n808), .B(n807), .Z(swire[107]) );
  XOR U1161 ( .A(sreg[235]), .B(n806), .Z(n807) );
  XOR U1162 ( .A(n813), .B(n838), .Z(n808) );
  XNOR U1163 ( .A(n812), .B(n806), .Z(n838) );
  XOR U1164 ( .A(n839), .B(n840), .Z(n806) );
  NOR U1165 ( .A(n841), .B(n842), .Z(n839) );
  NANDN U1166 ( .A(n187), .B(a[107]), .Z(n812) );
  XNOR U1167 ( .A(n831), .B(n832), .Z(n813) );
  XOR U1168 ( .A(n829), .B(n843), .Z(n832) );
  NAND U1169 ( .A(b[1]), .B(a[106]), .Z(n843) );
  XOR U1170 ( .A(n837), .B(n844), .Z(n831) );
  XOR U1171 ( .A(n829), .B(n836), .Z(n844) );
  XNOR U1172 ( .A(n845), .B(n835), .Z(n836) );
  AND U1173 ( .A(b[2]), .B(a[105]), .Z(n845) );
  NANDN U1174 ( .A(n846), .B(n847), .Z(n829) );
  XNOR U1175 ( .A(n835), .B(n828), .Z(n848) );
  XOR U1176 ( .A(n849), .B(n850), .Z(n828) );
  XOR U1177 ( .A(n826), .B(n851), .Z(n850) );
  XOR U1178 ( .A(n852), .B(n853), .Z(n851) );
  XOR U1179 ( .A(n854), .B(n855), .Z(n853) );
  XOR U1180 ( .A(n856), .B(n857), .Z(n855) );
  XOR U1181 ( .A(n858), .B(n859), .Z(n857) );
  NAND U1182 ( .A(b[6]), .B(a[101]), .Z(n859) );
  AND U1183 ( .A(b[7]), .B(a[100]), .Z(n858) );
  XOR U1184 ( .A(n860), .B(n856), .Z(n852) );
  XOR U1185 ( .A(n861), .B(n862), .Z(n856) );
  NOR U1186 ( .A(n863), .B(n864), .Z(n861) );
  AND U1187 ( .A(b[5]), .B(a[102]), .Z(n860) );
  XOR U1188 ( .A(n865), .B(n854), .Z(n849) );
  XOR U1189 ( .A(n866), .B(n867), .Z(n854) );
  ANDN U1190 ( .B(n868), .A(n869), .Z(n866) );
  AND U1191 ( .A(b[4]), .B(a[103]), .Z(n865) );
  XNOR U1192 ( .A(n870), .B(n871), .Z(n835) );
  NANDN U1193 ( .A(n872), .B(n873), .Z(n871) );
  XNOR U1194 ( .A(n874), .B(n826), .Z(n827) );
  XNOR U1195 ( .A(n875), .B(n876), .Z(n826) );
  AND U1196 ( .A(n877), .B(n878), .Z(n875) );
  AND U1197 ( .A(b[3]), .B(a[104]), .Z(n874) );
  XOR U1198 ( .A(n842), .B(n841), .Z(swire[106]) );
  XOR U1199 ( .A(sreg[234]), .B(n840), .Z(n841) );
  XOR U1200 ( .A(n847), .B(n879), .Z(n842) );
  XNOR U1201 ( .A(n846), .B(n840), .Z(n879) );
  XOR U1202 ( .A(n880), .B(n881), .Z(n840) );
  NOR U1203 ( .A(n882), .B(n883), .Z(n880) );
  NANDN U1204 ( .A(n187), .B(a[106]), .Z(n846) );
  XNOR U1205 ( .A(n872), .B(n873), .Z(n847) );
  XOR U1206 ( .A(n870), .B(n884), .Z(n873) );
  NAND U1207 ( .A(b[1]), .B(a[105]), .Z(n884) );
  XOR U1208 ( .A(n878), .B(n885), .Z(n872) );
  XOR U1209 ( .A(n870), .B(n877), .Z(n885) );
  XNOR U1210 ( .A(n886), .B(n876), .Z(n877) );
  AND U1211 ( .A(b[2]), .B(a[104]), .Z(n886) );
  NANDN U1212 ( .A(n887), .B(n888), .Z(n870) );
  XOR U1213 ( .A(n876), .B(n868), .Z(n889) );
  XOR U1214 ( .A(n867), .B(n864), .Z(n890) );
  XOR U1215 ( .A(n891), .B(n892), .Z(n864) );
  XOR U1216 ( .A(n862), .B(n893), .Z(n892) );
  XOR U1217 ( .A(n894), .B(n895), .Z(n893) );
  XOR U1218 ( .A(n896), .B(n897), .Z(n895) );
  NAND U1219 ( .A(b[6]), .B(a[100]), .Z(n897) );
  AND U1220 ( .A(b[7]), .B(a[99]), .Z(n896) );
  XOR U1221 ( .A(n898), .B(n894), .Z(n891) );
  XOR U1222 ( .A(n899), .B(n900), .Z(n894) );
  NOR U1223 ( .A(n901), .B(n902), .Z(n899) );
  AND U1224 ( .A(b[5]), .B(a[101]), .Z(n898) );
  XNOR U1225 ( .A(n903), .B(n862), .Z(n863) );
  XOR U1226 ( .A(n904), .B(n905), .Z(n862) );
  ANDN U1227 ( .B(n906), .A(n907), .Z(n904) );
  AND U1228 ( .A(b[4]), .B(a[102]), .Z(n903) );
  XNOR U1229 ( .A(n908), .B(n909), .Z(n876) );
  NANDN U1230 ( .A(n910), .B(n911), .Z(n909) );
  XNOR U1231 ( .A(n912), .B(n867), .Z(n869) );
  XNOR U1232 ( .A(n913), .B(n914), .Z(n867) );
  AND U1233 ( .A(n915), .B(n916), .Z(n913) );
  AND U1234 ( .A(b[3]), .B(a[103]), .Z(n912) );
  XOR U1235 ( .A(n883), .B(n882), .Z(swire[105]) );
  XOR U1236 ( .A(sreg[233]), .B(n881), .Z(n882) );
  XOR U1237 ( .A(n888), .B(n917), .Z(n883) );
  XNOR U1238 ( .A(n887), .B(n881), .Z(n917) );
  XOR U1239 ( .A(n918), .B(n919), .Z(n881) );
  NOR U1240 ( .A(n920), .B(n921), .Z(n918) );
  NANDN U1241 ( .A(n187), .B(a[105]), .Z(n887) );
  XNOR U1242 ( .A(n910), .B(n911), .Z(n888) );
  XOR U1243 ( .A(n908), .B(n922), .Z(n911) );
  NAND U1244 ( .A(b[1]), .B(a[104]), .Z(n922) );
  XOR U1245 ( .A(n916), .B(n923), .Z(n910) );
  XOR U1246 ( .A(n908), .B(n915), .Z(n923) );
  XNOR U1247 ( .A(n924), .B(n914), .Z(n915) );
  AND U1248 ( .A(b[2]), .B(a[103]), .Z(n924) );
  NANDN U1249 ( .A(n925), .B(n926), .Z(n908) );
  XOR U1250 ( .A(n914), .B(n906), .Z(n927) );
  XOR U1251 ( .A(n905), .B(n902), .Z(n928) );
  XOR U1252 ( .A(n929), .B(n930), .Z(n902) );
  XOR U1253 ( .A(n900), .B(n931), .Z(n930) );
  XOR U1254 ( .A(n932), .B(n933), .Z(n931) );
  XOR U1255 ( .A(n934), .B(n935), .Z(n933) );
  NAND U1256 ( .A(b[6]), .B(a[99]), .Z(n935) );
  AND U1257 ( .A(b[7]), .B(a[98]), .Z(n934) );
  XOR U1258 ( .A(n936), .B(n932), .Z(n929) );
  XOR U1259 ( .A(n937), .B(n938), .Z(n932) );
  NOR U1260 ( .A(n939), .B(n940), .Z(n937) );
  AND U1261 ( .A(b[5]), .B(a[100]), .Z(n936) );
  XNOR U1262 ( .A(n941), .B(n900), .Z(n901) );
  XOR U1263 ( .A(n942), .B(n943), .Z(n900) );
  ANDN U1264 ( .B(n944), .A(n945), .Z(n942) );
  AND U1265 ( .A(b[4]), .B(a[101]), .Z(n941) );
  XNOR U1266 ( .A(n946), .B(n947), .Z(n914) );
  NANDN U1267 ( .A(n948), .B(n949), .Z(n947) );
  XNOR U1268 ( .A(n950), .B(n905), .Z(n907) );
  XNOR U1269 ( .A(n951), .B(n952), .Z(n905) );
  AND U1270 ( .A(n953), .B(n954), .Z(n951) );
  AND U1271 ( .A(b[3]), .B(a[102]), .Z(n950) );
  XOR U1272 ( .A(n921), .B(n920), .Z(swire[104]) );
  XOR U1273 ( .A(sreg[232]), .B(n919), .Z(n920) );
  XOR U1274 ( .A(n926), .B(n955), .Z(n921) );
  XNOR U1275 ( .A(n925), .B(n919), .Z(n955) );
  XOR U1276 ( .A(n956), .B(n957), .Z(n919) );
  NOR U1277 ( .A(n958), .B(n959), .Z(n956) );
  NANDN U1278 ( .A(n187), .B(a[104]), .Z(n925) );
  XNOR U1279 ( .A(n948), .B(n949), .Z(n926) );
  XOR U1280 ( .A(n946), .B(n960), .Z(n949) );
  NAND U1281 ( .A(b[1]), .B(a[103]), .Z(n960) );
  XOR U1282 ( .A(n954), .B(n961), .Z(n948) );
  XOR U1283 ( .A(n946), .B(n953), .Z(n961) );
  XNOR U1284 ( .A(n962), .B(n952), .Z(n953) );
  AND U1285 ( .A(b[2]), .B(a[102]), .Z(n962) );
  NANDN U1286 ( .A(n963), .B(n964), .Z(n946) );
  XOR U1287 ( .A(n952), .B(n944), .Z(n965) );
  XOR U1288 ( .A(n943), .B(n940), .Z(n966) );
  XOR U1289 ( .A(n967), .B(n968), .Z(n940) );
  XOR U1290 ( .A(n938), .B(n969), .Z(n968) );
  XOR U1291 ( .A(n970), .B(n971), .Z(n969) );
  XOR U1292 ( .A(n972), .B(n973), .Z(n971) );
  NAND U1293 ( .A(b[6]), .B(a[98]), .Z(n973) );
  AND U1294 ( .A(b[7]), .B(a[97]), .Z(n972) );
  XOR U1295 ( .A(n974), .B(n970), .Z(n967) );
  XOR U1296 ( .A(n975), .B(n976), .Z(n970) );
  NOR U1297 ( .A(n977), .B(n978), .Z(n975) );
  AND U1298 ( .A(b[5]), .B(a[99]), .Z(n974) );
  XNOR U1299 ( .A(n979), .B(n938), .Z(n939) );
  XOR U1300 ( .A(n980), .B(n981), .Z(n938) );
  ANDN U1301 ( .B(n982), .A(n983), .Z(n980) );
  AND U1302 ( .A(b[4]), .B(a[100]), .Z(n979) );
  XNOR U1303 ( .A(n984), .B(n985), .Z(n952) );
  NANDN U1304 ( .A(n986), .B(n987), .Z(n985) );
  XNOR U1305 ( .A(n988), .B(n943), .Z(n945) );
  XNOR U1306 ( .A(n989), .B(n990), .Z(n943) );
  AND U1307 ( .A(n991), .B(n992), .Z(n989) );
  AND U1308 ( .A(b[3]), .B(a[101]), .Z(n988) );
  XOR U1309 ( .A(n959), .B(n958), .Z(swire[103]) );
  XOR U1310 ( .A(sreg[231]), .B(n957), .Z(n958) );
  XOR U1311 ( .A(n964), .B(n993), .Z(n959) );
  XNOR U1312 ( .A(n963), .B(n957), .Z(n993) );
  XOR U1313 ( .A(n994), .B(n995), .Z(n957) );
  NOR U1314 ( .A(n996), .B(n997), .Z(n994) );
  NANDN U1315 ( .A(n187), .B(a[103]), .Z(n963) );
  XNOR U1316 ( .A(n986), .B(n987), .Z(n964) );
  XOR U1317 ( .A(n984), .B(n998), .Z(n987) );
  NAND U1318 ( .A(b[1]), .B(a[102]), .Z(n998) );
  XOR U1319 ( .A(n992), .B(n999), .Z(n986) );
  XOR U1320 ( .A(n984), .B(n991), .Z(n999) );
  XNOR U1321 ( .A(n1000), .B(n990), .Z(n991) );
  AND U1322 ( .A(b[2]), .B(a[101]), .Z(n1000) );
  NANDN U1323 ( .A(n1001), .B(n1002), .Z(n984) );
  XOR U1324 ( .A(n990), .B(n982), .Z(n1003) );
  XOR U1325 ( .A(n981), .B(n978), .Z(n1004) );
  XOR U1326 ( .A(n1005), .B(n1006), .Z(n978) );
  XOR U1327 ( .A(n976), .B(n1007), .Z(n1006) );
  XOR U1328 ( .A(n1008), .B(n1009), .Z(n1007) );
  XOR U1329 ( .A(n1010), .B(n1011), .Z(n1009) );
  NAND U1330 ( .A(b[6]), .B(a[97]), .Z(n1011) );
  AND U1331 ( .A(b[7]), .B(a[96]), .Z(n1010) );
  XOR U1332 ( .A(n1012), .B(n1008), .Z(n1005) );
  XOR U1333 ( .A(n1013), .B(n1014), .Z(n1008) );
  NOR U1334 ( .A(n1015), .B(n1016), .Z(n1013) );
  AND U1335 ( .A(b[5]), .B(a[98]), .Z(n1012) );
  XNOR U1336 ( .A(n1017), .B(n976), .Z(n977) );
  XOR U1337 ( .A(n1018), .B(n1019), .Z(n976) );
  ANDN U1338 ( .B(n1020), .A(n1021), .Z(n1018) );
  AND U1339 ( .A(b[4]), .B(a[99]), .Z(n1017) );
  XNOR U1340 ( .A(n1022), .B(n1023), .Z(n990) );
  NANDN U1341 ( .A(n1024), .B(n1025), .Z(n1023) );
  XNOR U1342 ( .A(n1026), .B(n981), .Z(n983) );
  XNOR U1343 ( .A(n1027), .B(n1028), .Z(n981) );
  AND U1344 ( .A(n1029), .B(n1030), .Z(n1027) );
  AND U1345 ( .A(b[3]), .B(a[100]), .Z(n1026) );
  XOR U1346 ( .A(n997), .B(n996), .Z(swire[102]) );
  XOR U1347 ( .A(sreg[230]), .B(n995), .Z(n996) );
  XOR U1348 ( .A(n1002), .B(n1031), .Z(n997) );
  XNOR U1349 ( .A(n1001), .B(n995), .Z(n1031) );
  XOR U1350 ( .A(n1032), .B(n1033), .Z(n995) );
  NOR U1351 ( .A(n1034), .B(n1035), .Z(n1032) );
  NANDN U1352 ( .A(n187), .B(a[102]), .Z(n1001) );
  XNOR U1353 ( .A(n1024), .B(n1025), .Z(n1002) );
  XOR U1354 ( .A(n1022), .B(n1036), .Z(n1025) );
  NAND U1355 ( .A(b[1]), .B(a[101]), .Z(n1036) );
  XOR U1356 ( .A(n1030), .B(n1037), .Z(n1024) );
  XOR U1357 ( .A(n1022), .B(n1029), .Z(n1037) );
  XNOR U1358 ( .A(n1038), .B(n1028), .Z(n1029) );
  AND U1359 ( .A(b[2]), .B(a[100]), .Z(n1038) );
  NANDN U1360 ( .A(n1039), .B(n1040), .Z(n1022) );
  XOR U1361 ( .A(n1028), .B(n1020), .Z(n1041) );
  XOR U1362 ( .A(n1019), .B(n1016), .Z(n1042) );
  XOR U1363 ( .A(n1043), .B(n1044), .Z(n1016) );
  XOR U1364 ( .A(n1014), .B(n1045), .Z(n1044) );
  XOR U1365 ( .A(n1046), .B(n1047), .Z(n1045) );
  XOR U1366 ( .A(n1048), .B(n1049), .Z(n1047) );
  NAND U1367 ( .A(b[6]), .B(a[96]), .Z(n1049) );
  AND U1368 ( .A(b[7]), .B(a[95]), .Z(n1048) );
  XOR U1369 ( .A(n1050), .B(n1046), .Z(n1043) );
  XOR U1370 ( .A(n1051), .B(n1052), .Z(n1046) );
  NOR U1371 ( .A(n1053), .B(n1054), .Z(n1051) );
  AND U1372 ( .A(b[5]), .B(a[97]), .Z(n1050) );
  XNOR U1373 ( .A(n1055), .B(n1014), .Z(n1015) );
  XOR U1374 ( .A(n1056), .B(n1057), .Z(n1014) );
  ANDN U1375 ( .B(n1058), .A(n1059), .Z(n1056) );
  AND U1376 ( .A(b[4]), .B(a[98]), .Z(n1055) );
  XNOR U1377 ( .A(n1060), .B(n1061), .Z(n1028) );
  NANDN U1378 ( .A(n1062), .B(n1063), .Z(n1061) );
  XNOR U1379 ( .A(n1064), .B(n1019), .Z(n1021) );
  XNOR U1380 ( .A(n1065), .B(n1066), .Z(n1019) );
  AND U1381 ( .A(n1067), .B(n1068), .Z(n1065) );
  AND U1382 ( .A(b[3]), .B(a[99]), .Z(n1064) );
  XOR U1383 ( .A(n1035), .B(n1034), .Z(swire[101]) );
  XOR U1384 ( .A(sreg[229]), .B(n1033), .Z(n1034) );
  XOR U1385 ( .A(n1040), .B(n1069), .Z(n1035) );
  XNOR U1386 ( .A(n1039), .B(n1033), .Z(n1069) );
  XOR U1387 ( .A(n1070), .B(n1071), .Z(n1033) );
  NOR U1388 ( .A(n1072), .B(n1073), .Z(n1070) );
  NANDN U1389 ( .A(n187), .B(a[101]), .Z(n1039) );
  XNOR U1390 ( .A(n1062), .B(n1063), .Z(n1040) );
  XOR U1391 ( .A(n1060), .B(n1074), .Z(n1063) );
  NAND U1392 ( .A(b[1]), .B(a[100]), .Z(n1074) );
  XOR U1393 ( .A(n1068), .B(n1075), .Z(n1062) );
  XOR U1394 ( .A(n1060), .B(n1067), .Z(n1075) );
  XNOR U1395 ( .A(n1076), .B(n1066), .Z(n1067) );
  AND U1396 ( .A(b[2]), .B(a[99]), .Z(n1076) );
  NANDN U1397 ( .A(n1077), .B(n1078), .Z(n1060) );
  XOR U1398 ( .A(n1066), .B(n1058), .Z(n1079) );
  XOR U1399 ( .A(n1057), .B(n1054), .Z(n1080) );
  XOR U1400 ( .A(n1081), .B(n1082), .Z(n1054) );
  XOR U1401 ( .A(n1052), .B(n1083), .Z(n1082) );
  XOR U1402 ( .A(n1084), .B(n1085), .Z(n1083) );
  XOR U1403 ( .A(n1086), .B(n1087), .Z(n1085) );
  NAND U1404 ( .A(b[6]), .B(a[95]), .Z(n1087) );
  AND U1405 ( .A(b[7]), .B(a[94]), .Z(n1086) );
  XOR U1406 ( .A(n1088), .B(n1084), .Z(n1081) );
  XOR U1407 ( .A(n1089), .B(n1090), .Z(n1084) );
  NOR U1408 ( .A(n1091), .B(n1092), .Z(n1089) );
  AND U1409 ( .A(b[5]), .B(a[96]), .Z(n1088) );
  XNOR U1410 ( .A(n1093), .B(n1052), .Z(n1053) );
  XOR U1411 ( .A(n1094), .B(n1095), .Z(n1052) );
  ANDN U1412 ( .B(n1096), .A(n1097), .Z(n1094) );
  AND U1413 ( .A(b[4]), .B(a[97]), .Z(n1093) );
  XNOR U1414 ( .A(n1098), .B(n1099), .Z(n1066) );
  NANDN U1415 ( .A(n1100), .B(n1101), .Z(n1099) );
  XNOR U1416 ( .A(n1102), .B(n1057), .Z(n1059) );
  XNOR U1417 ( .A(n1103), .B(n1104), .Z(n1057) );
  AND U1418 ( .A(n1105), .B(n1106), .Z(n1103) );
  AND U1419 ( .A(b[3]), .B(a[98]), .Z(n1102) );
  XOR U1420 ( .A(n1073), .B(n1072), .Z(swire[100]) );
  XOR U1421 ( .A(sreg[228]), .B(n1071), .Z(n1072) );
  XOR U1422 ( .A(n1078), .B(n1107), .Z(n1073) );
  XNOR U1423 ( .A(n1077), .B(n1071), .Z(n1107) );
  XOR U1424 ( .A(n1108), .B(n1109), .Z(n1071) );
  ANDN U1425 ( .B(n4), .A(n3), .Z(n1108) );
  XOR U1426 ( .A(sreg[227]), .B(n1109), .Z(n3) );
  XOR U1427 ( .A(n1110), .B(n1111), .Z(n4) );
  XNOR U1428 ( .A(n1112), .B(n1109), .Z(n1111) );
  XOR U1429 ( .A(n1113), .B(n1114), .Z(n1109) );
  ANDN U1430 ( .B(n5), .A(n6), .Z(n1113) );
  XOR U1431 ( .A(sreg[226]), .B(n1114), .Z(n6) );
  XOR U1432 ( .A(n1115), .B(n1116), .Z(n5) );
  XNOR U1433 ( .A(n1117), .B(n1114), .Z(n1116) );
  XOR U1434 ( .A(n1118), .B(n1119), .Z(n1114) );
  ANDN U1435 ( .B(n7), .A(n8), .Z(n1118) );
  XOR U1436 ( .A(sreg[225]), .B(n1119), .Z(n8) );
  XOR U1437 ( .A(n1120), .B(n1121), .Z(n7) );
  XNOR U1438 ( .A(n1122), .B(n1119), .Z(n1121) );
  XOR U1439 ( .A(n1123), .B(n1124), .Z(n1119) );
  ANDN U1440 ( .B(n9), .A(n10), .Z(n1123) );
  XOR U1441 ( .A(sreg[224]), .B(n1124), .Z(n10) );
  XOR U1442 ( .A(n1125), .B(n1126), .Z(n9) );
  XNOR U1443 ( .A(n1127), .B(n1124), .Z(n1126) );
  XOR U1444 ( .A(n1128), .B(n1129), .Z(n1124) );
  ANDN U1445 ( .B(n11), .A(n12), .Z(n1128) );
  XOR U1446 ( .A(sreg[223]), .B(n1129), .Z(n12) );
  XOR U1447 ( .A(n1130), .B(n1131), .Z(n11) );
  XNOR U1448 ( .A(n1132), .B(n1129), .Z(n1131) );
  XOR U1449 ( .A(n1133), .B(n1134), .Z(n1129) );
  ANDN U1450 ( .B(n13), .A(n14), .Z(n1133) );
  XOR U1451 ( .A(sreg[222]), .B(n1134), .Z(n14) );
  XOR U1452 ( .A(n1135), .B(n1136), .Z(n13) );
  XNOR U1453 ( .A(n1137), .B(n1134), .Z(n1136) );
  XOR U1454 ( .A(n1138), .B(n1139), .Z(n1134) );
  ANDN U1455 ( .B(n15), .A(n16), .Z(n1138) );
  XOR U1456 ( .A(sreg[221]), .B(n1139), .Z(n16) );
  XOR U1457 ( .A(n1140), .B(n1141), .Z(n15) );
  XNOR U1458 ( .A(n1142), .B(n1139), .Z(n1141) );
  XOR U1459 ( .A(n1143), .B(n1144), .Z(n1139) );
  ANDN U1460 ( .B(n17), .A(n18), .Z(n1143) );
  XOR U1461 ( .A(sreg[220]), .B(n1144), .Z(n18) );
  XOR U1462 ( .A(n1145), .B(n1146), .Z(n17) );
  XNOR U1463 ( .A(n1147), .B(n1144), .Z(n1146) );
  XOR U1464 ( .A(n1148), .B(n1149), .Z(n1144) );
  ANDN U1465 ( .B(n19), .A(n20), .Z(n1148) );
  XOR U1466 ( .A(sreg[219]), .B(n1149), .Z(n20) );
  XOR U1467 ( .A(n1150), .B(n1151), .Z(n19) );
  XNOR U1468 ( .A(n1152), .B(n1149), .Z(n1151) );
  XOR U1469 ( .A(n1153), .B(n1154), .Z(n1149) );
  ANDN U1470 ( .B(n21), .A(n22), .Z(n1153) );
  XOR U1471 ( .A(sreg[218]), .B(n1154), .Z(n22) );
  XOR U1472 ( .A(n1155), .B(n1156), .Z(n21) );
  XNOR U1473 ( .A(n1157), .B(n1154), .Z(n1156) );
  XOR U1474 ( .A(n1158), .B(n1159), .Z(n1154) );
  ANDN U1475 ( .B(n25), .A(n26), .Z(n1158) );
  XOR U1476 ( .A(sreg[217]), .B(n1159), .Z(n26) );
  XOR U1477 ( .A(n1160), .B(n1161), .Z(n25) );
  XNOR U1478 ( .A(n1162), .B(n1159), .Z(n1161) );
  XOR U1479 ( .A(n1163), .B(n1164), .Z(n1159) );
  ANDN U1480 ( .B(n27), .A(n28), .Z(n1163) );
  XOR U1481 ( .A(sreg[216]), .B(n1164), .Z(n28) );
  XOR U1482 ( .A(n1165), .B(n1166), .Z(n27) );
  XNOR U1483 ( .A(n1167), .B(n1164), .Z(n1166) );
  XOR U1484 ( .A(n1168), .B(n1169), .Z(n1164) );
  ANDN U1485 ( .B(n29), .A(n30), .Z(n1168) );
  XOR U1486 ( .A(sreg[215]), .B(n1169), .Z(n30) );
  XOR U1487 ( .A(n1170), .B(n1171), .Z(n29) );
  XNOR U1488 ( .A(n1172), .B(n1169), .Z(n1171) );
  XOR U1489 ( .A(n1173), .B(n1174), .Z(n1169) );
  ANDN U1490 ( .B(n31), .A(n32), .Z(n1173) );
  XOR U1491 ( .A(sreg[214]), .B(n1174), .Z(n32) );
  XOR U1492 ( .A(n1175), .B(n1176), .Z(n31) );
  XNOR U1493 ( .A(n1177), .B(n1174), .Z(n1176) );
  XOR U1494 ( .A(n1178), .B(n1179), .Z(n1174) );
  ANDN U1495 ( .B(n33), .A(n34), .Z(n1178) );
  XOR U1496 ( .A(sreg[213]), .B(n1179), .Z(n34) );
  XOR U1497 ( .A(n1180), .B(n1181), .Z(n33) );
  XNOR U1498 ( .A(n1182), .B(n1179), .Z(n1181) );
  XOR U1499 ( .A(n1183), .B(n1184), .Z(n1179) );
  ANDN U1500 ( .B(n35), .A(n36), .Z(n1183) );
  XOR U1501 ( .A(sreg[212]), .B(n1184), .Z(n36) );
  XOR U1502 ( .A(n1185), .B(n1186), .Z(n35) );
  XNOR U1503 ( .A(n1187), .B(n1184), .Z(n1186) );
  XOR U1504 ( .A(n1188), .B(n1189), .Z(n1184) );
  ANDN U1505 ( .B(n37), .A(n38), .Z(n1188) );
  XOR U1506 ( .A(sreg[211]), .B(n1189), .Z(n38) );
  XOR U1507 ( .A(n1190), .B(n1191), .Z(n37) );
  XNOR U1508 ( .A(n1192), .B(n1189), .Z(n1191) );
  XOR U1509 ( .A(n1193), .B(n1194), .Z(n1189) );
  ANDN U1510 ( .B(n39), .A(n40), .Z(n1193) );
  XOR U1511 ( .A(sreg[210]), .B(n1194), .Z(n40) );
  XOR U1512 ( .A(n1195), .B(n1196), .Z(n39) );
  XNOR U1513 ( .A(n1197), .B(n1194), .Z(n1196) );
  XOR U1514 ( .A(n1198), .B(n1199), .Z(n1194) );
  ANDN U1515 ( .B(n41), .A(n42), .Z(n1198) );
  XOR U1516 ( .A(sreg[209]), .B(n1199), .Z(n42) );
  XOR U1517 ( .A(n1200), .B(n1201), .Z(n41) );
  XNOR U1518 ( .A(n1202), .B(n1199), .Z(n1201) );
  XOR U1519 ( .A(n1203), .B(n1204), .Z(n1199) );
  ANDN U1520 ( .B(n43), .A(n44), .Z(n1203) );
  XOR U1521 ( .A(sreg[208]), .B(n1204), .Z(n44) );
  XOR U1522 ( .A(n1205), .B(n1206), .Z(n43) );
  XNOR U1523 ( .A(n1207), .B(n1204), .Z(n1206) );
  XOR U1524 ( .A(n1208), .B(n1209), .Z(n1204) );
  ANDN U1525 ( .B(n45), .A(n46), .Z(n1208) );
  XOR U1526 ( .A(sreg[207]), .B(n1209), .Z(n46) );
  XOR U1527 ( .A(n1210), .B(n1211), .Z(n45) );
  XNOR U1528 ( .A(n1212), .B(n1209), .Z(n1211) );
  XOR U1529 ( .A(n1213), .B(n1214), .Z(n1209) );
  ANDN U1530 ( .B(n47), .A(n48), .Z(n1213) );
  XOR U1531 ( .A(sreg[206]), .B(n1214), .Z(n48) );
  XOR U1532 ( .A(n1215), .B(n1216), .Z(n47) );
  XNOR U1533 ( .A(n1217), .B(n1214), .Z(n1216) );
  XOR U1534 ( .A(n1218), .B(n1219), .Z(n1214) );
  ANDN U1535 ( .B(n49), .A(n50), .Z(n1218) );
  XOR U1536 ( .A(sreg[205]), .B(n1219), .Z(n50) );
  XOR U1537 ( .A(n1220), .B(n1221), .Z(n49) );
  XNOR U1538 ( .A(n1222), .B(n1219), .Z(n1221) );
  XOR U1539 ( .A(n1223), .B(n1224), .Z(n1219) );
  ANDN U1540 ( .B(n51), .A(n52), .Z(n1223) );
  XOR U1541 ( .A(sreg[204]), .B(n1224), .Z(n52) );
  XOR U1542 ( .A(n1225), .B(n1226), .Z(n51) );
  XNOR U1543 ( .A(n1227), .B(n1224), .Z(n1226) );
  XOR U1544 ( .A(n1228), .B(n1229), .Z(n1224) );
  ANDN U1545 ( .B(n53), .A(n54), .Z(n1228) );
  XOR U1546 ( .A(sreg[203]), .B(n1229), .Z(n54) );
  XOR U1547 ( .A(n1230), .B(n1231), .Z(n53) );
  XNOR U1548 ( .A(n1232), .B(n1229), .Z(n1231) );
  XOR U1549 ( .A(n1233), .B(n1234), .Z(n1229) );
  ANDN U1550 ( .B(n55), .A(n56), .Z(n1233) );
  XOR U1551 ( .A(sreg[202]), .B(n1234), .Z(n56) );
  XOR U1552 ( .A(n1235), .B(n1236), .Z(n55) );
  XNOR U1553 ( .A(n1237), .B(n1234), .Z(n1236) );
  XOR U1554 ( .A(n1238), .B(n1239), .Z(n1234) );
  ANDN U1555 ( .B(n57), .A(n58), .Z(n1238) );
  XOR U1556 ( .A(sreg[201]), .B(n1239), .Z(n58) );
  XOR U1557 ( .A(n1240), .B(n1241), .Z(n57) );
  XNOR U1558 ( .A(n1242), .B(n1239), .Z(n1241) );
  XOR U1559 ( .A(n1243), .B(n1244), .Z(n1239) );
  ANDN U1560 ( .B(n59), .A(n60), .Z(n1243) );
  XOR U1561 ( .A(sreg[200]), .B(n1244), .Z(n60) );
  XOR U1562 ( .A(n1245), .B(n1246), .Z(n59) );
  XNOR U1563 ( .A(n1247), .B(n1244), .Z(n1246) );
  XOR U1564 ( .A(n1248), .B(n1249), .Z(n1244) );
  ANDN U1565 ( .B(n61), .A(n62), .Z(n1248) );
  XOR U1566 ( .A(sreg[199]), .B(n1249), .Z(n62) );
  XOR U1567 ( .A(n1250), .B(n1251), .Z(n61) );
  XNOR U1568 ( .A(n1252), .B(n1249), .Z(n1251) );
  XOR U1569 ( .A(n1253), .B(n1254), .Z(n1249) );
  ANDN U1570 ( .B(n63), .A(n64), .Z(n1253) );
  XOR U1571 ( .A(sreg[198]), .B(n1254), .Z(n64) );
  XOR U1572 ( .A(n1255), .B(n1256), .Z(n63) );
  XNOR U1573 ( .A(n1257), .B(n1254), .Z(n1256) );
  XOR U1574 ( .A(n1258), .B(n1259), .Z(n1254) );
  ANDN U1575 ( .B(n65), .A(n66), .Z(n1258) );
  XOR U1576 ( .A(sreg[197]), .B(n1259), .Z(n66) );
  XOR U1577 ( .A(n1260), .B(n1261), .Z(n65) );
  XNOR U1578 ( .A(n1262), .B(n1259), .Z(n1261) );
  XOR U1579 ( .A(n1263), .B(n1264), .Z(n1259) );
  ANDN U1580 ( .B(n67), .A(n68), .Z(n1263) );
  XOR U1581 ( .A(sreg[196]), .B(n1264), .Z(n68) );
  XOR U1582 ( .A(n1265), .B(n1266), .Z(n67) );
  XNOR U1583 ( .A(n1267), .B(n1264), .Z(n1266) );
  XOR U1584 ( .A(n1268), .B(n1269), .Z(n1264) );
  ANDN U1585 ( .B(n69), .A(n70), .Z(n1268) );
  XOR U1586 ( .A(sreg[195]), .B(n1269), .Z(n70) );
  XOR U1587 ( .A(n1270), .B(n1271), .Z(n69) );
  XNOR U1588 ( .A(n1272), .B(n1269), .Z(n1271) );
  XOR U1589 ( .A(n1273), .B(n1274), .Z(n1269) );
  ANDN U1590 ( .B(n71), .A(n72), .Z(n1273) );
  XOR U1591 ( .A(sreg[194]), .B(n1274), .Z(n72) );
  XOR U1592 ( .A(n1275), .B(n1276), .Z(n71) );
  XNOR U1593 ( .A(n1277), .B(n1274), .Z(n1276) );
  XOR U1594 ( .A(n1278), .B(n1279), .Z(n1274) );
  ANDN U1595 ( .B(n73), .A(n74), .Z(n1278) );
  XOR U1596 ( .A(sreg[193]), .B(n1279), .Z(n74) );
  XOR U1597 ( .A(n1280), .B(n1281), .Z(n73) );
  XNOR U1598 ( .A(n1282), .B(n1279), .Z(n1281) );
  XOR U1599 ( .A(n1283), .B(n1284), .Z(n1279) );
  ANDN U1600 ( .B(n75), .A(n76), .Z(n1283) );
  XOR U1601 ( .A(sreg[192]), .B(n1284), .Z(n76) );
  XOR U1602 ( .A(n1285), .B(n1286), .Z(n75) );
  XNOR U1603 ( .A(n1287), .B(n1284), .Z(n1286) );
  XOR U1604 ( .A(n1288), .B(n1289), .Z(n1284) );
  ANDN U1605 ( .B(n77), .A(n78), .Z(n1288) );
  XOR U1606 ( .A(sreg[191]), .B(n1289), .Z(n78) );
  XOR U1607 ( .A(n1290), .B(n1291), .Z(n77) );
  XNOR U1608 ( .A(n1292), .B(n1289), .Z(n1291) );
  XOR U1609 ( .A(n1293), .B(n1294), .Z(n1289) );
  ANDN U1610 ( .B(n79), .A(n80), .Z(n1293) );
  XOR U1611 ( .A(sreg[190]), .B(n1294), .Z(n80) );
  XOR U1612 ( .A(n1295), .B(n1296), .Z(n79) );
  XNOR U1613 ( .A(n1297), .B(n1294), .Z(n1296) );
  XOR U1614 ( .A(n1298), .B(n1299), .Z(n1294) );
  ANDN U1615 ( .B(n81), .A(n82), .Z(n1298) );
  XOR U1616 ( .A(sreg[189]), .B(n1299), .Z(n82) );
  XOR U1617 ( .A(n1300), .B(n1301), .Z(n81) );
  XNOR U1618 ( .A(n1302), .B(n1299), .Z(n1301) );
  XOR U1619 ( .A(n1303), .B(n1304), .Z(n1299) );
  ANDN U1620 ( .B(n83), .A(n84), .Z(n1303) );
  XOR U1621 ( .A(sreg[188]), .B(n1304), .Z(n84) );
  XOR U1622 ( .A(n1305), .B(n1306), .Z(n83) );
  XNOR U1623 ( .A(n1307), .B(n1304), .Z(n1306) );
  XOR U1624 ( .A(n1308), .B(n1309), .Z(n1304) );
  ANDN U1625 ( .B(n85), .A(n86), .Z(n1308) );
  XOR U1626 ( .A(sreg[187]), .B(n1309), .Z(n86) );
  XOR U1627 ( .A(n1310), .B(n1311), .Z(n85) );
  XNOR U1628 ( .A(n1312), .B(n1309), .Z(n1311) );
  XOR U1629 ( .A(n1313), .B(n1314), .Z(n1309) );
  ANDN U1630 ( .B(n87), .A(n88), .Z(n1313) );
  XOR U1631 ( .A(sreg[186]), .B(n1314), .Z(n88) );
  XOR U1632 ( .A(n1315), .B(n1316), .Z(n87) );
  XNOR U1633 ( .A(n1317), .B(n1314), .Z(n1316) );
  XOR U1634 ( .A(n1318), .B(n1319), .Z(n1314) );
  ANDN U1635 ( .B(n89), .A(n90), .Z(n1318) );
  XOR U1636 ( .A(sreg[185]), .B(n1319), .Z(n90) );
  XOR U1637 ( .A(n1320), .B(n1321), .Z(n89) );
  XNOR U1638 ( .A(n1322), .B(n1319), .Z(n1321) );
  XOR U1639 ( .A(n1323), .B(n1324), .Z(n1319) );
  ANDN U1640 ( .B(n91), .A(n92), .Z(n1323) );
  XOR U1641 ( .A(sreg[184]), .B(n1324), .Z(n92) );
  XOR U1642 ( .A(n1325), .B(n1326), .Z(n91) );
  XNOR U1643 ( .A(n1327), .B(n1324), .Z(n1326) );
  XOR U1644 ( .A(n1328), .B(n1329), .Z(n1324) );
  ANDN U1645 ( .B(n93), .A(n94), .Z(n1328) );
  XOR U1646 ( .A(sreg[183]), .B(n1329), .Z(n94) );
  XOR U1647 ( .A(n1330), .B(n1331), .Z(n93) );
  XNOR U1648 ( .A(n1332), .B(n1329), .Z(n1331) );
  XOR U1649 ( .A(n1333), .B(n1334), .Z(n1329) );
  ANDN U1650 ( .B(n95), .A(n96), .Z(n1333) );
  XOR U1651 ( .A(sreg[182]), .B(n1334), .Z(n96) );
  XOR U1652 ( .A(n1335), .B(n1336), .Z(n95) );
  XNOR U1653 ( .A(n1337), .B(n1334), .Z(n1336) );
  XOR U1654 ( .A(n1338), .B(n1339), .Z(n1334) );
  ANDN U1655 ( .B(n97), .A(n98), .Z(n1338) );
  XOR U1656 ( .A(sreg[181]), .B(n1339), .Z(n98) );
  XOR U1657 ( .A(n1340), .B(n1341), .Z(n97) );
  XNOR U1658 ( .A(n1342), .B(n1339), .Z(n1341) );
  XOR U1659 ( .A(n1343), .B(n1344), .Z(n1339) );
  ANDN U1660 ( .B(n99), .A(n100), .Z(n1343) );
  XOR U1661 ( .A(sreg[180]), .B(n1344), .Z(n100) );
  XOR U1662 ( .A(n1345), .B(n1346), .Z(n99) );
  XNOR U1663 ( .A(n1347), .B(n1344), .Z(n1346) );
  XOR U1664 ( .A(n1348), .B(n1349), .Z(n1344) );
  ANDN U1665 ( .B(n101), .A(n102), .Z(n1348) );
  XOR U1666 ( .A(sreg[179]), .B(n1349), .Z(n102) );
  XOR U1667 ( .A(n1350), .B(n1351), .Z(n101) );
  XNOR U1668 ( .A(n1352), .B(n1349), .Z(n1351) );
  XOR U1669 ( .A(n1353), .B(n1354), .Z(n1349) );
  ANDN U1670 ( .B(n103), .A(n104), .Z(n1353) );
  XOR U1671 ( .A(sreg[178]), .B(n1354), .Z(n104) );
  XOR U1672 ( .A(n1355), .B(n1356), .Z(n103) );
  XNOR U1673 ( .A(n1357), .B(n1354), .Z(n1356) );
  XOR U1674 ( .A(n1358), .B(n1359), .Z(n1354) );
  ANDN U1675 ( .B(n105), .A(n106), .Z(n1358) );
  XOR U1676 ( .A(sreg[177]), .B(n1359), .Z(n106) );
  XOR U1677 ( .A(n1360), .B(n1361), .Z(n105) );
  XNOR U1678 ( .A(n1362), .B(n1359), .Z(n1361) );
  XOR U1679 ( .A(n1363), .B(n1364), .Z(n1359) );
  ANDN U1680 ( .B(n107), .A(n108), .Z(n1363) );
  XOR U1681 ( .A(sreg[176]), .B(n1364), .Z(n108) );
  XOR U1682 ( .A(n1365), .B(n1366), .Z(n107) );
  XNOR U1683 ( .A(n1367), .B(n1364), .Z(n1366) );
  XOR U1684 ( .A(n1368), .B(n1369), .Z(n1364) );
  ANDN U1685 ( .B(n109), .A(n110), .Z(n1368) );
  XOR U1686 ( .A(sreg[175]), .B(n1369), .Z(n110) );
  XOR U1687 ( .A(n1370), .B(n1371), .Z(n109) );
  XNOR U1688 ( .A(n1372), .B(n1369), .Z(n1371) );
  XOR U1689 ( .A(n1373), .B(n1374), .Z(n1369) );
  ANDN U1690 ( .B(n111), .A(n112), .Z(n1373) );
  XOR U1691 ( .A(sreg[174]), .B(n1374), .Z(n112) );
  XOR U1692 ( .A(n1375), .B(n1376), .Z(n111) );
  XNOR U1693 ( .A(n1377), .B(n1374), .Z(n1376) );
  XOR U1694 ( .A(n1378), .B(n1379), .Z(n1374) );
  ANDN U1695 ( .B(n113), .A(n114), .Z(n1378) );
  XOR U1696 ( .A(sreg[173]), .B(n1379), .Z(n114) );
  XOR U1697 ( .A(n1380), .B(n1381), .Z(n113) );
  XNOR U1698 ( .A(n1382), .B(n1379), .Z(n1381) );
  XOR U1699 ( .A(n1383), .B(n1384), .Z(n1379) );
  ANDN U1700 ( .B(n115), .A(n116), .Z(n1383) );
  XOR U1701 ( .A(sreg[172]), .B(n1384), .Z(n116) );
  XOR U1702 ( .A(n1385), .B(n1386), .Z(n115) );
  XNOR U1703 ( .A(n1387), .B(n1384), .Z(n1386) );
  XOR U1704 ( .A(n1388), .B(n1389), .Z(n1384) );
  ANDN U1705 ( .B(n117), .A(n118), .Z(n1388) );
  XOR U1706 ( .A(sreg[171]), .B(n1389), .Z(n118) );
  XOR U1707 ( .A(n1390), .B(n1391), .Z(n117) );
  XNOR U1708 ( .A(n1392), .B(n1389), .Z(n1391) );
  XOR U1709 ( .A(n1393), .B(n1394), .Z(n1389) );
  ANDN U1710 ( .B(n119), .A(n120), .Z(n1393) );
  XOR U1711 ( .A(sreg[170]), .B(n1394), .Z(n120) );
  XOR U1712 ( .A(n1395), .B(n1396), .Z(n119) );
  XNOR U1713 ( .A(n1397), .B(n1394), .Z(n1396) );
  XOR U1714 ( .A(n1398), .B(n1399), .Z(n1394) );
  ANDN U1715 ( .B(n121), .A(n122), .Z(n1398) );
  XOR U1716 ( .A(sreg[169]), .B(n1399), .Z(n122) );
  XOR U1717 ( .A(n1400), .B(n1401), .Z(n121) );
  XNOR U1718 ( .A(n1402), .B(n1399), .Z(n1401) );
  XOR U1719 ( .A(n1403), .B(n1404), .Z(n1399) );
  ANDN U1720 ( .B(n123), .A(n124), .Z(n1403) );
  XOR U1721 ( .A(sreg[168]), .B(n1404), .Z(n124) );
  XOR U1722 ( .A(n1405), .B(n1406), .Z(n123) );
  XNOR U1723 ( .A(n1407), .B(n1404), .Z(n1406) );
  XOR U1724 ( .A(n1408), .B(n1409), .Z(n1404) );
  ANDN U1725 ( .B(n125), .A(n126), .Z(n1408) );
  XOR U1726 ( .A(sreg[167]), .B(n1409), .Z(n126) );
  XOR U1727 ( .A(n1410), .B(n1411), .Z(n125) );
  XNOR U1728 ( .A(n1412), .B(n1409), .Z(n1411) );
  XOR U1729 ( .A(n1413), .B(n1414), .Z(n1409) );
  ANDN U1730 ( .B(n127), .A(n128), .Z(n1413) );
  XOR U1731 ( .A(sreg[166]), .B(n1414), .Z(n128) );
  XOR U1732 ( .A(n1415), .B(n1416), .Z(n127) );
  XNOR U1733 ( .A(n1417), .B(n1414), .Z(n1416) );
  XOR U1734 ( .A(n1418), .B(n1419), .Z(n1414) );
  ANDN U1735 ( .B(n129), .A(n130), .Z(n1418) );
  XOR U1736 ( .A(sreg[165]), .B(n1419), .Z(n130) );
  XOR U1737 ( .A(n1420), .B(n1421), .Z(n129) );
  XNOR U1738 ( .A(n1422), .B(n1419), .Z(n1421) );
  XOR U1739 ( .A(n1423), .B(n1424), .Z(n1419) );
  ANDN U1740 ( .B(n131), .A(n132), .Z(n1423) );
  XOR U1741 ( .A(sreg[164]), .B(n1424), .Z(n132) );
  XOR U1742 ( .A(n1425), .B(n1426), .Z(n131) );
  XNOR U1743 ( .A(n1427), .B(n1424), .Z(n1426) );
  XOR U1744 ( .A(n1428), .B(n1429), .Z(n1424) );
  ANDN U1745 ( .B(n133), .A(n134), .Z(n1428) );
  XOR U1746 ( .A(sreg[163]), .B(n1429), .Z(n134) );
  XOR U1747 ( .A(n1430), .B(n1431), .Z(n133) );
  XNOR U1748 ( .A(n1432), .B(n1429), .Z(n1431) );
  XOR U1749 ( .A(n1433), .B(n1434), .Z(n1429) );
  ANDN U1750 ( .B(n135), .A(n136), .Z(n1433) );
  XOR U1751 ( .A(sreg[162]), .B(n1434), .Z(n136) );
  XOR U1752 ( .A(n1435), .B(n1436), .Z(n135) );
  XNOR U1753 ( .A(n1437), .B(n1434), .Z(n1436) );
  XOR U1754 ( .A(n1438), .B(n1439), .Z(n1434) );
  ANDN U1755 ( .B(n137), .A(n138), .Z(n1438) );
  XOR U1756 ( .A(sreg[161]), .B(n1439), .Z(n138) );
  XOR U1757 ( .A(n1440), .B(n1441), .Z(n137) );
  XNOR U1758 ( .A(n1442), .B(n1439), .Z(n1441) );
  XOR U1759 ( .A(n1443), .B(n1444), .Z(n1439) );
  ANDN U1760 ( .B(n139), .A(n140), .Z(n1443) );
  XOR U1761 ( .A(sreg[160]), .B(n1444), .Z(n140) );
  XOR U1762 ( .A(n1445), .B(n1446), .Z(n139) );
  XNOR U1763 ( .A(n1447), .B(n1444), .Z(n1446) );
  XOR U1764 ( .A(n1448), .B(n1449), .Z(n1444) );
  ANDN U1765 ( .B(n141), .A(n142), .Z(n1448) );
  XOR U1766 ( .A(sreg[159]), .B(n1449), .Z(n142) );
  XOR U1767 ( .A(n1450), .B(n1451), .Z(n141) );
  XNOR U1768 ( .A(n1452), .B(n1449), .Z(n1451) );
  XOR U1769 ( .A(n1453), .B(n1454), .Z(n1449) );
  ANDN U1770 ( .B(n143), .A(n144), .Z(n1453) );
  XOR U1771 ( .A(sreg[158]), .B(n1454), .Z(n144) );
  XOR U1772 ( .A(n1455), .B(n1456), .Z(n143) );
  XNOR U1773 ( .A(n1457), .B(n1454), .Z(n1456) );
  XOR U1774 ( .A(n1458), .B(n1459), .Z(n1454) );
  ANDN U1775 ( .B(n145), .A(n146), .Z(n1458) );
  XOR U1776 ( .A(sreg[157]), .B(n1459), .Z(n146) );
  XOR U1777 ( .A(n1460), .B(n1461), .Z(n145) );
  XNOR U1778 ( .A(n1462), .B(n1459), .Z(n1461) );
  XOR U1779 ( .A(n1463), .B(n1464), .Z(n1459) );
  ANDN U1780 ( .B(n147), .A(n148), .Z(n1463) );
  XOR U1781 ( .A(sreg[156]), .B(n1464), .Z(n148) );
  XOR U1782 ( .A(n1465), .B(n1466), .Z(n147) );
  XNOR U1783 ( .A(n1467), .B(n1464), .Z(n1466) );
  XOR U1784 ( .A(n1468), .B(n1469), .Z(n1464) );
  ANDN U1785 ( .B(n149), .A(n150), .Z(n1468) );
  XOR U1786 ( .A(sreg[155]), .B(n1469), .Z(n150) );
  XOR U1787 ( .A(n1470), .B(n1471), .Z(n149) );
  XNOR U1788 ( .A(n1472), .B(n1469), .Z(n1471) );
  XOR U1789 ( .A(n1473), .B(n1474), .Z(n1469) );
  ANDN U1790 ( .B(n151), .A(n152), .Z(n1473) );
  XOR U1791 ( .A(sreg[154]), .B(n1474), .Z(n152) );
  XOR U1792 ( .A(n1475), .B(n1476), .Z(n151) );
  XNOR U1793 ( .A(n1477), .B(n1474), .Z(n1476) );
  XOR U1794 ( .A(n1478), .B(n1479), .Z(n1474) );
  ANDN U1795 ( .B(n153), .A(n154), .Z(n1478) );
  XOR U1796 ( .A(sreg[153]), .B(n1479), .Z(n154) );
  XOR U1797 ( .A(n1480), .B(n1481), .Z(n153) );
  XNOR U1798 ( .A(n1482), .B(n1479), .Z(n1481) );
  XOR U1799 ( .A(n1483), .B(n1484), .Z(n1479) );
  ANDN U1800 ( .B(n155), .A(n156), .Z(n1483) );
  XOR U1801 ( .A(sreg[152]), .B(n1484), .Z(n156) );
  XOR U1802 ( .A(n1485), .B(n1486), .Z(n155) );
  XNOR U1803 ( .A(n1487), .B(n1484), .Z(n1486) );
  XOR U1804 ( .A(n1488), .B(n1489), .Z(n1484) );
  ANDN U1805 ( .B(n157), .A(n158), .Z(n1488) );
  XOR U1806 ( .A(sreg[151]), .B(n1489), .Z(n158) );
  XOR U1807 ( .A(n1490), .B(n1491), .Z(n157) );
  XNOR U1808 ( .A(n1492), .B(n1489), .Z(n1491) );
  XOR U1809 ( .A(n1493), .B(n1494), .Z(n1489) );
  ANDN U1810 ( .B(n159), .A(n160), .Z(n1493) );
  XOR U1811 ( .A(sreg[150]), .B(n1494), .Z(n160) );
  XOR U1812 ( .A(n1495), .B(n1496), .Z(n159) );
  XNOR U1813 ( .A(n1497), .B(n1494), .Z(n1496) );
  XOR U1814 ( .A(n1498), .B(n1499), .Z(n1494) );
  ANDN U1815 ( .B(n161), .A(n162), .Z(n1498) );
  XOR U1816 ( .A(sreg[149]), .B(n1499), .Z(n162) );
  XOR U1817 ( .A(n1500), .B(n1501), .Z(n161) );
  XNOR U1818 ( .A(n1502), .B(n1499), .Z(n1501) );
  XOR U1819 ( .A(n1503), .B(n1504), .Z(n1499) );
  ANDN U1820 ( .B(n163), .A(n164), .Z(n1503) );
  XOR U1821 ( .A(sreg[148]), .B(n1504), .Z(n164) );
  XOR U1822 ( .A(n1505), .B(n1506), .Z(n163) );
  XNOR U1823 ( .A(n1507), .B(n1504), .Z(n1506) );
  XOR U1824 ( .A(n1508), .B(n1509), .Z(n1504) );
  ANDN U1825 ( .B(n165), .A(n166), .Z(n1508) );
  XOR U1826 ( .A(sreg[147]), .B(n1509), .Z(n166) );
  XOR U1827 ( .A(n1510), .B(n1511), .Z(n165) );
  XNOR U1828 ( .A(n1512), .B(n1509), .Z(n1511) );
  XOR U1829 ( .A(n1513), .B(n1514), .Z(n1509) );
  ANDN U1830 ( .B(n167), .A(n168), .Z(n1513) );
  XOR U1831 ( .A(sreg[146]), .B(n1514), .Z(n168) );
  XOR U1832 ( .A(n1515), .B(n1516), .Z(n167) );
  XNOR U1833 ( .A(n1517), .B(n1514), .Z(n1516) );
  XOR U1834 ( .A(n1518), .B(n1519), .Z(n1514) );
  ANDN U1835 ( .B(n169), .A(n170), .Z(n1518) );
  XOR U1836 ( .A(sreg[145]), .B(n1519), .Z(n170) );
  XOR U1837 ( .A(n1520), .B(n1521), .Z(n169) );
  XNOR U1838 ( .A(n1522), .B(n1519), .Z(n1521) );
  XOR U1839 ( .A(n1523), .B(n1524), .Z(n1519) );
  ANDN U1840 ( .B(n171), .A(n172), .Z(n1523) );
  XOR U1841 ( .A(sreg[144]), .B(n1524), .Z(n172) );
  XOR U1842 ( .A(n1525), .B(n1526), .Z(n171) );
  XNOR U1843 ( .A(n1527), .B(n1524), .Z(n1526) );
  XOR U1844 ( .A(n1528), .B(n1529), .Z(n1524) );
  ANDN U1845 ( .B(n173), .A(n174), .Z(n1528) );
  XOR U1846 ( .A(sreg[143]), .B(n1529), .Z(n174) );
  XOR U1847 ( .A(n1530), .B(n1531), .Z(n173) );
  XNOR U1848 ( .A(n1532), .B(n1529), .Z(n1531) );
  XOR U1849 ( .A(n1533), .B(n1534), .Z(n1529) );
  ANDN U1850 ( .B(n175), .A(n176), .Z(n1533) );
  XOR U1851 ( .A(sreg[142]), .B(n1534), .Z(n176) );
  XOR U1852 ( .A(n1535), .B(n1536), .Z(n175) );
  XNOR U1853 ( .A(n1537), .B(n1534), .Z(n1536) );
  XOR U1854 ( .A(n1538), .B(n1539), .Z(n1534) );
  ANDN U1855 ( .B(n177), .A(n178), .Z(n1538) );
  XOR U1856 ( .A(sreg[141]), .B(n1539), .Z(n178) );
  XOR U1857 ( .A(n1540), .B(n1541), .Z(n177) );
  XNOR U1858 ( .A(n1542), .B(n1539), .Z(n1541) );
  XOR U1859 ( .A(n1543), .B(n1544), .Z(n1539) );
  ANDN U1860 ( .B(n179), .A(n180), .Z(n1543) );
  XOR U1861 ( .A(sreg[140]), .B(n1544), .Z(n180) );
  XOR U1862 ( .A(n1545), .B(n1546), .Z(n179) );
  XNOR U1863 ( .A(n1547), .B(n1544), .Z(n1546) );
  XOR U1864 ( .A(n1548), .B(n1549), .Z(n1544) );
  ANDN U1865 ( .B(n426), .A(n427), .Z(n1548) );
  XOR U1866 ( .A(sreg[139]), .B(n1549), .Z(n427) );
  XOR U1867 ( .A(n1550), .B(n1551), .Z(n426) );
  XNOR U1868 ( .A(n1552), .B(n1549), .Z(n1551) );
  XOR U1869 ( .A(n1553), .B(n1554), .Z(n1549) );
  ANDN U1870 ( .B(n768), .A(n769), .Z(n1553) );
  XOR U1871 ( .A(sreg[138]), .B(n1554), .Z(n769) );
  XOR U1872 ( .A(n1555), .B(n1556), .Z(n768) );
  XNOR U1873 ( .A(n1557), .B(n1554), .Z(n1556) );
  XOR U1874 ( .A(n1558), .B(n1559), .Z(n1554) );
  ANDN U1875 ( .B(n2), .A(n1), .Z(n1558) );
  XOR U1876 ( .A(sreg[137]), .B(n1559), .Z(n1) );
  XOR U1877 ( .A(n1560), .B(n1561), .Z(n2) );
  XNOR U1878 ( .A(n1562), .B(n1559), .Z(n1561) );
  XOR U1879 ( .A(n1563), .B(n1564), .Z(n1559) );
  ANDN U1880 ( .B(n23), .A(n24), .Z(n1563) );
  XOR U1881 ( .A(sreg[136]), .B(n1564), .Z(n24) );
  XOR U1882 ( .A(n1565), .B(n1566), .Z(n23) );
  XNOR U1883 ( .A(n1567), .B(n1564), .Z(n1566) );
  XOR U1884 ( .A(n1568), .B(n1569), .Z(n1564) );
  ANDN U1885 ( .B(n1570), .A(n1571), .Z(n1568) );
  NANDN U1886 ( .A(n187), .B(a[100]), .Z(n1077) );
  XNOR U1887 ( .A(n1100), .B(n1101), .Z(n1078) );
  XOR U1888 ( .A(n1098), .B(n1572), .Z(n1101) );
  NAND U1889 ( .A(b[1]), .B(a[99]), .Z(n1572) );
  XOR U1890 ( .A(n1106), .B(n1573), .Z(n1100) );
  XOR U1891 ( .A(n1098), .B(n1105), .Z(n1573) );
  XNOR U1892 ( .A(n1574), .B(n1104), .Z(n1105) );
  AND U1893 ( .A(b[2]), .B(a[98]), .Z(n1574) );
  OR U1894 ( .A(n1112), .B(n1110), .Z(n1098) );
  XOR U1895 ( .A(n1575), .B(n1576), .Z(n1110) );
  NANDN U1896 ( .A(n187), .B(a[99]), .Z(n1112) );
  XOR U1897 ( .A(n1104), .B(n1096), .Z(n1577) );
  XOR U1898 ( .A(n1095), .B(n1092), .Z(n1578) );
  XOR U1899 ( .A(n1579), .B(n1580), .Z(n1092) );
  XOR U1900 ( .A(n1090), .B(n1581), .Z(n1580) );
  XNOR U1901 ( .A(n1582), .B(n1583), .Z(n1581) );
  XOR U1902 ( .A(n1584), .B(n1585), .Z(n1583) );
  NAND U1903 ( .A(b[6]), .B(a[94]), .Z(n1585) );
  AND U1904 ( .A(b[7]), .B(a[93]), .Z(n1584) );
  XNOR U1905 ( .A(n1586), .B(n1582), .Z(n1579) );
  XOR U1906 ( .A(n1587), .B(n1588), .Z(n1582) );
  NOR U1907 ( .A(n1589), .B(n1590), .Z(n1587) );
  AND U1908 ( .A(b[5]), .B(a[95]), .Z(n1586) );
  XNOR U1909 ( .A(n1591), .B(n1090), .Z(n1091) );
  XNOR U1910 ( .A(n1592), .B(n1593), .Z(n1090) );
  ANDN U1911 ( .B(n1594), .A(n1595), .Z(n1592) );
  AND U1912 ( .A(b[4]), .B(a[96]), .Z(n1591) );
  XNOR U1913 ( .A(n1596), .B(n1597), .Z(n1104) );
  NANDN U1914 ( .A(n1576), .B(n1575), .Z(n1597) );
  XOR U1915 ( .A(n1596), .B(n1598), .Z(n1575) );
  NAND U1916 ( .A(b[1]), .B(a[98]), .Z(n1598) );
  XOR U1917 ( .A(n1596), .B(n1600), .Z(n1599) );
  OR U1918 ( .A(n1117), .B(n1115), .Z(n1596) );
  XOR U1919 ( .A(n1602), .B(n1603), .Z(n1115) );
  NANDN U1920 ( .A(n187), .B(a[98]), .Z(n1117) );
  XNOR U1921 ( .A(n1604), .B(n1095), .Z(n1097) );
  XNOR U1922 ( .A(n1605), .B(n1606), .Z(n1095) );
  ANDN U1923 ( .B(n1600), .A(n1601), .Z(n1605) );
  XOR U1924 ( .A(n1607), .B(n1606), .Z(n1601) );
  IV U1925 ( .A(n1608), .Z(n1606) );
  AND U1926 ( .A(b[2]), .B(a[97]), .Z(n1607) );
  XNOR U1927 ( .A(n1594), .B(n1608), .Z(n1609) );
  XOR U1928 ( .A(n1610), .B(n1611), .Z(n1608) );
  NANDN U1929 ( .A(n1603), .B(n1602), .Z(n1611) );
  XOR U1930 ( .A(n1610), .B(n1612), .Z(n1602) );
  NAND U1931 ( .A(b[1]), .B(a[97]), .Z(n1612) );
  XOR U1932 ( .A(n1610), .B(n1614), .Z(n1613) );
  OR U1933 ( .A(n1122), .B(n1120), .Z(n1610) );
  XOR U1934 ( .A(n1616), .B(n1617), .Z(n1120) );
  NANDN U1935 ( .A(n187), .B(a[97]), .Z(n1122) );
  XOR U1936 ( .A(n1590), .B(n1619), .Z(n1618) );
  XOR U1937 ( .A(n1620), .B(n1621), .Z(n1590) );
  XNOR U1938 ( .A(n1622), .B(n1623), .Z(n1621) );
  XNOR U1939 ( .A(n1624), .B(n1625), .Z(n1622) );
  XOR U1940 ( .A(n1626), .B(n1627), .Z(n1625) );
  AND U1941 ( .A(b[7]), .B(a[92]), .Z(n1627) );
  AND U1942 ( .A(b[6]), .B(a[93]), .Z(n1626) );
  XNOR U1943 ( .A(n1628), .B(n1624), .Z(n1620) );
  XOR U1944 ( .A(n1629), .B(n1630), .Z(n1624) );
  NOR U1945 ( .A(n1631), .B(n1632), .Z(n1629) );
  AND U1946 ( .A(b[5]), .B(a[94]), .Z(n1628) );
  XOR U1947 ( .A(n1633), .B(n1588), .Z(n1589) );
  IV U1948 ( .A(n1623), .Z(n1588) );
  XOR U1949 ( .A(n1634), .B(n1635), .Z(n1623) );
  ANDN U1950 ( .B(n1636), .A(n1637), .Z(n1634) );
  AND U1951 ( .A(b[4]), .B(a[95]), .Z(n1633) );
  XOR U1952 ( .A(n1638), .B(n1593), .Z(n1595) );
  IV U1953 ( .A(n1619), .Z(n1593) );
  XOR U1954 ( .A(n1639), .B(n1640), .Z(n1619) );
  ANDN U1955 ( .B(n1614), .A(n1615), .Z(n1639) );
  AND U1956 ( .A(b[2]), .B(a[96]), .Z(n1641) );
  XNOR U1957 ( .A(n1636), .B(n1640), .Z(n1642) );
  XOR U1958 ( .A(n1643), .B(n1644), .Z(n1640) );
  NANDN U1959 ( .A(n1617), .B(n1616), .Z(n1644) );
  XOR U1960 ( .A(n1643), .B(n1645), .Z(n1616) );
  NAND U1961 ( .A(b[1]), .B(a[96]), .Z(n1645) );
  XOR U1962 ( .A(n1643), .B(n1647), .Z(n1646) );
  OR U1963 ( .A(n1127), .B(n1125), .Z(n1643) );
  XOR U1964 ( .A(n1649), .B(n1650), .Z(n1125) );
  NANDN U1965 ( .A(n187), .B(a[96]), .Z(n1127) );
  XOR U1966 ( .A(n1632), .B(n1635), .Z(n1651) );
  XOR U1967 ( .A(n1652), .B(n1653), .Z(n1632) );
  XNOR U1968 ( .A(n1654), .B(n1655), .Z(n1653) );
  XNOR U1969 ( .A(n1656), .B(n1657), .Z(n1654) );
  XOR U1970 ( .A(n1658), .B(n1659), .Z(n1657) );
  AND U1971 ( .A(b[6]), .B(a[92]), .Z(n1659) );
  AND U1972 ( .A(b[7]), .B(a[91]), .Z(n1658) );
  XNOR U1973 ( .A(n1660), .B(n1656), .Z(n1652) );
  XOR U1974 ( .A(n1661), .B(n1662), .Z(n1656) );
  NOR U1975 ( .A(n1663), .B(n1664), .Z(n1661) );
  AND U1976 ( .A(b[5]), .B(a[93]), .Z(n1660) );
  XOR U1977 ( .A(n1665), .B(n1630), .Z(n1631) );
  IV U1978 ( .A(n1655), .Z(n1630) );
  XOR U1979 ( .A(n1666), .B(n1667), .Z(n1655) );
  ANDN U1980 ( .B(n1668), .A(n1669), .Z(n1666) );
  AND U1981 ( .A(b[4]), .B(a[94]), .Z(n1665) );
  XOR U1982 ( .A(n1671), .B(n1672), .Z(n1635) );
  ANDN U1983 ( .B(n1647), .A(n1648), .Z(n1671) );
  AND U1984 ( .A(b[2]), .B(a[95]), .Z(n1673) );
  XNOR U1985 ( .A(n1668), .B(n1672), .Z(n1674) );
  XOR U1986 ( .A(n1675), .B(n1676), .Z(n1672) );
  NANDN U1987 ( .A(n1650), .B(n1649), .Z(n1676) );
  XOR U1988 ( .A(n1675), .B(n1677), .Z(n1649) );
  NAND U1989 ( .A(b[1]), .B(a[95]), .Z(n1677) );
  XOR U1990 ( .A(n1675), .B(n1679), .Z(n1678) );
  OR U1991 ( .A(n1132), .B(n1130), .Z(n1675) );
  XOR U1992 ( .A(n1681), .B(n1682), .Z(n1130) );
  NANDN U1993 ( .A(n187), .B(a[95]), .Z(n1132) );
  XOR U1994 ( .A(n1664), .B(n1667), .Z(n1683) );
  XOR U1995 ( .A(n1684), .B(n1685), .Z(n1664) );
  XNOR U1996 ( .A(n1686), .B(n1687), .Z(n1685) );
  XOR U1997 ( .A(n1688), .B(n1689), .Z(n1686) );
  AND U1998 ( .A(b[5]), .B(a[92]), .Z(n1688) );
  XOR U1999 ( .A(n1689), .B(n1690), .Z(n1684) );
  XOR U2000 ( .A(n1691), .B(n1692), .Z(n1690) );
  AND U2001 ( .A(b[6]), .B(a[91]), .Z(n1692) );
  AND U2002 ( .A(b[7]), .B(a[90]), .Z(n1691) );
  XOR U2003 ( .A(n1693), .B(n1694), .Z(n1689) );
  ANDN U2004 ( .B(n1695), .A(n1696), .Z(n1693) );
  XOR U2005 ( .A(n1697), .B(n1662), .Z(n1663) );
  IV U2006 ( .A(n1687), .Z(n1662) );
  XOR U2007 ( .A(n1698), .B(n1699), .Z(n1687) );
  NOR U2008 ( .A(n1700), .B(n1701), .Z(n1698) );
  AND U2009 ( .A(b[4]), .B(a[93]), .Z(n1697) );
  XOR U2010 ( .A(n1703), .B(n1704), .Z(n1667) );
  ANDN U2011 ( .B(n1679), .A(n1680), .Z(n1703) );
  AND U2012 ( .A(b[2]), .B(a[94]), .Z(n1705) );
  XOR U2013 ( .A(n1701), .B(n1704), .Z(n1706) );
  XOR U2014 ( .A(n1707), .B(n1708), .Z(n1704) );
  NANDN U2015 ( .A(n1682), .B(n1681), .Z(n1708) );
  XOR U2016 ( .A(n1707), .B(n1709), .Z(n1681) );
  NAND U2017 ( .A(b[1]), .B(a[94]), .Z(n1709) );
  XOR U2018 ( .A(n1707), .B(n1711), .Z(n1710) );
  OR U2019 ( .A(n1137), .B(n1135), .Z(n1707) );
  XOR U2020 ( .A(n1713), .B(n1714), .Z(n1135) );
  NANDN U2021 ( .A(n187), .B(a[94]), .Z(n1137) );
  XNOR U2022 ( .A(n1696), .B(n1715), .Z(n1701) );
  XNOR U2023 ( .A(n1695), .B(n1699), .Z(n1715) );
  XOR U2024 ( .A(n1716), .B(n1694), .Z(n1695) );
  AND U2025 ( .A(b[4]), .B(a[92]), .Z(n1716) );
  XOR U2026 ( .A(n1717), .B(n1718), .Z(n1696) );
  XOR U2027 ( .A(n1694), .B(n1719), .Z(n1718) );
  XOR U2028 ( .A(n1720), .B(n1721), .Z(n1719) );
  XOR U2029 ( .A(n1722), .B(n1723), .Z(n1721) );
  NAND U2030 ( .A(b[6]), .B(a[90]), .Z(n1723) );
  AND U2031 ( .A(b[7]), .B(a[89]), .Z(n1722) );
  XOR U2032 ( .A(n1724), .B(n1725), .Z(n1694) );
  ANDN U2033 ( .B(n1726), .A(n1727), .Z(n1724) );
  XOR U2034 ( .A(n1728), .B(n1720), .Z(n1717) );
  XOR U2035 ( .A(n1729), .B(n1730), .Z(n1720) );
  NOR U2036 ( .A(n1731), .B(n1732), .Z(n1729) );
  AND U2037 ( .A(b[5]), .B(a[91]), .Z(n1728) );
  XOR U2038 ( .A(n1734), .B(n1735), .Z(n1699) );
  ANDN U2039 ( .B(n1711), .A(n1712), .Z(n1734) );
  AND U2040 ( .A(b[2]), .B(a[93]), .Z(n1736) );
  XNOR U2041 ( .A(n1726), .B(n1735), .Z(n1737) );
  XOR U2042 ( .A(n1738), .B(n1739), .Z(n1735) );
  NANDN U2043 ( .A(n1714), .B(n1713), .Z(n1739) );
  XOR U2044 ( .A(n1738), .B(n1740), .Z(n1713) );
  NAND U2045 ( .A(b[1]), .B(a[93]), .Z(n1740) );
  XNOR U2046 ( .A(n1738), .B(n1742), .Z(n1741) );
  OR U2047 ( .A(n1142), .B(n1140), .Z(n1738) );
  NANDN U2048 ( .A(n187), .B(a[93]), .Z(n1142) );
  XOR U2049 ( .A(n1746), .B(n1725), .Z(n1726) );
  AND U2050 ( .A(b[3]), .B(a[92]), .Z(n1746) );
  XOR U2051 ( .A(n1725), .B(n1732), .Z(n1747) );
  XOR U2052 ( .A(n1748), .B(n1749), .Z(n1732) );
  XOR U2053 ( .A(n1730), .B(n1750), .Z(n1749) );
  XOR U2054 ( .A(n1751), .B(n1752), .Z(n1750) );
  XOR U2055 ( .A(n1753), .B(n1754), .Z(n1752) );
  NAND U2056 ( .A(b[6]), .B(a[89]), .Z(n1754) );
  AND U2057 ( .A(b[7]), .B(a[88]), .Z(n1753) );
  XOR U2058 ( .A(n1755), .B(n1751), .Z(n1748) );
  XOR U2059 ( .A(n1756), .B(n1757), .Z(n1751) );
  NOR U2060 ( .A(n1758), .B(n1759), .Z(n1756) );
  AND U2061 ( .A(b[5]), .B(a[90]), .Z(n1755) );
  XNOR U2062 ( .A(n1760), .B(n1761), .Z(n1725) );
  NOR U2063 ( .A(n1743), .B(n1742), .Z(n1760) );
  XOR U2064 ( .A(n1762), .B(n1761), .Z(n1742) );
  AND U2065 ( .A(b[2]), .B(a[92]), .Z(n1762) );
  XOR U2066 ( .A(n1761), .B(n1764), .Z(n1763) );
  XNOR U2067 ( .A(n1765), .B(n1766), .Z(n1761) );
  OR U2068 ( .A(n1744), .B(n1745), .Z(n1766) );
  XNOR U2069 ( .A(n1765), .B(n1768), .Z(n1767) );
  XNOR U2070 ( .A(n1765), .B(n1770), .Z(n1744) );
  NAND U2071 ( .A(b[1]), .B(a[92]), .Z(n1770) );
  OR U2072 ( .A(n1147), .B(n1145), .Z(n1765) );
  XOR U2073 ( .A(n1771), .B(n1772), .Z(n1145) );
  NANDN U2074 ( .A(n187), .B(a[92]), .Z(n1147) );
  XNOR U2075 ( .A(n1774), .B(n1730), .Z(n1731) );
  XOR U2076 ( .A(n1775), .B(n1776), .Z(n1730) );
  ANDN U2077 ( .B(n1764), .A(n1773), .Z(n1775) );
  XNOR U2078 ( .A(n1777), .B(n1776), .Z(n1773) );
  AND U2079 ( .A(b[3]), .B(a[91]), .Z(n1777) );
  XOR U2080 ( .A(n1776), .B(n1759), .Z(n1778) );
  XOR U2081 ( .A(n1779), .B(n1780), .Z(n1759) );
  XOR U2082 ( .A(n1757), .B(n1781), .Z(n1780) );
  XOR U2083 ( .A(n1782), .B(n1783), .Z(n1781) );
  XOR U2084 ( .A(n1784), .B(n1785), .Z(n1783) );
  NAND U2085 ( .A(b[6]), .B(a[88]), .Z(n1785) );
  AND U2086 ( .A(b[7]), .B(a[87]), .Z(n1784) );
  XOR U2087 ( .A(n1786), .B(n1782), .Z(n1779) );
  XOR U2088 ( .A(n1787), .B(n1788), .Z(n1782) );
  NOR U2089 ( .A(n1789), .B(n1790), .Z(n1787) );
  AND U2090 ( .A(b[5]), .B(a[89]), .Z(n1786) );
  XNOR U2091 ( .A(n1791), .B(n1792), .Z(n1776) );
  NOR U2092 ( .A(n1769), .B(n1768), .Z(n1791) );
  XOR U2093 ( .A(n1793), .B(n1792), .Z(n1768) );
  AND U2094 ( .A(b[2]), .B(a[91]), .Z(n1793) );
  XOR U2095 ( .A(n1792), .B(n1795), .Z(n1794) );
  XNOR U2096 ( .A(n1796), .B(n1797), .Z(n1792) );
  NANDN U2097 ( .A(n1772), .B(n1771), .Z(n1797) );
  XOR U2098 ( .A(n1796), .B(n1798), .Z(n1771) );
  NAND U2099 ( .A(b[1]), .B(a[91]), .Z(n1798) );
  XOR U2100 ( .A(n1796), .B(n1800), .Z(n1799) );
  OR U2101 ( .A(n1152), .B(n1150), .Z(n1796) );
  XOR U2102 ( .A(n1802), .B(n1803), .Z(n1150) );
  NANDN U2103 ( .A(n187), .B(a[91]), .Z(n1152) );
  XNOR U2104 ( .A(n1805), .B(n1757), .Z(n1758) );
  XOR U2105 ( .A(n1806), .B(n1807), .Z(n1757) );
  ANDN U2106 ( .B(n1795), .A(n1804), .Z(n1806) );
  XNOR U2107 ( .A(n1808), .B(n1807), .Z(n1804) );
  AND U2108 ( .A(b[3]), .B(a[90]), .Z(n1808) );
  XOR U2109 ( .A(n1807), .B(n1790), .Z(n1809) );
  XOR U2110 ( .A(n1810), .B(n1811), .Z(n1790) );
  XOR U2111 ( .A(n1788), .B(n1812), .Z(n1811) );
  XNOR U2112 ( .A(n1813), .B(n1814), .Z(n1812) );
  XOR U2113 ( .A(n1815), .B(n1816), .Z(n1814) );
  NAND U2114 ( .A(b[6]), .B(a[87]), .Z(n1816) );
  AND U2115 ( .A(b[7]), .B(a[86]), .Z(n1815) );
  XNOR U2116 ( .A(n1817), .B(n1813), .Z(n1810) );
  XOR U2117 ( .A(n1818), .B(n1819), .Z(n1813) );
  NOR U2118 ( .A(n1820), .B(n1821), .Z(n1818) );
  AND U2119 ( .A(b[5]), .B(a[88]), .Z(n1817) );
  XNOR U2120 ( .A(n1822), .B(n1823), .Z(n1807) );
  ANDN U2121 ( .B(n1800), .A(n1801), .Z(n1822) );
  XOR U2122 ( .A(n1824), .B(n1823), .Z(n1801) );
  IV U2123 ( .A(n1825), .Z(n1823) );
  AND U2124 ( .A(b[2]), .B(a[90]), .Z(n1824) );
  XNOR U2125 ( .A(n1827), .B(n1825), .Z(n1826) );
  XOR U2126 ( .A(n1828), .B(n1829), .Z(n1825) );
  NANDN U2127 ( .A(n1803), .B(n1802), .Z(n1829) );
  XOR U2128 ( .A(n1828), .B(n1830), .Z(n1802) );
  NAND U2129 ( .A(b[1]), .B(a[90]), .Z(n1830) );
  XOR U2130 ( .A(n1828), .B(n1832), .Z(n1831) );
  OR U2131 ( .A(n1157), .B(n1155), .Z(n1828) );
  XOR U2132 ( .A(n1834), .B(n1835), .Z(n1155) );
  NANDN U2133 ( .A(n187), .B(a[90]), .Z(n1157) );
  XNOR U2134 ( .A(n1837), .B(n1788), .Z(n1789) );
  XNOR U2135 ( .A(n1838), .B(n1839), .Z(n1788) );
  ANDN U2136 ( .B(n1827), .A(n1836), .Z(n1838) );
  XOR U2137 ( .A(n1840), .B(n1839), .Z(n1836) );
  IV U2138 ( .A(n1841), .Z(n1839) );
  AND U2139 ( .A(b[3]), .B(a[89]), .Z(n1840) );
  XOR U2140 ( .A(n1821), .B(n1841), .Z(n1842) );
  XOR U2141 ( .A(n1843), .B(n1844), .Z(n1841) );
  ANDN U2142 ( .B(n1832), .A(n1833), .Z(n1843) );
  AND U2143 ( .A(b[2]), .B(a[89]), .Z(n1845) );
  XNOR U2144 ( .A(n1847), .B(n1844), .Z(n1846) );
  XOR U2145 ( .A(n1848), .B(n1849), .Z(n1844) );
  NANDN U2146 ( .A(n1835), .B(n1834), .Z(n1849) );
  XOR U2147 ( .A(n1848), .B(n1850), .Z(n1834) );
  NAND U2148 ( .A(b[1]), .B(a[89]), .Z(n1850) );
  XOR U2149 ( .A(n1848), .B(n1852), .Z(n1851) );
  OR U2150 ( .A(n1162), .B(n1160), .Z(n1848) );
  XOR U2151 ( .A(n1854), .B(n1855), .Z(n1160) );
  NANDN U2152 ( .A(n187), .B(a[89]), .Z(n1162) );
  XOR U2153 ( .A(n1857), .B(n1858), .Z(n1821) );
  XNOR U2154 ( .A(n1859), .B(n1860), .Z(n1858) );
  XNOR U2155 ( .A(n1861), .B(n1862), .Z(n1859) );
  XOR U2156 ( .A(n1863), .B(n1864), .Z(n1862) );
  AND U2157 ( .A(b[7]), .B(a[85]), .Z(n1864) );
  AND U2158 ( .A(b[6]), .B(a[86]), .Z(n1863) );
  XNOR U2159 ( .A(n1865), .B(n1861), .Z(n1857) );
  XOR U2160 ( .A(n1866), .B(n1867), .Z(n1861) );
  NOR U2161 ( .A(n1868), .B(n1869), .Z(n1866) );
  AND U2162 ( .A(b[5]), .B(a[87]), .Z(n1865) );
  XOR U2163 ( .A(n1870), .B(n1819), .Z(n1820) );
  IV U2164 ( .A(n1860), .Z(n1819) );
  XOR U2165 ( .A(n1871), .B(n1872), .Z(n1860) );
  ANDN U2166 ( .B(n1847), .A(n1856), .Z(n1871) );
  AND U2167 ( .A(b[3]), .B(a[88]), .Z(n1873) );
  XOR U2168 ( .A(n1869), .B(n1872), .Z(n1874) );
  XOR U2169 ( .A(n1875), .B(n1876), .Z(n1872) );
  ANDN U2170 ( .B(n1852), .A(n1853), .Z(n1875) );
  AND U2171 ( .A(b[2]), .B(a[88]), .Z(n1877) );
  XNOR U2172 ( .A(n1879), .B(n1876), .Z(n1878) );
  XOR U2173 ( .A(n1880), .B(n1881), .Z(n1876) );
  NANDN U2174 ( .A(n1855), .B(n1854), .Z(n1881) );
  XOR U2175 ( .A(n1880), .B(n1882), .Z(n1854) );
  NAND U2176 ( .A(b[1]), .B(a[88]), .Z(n1882) );
  XOR U2177 ( .A(n1880), .B(n1884), .Z(n1883) );
  OR U2178 ( .A(n1167), .B(n1165), .Z(n1880) );
  XOR U2179 ( .A(n1886), .B(n1887), .Z(n1165) );
  NANDN U2180 ( .A(n187), .B(a[88]), .Z(n1167) );
  XOR U2181 ( .A(n1889), .B(n1890), .Z(n1869) );
  XNOR U2182 ( .A(n1891), .B(n1892), .Z(n1890) );
  XNOR U2183 ( .A(n1893), .B(n1894), .Z(n1891) );
  XOR U2184 ( .A(n1895), .B(n1896), .Z(n1894) );
  AND U2185 ( .A(b[6]), .B(a[85]), .Z(n1896) );
  AND U2186 ( .A(b[7]), .B(a[84]), .Z(n1895) );
  XNOR U2187 ( .A(n1897), .B(n1893), .Z(n1889) );
  XOR U2188 ( .A(n1898), .B(n1899), .Z(n1893) );
  NOR U2189 ( .A(n1900), .B(n1901), .Z(n1898) );
  AND U2190 ( .A(b[5]), .B(a[86]), .Z(n1897) );
  XOR U2191 ( .A(n1902), .B(n1867), .Z(n1868) );
  IV U2192 ( .A(n1892), .Z(n1867) );
  XOR U2193 ( .A(n1903), .B(n1904), .Z(n1892) );
  ANDN U2194 ( .B(n1879), .A(n1888), .Z(n1903) );
  AND U2195 ( .A(b[3]), .B(a[87]), .Z(n1905) );
  XOR U2196 ( .A(n1901), .B(n1904), .Z(n1906) );
  XOR U2197 ( .A(n1907), .B(n1908), .Z(n1904) );
  ANDN U2198 ( .B(n1884), .A(n1885), .Z(n1907) );
  AND U2199 ( .A(b[2]), .B(a[87]), .Z(n1909) );
  XOR U2200 ( .A(n1911), .B(n1908), .Z(n1910) );
  XOR U2201 ( .A(n1912), .B(n1913), .Z(n1908) );
  NANDN U2202 ( .A(n1887), .B(n1886), .Z(n1913) );
  XOR U2203 ( .A(n1912), .B(n1914), .Z(n1886) );
  NAND U2204 ( .A(b[1]), .B(a[87]), .Z(n1914) );
  XOR U2205 ( .A(n1912), .B(n1916), .Z(n1915) );
  OR U2206 ( .A(n1172), .B(n1170), .Z(n1912) );
  XOR U2207 ( .A(n1918), .B(n1919), .Z(n1170) );
  NANDN U2208 ( .A(n187), .B(a[87]), .Z(n1172) );
  XOR U2209 ( .A(n1921), .B(n1922), .Z(n1901) );
  XNOR U2210 ( .A(n1923), .B(n1924), .Z(n1922) );
  XOR U2211 ( .A(n1925), .B(n1926), .Z(n1923) );
  AND U2212 ( .A(b[5]), .B(a[85]), .Z(n1925) );
  XOR U2213 ( .A(n1926), .B(n1927), .Z(n1921) );
  XOR U2214 ( .A(n1928), .B(n1929), .Z(n1927) );
  AND U2215 ( .A(b[6]), .B(a[84]), .Z(n1929) );
  AND U2216 ( .A(b[7]), .B(a[83]), .Z(n1928) );
  XOR U2217 ( .A(n1930), .B(n1931), .Z(n1926) );
  ANDN U2218 ( .B(n1932), .A(n1933), .Z(n1930) );
  XOR U2219 ( .A(n1934), .B(n1899), .Z(n1900) );
  IV U2220 ( .A(n1924), .Z(n1899) );
  XOR U2221 ( .A(n1935), .B(n1936), .Z(n1924) );
  NOR U2222 ( .A(n1920), .B(n1911), .Z(n1935) );
  XNOR U2223 ( .A(n1933), .B(n1937), .Z(n1911) );
  XNOR U2224 ( .A(n1932), .B(n1936), .Z(n1937) );
  XOR U2225 ( .A(n1938), .B(n1931), .Z(n1932) );
  AND U2226 ( .A(b[4]), .B(a[85]), .Z(n1938) );
  XOR U2227 ( .A(n1939), .B(n1940), .Z(n1933) );
  XOR U2228 ( .A(n1931), .B(n1941), .Z(n1940) );
  XOR U2229 ( .A(n1942), .B(n1943), .Z(n1941) );
  XOR U2230 ( .A(n1944), .B(n1945), .Z(n1943) );
  NAND U2231 ( .A(b[6]), .B(a[83]), .Z(n1945) );
  AND U2232 ( .A(b[7]), .B(a[82]), .Z(n1944) );
  XOR U2233 ( .A(n1946), .B(n1947), .Z(n1931) );
  ANDN U2234 ( .B(n1948), .A(n1949), .Z(n1946) );
  XOR U2235 ( .A(n1950), .B(n1942), .Z(n1939) );
  XOR U2236 ( .A(n1951), .B(n1952), .Z(n1942) );
  NOR U2237 ( .A(n1953), .B(n1954), .Z(n1951) );
  AND U2238 ( .A(b[5]), .B(a[84]), .Z(n1950) );
  XOR U2239 ( .A(n1956), .B(n1957), .Z(n1936) );
  ANDN U2240 ( .B(n1916), .A(n1917), .Z(n1956) );
  AND U2241 ( .A(b[2]), .B(a[86]), .Z(n1958) );
  XNOR U2242 ( .A(n1948), .B(n1957), .Z(n1959) );
  XOR U2243 ( .A(n1960), .B(n1961), .Z(n1957) );
  NANDN U2244 ( .A(n1919), .B(n1918), .Z(n1961) );
  XOR U2245 ( .A(n1960), .B(n1962), .Z(n1918) );
  NAND U2246 ( .A(b[1]), .B(a[86]), .Z(n1962) );
  XNOR U2247 ( .A(n1960), .B(n1964), .Z(n1963) );
  OR U2248 ( .A(n1177), .B(n1175), .Z(n1960) );
  NANDN U2249 ( .A(n187), .B(a[86]), .Z(n1177) );
  XOR U2250 ( .A(n1968), .B(n1947), .Z(n1948) );
  AND U2251 ( .A(b[3]), .B(a[85]), .Z(n1968) );
  XOR U2252 ( .A(n1947), .B(n1954), .Z(n1969) );
  XOR U2253 ( .A(n1970), .B(n1971), .Z(n1954) );
  XOR U2254 ( .A(n1952), .B(n1972), .Z(n1971) );
  XOR U2255 ( .A(n1973), .B(n1974), .Z(n1972) );
  XOR U2256 ( .A(n1975), .B(n1976), .Z(n1974) );
  NAND U2257 ( .A(b[6]), .B(a[82]), .Z(n1976) );
  AND U2258 ( .A(b[7]), .B(a[81]), .Z(n1975) );
  XOR U2259 ( .A(n1977), .B(n1973), .Z(n1970) );
  XOR U2260 ( .A(n1978), .B(n1979), .Z(n1973) );
  NOR U2261 ( .A(n1980), .B(n1981), .Z(n1978) );
  AND U2262 ( .A(b[5]), .B(a[83]), .Z(n1977) );
  XNOR U2263 ( .A(n1982), .B(n1983), .Z(n1947) );
  NOR U2264 ( .A(n1965), .B(n1964), .Z(n1982) );
  XOR U2265 ( .A(n1984), .B(n1983), .Z(n1964) );
  AND U2266 ( .A(b[2]), .B(a[85]), .Z(n1984) );
  XOR U2267 ( .A(n1983), .B(n1986), .Z(n1985) );
  XNOR U2268 ( .A(n1987), .B(n1988), .Z(n1983) );
  OR U2269 ( .A(n1966), .B(n1967), .Z(n1988) );
  XNOR U2270 ( .A(n1987), .B(n1990), .Z(n1989) );
  XNOR U2271 ( .A(n1987), .B(n1992), .Z(n1966) );
  NAND U2272 ( .A(b[1]), .B(a[85]), .Z(n1992) );
  OR U2273 ( .A(n1182), .B(n1180), .Z(n1987) );
  XOR U2274 ( .A(n1993), .B(n1994), .Z(n1180) );
  NANDN U2275 ( .A(n187), .B(a[85]), .Z(n1182) );
  XNOR U2276 ( .A(n1996), .B(n1952), .Z(n1953) );
  XOR U2277 ( .A(n1997), .B(n1998), .Z(n1952) );
  ANDN U2278 ( .B(n1986), .A(n1995), .Z(n1997) );
  XNOR U2279 ( .A(n1999), .B(n1998), .Z(n1995) );
  AND U2280 ( .A(b[3]), .B(a[84]), .Z(n1999) );
  XOR U2281 ( .A(n1998), .B(n1981), .Z(n2000) );
  XOR U2282 ( .A(n2001), .B(n2002), .Z(n1981) );
  XOR U2283 ( .A(n1979), .B(n2003), .Z(n2002) );
  XOR U2284 ( .A(n2004), .B(n2005), .Z(n2003) );
  XOR U2285 ( .A(n2006), .B(n2007), .Z(n2005) );
  NAND U2286 ( .A(b[6]), .B(a[81]), .Z(n2007) );
  AND U2287 ( .A(b[7]), .B(a[80]), .Z(n2006) );
  XOR U2288 ( .A(n2008), .B(n2004), .Z(n2001) );
  XOR U2289 ( .A(n2009), .B(n2010), .Z(n2004) );
  NOR U2290 ( .A(n2011), .B(n2012), .Z(n2009) );
  AND U2291 ( .A(b[5]), .B(a[82]), .Z(n2008) );
  XNOR U2292 ( .A(n2013), .B(n2014), .Z(n1998) );
  NOR U2293 ( .A(n1991), .B(n1990), .Z(n2013) );
  XOR U2294 ( .A(n2015), .B(n2014), .Z(n1990) );
  AND U2295 ( .A(b[2]), .B(a[84]), .Z(n2015) );
  XOR U2296 ( .A(n2014), .B(n2017), .Z(n2016) );
  XNOR U2297 ( .A(n2018), .B(n2019), .Z(n2014) );
  NANDN U2298 ( .A(n1994), .B(n1993), .Z(n2019) );
  XOR U2299 ( .A(n2018), .B(n2020), .Z(n1993) );
  NAND U2300 ( .A(b[1]), .B(a[84]), .Z(n2020) );
  XOR U2301 ( .A(n2018), .B(n2022), .Z(n2021) );
  OR U2302 ( .A(n1187), .B(n1185), .Z(n2018) );
  XOR U2303 ( .A(n2024), .B(n2025), .Z(n1185) );
  NANDN U2304 ( .A(n187), .B(a[84]), .Z(n1187) );
  XNOR U2305 ( .A(n2027), .B(n1979), .Z(n1980) );
  XOR U2306 ( .A(n2028), .B(n2029), .Z(n1979) );
  ANDN U2307 ( .B(n2017), .A(n2026), .Z(n2028) );
  XNOR U2308 ( .A(n2030), .B(n2029), .Z(n2026) );
  AND U2309 ( .A(b[3]), .B(a[83]), .Z(n2030) );
  XOR U2310 ( .A(n2029), .B(n2012), .Z(n2031) );
  XOR U2311 ( .A(n2032), .B(n2033), .Z(n2012) );
  XOR U2312 ( .A(n2010), .B(n2034), .Z(n2033) );
  XNOR U2313 ( .A(n2035), .B(n2036), .Z(n2034) );
  XOR U2314 ( .A(n2037), .B(n2038), .Z(n2036) );
  NAND U2315 ( .A(b[6]), .B(a[80]), .Z(n2038) );
  AND U2316 ( .A(b[7]), .B(a[79]), .Z(n2037) );
  XNOR U2317 ( .A(n2039), .B(n2035), .Z(n2032) );
  XOR U2318 ( .A(n2040), .B(n2041), .Z(n2035) );
  NOR U2319 ( .A(n2042), .B(n2043), .Z(n2040) );
  AND U2320 ( .A(b[5]), .B(a[81]), .Z(n2039) );
  XNOR U2321 ( .A(n2044), .B(n2045), .Z(n2029) );
  ANDN U2322 ( .B(n2022), .A(n2023), .Z(n2044) );
  XOR U2323 ( .A(n2046), .B(n2045), .Z(n2023) );
  IV U2324 ( .A(n2047), .Z(n2045) );
  AND U2325 ( .A(b[2]), .B(a[83]), .Z(n2046) );
  XNOR U2326 ( .A(n2049), .B(n2047), .Z(n2048) );
  XOR U2327 ( .A(n2050), .B(n2051), .Z(n2047) );
  NANDN U2328 ( .A(n2025), .B(n2024), .Z(n2051) );
  XOR U2329 ( .A(n2050), .B(n2052), .Z(n2024) );
  NAND U2330 ( .A(b[1]), .B(a[83]), .Z(n2052) );
  XOR U2331 ( .A(n2050), .B(n2054), .Z(n2053) );
  OR U2332 ( .A(n1192), .B(n1190), .Z(n2050) );
  XOR U2333 ( .A(n2056), .B(n2057), .Z(n1190) );
  NANDN U2334 ( .A(n187), .B(a[83]), .Z(n1192) );
  XNOR U2335 ( .A(n2059), .B(n2010), .Z(n2011) );
  XNOR U2336 ( .A(n2060), .B(n2061), .Z(n2010) );
  ANDN U2337 ( .B(n2049), .A(n2058), .Z(n2060) );
  XOR U2338 ( .A(n2062), .B(n2061), .Z(n2058) );
  IV U2339 ( .A(n2063), .Z(n2061) );
  AND U2340 ( .A(b[3]), .B(a[82]), .Z(n2062) );
  XOR U2341 ( .A(n2043), .B(n2063), .Z(n2064) );
  XOR U2342 ( .A(n2065), .B(n2066), .Z(n2063) );
  ANDN U2343 ( .B(n2054), .A(n2055), .Z(n2065) );
  AND U2344 ( .A(b[2]), .B(a[82]), .Z(n2067) );
  XNOR U2345 ( .A(n2069), .B(n2066), .Z(n2068) );
  XOR U2346 ( .A(n2070), .B(n2071), .Z(n2066) );
  NANDN U2347 ( .A(n2057), .B(n2056), .Z(n2071) );
  XOR U2348 ( .A(n2070), .B(n2072), .Z(n2056) );
  NAND U2349 ( .A(b[1]), .B(a[82]), .Z(n2072) );
  XOR U2350 ( .A(n2070), .B(n2074), .Z(n2073) );
  OR U2351 ( .A(n1197), .B(n1195), .Z(n2070) );
  XOR U2352 ( .A(n2076), .B(n2077), .Z(n1195) );
  NANDN U2353 ( .A(n187), .B(a[82]), .Z(n1197) );
  XOR U2354 ( .A(n2079), .B(n2080), .Z(n2043) );
  XNOR U2355 ( .A(n2081), .B(n2082), .Z(n2080) );
  XNOR U2356 ( .A(n2083), .B(n2084), .Z(n2081) );
  XOR U2357 ( .A(n2085), .B(n2086), .Z(n2084) );
  AND U2358 ( .A(b[7]), .B(a[78]), .Z(n2086) );
  AND U2359 ( .A(b[6]), .B(a[79]), .Z(n2085) );
  XNOR U2360 ( .A(n2087), .B(n2083), .Z(n2079) );
  XOR U2361 ( .A(n2088), .B(n2089), .Z(n2083) );
  NOR U2362 ( .A(n2090), .B(n2091), .Z(n2088) );
  AND U2363 ( .A(b[5]), .B(a[80]), .Z(n2087) );
  XOR U2364 ( .A(n2092), .B(n2041), .Z(n2042) );
  IV U2365 ( .A(n2082), .Z(n2041) );
  XOR U2366 ( .A(n2093), .B(n2094), .Z(n2082) );
  ANDN U2367 ( .B(n2069), .A(n2078), .Z(n2093) );
  AND U2368 ( .A(b[3]), .B(a[81]), .Z(n2095) );
  XOR U2369 ( .A(n2091), .B(n2094), .Z(n2096) );
  XOR U2370 ( .A(n2097), .B(n2098), .Z(n2094) );
  ANDN U2371 ( .B(n2074), .A(n2075), .Z(n2097) );
  AND U2372 ( .A(b[2]), .B(a[81]), .Z(n2099) );
  XNOR U2373 ( .A(n2101), .B(n2098), .Z(n2100) );
  XOR U2374 ( .A(n2102), .B(n2103), .Z(n2098) );
  NANDN U2375 ( .A(n2077), .B(n2076), .Z(n2103) );
  XOR U2376 ( .A(n2102), .B(n2104), .Z(n2076) );
  NAND U2377 ( .A(b[1]), .B(a[81]), .Z(n2104) );
  XOR U2378 ( .A(n2102), .B(n2106), .Z(n2105) );
  OR U2379 ( .A(n1202), .B(n1200), .Z(n2102) );
  XOR U2380 ( .A(n2108), .B(n2109), .Z(n1200) );
  NANDN U2381 ( .A(n187), .B(a[81]), .Z(n1202) );
  XOR U2382 ( .A(n2111), .B(n2112), .Z(n2091) );
  XNOR U2383 ( .A(n2113), .B(n2114), .Z(n2112) );
  XNOR U2384 ( .A(n2115), .B(n2116), .Z(n2113) );
  XOR U2385 ( .A(n2117), .B(n2118), .Z(n2116) );
  AND U2386 ( .A(b[6]), .B(a[78]), .Z(n2118) );
  AND U2387 ( .A(b[7]), .B(a[77]), .Z(n2117) );
  XNOR U2388 ( .A(n2119), .B(n2115), .Z(n2111) );
  XOR U2389 ( .A(n2120), .B(n2121), .Z(n2115) );
  NOR U2390 ( .A(n2122), .B(n2123), .Z(n2120) );
  AND U2391 ( .A(b[5]), .B(a[79]), .Z(n2119) );
  XOR U2392 ( .A(n2124), .B(n2089), .Z(n2090) );
  IV U2393 ( .A(n2114), .Z(n2089) );
  XOR U2394 ( .A(n2125), .B(n2126), .Z(n2114) );
  ANDN U2395 ( .B(n2101), .A(n2110), .Z(n2125) );
  AND U2396 ( .A(b[3]), .B(a[80]), .Z(n2127) );
  XOR U2397 ( .A(n2123), .B(n2126), .Z(n2128) );
  XOR U2398 ( .A(n2129), .B(n2130), .Z(n2126) );
  ANDN U2399 ( .B(n2106), .A(n2107), .Z(n2129) );
  AND U2400 ( .A(b[2]), .B(a[80]), .Z(n2131) );
  XOR U2401 ( .A(n2133), .B(n2130), .Z(n2132) );
  XOR U2402 ( .A(n2134), .B(n2135), .Z(n2130) );
  NANDN U2403 ( .A(n2109), .B(n2108), .Z(n2135) );
  XOR U2404 ( .A(n2134), .B(n2136), .Z(n2108) );
  NAND U2405 ( .A(b[1]), .B(a[80]), .Z(n2136) );
  XOR U2406 ( .A(n2134), .B(n2138), .Z(n2137) );
  OR U2407 ( .A(n1207), .B(n1205), .Z(n2134) );
  XOR U2408 ( .A(n2140), .B(n2141), .Z(n1205) );
  NANDN U2409 ( .A(n187), .B(a[80]), .Z(n1207) );
  XOR U2410 ( .A(n2143), .B(n2144), .Z(n2123) );
  XNOR U2411 ( .A(n2145), .B(n2146), .Z(n2144) );
  XOR U2412 ( .A(n2147), .B(n2148), .Z(n2145) );
  AND U2413 ( .A(b[5]), .B(a[78]), .Z(n2147) );
  XOR U2414 ( .A(n2148), .B(n2149), .Z(n2143) );
  XOR U2415 ( .A(n2150), .B(n2151), .Z(n2149) );
  AND U2416 ( .A(b[6]), .B(a[77]), .Z(n2151) );
  AND U2417 ( .A(b[7]), .B(a[76]), .Z(n2150) );
  XOR U2418 ( .A(n2152), .B(n2153), .Z(n2148) );
  ANDN U2419 ( .B(n2154), .A(n2155), .Z(n2152) );
  XOR U2420 ( .A(n2156), .B(n2121), .Z(n2122) );
  IV U2421 ( .A(n2146), .Z(n2121) );
  XOR U2422 ( .A(n2157), .B(n2158), .Z(n2146) );
  NOR U2423 ( .A(n2142), .B(n2133), .Z(n2157) );
  XNOR U2424 ( .A(n2155), .B(n2159), .Z(n2133) );
  XNOR U2425 ( .A(n2154), .B(n2158), .Z(n2159) );
  XOR U2426 ( .A(n2160), .B(n2153), .Z(n2154) );
  AND U2427 ( .A(b[4]), .B(a[78]), .Z(n2160) );
  XOR U2428 ( .A(n2161), .B(n2162), .Z(n2155) );
  XOR U2429 ( .A(n2153), .B(n2163), .Z(n2162) );
  XOR U2430 ( .A(n2164), .B(n2165), .Z(n2163) );
  XOR U2431 ( .A(n2166), .B(n2167), .Z(n2165) );
  NAND U2432 ( .A(b[6]), .B(a[76]), .Z(n2167) );
  AND U2433 ( .A(b[7]), .B(a[75]), .Z(n2166) );
  XOR U2434 ( .A(n2168), .B(n2169), .Z(n2153) );
  ANDN U2435 ( .B(n2170), .A(n2171), .Z(n2168) );
  XOR U2436 ( .A(n2172), .B(n2164), .Z(n2161) );
  XOR U2437 ( .A(n2173), .B(n2174), .Z(n2164) );
  NOR U2438 ( .A(n2175), .B(n2176), .Z(n2173) );
  AND U2439 ( .A(b[5]), .B(a[77]), .Z(n2172) );
  XOR U2440 ( .A(n2178), .B(n2179), .Z(n2158) );
  ANDN U2441 ( .B(n2138), .A(n2139), .Z(n2178) );
  AND U2442 ( .A(b[2]), .B(a[79]), .Z(n2180) );
  XNOR U2443 ( .A(n2170), .B(n2179), .Z(n2181) );
  XOR U2444 ( .A(n2182), .B(n2183), .Z(n2179) );
  NANDN U2445 ( .A(n2141), .B(n2140), .Z(n2183) );
  XOR U2446 ( .A(n2182), .B(n2184), .Z(n2140) );
  NAND U2447 ( .A(b[1]), .B(a[79]), .Z(n2184) );
  XNOR U2448 ( .A(n2182), .B(n2186), .Z(n2185) );
  OR U2449 ( .A(n1212), .B(n1210), .Z(n2182) );
  NANDN U2450 ( .A(n187), .B(a[79]), .Z(n1212) );
  XOR U2451 ( .A(n2190), .B(n2169), .Z(n2170) );
  AND U2452 ( .A(b[3]), .B(a[78]), .Z(n2190) );
  XOR U2453 ( .A(n2169), .B(n2176), .Z(n2191) );
  XOR U2454 ( .A(n2192), .B(n2193), .Z(n2176) );
  XOR U2455 ( .A(n2174), .B(n2194), .Z(n2193) );
  XOR U2456 ( .A(n2195), .B(n2196), .Z(n2194) );
  XOR U2457 ( .A(n2197), .B(n2198), .Z(n2196) );
  NAND U2458 ( .A(b[6]), .B(a[75]), .Z(n2198) );
  AND U2459 ( .A(b[7]), .B(a[74]), .Z(n2197) );
  XOR U2460 ( .A(n2199), .B(n2195), .Z(n2192) );
  XOR U2461 ( .A(n2200), .B(n2201), .Z(n2195) );
  NOR U2462 ( .A(n2202), .B(n2203), .Z(n2200) );
  AND U2463 ( .A(b[5]), .B(a[76]), .Z(n2199) );
  XNOR U2464 ( .A(n2204), .B(n2205), .Z(n2169) );
  NOR U2465 ( .A(n2187), .B(n2186), .Z(n2204) );
  XOR U2466 ( .A(n2206), .B(n2205), .Z(n2186) );
  AND U2467 ( .A(b[2]), .B(a[78]), .Z(n2206) );
  XOR U2468 ( .A(n2205), .B(n2208), .Z(n2207) );
  XNOR U2469 ( .A(n2209), .B(n2210), .Z(n2205) );
  OR U2470 ( .A(n2188), .B(n2189), .Z(n2210) );
  XNOR U2471 ( .A(n2209), .B(n2212), .Z(n2211) );
  XNOR U2472 ( .A(n2209), .B(n2214), .Z(n2188) );
  NAND U2473 ( .A(b[1]), .B(a[78]), .Z(n2214) );
  OR U2474 ( .A(n1217), .B(n1215), .Z(n2209) );
  XOR U2475 ( .A(n2215), .B(n2216), .Z(n1215) );
  NANDN U2476 ( .A(n187), .B(a[78]), .Z(n1217) );
  XNOR U2477 ( .A(n2218), .B(n2174), .Z(n2175) );
  XOR U2478 ( .A(n2219), .B(n2220), .Z(n2174) );
  ANDN U2479 ( .B(n2208), .A(n2217), .Z(n2219) );
  XNOR U2480 ( .A(n2221), .B(n2220), .Z(n2217) );
  AND U2481 ( .A(b[3]), .B(a[77]), .Z(n2221) );
  XOR U2482 ( .A(n2220), .B(n2203), .Z(n2222) );
  XOR U2483 ( .A(n2223), .B(n2224), .Z(n2203) );
  XOR U2484 ( .A(n2201), .B(n2225), .Z(n2224) );
  XOR U2485 ( .A(n2226), .B(n2227), .Z(n2225) );
  XOR U2486 ( .A(n2228), .B(n2229), .Z(n2227) );
  NAND U2487 ( .A(b[6]), .B(a[74]), .Z(n2229) );
  AND U2488 ( .A(b[7]), .B(a[73]), .Z(n2228) );
  XOR U2489 ( .A(n2230), .B(n2226), .Z(n2223) );
  XOR U2490 ( .A(n2231), .B(n2232), .Z(n2226) );
  NOR U2491 ( .A(n2233), .B(n2234), .Z(n2231) );
  AND U2492 ( .A(b[5]), .B(a[75]), .Z(n2230) );
  XNOR U2493 ( .A(n2235), .B(n2236), .Z(n2220) );
  NOR U2494 ( .A(n2213), .B(n2212), .Z(n2235) );
  XOR U2495 ( .A(n2237), .B(n2236), .Z(n2212) );
  AND U2496 ( .A(b[2]), .B(a[77]), .Z(n2237) );
  XOR U2497 ( .A(n2236), .B(n2239), .Z(n2238) );
  XNOR U2498 ( .A(n2240), .B(n2241), .Z(n2236) );
  NANDN U2499 ( .A(n2216), .B(n2215), .Z(n2241) );
  XOR U2500 ( .A(n2240), .B(n2242), .Z(n2215) );
  NAND U2501 ( .A(b[1]), .B(a[77]), .Z(n2242) );
  XOR U2502 ( .A(n2240), .B(n2244), .Z(n2243) );
  OR U2503 ( .A(n1222), .B(n1220), .Z(n2240) );
  XOR U2504 ( .A(n2246), .B(n2247), .Z(n1220) );
  NANDN U2505 ( .A(n187), .B(a[77]), .Z(n1222) );
  XNOR U2506 ( .A(n2249), .B(n2201), .Z(n2202) );
  XOR U2507 ( .A(n2250), .B(n2251), .Z(n2201) );
  ANDN U2508 ( .B(n2239), .A(n2248), .Z(n2250) );
  XNOR U2509 ( .A(n2252), .B(n2251), .Z(n2248) );
  AND U2510 ( .A(b[3]), .B(a[76]), .Z(n2252) );
  XOR U2511 ( .A(n2251), .B(n2234), .Z(n2253) );
  XOR U2512 ( .A(n2254), .B(n2255), .Z(n2234) );
  XOR U2513 ( .A(n2232), .B(n2256), .Z(n2255) );
  XNOR U2514 ( .A(n2257), .B(n2258), .Z(n2256) );
  XOR U2515 ( .A(n2259), .B(n2260), .Z(n2258) );
  NAND U2516 ( .A(b[6]), .B(a[73]), .Z(n2260) );
  AND U2517 ( .A(b[7]), .B(a[72]), .Z(n2259) );
  XNOR U2518 ( .A(n2261), .B(n2257), .Z(n2254) );
  XOR U2519 ( .A(n2262), .B(n2263), .Z(n2257) );
  NOR U2520 ( .A(n2264), .B(n2265), .Z(n2262) );
  AND U2521 ( .A(b[5]), .B(a[74]), .Z(n2261) );
  XNOR U2522 ( .A(n2266), .B(n2267), .Z(n2251) );
  ANDN U2523 ( .B(n2244), .A(n2245), .Z(n2266) );
  XOR U2524 ( .A(n2268), .B(n2267), .Z(n2245) );
  IV U2525 ( .A(n2269), .Z(n2267) );
  AND U2526 ( .A(b[2]), .B(a[76]), .Z(n2268) );
  XNOR U2527 ( .A(n2271), .B(n2269), .Z(n2270) );
  XOR U2528 ( .A(n2272), .B(n2273), .Z(n2269) );
  NANDN U2529 ( .A(n2247), .B(n2246), .Z(n2273) );
  XOR U2530 ( .A(n2272), .B(n2274), .Z(n2246) );
  NAND U2531 ( .A(b[1]), .B(a[76]), .Z(n2274) );
  XOR U2532 ( .A(n2272), .B(n2276), .Z(n2275) );
  OR U2533 ( .A(n1227), .B(n1225), .Z(n2272) );
  XOR U2534 ( .A(n2278), .B(n2279), .Z(n1225) );
  NANDN U2535 ( .A(n187), .B(a[76]), .Z(n1227) );
  XNOR U2536 ( .A(n2281), .B(n2232), .Z(n2233) );
  XNOR U2537 ( .A(n2282), .B(n2283), .Z(n2232) );
  ANDN U2538 ( .B(n2271), .A(n2280), .Z(n2282) );
  XOR U2539 ( .A(n2284), .B(n2283), .Z(n2280) );
  IV U2540 ( .A(n2285), .Z(n2283) );
  AND U2541 ( .A(b[3]), .B(a[75]), .Z(n2284) );
  XOR U2542 ( .A(n2265), .B(n2285), .Z(n2286) );
  XOR U2543 ( .A(n2287), .B(n2288), .Z(n2285) );
  ANDN U2544 ( .B(n2276), .A(n2277), .Z(n2287) );
  AND U2545 ( .A(b[2]), .B(a[75]), .Z(n2289) );
  XNOR U2546 ( .A(n2291), .B(n2288), .Z(n2290) );
  XOR U2547 ( .A(n2292), .B(n2293), .Z(n2288) );
  NANDN U2548 ( .A(n2279), .B(n2278), .Z(n2293) );
  XOR U2549 ( .A(n2292), .B(n2294), .Z(n2278) );
  NAND U2550 ( .A(b[1]), .B(a[75]), .Z(n2294) );
  XOR U2551 ( .A(n2292), .B(n2296), .Z(n2295) );
  OR U2552 ( .A(n1232), .B(n1230), .Z(n2292) );
  XOR U2553 ( .A(n2298), .B(n2299), .Z(n1230) );
  NANDN U2554 ( .A(n187), .B(a[75]), .Z(n1232) );
  XOR U2555 ( .A(n2301), .B(n2302), .Z(n2265) );
  XNOR U2556 ( .A(n2303), .B(n2304), .Z(n2302) );
  XNOR U2557 ( .A(n2305), .B(n2306), .Z(n2303) );
  XOR U2558 ( .A(n2307), .B(n2308), .Z(n2306) );
  AND U2559 ( .A(b[7]), .B(a[71]), .Z(n2308) );
  AND U2560 ( .A(b[6]), .B(a[72]), .Z(n2307) );
  XNOR U2561 ( .A(n2309), .B(n2305), .Z(n2301) );
  XOR U2562 ( .A(n2310), .B(n2311), .Z(n2305) );
  NOR U2563 ( .A(n2312), .B(n2313), .Z(n2310) );
  AND U2564 ( .A(b[5]), .B(a[73]), .Z(n2309) );
  XOR U2565 ( .A(n2314), .B(n2263), .Z(n2264) );
  IV U2566 ( .A(n2304), .Z(n2263) );
  XOR U2567 ( .A(n2315), .B(n2316), .Z(n2304) );
  ANDN U2568 ( .B(n2291), .A(n2300), .Z(n2315) );
  AND U2569 ( .A(b[3]), .B(a[74]), .Z(n2317) );
  XOR U2570 ( .A(n2313), .B(n2316), .Z(n2318) );
  XOR U2571 ( .A(n2319), .B(n2320), .Z(n2316) );
  ANDN U2572 ( .B(n2296), .A(n2297), .Z(n2319) );
  AND U2573 ( .A(b[2]), .B(a[74]), .Z(n2321) );
  XNOR U2574 ( .A(n2323), .B(n2320), .Z(n2322) );
  XOR U2575 ( .A(n2324), .B(n2325), .Z(n2320) );
  NANDN U2576 ( .A(n2299), .B(n2298), .Z(n2325) );
  XOR U2577 ( .A(n2324), .B(n2326), .Z(n2298) );
  NAND U2578 ( .A(b[1]), .B(a[74]), .Z(n2326) );
  XOR U2579 ( .A(n2324), .B(n2328), .Z(n2327) );
  OR U2580 ( .A(n1237), .B(n1235), .Z(n2324) );
  XOR U2581 ( .A(n2330), .B(n2331), .Z(n1235) );
  NANDN U2582 ( .A(n187), .B(a[74]), .Z(n1237) );
  XOR U2583 ( .A(n2333), .B(n2334), .Z(n2313) );
  XNOR U2584 ( .A(n2335), .B(n2336), .Z(n2334) );
  XNOR U2585 ( .A(n2337), .B(n2338), .Z(n2335) );
  XOR U2586 ( .A(n2339), .B(n2340), .Z(n2338) );
  AND U2587 ( .A(b[6]), .B(a[71]), .Z(n2340) );
  AND U2588 ( .A(b[7]), .B(a[70]), .Z(n2339) );
  XNOR U2589 ( .A(n2341), .B(n2337), .Z(n2333) );
  XOR U2590 ( .A(n2342), .B(n2343), .Z(n2337) );
  NOR U2591 ( .A(n2344), .B(n2345), .Z(n2342) );
  AND U2592 ( .A(b[5]), .B(a[72]), .Z(n2341) );
  XOR U2593 ( .A(n2346), .B(n2311), .Z(n2312) );
  IV U2594 ( .A(n2336), .Z(n2311) );
  XOR U2595 ( .A(n2347), .B(n2348), .Z(n2336) );
  ANDN U2596 ( .B(n2323), .A(n2332), .Z(n2347) );
  AND U2597 ( .A(b[3]), .B(a[73]), .Z(n2349) );
  XOR U2598 ( .A(n2345), .B(n2348), .Z(n2350) );
  XOR U2599 ( .A(n2351), .B(n2352), .Z(n2348) );
  ANDN U2600 ( .B(n2328), .A(n2329), .Z(n2351) );
  AND U2601 ( .A(b[2]), .B(a[73]), .Z(n2353) );
  XOR U2602 ( .A(n2355), .B(n2352), .Z(n2354) );
  XOR U2603 ( .A(n2356), .B(n2357), .Z(n2352) );
  NANDN U2604 ( .A(n2331), .B(n2330), .Z(n2357) );
  XOR U2605 ( .A(n2356), .B(n2358), .Z(n2330) );
  NAND U2606 ( .A(b[1]), .B(a[73]), .Z(n2358) );
  XOR U2607 ( .A(n2356), .B(n2360), .Z(n2359) );
  OR U2608 ( .A(n1242), .B(n1240), .Z(n2356) );
  XOR U2609 ( .A(n2362), .B(n2363), .Z(n1240) );
  NANDN U2610 ( .A(n187), .B(a[73]), .Z(n1242) );
  XOR U2611 ( .A(n2365), .B(n2366), .Z(n2345) );
  XNOR U2612 ( .A(n2367), .B(n2368), .Z(n2366) );
  XOR U2613 ( .A(n2369), .B(n2370), .Z(n2367) );
  AND U2614 ( .A(b[5]), .B(a[71]), .Z(n2369) );
  XOR U2615 ( .A(n2370), .B(n2371), .Z(n2365) );
  XOR U2616 ( .A(n2372), .B(n2373), .Z(n2371) );
  AND U2617 ( .A(b[6]), .B(a[70]), .Z(n2373) );
  AND U2618 ( .A(b[7]), .B(a[69]), .Z(n2372) );
  XOR U2619 ( .A(n2374), .B(n2375), .Z(n2370) );
  ANDN U2620 ( .B(n2376), .A(n2377), .Z(n2374) );
  XOR U2621 ( .A(n2378), .B(n2343), .Z(n2344) );
  IV U2622 ( .A(n2368), .Z(n2343) );
  XOR U2623 ( .A(n2379), .B(n2380), .Z(n2368) );
  NOR U2624 ( .A(n2364), .B(n2355), .Z(n2379) );
  XNOR U2625 ( .A(n2377), .B(n2381), .Z(n2355) );
  XNOR U2626 ( .A(n2376), .B(n2380), .Z(n2381) );
  XOR U2627 ( .A(n2382), .B(n2375), .Z(n2376) );
  AND U2628 ( .A(b[4]), .B(a[71]), .Z(n2382) );
  XOR U2629 ( .A(n2383), .B(n2384), .Z(n2377) );
  XOR U2630 ( .A(n2375), .B(n2385), .Z(n2384) );
  XOR U2631 ( .A(n2386), .B(n2387), .Z(n2385) );
  XOR U2632 ( .A(n2388), .B(n2389), .Z(n2387) );
  NAND U2633 ( .A(b[6]), .B(a[69]), .Z(n2389) );
  AND U2634 ( .A(b[7]), .B(a[68]), .Z(n2388) );
  XOR U2635 ( .A(n2390), .B(n2391), .Z(n2375) );
  ANDN U2636 ( .B(n2392), .A(n2393), .Z(n2390) );
  XOR U2637 ( .A(n2394), .B(n2386), .Z(n2383) );
  XOR U2638 ( .A(n2395), .B(n2396), .Z(n2386) );
  NOR U2639 ( .A(n2397), .B(n2398), .Z(n2395) );
  AND U2640 ( .A(b[5]), .B(a[70]), .Z(n2394) );
  XOR U2641 ( .A(n2400), .B(n2401), .Z(n2380) );
  ANDN U2642 ( .B(n2360), .A(n2361), .Z(n2400) );
  AND U2643 ( .A(b[2]), .B(a[72]), .Z(n2402) );
  XNOR U2644 ( .A(n2392), .B(n2401), .Z(n2403) );
  XOR U2645 ( .A(n2404), .B(n2405), .Z(n2401) );
  NANDN U2646 ( .A(n2363), .B(n2362), .Z(n2405) );
  XOR U2647 ( .A(n2404), .B(n2406), .Z(n2362) );
  NAND U2648 ( .A(b[1]), .B(a[72]), .Z(n2406) );
  XNOR U2649 ( .A(n2404), .B(n2408), .Z(n2407) );
  OR U2650 ( .A(n1247), .B(n1245), .Z(n2404) );
  NANDN U2651 ( .A(n187), .B(a[72]), .Z(n1247) );
  XOR U2652 ( .A(n2412), .B(n2391), .Z(n2392) );
  AND U2653 ( .A(b[3]), .B(a[71]), .Z(n2412) );
  XOR U2654 ( .A(n2391), .B(n2398), .Z(n2413) );
  XOR U2655 ( .A(n2414), .B(n2415), .Z(n2398) );
  XOR U2656 ( .A(n2396), .B(n2416), .Z(n2415) );
  XOR U2657 ( .A(n2417), .B(n2418), .Z(n2416) );
  XOR U2658 ( .A(n2419), .B(n2420), .Z(n2418) );
  NAND U2659 ( .A(b[6]), .B(a[68]), .Z(n2420) );
  AND U2660 ( .A(b[7]), .B(a[67]), .Z(n2419) );
  XOR U2661 ( .A(n2421), .B(n2417), .Z(n2414) );
  XOR U2662 ( .A(n2422), .B(n2423), .Z(n2417) );
  NOR U2663 ( .A(n2424), .B(n2425), .Z(n2422) );
  AND U2664 ( .A(b[5]), .B(a[69]), .Z(n2421) );
  XNOR U2665 ( .A(n2426), .B(n2427), .Z(n2391) );
  NOR U2666 ( .A(n2409), .B(n2408), .Z(n2426) );
  XOR U2667 ( .A(n2428), .B(n2427), .Z(n2408) );
  AND U2668 ( .A(b[2]), .B(a[71]), .Z(n2428) );
  XOR U2669 ( .A(n2427), .B(n2430), .Z(n2429) );
  XNOR U2670 ( .A(n2431), .B(n2432), .Z(n2427) );
  OR U2671 ( .A(n2410), .B(n2411), .Z(n2432) );
  XNOR U2672 ( .A(n2431), .B(n2434), .Z(n2433) );
  XNOR U2673 ( .A(n2431), .B(n2436), .Z(n2410) );
  NAND U2674 ( .A(b[1]), .B(a[71]), .Z(n2436) );
  OR U2675 ( .A(n1252), .B(n1250), .Z(n2431) );
  XOR U2676 ( .A(n2437), .B(n2438), .Z(n1250) );
  NANDN U2677 ( .A(n187), .B(a[71]), .Z(n1252) );
  XNOR U2678 ( .A(n2440), .B(n2396), .Z(n2397) );
  XOR U2679 ( .A(n2441), .B(n2442), .Z(n2396) );
  ANDN U2680 ( .B(n2430), .A(n2439), .Z(n2441) );
  XNOR U2681 ( .A(n2443), .B(n2442), .Z(n2439) );
  AND U2682 ( .A(b[3]), .B(a[70]), .Z(n2443) );
  XOR U2683 ( .A(n2442), .B(n2425), .Z(n2444) );
  XOR U2684 ( .A(n2445), .B(n2446), .Z(n2425) );
  XOR U2685 ( .A(n2423), .B(n2447), .Z(n2446) );
  XOR U2686 ( .A(n2448), .B(n2449), .Z(n2447) );
  XOR U2687 ( .A(n2450), .B(n2451), .Z(n2449) );
  NAND U2688 ( .A(b[6]), .B(a[67]), .Z(n2451) );
  AND U2689 ( .A(b[7]), .B(a[66]), .Z(n2450) );
  XOR U2690 ( .A(n2452), .B(n2448), .Z(n2445) );
  XOR U2691 ( .A(n2453), .B(n2454), .Z(n2448) );
  NOR U2692 ( .A(n2455), .B(n2456), .Z(n2453) );
  AND U2693 ( .A(b[5]), .B(a[68]), .Z(n2452) );
  XNOR U2694 ( .A(n2457), .B(n2458), .Z(n2442) );
  NOR U2695 ( .A(n2435), .B(n2434), .Z(n2457) );
  XOR U2696 ( .A(n2459), .B(n2458), .Z(n2434) );
  AND U2697 ( .A(b[2]), .B(a[70]), .Z(n2459) );
  XOR U2698 ( .A(n2458), .B(n2461), .Z(n2460) );
  XNOR U2699 ( .A(n2462), .B(n2463), .Z(n2458) );
  NANDN U2700 ( .A(n2438), .B(n2437), .Z(n2463) );
  XOR U2701 ( .A(n2462), .B(n2464), .Z(n2437) );
  NAND U2702 ( .A(b[1]), .B(a[70]), .Z(n2464) );
  XOR U2703 ( .A(n2462), .B(n2466), .Z(n2465) );
  OR U2704 ( .A(n1257), .B(n1255), .Z(n2462) );
  XOR U2705 ( .A(n2468), .B(n2469), .Z(n1255) );
  NANDN U2706 ( .A(n187), .B(a[70]), .Z(n1257) );
  XNOR U2707 ( .A(n2471), .B(n2423), .Z(n2424) );
  XOR U2708 ( .A(n2472), .B(n2473), .Z(n2423) );
  ANDN U2709 ( .B(n2461), .A(n2470), .Z(n2472) );
  XNOR U2710 ( .A(n2474), .B(n2473), .Z(n2470) );
  AND U2711 ( .A(b[3]), .B(a[69]), .Z(n2474) );
  XOR U2712 ( .A(n2473), .B(n2456), .Z(n2475) );
  XOR U2713 ( .A(n2476), .B(n2477), .Z(n2456) );
  XOR U2714 ( .A(n2454), .B(n2478), .Z(n2477) );
  XNOR U2715 ( .A(n2479), .B(n2480), .Z(n2478) );
  XOR U2716 ( .A(n2481), .B(n2482), .Z(n2480) );
  NAND U2717 ( .A(b[6]), .B(a[66]), .Z(n2482) );
  AND U2718 ( .A(b[7]), .B(a[65]), .Z(n2481) );
  XNOR U2719 ( .A(n2483), .B(n2479), .Z(n2476) );
  XOR U2720 ( .A(n2484), .B(n2485), .Z(n2479) );
  NOR U2721 ( .A(n2486), .B(n2487), .Z(n2484) );
  AND U2722 ( .A(b[5]), .B(a[67]), .Z(n2483) );
  XNOR U2723 ( .A(n2488), .B(n2489), .Z(n2473) );
  ANDN U2724 ( .B(n2466), .A(n2467), .Z(n2488) );
  XOR U2725 ( .A(n2490), .B(n2489), .Z(n2467) );
  IV U2726 ( .A(n2491), .Z(n2489) );
  AND U2727 ( .A(b[2]), .B(a[69]), .Z(n2490) );
  XNOR U2728 ( .A(n2493), .B(n2491), .Z(n2492) );
  XOR U2729 ( .A(n2494), .B(n2495), .Z(n2491) );
  NANDN U2730 ( .A(n2469), .B(n2468), .Z(n2495) );
  XOR U2731 ( .A(n2494), .B(n2496), .Z(n2468) );
  NAND U2732 ( .A(b[1]), .B(a[69]), .Z(n2496) );
  XOR U2733 ( .A(n2494), .B(n2498), .Z(n2497) );
  OR U2734 ( .A(n1262), .B(n1260), .Z(n2494) );
  XOR U2735 ( .A(n2500), .B(n2501), .Z(n1260) );
  NANDN U2736 ( .A(n187), .B(a[69]), .Z(n1262) );
  XNOR U2737 ( .A(n2503), .B(n2454), .Z(n2455) );
  XNOR U2738 ( .A(n2504), .B(n2505), .Z(n2454) );
  ANDN U2739 ( .B(n2493), .A(n2502), .Z(n2504) );
  XOR U2740 ( .A(n2506), .B(n2505), .Z(n2502) );
  IV U2741 ( .A(n2507), .Z(n2505) );
  AND U2742 ( .A(b[3]), .B(a[68]), .Z(n2506) );
  XOR U2743 ( .A(n2487), .B(n2507), .Z(n2508) );
  XOR U2744 ( .A(n2509), .B(n2510), .Z(n2507) );
  ANDN U2745 ( .B(n2498), .A(n2499), .Z(n2509) );
  AND U2746 ( .A(b[2]), .B(a[68]), .Z(n2511) );
  XNOR U2747 ( .A(n2513), .B(n2510), .Z(n2512) );
  XOR U2748 ( .A(n2514), .B(n2515), .Z(n2510) );
  NANDN U2749 ( .A(n2501), .B(n2500), .Z(n2515) );
  XOR U2750 ( .A(n2514), .B(n2516), .Z(n2500) );
  NAND U2751 ( .A(b[1]), .B(a[68]), .Z(n2516) );
  XOR U2752 ( .A(n2514), .B(n2518), .Z(n2517) );
  OR U2753 ( .A(n1267), .B(n1265), .Z(n2514) );
  XOR U2754 ( .A(n2520), .B(n2521), .Z(n1265) );
  NANDN U2755 ( .A(n187), .B(a[68]), .Z(n1267) );
  XOR U2756 ( .A(n2523), .B(n2524), .Z(n2487) );
  XNOR U2757 ( .A(n2525), .B(n2526), .Z(n2524) );
  XNOR U2758 ( .A(n2527), .B(n2528), .Z(n2525) );
  XOR U2759 ( .A(n2529), .B(n2530), .Z(n2528) );
  AND U2760 ( .A(b[7]), .B(a[64]), .Z(n2530) );
  AND U2761 ( .A(b[6]), .B(a[65]), .Z(n2529) );
  XNOR U2762 ( .A(n2531), .B(n2527), .Z(n2523) );
  XOR U2763 ( .A(n2532), .B(n2533), .Z(n2527) );
  NOR U2764 ( .A(n2534), .B(n2535), .Z(n2532) );
  AND U2765 ( .A(b[5]), .B(a[66]), .Z(n2531) );
  XOR U2766 ( .A(n2536), .B(n2485), .Z(n2486) );
  IV U2767 ( .A(n2526), .Z(n2485) );
  XOR U2768 ( .A(n2537), .B(n2538), .Z(n2526) );
  ANDN U2769 ( .B(n2513), .A(n2522), .Z(n2537) );
  AND U2770 ( .A(b[3]), .B(a[67]), .Z(n2539) );
  XOR U2771 ( .A(n2535), .B(n2538), .Z(n2540) );
  XOR U2772 ( .A(n2541), .B(n2542), .Z(n2538) );
  ANDN U2773 ( .B(n2518), .A(n2519), .Z(n2541) );
  AND U2774 ( .A(b[2]), .B(a[67]), .Z(n2543) );
  XNOR U2775 ( .A(n2545), .B(n2542), .Z(n2544) );
  XOR U2776 ( .A(n2546), .B(n2547), .Z(n2542) );
  NANDN U2777 ( .A(n2521), .B(n2520), .Z(n2547) );
  XOR U2778 ( .A(n2546), .B(n2548), .Z(n2520) );
  NAND U2779 ( .A(b[1]), .B(a[67]), .Z(n2548) );
  XOR U2780 ( .A(n2546), .B(n2550), .Z(n2549) );
  OR U2781 ( .A(n1272), .B(n1270), .Z(n2546) );
  XOR U2782 ( .A(n2552), .B(n2553), .Z(n1270) );
  NANDN U2783 ( .A(n187), .B(a[67]), .Z(n1272) );
  XOR U2784 ( .A(n2555), .B(n2556), .Z(n2535) );
  XNOR U2785 ( .A(n2557), .B(n2558), .Z(n2556) );
  XNOR U2786 ( .A(n2559), .B(n2560), .Z(n2557) );
  XOR U2787 ( .A(n2561), .B(n2562), .Z(n2560) );
  AND U2788 ( .A(b[6]), .B(a[64]), .Z(n2562) );
  AND U2789 ( .A(b[7]), .B(a[63]), .Z(n2561) );
  XNOR U2790 ( .A(n2563), .B(n2559), .Z(n2555) );
  XOR U2791 ( .A(n2564), .B(n2565), .Z(n2559) );
  NOR U2792 ( .A(n2566), .B(n2567), .Z(n2564) );
  AND U2793 ( .A(b[5]), .B(a[65]), .Z(n2563) );
  XOR U2794 ( .A(n2568), .B(n2533), .Z(n2534) );
  IV U2795 ( .A(n2558), .Z(n2533) );
  XOR U2796 ( .A(n2569), .B(n2570), .Z(n2558) );
  ANDN U2797 ( .B(n2545), .A(n2554), .Z(n2569) );
  AND U2798 ( .A(b[3]), .B(a[66]), .Z(n2571) );
  XOR U2799 ( .A(n2567), .B(n2570), .Z(n2572) );
  XOR U2800 ( .A(n2573), .B(n2574), .Z(n2570) );
  ANDN U2801 ( .B(n2550), .A(n2551), .Z(n2573) );
  AND U2802 ( .A(b[2]), .B(a[66]), .Z(n2575) );
  XOR U2803 ( .A(n2577), .B(n2574), .Z(n2576) );
  XOR U2804 ( .A(n2578), .B(n2579), .Z(n2574) );
  NANDN U2805 ( .A(n2553), .B(n2552), .Z(n2579) );
  XOR U2806 ( .A(n2578), .B(n2580), .Z(n2552) );
  NAND U2807 ( .A(b[1]), .B(a[66]), .Z(n2580) );
  XOR U2808 ( .A(n2578), .B(n2582), .Z(n2581) );
  OR U2809 ( .A(n1277), .B(n1275), .Z(n2578) );
  XOR U2810 ( .A(n2584), .B(n2585), .Z(n1275) );
  NANDN U2811 ( .A(n187), .B(a[66]), .Z(n1277) );
  XOR U2812 ( .A(n2587), .B(n2588), .Z(n2567) );
  XNOR U2813 ( .A(n2589), .B(n2590), .Z(n2588) );
  XOR U2814 ( .A(n2591), .B(n2592), .Z(n2589) );
  AND U2815 ( .A(b[5]), .B(a[64]), .Z(n2591) );
  XOR U2816 ( .A(n2592), .B(n2593), .Z(n2587) );
  XOR U2817 ( .A(n2594), .B(n2595), .Z(n2593) );
  AND U2818 ( .A(b[6]), .B(a[63]), .Z(n2595) );
  AND U2819 ( .A(b[7]), .B(a[62]), .Z(n2594) );
  XOR U2820 ( .A(n2596), .B(n2597), .Z(n2592) );
  ANDN U2821 ( .B(n2598), .A(n2599), .Z(n2596) );
  XOR U2822 ( .A(n2600), .B(n2565), .Z(n2566) );
  IV U2823 ( .A(n2590), .Z(n2565) );
  XOR U2824 ( .A(n2601), .B(n2602), .Z(n2590) );
  NOR U2825 ( .A(n2586), .B(n2577), .Z(n2601) );
  XNOR U2826 ( .A(n2599), .B(n2603), .Z(n2577) );
  XNOR U2827 ( .A(n2598), .B(n2602), .Z(n2603) );
  XOR U2828 ( .A(n2604), .B(n2597), .Z(n2598) );
  AND U2829 ( .A(b[4]), .B(a[64]), .Z(n2604) );
  XOR U2830 ( .A(n2605), .B(n2606), .Z(n2599) );
  XOR U2831 ( .A(n2597), .B(n2607), .Z(n2606) );
  XOR U2832 ( .A(n2608), .B(n2609), .Z(n2607) );
  XOR U2833 ( .A(n2610), .B(n2611), .Z(n2609) );
  NAND U2834 ( .A(b[6]), .B(a[62]), .Z(n2611) );
  AND U2835 ( .A(b[7]), .B(a[61]), .Z(n2610) );
  XOR U2836 ( .A(n2612), .B(n2613), .Z(n2597) );
  ANDN U2837 ( .B(n2614), .A(n2615), .Z(n2612) );
  XOR U2838 ( .A(n2616), .B(n2608), .Z(n2605) );
  XOR U2839 ( .A(n2617), .B(n2618), .Z(n2608) );
  NOR U2840 ( .A(n2619), .B(n2620), .Z(n2617) );
  AND U2841 ( .A(b[5]), .B(a[63]), .Z(n2616) );
  XOR U2842 ( .A(n2622), .B(n2623), .Z(n2602) );
  ANDN U2843 ( .B(n2582), .A(n2583), .Z(n2622) );
  AND U2844 ( .A(b[2]), .B(a[65]), .Z(n2624) );
  XNOR U2845 ( .A(n2614), .B(n2623), .Z(n2625) );
  XOR U2846 ( .A(n2626), .B(n2627), .Z(n2623) );
  NANDN U2847 ( .A(n2585), .B(n2584), .Z(n2627) );
  XOR U2848 ( .A(n2626), .B(n2628), .Z(n2584) );
  NAND U2849 ( .A(b[1]), .B(a[65]), .Z(n2628) );
  XNOR U2850 ( .A(n2626), .B(n2630), .Z(n2629) );
  OR U2851 ( .A(n1282), .B(n1280), .Z(n2626) );
  NANDN U2852 ( .A(n187), .B(a[65]), .Z(n1282) );
  XOR U2853 ( .A(n2634), .B(n2613), .Z(n2614) );
  AND U2854 ( .A(b[3]), .B(a[64]), .Z(n2634) );
  XOR U2855 ( .A(n2613), .B(n2620), .Z(n2635) );
  XOR U2856 ( .A(n2636), .B(n2637), .Z(n2620) );
  XOR U2857 ( .A(n2618), .B(n2638), .Z(n2637) );
  XOR U2858 ( .A(n2639), .B(n2640), .Z(n2638) );
  XOR U2859 ( .A(n2641), .B(n2642), .Z(n2640) );
  NAND U2860 ( .A(b[6]), .B(a[61]), .Z(n2642) );
  AND U2861 ( .A(b[7]), .B(a[60]), .Z(n2641) );
  XOR U2862 ( .A(n2643), .B(n2639), .Z(n2636) );
  XOR U2863 ( .A(n2644), .B(n2645), .Z(n2639) );
  NOR U2864 ( .A(n2646), .B(n2647), .Z(n2644) );
  AND U2865 ( .A(b[5]), .B(a[62]), .Z(n2643) );
  XNOR U2866 ( .A(n2648), .B(n2649), .Z(n2613) );
  NOR U2867 ( .A(n2631), .B(n2630), .Z(n2648) );
  XOR U2868 ( .A(n2650), .B(n2649), .Z(n2630) );
  AND U2869 ( .A(b[2]), .B(a[64]), .Z(n2650) );
  XOR U2870 ( .A(n2649), .B(n2652), .Z(n2651) );
  XNOR U2871 ( .A(n2653), .B(n2654), .Z(n2649) );
  OR U2872 ( .A(n2632), .B(n2633), .Z(n2654) );
  XNOR U2873 ( .A(n2653), .B(n2656), .Z(n2655) );
  XNOR U2874 ( .A(n2653), .B(n2658), .Z(n2632) );
  NAND U2875 ( .A(b[1]), .B(a[64]), .Z(n2658) );
  OR U2876 ( .A(n1287), .B(n1285), .Z(n2653) );
  XOR U2877 ( .A(n2659), .B(n2660), .Z(n1285) );
  NANDN U2878 ( .A(n187), .B(a[64]), .Z(n1287) );
  XNOR U2879 ( .A(n2662), .B(n2618), .Z(n2619) );
  XOR U2880 ( .A(n2663), .B(n2664), .Z(n2618) );
  ANDN U2881 ( .B(n2652), .A(n2661), .Z(n2663) );
  XNOR U2882 ( .A(n2665), .B(n2664), .Z(n2661) );
  AND U2883 ( .A(b[3]), .B(a[63]), .Z(n2665) );
  XOR U2884 ( .A(n2664), .B(n2647), .Z(n2666) );
  XOR U2885 ( .A(n2667), .B(n2668), .Z(n2647) );
  XOR U2886 ( .A(n2645), .B(n2669), .Z(n2668) );
  XOR U2887 ( .A(n2670), .B(n2671), .Z(n2669) );
  XOR U2888 ( .A(n2672), .B(n2673), .Z(n2671) );
  NAND U2889 ( .A(b[6]), .B(a[60]), .Z(n2673) );
  AND U2890 ( .A(b[7]), .B(a[59]), .Z(n2672) );
  XOR U2891 ( .A(n2674), .B(n2670), .Z(n2667) );
  XOR U2892 ( .A(n2675), .B(n2676), .Z(n2670) );
  NOR U2893 ( .A(n2677), .B(n2678), .Z(n2675) );
  AND U2894 ( .A(b[5]), .B(a[61]), .Z(n2674) );
  XNOR U2895 ( .A(n2679), .B(n2680), .Z(n2664) );
  NOR U2896 ( .A(n2657), .B(n2656), .Z(n2679) );
  XOR U2897 ( .A(n2681), .B(n2680), .Z(n2656) );
  AND U2898 ( .A(b[2]), .B(a[63]), .Z(n2681) );
  XOR U2899 ( .A(n2680), .B(n2683), .Z(n2682) );
  XNOR U2900 ( .A(n2684), .B(n2685), .Z(n2680) );
  NANDN U2901 ( .A(n2660), .B(n2659), .Z(n2685) );
  XOR U2902 ( .A(n2684), .B(n2686), .Z(n2659) );
  NAND U2903 ( .A(b[1]), .B(a[63]), .Z(n2686) );
  XOR U2904 ( .A(n2684), .B(n2688), .Z(n2687) );
  OR U2905 ( .A(n1292), .B(n1290), .Z(n2684) );
  XOR U2906 ( .A(n2690), .B(n2691), .Z(n1290) );
  NANDN U2907 ( .A(n187), .B(a[63]), .Z(n1292) );
  XNOR U2908 ( .A(n2693), .B(n2645), .Z(n2646) );
  XOR U2909 ( .A(n2694), .B(n2695), .Z(n2645) );
  ANDN U2910 ( .B(n2683), .A(n2692), .Z(n2694) );
  XNOR U2911 ( .A(n2696), .B(n2695), .Z(n2692) );
  AND U2912 ( .A(b[3]), .B(a[62]), .Z(n2696) );
  XOR U2913 ( .A(n2695), .B(n2678), .Z(n2697) );
  XOR U2914 ( .A(n2698), .B(n2699), .Z(n2678) );
  XOR U2915 ( .A(n2676), .B(n2700), .Z(n2699) );
  XNOR U2916 ( .A(n2701), .B(n2702), .Z(n2700) );
  XOR U2917 ( .A(n2703), .B(n2704), .Z(n2702) );
  NAND U2918 ( .A(b[6]), .B(a[59]), .Z(n2704) );
  AND U2919 ( .A(b[7]), .B(a[58]), .Z(n2703) );
  XNOR U2920 ( .A(n2705), .B(n2701), .Z(n2698) );
  XOR U2921 ( .A(n2706), .B(n2707), .Z(n2701) );
  NOR U2922 ( .A(n2708), .B(n2709), .Z(n2706) );
  AND U2923 ( .A(b[5]), .B(a[60]), .Z(n2705) );
  XNOR U2924 ( .A(n2710), .B(n2711), .Z(n2695) );
  ANDN U2925 ( .B(n2688), .A(n2689), .Z(n2710) );
  XOR U2926 ( .A(n2712), .B(n2711), .Z(n2689) );
  IV U2927 ( .A(n2713), .Z(n2711) );
  AND U2928 ( .A(b[2]), .B(a[62]), .Z(n2712) );
  XNOR U2929 ( .A(n2715), .B(n2713), .Z(n2714) );
  XOR U2930 ( .A(n2716), .B(n2717), .Z(n2713) );
  NANDN U2931 ( .A(n2691), .B(n2690), .Z(n2717) );
  XOR U2932 ( .A(n2716), .B(n2718), .Z(n2690) );
  NAND U2933 ( .A(b[1]), .B(a[62]), .Z(n2718) );
  XOR U2934 ( .A(n2716), .B(n2720), .Z(n2719) );
  OR U2935 ( .A(n1297), .B(n1295), .Z(n2716) );
  XOR U2936 ( .A(n2722), .B(n2723), .Z(n1295) );
  NANDN U2937 ( .A(n187), .B(a[62]), .Z(n1297) );
  XNOR U2938 ( .A(n2725), .B(n2676), .Z(n2677) );
  XNOR U2939 ( .A(n2726), .B(n2727), .Z(n2676) );
  ANDN U2940 ( .B(n2715), .A(n2724), .Z(n2726) );
  XOR U2941 ( .A(n2728), .B(n2727), .Z(n2724) );
  IV U2942 ( .A(n2729), .Z(n2727) );
  AND U2943 ( .A(b[3]), .B(a[61]), .Z(n2728) );
  XOR U2944 ( .A(n2709), .B(n2729), .Z(n2730) );
  XOR U2945 ( .A(n2731), .B(n2732), .Z(n2729) );
  ANDN U2946 ( .B(n2720), .A(n2721), .Z(n2731) );
  AND U2947 ( .A(b[2]), .B(a[61]), .Z(n2733) );
  XNOR U2948 ( .A(n2735), .B(n2732), .Z(n2734) );
  XOR U2949 ( .A(n2736), .B(n2737), .Z(n2732) );
  NANDN U2950 ( .A(n2723), .B(n2722), .Z(n2737) );
  XOR U2951 ( .A(n2736), .B(n2738), .Z(n2722) );
  NAND U2952 ( .A(b[1]), .B(a[61]), .Z(n2738) );
  XOR U2953 ( .A(n2736), .B(n2740), .Z(n2739) );
  OR U2954 ( .A(n1302), .B(n1300), .Z(n2736) );
  XOR U2955 ( .A(n2742), .B(n2743), .Z(n1300) );
  NANDN U2956 ( .A(n187), .B(a[61]), .Z(n1302) );
  XOR U2957 ( .A(n2745), .B(n2746), .Z(n2709) );
  XNOR U2958 ( .A(n2747), .B(n2748), .Z(n2746) );
  XNOR U2959 ( .A(n2749), .B(n2750), .Z(n2747) );
  XOR U2960 ( .A(n2751), .B(n2752), .Z(n2750) );
  AND U2961 ( .A(b[7]), .B(a[57]), .Z(n2752) );
  AND U2962 ( .A(b[6]), .B(a[58]), .Z(n2751) );
  XNOR U2963 ( .A(n2753), .B(n2749), .Z(n2745) );
  XOR U2964 ( .A(n2754), .B(n2755), .Z(n2749) );
  NOR U2965 ( .A(n2756), .B(n2757), .Z(n2754) );
  AND U2966 ( .A(b[5]), .B(a[59]), .Z(n2753) );
  XOR U2967 ( .A(n2758), .B(n2707), .Z(n2708) );
  IV U2968 ( .A(n2748), .Z(n2707) );
  XOR U2969 ( .A(n2759), .B(n2760), .Z(n2748) );
  ANDN U2970 ( .B(n2735), .A(n2744), .Z(n2759) );
  AND U2971 ( .A(b[3]), .B(a[60]), .Z(n2761) );
  XOR U2972 ( .A(n2757), .B(n2760), .Z(n2762) );
  XOR U2973 ( .A(n2763), .B(n2764), .Z(n2760) );
  ANDN U2974 ( .B(n2740), .A(n2741), .Z(n2763) );
  AND U2975 ( .A(b[2]), .B(a[60]), .Z(n2765) );
  XNOR U2976 ( .A(n2767), .B(n2764), .Z(n2766) );
  XOR U2977 ( .A(n2768), .B(n2769), .Z(n2764) );
  NANDN U2978 ( .A(n2743), .B(n2742), .Z(n2769) );
  XOR U2979 ( .A(n2768), .B(n2770), .Z(n2742) );
  NAND U2980 ( .A(b[1]), .B(a[60]), .Z(n2770) );
  XOR U2981 ( .A(n2768), .B(n2772), .Z(n2771) );
  OR U2982 ( .A(n1307), .B(n1305), .Z(n2768) );
  XOR U2983 ( .A(n2774), .B(n2775), .Z(n1305) );
  NANDN U2984 ( .A(n187), .B(a[60]), .Z(n1307) );
  XOR U2985 ( .A(n2777), .B(n2778), .Z(n2757) );
  XNOR U2986 ( .A(n2779), .B(n2780), .Z(n2778) );
  XNOR U2987 ( .A(n2781), .B(n2782), .Z(n2779) );
  XOR U2988 ( .A(n2783), .B(n2784), .Z(n2782) );
  AND U2989 ( .A(b[6]), .B(a[57]), .Z(n2784) );
  AND U2990 ( .A(b[7]), .B(a[56]), .Z(n2783) );
  XNOR U2991 ( .A(n2785), .B(n2781), .Z(n2777) );
  XOR U2992 ( .A(n2786), .B(n2787), .Z(n2781) );
  NOR U2993 ( .A(n2788), .B(n2789), .Z(n2786) );
  AND U2994 ( .A(b[5]), .B(a[58]), .Z(n2785) );
  XOR U2995 ( .A(n2790), .B(n2755), .Z(n2756) );
  IV U2996 ( .A(n2780), .Z(n2755) );
  XOR U2997 ( .A(n2791), .B(n2792), .Z(n2780) );
  ANDN U2998 ( .B(n2767), .A(n2776), .Z(n2791) );
  AND U2999 ( .A(b[3]), .B(a[59]), .Z(n2793) );
  XOR U3000 ( .A(n2789), .B(n2792), .Z(n2794) );
  XOR U3001 ( .A(n2795), .B(n2796), .Z(n2792) );
  ANDN U3002 ( .B(n2772), .A(n2773), .Z(n2795) );
  AND U3003 ( .A(b[2]), .B(a[59]), .Z(n2797) );
  XOR U3004 ( .A(n2799), .B(n2796), .Z(n2798) );
  XOR U3005 ( .A(n2800), .B(n2801), .Z(n2796) );
  NANDN U3006 ( .A(n2775), .B(n2774), .Z(n2801) );
  XOR U3007 ( .A(n2800), .B(n2802), .Z(n2774) );
  NAND U3008 ( .A(b[1]), .B(a[59]), .Z(n2802) );
  XOR U3009 ( .A(n2800), .B(n2804), .Z(n2803) );
  OR U3010 ( .A(n1312), .B(n1310), .Z(n2800) );
  XOR U3011 ( .A(n2806), .B(n2807), .Z(n1310) );
  NANDN U3012 ( .A(n187), .B(a[59]), .Z(n1312) );
  XOR U3013 ( .A(n2809), .B(n2810), .Z(n2789) );
  XNOR U3014 ( .A(n2811), .B(n2812), .Z(n2810) );
  XOR U3015 ( .A(n2813), .B(n2814), .Z(n2811) );
  AND U3016 ( .A(b[5]), .B(a[57]), .Z(n2813) );
  XOR U3017 ( .A(n2814), .B(n2815), .Z(n2809) );
  XOR U3018 ( .A(n2816), .B(n2817), .Z(n2815) );
  AND U3019 ( .A(b[6]), .B(a[56]), .Z(n2817) );
  AND U3020 ( .A(b[7]), .B(a[55]), .Z(n2816) );
  XOR U3021 ( .A(n2818), .B(n2819), .Z(n2814) );
  ANDN U3022 ( .B(n2820), .A(n2821), .Z(n2818) );
  XOR U3023 ( .A(n2822), .B(n2787), .Z(n2788) );
  IV U3024 ( .A(n2812), .Z(n2787) );
  XOR U3025 ( .A(n2823), .B(n2824), .Z(n2812) );
  NOR U3026 ( .A(n2808), .B(n2799), .Z(n2823) );
  XNOR U3027 ( .A(n2821), .B(n2825), .Z(n2799) );
  XNOR U3028 ( .A(n2820), .B(n2824), .Z(n2825) );
  XOR U3029 ( .A(n2826), .B(n2819), .Z(n2820) );
  AND U3030 ( .A(b[4]), .B(a[57]), .Z(n2826) );
  XOR U3031 ( .A(n2827), .B(n2828), .Z(n2821) );
  XOR U3032 ( .A(n2819), .B(n2829), .Z(n2828) );
  XOR U3033 ( .A(n2830), .B(n2831), .Z(n2829) );
  XOR U3034 ( .A(n2832), .B(n2833), .Z(n2831) );
  NAND U3035 ( .A(b[6]), .B(a[55]), .Z(n2833) );
  AND U3036 ( .A(b[7]), .B(a[54]), .Z(n2832) );
  XOR U3037 ( .A(n2834), .B(n2835), .Z(n2819) );
  ANDN U3038 ( .B(n2836), .A(n2837), .Z(n2834) );
  XOR U3039 ( .A(n2838), .B(n2830), .Z(n2827) );
  XOR U3040 ( .A(n2839), .B(n2840), .Z(n2830) );
  NOR U3041 ( .A(n2841), .B(n2842), .Z(n2839) );
  AND U3042 ( .A(b[5]), .B(a[56]), .Z(n2838) );
  XOR U3043 ( .A(n2844), .B(n2845), .Z(n2824) );
  ANDN U3044 ( .B(n2804), .A(n2805), .Z(n2844) );
  AND U3045 ( .A(b[2]), .B(a[58]), .Z(n2846) );
  XNOR U3046 ( .A(n2836), .B(n2845), .Z(n2847) );
  XOR U3047 ( .A(n2848), .B(n2849), .Z(n2845) );
  NANDN U3048 ( .A(n2807), .B(n2806), .Z(n2849) );
  XOR U3049 ( .A(n2848), .B(n2850), .Z(n2806) );
  NAND U3050 ( .A(b[1]), .B(a[58]), .Z(n2850) );
  XNOR U3051 ( .A(n2848), .B(n2852), .Z(n2851) );
  OR U3052 ( .A(n1317), .B(n1315), .Z(n2848) );
  NANDN U3053 ( .A(n187), .B(a[58]), .Z(n1317) );
  XOR U3054 ( .A(n2856), .B(n2835), .Z(n2836) );
  AND U3055 ( .A(b[3]), .B(a[57]), .Z(n2856) );
  XOR U3056 ( .A(n2835), .B(n2842), .Z(n2857) );
  XOR U3057 ( .A(n2858), .B(n2859), .Z(n2842) );
  XOR U3058 ( .A(n2840), .B(n2860), .Z(n2859) );
  XOR U3059 ( .A(n2861), .B(n2862), .Z(n2860) );
  XOR U3060 ( .A(n2863), .B(n2864), .Z(n2862) );
  NAND U3061 ( .A(b[6]), .B(a[54]), .Z(n2864) );
  AND U3062 ( .A(b[7]), .B(a[53]), .Z(n2863) );
  XOR U3063 ( .A(n2865), .B(n2861), .Z(n2858) );
  XOR U3064 ( .A(n2866), .B(n2867), .Z(n2861) );
  NOR U3065 ( .A(n2868), .B(n2869), .Z(n2866) );
  AND U3066 ( .A(b[5]), .B(a[55]), .Z(n2865) );
  XNOR U3067 ( .A(n2870), .B(n2871), .Z(n2835) );
  NOR U3068 ( .A(n2853), .B(n2852), .Z(n2870) );
  XOR U3069 ( .A(n2872), .B(n2871), .Z(n2852) );
  AND U3070 ( .A(b[2]), .B(a[57]), .Z(n2872) );
  XOR U3071 ( .A(n2871), .B(n2874), .Z(n2873) );
  XNOR U3072 ( .A(n2875), .B(n2876), .Z(n2871) );
  OR U3073 ( .A(n2854), .B(n2855), .Z(n2876) );
  XNOR U3074 ( .A(n2875), .B(n2878), .Z(n2877) );
  XNOR U3075 ( .A(n2875), .B(n2880), .Z(n2854) );
  NAND U3076 ( .A(b[1]), .B(a[57]), .Z(n2880) );
  OR U3077 ( .A(n1322), .B(n1320), .Z(n2875) );
  XOR U3078 ( .A(n2881), .B(n2882), .Z(n1320) );
  NANDN U3079 ( .A(n187), .B(a[57]), .Z(n1322) );
  XNOR U3080 ( .A(n2884), .B(n2840), .Z(n2841) );
  XOR U3081 ( .A(n2885), .B(n2886), .Z(n2840) );
  ANDN U3082 ( .B(n2874), .A(n2883), .Z(n2885) );
  XNOR U3083 ( .A(n2887), .B(n2886), .Z(n2883) );
  AND U3084 ( .A(b[3]), .B(a[56]), .Z(n2887) );
  XOR U3085 ( .A(n2886), .B(n2869), .Z(n2888) );
  XOR U3086 ( .A(n2889), .B(n2890), .Z(n2869) );
  XOR U3087 ( .A(n2867), .B(n2891), .Z(n2890) );
  XOR U3088 ( .A(n2892), .B(n2893), .Z(n2891) );
  XOR U3089 ( .A(n2894), .B(n2895), .Z(n2893) );
  NAND U3090 ( .A(b[6]), .B(a[53]), .Z(n2895) );
  AND U3091 ( .A(b[7]), .B(a[52]), .Z(n2894) );
  XOR U3092 ( .A(n2896), .B(n2892), .Z(n2889) );
  XOR U3093 ( .A(n2897), .B(n2898), .Z(n2892) );
  NOR U3094 ( .A(n2899), .B(n2900), .Z(n2897) );
  AND U3095 ( .A(b[5]), .B(a[54]), .Z(n2896) );
  XNOR U3096 ( .A(n2901), .B(n2902), .Z(n2886) );
  NOR U3097 ( .A(n2879), .B(n2878), .Z(n2901) );
  XOR U3098 ( .A(n2903), .B(n2902), .Z(n2878) );
  AND U3099 ( .A(b[2]), .B(a[56]), .Z(n2903) );
  XOR U3100 ( .A(n2902), .B(n2905), .Z(n2904) );
  XNOR U3101 ( .A(n2906), .B(n2907), .Z(n2902) );
  NANDN U3102 ( .A(n2882), .B(n2881), .Z(n2907) );
  XOR U3103 ( .A(n2906), .B(n2908), .Z(n2881) );
  NAND U3104 ( .A(b[1]), .B(a[56]), .Z(n2908) );
  XOR U3105 ( .A(n2906), .B(n2910), .Z(n2909) );
  OR U3106 ( .A(n1327), .B(n1325), .Z(n2906) );
  XOR U3107 ( .A(n2912), .B(n2913), .Z(n1325) );
  NANDN U3108 ( .A(n187), .B(a[56]), .Z(n1327) );
  XNOR U3109 ( .A(n2915), .B(n2867), .Z(n2868) );
  XOR U3110 ( .A(n2916), .B(n2917), .Z(n2867) );
  ANDN U3111 ( .B(n2905), .A(n2914), .Z(n2916) );
  XNOR U3112 ( .A(n2918), .B(n2917), .Z(n2914) );
  AND U3113 ( .A(b[3]), .B(a[55]), .Z(n2918) );
  XOR U3114 ( .A(n2917), .B(n2900), .Z(n2919) );
  XOR U3115 ( .A(n2920), .B(n2921), .Z(n2900) );
  XOR U3116 ( .A(n2898), .B(n2922), .Z(n2921) );
  XNOR U3117 ( .A(n2923), .B(n2924), .Z(n2922) );
  XOR U3118 ( .A(n2925), .B(n2926), .Z(n2924) );
  NAND U3119 ( .A(b[6]), .B(a[52]), .Z(n2926) );
  AND U3120 ( .A(b[7]), .B(a[51]), .Z(n2925) );
  XNOR U3121 ( .A(n2927), .B(n2923), .Z(n2920) );
  XOR U3122 ( .A(n2928), .B(n2929), .Z(n2923) );
  NOR U3123 ( .A(n2930), .B(n2931), .Z(n2928) );
  AND U3124 ( .A(b[5]), .B(a[53]), .Z(n2927) );
  XNOR U3125 ( .A(n2932), .B(n2933), .Z(n2917) );
  ANDN U3126 ( .B(n2910), .A(n2911), .Z(n2932) );
  XOR U3127 ( .A(n2934), .B(n2933), .Z(n2911) );
  IV U3128 ( .A(n2935), .Z(n2933) );
  AND U3129 ( .A(b[2]), .B(a[55]), .Z(n2934) );
  XNOR U3130 ( .A(n2937), .B(n2935), .Z(n2936) );
  XOR U3131 ( .A(n2938), .B(n2939), .Z(n2935) );
  NANDN U3132 ( .A(n2913), .B(n2912), .Z(n2939) );
  XOR U3133 ( .A(n2938), .B(n2940), .Z(n2912) );
  NAND U3134 ( .A(b[1]), .B(a[55]), .Z(n2940) );
  XOR U3135 ( .A(n2938), .B(n2942), .Z(n2941) );
  OR U3136 ( .A(n1332), .B(n1330), .Z(n2938) );
  XOR U3137 ( .A(n2944), .B(n2945), .Z(n1330) );
  NANDN U3138 ( .A(n187), .B(a[55]), .Z(n1332) );
  XNOR U3139 ( .A(n2947), .B(n2898), .Z(n2899) );
  XNOR U3140 ( .A(n2948), .B(n2949), .Z(n2898) );
  ANDN U3141 ( .B(n2937), .A(n2946), .Z(n2948) );
  XOR U3142 ( .A(n2950), .B(n2949), .Z(n2946) );
  IV U3143 ( .A(n2951), .Z(n2949) );
  AND U3144 ( .A(b[3]), .B(a[54]), .Z(n2950) );
  XOR U3145 ( .A(n2931), .B(n2951), .Z(n2952) );
  XOR U3146 ( .A(n2953), .B(n2954), .Z(n2951) );
  ANDN U3147 ( .B(n2942), .A(n2943), .Z(n2953) );
  AND U3148 ( .A(b[2]), .B(a[54]), .Z(n2955) );
  XNOR U3149 ( .A(n2957), .B(n2954), .Z(n2956) );
  XOR U3150 ( .A(n2958), .B(n2959), .Z(n2954) );
  NANDN U3151 ( .A(n2945), .B(n2944), .Z(n2959) );
  XOR U3152 ( .A(n2958), .B(n2960), .Z(n2944) );
  NAND U3153 ( .A(b[1]), .B(a[54]), .Z(n2960) );
  XOR U3154 ( .A(n2958), .B(n2962), .Z(n2961) );
  OR U3155 ( .A(n1337), .B(n1335), .Z(n2958) );
  XOR U3156 ( .A(n2964), .B(n2965), .Z(n1335) );
  NANDN U3157 ( .A(n187), .B(a[54]), .Z(n1337) );
  XOR U3158 ( .A(n2967), .B(n2968), .Z(n2931) );
  XNOR U3159 ( .A(n2969), .B(n2970), .Z(n2968) );
  XNOR U3160 ( .A(n2971), .B(n2972), .Z(n2969) );
  XOR U3161 ( .A(n2973), .B(n2974), .Z(n2972) );
  AND U3162 ( .A(b[7]), .B(a[50]), .Z(n2974) );
  AND U3163 ( .A(b[6]), .B(a[51]), .Z(n2973) );
  XNOR U3164 ( .A(n2975), .B(n2971), .Z(n2967) );
  XOR U3165 ( .A(n2976), .B(n2977), .Z(n2971) );
  NOR U3166 ( .A(n2978), .B(n2979), .Z(n2976) );
  AND U3167 ( .A(b[5]), .B(a[52]), .Z(n2975) );
  XOR U3168 ( .A(n2980), .B(n2929), .Z(n2930) );
  IV U3169 ( .A(n2970), .Z(n2929) );
  XOR U3170 ( .A(n2981), .B(n2982), .Z(n2970) );
  ANDN U3171 ( .B(n2957), .A(n2966), .Z(n2981) );
  AND U3172 ( .A(b[3]), .B(a[53]), .Z(n2983) );
  XOR U3173 ( .A(n2979), .B(n2982), .Z(n2984) );
  XOR U3174 ( .A(n2985), .B(n2986), .Z(n2982) );
  ANDN U3175 ( .B(n2962), .A(n2963), .Z(n2985) );
  AND U3176 ( .A(b[2]), .B(a[53]), .Z(n2987) );
  XNOR U3177 ( .A(n2989), .B(n2986), .Z(n2988) );
  XOR U3178 ( .A(n2990), .B(n2991), .Z(n2986) );
  NANDN U3179 ( .A(n2965), .B(n2964), .Z(n2991) );
  XOR U3180 ( .A(n2990), .B(n2992), .Z(n2964) );
  NAND U3181 ( .A(b[1]), .B(a[53]), .Z(n2992) );
  XOR U3182 ( .A(n2990), .B(n2994), .Z(n2993) );
  OR U3183 ( .A(n1342), .B(n1340), .Z(n2990) );
  XOR U3184 ( .A(n2996), .B(n2997), .Z(n1340) );
  NANDN U3185 ( .A(n187), .B(a[53]), .Z(n1342) );
  XOR U3186 ( .A(n2999), .B(n3000), .Z(n2979) );
  XNOR U3187 ( .A(n3001), .B(n3002), .Z(n3000) );
  XNOR U3188 ( .A(n3003), .B(n3004), .Z(n3001) );
  XOR U3189 ( .A(n3005), .B(n3006), .Z(n3004) );
  AND U3190 ( .A(b[6]), .B(a[50]), .Z(n3006) );
  AND U3191 ( .A(b[7]), .B(a[49]), .Z(n3005) );
  XNOR U3192 ( .A(n3007), .B(n3003), .Z(n2999) );
  XOR U3193 ( .A(n3008), .B(n3009), .Z(n3003) );
  NOR U3194 ( .A(n3010), .B(n3011), .Z(n3008) );
  AND U3195 ( .A(b[5]), .B(a[51]), .Z(n3007) );
  XOR U3196 ( .A(n3012), .B(n2977), .Z(n2978) );
  IV U3197 ( .A(n3002), .Z(n2977) );
  XOR U3198 ( .A(n3013), .B(n3014), .Z(n3002) );
  ANDN U3199 ( .B(n2989), .A(n2998), .Z(n3013) );
  AND U3200 ( .A(b[3]), .B(a[52]), .Z(n3015) );
  XOR U3201 ( .A(n3011), .B(n3014), .Z(n3016) );
  XOR U3202 ( .A(n3017), .B(n3018), .Z(n3014) );
  ANDN U3203 ( .B(n2994), .A(n2995), .Z(n3017) );
  AND U3204 ( .A(b[2]), .B(a[52]), .Z(n3019) );
  XOR U3205 ( .A(n3021), .B(n3018), .Z(n3020) );
  XOR U3206 ( .A(n3022), .B(n3023), .Z(n3018) );
  NANDN U3207 ( .A(n2997), .B(n2996), .Z(n3023) );
  XOR U3208 ( .A(n3022), .B(n3024), .Z(n2996) );
  NAND U3209 ( .A(b[1]), .B(a[52]), .Z(n3024) );
  XOR U3210 ( .A(n3022), .B(n3026), .Z(n3025) );
  OR U3211 ( .A(n1347), .B(n1345), .Z(n3022) );
  XOR U3212 ( .A(n3028), .B(n3029), .Z(n1345) );
  NANDN U3213 ( .A(n187), .B(a[52]), .Z(n1347) );
  XOR U3214 ( .A(n3031), .B(n3032), .Z(n3011) );
  XNOR U3215 ( .A(n3033), .B(n3034), .Z(n3032) );
  XOR U3216 ( .A(n3035), .B(n3036), .Z(n3033) );
  AND U3217 ( .A(b[5]), .B(a[50]), .Z(n3035) );
  XOR U3218 ( .A(n3036), .B(n3037), .Z(n3031) );
  XOR U3219 ( .A(n3038), .B(n3039), .Z(n3037) );
  AND U3220 ( .A(b[6]), .B(a[49]), .Z(n3039) );
  AND U3221 ( .A(b[7]), .B(a[48]), .Z(n3038) );
  XOR U3222 ( .A(n3040), .B(n3041), .Z(n3036) );
  ANDN U3223 ( .B(n3042), .A(n3043), .Z(n3040) );
  XOR U3224 ( .A(n3044), .B(n3009), .Z(n3010) );
  IV U3225 ( .A(n3034), .Z(n3009) );
  XOR U3226 ( .A(n3045), .B(n3046), .Z(n3034) );
  NOR U3227 ( .A(n3030), .B(n3021), .Z(n3045) );
  XNOR U3228 ( .A(n3043), .B(n3047), .Z(n3021) );
  XNOR U3229 ( .A(n3042), .B(n3046), .Z(n3047) );
  XOR U3230 ( .A(n3048), .B(n3041), .Z(n3042) );
  AND U3231 ( .A(b[4]), .B(a[50]), .Z(n3048) );
  XOR U3232 ( .A(n3049), .B(n3050), .Z(n3043) );
  XOR U3233 ( .A(n3041), .B(n3051), .Z(n3050) );
  XOR U3234 ( .A(n3052), .B(n3053), .Z(n3051) );
  XOR U3235 ( .A(n3054), .B(n3055), .Z(n3053) );
  NAND U3236 ( .A(b[6]), .B(a[48]), .Z(n3055) );
  AND U3237 ( .A(b[7]), .B(a[47]), .Z(n3054) );
  XOR U3238 ( .A(n3056), .B(n3057), .Z(n3041) );
  ANDN U3239 ( .B(n3058), .A(n3059), .Z(n3056) );
  XOR U3240 ( .A(n3060), .B(n3052), .Z(n3049) );
  XOR U3241 ( .A(n3061), .B(n3062), .Z(n3052) );
  NOR U3242 ( .A(n3063), .B(n3064), .Z(n3061) );
  AND U3243 ( .A(b[5]), .B(a[49]), .Z(n3060) );
  XOR U3244 ( .A(n3066), .B(n3067), .Z(n3046) );
  ANDN U3245 ( .B(n3026), .A(n3027), .Z(n3066) );
  AND U3246 ( .A(b[2]), .B(a[51]), .Z(n3068) );
  XNOR U3247 ( .A(n3058), .B(n3067), .Z(n3069) );
  XOR U3248 ( .A(n3070), .B(n3071), .Z(n3067) );
  NANDN U3249 ( .A(n3029), .B(n3028), .Z(n3071) );
  XOR U3250 ( .A(n3070), .B(n3072), .Z(n3028) );
  NAND U3251 ( .A(b[1]), .B(a[51]), .Z(n3072) );
  XNOR U3252 ( .A(n3070), .B(n3074), .Z(n3073) );
  OR U3253 ( .A(n1352), .B(n1350), .Z(n3070) );
  NANDN U3254 ( .A(n187), .B(a[51]), .Z(n1352) );
  XOR U3255 ( .A(n3078), .B(n3057), .Z(n3058) );
  AND U3256 ( .A(b[3]), .B(a[50]), .Z(n3078) );
  XOR U3257 ( .A(n3057), .B(n3064), .Z(n3079) );
  XOR U3258 ( .A(n3080), .B(n3081), .Z(n3064) );
  XOR U3259 ( .A(n3062), .B(n3082), .Z(n3081) );
  XOR U3260 ( .A(n3083), .B(n3084), .Z(n3082) );
  XOR U3261 ( .A(n3085), .B(n3086), .Z(n3084) );
  NAND U3262 ( .A(b[6]), .B(a[47]), .Z(n3086) );
  AND U3263 ( .A(b[7]), .B(a[46]), .Z(n3085) );
  XOR U3264 ( .A(n3087), .B(n3083), .Z(n3080) );
  XOR U3265 ( .A(n3088), .B(n3089), .Z(n3083) );
  NOR U3266 ( .A(n3090), .B(n3091), .Z(n3088) );
  AND U3267 ( .A(b[5]), .B(a[48]), .Z(n3087) );
  XNOR U3268 ( .A(n3092), .B(n3093), .Z(n3057) );
  NOR U3269 ( .A(n3075), .B(n3074), .Z(n3092) );
  XOR U3270 ( .A(n3094), .B(n3093), .Z(n3074) );
  AND U3271 ( .A(b[2]), .B(a[50]), .Z(n3094) );
  XOR U3272 ( .A(n3093), .B(n3096), .Z(n3095) );
  XNOR U3273 ( .A(n3097), .B(n3098), .Z(n3093) );
  OR U3274 ( .A(n3076), .B(n3077), .Z(n3098) );
  XNOR U3275 ( .A(n3097), .B(n3100), .Z(n3099) );
  XNOR U3276 ( .A(n3097), .B(n3102), .Z(n3076) );
  NAND U3277 ( .A(b[1]), .B(a[50]), .Z(n3102) );
  OR U3278 ( .A(n1357), .B(n1355), .Z(n3097) );
  XOR U3279 ( .A(n3103), .B(n3104), .Z(n1355) );
  NANDN U3280 ( .A(n187), .B(a[50]), .Z(n1357) );
  XNOR U3281 ( .A(n3106), .B(n3062), .Z(n3063) );
  XOR U3282 ( .A(n3107), .B(n3108), .Z(n3062) );
  ANDN U3283 ( .B(n3096), .A(n3105), .Z(n3107) );
  XNOR U3284 ( .A(n3109), .B(n3108), .Z(n3105) );
  AND U3285 ( .A(b[3]), .B(a[49]), .Z(n3109) );
  XOR U3286 ( .A(n3108), .B(n3091), .Z(n3110) );
  XOR U3287 ( .A(n3111), .B(n3112), .Z(n3091) );
  XOR U3288 ( .A(n3089), .B(n3113), .Z(n3112) );
  XOR U3289 ( .A(n3114), .B(n3115), .Z(n3113) );
  XOR U3290 ( .A(n3116), .B(n3117), .Z(n3115) );
  NAND U3291 ( .A(b[6]), .B(a[46]), .Z(n3117) );
  AND U3292 ( .A(b[7]), .B(a[45]), .Z(n3116) );
  XOR U3293 ( .A(n3118), .B(n3114), .Z(n3111) );
  XOR U3294 ( .A(n3119), .B(n3120), .Z(n3114) );
  NOR U3295 ( .A(n3121), .B(n3122), .Z(n3119) );
  AND U3296 ( .A(b[5]), .B(a[47]), .Z(n3118) );
  XNOR U3297 ( .A(n3123), .B(n3124), .Z(n3108) );
  NOR U3298 ( .A(n3101), .B(n3100), .Z(n3123) );
  XOR U3299 ( .A(n3125), .B(n3124), .Z(n3100) );
  AND U3300 ( .A(b[2]), .B(a[49]), .Z(n3125) );
  XOR U3301 ( .A(n3124), .B(n3127), .Z(n3126) );
  XNOR U3302 ( .A(n3128), .B(n3129), .Z(n3124) );
  NANDN U3303 ( .A(n3104), .B(n3103), .Z(n3129) );
  XOR U3304 ( .A(n3128), .B(n3130), .Z(n3103) );
  NAND U3305 ( .A(b[1]), .B(a[49]), .Z(n3130) );
  XOR U3306 ( .A(n3128), .B(n3132), .Z(n3131) );
  OR U3307 ( .A(n1362), .B(n1360), .Z(n3128) );
  XOR U3308 ( .A(n3134), .B(n3135), .Z(n1360) );
  NANDN U3309 ( .A(n187), .B(a[49]), .Z(n1362) );
  XNOR U3310 ( .A(n3137), .B(n3089), .Z(n3090) );
  XOR U3311 ( .A(n3138), .B(n3139), .Z(n3089) );
  ANDN U3312 ( .B(n3127), .A(n3136), .Z(n3138) );
  XNOR U3313 ( .A(n3140), .B(n3139), .Z(n3136) );
  AND U3314 ( .A(b[3]), .B(a[48]), .Z(n3140) );
  XOR U3315 ( .A(n3139), .B(n3122), .Z(n3141) );
  XOR U3316 ( .A(n3142), .B(n3143), .Z(n3122) );
  XOR U3317 ( .A(n3120), .B(n3144), .Z(n3143) );
  XNOR U3318 ( .A(n3145), .B(n3146), .Z(n3144) );
  XOR U3319 ( .A(n3147), .B(n3148), .Z(n3146) );
  NAND U3320 ( .A(b[6]), .B(a[45]), .Z(n3148) );
  AND U3321 ( .A(b[7]), .B(a[44]), .Z(n3147) );
  XNOR U3322 ( .A(n3149), .B(n3145), .Z(n3142) );
  XOR U3323 ( .A(n3150), .B(n3151), .Z(n3145) );
  NOR U3324 ( .A(n3152), .B(n3153), .Z(n3150) );
  AND U3325 ( .A(b[5]), .B(a[46]), .Z(n3149) );
  XNOR U3326 ( .A(n3154), .B(n3155), .Z(n3139) );
  ANDN U3327 ( .B(n3132), .A(n3133), .Z(n3154) );
  XOR U3328 ( .A(n3156), .B(n3155), .Z(n3133) );
  IV U3329 ( .A(n3157), .Z(n3155) );
  AND U3330 ( .A(b[2]), .B(a[48]), .Z(n3156) );
  XNOR U3331 ( .A(n3159), .B(n3157), .Z(n3158) );
  XOR U3332 ( .A(n3160), .B(n3161), .Z(n3157) );
  NANDN U3333 ( .A(n3135), .B(n3134), .Z(n3161) );
  XOR U3334 ( .A(n3160), .B(n3162), .Z(n3134) );
  NAND U3335 ( .A(b[1]), .B(a[48]), .Z(n3162) );
  XOR U3336 ( .A(n3160), .B(n3164), .Z(n3163) );
  OR U3337 ( .A(n1367), .B(n1365), .Z(n3160) );
  XOR U3338 ( .A(n3166), .B(n3167), .Z(n1365) );
  NANDN U3339 ( .A(n187), .B(a[48]), .Z(n1367) );
  XNOR U3340 ( .A(n3169), .B(n3120), .Z(n3121) );
  XNOR U3341 ( .A(n3170), .B(n3171), .Z(n3120) );
  ANDN U3342 ( .B(n3159), .A(n3168), .Z(n3170) );
  XOR U3343 ( .A(n3172), .B(n3171), .Z(n3168) );
  IV U3344 ( .A(n3173), .Z(n3171) );
  AND U3345 ( .A(b[3]), .B(a[47]), .Z(n3172) );
  XOR U3346 ( .A(n3153), .B(n3173), .Z(n3174) );
  XOR U3347 ( .A(n3175), .B(n3176), .Z(n3173) );
  ANDN U3348 ( .B(n3164), .A(n3165), .Z(n3175) );
  AND U3349 ( .A(b[2]), .B(a[47]), .Z(n3177) );
  XNOR U3350 ( .A(n3179), .B(n3176), .Z(n3178) );
  XOR U3351 ( .A(n3180), .B(n3181), .Z(n3176) );
  NANDN U3352 ( .A(n3167), .B(n3166), .Z(n3181) );
  XOR U3353 ( .A(n3180), .B(n3182), .Z(n3166) );
  NAND U3354 ( .A(b[1]), .B(a[47]), .Z(n3182) );
  XOR U3355 ( .A(n3180), .B(n3184), .Z(n3183) );
  OR U3356 ( .A(n1372), .B(n1370), .Z(n3180) );
  XOR U3357 ( .A(n3186), .B(n3187), .Z(n1370) );
  NANDN U3358 ( .A(n187), .B(a[47]), .Z(n1372) );
  XOR U3359 ( .A(n3189), .B(n3190), .Z(n3153) );
  XNOR U3360 ( .A(n3191), .B(n3192), .Z(n3190) );
  XNOR U3361 ( .A(n3193), .B(n3194), .Z(n3191) );
  XOR U3362 ( .A(n3195), .B(n3196), .Z(n3194) );
  AND U3363 ( .A(b[7]), .B(a[43]), .Z(n3196) );
  AND U3364 ( .A(b[6]), .B(a[44]), .Z(n3195) );
  XNOR U3365 ( .A(n3197), .B(n3193), .Z(n3189) );
  XOR U3366 ( .A(n3198), .B(n3199), .Z(n3193) );
  NOR U3367 ( .A(n3200), .B(n3201), .Z(n3198) );
  AND U3368 ( .A(b[5]), .B(a[45]), .Z(n3197) );
  XOR U3369 ( .A(n3202), .B(n3151), .Z(n3152) );
  IV U3370 ( .A(n3192), .Z(n3151) );
  XOR U3371 ( .A(n3203), .B(n3204), .Z(n3192) );
  ANDN U3372 ( .B(n3179), .A(n3188), .Z(n3203) );
  AND U3373 ( .A(b[3]), .B(a[46]), .Z(n3205) );
  XOR U3374 ( .A(n3201), .B(n3204), .Z(n3206) );
  XOR U3375 ( .A(n3207), .B(n3208), .Z(n3204) );
  ANDN U3376 ( .B(n3184), .A(n3185), .Z(n3207) );
  AND U3377 ( .A(b[2]), .B(a[46]), .Z(n3209) );
  XNOR U3378 ( .A(n3211), .B(n3208), .Z(n3210) );
  XOR U3379 ( .A(n3212), .B(n3213), .Z(n3208) );
  NANDN U3380 ( .A(n3187), .B(n3186), .Z(n3213) );
  XOR U3381 ( .A(n3212), .B(n3214), .Z(n3186) );
  NAND U3382 ( .A(b[1]), .B(a[46]), .Z(n3214) );
  XOR U3383 ( .A(n3212), .B(n3216), .Z(n3215) );
  OR U3384 ( .A(n1377), .B(n1375), .Z(n3212) );
  XOR U3385 ( .A(n3218), .B(n3219), .Z(n1375) );
  NANDN U3386 ( .A(n187), .B(a[46]), .Z(n1377) );
  XOR U3387 ( .A(n3221), .B(n3222), .Z(n3201) );
  XNOR U3388 ( .A(n3223), .B(n3224), .Z(n3222) );
  XNOR U3389 ( .A(n3225), .B(n3226), .Z(n3223) );
  XOR U3390 ( .A(n3227), .B(n3228), .Z(n3226) );
  AND U3391 ( .A(b[6]), .B(a[43]), .Z(n3228) );
  AND U3392 ( .A(b[7]), .B(a[42]), .Z(n3227) );
  XNOR U3393 ( .A(n3229), .B(n3225), .Z(n3221) );
  XOR U3394 ( .A(n3230), .B(n3231), .Z(n3225) );
  NOR U3395 ( .A(n3232), .B(n3233), .Z(n3230) );
  AND U3396 ( .A(b[5]), .B(a[44]), .Z(n3229) );
  XOR U3397 ( .A(n3234), .B(n3199), .Z(n3200) );
  IV U3398 ( .A(n3224), .Z(n3199) );
  XOR U3399 ( .A(n3235), .B(n3236), .Z(n3224) );
  ANDN U3400 ( .B(n3211), .A(n3220), .Z(n3235) );
  AND U3401 ( .A(b[3]), .B(a[45]), .Z(n3237) );
  XOR U3402 ( .A(n3233), .B(n3236), .Z(n3238) );
  XOR U3403 ( .A(n3239), .B(n3240), .Z(n3236) );
  ANDN U3404 ( .B(n3216), .A(n3217), .Z(n3239) );
  AND U3405 ( .A(b[2]), .B(a[45]), .Z(n3241) );
  XOR U3406 ( .A(n3243), .B(n3240), .Z(n3242) );
  XOR U3407 ( .A(n3244), .B(n3245), .Z(n3240) );
  NANDN U3408 ( .A(n3219), .B(n3218), .Z(n3245) );
  XOR U3409 ( .A(n3244), .B(n3246), .Z(n3218) );
  NAND U3410 ( .A(b[1]), .B(a[45]), .Z(n3246) );
  XOR U3411 ( .A(n3244), .B(n3248), .Z(n3247) );
  OR U3412 ( .A(n1382), .B(n1380), .Z(n3244) );
  XOR U3413 ( .A(n3250), .B(n3251), .Z(n1380) );
  NANDN U3414 ( .A(n187), .B(a[45]), .Z(n1382) );
  XOR U3415 ( .A(n3253), .B(n3254), .Z(n3233) );
  XNOR U3416 ( .A(n3255), .B(n3256), .Z(n3254) );
  XOR U3417 ( .A(n3257), .B(n3258), .Z(n3255) );
  AND U3418 ( .A(b[5]), .B(a[43]), .Z(n3257) );
  XOR U3419 ( .A(n3258), .B(n3259), .Z(n3253) );
  XOR U3420 ( .A(n3260), .B(n3261), .Z(n3259) );
  AND U3421 ( .A(b[6]), .B(a[42]), .Z(n3261) );
  AND U3422 ( .A(b[7]), .B(a[41]), .Z(n3260) );
  XOR U3423 ( .A(n3262), .B(n3263), .Z(n3258) );
  ANDN U3424 ( .B(n3264), .A(n3265), .Z(n3262) );
  XOR U3425 ( .A(n3266), .B(n3231), .Z(n3232) );
  IV U3426 ( .A(n3256), .Z(n3231) );
  XOR U3427 ( .A(n3267), .B(n3268), .Z(n3256) );
  NOR U3428 ( .A(n3252), .B(n3243), .Z(n3267) );
  XNOR U3429 ( .A(n3265), .B(n3269), .Z(n3243) );
  XNOR U3430 ( .A(n3264), .B(n3268), .Z(n3269) );
  XOR U3431 ( .A(n3270), .B(n3263), .Z(n3264) );
  AND U3432 ( .A(b[4]), .B(a[43]), .Z(n3270) );
  XOR U3433 ( .A(n3271), .B(n3272), .Z(n3265) );
  XOR U3434 ( .A(n3263), .B(n3273), .Z(n3272) );
  XOR U3435 ( .A(n3274), .B(n3275), .Z(n3273) );
  XOR U3436 ( .A(n3276), .B(n3277), .Z(n3275) );
  NAND U3437 ( .A(b[6]), .B(a[41]), .Z(n3277) );
  AND U3438 ( .A(b[7]), .B(a[40]), .Z(n3276) );
  XOR U3439 ( .A(n3278), .B(n3279), .Z(n3263) );
  ANDN U3440 ( .B(n3280), .A(n3281), .Z(n3278) );
  XOR U3441 ( .A(n3282), .B(n3274), .Z(n3271) );
  XOR U3442 ( .A(n3283), .B(n3284), .Z(n3274) );
  NOR U3443 ( .A(n3285), .B(n3286), .Z(n3283) );
  AND U3444 ( .A(b[5]), .B(a[42]), .Z(n3282) );
  XOR U3445 ( .A(n3288), .B(n3289), .Z(n3268) );
  ANDN U3446 ( .B(n3248), .A(n3249), .Z(n3288) );
  AND U3447 ( .A(b[2]), .B(a[44]), .Z(n3290) );
  XNOR U3448 ( .A(n3280), .B(n3289), .Z(n3291) );
  XOR U3449 ( .A(n3292), .B(n3293), .Z(n3289) );
  NANDN U3450 ( .A(n3251), .B(n3250), .Z(n3293) );
  XOR U3451 ( .A(n3292), .B(n3294), .Z(n3250) );
  NAND U3452 ( .A(b[1]), .B(a[44]), .Z(n3294) );
  XNOR U3453 ( .A(n3292), .B(n3296), .Z(n3295) );
  OR U3454 ( .A(n1387), .B(n1385), .Z(n3292) );
  NANDN U3455 ( .A(n187), .B(a[44]), .Z(n1387) );
  XOR U3456 ( .A(n3300), .B(n3279), .Z(n3280) );
  AND U3457 ( .A(b[3]), .B(a[43]), .Z(n3300) );
  XOR U3458 ( .A(n3279), .B(n3286), .Z(n3301) );
  XOR U3459 ( .A(n3302), .B(n3303), .Z(n3286) );
  XOR U3460 ( .A(n3284), .B(n3304), .Z(n3303) );
  XOR U3461 ( .A(n3305), .B(n3306), .Z(n3304) );
  XOR U3462 ( .A(n3307), .B(n3308), .Z(n3306) );
  NAND U3463 ( .A(b[6]), .B(a[40]), .Z(n3308) );
  AND U3464 ( .A(b[7]), .B(a[39]), .Z(n3307) );
  XOR U3465 ( .A(n3309), .B(n3305), .Z(n3302) );
  XOR U3466 ( .A(n3310), .B(n3311), .Z(n3305) );
  NOR U3467 ( .A(n3312), .B(n3313), .Z(n3310) );
  AND U3468 ( .A(b[5]), .B(a[41]), .Z(n3309) );
  XNOR U3469 ( .A(n3314), .B(n3315), .Z(n3279) );
  NOR U3470 ( .A(n3297), .B(n3296), .Z(n3314) );
  XOR U3471 ( .A(n3316), .B(n3315), .Z(n3296) );
  AND U3472 ( .A(b[2]), .B(a[43]), .Z(n3316) );
  XOR U3473 ( .A(n3315), .B(n3318), .Z(n3317) );
  XNOR U3474 ( .A(n3319), .B(n3320), .Z(n3315) );
  OR U3475 ( .A(n3298), .B(n3299), .Z(n3320) );
  XNOR U3476 ( .A(n3319), .B(n3322), .Z(n3321) );
  XNOR U3477 ( .A(n3319), .B(n3324), .Z(n3298) );
  NAND U3478 ( .A(b[1]), .B(a[43]), .Z(n3324) );
  OR U3479 ( .A(n1392), .B(n1390), .Z(n3319) );
  XOR U3480 ( .A(n3325), .B(n3326), .Z(n1390) );
  NANDN U3481 ( .A(n187), .B(a[43]), .Z(n1392) );
  XNOR U3482 ( .A(n3328), .B(n3284), .Z(n3285) );
  XOR U3483 ( .A(n3329), .B(n3330), .Z(n3284) );
  ANDN U3484 ( .B(n3318), .A(n3327), .Z(n3329) );
  XNOR U3485 ( .A(n3331), .B(n3330), .Z(n3327) );
  AND U3486 ( .A(b[3]), .B(a[42]), .Z(n3331) );
  XOR U3487 ( .A(n3330), .B(n3313), .Z(n3332) );
  XOR U3488 ( .A(n3333), .B(n3334), .Z(n3313) );
  XOR U3489 ( .A(n3311), .B(n3335), .Z(n3334) );
  XOR U3490 ( .A(n3336), .B(n3337), .Z(n3335) );
  XOR U3491 ( .A(n3338), .B(n3339), .Z(n3337) );
  NAND U3492 ( .A(b[6]), .B(a[39]), .Z(n3339) );
  AND U3493 ( .A(b[7]), .B(a[38]), .Z(n3338) );
  XOR U3494 ( .A(n3340), .B(n3336), .Z(n3333) );
  XOR U3495 ( .A(n3341), .B(n3342), .Z(n3336) );
  NOR U3496 ( .A(n3343), .B(n3344), .Z(n3341) );
  AND U3497 ( .A(b[5]), .B(a[40]), .Z(n3340) );
  XNOR U3498 ( .A(n3345), .B(n3346), .Z(n3330) );
  NOR U3499 ( .A(n3323), .B(n3322), .Z(n3345) );
  XOR U3500 ( .A(n3347), .B(n3346), .Z(n3322) );
  AND U3501 ( .A(b[2]), .B(a[42]), .Z(n3347) );
  XOR U3502 ( .A(n3346), .B(n3349), .Z(n3348) );
  XNOR U3503 ( .A(n3350), .B(n3351), .Z(n3346) );
  NANDN U3504 ( .A(n3326), .B(n3325), .Z(n3351) );
  XOR U3505 ( .A(n3350), .B(n3352), .Z(n3325) );
  NAND U3506 ( .A(b[1]), .B(a[42]), .Z(n3352) );
  XOR U3507 ( .A(n3350), .B(n3354), .Z(n3353) );
  OR U3508 ( .A(n1397), .B(n1395), .Z(n3350) );
  XOR U3509 ( .A(n3356), .B(n3357), .Z(n1395) );
  NANDN U3510 ( .A(n187), .B(a[42]), .Z(n1397) );
  XNOR U3511 ( .A(n3359), .B(n3311), .Z(n3312) );
  XOR U3512 ( .A(n3360), .B(n3361), .Z(n3311) );
  ANDN U3513 ( .B(n3349), .A(n3358), .Z(n3360) );
  XNOR U3514 ( .A(n3362), .B(n3361), .Z(n3358) );
  AND U3515 ( .A(b[3]), .B(a[41]), .Z(n3362) );
  XOR U3516 ( .A(n3361), .B(n3344), .Z(n3363) );
  XOR U3517 ( .A(n3364), .B(n3365), .Z(n3344) );
  XOR U3518 ( .A(n3342), .B(n3366), .Z(n3365) );
  XNOR U3519 ( .A(n3367), .B(n3368), .Z(n3366) );
  XOR U3520 ( .A(n3369), .B(n3370), .Z(n3368) );
  NAND U3521 ( .A(b[6]), .B(a[38]), .Z(n3370) );
  AND U3522 ( .A(b[7]), .B(a[37]), .Z(n3369) );
  XNOR U3523 ( .A(n3371), .B(n3367), .Z(n3364) );
  XOR U3524 ( .A(n3372), .B(n3373), .Z(n3367) );
  NOR U3525 ( .A(n3374), .B(n3375), .Z(n3372) );
  AND U3526 ( .A(b[5]), .B(a[39]), .Z(n3371) );
  XNOR U3527 ( .A(n3376), .B(n3377), .Z(n3361) );
  ANDN U3528 ( .B(n3354), .A(n3355), .Z(n3376) );
  XOR U3529 ( .A(n3378), .B(n3377), .Z(n3355) );
  IV U3530 ( .A(n3379), .Z(n3377) );
  AND U3531 ( .A(b[2]), .B(a[41]), .Z(n3378) );
  XNOR U3532 ( .A(n3381), .B(n3379), .Z(n3380) );
  XOR U3533 ( .A(n3382), .B(n3383), .Z(n3379) );
  NANDN U3534 ( .A(n3357), .B(n3356), .Z(n3383) );
  XOR U3535 ( .A(n3382), .B(n3384), .Z(n3356) );
  NAND U3536 ( .A(b[1]), .B(a[41]), .Z(n3384) );
  XOR U3537 ( .A(n3382), .B(n3386), .Z(n3385) );
  OR U3538 ( .A(n1402), .B(n1400), .Z(n3382) );
  XOR U3539 ( .A(n3388), .B(n3389), .Z(n1400) );
  NANDN U3540 ( .A(n187), .B(a[41]), .Z(n1402) );
  XNOR U3541 ( .A(n3391), .B(n3342), .Z(n3343) );
  XNOR U3542 ( .A(n3392), .B(n3393), .Z(n3342) );
  ANDN U3543 ( .B(n3381), .A(n3390), .Z(n3392) );
  XOR U3544 ( .A(n3394), .B(n3393), .Z(n3390) );
  IV U3545 ( .A(n3395), .Z(n3393) );
  AND U3546 ( .A(b[3]), .B(a[40]), .Z(n3394) );
  XOR U3547 ( .A(n3375), .B(n3395), .Z(n3396) );
  XOR U3548 ( .A(n3397), .B(n3398), .Z(n3395) );
  ANDN U3549 ( .B(n3386), .A(n3387), .Z(n3397) );
  AND U3550 ( .A(b[2]), .B(a[40]), .Z(n3399) );
  XNOR U3551 ( .A(n3401), .B(n3398), .Z(n3400) );
  XOR U3552 ( .A(n3402), .B(n3403), .Z(n3398) );
  NANDN U3553 ( .A(n3389), .B(n3388), .Z(n3403) );
  XOR U3554 ( .A(n3402), .B(n3404), .Z(n3388) );
  NAND U3555 ( .A(b[1]), .B(a[40]), .Z(n3404) );
  XOR U3556 ( .A(n3402), .B(n3406), .Z(n3405) );
  OR U3557 ( .A(n1407), .B(n1405), .Z(n3402) );
  XOR U3558 ( .A(n3408), .B(n3409), .Z(n1405) );
  NANDN U3559 ( .A(n187), .B(a[40]), .Z(n1407) );
  XOR U3560 ( .A(n3411), .B(n3412), .Z(n3375) );
  XNOR U3561 ( .A(n3413), .B(n3414), .Z(n3412) );
  XNOR U3562 ( .A(n3415), .B(n3416), .Z(n3413) );
  XOR U3563 ( .A(n3417), .B(n3418), .Z(n3416) );
  AND U3564 ( .A(b[7]), .B(a[36]), .Z(n3418) );
  AND U3565 ( .A(b[6]), .B(a[37]), .Z(n3417) );
  XNOR U3566 ( .A(n3419), .B(n3415), .Z(n3411) );
  XOR U3567 ( .A(n3420), .B(n3421), .Z(n3415) );
  NOR U3568 ( .A(n3422), .B(n3423), .Z(n3420) );
  AND U3569 ( .A(b[5]), .B(a[38]), .Z(n3419) );
  XOR U3570 ( .A(n3424), .B(n3373), .Z(n3374) );
  IV U3571 ( .A(n3414), .Z(n3373) );
  XOR U3572 ( .A(n3425), .B(n3426), .Z(n3414) );
  ANDN U3573 ( .B(n3401), .A(n3410), .Z(n3425) );
  AND U3574 ( .A(b[3]), .B(a[39]), .Z(n3427) );
  XOR U3575 ( .A(n3423), .B(n3426), .Z(n3428) );
  XOR U3576 ( .A(n3429), .B(n3430), .Z(n3426) );
  ANDN U3577 ( .B(n3406), .A(n3407), .Z(n3429) );
  AND U3578 ( .A(b[2]), .B(a[39]), .Z(n3431) );
  XNOR U3579 ( .A(n3433), .B(n3430), .Z(n3432) );
  XOR U3580 ( .A(n3434), .B(n3435), .Z(n3430) );
  NANDN U3581 ( .A(n3409), .B(n3408), .Z(n3435) );
  XOR U3582 ( .A(n3434), .B(n3436), .Z(n3408) );
  NAND U3583 ( .A(b[1]), .B(a[39]), .Z(n3436) );
  XOR U3584 ( .A(n3434), .B(n3438), .Z(n3437) );
  OR U3585 ( .A(n1412), .B(n1410), .Z(n3434) );
  XOR U3586 ( .A(n3440), .B(n3441), .Z(n1410) );
  NANDN U3587 ( .A(n187), .B(a[39]), .Z(n1412) );
  XOR U3588 ( .A(n3443), .B(n3444), .Z(n3423) );
  XNOR U3589 ( .A(n3445), .B(n3446), .Z(n3444) );
  XNOR U3590 ( .A(n3447), .B(n3448), .Z(n3445) );
  XOR U3591 ( .A(n3449), .B(n3450), .Z(n3448) );
  AND U3592 ( .A(b[6]), .B(a[36]), .Z(n3450) );
  AND U3593 ( .A(b[7]), .B(a[35]), .Z(n3449) );
  XNOR U3594 ( .A(n3451), .B(n3447), .Z(n3443) );
  XOR U3595 ( .A(n3452), .B(n3453), .Z(n3447) );
  NOR U3596 ( .A(n3454), .B(n3455), .Z(n3452) );
  AND U3597 ( .A(b[5]), .B(a[37]), .Z(n3451) );
  XOR U3598 ( .A(n3456), .B(n3421), .Z(n3422) );
  IV U3599 ( .A(n3446), .Z(n3421) );
  XOR U3600 ( .A(n3457), .B(n3458), .Z(n3446) );
  ANDN U3601 ( .B(n3433), .A(n3442), .Z(n3457) );
  AND U3602 ( .A(b[3]), .B(a[38]), .Z(n3459) );
  XOR U3603 ( .A(n3455), .B(n3458), .Z(n3460) );
  XOR U3604 ( .A(n3461), .B(n3462), .Z(n3458) );
  ANDN U3605 ( .B(n3438), .A(n3439), .Z(n3461) );
  AND U3606 ( .A(b[2]), .B(a[38]), .Z(n3463) );
  XOR U3607 ( .A(n3465), .B(n3462), .Z(n3464) );
  XOR U3608 ( .A(n3466), .B(n3467), .Z(n3462) );
  NANDN U3609 ( .A(n3441), .B(n3440), .Z(n3467) );
  XOR U3610 ( .A(n3466), .B(n3468), .Z(n3440) );
  NAND U3611 ( .A(b[1]), .B(a[38]), .Z(n3468) );
  XOR U3612 ( .A(n3466), .B(n3470), .Z(n3469) );
  OR U3613 ( .A(n1417), .B(n1415), .Z(n3466) );
  XOR U3614 ( .A(n3472), .B(n3473), .Z(n1415) );
  NANDN U3615 ( .A(n187), .B(a[38]), .Z(n1417) );
  XOR U3616 ( .A(n3475), .B(n3476), .Z(n3455) );
  XNOR U3617 ( .A(n3477), .B(n3478), .Z(n3476) );
  XOR U3618 ( .A(n3479), .B(n3480), .Z(n3477) );
  AND U3619 ( .A(b[5]), .B(a[36]), .Z(n3479) );
  XOR U3620 ( .A(n3480), .B(n3481), .Z(n3475) );
  XOR U3621 ( .A(n3482), .B(n3483), .Z(n3481) );
  AND U3622 ( .A(b[6]), .B(a[35]), .Z(n3483) );
  AND U3623 ( .A(b[7]), .B(a[34]), .Z(n3482) );
  XOR U3624 ( .A(n3484), .B(n3485), .Z(n3480) );
  ANDN U3625 ( .B(n3486), .A(n3487), .Z(n3484) );
  XOR U3626 ( .A(n3488), .B(n3453), .Z(n3454) );
  IV U3627 ( .A(n3478), .Z(n3453) );
  XOR U3628 ( .A(n3489), .B(n3490), .Z(n3478) );
  NOR U3629 ( .A(n3474), .B(n3465), .Z(n3489) );
  XNOR U3630 ( .A(n3487), .B(n3491), .Z(n3465) );
  XNOR U3631 ( .A(n3486), .B(n3490), .Z(n3491) );
  XOR U3632 ( .A(n3492), .B(n3485), .Z(n3486) );
  AND U3633 ( .A(b[4]), .B(a[36]), .Z(n3492) );
  XOR U3634 ( .A(n3493), .B(n3494), .Z(n3487) );
  XOR U3635 ( .A(n3485), .B(n3495), .Z(n3494) );
  XOR U3636 ( .A(n3496), .B(n3497), .Z(n3495) );
  XOR U3637 ( .A(n3498), .B(n3499), .Z(n3497) );
  NAND U3638 ( .A(b[6]), .B(a[34]), .Z(n3499) );
  AND U3639 ( .A(b[7]), .B(a[33]), .Z(n3498) );
  XOR U3640 ( .A(n3500), .B(n3501), .Z(n3485) );
  ANDN U3641 ( .B(n3502), .A(n3503), .Z(n3500) );
  XOR U3642 ( .A(n3504), .B(n3496), .Z(n3493) );
  XOR U3643 ( .A(n3505), .B(n3506), .Z(n3496) );
  NOR U3644 ( .A(n3507), .B(n3508), .Z(n3505) );
  AND U3645 ( .A(b[5]), .B(a[35]), .Z(n3504) );
  XOR U3646 ( .A(n3510), .B(n3511), .Z(n3490) );
  ANDN U3647 ( .B(n3470), .A(n3471), .Z(n3510) );
  AND U3648 ( .A(b[2]), .B(a[37]), .Z(n3512) );
  XNOR U3649 ( .A(n3502), .B(n3511), .Z(n3513) );
  XOR U3650 ( .A(n3514), .B(n3515), .Z(n3511) );
  NANDN U3651 ( .A(n3473), .B(n3472), .Z(n3515) );
  XOR U3652 ( .A(n3514), .B(n3516), .Z(n3472) );
  NAND U3653 ( .A(b[1]), .B(a[37]), .Z(n3516) );
  XNOR U3654 ( .A(n3514), .B(n3518), .Z(n3517) );
  OR U3655 ( .A(n1422), .B(n1420), .Z(n3514) );
  NANDN U3656 ( .A(n187), .B(a[37]), .Z(n1422) );
  XOR U3657 ( .A(n3522), .B(n3501), .Z(n3502) );
  AND U3658 ( .A(b[3]), .B(a[36]), .Z(n3522) );
  XOR U3659 ( .A(n3501), .B(n3508), .Z(n3523) );
  XOR U3660 ( .A(n3524), .B(n3525), .Z(n3508) );
  XOR U3661 ( .A(n3506), .B(n3526), .Z(n3525) );
  XOR U3662 ( .A(n3527), .B(n3528), .Z(n3526) );
  XOR U3663 ( .A(n3529), .B(n3530), .Z(n3528) );
  NAND U3664 ( .A(b[6]), .B(a[33]), .Z(n3530) );
  AND U3665 ( .A(b[7]), .B(a[32]), .Z(n3529) );
  XOR U3666 ( .A(n3531), .B(n3527), .Z(n3524) );
  XOR U3667 ( .A(n3532), .B(n3533), .Z(n3527) );
  NOR U3668 ( .A(n3534), .B(n3535), .Z(n3532) );
  AND U3669 ( .A(b[5]), .B(a[34]), .Z(n3531) );
  XNOR U3670 ( .A(n3536), .B(n3537), .Z(n3501) );
  NOR U3671 ( .A(n3519), .B(n3518), .Z(n3536) );
  XOR U3672 ( .A(n3538), .B(n3537), .Z(n3518) );
  AND U3673 ( .A(b[2]), .B(a[36]), .Z(n3538) );
  XOR U3674 ( .A(n3537), .B(n3540), .Z(n3539) );
  XNOR U3675 ( .A(n3541), .B(n3542), .Z(n3537) );
  OR U3676 ( .A(n3520), .B(n3521), .Z(n3542) );
  XNOR U3677 ( .A(n3541), .B(n3544), .Z(n3543) );
  XNOR U3678 ( .A(n3541), .B(n3546), .Z(n3520) );
  NAND U3679 ( .A(b[1]), .B(a[36]), .Z(n3546) );
  OR U3680 ( .A(n1427), .B(n1425), .Z(n3541) );
  XOR U3681 ( .A(n3547), .B(n3548), .Z(n1425) );
  NANDN U3682 ( .A(n187), .B(a[36]), .Z(n1427) );
  XNOR U3683 ( .A(n3550), .B(n3506), .Z(n3507) );
  XOR U3684 ( .A(n3551), .B(n3552), .Z(n3506) );
  ANDN U3685 ( .B(n3540), .A(n3549), .Z(n3551) );
  XNOR U3686 ( .A(n3553), .B(n3552), .Z(n3549) );
  AND U3687 ( .A(b[3]), .B(a[35]), .Z(n3553) );
  XOR U3688 ( .A(n3552), .B(n3535), .Z(n3554) );
  XOR U3689 ( .A(n3555), .B(n3556), .Z(n3535) );
  XOR U3690 ( .A(n3533), .B(n3557), .Z(n3556) );
  XOR U3691 ( .A(n3558), .B(n3559), .Z(n3557) );
  XOR U3692 ( .A(n3560), .B(n3561), .Z(n3559) );
  NAND U3693 ( .A(b[6]), .B(a[32]), .Z(n3561) );
  AND U3694 ( .A(b[7]), .B(a[31]), .Z(n3560) );
  XOR U3695 ( .A(n3562), .B(n3558), .Z(n3555) );
  XOR U3696 ( .A(n3563), .B(n3564), .Z(n3558) );
  NOR U3697 ( .A(n3565), .B(n3566), .Z(n3563) );
  AND U3698 ( .A(b[5]), .B(a[33]), .Z(n3562) );
  XNOR U3699 ( .A(n3567), .B(n3568), .Z(n3552) );
  NOR U3700 ( .A(n3545), .B(n3544), .Z(n3567) );
  XOR U3701 ( .A(n3569), .B(n3568), .Z(n3544) );
  AND U3702 ( .A(b[2]), .B(a[35]), .Z(n3569) );
  XOR U3703 ( .A(n3568), .B(n3571), .Z(n3570) );
  XNOR U3704 ( .A(n3572), .B(n3573), .Z(n3568) );
  NANDN U3705 ( .A(n3548), .B(n3547), .Z(n3573) );
  XOR U3706 ( .A(n3572), .B(n3574), .Z(n3547) );
  NAND U3707 ( .A(b[1]), .B(a[35]), .Z(n3574) );
  XOR U3708 ( .A(n3572), .B(n3576), .Z(n3575) );
  OR U3709 ( .A(n1432), .B(n1430), .Z(n3572) );
  XOR U3710 ( .A(n3578), .B(n3579), .Z(n1430) );
  NANDN U3711 ( .A(n187), .B(a[35]), .Z(n1432) );
  XNOR U3712 ( .A(n3581), .B(n3533), .Z(n3534) );
  XOR U3713 ( .A(n3582), .B(n3583), .Z(n3533) );
  ANDN U3714 ( .B(n3571), .A(n3580), .Z(n3582) );
  XNOR U3715 ( .A(n3584), .B(n3583), .Z(n3580) );
  AND U3716 ( .A(b[3]), .B(a[34]), .Z(n3584) );
  XOR U3717 ( .A(n3583), .B(n3566), .Z(n3585) );
  XOR U3718 ( .A(n3586), .B(n3587), .Z(n3566) );
  XOR U3719 ( .A(n3564), .B(n3588), .Z(n3587) );
  XNOR U3720 ( .A(n3589), .B(n3590), .Z(n3588) );
  XOR U3721 ( .A(n3591), .B(n3592), .Z(n3590) );
  NAND U3722 ( .A(b[6]), .B(a[31]), .Z(n3592) );
  AND U3723 ( .A(b[7]), .B(a[30]), .Z(n3591) );
  XNOR U3724 ( .A(n3593), .B(n3589), .Z(n3586) );
  XOR U3725 ( .A(n3594), .B(n3595), .Z(n3589) );
  NOR U3726 ( .A(n3596), .B(n3597), .Z(n3594) );
  AND U3727 ( .A(b[5]), .B(a[32]), .Z(n3593) );
  XNOR U3728 ( .A(n3598), .B(n3599), .Z(n3583) );
  ANDN U3729 ( .B(n3576), .A(n3577), .Z(n3598) );
  XOR U3730 ( .A(n3600), .B(n3599), .Z(n3577) );
  IV U3731 ( .A(n3601), .Z(n3599) );
  AND U3732 ( .A(b[2]), .B(a[34]), .Z(n3600) );
  XNOR U3733 ( .A(n3603), .B(n3601), .Z(n3602) );
  XOR U3734 ( .A(n3604), .B(n3605), .Z(n3601) );
  NANDN U3735 ( .A(n3579), .B(n3578), .Z(n3605) );
  XOR U3736 ( .A(n3604), .B(n3606), .Z(n3578) );
  NAND U3737 ( .A(b[1]), .B(a[34]), .Z(n3606) );
  XOR U3738 ( .A(n3604), .B(n3608), .Z(n3607) );
  OR U3739 ( .A(n1437), .B(n1435), .Z(n3604) );
  XOR U3740 ( .A(n3610), .B(n3611), .Z(n1435) );
  NANDN U3741 ( .A(n187), .B(a[34]), .Z(n1437) );
  XNOR U3742 ( .A(n3613), .B(n3564), .Z(n3565) );
  XNOR U3743 ( .A(n3614), .B(n3615), .Z(n3564) );
  ANDN U3744 ( .B(n3603), .A(n3612), .Z(n3614) );
  XOR U3745 ( .A(n3616), .B(n3615), .Z(n3612) );
  IV U3746 ( .A(n3617), .Z(n3615) );
  AND U3747 ( .A(b[3]), .B(a[33]), .Z(n3616) );
  XOR U3748 ( .A(n3597), .B(n3617), .Z(n3618) );
  XOR U3749 ( .A(n3619), .B(n3620), .Z(n3617) );
  ANDN U3750 ( .B(n3608), .A(n3609), .Z(n3619) );
  AND U3751 ( .A(b[2]), .B(a[33]), .Z(n3621) );
  XNOR U3752 ( .A(n3623), .B(n3620), .Z(n3622) );
  XOR U3753 ( .A(n3624), .B(n3625), .Z(n3620) );
  NANDN U3754 ( .A(n3611), .B(n3610), .Z(n3625) );
  XOR U3755 ( .A(n3624), .B(n3626), .Z(n3610) );
  NAND U3756 ( .A(b[1]), .B(a[33]), .Z(n3626) );
  XOR U3757 ( .A(n3624), .B(n3628), .Z(n3627) );
  OR U3758 ( .A(n1442), .B(n1440), .Z(n3624) );
  XOR U3759 ( .A(n3630), .B(n3631), .Z(n1440) );
  NANDN U3760 ( .A(n187), .B(a[33]), .Z(n1442) );
  XOR U3761 ( .A(n3633), .B(n3634), .Z(n3597) );
  XNOR U3762 ( .A(n3635), .B(n3636), .Z(n3634) );
  XNOR U3763 ( .A(n3637), .B(n3638), .Z(n3635) );
  XOR U3764 ( .A(n3639), .B(n3640), .Z(n3638) );
  AND U3765 ( .A(b[7]), .B(a[29]), .Z(n3640) );
  AND U3766 ( .A(b[6]), .B(a[30]), .Z(n3639) );
  XNOR U3767 ( .A(n3641), .B(n3637), .Z(n3633) );
  XOR U3768 ( .A(n3642), .B(n3643), .Z(n3637) );
  NOR U3769 ( .A(n3644), .B(n3645), .Z(n3642) );
  AND U3770 ( .A(b[5]), .B(a[31]), .Z(n3641) );
  XOR U3771 ( .A(n3646), .B(n3595), .Z(n3596) );
  IV U3772 ( .A(n3636), .Z(n3595) );
  XOR U3773 ( .A(n3647), .B(n3648), .Z(n3636) );
  ANDN U3774 ( .B(n3623), .A(n3632), .Z(n3647) );
  AND U3775 ( .A(b[3]), .B(a[32]), .Z(n3649) );
  XOR U3776 ( .A(n3645), .B(n3648), .Z(n3650) );
  XOR U3777 ( .A(n3651), .B(n3652), .Z(n3648) );
  ANDN U3778 ( .B(n3628), .A(n3629), .Z(n3651) );
  AND U3779 ( .A(b[2]), .B(a[32]), .Z(n3653) );
  XNOR U3780 ( .A(n3655), .B(n3652), .Z(n3654) );
  XOR U3781 ( .A(n3656), .B(n3657), .Z(n3652) );
  NANDN U3782 ( .A(n3631), .B(n3630), .Z(n3657) );
  XOR U3783 ( .A(n3656), .B(n3658), .Z(n3630) );
  NAND U3784 ( .A(b[1]), .B(a[32]), .Z(n3658) );
  XOR U3785 ( .A(n3656), .B(n3660), .Z(n3659) );
  OR U3786 ( .A(n1447), .B(n1445), .Z(n3656) );
  XOR U3787 ( .A(n3662), .B(n3663), .Z(n1445) );
  NANDN U3788 ( .A(n187), .B(a[32]), .Z(n1447) );
  XOR U3789 ( .A(n3665), .B(n3666), .Z(n3645) );
  XNOR U3790 ( .A(n3667), .B(n3668), .Z(n3666) );
  XNOR U3791 ( .A(n3669), .B(n3670), .Z(n3667) );
  XOR U3792 ( .A(n3671), .B(n3672), .Z(n3670) );
  AND U3793 ( .A(b[6]), .B(a[29]), .Z(n3672) );
  AND U3794 ( .A(b[7]), .B(a[28]), .Z(n3671) );
  XNOR U3795 ( .A(n3673), .B(n3669), .Z(n3665) );
  XOR U3796 ( .A(n3674), .B(n3675), .Z(n3669) );
  NOR U3797 ( .A(n3676), .B(n3677), .Z(n3674) );
  AND U3798 ( .A(b[5]), .B(a[30]), .Z(n3673) );
  XOR U3799 ( .A(n3678), .B(n3643), .Z(n3644) );
  IV U3800 ( .A(n3668), .Z(n3643) );
  XOR U3801 ( .A(n3679), .B(n3680), .Z(n3668) );
  ANDN U3802 ( .B(n3655), .A(n3664), .Z(n3679) );
  AND U3803 ( .A(b[3]), .B(a[31]), .Z(n3681) );
  XOR U3804 ( .A(n3677), .B(n3680), .Z(n3682) );
  XOR U3805 ( .A(n3683), .B(n3684), .Z(n3680) );
  ANDN U3806 ( .B(n3660), .A(n3661), .Z(n3683) );
  AND U3807 ( .A(b[2]), .B(a[31]), .Z(n3685) );
  XOR U3808 ( .A(n3687), .B(n3684), .Z(n3686) );
  XOR U3809 ( .A(n3688), .B(n3689), .Z(n3684) );
  NANDN U3810 ( .A(n3663), .B(n3662), .Z(n3689) );
  XOR U3811 ( .A(n3688), .B(n3690), .Z(n3662) );
  NAND U3812 ( .A(b[1]), .B(a[31]), .Z(n3690) );
  XOR U3813 ( .A(n3688), .B(n3692), .Z(n3691) );
  OR U3814 ( .A(n1452), .B(n1450), .Z(n3688) );
  XOR U3815 ( .A(n3694), .B(n3695), .Z(n1450) );
  NANDN U3816 ( .A(n187), .B(a[31]), .Z(n1452) );
  XOR U3817 ( .A(n3697), .B(n3698), .Z(n3677) );
  XNOR U3818 ( .A(n3699), .B(n3700), .Z(n3698) );
  XOR U3819 ( .A(n3701), .B(n3702), .Z(n3699) );
  AND U3820 ( .A(b[5]), .B(a[29]), .Z(n3701) );
  XOR U3821 ( .A(n3702), .B(n3703), .Z(n3697) );
  XOR U3822 ( .A(n3704), .B(n3705), .Z(n3703) );
  AND U3823 ( .A(b[6]), .B(a[28]), .Z(n3705) );
  AND U3824 ( .A(b[7]), .B(a[27]), .Z(n3704) );
  XOR U3825 ( .A(n3706), .B(n3707), .Z(n3702) );
  ANDN U3826 ( .B(n3708), .A(n3709), .Z(n3706) );
  XOR U3827 ( .A(n3710), .B(n3675), .Z(n3676) );
  IV U3828 ( .A(n3700), .Z(n3675) );
  XOR U3829 ( .A(n3711), .B(n3712), .Z(n3700) );
  NOR U3830 ( .A(n3696), .B(n3687), .Z(n3711) );
  XNOR U3831 ( .A(n3709), .B(n3713), .Z(n3687) );
  XNOR U3832 ( .A(n3708), .B(n3712), .Z(n3713) );
  XOR U3833 ( .A(n3714), .B(n3707), .Z(n3708) );
  AND U3834 ( .A(b[4]), .B(a[29]), .Z(n3714) );
  XOR U3835 ( .A(n3715), .B(n3716), .Z(n3709) );
  XOR U3836 ( .A(n3707), .B(n3717), .Z(n3716) );
  XOR U3837 ( .A(n3718), .B(n3719), .Z(n3717) );
  XOR U3838 ( .A(n3720), .B(n3721), .Z(n3719) );
  NAND U3839 ( .A(b[6]), .B(a[27]), .Z(n3721) );
  AND U3840 ( .A(b[7]), .B(a[26]), .Z(n3720) );
  XOR U3841 ( .A(n3722), .B(n3723), .Z(n3707) );
  ANDN U3842 ( .B(n3724), .A(n3725), .Z(n3722) );
  XOR U3843 ( .A(n3726), .B(n3718), .Z(n3715) );
  XOR U3844 ( .A(n3727), .B(n3728), .Z(n3718) );
  NOR U3845 ( .A(n3729), .B(n3730), .Z(n3727) );
  AND U3846 ( .A(b[5]), .B(a[28]), .Z(n3726) );
  XOR U3847 ( .A(n3732), .B(n3733), .Z(n3712) );
  ANDN U3848 ( .B(n3692), .A(n3693), .Z(n3732) );
  AND U3849 ( .A(b[2]), .B(a[30]), .Z(n3734) );
  XNOR U3850 ( .A(n3724), .B(n3733), .Z(n3735) );
  XOR U3851 ( .A(n3736), .B(n3737), .Z(n3733) );
  NANDN U3852 ( .A(n3695), .B(n3694), .Z(n3737) );
  XOR U3853 ( .A(n3736), .B(n3738), .Z(n3694) );
  NAND U3854 ( .A(b[1]), .B(a[30]), .Z(n3738) );
  XNOR U3855 ( .A(n3736), .B(n3740), .Z(n3739) );
  OR U3856 ( .A(n1457), .B(n1455), .Z(n3736) );
  NANDN U3857 ( .A(n187), .B(a[30]), .Z(n1457) );
  XOR U3858 ( .A(n3744), .B(n3723), .Z(n3724) );
  AND U3859 ( .A(b[3]), .B(a[29]), .Z(n3744) );
  XOR U3860 ( .A(n3723), .B(n3730), .Z(n3745) );
  XOR U3861 ( .A(n3746), .B(n3747), .Z(n3730) );
  XOR U3862 ( .A(n3728), .B(n3748), .Z(n3747) );
  XOR U3863 ( .A(n3749), .B(n3750), .Z(n3748) );
  XOR U3864 ( .A(n3751), .B(n3752), .Z(n3750) );
  NAND U3865 ( .A(b[6]), .B(a[26]), .Z(n3752) );
  AND U3866 ( .A(b[7]), .B(a[25]), .Z(n3751) );
  XOR U3867 ( .A(n3753), .B(n3749), .Z(n3746) );
  XOR U3868 ( .A(n3754), .B(n3755), .Z(n3749) );
  NOR U3869 ( .A(n3756), .B(n3757), .Z(n3754) );
  AND U3870 ( .A(b[5]), .B(a[27]), .Z(n3753) );
  XNOR U3871 ( .A(n3758), .B(n3759), .Z(n3723) );
  NOR U3872 ( .A(n3741), .B(n3740), .Z(n3758) );
  XOR U3873 ( .A(n3760), .B(n3759), .Z(n3740) );
  AND U3874 ( .A(b[2]), .B(a[29]), .Z(n3760) );
  XOR U3875 ( .A(n3759), .B(n3762), .Z(n3761) );
  XNOR U3876 ( .A(n3763), .B(n3764), .Z(n3759) );
  OR U3877 ( .A(n3742), .B(n3743), .Z(n3764) );
  XNOR U3878 ( .A(n3763), .B(n3766), .Z(n3765) );
  XNOR U3879 ( .A(n3763), .B(n3768), .Z(n3742) );
  NAND U3880 ( .A(b[1]), .B(a[29]), .Z(n3768) );
  OR U3881 ( .A(n1462), .B(n1460), .Z(n3763) );
  XOR U3882 ( .A(n3769), .B(n3770), .Z(n1460) );
  NANDN U3883 ( .A(n187), .B(a[29]), .Z(n1462) );
  XNOR U3884 ( .A(n3772), .B(n3728), .Z(n3729) );
  XOR U3885 ( .A(n3773), .B(n3774), .Z(n3728) );
  ANDN U3886 ( .B(n3762), .A(n3771), .Z(n3773) );
  XNOR U3887 ( .A(n3775), .B(n3774), .Z(n3771) );
  AND U3888 ( .A(b[3]), .B(a[28]), .Z(n3775) );
  XOR U3889 ( .A(n3774), .B(n3757), .Z(n3776) );
  XOR U3890 ( .A(n3777), .B(n3778), .Z(n3757) );
  XOR U3891 ( .A(n3755), .B(n3779), .Z(n3778) );
  XOR U3892 ( .A(n3780), .B(n3781), .Z(n3779) );
  XOR U3893 ( .A(n3782), .B(n3783), .Z(n3781) );
  NAND U3894 ( .A(b[6]), .B(a[25]), .Z(n3783) );
  AND U3895 ( .A(b[7]), .B(a[24]), .Z(n3782) );
  XOR U3896 ( .A(n3784), .B(n3780), .Z(n3777) );
  XOR U3897 ( .A(n3785), .B(n3786), .Z(n3780) );
  NOR U3898 ( .A(n3787), .B(n3788), .Z(n3785) );
  AND U3899 ( .A(b[5]), .B(a[26]), .Z(n3784) );
  XNOR U3900 ( .A(n3789), .B(n3790), .Z(n3774) );
  NOR U3901 ( .A(n3767), .B(n3766), .Z(n3789) );
  XOR U3902 ( .A(n3791), .B(n3790), .Z(n3766) );
  AND U3903 ( .A(b[2]), .B(a[28]), .Z(n3791) );
  XOR U3904 ( .A(n3790), .B(n3793), .Z(n3792) );
  XNOR U3905 ( .A(n3794), .B(n3795), .Z(n3790) );
  NANDN U3906 ( .A(n3770), .B(n3769), .Z(n3795) );
  XOR U3907 ( .A(n3794), .B(n3796), .Z(n3769) );
  NAND U3908 ( .A(b[1]), .B(a[28]), .Z(n3796) );
  XOR U3909 ( .A(n3794), .B(n3798), .Z(n3797) );
  OR U3910 ( .A(n1467), .B(n1465), .Z(n3794) );
  XOR U3911 ( .A(n3800), .B(n3801), .Z(n1465) );
  NANDN U3912 ( .A(n187), .B(a[28]), .Z(n1467) );
  XNOR U3913 ( .A(n3803), .B(n3755), .Z(n3756) );
  XOR U3914 ( .A(n3804), .B(n3805), .Z(n3755) );
  ANDN U3915 ( .B(n3793), .A(n3802), .Z(n3804) );
  XNOR U3916 ( .A(n3806), .B(n3805), .Z(n3802) );
  AND U3917 ( .A(b[3]), .B(a[27]), .Z(n3806) );
  XOR U3918 ( .A(n3805), .B(n3788), .Z(n3807) );
  XOR U3919 ( .A(n3808), .B(n3809), .Z(n3788) );
  XOR U3920 ( .A(n3786), .B(n3810), .Z(n3809) );
  XNOR U3921 ( .A(n3811), .B(n3812), .Z(n3810) );
  XOR U3922 ( .A(n3813), .B(n3814), .Z(n3812) );
  NAND U3923 ( .A(b[6]), .B(a[24]), .Z(n3814) );
  AND U3924 ( .A(b[7]), .B(a[23]), .Z(n3813) );
  XNOR U3925 ( .A(n3815), .B(n3811), .Z(n3808) );
  XOR U3926 ( .A(n3816), .B(n3817), .Z(n3811) );
  NOR U3927 ( .A(n3818), .B(n3819), .Z(n3816) );
  AND U3928 ( .A(b[5]), .B(a[25]), .Z(n3815) );
  XNOR U3929 ( .A(n3820), .B(n3821), .Z(n3805) );
  ANDN U3930 ( .B(n3798), .A(n3799), .Z(n3820) );
  XOR U3931 ( .A(n3822), .B(n3821), .Z(n3799) );
  IV U3932 ( .A(n3823), .Z(n3821) );
  AND U3933 ( .A(b[2]), .B(a[27]), .Z(n3822) );
  XNOR U3934 ( .A(n3825), .B(n3823), .Z(n3824) );
  XOR U3935 ( .A(n3826), .B(n3827), .Z(n3823) );
  NANDN U3936 ( .A(n3801), .B(n3800), .Z(n3827) );
  XOR U3937 ( .A(n3826), .B(n3828), .Z(n3800) );
  NAND U3938 ( .A(b[1]), .B(a[27]), .Z(n3828) );
  XOR U3939 ( .A(n3826), .B(n3830), .Z(n3829) );
  OR U3940 ( .A(n1472), .B(n1470), .Z(n3826) );
  XOR U3941 ( .A(n3832), .B(n3833), .Z(n1470) );
  NANDN U3942 ( .A(n187), .B(a[27]), .Z(n1472) );
  XNOR U3943 ( .A(n3835), .B(n3786), .Z(n3787) );
  XNOR U3944 ( .A(n3836), .B(n3837), .Z(n3786) );
  ANDN U3945 ( .B(n3825), .A(n3834), .Z(n3836) );
  XOR U3946 ( .A(n3838), .B(n3837), .Z(n3834) );
  IV U3947 ( .A(n3839), .Z(n3837) );
  AND U3948 ( .A(b[3]), .B(a[26]), .Z(n3838) );
  XOR U3949 ( .A(n3819), .B(n3839), .Z(n3840) );
  XOR U3950 ( .A(n3841), .B(n3842), .Z(n3839) );
  ANDN U3951 ( .B(n3830), .A(n3831), .Z(n3841) );
  AND U3952 ( .A(b[2]), .B(a[26]), .Z(n3843) );
  XNOR U3953 ( .A(n3845), .B(n3842), .Z(n3844) );
  XOR U3954 ( .A(n3846), .B(n3847), .Z(n3842) );
  NANDN U3955 ( .A(n3833), .B(n3832), .Z(n3847) );
  XOR U3956 ( .A(n3846), .B(n3848), .Z(n3832) );
  NAND U3957 ( .A(b[1]), .B(a[26]), .Z(n3848) );
  XOR U3958 ( .A(n3846), .B(n3850), .Z(n3849) );
  OR U3959 ( .A(n1477), .B(n1475), .Z(n3846) );
  XOR U3960 ( .A(n3852), .B(n3853), .Z(n1475) );
  NANDN U3961 ( .A(n187), .B(a[26]), .Z(n1477) );
  XOR U3962 ( .A(n3855), .B(n3856), .Z(n3819) );
  XNOR U3963 ( .A(n3857), .B(n3858), .Z(n3856) );
  XNOR U3964 ( .A(n3859), .B(n3860), .Z(n3857) );
  XOR U3965 ( .A(n3861), .B(n3862), .Z(n3860) );
  AND U3966 ( .A(b[7]), .B(a[22]), .Z(n3862) );
  AND U3967 ( .A(b[6]), .B(a[23]), .Z(n3861) );
  XNOR U3968 ( .A(n3863), .B(n3859), .Z(n3855) );
  XOR U3969 ( .A(n3864), .B(n3865), .Z(n3859) );
  NOR U3970 ( .A(n3866), .B(n3867), .Z(n3864) );
  AND U3971 ( .A(b[5]), .B(a[24]), .Z(n3863) );
  XOR U3972 ( .A(n3868), .B(n3817), .Z(n3818) );
  IV U3973 ( .A(n3858), .Z(n3817) );
  XOR U3974 ( .A(n3869), .B(n3870), .Z(n3858) );
  ANDN U3975 ( .B(n3845), .A(n3854), .Z(n3869) );
  AND U3976 ( .A(b[3]), .B(a[25]), .Z(n3871) );
  XOR U3977 ( .A(n3867), .B(n3870), .Z(n3872) );
  XOR U3978 ( .A(n3873), .B(n3874), .Z(n3870) );
  ANDN U3979 ( .B(n3850), .A(n3851), .Z(n3873) );
  AND U3980 ( .A(b[2]), .B(a[25]), .Z(n3875) );
  XNOR U3981 ( .A(n3877), .B(n3874), .Z(n3876) );
  XOR U3982 ( .A(n3878), .B(n3879), .Z(n3874) );
  NANDN U3983 ( .A(n3853), .B(n3852), .Z(n3879) );
  XOR U3984 ( .A(n3878), .B(n3880), .Z(n3852) );
  NAND U3985 ( .A(b[1]), .B(a[25]), .Z(n3880) );
  XOR U3986 ( .A(n3878), .B(n3882), .Z(n3881) );
  OR U3987 ( .A(n1482), .B(n1480), .Z(n3878) );
  XOR U3988 ( .A(n3884), .B(n3885), .Z(n1480) );
  NANDN U3989 ( .A(n187), .B(a[25]), .Z(n1482) );
  XOR U3990 ( .A(n3887), .B(n3888), .Z(n3867) );
  XNOR U3991 ( .A(n3889), .B(n3890), .Z(n3888) );
  XNOR U3992 ( .A(n3891), .B(n3892), .Z(n3889) );
  XOR U3993 ( .A(n3893), .B(n3894), .Z(n3892) );
  AND U3994 ( .A(b[6]), .B(a[22]), .Z(n3894) );
  AND U3995 ( .A(b[7]), .B(a[21]), .Z(n3893) );
  XNOR U3996 ( .A(n3895), .B(n3891), .Z(n3887) );
  XOR U3997 ( .A(n3896), .B(n3897), .Z(n3891) );
  NOR U3998 ( .A(n3898), .B(n3899), .Z(n3896) );
  AND U3999 ( .A(b[5]), .B(a[23]), .Z(n3895) );
  XOR U4000 ( .A(n3900), .B(n3865), .Z(n3866) );
  IV U4001 ( .A(n3890), .Z(n3865) );
  XOR U4002 ( .A(n3901), .B(n3902), .Z(n3890) );
  ANDN U4003 ( .B(n3877), .A(n3886), .Z(n3901) );
  AND U4004 ( .A(b[3]), .B(a[24]), .Z(n3903) );
  XOR U4005 ( .A(n3899), .B(n3902), .Z(n3904) );
  XOR U4006 ( .A(n3905), .B(n3906), .Z(n3902) );
  ANDN U4007 ( .B(n3882), .A(n3883), .Z(n3905) );
  AND U4008 ( .A(b[2]), .B(a[24]), .Z(n3907) );
  XOR U4009 ( .A(n3909), .B(n3906), .Z(n3908) );
  XOR U4010 ( .A(n3910), .B(n3911), .Z(n3906) );
  NANDN U4011 ( .A(n3885), .B(n3884), .Z(n3911) );
  XOR U4012 ( .A(n3910), .B(n3912), .Z(n3884) );
  NAND U4013 ( .A(b[1]), .B(a[24]), .Z(n3912) );
  XOR U4014 ( .A(n3910), .B(n3914), .Z(n3913) );
  OR U4015 ( .A(n1487), .B(n1485), .Z(n3910) );
  XOR U4016 ( .A(n3916), .B(n3917), .Z(n1485) );
  NANDN U4017 ( .A(n187), .B(a[24]), .Z(n1487) );
  XOR U4018 ( .A(n3919), .B(n3920), .Z(n3899) );
  XNOR U4019 ( .A(n3921), .B(n3922), .Z(n3920) );
  XOR U4020 ( .A(n3923), .B(n3924), .Z(n3921) );
  AND U4021 ( .A(b[5]), .B(a[22]), .Z(n3923) );
  XOR U4022 ( .A(n3924), .B(n3925), .Z(n3919) );
  XOR U4023 ( .A(n3926), .B(n3927), .Z(n3925) );
  AND U4024 ( .A(b[6]), .B(a[21]), .Z(n3927) );
  AND U4025 ( .A(b[7]), .B(a[20]), .Z(n3926) );
  XOR U4026 ( .A(n3928), .B(n3929), .Z(n3924) );
  ANDN U4027 ( .B(n3930), .A(n3931), .Z(n3928) );
  XOR U4028 ( .A(n3932), .B(n3897), .Z(n3898) );
  IV U4029 ( .A(n3922), .Z(n3897) );
  XOR U4030 ( .A(n3933), .B(n3934), .Z(n3922) );
  NOR U4031 ( .A(n3918), .B(n3909), .Z(n3933) );
  XNOR U4032 ( .A(n3931), .B(n3935), .Z(n3909) );
  XNOR U4033 ( .A(n3930), .B(n3934), .Z(n3935) );
  XOR U4034 ( .A(n3936), .B(n3929), .Z(n3930) );
  AND U4035 ( .A(b[4]), .B(a[22]), .Z(n3936) );
  XOR U4036 ( .A(n3937), .B(n3938), .Z(n3931) );
  XOR U4037 ( .A(n3929), .B(n3939), .Z(n3938) );
  XOR U4038 ( .A(n3940), .B(n3941), .Z(n3939) );
  XOR U4039 ( .A(n3942), .B(n3943), .Z(n3941) );
  NAND U4040 ( .A(b[6]), .B(a[20]), .Z(n3943) );
  AND U4041 ( .A(b[7]), .B(a[19]), .Z(n3942) );
  XOR U4042 ( .A(n3944), .B(n3945), .Z(n3929) );
  ANDN U4043 ( .B(n3946), .A(n3947), .Z(n3944) );
  XOR U4044 ( .A(n3948), .B(n3940), .Z(n3937) );
  XOR U4045 ( .A(n3949), .B(n3950), .Z(n3940) );
  NOR U4046 ( .A(n3951), .B(n3952), .Z(n3949) );
  AND U4047 ( .A(b[5]), .B(a[21]), .Z(n3948) );
  XOR U4048 ( .A(n3954), .B(n3955), .Z(n3934) );
  ANDN U4049 ( .B(n3914), .A(n3915), .Z(n3954) );
  AND U4050 ( .A(b[2]), .B(a[23]), .Z(n3956) );
  XNOR U4051 ( .A(n3946), .B(n3955), .Z(n3957) );
  XOR U4052 ( .A(n3958), .B(n3959), .Z(n3955) );
  NANDN U4053 ( .A(n3917), .B(n3916), .Z(n3959) );
  XOR U4054 ( .A(n3958), .B(n3960), .Z(n3916) );
  NAND U4055 ( .A(b[1]), .B(a[23]), .Z(n3960) );
  XNOR U4056 ( .A(n3958), .B(n3962), .Z(n3961) );
  OR U4057 ( .A(n1492), .B(n1490), .Z(n3958) );
  NANDN U4058 ( .A(n187), .B(a[23]), .Z(n1492) );
  XOR U4059 ( .A(n3966), .B(n3945), .Z(n3946) );
  AND U4060 ( .A(b[3]), .B(a[22]), .Z(n3966) );
  XOR U4061 ( .A(n3945), .B(n3952), .Z(n3967) );
  XOR U4062 ( .A(n3968), .B(n3969), .Z(n3952) );
  XOR U4063 ( .A(n3950), .B(n3970), .Z(n3969) );
  XOR U4064 ( .A(n3971), .B(n3972), .Z(n3970) );
  XOR U4065 ( .A(n3973), .B(n3974), .Z(n3972) );
  NAND U4066 ( .A(b[6]), .B(a[19]), .Z(n3974) );
  AND U4067 ( .A(b[7]), .B(a[18]), .Z(n3973) );
  XOR U4068 ( .A(n3975), .B(n3971), .Z(n3968) );
  XOR U4069 ( .A(n3976), .B(n3977), .Z(n3971) );
  NOR U4070 ( .A(n3978), .B(n3979), .Z(n3976) );
  AND U4071 ( .A(b[5]), .B(a[20]), .Z(n3975) );
  XNOR U4072 ( .A(n3980), .B(n3981), .Z(n3945) );
  NOR U4073 ( .A(n3963), .B(n3962), .Z(n3980) );
  XOR U4074 ( .A(n3982), .B(n3981), .Z(n3962) );
  AND U4075 ( .A(b[2]), .B(a[22]), .Z(n3982) );
  XOR U4076 ( .A(n3981), .B(n3984), .Z(n3983) );
  XNOR U4077 ( .A(n3985), .B(n3986), .Z(n3981) );
  OR U4078 ( .A(n3964), .B(n3965), .Z(n3986) );
  XNOR U4079 ( .A(n3985), .B(n3988), .Z(n3987) );
  XNOR U4080 ( .A(n3985), .B(n3990), .Z(n3964) );
  NAND U4081 ( .A(b[1]), .B(a[22]), .Z(n3990) );
  OR U4082 ( .A(n1497), .B(n1495), .Z(n3985) );
  XOR U4083 ( .A(n3991), .B(n3992), .Z(n1495) );
  NANDN U4084 ( .A(n187), .B(a[22]), .Z(n1497) );
  XNOR U4085 ( .A(n3994), .B(n3950), .Z(n3951) );
  XOR U4086 ( .A(n3995), .B(n3996), .Z(n3950) );
  ANDN U4087 ( .B(n3984), .A(n3993), .Z(n3995) );
  XNOR U4088 ( .A(n3997), .B(n3996), .Z(n3993) );
  AND U4089 ( .A(b[3]), .B(a[21]), .Z(n3997) );
  XOR U4090 ( .A(n3996), .B(n3979), .Z(n3998) );
  XOR U4091 ( .A(n3999), .B(n4000), .Z(n3979) );
  XOR U4092 ( .A(n3977), .B(n4001), .Z(n4000) );
  XOR U4093 ( .A(n4002), .B(n4003), .Z(n4001) );
  XOR U4094 ( .A(n4004), .B(n4005), .Z(n4003) );
  NAND U4095 ( .A(b[6]), .B(a[18]), .Z(n4005) );
  AND U4096 ( .A(b[7]), .B(a[17]), .Z(n4004) );
  XOR U4097 ( .A(n4006), .B(n4002), .Z(n3999) );
  XOR U4098 ( .A(n4007), .B(n4008), .Z(n4002) );
  NOR U4099 ( .A(n4009), .B(n4010), .Z(n4007) );
  AND U4100 ( .A(b[5]), .B(a[19]), .Z(n4006) );
  XNOR U4101 ( .A(n4011), .B(n4012), .Z(n3996) );
  NOR U4102 ( .A(n3989), .B(n3988), .Z(n4011) );
  XOR U4103 ( .A(n4013), .B(n4012), .Z(n3988) );
  AND U4104 ( .A(b[2]), .B(a[21]), .Z(n4013) );
  XOR U4105 ( .A(n4012), .B(n4015), .Z(n4014) );
  XNOR U4106 ( .A(n4016), .B(n4017), .Z(n4012) );
  NANDN U4107 ( .A(n3992), .B(n3991), .Z(n4017) );
  XOR U4108 ( .A(n4016), .B(n4018), .Z(n3991) );
  NAND U4109 ( .A(b[1]), .B(a[21]), .Z(n4018) );
  XOR U4110 ( .A(n4016), .B(n4020), .Z(n4019) );
  OR U4111 ( .A(n1502), .B(n1500), .Z(n4016) );
  XOR U4112 ( .A(n4022), .B(n4023), .Z(n1500) );
  NANDN U4113 ( .A(n187), .B(a[21]), .Z(n1502) );
  XNOR U4114 ( .A(n4025), .B(n3977), .Z(n3978) );
  XOR U4115 ( .A(n4026), .B(n4027), .Z(n3977) );
  ANDN U4116 ( .B(n4015), .A(n4024), .Z(n4026) );
  XNOR U4117 ( .A(n4028), .B(n4027), .Z(n4024) );
  AND U4118 ( .A(b[3]), .B(a[20]), .Z(n4028) );
  XOR U4119 ( .A(n4027), .B(n4010), .Z(n4029) );
  XOR U4120 ( .A(n4030), .B(n4031), .Z(n4010) );
  XOR U4121 ( .A(n4008), .B(n4032), .Z(n4031) );
  XNOR U4122 ( .A(n4033), .B(n4034), .Z(n4032) );
  XOR U4123 ( .A(n4035), .B(n4036), .Z(n4034) );
  NAND U4124 ( .A(b[6]), .B(a[17]), .Z(n4036) );
  AND U4125 ( .A(b[7]), .B(a[16]), .Z(n4035) );
  XNOR U4126 ( .A(n4037), .B(n4033), .Z(n4030) );
  XOR U4127 ( .A(n4038), .B(n4039), .Z(n4033) );
  NOR U4128 ( .A(n4040), .B(n4041), .Z(n4038) );
  AND U4129 ( .A(b[5]), .B(a[18]), .Z(n4037) );
  XNOR U4130 ( .A(n4042), .B(n4043), .Z(n4027) );
  ANDN U4131 ( .B(n4020), .A(n4021), .Z(n4042) );
  XOR U4132 ( .A(n4044), .B(n4043), .Z(n4021) );
  IV U4133 ( .A(n4045), .Z(n4043) );
  AND U4134 ( .A(b[2]), .B(a[20]), .Z(n4044) );
  XNOR U4135 ( .A(n4047), .B(n4045), .Z(n4046) );
  XOR U4136 ( .A(n4048), .B(n4049), .Z(n4045) );
  NANDN U4137 ( .A(n4023), .B(n4022), .Z(n4049) );
  XOR U4138 ( .A(n4048), .B(n4050), .Z(n4022) );
  NAND U4139 ( .A(b[1]), .B(a[20]), .Z(n4050) );
  XOR U4140 ( .A(n4048), .B(n4052), .Z(n4051) );
  OR U4141 ( .A(n1507), .B(n1505), .Z(n4048) );
  XOR U4142 ( .A(n4054), .B(n4055), .Z(n1505) );
  NANDN U4143 ( .A(n187), .B(a[20]), .Z(n1507) );
  XNOR U4144 ( .A(n4057), .B(n4008), .Z(n4009) );
  XNOR U4145 ( .A(n4058), .B(n4059), .Z(n4008) );
  ANDN U4146 ( .B(n4047), .A(n4056), .Z(n4058) );
  XOR U4147 ( .A(n4060), .B(n4059), .Z(n4056) );
  IV U4148 ( .A(n4061), .Z(n4059) );
  AND U4149 ( .A(b[3]), .B(a[19]), .Z(n4060) );
  XOR U4150 ( .A(n4041), .B(n4061), .Z(n4062) );
  XOR U4151 ( .A(n4063), .B(n4064), .Z(n4061) );
  ANDN U4152 ( .B(n4052), .A(n4053), .Z(n4063) );
  AND U4153 ( .A(b[2]), .B(a[19]), .Z(n4065) );
  XNOR U4154 ( .A(n4067), .B(n4064), .Z(n4066) );
  XOR U4155 ( .A(n4068), .B(n4069), .Z(n4064) );
  NANDN U4156 ( .A(n4055), .B(n4054), .Z(n4069) );
  XOR U4157 ( .A(n4068), .B(n4070), .Z(n4054) );
  NAND U4158 ( .A(b[1]), .B(a[19]), .Z(n4070) );
  XOR U4159 ( .A(n4068), .B(n4072), .Z(n4071) );
  OR U4160 ( .A(n1512), .B(n1510), .Z(n4068) );
  XOR U4161 ( .A(n4074), .B(n4075), .Z(n1510) );
  NANDN U4162 ( .A(n187), .B(a[19]), .Z(n1512) );
  XOR U4163 ( .A(n4077), .B(n4078), .Z(n4041) );
  XNOR U4164 ( .A(n4079), .B(n4080), .Z(n4078) );
  XNOR U4165 ( .A(n4081), .B(n4082), .Z(n4079) );
  XOR U4166 ( .A(n4083), .B(n4084), .Z(n4082) );
  AND U4167 ( .A(b[7]), .B(a[15]), .Z(n4084) );
  AND U4168 ( .A(b[6]), .B(a[16]), .Z(n4083) );
  XNOR U4169 ( .A(n4085), .B(n4081), .Z(n4077) );
  XOR U4170 ( .A(n4086), .B(n4087), .Z(n4081) );
  NOR U4171 ( .A(n4088), .B(n4089), .Z(n4086) );
  AND U4172 ( .A(b[5]), .B(a[17]), .Z(n4085) );
  XOR U4173 ( .A(n4090), .B(n4039), .Z(n4040) );
  IV U4174 ( .A(n4080), .Z(n4039) );
  XOR U4175 ( .A(n4091), .B(n4092), .Z(n4080) );
  ANDN U4176 ( .B(n4067), .A(n4076), .Z(n4091) );
  AND U4177 ( .A(b[3]), .B(a[18]), .Z(n4093) );
  XOR U4178 ( .A(n4089), .B(n4092), .Z(n4094) );
  XOR U4179 ( .A(n4095), .B(n4096), .Z(n4092) );
  ANDN U4180 ( .B(n4072), .A(n4073), .Z(n4095) );
  AND U4181 ( .A(b[2]), .B(a[18]), .Z(n4097) );
  XNOR U4182 ( .A(n4099), .B(n4096), .Z(n4098) );
  XOR U4183 ( .A(n4100), .B(n4101), .Z(n4096) );
  NANDN U4184 ( .A(n4075), .B(n4074), .Z(n4101) );
  XOR U4185 ( .A(n4100), .B(n4102), .Z(n4074) );
  NAND U4186 ( .A(b[1]), .B(a[18]), .Z(n4102) );
  XOR U4187 ( .A(n4100), .B(n4104), .Z(n4103) );
  OR U4188 ( .A(n1517), .B(n1515), .Z(n4100) );
  XOR U4189 ( .A(n4106), .B(n4107), .Z(n1515) );
  NANDN U4190 ( .A(n187), .B(a[18]), .Z(n1517) );
  XOR U4191 ( .A(n4109), .B(n4110), .Z(n4089) );
  XNOR U4192 ( .A(n4111), .B(n4112), .Z(n4110) );
  XNOR U4193 ( .A(n4113), .B(n4114), .Z(n4111) );
  XOR U4194 ( .A(n4115), .B(n4116), .Z(n4114) );
  AND U4195 ( .A(b[6]), .B(a[15]), .Z(n4116) );
  AND U4196 ( .A(b[7]), .B(a[14]), .Z(n4115) );
  XNOR U4197 ( .A(n4117), .B(n4113), .Z(n4109) );
  XOR U4198 ( .A(n4118), .B(n4119), .Z(n4113) );
  NOR U4199 ( .A(n4120), .B(n4121), .Z(n4118) );
  AND U4200 ( .A(b[5]), .B(a[16]), .Z(n4117) );
  XOR U4201 ( .A(n4122), .B(n4087), .Z(n4088) );
  IV U4202 ( .A(n4112), .Z(n4087) );
  XOR U4203 ( .A(n4123), .B(n4124), .Z(n4112) );
  ANDN U4204 ( .B(n4099), .A(n4108), .Z(n4123) );
  AND U4205 ( .A(b[3]), .B(a[17]), .Z(n4125) );
  XOR U4206 ( .A(n4121), .B(n4124), .Z(n4126) );
  XOR U4207 ( .A(n4127), .B(n4128), .Z(n4124) );
  ANDN U4208 ( .B(n4104), .A(n4105), .Z(n4127) );
  AND U4209 ( .A(b[2]), .B(a[17]), .Z(n4129) );
  XOR U4210 ( .A(n4131), .B(n4128), .Z(n4130) );
  XOR U4211 ( .A(n4132), .B(n4133), .Z(n4128) );
  NANDN U4212 ( .A(n4107), .B(n4106), .Z(n4133) );
  XOR U4213 ( .A(n4132), .B(n4134), .Z(n4106) );
  NAND U4214 ( .A(b[1]), .B(a[17]), .Z(n4134) );
  XOR U4215 ( .A(n4132), .B(n4136), .Z(n4135) );
  OR U4216 ( .A(n1522), .B(n1520), .Z(n4132) );
  XOR U4217 ( .A(n4138), .B(n4139), .Z(n1520) );
  NANDN U4218 ( .A(n187), .B(a[17]), .Z(n1522) );
  XOR U4219 ( .A(n4141), .B(n4142), .Z(n4121) );
  XNOR U4220 ( .A(n4143), .B(n4144), .Z(n4142) );
  XOR U4221 ( .A(n4145), .B(n4146), .Z(n4143) );
  AND U4222 ( .A(b[5]), .B(a[15]), .Z(n4145) );
  XOR U4223 ( .A(n4146), .B(n4147), .Z(n4141) );
  XOR U4224 ( .A(n4148), .B(n4149), .Z(n4147) );
  AND U4225 ( .A(b[6]), .B(a[14]), .Z(n4149) );
  AND U4226 ( .A(b[7]), .B(a[13]), .Z(n4148) );
  XOR U4227 ( .A(n4150), .B(n4151), .Z(n4146) );
  ANDN U4228 ( .B(n4152), .A(n4153), .Z(n4150) );
  XOR U4229 ( .A(n4154), .B(n4119), .Z(n4120) );
  IV U4230 ( .A(n4144), .Z(n4119) );
  XOR U4231 ( .A(n4155), .B(n4156), .Z(n4144) );
  NOR U4232 ( .A(n4140), .B(n4131), .Z(n4155) );
  XNOR U4233 ( .A(n4153), .B(n4157), .Z(n4131) );
  XNOR U4234 ( .A(n4152), .B(n4156), .Z(n4157) );
  XOR U4235 ( .A(n4158), .B(n4151), .Z(n4152) );
  AND U4236 ( .A(b[4]), .B(a[15]), .Z(n4158) );
  XOR U4237 ( .A(n4159), .B(n4160), .Z(n4153) );
  XOR U4238 ( .A(n4151), .B(n4161), .Z(n4160) );
  XOR U4239 ( .A(n4162), .B(n4163), .Z(n4161) );
  XOR U4240 ( .A(n4164), .B(n4165), .Z(n4163) );
  NAND U4241 ( .A(b[6]), .B(a[13]), .Z(n4165) );
  AND U4242 ( .A(b[7]), .B(a[12]), .Z(n4164) );
  XOR U4243 ( .A(n4166), .B(n4167), .Z(n4151) );
  ANDN U4244 ( .B(n4168), .A(n4169), .Z(n4166) );
  XOR U4245 ( .A(n4170), .B(n4162), .Z(n4159) );
  XOR U4246 ( .A(n4171), .B(n4172), .Z(n4162) );
  NOR U4247 ( .A(n4173), .B(n4174), .Z(n4171) );
  AND U4248 ( .A(b[5]), .B(a[14]), .Z(n4170) );
  XOR U4249 ( .A(n4176), .B(n4177), .Z(n4156) );
  ANDN U4250 ( .B(n4136), .A(n4137), .Z(n4176) );
  AND U4251 ( .A(b[2]), .B(a[16]), .Z(n4178) );
  XNOR U4252 ( .A(n4168), .B(n4177), .Z(n4179) );
  XOR U4253 ( .A(n4180), .B(n4181), .Z(n4177) );
  NANDN U4254 ( .A(n4139), .B(n4138), .Z(n4181) );
  XOR U4255 ( .A(n4180), .B(n4182), .Z(n4138) );
  NAND U4256 ( .A(b[1]), .B(a[16]), .Z(n4182) );
  XNOR U4257 ( .A(n4180), .B(n4184), .Z(n4183) );
  OR U4258 ( .A(n1527), .B(n1525), .Z(n4180) );
  NANDN U4259 ( .A(n187), .B(a[16]), .Z(n1527) );
  XOR U4260 ( .A(n4188), .B(n4167), .Z(n4168) );
  AND U4261 ( .A(b[3]), .B(a[15]), .Z(n4188) );
  XOR U4262 ( .A(n4167), .B(n4174), .Z(n4189) );
  XOR U4263 ( .A(n4190), .B(n4191), .Z(n4174) );
  XOR U4264 ( .A(n4172), .B(n4192), .Z(n4191) );
  XOR U4265 ( .A(n4193), .B(n4194), .Z(n4192) );
  XOR U4266 ( .A(n4195), .B(n4196), .Z(n4194) );
  NAND U4267 ( .A(b[6]), .B(a[12]), .Z(n4196) );
  AND U4268 ( .A(b[7]), .B(a[11]), .Z(n4195) );
  XOR U4269 ( .A(n4197), .B(n4193), .Z(n4190) );
  XOR U4270 ( .A(n4198), .B(n4199), .Z(n4193) );
  NOR U4271 ( .A(n4200), .B(n4201), .Z(n4198) );
  AND U4272 ( .A(b[5]), .B(a[13]), .Z(n4197) );
  XNOR U4273 ( .A(n4202), .B(n4203), .Z(n4167) );
  NOR U4274 ( .A(n4185), .B(n4184), .Z(n4202) );
  XOR U4275 ( .A(n4204), .B(n4203), .Z(n4184) );
  AND U4276 ( .A(b[2]), .B(a[15]), .Z(n4204) );
  XOR U4277 ( .A(n4203), .B(n4206), .Z(n4205) );
  XNOR U4278 ( .A(n4207), .B(n4208), .Z(n4203) );
  OR U4279 ( .A(n4186), .B(n4187), .Z(n4208) );
  XNOR U4280 ( .A(n4207), .B(n4210), .Z(n4209) );
  XNOR U4281 ( .A(n4207), .B(n4212), .Z(n4186) );
  NAND U4282 ( .A(b[1]), .B(a[15]), .Z(n4212) );
  OR U4283 ( .A(n1532), .B(n1530), .Z(n4207) );
  XOR U4284 ( .A(n4213), .B(n4214), .Z(n1530) );
  NANDN U4285 ( .A(n187), .B(a[15]), .Z(n1532) );
  XNOR U4286 ( .A(n4216), .B(n4172), .Z(n4173) );
  XOR U4287 ( .A(n4217), .B(n4218), .Z(n4172) );
  ANDN U4288 ( .B(n4206), .A(n4215), .Z(n4217) );
  XNOR U4289 ( .A(n4219), .B(n4218), .Z(n4215) );
  AND U4290 ( .A(b[3]), .B(a[14]), .Z(n4219) );
  XOR U4291 ( .A(n4218), .B(n4201), .Z(n4220) );
  XOR U4292 ( .A(n4221), .B(n4222), .Z(n4201) );
  XOR U4293 ( .A(n4199), .B(n4223), .Z(n4222) );
  XOR U4294 ( .A(n4224), .B(n4225), .Z(n4223) );
  XOR U4295 ( .A(n4226), .B(n4227), .Z(n4225) );
  NAND U4296 ( .A(b[6]), .B(a[11]), .Z(n4227) );
  AND U4297 ( .A(b[7]), .B(a[10]), .Z(n4226) );
  XOR U4298 ( .A(n4228), .B(n4224), .Z(n4221) );
  XOR U4299 ( .A(n4229), .B(n4230), .Z(n4224) );
  NOR U4300 ( .A(n4231), .B(n4232), .Z(n4229) );
  AND U4301 ( .A(b[5]), .B(a[12]), .Z(n4228) );
  XNOR U4302 ( .A(n4233), .B(n4234), .Z(n4218) );
  NOR U4303 ( .A(n4211), .B(n4210), .Z(n4233) );
  XOR U4304 ( .A(n4235), .B(n4234), .Z(n4210) );
  AND U4305 ( .A(b[2]), .B(a[14]), .Z(n4235) );
  XOR U4306 ( .A(n4234), .B(n4237), .Z(n4236) );
  XNOR U4307 ( .A(n4238), .B(n4239), .Z(n4234) );
  NANDN U4308 ( .A(n4214), .B(n4213), .Z(n4239) );
  XOR U4309 ( .A(n4238), .B(n4240), .Z(n4213) );
  NAND U4310 ( .A(b[1]), .B(a[14]), .Z(n4240) );
  XOR U4311 ( .A(n4238), .B(n4242), .Z(n4241) );
  OR U4312 ( .A(n1537), .B(n1535), .Z(n4238) );
  XOR U4313 ( .A(n4244), .B(n4245), .Z(n1535) );
  NANDN U4314 ( .A(n187), .B(a[14]), .Z(n1537) );
  XNOR U4315 ( .A(n4247), .B(n4199), .Z(n4200) );
  XOR U4316 ( .A(n4248), .B(n4249), .Z(n4199) );
  ANDN U4317 ( .B(n4237), .A(n4246), .Z(n4248) );
  XNOR U4318 ( .A(n4250), .B(n4249), .Z(n4246) );
  AND U4319 ( .A(b[3]), .B(a[13]), .Z(n4250) );
  XOR U4320 ( .A(n4249), .B(n4232), .Z(n4251) );
  XOR U4321 ( .A(n4252), .B(n4253), .Z(n4232) );
  XOR U4322 ( .A(n4230), .B(n4254), .Z(n4253) );
  XNOR U4323 ( .A(n4255), .B(n4256), .Z(n4254) );
  XOR U4324 ( .A(n4257), .B(n4258), .Z(n4256) );
  NAND U4325 ( .A(b[6]), .B(a[10]), .Z(n4258) );
  AND U4326 ( .A(b[7]), .B(a[9]), .Z(n4257) );
  XNOR U4327 ( .A(n4259), .B(n4255), .Z(n4252) );
  XOR U4328 ( .A(n4260), .B(n4261), .Z(n4255) );
  NOR U4329 ( .A(n4262), .B(n4263), .Z(n4260) );
  AND U4330 ( .A(b[5]), .B(a[11]), .Z(n4259) );
  XNOR U4331 ( .A(n4264), .B(n4265), .Z(n4249) );
  ANDN U4332 ( .B(n4242), .A(n4243), .Z(n4264) );
  XOR U4333 ( .A(n4266), .B(n4265), .Z(n4243) );
  IV U4334 ( .A(n4267), .Z(n4265) );
  AND U4335 ( .A(b[2]), .B(a[13]), .Z(n4266) );
  XNOR U4336 ( .A(n4269), .B(n4267), .Z(n4268) );
  XOR U4337 ( .A(n4270), .B(n4271), .Z(n4267) );
  NANDN U4338 ( .A(n4245), .B(n4244), .Z(n4271) );
  XOR U4339 ( .A(n4270), .B(n4272), .Z(n4244) );
  NAND U4340 ( .A(b[1]), .B(a[13]), .Z(n4272) );
  XOR U4341 ( .A(n4270), .B(n4274), .Z(n4273) );
  OR U4342 ( .A(n1542), .B(n1540), .Z(n4270) );
  XOR U4343 ( .A(n4276), .B(n4277), .Z(n1540) );
  NANDN U4344 ( .A(n187), .B(a[13]), .Z(n1542) );
  XNOR U4345 ( .A(n4279), .B(n4230), .Z(n4231) );
  XNOR U4346 ( .A(n4280), .B(n4281), .Z(n4230) );
  ANDN U4347 ( .B(n4269), .A(n4278), .Z(n4280) );
  XOR U4348 ( .A(n4282), .B(n4281), .Z(n4278) );
  IV U4349 ( .A(n4283), .Z(n4281) );
  AND U4350 ( .A(b[3]), .B(a[12]), .Z(n4282) );
  XOR U4351 ( .A(n4263), .B(n4283), .Z(n4284) );
  XOR U4352 ( .A(n4285), .B(n4286), .Z(n4283) );
  ANDN U4353 ( .B(n4274), .A(n4275), .Z(n4285) );
  AND U4354 ( .A(b[2]), .B(a[12]), .Z(n4287) );
  XNOR U4355 ( .A(n4289), .B(n4286), .Z(n4288) );
  XOR U4356 ( .A(n4290), .B(n4291), .Z(n4286) );
  NANDN U4357 ( .A(n4277), .B(n4276), .Z(n4291) );
  XOR U4358 ( .A(n4290), .B(n4292), .Z(n4276) );
  NAND U4359 ( .A(b[1]), .B(a[12]), .Z(n4292) );
  XOR U4360 ( .A(n4290), .B(n4294), .Z(n4293) );
  OR U4361 ( .A(n1547), .B(n1545), .Z(n4290) );
  XOR U4362 ( .A(n4296), .B(n4297), .Z(n1545) );
  NANDN U4363 ( .A(n187), .B(a[12]), .Z(n1547) );
  XOR U4364 ( .A(n4299), .B(n4300), .Z(n4263) );
  XNOR U4365 ( .A(n4301), .B(n4302), .Z(n4300) );
  XNOR U4366 ( .A(n4303), .B(n4304), .Z(n4301) );
  XOR U4367 ( .A(n4305), .B(n4306), .Z(n4304) );
  AND U4368 ( .A(b[7]), .B(a[8]), .Z(n4306) );
  AND U4369 ( .A(b[6]), .B(a[9]), .Z(n4305) );
  XNOR U4370 ( .A(n4307), .B(n4303), .Z(n4299) );
  XOR U4371 ( .A(n4308), .B(n4309), .Z(n4303) );
  NOR U4372 ( .A(n4310), .B(n4311), .Z(n4308) );
  AND U4373 ( .A(b[5]), .B(a[10]), .Z(n4307) );
  XOR U4374 ( .A(n4312), .B(n4261), .Z(n4262) );
  IV U4375 ( .A(n4302), .Z(n4261) );
  XOR U4376 ( .A(n4313), .B(n4314), .Z(n4302) );
  ANDN U4377 ( .B(n4289), .A(n4298), .Z(n4313) );
  AND U4378 ( .A(b[3]), .B(a[11]), .Z(n4315) );
  XOR U4379 ( .A(n4311), .B(n4314), .Z(n4316) );
  XOR U4380 ( .A(n4317), .B(n4318), .Z(n4314) );
  ANDN U4381 ( .B(n4294), .A(n4295), .Z(n4317) );
  AND U4382 ( .A(b[2]), .B(a[11]), .Z(n4319) );
  XNOR U4383 ( .A(n4321), .B(n4318), .Z(n4320) );
  XOR U4384 ( .A(n4322), .B(n4323), .Z(n4318) );
  NANDN U4385 ( .A(n4297), .B(n4296), .Z(n4323) );
  XOR U4386 ( .A(n4322), .B(n4324), .Z(n4296) );
  NAND U4387 ( .A(b[1]), .B(a[11]), .Z(n4324) );
  XOR U4388 ( .A(n4322), .B(n4326), .Z(n4325) );
  OR U4389 ( .A(n1552), .B(n1550), .Z(n4322) );
  XOR U4390 ( .A(n4328), .B(n4329), .Z(n1550) );
  NANDN U4391 ( .A(n187), .B(a[11]), .Z(n1552) );
  XOR U4392 ( .A(n4331), .B(n4332), .Z(n4311) );
  XNOR U4393 ( .A(n4333), .B(n4334), .Z(n4332) );
  XNOR U4394 ( .A(n4335), .B(n4336), .Z(n4333) );
  XOR U4395 ( .A(n4337), .B(n4338), .Z(n4336) );
  AND U4396 ( .A(b[6]), .B(a[8]), .Z(n4338) );
  AND U4397 ( .A(a[7]), .B(b[7]), .Z(n4337) );
  XNOR U4398 ( .A(n4339), .B(n4335), .Z(n4331) );
  XOR U4399 ( .A(n4340), .B(n4341), .Z(n4335) );
  NOR U4400 ( .A(n4342), .B(n4343), .Z(n4340) );
  AND U4401 ( .A(b[5]), .B(a[9]), .Z(n4339) );
  XOR U4402 ( .A(n4344), .B(n4309), .Z(n4310) );
  IV U4403 ( .A(n4334), .Z(n4309) );
  XOR U4404 ( .A(n4345), .B(n4346), .Z(n4334) );
  ANDN U4405 ( .B(n4321), .A(n4330), .Z(n4345) );
  AND U4406 ( .A(b[3]), .B(a[10]), .Z(n4347) );
  XOR U4407 ( .A(n4343), .B(n4346), .Z(n4348) );
  XOR U4408 ( .A(n4349), .B(n4350), .Z(n4346) );
  ANDN U4409 ( .B(n4326), .A(n4327), .Z(n4349) );
  AND U4410 ( .A(b[2]), .B(a[10]), .Z(n4351) );
  XOR U4411 ( .A(n4353), .B(n4350), .Z(n4352) );
  XOR U4412 ( .A(n4354), .B(n4355), .Z(n4350) );
  NANDN U4413 ( .A(n4329), .B(n4328), .Z(n4355) );
  XOR U4414 ( .A(n4354), .B(n4356), .Z(n4328) );
  NAND U4415 ( .A(b[1]), .B(a[10]), .Z(n4356) );
  XOR U4416 ( .A(n4354), .B(n4358), .Z(n4357) );
  OR U4417 ( .A(n1557), .B(n1555), .Z(n4354) );
  XOR U4418 ( .A(n4360), .B(n4361), .Z(n1555) );
  NANDN U4419 ( .A(n187), .B(a[10]), .Z(n1557) );
  XOR U4420 ( .A(n4363), .B(n4364), .Z(n4343) );
  XNOR U4421 ( .A(n4365), .B(n4366), .Z(n4364) );
  XOR U4422 ( .A(n4367), .B(n4368), .Z(n4365) );
  AND U4423 ( .A(b[5]), .B(a[8]), .Z(n4367) );
  XOR U4424 ( .A(n4368), .B(n4369), .Z(n4363) );
  XOR U4425 ( .A(n4370), .B(n4371), .Z(n4369) );
  AND U4426 ( .A(a[7]), .B(b[6]), .Z(n4371) );
  AND U4427 ( .A(a[6]), .B(b[7]), .Z(n4370) );
  XOR U4428 ( .A(n4372), .B(n4373), .Z(n4368) );
  ANDN U4429 ( .B(n4374), .A(n4375), .Z(n4372) );
  XOR U4430 ( .A(n4376), .B(n4341), .Z(n4342) );
  IV U4431 ( .A(n4366), .Z(n4341) );
  XOR U4432 ( .A(n4377), .B(n4378), .Z(n4366) );
  NOR U4433 ( .A(n4362), .B(n4353), .Z(n4377) );
  XNOR U4434 ( .A(n4375), .B(n4379), .Z(n4353) );
  XNOR U4435 ( .A(n4374), .B(n4378), .Z(n4379) );
  XOR U4436 ( .A(n4380), .B(n4373), .Z(n4374) );
  AND U4437 ( .A(b[4]), .B(a[8]), .Z(n4380) );
  XOR U4438 ( .A(n4381), .B(n4382), .Z(n4375) );
  XOR U4439 ( .A(n4373), .B(n4383), .Z(n4382) );
  XOR U4440 ( .A(n4384), .B(n4385), .Z(n4383) );
  XOR U4441 ( .A(n4386), .B(n4387), .Z(n4385) );
  NAND U4442 ( .A(b[6]), .B(a[6]), .Z(n4387) );
  AND U4443 ( .A(a[5]), .B(b[7]), .Z(n4386) );
  XOR U4444 ( .A(n4388), .B(n4389), .Z(n4373) );
  ANDN U4445 ( .B(n4390), .A(n4391), .Z(n4388) );
  XOR U4446 ( .A(n4392), .B(n4384), .Z(n4381) );
  XOR U4447 ( .A(n4393), .B(n4394), .Z(n4384) );
  NOR U4448 ( .A(n4395), .B(n4396), .Z(n4393) );
  AND U4449 ( .A(a[7]), .B(b[5]), .Z(n4392) );
  XOR U4450 ( .A(n4398), .B(n4399), .Z(n4378) );
  ANDN U4451 ( .B(n4358), .A(n4359), .Z(n4398) );
  AND U4452 ( .A(b[2]), .B(a[9]), .Z(n4400) );
  XNOR U4453 ( .A(n4390), .B(n4399), .Z(n4401) );
  XOR U4454 ( .A(n4402), .B(n4403), .Z(n4399) );
  NANDN U4455 ( .A(n4361), .B(n4360), .Z(n4403) );
  XOR U4456 ( .A(n4402), .B(n4404), .Z(n4360) );
  NAND U4457 ( .A(b[1]), .B(a[9]), .Z(n4404) );
  XNOR U4458 ( .A(n4402), .B(n4406), .Z(n4405) );
  OR U4459 ( .A(n1562), .B(n1560), .Z(n4402) );
  NANDN U4460 ( .A(n187), .B(a[9]), .Z(n1562) );
  XOR U4461 ( .A(n4410), .B(n4389), .Z(n4390) );
  AND U4462 ( .A(b[3]), .B(a[8]), .Z(n4410) );
  XOR U4463 ( .A(n4389), .B(n4396), .Z(n4411) );
  XOR U4464 ( .A(n4412), .B(n4413), .Z(n4396) );
  XOR U4465 ( .A(n4394), .B(n4414), .Z(n4413) );
  XOR U4466 ( .A(n4415), .B(n4416), .Z(n4414) );
  XOR U4467 ( .A(n4417), .B(n4418), .Z(n4416) );
  NAND U4468 ( .A(a[5]), .B(b[6]), .Z(n4418) );
  AND U4469 ( .A(a[4]), .B(b[7]), .Z(n4417) );
  XOR U4470 ( .A(n4419), .B(n4415), .Z(n4412) );
  XOR U4471 ( .A(n4420), .B(n4421), .Z(n4415) );
  NOR U4472 ( .A(n4422), .B(n4423), .Z(n4420) );
  AND U4473 ( .A(b[5]), .B(a[6]), .Z(n4419) );
  XNOR U4474 ( .A(n4424), .B(n4425), .Z(n4389) );
  NOR U4475 ( .A(n4407), .B(n4406), .Z(n4424) );
  XOR U4476 ( .A(n4426), .B(n4425), .Z(n4406) );
  AND U4477 ( .A(b[2]), .B(a[8]), .Z(n4426) );
  XOR U4478 ( .A(n4425), .B(n4428), .Z(n4427) );
  XNOR U4479 ( .A(n4429), .B(n4430), .Z(n4425) );
  OR U4480 ( .A(n4408), .B(n4409), .Z(n4430) );
  XNOR U4481 ( .A(n4429), .B(n4432), .Z(n4431) );
  XNOR U4482 ( .A(n4429), .B(n4434), .Z(n4408) );
  NAND U4483 ( .A(b[1]), .B(a[8]), .Z(n4434) );
  OR U4484 ( .A(n1567), .B(n1565), .Z(n4429) );
  XOR U4485 ( .A(n4435), .B(n4436), .Z(n1565) );
  NANDN U4486 ( .A(n187), .B(a[8]), .Z(n1567) );
  XNOR U4487 ( .A(n4438), .B(n4394), .Z(n4395) );
  XOR U4488 ( .A(n4439), .B(n4440), .Z(n4394) );
  ANDN U4489 ( .B(n4428), .A(n4437), .Z(n4439) );
  XNOR U4490 ( .A(n4441), .B(n4440), .Z(n4437) );
  AND U4491 ( .A(a[7]), .B(b[3]), .Z(n4441) );
  XOR U4492 ( .A(n4440), .B(n4423), .Z(n4442) );
  XOR U4493 ( .A(n4443), .B(n4444), .Z(n4423) );
  XOR U4494 ( .A(n4421), .B(n4445), .Z(n4444) );
  XOR U4495 ( .A(n4446), .B(n4447), .Z(n4445) );
  XOR U4496 ( .A(n4448), .B(n4449), .Z(n4447) );
  NAND U4497 ( .A(a[4]), .B(b[6]), .Z(n4449) );
  AND U4498 ( .A(a[3]), .B(b[7]), .Z(n4448) );
  XOR U4499 ( .A(n4450), .B(n4446), .Z(n4443) );
  XOR U4500 ( .A(n4451), .B(n4452), .Z(n4446) );
  NOR U4501 ( .A(n4453), .B(n4454), .Z(n4451) );
  AND U4502 ( .A(a[5]), .B(b[5]), .Z(n4450) );
  XNOR U4503 ( .A(n4455), .B(n4456), .Z(n4440) );
  NOR U4504 ( .A(n4433), .B(n4432), .Z(n4455) );
  XOR U4505 ( .A(n4457), .B(n4456), .Z(n4432) );
  AND U4506 ( .A(a[7]), .B(b[2]), .Z(n4457) );
  XOR U4507 ( .A(n4456), .B(n4459), .Z(n4458) );
  XNOR U4508 ( .A(n4460), .B(n4461), .Z(n4456) );
  NANDN U4509 ( .A(n4436), .B(n4435), .Z(n4461) );
  XOR U4510 ( .A(n4460), .B(n4462), .Z(n4435) );
  NAND U4511 ( .A(a[7]), .B(b[1]), .Z(n4462) );
  XOR U4512 ( .A(n4460), .B(n4464), .Z(n4463) );
  OR U4513 ( .A(n4466), .B(n4467), .Z(n4460) );
  XNOR U4514 ( .A(n4469), .B(n4421), .Z(n4422) );
  XOR U4515 ( .A(n4470), .B(n4471), .Z(n4421) );
  ANDN U4516 ( .B(n4459), .A(n4468), .Z(n4470) );
  XNOR U4517 ( .A(n4472), .B(n4471), .Z(n4468) );
  AND U4518 ( .A(b[3]), .B(a[6]), .Z(n4472) );
  XOR U4519 ( .A(n4471), .B(n4454), .Z(n4473) );
  XOR U4520 ( .A(n4474), .B(n4475), .Z(n4454) );
  XOR U4521 ( .A(n4452), .B(n4476), .Z(n4475) );
  XNOR U4522 ( .A(n4477), .B(n4478), .Z(n4476) );
  XOR U4523 ( .A(n4479), .B(n4480), .Z(n4478) );
  NAND U4524 ( .A(a[3]), .B(b[6]), .Z(n4480) );
  AND U4525 ( .A(a[2]), .B(b[7]), .Z(n4479) );
  XNOR U4526 ( .A(n4481), .B(n4477), .Z(n4474) );
  XNOR U4527 ( .A(n4482), .B(n4483), .Z(n4477) );
  NOR U4528 ( .A(n4484), .B(n4485), .Z(n4482) );
  AND U4529 ( .A(a[4]), .B(b[5]), .Z(n4481) );
  XNOR U4530 ( .A(n4486), .B(n4487), .Z(n4471) );
  ANDN U4531 ( .B(n4464), .A(n4465), .Z(n4486) );
  XOR U4532 ( .A(n4488), .B(n4487), .Z(n4465) );
  IV U4533 ( .A(n4489), .Z(n4487) );
  AND U4534 ( .A(b[2]), .B(a[6]), .Z(n4488) );
  XNOR U4535 ( .A(n4491), .B(n4489), .Z(n4490) );
  XOR U4536 ( .A(n4492), .B(n4493), .Z(n4489) );
  OR U4537 ( .A(n4494), .B(n4495), .Z(n4493) );
  XNOR U4538 ( .A(n4497), .B(n4452), .Z(n4453) );
  XOR U4539 ( .A(n4498), .B(n4499), .Z(n4452) );
  ANDN U4540 ( .B(n4491), .A(n4496), .Z(n4498) );
  XNOR U4541 ( .A(n4500), .B(n4499), .Z(n4496) );
  AND U4542 ( .A(a[5]), .B(b[3]), .Z(n4500) );
  XOR U4543 ( .A(n4485), .B(n4499), .Z(n4501) );
  XNOR U4544 ( .A(n4502), .B(n4503), .Z(n4499) );
  NOR U4545 ( .A(n4504), .B(n4505), .Z(n4502) );
  XOR U4546 ( .A(n4506), .B(n4507), .Z(n4485) );
  XNOR U4547 ( .A(n4508), .B(n4483), .Z(n4507) );
  XOR U4548 ( .A(n4509), .B(n4510), .Z(n4508) );
  XOR U4549 ( .A(n4511), .B(n4512), .Z(n4510) );
  AND U4550 ( .A(a[1]), .B(b[7]), .Z(n4512) );
  AND U4551 ( .A(a[2]), .B(b[6]), .Z(n4511) );
  XOR U4552 ( .A(n4513), .B(n4509), .Z(n4506) );
  XOR U4553 ( .A(n4514), .B(n4515), .Z(n4509) );
  NOR U4554 ( .A(n4516), .B(n4517), .Z(n4514) );
  AND U4555 ( .A(a[3]), .B(b[5]), .Z(n4513) );
  XNOR U4556 ( .A(n4518), .B(n4483), .Z(n4484) );
  XOR U4557 ( .A(n4519), .B(n4520), .Z(n4483) );
  ANDN U4558 ( .B(n4521), .A(n4522), .Z(n4519) );
  AND U4559 ( .A(b[4]), .B(a[4]), .Z(n4518) );
  AND U4560 ( .A(a[5]), .B(b[4]), .Z(n4497) );
  AND U4561 ( .A(b[4]), .B(a[6]), .Z(n4469) );
  AND U4562 ( .A(a[7]), .B(b[4]), .Z(n4438) );
  AND U4563 ( .A(b[3]), .B(a[9]), .Z(n4397) );
  AND U4564 ( .A(b[4]), .B(a[9]), .Z(n4376) );
  AND U4565 ( .A(b[4]), .B(a[10]), .Z(n4344) );
  AND U4566 ( .A(b[4]), .B(a[11]), .Z(n4312) );
  AND U4567 ( .A(b[4]), .B(a[12]), .Z(n4279) );
  AND U4568 ( .A(b[4]), .B(a[13]), .Z(n4247) );
  AND U4569 ( .A(b[4]), .B(a[14]), .Z(n4216) );
  AND U4570 ( .A(b[3]), .B(a[16]), .Z(n4175) );
  AND U4571 ( .A(b[4]), .B(a[16]), .Z(n4154) );
  AND U4572 ( .A(b[4]), .B(a[17]), .Z(n4122) );
  AND U4573 ( .A(b[4]), .B(a[18]), .Z(n4090) );
  AND U4574 ( .A(b[4]), .B(a[19]), .Z(n4057) );
  AND U4575 ( .A(b[4]), .B(a[20]), .Z(n4025) );
  AND U4576 ( .A(b[4]), .B(a[21]), .Z(n3994) );
  AND U4577 ( .A(b[3]), .B(a[23]), .Z(n3953) );
  AND U4578 ( .A(b[4]), .B(a[23]), .Z(n3932) );
  AND U4579 ( .A(b[4]), .B(a[24]), .Z(n3900) );
  AND U4580 ( .A(b[4]), .B(a[25]), .Z(n3868) );
  AND U4581 ( .A(b[4]), .B(a[26]), .Z(n3835) );
  AND U4582 ( .A(b[4]), .B(a[27]), .Z(n3803) );
  AND U4583 ( .A(b[4]), .B(a[28]), .Z(n3772) );
  AND U4584 ( .A(b[3]), .B(a[30]), .Z(n3731) );
  AND U4585 ( .A(b[4]), .B(a[30]), .Z(n3710) );
  AND U4586 ( .A(b[4]), .B(a[31]), .Z(n3678) );
  AND U4587 ( .A(b[4]), .B(a[32]), .Z(n3646) );
  AND U4588 ( .A(b[4]), .B(a[33]), .Z(n3613) );
  AND U4589 ( .A(b[4]), .B(a[34]), .Z(n3581) );
  AND U4590 ( .A(b[4]), .B(a[35]), .Z(n3550) );
  AND U4591 ( .A(b[3]), .B(a[37]), .Z(n3509) );
  AND U4592 ( .A(b[4]), .B(a[37]), .Z(n3488) );
  AND U4593 ( .A(b[4]), .B(a[38]), .Z(n3456) );
  AND U4594 ( .A(b[4]), .B(a[39]), .Z(n3424) );
  AND U4595 ( .A(b[4]), .B(a[40]), .Z(n3391) );
  AND U4596 ( .A(b[4]), .B(a[41]), .Z(n3359) );
  AND U4597 ( .A(b[4]), .B(a[42]), .Z(n3328) );
  AND U4598 ( .A(b[3]), .B(a[44]), .Z(n3287) );
  AND U4599 ( .A(b[4]), .B(a[44]), .Z(n3266) );
  AND U4600 ( .A(b[4]), .B(a[45]), .Z(n3234) );
  AND U4601 ( .A(b[4]), .B(a[46]), .Z(n3202) );
  AND U4602 ( .A(b[4]), .B(a[47]), .Z(n3169) );
  AND U4603 ( .A(b[4]), .B(a[48]), .Z(n3137) );
  AND U4604 ( .A(b[4]), .B(a[49]), .Z(n3106) );
  AND U4605 ( .A(b[3]), .B(a[51]), .Z(n3065) );
  AND U4606 ( .A(b[4]), .B(a[51]), .Z(n3044) );
  AND U4607 ( .A(b[4]), .B(a[52]), .Z(n3012) );
  AND U4608 ( .A(b[4]), .B(a[53]), .Z(n2980) );
  AND U4609 ( .A(b[4]), .B(a[54]), .Z(n2947) );
  AND U4610 ( .A(b[4]), .B(a[55]), .Z(n2915) );
  AND U4611 ( .A(b[4]), .B(a[56]), .Z(n2884) );
  AND U4612 ( .A(b[3]), .B(a[58]), .Z(n2843) );
  AND U4613 ( .A(b[4]), .B(a[58]), .Z(n2822) );
  AND U4614 ( .A(b[4]), .B(a[59]), .Z(n2790) );
  AND U4615 ( .A(b[4]), .B(a[60]), .Z(n2758) );
  AND U4616 ( .A(b[4]), .B(a[61]), .Z(n2725) );
  AND U4617 ( .A(b[4]), .B(a[62]), .Z(n2693) );
  AND U4618 ( .A(b[4]), .B(a[63]), .Z(n2662) );
  AND U4619 ( .A(b[3]), .B(a[65]), .Z(n2621) );
  AND U4620 ( .A(b[4]), .B(a[65]), .Z(n2600) );
  AND U4621 ( .A(b[4]), .B(a[66]), .Z(n2568) );
  AND U4622 ( .A(b[4]), .B(a[67]), .Z(n2536) );
  AND U4623 ( .A(b[4]), .B(a[68]), .Z(n2503) );
  AND U4624 ( .A(b[4]), .B(a[69]), .Z(n2471) );
  AND U4625 ( .A(b[4]), .B(a[70]), .Z(n2440) );
  AND U4626 ( .A(b[3]), .B(a[72]), .Z(n2399) );
  AND U4627 ( .A(b[4]), .B(a[72]), .Z(n2378) );
  AND U4628 ( .A(b[4]), .B(a[73]), .Z(n2346) );
  AND U4629 ( .A(b[4]), .B(a[74]), .Z(n2314) );
  AND U4630 ( .A(b[4]), .B(a[75]), .Z(n2281) );
  AND U4631 ( .A(b[4]), .B(a[76]), .Z(n2249) );
  AND U4632 ( .A(b[4]), .B(a[77]), .Z(n2218) );
  AND U4633 ( .A(b[3]), .B(a[79]), .Z(n2177) );
  AND U4634 ( .A(b[4]), .B(a[79]), .Z(n2156) );
  AND U4635 ( .A(b[4]), .B(a[80]), .Z(n2124) );
  AND U4636 ( .A(b[4]), .B(a[81]), .Z(n2092) );
  AND U4637 ( .A(b[4]), .B(a[82]), .Z(n2059) );
  AND U4638 ( .A(b[4]), .B(a[83]), .Z(n2027) );
  AND U4639 ( .A(b[4]), .B(a[84]), .Z(n1996) );
  AND U4640 ( .A(b[3]), .B(a[86]), .Z(n1955) );
  AND U4641 ( .A(b[4]), .B(a[86]), .Z(n1934) );
  AND U4642 ( .A(b[4]), .B(a[87]), .Z(n1902) );
  AND U4643 ( .A(b[4]), .B(a[88]), .Z(n1870) );
  AND U4644 ( .A(b[4]), .B(a[89]), .Z(n1837) );
  AND U4645 ( .A(b[4]), .B(a[90]), .Z(n1805) );
  AND U4646 ( .A(b[4]), .B(a[91]), .Z(n1774) );
  AND U4647 ( .A(b[3]), .B(a[93]), .Z(n1733) );
  AND U4648 ( .A(b[3]), .B(a[94]), .Z(n1702) );
  AND U4649 ( .A(b[3]), .B(a[95]), .Z(n1670) );
  AND U4650 ( .A(b[3]), .B(a[96]), .Z(n1638) );
  AND U4651 ( .A(b[3]), .B(a[97]), .Z(n1604) );
  XNOR U4652 ( .A(n1570), .B(n1571), .Z(c[127]) );
  XOR U4653 ( .A(sreg[135]), .B(n1569), .Z(n1571) );
  XOR U4654 ( .A(n4467), .B(n4523), .Z(n1570) );
  XNOR U4655 ( .A(n4466), .B(n1569), .Z(n4523) );
  XOR U4656 ( .A(n4524), .B(n4525), .Z(n1569) );
  ANDN U4657 ( .B(n4526), .A(n4527), .Z(n4524) );
  NANDN U4658 ( .A(n187), .B(a[7]), .Z(n4466) );
  XNOR U4659 ( .A(n4492), .B(n4528), .Z(n4494) );
  NAND U4660 ( .A(b[1]), .B(a[6]), .Z(n4528) );
  XNOR U4661 ( .A(n4492), .B(n4505), .Z(n4529) );
  XOR U4662 ( .A(n4530), .B(n4503), .Z(n4505) );
  AND U4663 ( .A(a[5]), .B(b[2]), .Z(n4530) );
  OR U4664 ( .A(n4531), .B(n4532), .Z(n4492) );
  XOR U4665 ( .A(n4503), .B(n4521), .Z(n4533) );
  XOR U4666 ( .A(n4520), .B(n4517), .Z(n4534) );
  XOR U4667 ( .A(n4535), .B(n4536), .Z(n4517) );
  XOR U4668 ( .A(n4515), .B(n4537), .Z(n4536) );
  XOR U4669 ( .A(n4538), .B(n4539), .Z(n4537) );
  XOR U4670 ( .A(n4540), .B(n4541), .Z(n4539) );
  NAND U4671 ( .A(a[1]), .B(b[6]), .Z(n4541) );
  AND U4672 ( .A(a[0]), .B(b[7]), .Z(n4540) );
  XOR U4673 ( .A(n4542), .B(n4538), .Z(n4535) );
  XOR U4674 ( .A(n4543), .B(n4544), .Z(n4538) );
  NOR U4675 ( .A(n4545), .B(n4546), .Z(n4543) );
  AND U4676 ( .A(a[2]), .B(b[5]), .Z(n4542) );
  XNOR U4677 ( .A(n4547), .B(n4515), .Z(n4516) );
  XOR U4678 ( .A(n4548), .B(n4549), .Z(n4515) );
  ANDN U4679 ( .B(n4550), .A(n4551), .Z(n4548) );
  AND U4680 ( .A(a[3]), .B(b[4]), .Z(n4547) );
  XNOR U4681 ( .A(n4552), .B(n4553), .Z(n4503) );
  OR U4682 ( .A(n4554), .B(n4555), .Z(n4553) );
  XNOR U4683 ( .A(n4556), .B(n4520), .Z(n4522) );
  XNOR U4684 ( .A(n4557), .B(n4558), .Z(n4520) );
  NOR U4685 ( .A(n4559), .B(n4560), .Z(n4557) );
  AND U4686 ( .A(b[3]), .B(a[4]), .Z(n4556) );
  XNOR U4687 ( .A(n4526), .B(n4527), .Z(c[126]) );
  XOR U4688 ( .A(sreg[134]), .B(n4525), .Z(n4527) );
  XOR U4689 ( .A(n4532), .B(n4561), .Z(n4526) );
  XNOR U4690 ( .A(n4531), .B(n4525), .Z(n4561) );
  XOR U4691 ( .A(n4562), .B(n4563), .Z(n4525) );
  ANDN U4692 ( .B(n4564), .A(n4565), .Z(n4562) );
  NANDN U4693 ( .A(n187), .B(a[6]), .Z(n4531) );
  XNOR U4694 ( .A(n4552), .B(n4566), .Z(n4554) );
  NAND U4695 ( .A(a[5]), .B(b[1]), .Z(n4566) );
  XNOR U4696 ( .A(n4552), .B(n4560), .Z(n4567) );
  XOR U4697 ( .A(n4568), .B(n4558), .Z(n4560) );
  AND U4698 ( .A(b[2]), .B(a[4]), .Z(n4568) );
  OR U4699 ( .A(n4569), .B(n4570), .Z(n4552) );
  XOR U4700 ( .A(n4558), .B(n4550), .Z(n4571) );
  XOR U4701 ( .A(n4549), .B(n4546), .Z(n4572) );
  XOR U4702 ( .A(n4573), .B(n4574), .Z(n4546) );
  XOR U4703 ( .A(n4544), .B(n4575), .Z(n4574) );
  XOR U4704 ( .A(n4576), .B(n4577), .Z(n4575) );
  AND U4705 ( .A(a[0]), .B(b[6]), .Z(n4576) );
  XNOR U4706 ( .A(n4578), .B(n4577), .Z(n4573) );
  XOR U4707 ( .A(n4579), .B(n4580), .Z(n4577) );
  NOR U4708 ( .A(n4581), .B(n4582), .Z(n4579) );
  AND U4709 ( .A(a[1]), .B(b[5]), .Z(n4578) );
  XNOR U4710 ( .A(n4583), .B(n4544), .Z(n4545) );
  XOR U4711 ( .A(n4584), .B(n4585), .Z(n4544) );
  NOR U4712 ( .A(n4586), .B(n4587), .Z(n4584) );
  AND U4713 ( .A(a[2]), .B(b[4]), .Z(n4583) );
  XNOR U4714 ( .A(n4588), .B(n4589), .Z(n4558) );
  OR U4715 ( .A(n4590), .B(n4591), .Z(n4589) );
  XNOR U4716 ( .A(n4592), .B(n4549), .Z(n4551) );
  XNOR U4717 ( .A(n4593), .B(n4594), .Z(n4549) );
  NOR U4718 ( .A(n4595), .B(n4596), .Z(n4593) );
  AND U4719 ( .A(a[3]), .B(b[3]), .Z(n4592) );
  XNOR U4720 ( .A(n4564), .B(n4565), .Z(c[125]) );
  XOR U4721 ( .A(sreg[133]), .B(n4563), .Z(n4565) );
  XOR U4722 ( .A(n4570), .B(n4597), .Z(n4564) );
  XNOR U4723 ( .A(n4569), .B(n4563), .Z(n4597) );
  XOR U4724 ( .A(n4598), .B(n4599), .Z(n4563) );
  ANDN U4725 ( .B(n4600), .A(n4601), .Z(n4598) );
  NANDN U4726 ( .A(n187), .B(a[5]), .Z(n4569) );
  XNOR U4727 ( .A(n4588), .B(n4602), .Z(n4590) );
  NAND U4728 ( .A(b[1]), .B(a[4]), .Z(n4602) );
  XNOR U4729 ( .A(n4588), .B(n4596), .Z(n4603) );
  XOR U4730 ( .A(n4604), .B(n4594), .Z(n4596) );
  AND U4731 ( .A(b[2]), .B(a[3]), .Z(n4604) );
  OR U4732 ( .A(n4605), .B(n4606), .Z(n4588) );
  XNOR U4733 ( .A(n4594), .B(n4587), .Z(n4607) );
  XOR U4734 ( .A(n4581), .B(n4608), .Z(n4587) );
  XNOR U4735 ( .A(n4585), .B(n4582), .Z(n4608) );
  XNOR U4736 ( .A(n4609), .B(n4580), .Z(n4582) );
  AND U4737 ( .A(a[0]), .B(b[5]), .Z(n4609) );
  XNOR U4738 ( .A(n4610), .B(n4580), .Z(n4581) );
  XOR U4739 ( .A(n4611), .B(n4612), .Z(n4580) );
  NOR U4740 ( .A(n4613), .B(n4614), .Z(n4611) );
  AND U4741 ( .A(a[1]), .B(b[4]), .Z(n4610) );
  XNOR U4742 ( .A(n4615), .B(n4616), .Z(n4594) );
  OR U4743 ( .A(n4617), .B(n4618), .Z(n4616) );
  XNOR U4744 ( .A(n4619), .B(n4585), .Z(n4586) );
  XNOR U4745 ( .A(n4620), .B(n4621), .Z(n4585) );
  NOR U4746 ( .A(n4622), .B(n4623), .Z(n4620) );
  AND U4747 ( .A(a[2]), .B(b[3]), .Z(n4619) );
  XNOR U4748 ( .A(n4600), .B(n4601), .Z(c[124]) );
  XOR U4749 ( .A(sreg[132]), .B(n4599), .Z(n4601) );
  XOR U4750 ( .A(n4606), .B(n4624), .Z(n4600) );
  XNOR U4751 ( .A(n4605), .B(n4599), .Z(n4624) );
  XOR U4752 ( .A(n4625), .B(n4626), .Z(n4599) );
  ANDN U4753 ( .B(n4627), .A(n4628), .Z(n4625) );
  NANDN U4754 ( .A(n187), .B(a[4]), .Z(n4605) );
  XNOR U4755 ( .A(n4615), .B(n4629), .Z(n4617) );
  NAND U4756 ( .A(a[3]), .B(b[1]), .Z(n4629) );
  XNOR U4757 ( .A(n4615), .B(n4623), .Z(n4630) );
  XOR U4758 ( .A(n4631), .B(n4621), .Z(n4623) );
  AND U4759 ( .A(b[2]), .B(a[2]), .Z(n4631) );
  OR U4760 ( .A(n4632), .B(n4633), .Z(n4615) );
  XOR U4761 ( .A(n4613), .B(n4634), .Z(n4622) );
  XOR U4762 ( .A(n4621), .B(n4614), .Z(n4634) );
  XNOR U4763 ( .A(n4635), .B(n4612), .Z(n4614) );
  AND U4764 ( .A(a[0]), .B(b[4]), .Z(n4635) );
  XOR U4765 ( .A(n4636), .B(n4637), .Z(n4621) );
  OR U4766 ( .A(n4638), .B(n4639), .Z(n4637) );
  XNOR U4767 ( .A(n4640), .B(n4612), .Z(n4613) );
  XOR U4768 ( .A(n4641), .B(n4642), .Z(n4612) );
  NOR U4769 ( .A(n4643), .B(n4644), .Z(n4641) );
  AND U4770 ( .A(a[1]), .B(b[3]), .Z(n4640) );
  XNOR U4771 ( .A(n4627), .B(n4628), .Z(c[123]) );
  XOR U4772 ( .A(sreg[131]), .B(n4626), .Z(n4628) );
  XOR U4773 ( .A(n4633), .B(n4645), .Z(n4627) );
  XNOR U4774 ( .A(n4632), .B(n4626), .Z(n4645) );
  XNOR U4775 ( .A(n4646), .B(n4647), .Z(n4626) );
  ANDN U4776 ( .B(n4648), .A(n4649), .Z(n4646) );
  NANDN U4777 ( .A(n187), .B(a[3]), .Z(n4632) );
  XOR U4778 ( .A(n4636), .B(n4650), .Z(n4638) );
  NAND U4779 ( .A(b[1]), .B(a[2]), .Z(n4650) );
  XOR U4780 ( .A(n4643), .B(n4651), .Z(n4639) );
  XNOR U4781 ( .A(n4636), .B(n4644), .Z(n4651) );
  XNOR U4782 ( .A(n4652), .B(n4642), .Z(n4644) );
  AND U4783 ( .A(b[2]), .B(a[1]), .Z(n4652) );
  NOR U4784 ( .A(n4653), .B(n4654), .Z(n4636) );
  XNOR U4785 ( .A(n4655), .B(n4642), .Z(n4643) );
  NAND U4786 ( .A(n4656), .B(n4657), .Z(n4642) );
  OR U4787 ( .A(n4658), .B(n4659), .Z(n4657) );
  AND U4788 ( .A(a[0]), .B(b[3]), .Z(n4655) );
  XNOR U4789 ( .A(n4648), .B(n4649), .Z(c[122]) );
  XNOR U4790 ( .A(sreg[130]), .B(n4647), .Z(n4649) );
  XNOR U4791 ( .A(n4654), .B(n4661), .Z(n4660) );
  IV U4792 ( .A(n4647), .Z(n4661) );
  XNOR U4793 ( .A(n4662), .B(n4663), .Z(n4647) );
  NAND U4794 ( .A(n4664), .B(n4665), .Z(n4663) );
  NANDN U4795 ( .A(n187), .B(a[2]), .Z(n4654) );
  XOR U4796 ( .A(n4666), .B(n4656), .Z(n4659) );
  AND U4797 ( .A(b[2]), .B(a[0]), .Z(n4666) );
  NAND U4798 ( .A(n4667), .B(b[1]), .Z(n4658) );
  NANDN U4799 ( .A(n4668), .B(n4669), .Z(n4656) );
  XOR U4800 ( .A(n4664), .B(n4665), .Z(c[121]) );
  XOR U4801 ( .A(sreg[129]), .B(n4662), .Z(n4665) );
  XNOR U4802 ( .A(n4662), .B(n4670), .Z(n4664) );
  XOR U4803 ( .A(n4668), .B(n4669), .Z(n4670) );
  AND U4804 ( .A(a[1]), .B(b[0]), .Z(n4669) );
  NAND U4805 ( .A(b[1]), .B(a[0]), .Z(n4668) );
  ANDN U4806 ( .B(sreg[128]), .A(n4671), .Z(n4662) );
  XNOR U4807 ( .A(sreg[128]), .B(n4671), .Z(c[120]) );
  NANDN U4808 ( .A(n187), .B(a[0]), .Z(n4671) );
  IV U4809 ( .A(b[0]), .Z(n187) );
endmodule

