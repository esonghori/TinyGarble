
module sum_N1024_CC16 ( clk, rst, a, b, c );
  input [63:0] a;
  input [63:0] b;
  output [63:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .Q(carry_on) );
  XOR U3 ( .A(a[0]), .B(b[0]), .Z(n1) );
  XOR U4 ( .A(n1), .B(carry_on), .Z(c[0]) );
  XOR U5 ( .A(a[1]), .B(b[1]), .Z(n4) );
  NAND U6 ( .A(b[0]), .B(a[0]), .Z(n3) );
  NAND U7 ( .A(carry_on), .B(n1), .Z(n2) );
  AND U8 ( .A(n3), .B(n2), .Z(n5) );
  XNOR U9 ( .A(n4), .B(n5), .Z(c[1]) );
  XOR U10 ( .A(a[2]), .B(b[2]), .Z(n8) );
  NAND U11 ( .A(b[1]), .B(a[1]), .Z(n7) );
  NANDN U12 ( .A(n5), .B(n4), .Z(n6) );
  AND U13 ( .A(n7), .B(n6), .Z(n9) );
  XNOR U14 ( .A(n8), .B(n9), .Z(c[2]) );
  XOR U15 ( .A(a[3]), .B(b[3]), .Z(n12) );
  NAND U16 ( .A(b[2]), .B(a[2]), .Z(n11) );
  NANDN U17 ( .A(n9), .B(n8), .Z(n10) );
  AND U18 ( .A(n11), .B(n10), .Z(n13) );
  XNOR U19 ( .A(n12), .B(n13), .Z(c[3]) );
  XOR U20 ( .A(a[4]), .B(b[4]), .Z(n16) );
  NAND U21 ( .A(b[3]), .B(a[3]), .Z(n15) );
  NANDN U22 ( .A(n13), .B(n12), .Z(n14) );
  AND U23 ( .A(n15), .B(n14), .Z(n17) );
  XNOR U24 ( .A(n16), .B(n17), .Z(c[4]) );
  XOR U25 ( .A(a[5]), .B(b[5]), .Z(n20) );
  NAND U26 ( .A(b[4]), .B(a[4]), .Z(n19) );
  NANDN U27 ( .A(n17), .B(n16), .Z(n18) );
  AND U28 ( .A(n19), .B(n18), .Z(n21) );
  XNOR U29 ( .A(n20), .B(n21), .Z(c[5]) );
  XOR U30 ( .A(a[6]), .B(b[6]), .Z(n24) );
  NAND U31 ( .A(b[5]), .B(a[5]), .Z(n23) );
  NANDN U32 ( .A(n21), .B(n20), .Z(n22) );
  AND U33 ( .A(n23), .B(n22), .Z(n25) );
  XNOR U34 ( .A(n24), .B(n25), .Z(c[6]) );
  XOR U35 ( .A(a[7]), .B(b[7]), .Z(n28) );
  NAND U36 ( .A(b[6]), .B(a[6]), .Z(n27) );
  NANDN U37 ( .A(n25), .B(n24), .Z(n26) );
  AND U38 ( .A(n27), .B(n26), .Z(n29) );
  XNOR U39 ( .A(n28), .B(n29), .Z(c[7]) );
  XOR U40 ( .A(a[8]), .B(b[8]), .Z(n32) );
  NAND U41 ( .A(b[7]), .B(a[7]), .Z(n31) );
  NANDN U42 ( .A(n29), .B(n28), .Z(n30) );
  AND U43 ( .A(n31), .B(n30), .Z(n33) );
  XNOR U44 ( .A(n32), .B(n33), .Z(c[8]) );
  XOR U45 ( .A(a[9]), .B(b[9]), .Z(n36) );
  NAND U46 ( .A(b[8]), .B(a[8]), .Z(n35) );
  NANDN U47 ( .A(n33), .B(n32), .Z(n34) );
  AND U48 ( .A(n35), .B(n34), .Z(n37) );
  XNOR U49 ( .A(n36), .B(n37), .Z(c[9]) );
  XOR U50 ( .A(a[10]), .B(b[10]), .Z(n40) );
  NAND U51 ( .A(b[9]), .B(a[9]), .Z(n39) );
  NANDN U52 ( .A(n37), .B(n36), .Z(n38) );
  AND U53 ( .A(n39), .B(n38), .Z(n41) );
  XNOR U54 ( .A(n40), .B(n41), .Z(c[10]) );
  XOR U55 ( .A(a[11]), .B(b[11]), .Z(n44) );
  NAND U56 ( .A(b[10]), .B(a[10]), .Z(n43) );
  NANDN U57 ( .A(n41), .B(n40), .Z(n42) );
  AND U58 ( .A(n43), .B(n42), .Z(n45) );
  XNOR U59 ( .A(n44), .B(n45), .Z(c[11]) );
  XOR U60 ( .A(a[12]), .B(b[12]), .Z(n48) );
  NAND U61 ( .A(b[11]), .B(a[11]), .Z(n47) );
  NANDN U62 ( .A(n45), .B(n44), .Z(n46) );
  AND U63 ( .A(n47), .B(n46), .Z(n49) );
  XNOR U64 ( .A(n48), .B(n49), .Z(c[12]) );
  XOR U65 ( .A(a[13]), .B(b[13]), .Z(n52) );
  NAND U66 ( .A(b[12]), .B(a[12]), .Z(n51) );
  NANDN U67 ( .A(n49), .B(n48), .Z(n50) );
  AND U68 ( .A(n51), .B(n50), .Z(n53) );
  XNOR U69 ( .A(n52), .B(n53), .Z(c[13]) );
  XOR U70 ( .A(a[14]), .B(b[14]), .Z(n56) );
  NAND U71 ( .A(b[13]), .B(a[13]), .Z(n55) );
  NANDN U72 ( .A(n53), .B(n52), .Z(n54) );
  AND U73 ( .A(n55), .B(n54), .Z(n57) );
  XNOR U74 ( .A(n56), .B(n57), .Z(c[14]) );
  XOR U75 ( .A(a[15]), .B(b[15]), .Z(n60) );
  NAND U76 ( .A(b[14]), .B(a[14]), .Z(n59) );
  NANDN U77 ( .A(n57), .B(n56), .Z(n58) );
  AND U78 ( .A(n59), .B(n58), .Z(n61) );
  XNOR U79 ( .A(n60), .B(n61), .Z(c[15]) );
  XOR U80 ( .A(a[16]), .B(b[16]), .Z(n64) );
  NAND U81 ( .A(b[15]), .B(a[15]), .Z(n63) );
  NANDN U82 ( .A(n61), .B(n60), .Z(n62) );
  AND U83 ( .A(n63), .B(n62), .Z(n65) );
  XNOR U84 ( .A(n64), .B(n65), .Z(c[16]) );
  XOR U85 ( .A(a[17]), .B(b[17]), .Z(n68) );
  NAND U86 ( .A(b[16]), .B(a[16]), .Z(n67) );
  NANDN U87 ( .A(n65), .B(n64), .Z(n66) );
  AND U88 ( .A(n67), .B(n66), .Z(n69) );
  XNOR U89 ( .A(n68), .B(n69), .Z(c[17]) );
  XOR U90 ( .A(a[18]), .B(b[18]), .Z(n72) );
  NAND U91 ( .A(b[17]), .B(a[17]), .Z(n71) );
  NANDN U92 ( .A(n69), .B(n68), .Z(n70) );
  AND U93 ( .A(n71), .B(n70), .Z(n73) );
  XNOR U94 ( .A(n72), .B(n73), .Z(c[18]) );
  XOR U95 ( .A(a[19]), .B(b[19]), .Z(n76) );
  NAND U96 ( .A(b[18]), .B(a[18]), .Z(n75) );
  NANDN U97 ( .A(n73), .B(n72), .Z(n74) );
  AND U98 ( .A(n75), .B(n74), .Z(n77) );
  XNOR U99 ( .A(n76), .B(n77), .Z(c[19]) );
  XOR U100 ( .A(a[20]), .B(b[20]), .Z(n80) );
  NAND U101 ( .A(b[19]), .B(a[19]), .Z(n79) );
  NANDN U102 ( .A(n77), .B(n76), .Z(n78) );
  AND U103 ( .A(n79), .B(n78), .Z(n81) );
  XNOR U104 ( .A(n80), .B(n81), .Z(c[20]) );
  XOR U105 ( .A(a[21]), .B(b[21]), .Z(n84) );
  NAND U106 ( .A(b[20]), .B(a[20]), .Z(n83) );
  NANDN U107 ( .A(n81), .B(n80), .Z(n82) );
  AND U108 ( .A(n83), .B(n82), .Z(n85) );
  XNOR U109 ( .A(n84), .B(n85), .Z(c[21]) );
  XOR U110 ( .A(a[22]), .B(b[22]), .Z(n88) );
  NAND U111 ( .A(b[21]), .B(a[21]), .Z(n87) );
  NANDN U112 ( .A(n85), .B(n84), .Z(n86) );
  AND U113 ( .A(n87), .B(n86), .Z(n89) );
  XNOR U114 ( .A(n88), .B(n89), .Z(c[22]) );
  XOR U115 ( .A(a[23]), .B(b[23]), .Z(n92) );
  NAND U116 ( .A(b[22]), .B(a[22]), .Z(n91) );
  NANDN U117 ( .A(n89), .B(n88), .Z(n90) );
  AND U118 ( .A(n91), .B(n90), .Z(n93) );
  XNOR U119 ( .A(n92), .B(n93), .Z(c[23]) );
  XOR U120 ( .A(a[24]), .B(b[24]), .Z(n96) );
  NAND U121 ( .A(b[23]), .B(a[23]), .Z(n95) );
  NANDN U122 ( .A(n93), .B(n92), .Z(n94) );
  AND U123 ( .A(n95), .B(n94), .Z(n97) );
  XNOR U124 ( .A(n96), .B(n97), .Z(c[24]) );
  XOR U125 ( .A(a[25]), .B(b[25]), .Z(n100) );
  NAND U126 ( .A(b[24]), .B(a[24]), .Z(n99) );
  NANDN U127 ( .A(n97), .B(n96), .Z(n98) );
  AND U128 ( .A(n99), .B(n98), .Z(n101) );
  XNOR U129 ( .A(n100), .B(n101), .Z(c[25]) );
  XOR U130 ( .A(a[26]), .B(b[26]), .Z(n104) );
  NAND U131 ( .A(b[25]), .B(a[25]), .Z(n103) );
  NANDN U132 ( .A(n101), .B(n100), .Z(n102) );
  AND U133 ( .A(n103), .B(n102), .Z(n105) );
  XNOR U134 ( .A(n104), .B(n105), .Z(c[26]) );
  XOR U135 ( .A(a[27]), .B(b[27]), .Z(n108) );
  NAND U136 ( .A(b[26]), .B(a[26]), .Z(n107) );
  NANDN U137 ( .A(n105), .B(n104), .Z(n106) );
  AND U138 ( .A(n107), .B(n106), .Z(n109) );
  XNOR U139 ( .A(n108), .B(n109), .Z(c[27]) );
  XOR U140 ( .A(a[28]), .B(b[28]), .Z(n112) );
  NAND U141 ( .A(b[27]), .B(a[27]), .Z(n111) );
  NANDN U142 ( .A(n109), .B(n108), .Z(n110) );
  AND U143 ( .A(n111), .B(n110), .Z(n113) );
  XNOR U144 ( .A(n112), .B(n113), .Z(c[28]) );
  XOR U145 ( .A(a[29]), .B(b[29]), .Z(n116) );
  NAND U146 ( .A(b[28]), .B(a[28]), .Z(n115) );
  NANDN U147 ( .A(n113), .B(n112), .Z(n114) );
  AND U148 ( .A(n115), .B(n114), .Z(n117) );
  XNOR U149 ( .A(n116), .B(n117), .Z(c[29]) );
  XOR U150 ( .A(a[30]), .B(b[30]), .Z(n120) );
  NAND U151 ( .A(b[29]), .B(a[29]), .Z(n119) );
  NANDN U152 ( .A(n117), .B(n116), .Z(n118) );
  AND U153 ( .A(n119), .B(n118), .Z(n121) );
  XNOR U154 ( .A(n120), .B(n121), .Z(c[30]) );
  XOR U155 ( .A(a[31]), .B(b[31]), .Z(n124) );
  NAND U156 ( .A(b[30]), .B(a[30]), .Z(n123) );
  NANDN U157 ( .A(n121), .B(n120), .Z(n122) );
  AND U158 ( .A(n123), .B(n122), .Z(n125) );
  XNOR U159 ( .A(n124), .B(n125), .Z(c[31]) );
  XOR U160 ( .A(a[32]), .B(b[32]), .Z(n128) );
  NAND U161 ( .A(b[31]), .B(a[31]), .Z(n127) );
  NANDN U162 ( .A(n125), .B(n124), .Z(n126) );
  AND U163 ( .A(n127), .B(n126), .Z(n129) );
  XNOR U164 ( .A(n128), .B(n129), .Z(c[32]) );
  XOR U165 ( .A(a[33]), .B(b[33]), .Z(n132) );
  NAND U166 ( .A(b[32]), .B(a[32]), .Z(n131) );
  NANDN U167 ( .A(n129), .B(n128), .Z(n130) );
  AND U168 ( .A(n131), .B(n130), .Z(n133) );
  XNOR U169 ( .A(n132), .B(n133), .Z(c[33]) );
  XOR U170 ( .A(a[34]), .B(b[34]), .Z(n136) );
  NAND U171 ( .A(b[33]), .B(a[33]), .Z(n135) );
  NANDN U172 ( .A(n133), .B(n132), .Z(n134) );
  AND U173 ( .A(n135), .B(n134), .Z(n137) );
  XNOR U174 ( .A(n136), .B(n137), .Z(c[34]) );
  XOR U175 ( .A(a[35]), .B(b[35]), .Z(n140) );
  NAND U176 ( .A(b[34]), .B(a[34]), .Z(n139) );
  NANDN U177 ( .A(n137), .B(n136), .Z(n138) );
  AND U178 ( .A(n139), .B(n138), .Z(n141) );
  XNOR U179 ( .A(n140), .B(n141), .Z(c[35]) );
  XOR U180 ( .A(a[36]), .B(b[36]), .Z(n144) );
  NAND U181 ( .A(b[35]), .B(a[35]), .Z(n143) );
  NANDN U182 ( .A(n141), .B(n140), .Z(n142) );
  AND U183 ( .A(n143), .B(n142), .Z(n145) );
  XNOR U184 ( .A(n144), .B(n145), .Z(c[36]) );
  XOR U185 ( .A(a[37]), .B(b[37]), .Z(n148) );
  NAND U186 ( .A(b[36]), .B(a[36]), .Z(n147) );
  NANDN U187 ( .A(n145), .B(n144), .Z(n146) );
  AND U188 ( .A(n147), .B(n146), .Z(n149) );
  XNOR U189 ( .A(n148), .B(n149), .Z(c[37]) );
  XOR U190 ( .A(a[38]), .B(b[38]), .Z(n152) );
  NAND U191 ( .A(b[37]), .B(a[37]), .Z(n151) );
  NANDN U192 ( .A(n149), .B(n148), .Z(n150) );
  AND U193 ( .A(n151), .B(n150), .Z(n153) );
  XNOR U194 ( .A(n152), .B(n153), .Z(c[38]) );
  XOR U195 ( .A(a[39]), .B(b[39]), .Z(n156) );
  NAND U196 ( .A(b[38]), .B(a[38]), .Z(n155) );
  NANDN U197 ( .A(n153), .B(n152), .Z(n154) );
  AND U198 ( .A(n155), .B(n154), .Z(n157) );
  XNOR U199 ( .A(n156), .B(n157), .Z(c[39]) );
  XOR U200 ( .A(a[40]), .B(b[40]), .Z(n160) );
  NAND U201 ( .A(b[39]), .B(a[39]), .Z(n159) );
  NANDN U202 ( .A(n157), .B(n156), .Z(n158) );
  AND U203 ( .A(n159), .B(n158), .Z(n161) );
  XNOR U204 ( .A(n160), .B(n161), .Z(c[40]) );
  XOR U205 ( .A(a[41]), .B(b[41]), .Z(n164) );
  NAND U206 ( .A(b[40]), .B(a[40]), .Z(n163) );
  NANDN U207 ( .A(n161), .B(n160), .Z(n162) );
  AND U208 ( .A(n163), .B(n162), .Z(n165) );
  XNOR U209 ( .A(n164), .B(n165), .Z(c[41]) );
  XOR U210 ( .A(a[42]), .B(b[42]), .Z(n168) );
  NAND U211 ( .A(b[41]), .B(a[41]), .Z(n167) );
  NANDN U212 ( .A(n165), .B(n164), .Z(n166) );
  AND U213 ( .A(n167), .B(n166), .Z(n169) );
  XNOR U214 ( .A(n168), .B(n169), .Z(c[42]) );
  XOR U215 ( .A(a[43]), .B(b[43]), .Z(n172) );
  NAND U216 ( .A(b[42]), .B(a[42]), .Z(n171) );
  NANDN U217 ( .A(n169), .B(n168), .Z(n170) );
  AND U218 ( .A(n171), .B(n170), .Z(n173) );
  XNOR U219 ( .A(n172), .B(n173), .Z(c[43]) );
  XOR U220 ( .A(a[44]), .B(b[44]), .Z(n176) );
  NAND U221 ( .A(b[43]), .B(a[43]), .Z(n175) );
  NANDN U222 ( .A(n173), .B(n172), .Z(n174) );
  AND U223 ( .A(n175), .B(n174), .Z(n177) );
  XNOR U224 ( .A(n176), .B(n177), .Z(c[44]) );
  XOR U225 ( .A(a[45]), .B(b[45]), .Z(n180) );
  NAND U226 ( .A(b[44]), .B(a[44]), .Z(n179) );
  NANDN U227 ( .A(n177), .B(n176), .Z(n178) );
  AND U228 ( .A(n179), .B(n178), .Z(n181) );
  XNOR U229 ( .A(n180), .B(n181), .Z(c[45]) );
  XOR U230 ( .A(a[46]), .B(b[46]), .Z(n184) );
  NAND U231 ( .A(b[45]), .B(a[45]), .Z(n183) );
  NANDN U232 ( .A(n181), .B(n180), .Z(n182) );
  AND U233 ( .A(n183), .B(n182), .Z(n185) );
  XNOR U234 ( .A(n184), .B(n185), .Z(c[46]) );
  XOR U235 ( .A(a[47]), .B(b[47]), .Z(n188) );
  NAND U236 ( .A(b[46]), .B(a[46]), .Z(n187) );
  NANDN U237 ( .A(n185), .B(n184), .Z(n186) );
  AND U238 ( .A(n187), .B(n186), .Z(n189) );
  XNOR U239 ( .A(n188), .B(n189), .Z(c[47]) );
  XOR U240 ( .A(a[48]), .B(b[48]), .Z(n192) );
  NAND U241 ( .A(b[47]), .B(a[47]), .Z(n191) );
  NANDN U242 ( .A(n189), .B(n188), .Z(n190) );
  AND U243 ( .A(n191), .B(n190), .Z(n193) );
  XNOR U244 ( .A(n192), .B(n193), .Z(c[48]) );
  XOR U245 ( .A(a[49]), .B(b[49]), .Z(n196) );
  NAND U246 ( .A(b[48]), .B(a[48]), .Z(n195) );
  NANDN U247 ( .A(n193), .B(n192), .Z(n194) );
  AND U248 ( .A(n195), .B(n194), .Z(n197) );
  XNOR U249 ( .A(n196), .B(n197), .Z(c[49]) );
  XOR U250 ( .A(a[50]), .B(b[50]), .Z(n200) );
  NAND U251 ( .A(b[49]), .B(a[49]), .Z(n199) );
  NANDN U252 ( .A(n197), .B(n196), .Z(n198) );
  AND U253 ( .A(n199), .B(n198), .Z(n201) );
  XNOR U254 ( .A(n200), .B(n201), .Z(c[50]) );
  XOR U255 ( .A(a[51]), .B(b[51]), .Z(n204) );
  NAND U256 ( .A(b[50]), .B(a[50]), .Z(n203) );
  NANDN U257 ( .A(n201), .B(n200), .Z(n202) );
  AND U258 ( .A(n203), .B(n202), .Z(n205) );
  XNOR U259 ( .A(n204), .B(n205), .Z(c[51]) );
  XOR U260 ( .A(a[52]), .B(b[52]), .Z(n208) );
  NAND U261 ( .A(b[51]), .B(a[51]), .Z(n207) );
  NANDN U262 ( .A(n205), .B(n204), .Z(n206) );
  AND U263 ( .A(n207), .B(n206), .Z(n209) );
  XNOR U264 ( .A(n208), .B(n209), .Z(c[52]) );
  XOR U265 ( .A(a[53]), .B(b[53]), .Z(n212) );
  NAND U266 ( .A(b[52]), .B(a[52]), .Z(n211) );
  NANDN U267 ( .A(n209), .B(n208), .Z(n210) );
  AND U268 ( .A(n211), .B(n210), .Z(n213) );
  XNOR U269 ( .A(n212), .B(n213), .Z(c[53]) );
  XOR U270 ( .A(a[54]), .B(b[54]), .Z(n216) );
  NAND U271 ( .A(b[53]), .B(a[53]), .Z(n215) );
  NANDN U272 ( .A(n213), .B(n212), .Z(n214) );
  AND U273 ( .A(n215), .B(n214), .Z(n217) );
  XNOR U274 ( .A(n216), .B(n217), .Z(c[54]) );
  XOR U275 ( .A(a[55]), .B(b[55]), .Z(n220) );
  NAND U276 ( .A(b[54]), .B(a[54]), .Z(n219) );
  NANDN U277 ( .A(n217), .B(n216), .Z(n218) );
  AND U278 ( .A(n219), .B(n218), .Z(n221) );
  XNOR U279 ( .A(n220), .B(n221), .Z(c[55]) );
  XOR U280 ( .A(a[56]), .B(b[56]), .Z(n224) );
  NAND U281 ( .A(b[55]), .B(a[55]), .Z(n223) );
  NANDN U282 ( .A(n221), .B(n220), .Z(n222) );
  AND U283 ( .A(n223), .B(n222), .Z(n225) );
  XNOR U284 ( .A(n224), .B(n225), .Z(c[56]) );
  XOR U285 ( .A(a[57]), .B(b[57]), .Z(n228) );
  NAND U286 ( .A(b[56]), .B(a[56]), .Z(n227) );
  NANDN U287 ( .A(n225), .B(n224), .Z(n226) );
  AND U288 ( .A(n227), .B(n226), .Z(n229) );
  XNOR U289 ( .A(n228), .B(n229), .Z(c[57]) );
  XOR U290 ( .A(a[58]), .B(b[58]), .Z(n232) );
  NAND U291 ( .A(b[57]), .B(a[57]), .Z(n231) );
  NANDN U292 ( .A(n229), .B(n228), .Z(n230) );
  AND U293 ( .A(n231), .B(n230), .Z(n233) );
  XNOR U294 ( .A(n232), .B(n233), .Z(c[58]) );
  XOR U295 ( .A(a[59]), .B(b[59]), .Z(n236) );
  NAND U296 ( .A(b[58]), .B(a[58]), .Z(n235) );
  NANDN U297 ( .A(n233), .B(n232), .Z(n234) );
  AND U298 ( .A(n235), .B(n234), .Z(n237) );
  XNOR U299 ( .A(n236), .B(n237), .Z(c[59]) );
  XOR U300 ( .A(a[60]), .B(b[60]), .Z(n240) );
  NAND U301 ( .A(b[59]), .B(a[59]), .Z(n239) );
  NANDN U302 ( .A(n237), .B(n236), .Z(n238) );
  AND U303 ( .A(n239), .B(n238), .Z(n241) );
  XNOR U304 ( .A(n240), .B(n241), .Z(c[60]) );
  XOR U305 ( .A(a[61]), .B(b[61]), .Z(n244) );
  NAND U306 ( .A(b[60]), .B(a[60]), .Z(n243) );
  NANDN U307 ( .A(n241), .B(n240), .Z(n242) );
  AND U308 ( .A(n243), .B(n242), .Z(n245) );
  XNOR U309 ( .A(n244), .B(n245), .Z(c[61]) );
  XOR U310 ( .A(a[62]), .B(b[62]), .Z(n248) );
  NAND U311 ( .A(b[61]), .B(a[61]), .Z(n247) );
  NANDN U312 ( .A(n245), .B(n244), .Z(n246) );
  AND U313 ( .A(n247), .B(n246), .Z(n249) );
  XNOR U314 ( .A(n248), .B(n249), .Z(c[62]) );
  NAND U315 ( .A(b[62]), .B(a[62]), .Z(n251) );
  NANDN U316 ( .A(n249), .B(n248), .Z(n250) );
  NAND U317 ( .A(n251), .B(n250), .Z(n252) );
  XOR U318 ( .A(a[63]), .B(b[63]), .Z(n253) );
  XOR U319 ( .A(n252), .B(n253), .Z(c[63]) );
  NAND U320 ( .A(b[63]), .B(a[63]), .Z(n255) );
  NAND U321 ( .A(n253), .B(n252), .Z(n254) );
  NAND U322 ( .A(n255), .B(n254), .Z(carry_on_d) );
endmodule

