
module first_nns_comb_W7_N128 ( q, DB, min_val_out );
  input [6:0] q;
  input [895:0] DB;
  output [6:0] min_val_out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037;

  XOR U897 ( .A(DB[895]), .B(n1), .Z(min_val_out[6]) );
  AND U898 ( .A(n2), .B(n3), .Z(n1) );
  XOR U899 ( .A(n4), .B(n5), .Z(n3) );
  XOR U900 ( .A(DB[895]), .B(DB[888]), .Z(n5) );
  AND U901 ( .A(n6), .B(n7), .Z(n4) );
  XOR U902 ( .A(n8), .B(n9), .Z(n7) );
  XOR U903 ( .A(DB[888]), .B(DB[881]), .Z(n9) );
  AND U904 ( .A(n10), .B(n11), .Z(n8) );
  XOR U905 ( .A(n12), .B(n13), .Z(n11) );
  XOR U906 ( .A(DB[881]), .B(DB[874]), .Z(n13) );
  AND U907 ( .A(n14), .B(n15), .Z(n12) );
  XOR U908 ( .A(n16), .B(n17), .Z(n15) );
  XOR U909 ( .A(DB[874]), .B(DB[867]), .Z(n17) );
  AND U910 ( .A(n18), .B(n19), .Z(n16) );
  XOR U911 ( .A(n20), .B(n21), .Z(n19) );
  XOR U912 ( .A(DB[867]), .B(DB[860]), .Z(n21) );
  AND U913 ( .A(n22), .B(n23), .Z(n20) );
  XOR U914 ( .A(n24), .B(n25), .Z(n23) );
  XOR U915 ( .A(DB[860]), .B(DB[853]), .Z(n25) );
  AND U916 ( .A(n26), .B(n27), .Z(n24) );
  XOR U917 ( .A(n28), .B(n29), .Z(n27) );
  XOR U918 ( .A(DB[853]), .B(DB[846]), .Z(n29) );
  AND U919 ( .A(n30), .B(n31), .Z(n28) );
  XOR U920 ( .A(n32), .B(n33), .Z(n31) );
  XOR U921 ( .A(DB[846]), .B(DB[839]), .Z(n33) );
  AND U922 ( .A(n34), .B(n35), .Z(n32) );
  XOR U923 ( .A(n36), .B(n37), .Z(n35) );
  XOR U924 ( .A(DB[839]), .B(DB[832]), .Z(n37) );
  AND U925 ( .A(n38), .B(n39), .Z(n36) );
  XOR U926 ( .A(n40), .B(n41), .Z(n39) );
  XOR U927 ( .A(DB[832]), .B(DB[825]), .Z(n41) );
  AND U928 ( .A(n42), .B(n43), .Z(n40) );
  XOR U929 ( .A(n44), .B(n45), .Z(n43) );
  XOR U930 ( .A(DB[825]), .B(DB[818]), .Z(n45) );
  AND U931 ( .A(n46), .B(n47), .Z(n44) );
  XOR U932 ( .A(n48), .B(n49), .Z(n47) );
  XOR U933 ( .A(DB[818]), .B(DB[811]), .Z(n49) );
  AND U934 ( .A(n50), .B(n51), .Z(n48) );
  XOR U935 ( .A(n52), .B(n53), .Z(n51) );
  XOR U936 ( .A(DB[811]), .B(DB[804]), .Z(n53) );
  AND U937 ( .A(n54), .B(n55), .Z(n52) );
  XOR U938 ( .A(n56), .B(n57), .Z(n55) );
  XOR U939 ( .A(DB[804]), .B(DB[797]), .Z(n57) );
  AND U940 ( .A(n58), .B(n59), .Z(n56) );
  XOR U941 ( .A(n60), .B(n61), .Z(n59) );
  XOR U942 ( .A(DB[797]), .B(DB[790]), .Z(n61) );
  AND U943 ( .A(n62), .B(n63), .Z(n60) );
  XOR U944 ( .A(n64), .B(n65), .Z(n63) );
  XOR U945 ( .A(DB[790]), .B(DB[783]), .Z(n65) );
  AND U946 ( .A(n66), .B(n67), .Z(n64) );
  XOR U947 ( .A(n68), .B(n69), .Z(n67) );
  XOR U948 ( .A(DB[783]), .B(DB[776]), .Z(n69) );
  AND U949 ( .A(n70), .B(n71), .Z(n68) );
  XOR U950 ( .A(n72), .B(n73), .Z(n71) );
  XOR U951 ( .A(DB[776]), .B(DB[769]), .Z(n73) );
  AND U952 ( .A(n74), .B(n75), .Z(n72) );
  XOR U953 ( .A(n76), .B(n77), .Z(n75) );
  XOR U954 ( .A(DB[769]), .B(DB[762]), .Z(n77) );
  AND U955 ( .A(n78), .B(n79), .Z(n76) );
  XOR U956 ( .A(n80), .B(n81), .Z(n79) );
  XOR U957 ( .A(DB[762]), .B(DB[755]), .Z(n81) );
  AND U958 ( .A(n82), .B(n83), .Z(n80) );
  XOR U959 ( .A(n84), .B(n85), .Z(n83) );
  XOR U960 ( .A(DB[755]), .B(DB[748]), .Z(n85) );
  AND U961 ( .A(n86), .B(n87), .Z(n84) );
  XOR U962 ( .A(n88), .B(n89), .Z(n87) );
  XOR U963 ( .A(DB[748]), .B(DB[741]), .Z(n89) );
  AND U964 ( .A(n90), .B(n91), .Z(n88) );
  XOR U965 ( .A(n92), .B(n93), .Z(n91) );
  XOR U966 ( .A(DB[741]), .B(DB[734]), .Z(n93) );
  AND U967 ( .A(n94), .B(n95), .Z(n92) );
  XOR U968 ( .A(n96), .B(n97), .Z(n95) );
  XOR U969 ( .A(DB[734]), .B(DB[727]), .Z(n97) );
  AND U970 ( .A(n98), .B(n99), .Z(n96) );
  XOR U971 ( .A(n100), .B(n101), .Z(n99) );
  XOR U972 ( .A(DB[727]), .B(DB[720]), .Z(n101) );
  AND U973 ( .A(n102), .B(n103), .Z(n100) );
  XOR U974 ( .A(n104), .B(n105), .Z(n103) );
  XOR U975 ( .A(DB[720]), .B(DB[713]), .Z(n105) );
  AND U976 ( .A(n106), .B(n107), .Z(n104) );
  XOR U977 ( .A(n108), .B(n109), .Z(n107) );
  XOR U978 ( .A(DB[713]), .B(DB[706]), .Z(n109) );
  AND U979 ( .A(n110), .B(n111), .Z(n108) );
  XOR U980 ( .A(n112), .B(n113), .Z(n111) );
  XOR U981 ( .A(DB[706]), .B(DB[699]), .Z(n113) );
  AND U982 ( .A(n114), .B(n115), .Z(n112) );
  XOR U983 ( .A(n116), .B(n117), .Z(n115) );
  XOR U984 ( .A(DB[699]), .B(DB[692]), .Z(n117) );
  AND U985 ( .A(n118), .B(n119), .Z(n116) );
  XOR U986 ( .A(n120), .B(n121), .Z(n119) );
  XOR U987 ( .A(DB[692]), .B(DB[685]), .Z(n121) );
  AND U988 ( .A(n122), .B(n123), .Z(n120) );
  XOR U989 ( .A(n124), .B(n125), .Z(n123) );
  XOR U990 ( .A(DB[685]), .B(DB[678]), .Z(n125) );
  AND U991 ( .A(n126), .B(n127), .Z(n124) );
  XOR U992 ( .A(n128), .B(n129), .Z(n127) );
  XOR U993 ( .A(DB[678]), .B(DB[671]), .Z(n129) );
  AND U994 ( .A(n130), .B(n131), .Z(n128) );
  XOR U995 ( .A(n132), .B(n133), .Z(n131) );
  XOR U996 ( .A(DB[671]), .B(DB[664]), .Z(n133) );
  AND U997 ( .A(n134), .B(n135), .Z(n132) );
  XOR U998 ( .A(n136), .B(n137), .Z(n135) );
  XOR U999 ( .A(DB[664]), .B(DB[657]), .Z(n137) );
  AND U1000 ( .A(n138), .B(n139), .Z(n136) );
  XOR U1001 ( .A(n140), .B(n141), .Z(n139) );
  XOR U1002 ( .A(DB[657]), .B(DB[650]), .Z(n141) );
  AND U1003 ( .A(n142), .B(n143), .Z(n140) );
  XOR U1004 ( .A(n144), .B(n145), .Z(n143) );
  XOR U1005 ( .A(DB[650]), .B(DB[643]), .Z(n145) );
  AND U1006 ( .A(n146), .B(n147), .Z(n144) );
  XOR U1007 ( .A(n148), .B(n149), .Z(n147) );
  XOR U1008 ( .A(DB[643]), .B(DB[636]), .Z(n149) );
  AND U1009 ( .A(n150), .B(n151), .Z(n148) );
  XOR U1010 ( .A(n152), .B(n153), .Z(n151) );
  XOR U1011 ( .A(DB[636]), .B(DB[629]), .Z(n153) );
  AND U1012 ( .A(n154), .B(n155), .Z(n152) );
  XOR U1013 ( .A(n156), .B(n157), .Z(n155) );
  XOR U1014 ( .A(DB[629]), .B(DB[622]), .Z(n157) );
  AND U1015 ( .A(n158), .B(n159), .Z(n156) );
  XOR U1016 ( .A(n160), .B(n161), .Z(n159) );
  XOR U1017 ( .A(DB[622]), .B(DB[615]), .Z(n161) );
  AND U1018 ( .A(n162), .B(n163), .Z(n160) );
  XOR U1019 ( .A(n164), .B(n165), .Z(n163) );
  XOR U1020 ( .A(DB[615]), .B(DB[608]), .Z(n165) );
  AND U1021 ( .A(n166), .B(n167), .Z(n164) );
  XOR U1022 ( .A(n168), .B(n169), .Z(n167) );
  XOR U1023 ( .A(DB[608]), .B(DB[601]), .Z(n169) );
  AND U1024 ( .A(n170), .B(n171), .Z(n168) );
  XOR U1025 ( .A(n172), .B(n173), .Z(n171) );
  XOR U1026 ( .A(DB[601]), .B(DB[594]), .Z(n173) );
  AND U1027 ( .A(n174), .B(n175), .Z(n172) );
  XOR U1028 ( .A(n176), .B(n177), .Z(n175) );
  XOR U1029 ( .A(DB[594]), .B(DB[587]), .Z(n177) );
  AND U1030 ( .A(n178), .B(n179), .Z(n176) );
  XOR U1031 ( .A(n180), .B(n181), .Z(n179) );
  XOR U1032 ( .A(DB[587]), .B(DB[580]), .Z(n181) );
  AND U1033 ( .A(n182), .B(n183), .Z(n180) );
  XOR U1034 ( .A(n184), .B(n185), .Z(n183) );
  XOR U1035 ( .A(DB[580]), .B(DB[573]), .Z(n185) );
  AND U1036 ( .A(n186), .B(n187), .Z(n184) );
  XOR U1037 ( .A(n188), .B(n189), .Z(n187) );
  XOR U1038 ( .A(DB[573]), .B(DB[566]), .Z(n189) );
  AND U1039 ( .A(n190), .B(n191), .Z(n188) );
  XOR U1040 ( .A(n192), .B(n193), .Z(n191) );
  XOR U1041 ( .A(DB[566]), .B(DB[559]), .Z(n193) );
  AND U1042 ( .A(n194), .B(n195), .Z(n192) );
  XOR U1043 ( .A(n196), .B(n197), .Z(n195) );
  XOR U1044 ( .A(DB[559]), .B(DB[552]), .Z(n197) );
  AND U1045 ( .A(n198), .B(n199), .Z(n196) );
  XOR U1046 ( .A(n200), .B(n201), .Z(n199) );
  XOR U1047 ( .A(DB[552]), .B(DB[545]), .Z(n201) );
  AND U1048 ( .A(n202), .B(n203), .Z(n200) );
  XOR U1049 ( .A(n204), .B(n205), .Z(n203) );
  XOR U1050 ( .A(DB[545]), .B(DB[538]), .Z(n205) );
  AND U1051 ( .A(n206), .B(n207), .Z(n204) );
  XOR U1052 ( .A(n208), .B(n209), .Z(n207) );
  XOR U1053 ( .A(DB[538]), .B(DB[531]), .Z(n209) );
  AND U1054 ( .A(n210), .B(n211), .Z(n208) );
  XOR U1055 ( .A(n212), .B(n213), .Z(n211) );
  XOR U1056 ( .A(DB[531]), .B(DB[524]), .Z(n213) );
  AND U1057 ( .A(n214), .B(n215), .Z(n212) );
  XOR U1058 ( .A(n216), .B(n217), .Z(n215) );
  XOR U1059 ( .A(DB[524]), .B(DB[517]), .Z(n217) );
  AND U1060 ( .A(n218), .B(n219), .Z(n216) );
  XOR U1061 ( .A(n220), .B(n221), .Z(n219) );
  XOR U1062 ( .A(DB[517]), .B(DB[510]), .Z(n221) );
  AND U1063 ( .A(n222), .B(n223), .Z(n220) );
  XOR U1064 ( .A(n224), .B(n225), .Z(n223) );
  XOR U1065 ( .A(DB[510]), .B(DB[503]), .Z(n225) );
  AND U1066 ( .A(n226), .B(n227), .Z(n224) );
  XOR U1067 ( .A(n228), .B(n229), .Z(n227) );
  XOR U1068 ( .A(DB[503]), .B(DB[496]), .Z(n229) );
  AND U1069 ( .A(n230), .B(n231), .Z(n228) );
  XOR U1070 ( .A(n232), .B(n233), .Z(n231) );
  XOR U1071 ( .A(DB[496]), .B(DB[489]), .Z(n233) );
  AND U1072 ( .A(n234), .B(n235), .Z(n232) );
  XOR U1073 ( .A(n236), .B(n237), .Z(n235) );
  XOR U1074 ( .A(DB[489]), .B(DB[482]), .Z(n237) );
  AND U1075 ( .A(n238), .B(n239), .Z(n236) );
  XOR U1076 ( .A(n240), .B(n241), .Z(n239) );
  XOR U1077 ( .A(DB[482]), .B(DB[475]), .Z(n241) );
  AND U1078 ( .A(n242), .B(n243), .Z(n240) );
  XOR U1079 ( .A(n244), .B(n245), .Z(n243) );
  XOR U1080 ( .A(DB[475]), .B(DB[468]), .Z(n245) );
  AND U1081 ( .A(n246), .B(n247), .Z(n244) );
  XOR U1082 ( .A(n248), .B(n249), .Z(n247) );
  XOR U1083 ( .A(DB[468]), .B(DB[461]), .Z(n249) );
  AND U1084 ( .A(n250), .B(n251), .Z(n248) );
  XOR U1085 ( .A(n252), .B(n253), .Z(n251) );
  XOR U1086 ( .A(DB[461]), .B(DB[454]), .Z(n253) );
  AND U1087 ( .A(n254), .B(n255), .Z(n252) );
  XOR U1088 ( .A(n256), .B(n257), .Z(n255) );
  XOR U1089 ( .A(DB[454]), .B(DB[447]), .Z(n257) );
  AND U1090 ( .A(n258), .B(n259), .Z(n256) );
  XOR U1091 ( .A(n260), .B(n261), .Z(n259) );
  XOR U1092 ( .A(DB[447]), .B(DB[440]), .Z(n261) );
  AND U1093 ( .A(n262), .B(n263), .Z(n260) );
  XOR U1094 ( .A(n264), .B(n265), .Z(n263) );
  XOR U1095 ( .A(DB[440]), .B(DB[433]), .Z(n265) );
  AND U1096 ( .A(n266), .B(n267), .Z(n264) );
  XOR U1097 ( .A(n268), .B(n269), .Z(n267) );
  XOR U1098 ( .A(DB[433]), .B(DB[426]), .Z(n269) );
  AND U1099 ( .A(n270), .B(n271), .Z(n268) );
  XOR U1100 ( .A(n272), .B(n273), .Z(n271) );
  XOR U1101 ( .A(DB[426]), .B(DB[419]), .Z(n273) );
  AND U1102 ( .A(n274), .B(n275), .Z(n272) );
  XOR U1103 ( .A(n276), .B(n277), .Z(n275) );
  XOR U1104 ( .A(DB[419]), .B(DB[412]), .Z(n277) );
  AND U1105 ( .A(n278), .B(n279), .Z(n276) );
  XOR U1106 ( .A(n280), .B(n281), .Z(n279) );
  XOR U1107 ( .A(DB[412]), .B(DB[405]), .Z(n281) );
  AND U1108 ( .A(n282), .B(n283), .Z(n280) );
  XOR U1109 ( .A(n284), .B(n285), .Z(n283) );
  XOR U1110 ( .A(DB[405]), .B(DB[398]), .Z(n285) );
  AND U1111 ( .A(n286), .B(n287), .Z(n284) );
  XOR U1112 ( .A(n288), .B(n289), .Z(n287) );
  XOR U1113 ( .A(DB[398]), .B(DB[391]), .Z(n289) );
  AND U1114 ( .A(n290), .B(n291), .Z(n288) );
  XOR U1115 ( .A(n292), .B(n293), .Z(n291) );
  XOR U1116 ( .A(DB[391]), .B(DB[384]), .Z(n293) );
  AND U1117 ( .A(n294), .B(n295), .Z(n292) );
  XOR U1118 ( .A(n296), .B(n297), .Z(n295) );
  XOR U1119 ( .A(DB[384]), .B(DB[377]), .Z(n297) );
  AND U1120 ( .A(n298), .B(n299), .Z(n296) );
  XOR U1121 ( .A(n300), .B(n301), .Z(n299) );
  XOR U1122 ( .A(DB[377]), .B(DB[370]), .Z(n301) );
  AND U1123 ( .A(n302), .B(n303), .Z(n300) );
  XOR U1124 ( .A(n304), .B(n305), .Z(n303) );
  XOR U1125 ( .A(DB[370]), .B(DB[363]), .Z(n305) );
  AND U1126 ( .A(n306), .B(n307), .Z(n304) );
  XOR U1127 ( .A(n308), .B(n309), .Z(n307) );
  XOR U1128 ( .A(DB[363]), .B(DB[356]), .Z(n309) );
  AND U1129 ( .A(n310), .B(n311), .Z(n308) );
  XOR U1130 ( .A(n312), .B(n313), .Z(n311) );
  XOR U1131 ( .A(DB[356]), .B(DB[349]), .Z(n313) );
  AND U1132 ( .A(n314), .B(n315), .Z(n312) );
  XOR U1133 ( .A(n316), .B(n317), .Z(n315) );
  XOR U1134 ( .A(DB[349]), .B(DB[342]), .Z(n317) );
  AND U1135 ( .A(n318), .B(n319), .Z(n316) );
  XOR U1136 ( .A(n320), .B(n321), .Z(n319) );
  XOR U1137 ( .A(DB[342]), .B(DB[335]), .Z(n321) );
  AND U1138 ( .A(n322), .B(n323), .Z(n320) );
  XOR U1139 ( .A(n324), .B(n325), .Z(n323) );
  XOR U1140 ( .A(DB[335]), .B(DB[328]), .Z(n325) );
  AND U1141 ( .A(n326), .B(n327), .Z(n324) );
  XOR U1142 ( .A(n328), .B(n329), .Z(n327) );
  XOR U1143 ( .A(DB[328]), .B(DB[321]), .Z(n329) );
  AND U1144 ( .A(n330), .B(n331), .Z(n328) );
  XOR U1145 ( .A(n332), .B(n333), .Z(n331) );
  XOR U1146 ( .A(DB[321]), .B(DB[314]), .Z(n333) );
  AND U1147 ( .A(n334), .B(n335), .Z(n332) );
  XOR U1148 ( .A(n336), .B(n337), .Z(n335) );
  XOR U1149 ( .A(DB[314]), .B(DB[307]), .Z(n337) );
  AND U1150 ( .A(n338), .B(n339), .Z(n336) );
  XOR U1151 ( .A(n340), .B(n341), .Z(n339) );
  XOR U1152 ( .A(DB[307]), .B(DB[300]), .Z(n341) );
  AND U1153 ( .A(n342), .B(n343), .Z(n340) );
  XOR U1154 ( .A(n344), .B(n345), .Z(n343) );
  XOR U1155 ( .A(DB[300]), .B(DB[293]), .Z(n345) );
  AND U1156 ( .A(n346), .B(n347), .Z(n344) );
  XOR U1157 ( .A(n348), .B(n349), .Z(n347) );
  XOR U1158 ( .A(DB[293]), .B(DB[286]), .Z(n349) );
  AND U1159 ( .A(n350), .B(n351), .Z(n348) );
  XOR U1160 ( .A(n352), .B(n353), .Z(n351) );
  XOR U1161 ( .A(DB[286]), .B(DB[279]), .Z(n353) );
  AND U1162 ( .A(n354), .B(n355), .Z(n352) );
  XOR U1163 ( .A(n356), .B(n357), .Z(n355) );
  XOR U1164 ( .A(DB[279]), .B(DB[272]), .Z(n357) );
  AND U1165 ( .A(n358), .B(n359), .Z(n356) );
  XOR U1166 ( .A(n360), .B(n361), .Z(n359) );
  XOR U1167 ( .A(DB[272]), .B(DB[265]), .Z(n361) );
  AND U1168 ( .A(n362), .B(n363), .Z(n360) );
  XOR U1169 ( .A(n364), .B(n365), .Z(n363) );
  XOR U1170 ( .A(DB[265]), .B(DB[258]), .Z(n365) );
  AND U1171 ( .A(n366), .B(n367), .Z(n364) );
  XOR U1172 ( .A(n368), .B(n369), .Z(n367) );
  XOR U1173 ( .A(DB[258]), .B(DB[251]), .Z(n369) );
  AND U1174 ( .A(n370), .B(n371), .Z(n368) );
  XOR U1175 ( .A(n372), .B(n373), .Z(n371) );
  XOR U1176 ( .A(DB[251]), .B(DB[244]), .Z(n373) );
  AND U1177 ( .A(n374), .B(n375), .Z(n372) );
  XOR U1178 ( .A(n376), .B(n377), .Z(n375) );
  XOR U1179 ( .A(DB[244]), .B(DB[237]), .Z(n377) );
  AND U1180 ( .A(n378), .B(n379), .Z(n376) );
  XOR U1181 ( .A(n380), .B(n381), .Z(n379) );
  XOR U1182 ( .A(DB[237]), .B(DB[230]), .Z(n381) );
  AND U1183 ( .A(n382), .B(n383), .Z(n380) );
  XOR U1184 ( .A(n384), .B(n385), .Z(n383) );
  XOR U1185 ( .A(DB[230]), .B(DB[223]), .Z(n385) );
  AND U1186 ( .A(n386), .B(n387), .Z(n384) );
  XOR U1187 ( .A(n388), .B(n389), .Z(n387) );
  XOR U1188 ( .A(DB[223]), .B(DB[216]), .Z(n389) );
  AND U1189 ( .A(n390), .B(n391), .Z(n388) );
  XOR U1190 ( .A(n392), .B(n393), .Z(n391) );
  XOR U1191 ( .A(DB[216]), .B(DB[209]), .Z(n393) );
  AND U1192 ( .A(n394), .B(n395), .Z(n392) );
  XOR U1193 ( .A(n396), .B(n397), .Z(n395) );
  XOR U1194 ( .A(DB[209]), .B(DB[202]), .Z(n397) );
  AND U1195 ( .A(n398), .B(n399), .Z(n396) );
  XOR U1196 ( .A(n400), .B(n401), .Z(n399) );
  XOR U1197 ( .A(DB[202]), .B(DB[195]), .Z(n401) );
  AND U1198 ( .A(n402), .B(n403), .Z(n400) );
  XOR U1199 ( .A(n404), .B(n405), .Z(n403) );
  XOR U1200 ( .A(DB[195]), .B(DB[188]), .Z(n405) );
  AND U1201 ( .A(n406), .B(n407), .Z(n404) );
  XOR U1202 ( .A(n408), .B(n409), .Z(n407) );
  XOR U1203 ( .A(DB[188]), .B(DB[181]), .Z(n409) );
  AND U1204 ( .A(n410), .B(n411), .Z(n408) );
  XOR U1205 ( .A(n412), .B(n413), .Z(n411) );
  XOR U1206 ( .A(DB[181]), .B(DB[174]), .Z(n413) );
  AND U1207 ( .A(n414), .B(n415), .Z(n412) );
  XOR U1208 ( .A(n416), .B(n417), .Z(n415) );
  XOR U1209 ( .A(DB[174]), .B(DB[167]), .Z(n417) );
  AND U1210 ( .A(n418), .B(n419), .Z(n416) );
  XOR U1211 ( .A(n420), .B(n421), .Z(n419) );
  XOR U1212 ( .A(DB[167]), .B(DB[160]), .Z(n421) );
  AND U1213 ( .A(n422), .B(n423), .Z(n420) );
  XOR U1214 ( .A(n424), .B(n425), .Z(n423) );
  XOR U1215 ( .A(DB[160]), .B(DB[153]), .Z(n425) );
  AND U1216 ( .A(n426), .B(n427), .Z(n424) );
  XOR U1217 ( .A(n428), .B(n429), .Z(n427) );
  XOR U1218 ( .A(DB[153]), .B(DB[146]), .Z(n429) );
  AND U1219 ( .A(n430), .B(n431), .Z(n428) );
  XOR U1220 ( .A(n432), .B(n433), .Z(n431) );
  XOR U1221 ( .A(DB[146]), .B(DB[139]), .Z(n433) );
  AND U1222 ( .A(n434), .B(n435), .Z(n432) );
  XOR U1223 ( .A(n436), .B(n437), .Z(n435) );
  XOR U1224 ( .A(DB[139]), .B(DB[132]), .Z(n437) );
  AND U1225 ( .A(n438), .B(n439), .Z(n436) );
  XOR U1226 ( .A(n440), .B(n441), .Z(n439) );
  XOR U1227 ( .A(DB[132]), .B(DB[125]), .Z(n441) );
  AND U1228 ( .A(n442), .B(n443), .Z(n440) );
  XOR U1229 ( .A(n444), .B(n445), .Z(n443) );
  XOR U1230 ( .A(DB[125]), .B(DB[118]), .Z(n445) );
  AND U1231 ( .A(n446), .B(n447), .Z(n444) );
  XOR U1232 ( .A(n448), .B(n449), .Z(n447) );
  XOR U1233 ( .A(DB[118]), .B(DB[111]), .Z(n449) );
  AND U1234 ( .A(n450), .B(n451), .Z(n448) );
  XOR U1235 ( .A(n452), .B(n453), .Z(n451) );
  XOR U1236 ( .A(DB[111]), .B(DB[104]), .Z(n453) );
  AND U1237 ( .A(n454), .B(n455), .Z(n452) );
  XOR U1238 ( .A(n456), .B(n457), .Z(n455) );
  XOR U1239 ( .A(DB[97]), .B(DB[104]), .Z(n457) );
  AND U1240 ( .A(n458), .B(n459), .Z(n456) );
  XOR U1241 ( .A(n460), .B(n461), .Z(n459) );
  XOR U1242 ( .A(DB[97]), .B(DB[90]), .Z(n461) );
  AND U1243 ( .A(n462), .B(n463), .Z(n460) );
  XOR U1244 ( .A(n464), .B(n465), .Z(n463) );
  XOR U1245 ( .A(DB[90]), .B(DB[83]), .Z(n465) );
  AND U1246 ( .A(n466), .B(n467), .Z(n464) );
  XOR U1247 ( .A(n468), .B(n469), .Z(n467) );
  XOR U1248 ( .A(DB[83]), .B(DB[76]), .Z(n469) );
  AND U1249 ( .A(n470), .B(n471), .Z(n468) );
  XOR U1250 ( .A(n472), .B(n473), .Z(n471) );
  XOR U1251 ( .A(DB[76]), .B(DB[69]), .Z(n473) );
  AND U1252 ( .A(n474), .B(n475), .Z(n472) );
  XOR U1253 ( .A(n476), .B(n477), .Z(n475) );
  XOR U1254 ( .A(DB[69]), .B(DB[62]), .Z(n477) );
  AND U1255 ( .A(n478), .B(n479), .Z(n476) );
  XOR U1256 ( .A(n480), .B(n481), .Z(n479) );
  XOR U1257 ( .A(DB[62]), .B(DB[55]), .Z(n481) );
  AND U1258 ( .A(n482), .B(n483), .Z(n480) );
  XOR U1259 ( .A(n484), .B(n485), .Z(n483) );
  XOR U1260 ( .A(DB[55]), .B(DB[48]), .Z(n485) );
  AND U1261 ( .A(n486), .B(n487), .Z(n484) );
  XOR U1262 ( .A(n488), .B(n489), .Z(n487) );
  XOR U1263 ( .A(DB[48]), .B(DB[41]), .Z(n489) );
  AND U1264 ( .A(n490), .B(n491), .Z(n488) );
  XOR U1265 ( .A(n492), .B(n493), .Z(n491) );
  XOR U1266 ( .A(DB[41]), .B(DB[34]), .Z(n493) );
  AND U1267 ( .A(n494), .B(n495), .Z(n492) );
  XOR U1268 ( .A(n496), .B(n497), .Z(n495) );
  XOR U1269 ( .A(DB[34]), .B(DB[27]), .Z(n497) );
  AND U1270 ( .A(n498), .B(n499), .Z(n496) );
  XOR U1271 ( .A(n500), .B(n501), .Z(n499) );
  XOR U1272 ( .A(DB[27]), .B(DB[20]), .Z(n501) );
  AND U1273 ( .A(n502), .B(n503), .Z(n500) );
  XOR U1274 ( .A(n504), .B(n505), .Z(n503) );
  XOR U1275 ( .A(DB[20]), .B(DB[13]), .Z(n505) );
  AND U1276 ( .A(n506), .B(n507), .Z(n504) );
  XOR U1277 ( .A(DB[6]), .B(DB[13]), .Z(n507) );
  XOR U1278 ( .A(DB[894]), .B(n508), .Z(min_val_out[5]) );
  AND U1279 ( .A(n2), .B(n509), .Z(n508) );
  XOR U1280 ( .A(n510), .B(n511), .Z(n509) );
  XOR U1281 ( .A(DB[894]), .B(DB[887]), .Z(n511) );
  AND U1282 ( .A(n6), .B(n512), .Z(n510) );
  XOR U1283 ( .A(n513), .B(n514), .Z(n512) );
  XOR U1284 ( .A(DB[887]), .B(DB[880]), .Z(n514) );
  AND U1285 ( .A(n10), .B(n515), .Z(n513) );
  XOR U1286 ( .A(n516), .B(n517), .Z(n515) );
  XOR U1287 ( .A(DB[880]), .B(DB[873]), .Z(n517) );
  AND U1288 ( .A(n14), .B(n518), .Z(n516) );
  XOR U1289 ( .A(n519), .B(n520), .Z(n518) );
  XOR U1290 ( .A(DB[873]), .B(DB[866]), .Z(n520) );
  AND U1291 ( .A(n18), .B(n521), .Z(n519) );
  XOR U1292 ( .A(n522), .B(n523), .Z(n521) );
  XOR U1293 ( .A(DB[866]), .B(DB[859]), .Z(n523) );
  AND U1294 ( .A(n22), .B(n524), .Z(n522) );
  XOR U1295 ( .A(n525), .B(n526), .Z(n524) );
  XOR U1296 ( .A(DB[859]), .B(DB[852]), .Z(n526) );
  AND U1297 ( .A(n26), .B(n527), .Z(n525) );
  XOR U1298 ( .A(n528), .B(n529), .Z(n527) );
  XOR U1299 ( .A(DB[852]), .B(DB[845]), .Z(n529) );
  AND U1300 ( .A(n30), .B(n530), .Z(n528) );
  XOR U1301 ( .A(n531), .B(n532), .Z(n530) );
  XOR U1302 ( .A(DB[845]), .B(DB[838]), .Z(n532) );
  AND U1303 ( .A(n34), .B(n533), .Z(n531) );
  XOR U1304 ( .A(n534), .B(n535), .Z(n533) );
  XOR U1305 ( .A(DB[838]), .B(DB[831]), .Z(n535) );
  AND U1306 ( .A(n38), .B(n536), .Z(n534) );
  XOR U1307 ( .A(n537), .B(n538), .Z(n536) );
  XOR U1308 ( .A(DB[831]), .B(DB[824]), .Z(n538) );
  AND U1309 ( .A(n42), .B(n539), .Z(n537) );
  XOR U1310 ( .A(n540), .B(n541), .Z(n539) );
  XOR U1311 ( .A(DB[824]), .B(DB[817]), .Z(n541) );
  AND U1312 ( .A(n46), .B(n542), .Z(n540) );
  XOR U1313 ( .A(n543), .B(n544), .Z(n542) );
  XOR U1314 ( .A(DB[817]), .B(DB[810]), .Z(n544) );
  AND U1315 ( .A(n50), .B(n545), .Z(n543) );
  XOR U1316 ( .A(n546), .B(n547), .Z(n545) );
  XOR U1317 ( .A(DB[810]), .B(DB[803]), .Z(n547) );
  AND U1318 ( .A(n54), .B(n548), .Z(n546) );
  XOR U1319 ( .A(n549), .B(n550), .Z(n548) );
  XOR U1320 ( .A(DB[803]), .B(DB[796]), .Z(n550) );
  AND U1321 ( .A(n58), .B(n551), .Z(n549) );
  XOR U1322 ( .A(n552), .B(n553), .Z(n551) );
  XOR U1323 ( .A(DB[796]), .B(DB[789]), .Z(n553) );
  AND U1324 ( .A(n62), .B(n554), .Z(n552) );
  XOR U1325 ( .A(n555), .B(n556), .Z(n554) );
  XOR U1326 ( .A(DB[789]), .B(DB[782]), .Z(n556) );
  AND U1327 ( .A(n66), .B(n557), .Z(n555) );
  XOR U1328 ( .A(n558), .B(n559), .Z(n557) );
  XOR U1329 ( .A(DB[782]), .B(DB[775]), .Z(n559) );
  AND U1330 ( .A(n70), .B(n560), .Z(n558) );
  XOR U1331 ( .A(n561), .B(n562), .Z(n560) );
  XOR U1332 ( .A(DB[775]), .B(DB[768]), .Z(n562) );
  AND U1333 ( .A(n74), .B(n563), .Z(n561) );
  XOR U1334 ( .A(n564), .B(n565), .Z(n563) );
  XOR U1335 ( .A(DB[768]), .B(DB[761]), .Z(n565) );
  AND U1336 ( .A(n78), .B(n566), .Z(n564) );
  XOR U1337 ( .A(n567), .B(n568), .Z(n566) );
  XOR U1338 ( .A(DB[761]), .B(DB[754]), .Z(n568) );
  AND U1339 ( .A(n82), .B(n569), .Z(n567) );
  XOR U1340 ( .A(n570), .B(n571), .Z(n569) );
  XOR U1341 ( .A(DB[754]), .B(DB[747]), .Z(n571) );
  AND U1342 ( .A(n86), .B(n572), .Z(n570) );
  XOR U1343 ( .A(n573), .B(n574), .Z(n572) );
  XOR U1344 ( .A(DB[747]), .B(DB[740]), .Z(n574) );
  AND U1345 ( .A(n90), .B(n575), .Z(n573) );
  XOR U1346 ( .A(n576), .B(n577), .Z(n575) );
  XOR U1347 ( .A(DB[740]), .B(DB[733]), .Z(n577) );
  AND U1348 ( .A(n94), .B(n578), .Z(n576) );
  XOR U1349 ( .A(n579), .B(n580), .Z(n578) );
  XOR U1350 ( .A(DB[733]), .B(DB[726]), .Z(n580) );
  AND U1351 ( .A(n98), .B(n581), .Z(n579) );
  XOR U1352 ( .A(n582), .B(n583), .Z(n581) );
  XOR U1353 ( .A(DB[726]), .B(DB[719]), .Z(n583) );
  AND U1354 ( .A(n102), .B(n584), .Z(n582) );
  XOR U1355 ( .A(n585), .B(n586), .Z(n584) );
  XOR U1356 ( .A(DB[719]), .B(DB[712]), .Z(n586) );
  AND U1357 ( .A(n106), .B(n587), .Z(n585) );
  XOR U1358 ( .A(n588), .B(n589), .Z(n587) );
  XOR U1359 ( .A(DB[712]), .B(DB[705]), .Z(n589) );
  AND U1360 ( .A(n110), .B(n590), .Z(n588) );
  XOR U1361 ( .A(n591), .B(n592), .Z(n590) );
  XOR U1362 ( .A(DB[705]), .B(DB[698]), .Z(n592) );
  AND U1363 ( .A(n114), .B(n593), .Z(n591) );
  XOR U1364 ( .A(n594), .B(n595), .Z(n593) );
  XOR U1365 ( .A(DB[698]), .B(DB[691]), .Z(n595) );
  AND U1366 ( .A(n118), .B(n596), .Z(n594) );
  XOR U1367 ( .A(n597), .B(n598), .Z(n596) );
  XOR U1368 ( .A(DB[691]), .B(DB[684]), .Z(n598) );
  AND U1369 ( .A(n122), .B(n599), .Z(n597) );
  XOR U1370 ( .A(n600), .B(n601), .Z(n599) );
  XOR U1371 ( .A(DB[684]), .B(DB[677]), .Z(n601) );
  AND U1372 ( .A(n126), .B(n602), .Z(n600) );
  XOR U1373 ( .A(n603), .B(n604), .Z(n602) );
  XOR U1374 ( .A(DB[677]), .B(DB[670]), .Z(n604) );
  AND U1375 ( .A(n130), .B(n605), .Z(n603) );
  XOR U1376 ( .A(n606), .B(n607), .Z(n605) );
  XOR U1377 ( .A(DB[670]), .B(DB[663]), .Z(n607) );
  AND U1378 ( .A(n134), .B(n608), .Z(n606) );
  XOR U1379 ( .A(n609), .B(n610), .Z(n608) );
  XOR U1380 ( .A(DB[663]), .B(DB[656]), .Z(n610) );
  AND U1381 ( .A(n138), .B(n611), .Z(n609) );
  XOR U1382 ( .A(n612), .B(n613), .Z(n611) );
  XOR U1383 ( .A(DB[656]), .B(DB[649]), .Z(n613) );
  AND U1384 ( .A(n142), .B(n614), .Z(n612) );
  XOR U1385 ( .A(n615), .B(n616), .Z(n614) );
  XOR U1386 ( .A(DB[649]), .B(DB[642]), .Z(n616) );
  AND U1387 ( .A(n146), .B(n617), .Z(n615) );
  XOR U1388 ( .A(n618), .B(n619), .Z(n617) );
  XOR U1389 ( .A(DB[642]), .B(DB[635]), .Z(n619) );
  AND U1390 ( .A(n150), .B(n620), .Z(n618) );
  XOR U1391 ( .A(n621), .B(n622), .Z(n620) );
  XOR U1392 ( .A(DB[635]), .B(DB[628]), .Z(n622) );
  AND U1393 ( .A(n154), .B(n623), .Z(n621) );
  XOR U1394 ( .A(n624), .B(n625), .Z(n623) );
  XOR U1395 ( .A(DB[628]), .B(DB[621]), .Z(n625) );
  AND U1396 ( .A(n158), .B(n626), .Z(n624) );
  XOR U1397 ( .A(n627), .B(n628), .Z(n626) );
  XOR U1398 ( .A(DB[621]), .B(DB[614]), .Z(n628) );
  AND U1399 ( .A(n162), .B(n629), .Z(n627) );
  XOR U1400 ( .A(n630), .B(n631), .Z(n629) );
  XOR U1401 ( .A(DB[614]), .B(DB[607]), .Z(n631) );
  AND U1402 ( .A(n166), .B(n632), .Z(n630) );
  XOR U1403 ( .A(n633), .B(n634), .Z(n632) );
  XOR U1404 ( .A(DB[607]), .B(DB[600]), .Z(n634) );
  AND U1405 ( .A(n170), .B(n635), .Z(n633) );
  XOR U1406 ( .A(n636), .B(n637), .Z(n635) );
  XOR U1407 ( .A(DB[600]), .B(DB[593]), .Z(n637) );
  AND U1408 ( .A(n174), .B(n638), .Z(n636) );
  XOR U1409 ( .A(n639), .B(n640), .Z(n638) );
  XOR U1410 ( .A(DB[593]), .B(DB[586]), .Z(n640) );
  AND U1411 ( .A(n178), .B(n641), .Z(n639) );
  XOR U1412 ( .A(n642), .B(n643), .Z(n641) );
  XOR U1413 ( .A(DB[586]), .B(DB[579]), .Z(n643) );
  AND U1414 ( .A(n182), .B(n644), .Z(n642) );
  XOR U1415 ( .A(n645), .B(n646), .Z(n644) );
  XOR U1416 ( .A(DB[579]), .B(DB[572]), .Z(n646) );
  AND U1417 ( .A(n186), .B(n647), .Z(n645) );
  XOR U1418 ( .A(n648), .B(n649), .Z(n647) );
  XOR U1419 ( .A(DB[572]), .B(DB[565]), .Z(n649) );
  AND U1420 ( .A(n190), .B(n650), .Z(n648) );
  XOR U1421 ( .A(n651), .B(n652), .Z(n650) );
  XOR U1422 ( .A(DB[565]), .B(DB[558]), .Z(n652) );
  AND U1423 ( .A(n194), .B(n653), .Z(n651) );
  XOR U1424 ( .A(n654), .B(n655), .Z(n653) );
  XOR U1425 ( .A(DB[558]), .B(DB[551]), .Z(n655) );
  AND U1426 ( .A(n198), .B(n656), .Z(n654) );
  XOR U1427 ( .A(n657), .B(n658), .Z(n656) );
  XOR U1428 ( .A(DB[551]), .B(DB[544]), .Z(n658) );
  AND U1429 ( .A(n202), .B(n659), .Z(n657) );
  XOR U1430 ( .A(n660), .B(n661), .Z(n659) );
  XOR U1431 ( .A(DB[544]), .B(DB[537]), .Z(n661) );
  AND U1432 ( .A(n206), .B(n662), .Z(n660) );
  XOR U1433 ( .A(n663), .B(n664), .Z(n662) );
  XOR U1434 ( .A(DB[537]), .B(DB[530]), .Z(n664) );
  AND U1435 ( .A(n210), .B(n665), .Z(n663) );
  XOR U1436 ( .A(n666), .B(n667), .Z(n665) );
  XOR U1437 ( .A(DB[530]), .B(DB[523]), .Z(n667) );
  AND U1438 ( .A(n214), .B(n668), .Z(n666) );
  XOR U1439 ( .A(n669), .B(n670), .Z(n668) );
  XOR U1440 ( .A(DB[523]), .B(DB[516]), .Z(n670) );
  AND U1441 ( .A(n218), .B(n671), .Z(n669) );
  XOR U1442 ( .A(n672), .B(n673), .Z(n671) );
  XOR U1443 ( .A(DB[516]), .B(DB[509]), .Z(n673) );
  AND U1444 ( .A(n222), .B(n674), .Z(n672) );
  XOR U1445 ( .A(n675), .B(n676), .Z(n674) );
  XOR U1446 ( .A(DB[509]), .B(DB[502]), .Z(n676) );
  AND U1447 ( .A(n226), .B(n677), .Z(n675) );
  XOR U1448 ( .A(n678), .B(n679), .Z(n677) );
  XOR U1449 ( .A(DB[502]), .B(DB[495]), .Z(n679) );
  AND U1450 ( .A(n230), .B(n680), .Z(n678) );
  XOR U1451 ( .A(n681), .B(n682), .Z(n680) );
  XOR U1452 ( .A(DB[495]), .B(DB[488]), .Z(n682) );
  AND U1453 ( .A(n234), .B(n683), .Z(n681) );
  XOR U1454 ( .A(n684), .B(n685), .Z(n683) );
  XOR U1455 ( .A(DB[488]), .B(DB[481]), .Z(n685) );
  AND U1456 ( .A(n238), .B(n686), .Z(n684) );
  XOR U1457 ( .A(n687), .B(n688), .Z(n686) );
  XOR U1458 ( .A(DB[481]), .B(DB[474]), .Z(n688) );
  AND U1459 ( .A(n242), .B(n689), .Z(n687) );
  XOR U1460 ( .A(n690), .B(n691), .Z(n689) );
  XOR U1461 ( .A(DB[474]), .B(DB[467]), .Z(n691) );
  AND U1462 ( .A(n246), .B(n692), .Z(n690) );
  XOR U1463 ( .A(n693), .B(n694), .Z(n692) );
  XOR U1464 ( .A(DB[467]), .B(DB[460]), .Z(n694) );
  AND U1465 ( .A(n250), .B(n695), .Z(n693) );
  XOR U1466 ( .A(n696), .B(n697), .Z(n695) );
  XOR U1467 ( .A(DB[460]), .B(DB[453]), .Z(n697) );
  AND U1468 ( .A(n254), .B(n698), .Z(n696) );
  XOR U1469 ( .A(n699), .B(n700), .Z(n698) );
  XOR U1470 ( .A(DB[453]), .B(DB[446]), .Z(n700) );
  AND U1471 ( .A(n258), .B(n701), .Z(n699) );
  XOR U1472 ( .A(n702), .B(n703), .Z(n701) );
  XOR U1473 ( .A(DB[446]), .B(DB[439]), .Z(n703) );
  AND U1474 ( .A(n262), .B(n704), .Z(n702) );
  XOR U1475 ( .A(n705), .B(n706), .Z(n704) );
  XOR U1476 ( .A(DB[439]), .B(DB[432]), .Z(n706) );
  AND U1477 ( .A(n266), .B(n707), .Z(n705) );
  XOR U1478 ( .A(n708), .B(n709), .Z(n707) );
  XOR U1479 ( .A(DB[432]), .B(DB[425]), .Z(n709) );
  AND U1480 ( .A(n270), .B(n710), .Z(n708) );
  XOR U1481 ( .A(n711), .B(n712), .Z(n710) );
  XOR U1482 ( .A(DB[425]), .B(DB[418]), .Z(n712) );
  AND U1483 ( .A(n274), .B(n713), .Z(n711) );
  XOR U1484 ( .A(n714), .B(n715), .Z(n713) );
  XOR U1485 ( .A(DB[418]), .B(DB[411]), .Z(n715) );
  AND U1486 ( .A(n278), .B(n716), .Z(n714) );
  XOR U1487 ( .A(n717), .B(n718), .Z(n716) );
  XOR U1488 ( .A(DB[411]), .B(DB[404]), .Z(n718) );
  AND U1489 ( .A(n282), .B(n719), .Z(n717) );
  XOR U1490 ( .A(n720), .B(n721), .Z(n719) );
  XOR U1491 ( .A(DB[404]), .B(DB[397]), .Z(n721) );
  AND U1492 ( .A(n286), .B(n722), .Z(n720) );
  XOR U1493 ( .A(n723), .B(n724), .Z(n722) );
  XOR U1494 ( .A(DB[397]), .B(DB[390]), .Z(n724) );
  AND U1495 ( .A(n290), .B(n725), .Z(n723) );
  XOR U1496 ( .A(n726), .B(n727), .Z(n725) );
  XOR U1497 ( .A(DB[390]), .B(DB[383]), .Z(n727) );
  AND U1498 ( .A(n294), .B(n728), .Z(n726) );
  XOR U1499 ( .A(n729), .B(n730), .Z(n728) );
  XOR U1500 ( .A(DB[383]), .B(DB[376]), .Z(n730) );
  AND U1501 ( .A(n298), .B(n731), .Z(n729) );
  XOR U1502 ( .A(n732), .B(n733), .Z(n731) );
  XOR U1503 ( .A(DB[376]), .B(DB[369]), .Z(n733) );
  AND U1504 ( .A(n302), .B(n734), .Z(n732) );
  XOR U1505 ( .A(n735), .B(n736), .Z(n734) );
  XOR U1506 ( .A(DB[369]), .B(DB[362]), .Z(n736) );
  AND U1507 ( .A(n306), .B(n737), .Z(n735) );
  XOR U1508 ( .A(n738), .B(n739), .Z(n737) );
  XOR U1509 ( .A(DB[362]), .B(DB[355]), .Z(n739) );
  AND U1510 ( .A(n310), .B(n740), .Z(n738) );
  XOR U1511 ( .A(n741), .B(n742), .Z(n740) );
  XOR U1512 ( .A(DB[355]), .B(DB[348]), .Z(n742) );
  AND U1513 ( .A(n314), .B(n743), .Z(n741) );
  XOR U1514 ( .A(n744), .B(n745), .Z(n743) );
  XOR U1515 ( .A(DB[348]), .B(DB[341]), .Z(n745) );
  AND U1516 ( .A(n318), .B(n746), .Z(n744) );
  XOR U1517 ( .A(n747), .B(n748), .Z(n746) );
  XOR U1518 ( .A(DB[341]), .B(DB[334]), .Z(n748) );
  AND U1519 ( .A(n322), .B(n749), .Z(n747) );
  XOR U1520 ( .A(n750), .B(n751), .Z(n749) );
  XOR U1521 ( .A(DB[334]), .B(DB[327]), .Z(n751) );
  AND U1522 ( .A(n326), .B(n752), .Z(n750) );
  XOR U1523 ( .A(n753), .B(n754), .Z(n752) );
  XOR U1524 ( .A(DB[327]), .B(DB[320]), .Z(n754) );
  AND U1525 ( .A(n330), .B(n755), .Z(n753) );
  XOR U1526 ( .A(n756), .B(n757), .Z(n755) );
  XOR U1527 ( .A(DB[320]), .B(DB[313]), .Z(n757) );
  AND U1528 ( .A(n334), .B(n758), .Z(n756) );
  XOR U1529 ( .A(n759), .B(n760), .Z(n758) );
  XOR U1530 ( .A(DB[313]), .B(DB[306]), .Z(n760) );
  AND U1531 ( .A(n338), .B(n761), .Z(n759) );
  XOR U1532 ( .A(n762), .B(n763), .Z(n761) );
  XOR U1533 ( .A(DB[306]), .B(DB[299]), .Z(n763) );
  AND U1534 ( .A(n342), .B(n764), .Z(n762) );
  XOR U1535 ( .A(n765), .B(n766), .Z(n764) );
  XOR U1536 ( .A(DB[299]), .B(DB[292]), .Z(n766) );
  AND U1537 ( .A(n346), .B(n767), .Z(n765) );
  XOR U1538 ( .A(n768), .B(n769), .Z(n767) );
  XOR U1539 ( .A(DB[292]), .B(DB[285]), .Z(n769) );
  AND U1540 ( .A(n350), .B(n770), .Z(n768) );
  XOR U1541 ( .A(n771), .B(n772), .Z(n770) );
  XOR U1542 ( .A(DB[285]), .B(DB[278]), .Z(n772) );
  AND U1543 ( .A(n354), .B(n773), .Z(n771) );
  XOR U1544 ( .A(n774), .B(n775), .Z(n773) );
  XOR U1545 ( .A(DB[278]), .B(DB[271]), .Z(n775) );
  AND U1546 ( .A(n358), .B(n776), .Z(n774) );
  XOR U1547 ( .A(n777), .B(n778), .Z(n776) );
  XOR U1548 ( .A(DB[271]), .B(DB[264]), .Z(n778) );
  AND U1549 ( .A(n362), .B(n779), .Z(n777) );
  XOR U1550 ( .A(n780), .B(n781), .Z(n779) );
  XOR U1551 ( .A(DB[264]), .B(DB[257]), .Z(n781) );
  AND U1552 ( .A(n366), .B(n782), .Z(n780) );
  XOR U1553 ( .A(n783), .B(n784), .Z(n782) );
  XOR U1554 ( .A(DB[257]), .B(DB[250]), .Z(n784) );
  AND U1555 ( .A(n370), .B(n785), .Z(n783) );
  XOR U1556 ( .A(n786), .B(n787), .Z(n785) );
  XOR U1557 ( .A(DB[250]), .B(DB[243]), .Z(n787) );
  AND U1558 ( .A(n374), .B(n788), .Z(n786) );
  XOR U1559 ( .A(n789), .B(n790), .Z(n788) );
  XOR U1560 ( .A(DB[243]), .B(DB[236]), .Z(n790) );
  AND U1561 ( .A(n378), .B(n791), .Z(n789) );
  XOR U1562 ( .A(n792), .B(n793), .Z(n791) );
  XOR U1563 ( .A(DB[236]), .B(DB[229]), .Z(n793) );
  AND U1564 ( .A(n382), .B(n794), .Z(n792) );
  XOR U1565 ( .A(n795), .B(n796), .Z(n794) );
  XOR U1566 ( .A(DB[229]), .B(DB[222]), .Z(n796) );
  AND U1567 ( .A(n386), .B(n797), .Z(n795) );
  XOR U1568 ( .A(n798), .B(n799), .Z(n797) );
  XOR U1569 ( .A(DB[222]), .B(DB[215]), .Z(n799) );
  AND U1570 ( .A(n390), .B(n800), .Z(n798) );
  XOR U1571 ( .A(n801), .B(n802), .Z(n800) );
  XOR U1572 ( .A(DB[215]), .B(DB[208]), .Z(n802) );
  AND U1573 ( .A(n394), .B(n803), .Z(n801) );
  XOR U1574 ( .A(n804), .B(n805), .Z(n803) );
  XOR U1575 ( .A(DB[208]), .B(DB[201]), .Z(n805) );
  AND U1576 ( .A(n398), .B(n806), .Z(n804) );
  XOR U1577 ( .A(n807), .B(n808), .Z(n806) );
  XOR U1578 ( .A(DB[201]), .B(DB[194]), .Z(n808) );
  AND U1579 ( .A(n402), .B(n809), .Z(n807) );
  XOR U1580 ( .A(n810), .B(n811), .Z(n809) );
  XOR U1581 ( .A(DB[194]), .B(DB[187]), .Z(n811) );
  AND U1582 ( .A(n406), .B(n812), .Z(n810) );
  XOR U1583 ( .A(n813), .B(n814), .Z(n812) );
  XOR U1584 ( .A(DB[187]), .B(DB[180]), .Z(n814) );
  AND U1585 ( .A(n410), .B(n815), .Z(n813) );
  XOR U1586 ( .A(n816), .B(n817), .Z(n815) );
  XOR U1587 ( .A(DB[180]), .B(DB[173]), .Z(n817) );
  AND U1588 ( .A(n414), .B(n818), .Z(n816) );
  XOR U1589 ( .A(n819), .B(n820), .Z(n818) );
  XOR U1590 ( .A(DB[173]), .B(DB[166]), .Z(n820) );
  AND U1591 ( .A(n418), .B(n821), .Z(n819) );
  XOR U1592 ( .A(n822), .B(n823), .Z(n821) );
  XOR U1593 ( .A(DB[166]), .B(DB[159]), .Z(n823) );
  AND U1594 ( .A(n422), .B(n824), .Z(n822) );
  XOR U1595 ( .A(n825), .B(n826), .Z(n824) );
  XOR U1596 ( .A(DB[159]), .B(DB[152]), .Z(n826) );
  AND U1597 ( .A(n426), .B(n827), .Z(n825) );
  XOR U1598 ( .A(n828), .B(n829), .Z(n827) );
  XOR U1599 ( .A(DB[152]), .B(DB[145]), .Z(n829) );
  AND U1600 ( .A(n430), .B(n830), .Z(n828) );
  XOR U1601 ( .A(n831), .B(n832), .Z(n830) );
  XOR U1602 ( .A(DB[145]), .B(DB[138]), .Z(n832) );
  AND U1603 ( .A(n434), .B(n833), .Z(n831) );
  XOR U1604 ( .A(n834), .B(n835), .Z(n833) );
  XOR U1605 ( .A(DB[138]), .B(DB[131]), .Z(n835) );
  AND U1606 ( .A(n438), .B(n836), .Z(n834) );
  XOR U1607 ( .A(n837), .B(n838), .Z(n836) );
  XOR U1608 ( .A(DB[131]), .B(DB[124]), .Z(n838) );
  AND U1609 ( .A(n442), .B(n839), .Z(n837) );
  XOR U1610 ( .A(n840), .B(n841), .Z(n839) );
  XOR U1611 ( .A(DB[124]), .B(DB[117]), .Z(n841) );
  AND U1612 ( .A(n446), .B(n842), .Z(n840) );
  XOR U1613 ( .A(n843), .B(n844), .Z(n842) );
  XOR U1614 ( .A(DB[117]), .B(DB[110]), .Z(n844) );
  AND U1615 ( .A(n450), .B(n845), .Z(n843) );
  XOR U1616 ( .A(n846), .B(n847), .Z(n845) );
  XOR U1617 ( .A(DB[110]), .B(DB[103]), .Z(n847) );
  AND U1618 ( .A(n454), .B(n848), .Z(n846) );
  XOR U1619 ( .A(n849), .B(n850), .Z(n848) );
  XOR U1620 ( .A(DB[96]), .B(DB[103]), .Z(n850) );
  AND U1621 ( .A(n458), .B(n851), .Z(n849) );
  XOR U1622 ( .A(n852), .B(n853), .Z(n851) );
  XOR U1623 ( .A(DB[96]), .B(DB[89]), .Z(n853) );
  AND U1624 ( .A(n462), .B(n854), .Z(n852) );
  XOR U1625 ( .A(n855), .B(n856), .Z(n854) );
  XOR U1626 ( .A(DB[89]), .B(DB[82]), .Z(n856) );
  AND U1627 ( .A(n466), .B(n857), .Z(n855) );
  XOR U1628 ( .A(n858), .B(n859), .Z(n857) );
  XOR U1629 ( .A(DB[82]), .B(DB[75]), .Z(n859) );
  AND U1630 ( .A(n470), .B(n860), .Z(n858) );
  XOR U1631 ( .A(n861), .B(n862), .Z(n860) );
  XOR U1632 ( .A(DB[75]), .B(DB[68]), .Z(n862) );
  AND U1633 ( .A(n474), .B(n863), .Z(n861) );
  XOR U1634 ( .A(n864), .B(n865), .Z(n863) );
  XOR U1635 ( .A(DB[68]), .B(DB[61]), .Z(n865) );
  AND U1636 ( .A(n478), .B(n866), .Z(n864) );
  XOR U1637 ( .A(n867), .B(n868), .Z(n866) );
  XOR U1638 ( .A(DB[61]), .B(DB[54]), .Z(n868) );
  AND U1639 ( .A(n482), .B(n869), .Z(n867) );
  XOR U1640 ( .A(n870), .B(n871), .Z(n869) );
  XOR U1641 ( .A(DB[54]), .B(DB[47]), .Z(n871) );
  AND U1642 ( .A(n486), .B(n872), .Z(n870) );
  XOR U1643 ( .A(n873), .B(n874), .Z(n872) );
  XOR U1644 ( .A(DB[47]), .B(DB[40]), .Z(n874) );
  AND U1645 ( .A(n490), .B(n875), .Z(n873) );
  XOR U1646 ( .A(n876), .B(n877), .Z(n875) );
  XOR U1647 ( .A(DB[40]), .B(DB[33]), .Z(n877) );
  AND U1648 ( .A(n494), .B(n878), .Z(n876) );
  XOR U1649 ( .A(n879), .B(n880), .Z(n878) );
  XOR U1650 ( .A(DB[33]), .B(DB[26]), .Z(n880) );
  AND U1651 ( .A(n498), .B(n881), .Z(n879) );
  XOR U1652 ( .A(n882), .B(n883), .Z(n881) );
  XOR U1653 ( .A(DB[26]), .B(DB[19]), .Z(n883) );
  AND U1654 ( .A(n502), .B(n884), .Z(n882) );
  XOR U1655 ( .A(n885), .B(n886), .Z(n884) );
  XOR U1656 ( .A(DB[19]), .B(DB[12]), .Z(n886) );
  AND U1657 ( .A(n506), .B(n887), .Z(n885) );
  XOR U1658 ( .A(DB[5]), .B(DB[12]), .Z(n887) );
  XOR U1659 ( .A(DB[893]), .B(n888), .Z(min_val_out[4]) );
  AND U1660 ( .A(n2), .B(n889), .Z(n888) );
  XOR U1661 ( .A(n890), .B(n891), .Z(n889) );
  XOR U1662 ( .A(n892), .B(n893), .Z(n891) );
  IV U1663 ( .A(DB[893]), .Z(n892) );
  AND U1664 ( .A(n6), .B(n894), .Z(n890) );
  XOR U1665 ( .A(n895), .B(n896), .Z(n894) );
  XOR U1666 ( .A(DB[886]), .B(DB[879]), .Z(n896) );
  AND U1667 ( .A(n10), .B(n897), .Z(n895) );
  XOR U1668 ( .A(n898), .B(n899), .Z(n897) );
  XOR U1669 ( .A(DB[879]), .B(DB[872]), .Z(n899) );
  AND U1670 ( .A(n14), .B(n900), .Z(n898) );
  XOR U1671 ( .A(n901), .B(n902), .Z(n900) );
  XOR U1672 ( .A(DB[872]), .B(DB[865]), .Z(n902) );
  AND U1673 ( .A(n18), .B(n903), .Z(n901) );
  XOR U1674 ( .A(n904), .B(n905), .Z(n903) );
  XOR U1675 ( .A(DB[865]), .B(DB[858]), .Z(n905) );
  AND U1676 ( .A(n22), .B(n906), .Z(n904) );
  XOR U1677 ( .A(n907), .B(n908), .Z(n906) );
  XOR U1678 ( .A(DB[858]), .B(DB[851]), .Z(n908) );
  AND U1679 ( .A(n26), .B(n909), .Z(n907) );
  XOR U1680 ( .A(n910), .B(n911), .Z(n909) );
  XOR U1681 ( .A(DB[851]), .B(DB[844]), .Z(n911) );
  AND U1682 ( .A(n30), .B(n912), .Z(n910) );
  XOR U1683 ( .A(n913), .B(n914), .Z(n912) );
  XOR U1684 ( .A(DB[844]), .B(DB[837]), .Z(n914) );
  AND U1685 ( .A(n34), .B(n915), .Z(n913) );
  XOR U1686 ( .A(n916), .B(n917), .Z(n915) );
  XOR U1687 ( .A(DB[837]), .B(DB[830]), .Z(n917) );
  AND U1688 ( .A(n38), .B(n918), .Z(n916) );
  XOR U1689 ( .A(n919), .B(n920), .Z(n918) );
  XOR U1690 ( .A(DB[830]), .B(DB[823]), .Z(n920) );
  AND U1691 ( .A(n42), .B(n921), .Z(n919) );
  XOR U1692 ( .A(n922), .B(n923), .Z(n921) );
  XOR U1693 ( .A(DB[823]), .B(DB[816]), .Z(n923) );
  AND U1694 ( .A(n46), .B(n924), .Z(n922) );
  XOR U1695 ( .A(n925), .B(n926), .Z(n924) );
  XOR U1696 ( .A(DB[816]), .B(DB[809]), .Z(n926) );
  AND U1697 ( .A(n50), .B(n927), .Z(n925) );
  XOR U1698 ( .A(n928), .B(n929), .Z(n927) );
  XOR U1699 ( .A(DB[809]), .B(DB[802]), .Z(n929) );
  AND U1700 ( .A(n54), .B(n930), .Z(n928) );
  XOR U1701 ( .A(n931), .B(n932), .Z(n930) );
  XOR U1702 ( .A(DB[802]), .B(DB[795]), .Z(n932) );
  AND U1703 ( .A(n58), .B(n933), .Z(n931) );
  XOR U1704 ( .A(n934), .B(n935), .Z(n933) );
  XOR U1705 ( .A(DB[795]), .B(DB[788]), .Z(n935) );
  AND U1706 ( .A(n62), .B(n936), .Z(n934) );
  XOR U1707 ( .A(n937), .B(n938), .Z(n936) );
  XOR U1708 ( .A(DB[788]), .B(DB[781]), .Z(n938) );
  AND U1709 ( .A(n66), .B(n939), .Z(n937) );
  XOR U1710 ( .A(n940), .B(n941), .Z(n939) );
  XOR U1711 ( .A(DB[781]), .B(DB[774]), .Z(n941) );
  AND U1712 ( .A(n70), .B(n942), .Z(n940) );
  XOR U1713 ( .A(n943), .B(n944), .Z(n942) );
  XOR U1714 ( .A(DB[774]), .B(DB[767]), .Z(n944) );
  AND U1715 ( .A(n74), .B(n945), .Z(n943) );
  XOR U1716 ( .A(n946), .B(n947), .Z(n945) );
  XOR U1717 ( .A(DB[767]), .B(DB[760]), .Z(n947) );
  AND U1718 ( .A(n78), .B(n948), .Z(n946) );
  XOR U1719 ( .A(n949), .B(n950), .Z(n948) );
  XOR U1720 ( .A(DB[760]), .B(DB[753]), .Z(n950) );
  AND U1721 ( .A(n82), .B(n951), .Z(n949) );
  XOR U1722 ( .A(n952), .B(n953), .Z(n951) );
  XOR U1723 ( .A(DB[753]), .B(DB[746]), .Z(n953) );
  AND U1724 ( .A(n86), .B(n954), .Z(n952) );
  XOR U1725 ( .A(n955), .B(n956), .Z(n954) );
  XOR U1726 ( .A(DB[746]), .B(DB[739]), .Z(n956) );
  AND U1727 ( .A(n90), .B(n957), .Z(n955) );
  XOR U1728 ( .A(n958), .B(n959), .Z(n957) );
  XOR U1729 ( .A(DB[739]), .B(DB[732]), .Z(n959) );
  AND U1730 ( .A(n94), .B(n960), .Z(n958) );
  XOR U1731 ( .A(n961), .B(n962), .Z(n960) );
  XOR U1732 ( .A(DB[732]), .B(DB[725]), .Z(n962) );
  AND U1733 ( .A(n98), .B(n963), .Z(n961) );
  XOR U1734 ( .A(n964), .B(n965), .Z(n963) );
  XOR U1735 ( .A(DB[725]), .B(DB[718]), .Z(n965) );
  AND U1736 ( .A(n102), .B(n966), .Z(n964) );
  XOR U1737 ( .A(n967), .B(n968), .Z(n966) );
  XOR U1738 ( .A(DB[718]), .B(DB[711]), .Z(n968) );
  AND U1739 ( .A(n106), .B(n969), .Z(n967) );
  XOR U1740 ( .A(n970), .B(n971), .Z(n969) );
  XOR U1741 ( .A(DB[711]), .B(DB[704]), .Z(n971) );
  AND U1742 ( .A(n110), .B(n972), .Z(n970) );
  XOR U1743 ( .A(n973), .B(n974), .Z(n972) );
  XOR U1744 ( .A(DB[704]), .B(DB[697]), .Z(n974) );
  AND U1745 ( .A(n114), .B(n975), .Z(n973) );
  XOR U1746 ( .A(n976), .B(n977), .Z(n975) );
  XOR U1747 ( .A(DB[697]), .B(DB[690]), .Z(n977) );
  AND U1748 ( .A(n118), .B(n978), .Z(n976) );
  XOR U1749 ( .A(n979), .B(n980), .Z(n978) );
  XOR U1750 ( .A(DB[690]), .B(DB[683]), .Z(n980) );
  AND U1751 ( .A(n122), .B(n981), .Z(n979) );
  XOR U1752 ( .A(n982), .B(n983), .Z(n981) );
  XOR U1753 ( .A(DB[683]), .B(DB[676]), .Z(n983) );
  AND U1754 ( .A(n126), .B(n984), .Z(n982) );
  XOR U1755 ( .A(n985), .B(n986), .Z(n984) );
  XOR U1756 ( .A(DB[676]), .B(DB[669]), .Z(n986) );
  AND U1757 ( .A(n130), .B(n987), .Z(n985) );
  XOR U1758 ( .A(n988), .B(n989), .Z(n987) );
  XOR U1759 ( .A(DB[669]), .B(DB[662]), .Z(n989) );
  AND U1760 ( .A(n134), .B(n990), .Z(n988) );
  XOR U1761 ( .A(n991), .B(n992), .Z(n990) );
  XOR U1762 ( .A(DB[662]), .B(DB[655]), .Z(n992) );
  AND U1763 ( .A(n138), .B(n993), .Z(n991) );
  XOR U1764 ( .A(n994), .B(n995), .Z(n993) );
  XOR U1765 ( .A(DB[655]), .B(DB[648]), .Z(n995) );
  AND U1766 ( .A(n142), .B(n996), .Z(n994) );
  XOR U1767 ( .A(n997), .B(n998), .Z(n996) );
  XOR U1768 ( .A(DB[648]), .B(DB[641]), .Z(n998) );
  AND U1769 ( .A(n146), .B(n999), .Z(n997) );
  XOR U1770 ( .A(n1000), .B(n1001), .Z(n999) );
  XOR U1771 ( .A(DB[641]), .B(DB[634]), .Z(n1001) );
  AND U1772 ( .A(n150), .B(n1002), .Z(n1000) );
  XOR U1773 ( .A(n1003), .B(n1004), .Z(n1002) );
  XOR U1774 ( .A(DB[634]), .B(DB[627]), .Z(n1004) );
  AND U1775 ( .A(n154), .B(n1005), .Z(n1003) );
  XOR U1776 ( .A(n1006), .B(n1007), .Z(n1005) );
  XOR U1777 ( .A(DB[627]), .B(DB[620]), .Z(n1007) );
  AND U1778 ( .A(n158), .B(n1008), .Z(n1006) );
  XOR U1779 ( .A(n1009), .B(n1010), .Z(n1008) );
  XOR U1780 ( .A(DB[620]), .B(DB[613]), .Z(n1010) );
  AND U1781 ( .A(n162), .B(n1011), .Z(n1009) );
  XOR U1782 ( .A(n1012), .B(n1013), .Z(n1011) );
  XOR U1783 ( .A(DB[613]), .B(DB[606]), .Z(n1013) );
  AND U1784 ( .A(n166), .B(n1014), .Z(n1012) );
  XOR U1785 ( .A(n1015), .B(n1016), .Z(n1014) );
  XOR U1786 ( .A(DB[606]), .B(DB[599]), .Z(n1016) );
  AND U1787 ( .A(n170), .B(n1017), .Z(n1015) );
  XOR U1788 ( .A(n1018), .B(n1019), .Z(n1017) );
  XOR U1789 ( .A(DB[599]), .B(DB[592]), .Z(n1019) );
  AND U1790 ( .A(n174), .B(n1020), .Z(n1018) );
  XOR U1791 ( .A(n1021), .B(n1022), .Z(n1020) );
  XOR U1792 ( .A(DB[592]), .B(DB[585]), .Z(n1022) );
  AND U1793 ( .A(n178), .B(n1023), .Z(n1021) );
  XOR U1794 ( .A(n1024), .B(n1025), .Z(n1023) );
  XOR U1795 ( .A(DB[585]), .B(DB[578]), .Z(n1025) );
  AND U1796 ( .A(n182), .B(n1026), .Z(n1024) );
  XOR U1797 ( .A(n1027), .B(n1028), .Z(n1026) );
  XOR U1798 ( .A(DB[578]), .B(DB[571]), .Z(n1028) );
  AND U1799 ( .A(n186), .B(n1029), .Z(n1027) );
  XOR U1800 ( .A(n1030), .B(n1031), .Z(n1029) );
  XOR U1801 ( .A(DB[571]), .B(DB[564]), .Z(n1031) );
  AND U1802 ( .A(n190), .B(n1032), .Z(n1030) );
  XOR U1803 ( .A(n1033), .B(n1034), .Z(n1032) );
  XOR U1804 ( .A(DB[564]), .B(DB[557]), .Z(n1034) );
  AND U1805 ( .A(n194), .B(n1035), .Z(n1033) );
  XOR U1806 ( .A(n1036), .B(n1037), .Z(n1035) );
  XOR U1807 ( .A(DB[557]), .B(DB[550]), .Z(n1037) );
  AND U1808 ( .A(n198), .B(n1038), .Z(n1036) );
  XOR U1809 ( .A(n1039), .B(n1040), .Z(n1038) );
  XOR U1810 ( .A(DB[550]), .B(DB[543]), .Z(n1040) );
  AND U1811 ( .A(n202), .B(n1041), .Z(n1039) );
  XOR U1812 ( .A(n1042), .B(n1043), .Z(n1041) );
  XOR U1813 ( .A(DB[543]), .B(DB[536]), .Z(n1043) );
  AND U1814 ( .A(n206), .B(n1044), .Z(n1042) );
  XOR U1815 ( .A(n1045), .B(n1046), .Z(n1044) );
  XOR U1816 ( .A(DB[536]), .B(DB[529]), .Z(n1046) );
  AND U1817 ( .A(n210), .B(n1047), .Z(n1045) );
  XOR U1818 ( .A(n1048), .B(n1049), .Z(n1047) );
  XOR U1819 ( .A(DB[529]), .B(DB[522]), .Z(n1049) );
  AND U1820 ( .A(n214), .B(n1050), .Z(n1048) );
  XOR U1821 ( .A(n1051), .B(n1052), .Z(n1050) );
  XOR U1822 ( .A(DB[522]), .B(DB[515]), .Z(n1052) );
  AND U1823 ( .A(n218), .B(n1053), .Z(n1051) );
  XOR U1824 ( .A(n1054), .B(n1055), .Z(n1053) );
  XOR U1825 ( .A(DB[515]), .B(DB[508]), .Z(n1055) );
  AND U1826 ( .A(n222), .B(n1056), .Z(n1054) );
  XOR U1827 ( .A(n1057), .B(n1058), .Z(n1056) );
  XOR U1828 ( .A(DB[508]), .B(DB[501]), .Z(n1058) );
  AND U1829 ( .A(n226), .B(n1059), .Z(n1057) );
  XOR U1830 ( .A(n1060), .B(n1061), .Z(n1059) );
  XOR U1831 ( .A(DB[501]), .B(DB[494]), .Z(n1061) );
  AND U1832 ( .A(n230), .B(n1062), .Z(n1060) );
  XOR U1833 ( .A(n1063), .B(n1064), .Z(n1062) );
  XOR U1834 ( .A(DB[494]), .B(DB[487]), .Z(n1064) );
  AND U1835 ( .A(n234), .B(n1065), .Z(n1063) );
  XOR U1836 ( .A(n1066), .B(n1067), .Z(n1065) );
  XOR U1837 ( .A(DB[487]), .B(DB[480]), .Z(n1067) );
  AND U1838 ( .A(n238), .B(n1068), .Z(n1066) );
  XOR U1839 ( .A(n1069), .B(n1070), .Z(n1068) );
  XOR U1840 ( .A(DB[480]), .B(DB[473]), .Z(n1070) );
  AND U1841 ( .A(n242), .B(n1071), .Z(n1069) );
  XOR U1842 ( .A(n1072), .B(n1073), .Z(n1071) );
  XOR U1843 ( .A(DB[473]), .B(DB[466]), .Z(n1073) );
  AND U1844 ( .A(n246), .B(n1074), .Z(n1072) );
  XOR U1845 ( .A(n1075), .B(n1076), .Z(n1074) );
  XOR U1846 ( .A(DB[466]), .B(DB[459]), .Z(n1076) );
  AND U1847 ( .A(n250), .B(n1077), .Z(n1075) );
  XOR U1848 ( .A(n1078), .B(n1079), .Z(n1077) );
  XOR U1849 ( .A(DB[459]), .B(DB[452]), .Z(n1079) );
  AND U1850 ( .A(n254), .B(n1080), .Z(n1078) );
  XOR U1851 ( .A(n1081), .B(n1082), .Z(n1080) );
  XOR U1852 ( .A(DB[452]), .B(DB[445]), .Z(n1082) );
  AND U1853 ( .A(n258), .B(n1083), .Z(n1081) );
  XOR U1854 ( .A(n1084), .B(n1085), .Z(n1083) );
  XOR U1855 ( .A(DB[445]), .B(DB[438]), .Z(n1085) );
  AND U1856 ( .A(n262), .B(n1086), .Z(n1084) );
  XOR U1857 ( .A(n1087), .B(n1088), .Z(n1086) );
  XOR U1858 ( .A(DB[438]), .B(DB[431]), .Z(n1088) );
  AND U1859 ( .A(n266), .B(n1089), .Z(n1087) );
  XOR U1860 ( .A(n1090), .B(n1091), .Z(n1089) );
  XOR U1861 ( .A(DB[431]), .B(DB[424]), .Z(n1091) );
  AND U1862 ( .A(n270), .B(n1092), .Z(n1090) );
  XOR U1863 ( .A(n1093), .B(n1094), .Z(n1092) );
  XOR U1864 ( .A(DB[424]), .B(DB[417]), .Z(n1094) );
  AND U1865 ( .A(n274), .B(n1095), .Z(n1093) );
  XOR U1866 ( .A(n1096), .B(n1097), .Z(n1095) );
  XOR U1867 ( .A(DB[417]), .B(DB[410]), .Z(n1097) );
  AND U1868 ( .A(n278), .B(n1098), .Z(n1096) );
  XOR U1869 ( .A(n1099), .B(n1100), .Z(n1098) );
  XOR U1870 ( .A(DB[410]), .B(DB[403]), .Z(n1100) );
  AND U1871 ( .A(n282), .B(n1101), .Z(n1099) );
  XOR U1872 ( .A(n1102), .B(n1103), .Z(n1101) );
  XOR U1873 ( .A(DB[403]), .B(DB[396]), .Z(n1103) );
  AND U1874 ( .A(n286), .B(n1104), .Z(n1102) );
  XOR U1875 ( .A(n1105), .B(n1106), .Z(n1104) );
  XOR U1876 ( .A(DB[396]), .B(DB[389]), .Z(n1106) );
  AND U1877 ( .A(n290), .B(n1107), .Z(n1105) );
  XOR U1878 ( .A(n1108), .B(n1109), .Z(n1107) );
  XOR U1879 ( .A(DB[389]), .B(DB[382]), .Z(n1109) );
  AND U1880 ( .A(n294), .B(n1110), .Z(n1108) );
  XOR U1881 ( .A(n1111), .B(n1112), .Z(n1110) );
  XOR U1882 ( .A(DB[382]), .B(DB[375]), .Z(n1112) );
  AND U1883 ( .A(n298), .B(n1113), .Z(n1111) );
  XOR U1884 ( .A(n1114), .B(n1115), .Z(n1113) );
  XOR U1885 ( .A(DB[375]), .B(DB[368]), .Z(n1115) );
  AND U1886 ( .A(n302), .B(n1116), .Z(n1114) );
  XOR U1887 ( .A(n1117), .B(n1118), .Z(n1116) );
  XOR U1888 ( .A(DB[368]), .B(DB[361]), .Z(n1118) );
  AND U1889 ( .A(n306), .B(n1119), .Z(n1117) );
  XOR U1890 ( .A(n1120), .B(n1121), .Z(n1119) );
  XOR U1891 ( .A(DB[361]), .B(DB[354]), .Z(n1121) );
  AND U1892 ( .A(n310), .B(n1122), .Z(n1120) );
  XOR U1893 ( .A(n1123), .B(n1124), .Z(n1122) );
  XOR U1894 ( .A(DB[354]), .B(DB[347]), .Z(n1124) );
  AND U1895 ( .A(n314), .B(n1125), .Z(n1123) );
  XOR U1896 ( .A(n1126), .B(n1127), .Z(n1125) );
  XOR U1897 ( .A(DB[347]), .B(DB[340]), .Z(n1127) );
  AND U1898 ( .A(n318), .B(n1128), .Z(n1126) );
  XOR U1899 ( .A(n1129), .B(n1130), .Z(n1128) );
  XOR U1900 ( .A(DB[340]), .B(DB[333]), .Z(n1130) );
  AND U1901 ( .A(n322), .B(n1131), .Z(n1129) );
  XOR U1902 ( .A(n1132), .B(n1133), .Z(n1131) );
  XOR U1903 ( .A(DB[333]), .B(DB[326]), .Z(n1133) );
  AND U1904 ( .A(n326), .B(n1134), .Z(n1132) );
  XOR U1905 ( .A(n1135), .B(n1136), .Z(n1134) );
  XOR U1906 ( .A(DB[326]), .B(DB[319]), .Z(n1136) );
  AND U1907 ( .A(n330), .B(n1137), .Z(n1135) );
  XOR U1908 ( .A(n1138), .B(n1139), .Z(n1137) );
  XOR U1909 ( .A(DB[319]), .B(DB[312]), .Z(n1139) );
  AND U1910 ( .A(n334), .B(n1140), .Z(n1138) );
  XOR U1911 ( .A(n1141), .B(n1142), .Z(n1140) );
  XOR U1912 ( .A(DB[312]), .B(DB[305]), .Z(n1142) );
  AND U1913 ( .A(n338), .B(n1143), .Z(n1141) );
  XOR U1914 ( .A(n1144), .B(n1145), .Z(n1143) );
  XOR U1915 ( .A(DB[305]), .B(DB[298]), .Z(n1145) );
  AND U1916 ( .A(n342), .B(n1146), .Z(n1144) );
  XOR U1917 ( .A(n1147), .B(n1148), .Z(n1146) );
  XOR U1918 ( .A(DB[298]), .B(DB[291]), .Z(n1148) );
  AND U1919 ( .A(n346), .B(n1149), .Z(n1147) );
  XOR U1920 ( .A(n1150), .B(n1151), .Z(n1149) );
  XOR U1921 ( .A(DB[291]), .B(DB[284]), .Z(n1151) );
  AND U1922 ( .A(n350), .B(n1152), .Z(n1150) );
  XOR U1923 ( .A(n1153), .B(n1154), .Z(n1152) );
  XOR U1924 ( .A(DB[284]), .B(DB[277]), .Z(n1154) );
  AND U1925 ( .A(n354), .B(n1155), .Z(n1153) );
  XOR U1926 ( .A(n1156), .B(n1157), .Z(n1155) );
  XOR U1927 ( .A(DB[277]), .B(DB[270]), .Z(n1157) );
  AND U1928 ( .A(n358), .B(n1158), .Z(n1156) );
  XOR U1929 ( .A(n1159), .B(n1160), .Z(n1158) );
  XOR U1930 ( .A(DB[270]), .B(DB[263]), .Z(n1160) );
  AND U1931 ( .A(n362), .B(n1161), .Z(n1159) );
  XOR U1932 ( .A(n1162), .B(n1163), .Z(n1161) );
  XOR U1933 ( .A(DB[263]), .B(DB[256]), .Z(n1163) );
  AND U1934 ( .A(n366), .B(n1164), .Z(n1162) );
  XOR U1935 ( .A(n1165), .B(n1166), .Z(n1164) );
  XOR U1936 ( .A(DB[256]), .B(DB[249]), .Z(n1166) );
  AND U1937 ( .A(n370), .B(n1167), .Z(n1165) );
  XOR U1938 ( .A(n1168), .B(n1169), .Z(n1167) );
  XOR U1939 ( .A(DB[249]), .B(DB[242]), .Z(n1169) );
  AND U1940 ( .A(n374), .B(n1170), .Z(n1168) );
  XOR U1941 ( .A(n1171), .B(n1172), .Z(n1170) );
  XOR U1942 ( .A(DB[242]), .B(DB[235]), .Z(n1172) );
  AND U1943 ( .A(n378), .B(n1173), .Z(n1171) );
  XOR U1944 ( .A(n1174), .B(n1175), .Z(n1173) );
  XOR U1945 ( .A(DB[235]), .B(DB[228]), .Z(n1175) );
  AND U1946 ( .A(n382), .B(n1176), .Z(n1174) );
  XOR U1947 ( .A(n1177), .B(n1178), .Z(n1176) );
  XOR U1948 ( .A(DB[228]), .B(DB[221]), .Z(n1178) );
  AND U1949 ( .A(n386), .B(n1179), .Z(n1177) );
  XOR U1950 ( .A(n1180), .B(n1181), .Z(n1179) );
  XOR U1951 ( .A(DB[221]), .B(DB[214]), .Z(n1181) );
  AND U1952 ( .A(n390), .B(n1182), .Z(n1180) );
  XOR U1953 ( .A(n1183), .B(n1184), .Z(n1182) );
  XOR U1954 ( .A(DB[214]), .B(DB[207]), .Z(n1184) );
  AND U1955 ( .A(n394), .B(n1185), .Z(n1183) );
  XOR U1956 ( .A(n1186), .B(n1187), .Z(n1185) );
  XOR U1957 ( .A(DB[207]), .B(DB[200]), .Z(n1187) );
  AND U1958 ( .A(n398), .B(n1188), .Z(n1186) );
  XOR U1959 ( .A(n1189), .B(n1190), .Z(n1188) );
  XOR U1960 ( .A(DB[200]), .B(DB[193]), .Z(n1190) );
  AND U1961 ( .A(n402), .B(n1191), .Z(n1189) );
  XOR U1962 ( .A(n1192), .B(n1193), .Z(n1191) );
  XOR U1963 ( .A(DB[193]), .B(DB[186]), .Z(n1193) );
  AND U1964 ( .A(n406), .B(n1194), .Z(n1192) );
  XOR U1965 ( .A(n1195), .B(n1196), .Z(n1194) );
  XOR U1966 ( .A(DB[186]), .B(DB[179]), .Z(n1196) );
  AND U1967 ( .A(n410), .B(n1197), .Z(n1195) );
  XOR U1968 ( .A(n1198), .B(n1199), .Z(n1197) );
  XOR U1969 ( .A(DB[179]), .B(DB[172]), .Z(n1199) );
  AND U1970 ( .A(n414), .B(n1200), .Z(n1198) );
  XOR U1971 ( .A(n1201), .B(n1202), .Z(n1200) );
  XOR U1972 ( .A(DB[172]), .B(DB[165]), .Z(n1202) );
  AND U1973 ( .A(n418), .B(n1203), .Z(n1201) );
  XOR U1974 ( .A(n1204), .B(n1205), .Z(n1203) );
  XOR U1975 ( .A(DB[165]), .B(DB[158]), .Z(n1205) );
  AND U1976 ( .A(n422), .B(n1206), .Z(n1204) );
  XOR U1977 ( .A(n1207), .B(n1208), .Z(n1206) );
  XOR U1978 ( .A(DB[158]), .B(DB[151]), .Z(n1208) );
  AND U1979 ( .A(n426), .B(n1209), .Z(n1207) );
  XOR U1980 ( .A(n1210), .B(n1211), .Z(n1209) );
  XOR U1981 ( .A(DB[151]), .B(DB[144]), .Z(n1211) );
  AND U1982 ( .A(n430), .B(n1212), .Z(n1210) );
  XOR U1983 ( .A(n1213), .B(n1214), .Z(n1212) );
  XOR U1984 ( .A(DB[144]), .B(DB[137]), .Z(n1214) );
  AND U1985 ( .A(n434), .B(n1215), .Z(n1213) );
  XOR U1986 ( .A(n1216), .B(n1217), .Z(n1215) );
  XOR U1987 ( .A(DB[137]), .B(DB[130]), .Z(n1217) );
  AND U1988 ( .A(n438), .B(n1218), .Z(n1216) );
  XOR U1989 ( .A(n1219), .B(n1220), .Z(n1218) );
  XOR U1990 ( .A(DB[130]), .B(DB[123]), .Z(n1220) );
  AND U1991 ( .A(n442), .B(n1221), .Z(n1219) );
  XOR U1992 ( .A(n1222), .B(n1223), .Z(n1221) );
  XOR U1993 ( .A(DB[123]), .B(DB[116]), .Z(n1223) );
  AND U1994 ( .A(n446), .B(n1224), .Z(n1222) );
  XOR U1995 ( .A(n1225), .B(n1226), .Z(n1224) );
  XOR U1996 ( .A(DB[116]), .B(DB[109]), .Z(n1226) );
  AND U1997 ( .A(n450), .B(n1227), .Z(n1225) );
  XOR U1998 ( .A(n1228), .B(n1229), .Z(n1227) );
  XOR U1999 ( .A(DB[109]), .B(DB[102]), .Z(n1229) );
  AND U2000 ( .A(n454), .B(n1230), .Z(n1228) );
  XOR U2001 ( .A(n1231), .B(n1232), .Z(n1230) );
  XOR U2002 ( .A(DB[95]), .B(DB[102]), .Z(n1232) );
  AND U2003 ( .A(n458), .B(n1233), .Z(n1231) );
  XOR U2004 ( .A(n1234), .B(n1235), .Z(n1233) );
  XOR U2005 ( .A(DB[95]), .B(DB[88]), .Z(n1235) );
  AND U2006 ( .A(n462), .B(n1236), .Z(n1234) );
  XOR U2007 ( .A(n1237), .B(n1238), .Z(n1236) );
  XOR U2008 ( .A(DB[88]), .B(DB[81]), .Z(n1238) );
  AND U2009 ( .A(n466), .B(n1239), .Z(n1237) );
  XOR U2010 ( .A(n1240), .B(n1241), .Z(n1239) );
  XOR U2011 ( .A(DB[81]), .B(DB[74]), .Z(n1241) );
  AND U2012 ( .A(n470), .B(n1242), .Z(n1240) );
  XOR U2013 ( .A(n1243), .B(n1244), .Z(n1242) );
  XOR U2014 ( .A(DB[74]), .B(DB[67]), .Z(n1244) );
  AND U2015 ( .A(n474), .B(n1245), .Z(n1243) );
  XOR U2016 ( .A(n1246), .B(n1247), .Z(n1245) );
  XOR U2017 ( .A(DB[67]), .B(DB[60]), .Z(n1247) );
  AND U2018 ( .A(n478), .B(n1248), .Z(n1246) );
  XOR U2019 ( .A(n1249), .B(n1250), .Z(n1248) );
  XOR U2020 ( .A(DB[60]), .B(DB[53]), .Z(n1250) );
  AND U2021 ( .A(n482), .B(n1251), .Z(n1249) );
  XOR U2022 ( .A(n1252), .B(n1253), .Z(n1251) );
  XOR U2023 ( .A(DB[53]), .B(DB[46]), .Z(n1253) );
  AND U2024 ( .A(n486), .B(n1254), .Z(n1252) );
  XOR U2025 ( .A(n1255), .B(n1256), .Z(n1254) );
  XOR U2026 ( .A(DB[46]), .B(DB[39]), .Z(n1256) );
  AND U2027 ( .A(n490), .B(n1257), .Z(n1255) );
  XOR U2028 ( .A(n1258), .B(n1259), .Z(n1257) );
  XOR U2029 ( .A(DB[39]), .B(DB[32]), .Z(n1259) );
  AND U2030 ( .A(n494), .B(n1260), .Z(n1258) );
  XOR U2031 ( .A(n1261), .B(n1262), .Z(n1260) );
  XOR U2032 ( .A(DB[32]), .B(DB[25]), .Z(n1262) );
  AND U2033 ( .A(n498), .B(n1263), .Z(n1261) );
  XOR U2034 ( .A(n1264), .B(n1265), .Z(n1263) );
  XOR U2035 ( .A(DB[25]), .B(DB[18]), .Z(n1265) );
  AND U2036 ( .A(n502), .B(n1266), .Z(n1264) );
  XOR U2037 ( .A(n1267), .B(n1268), .Z(n1266) );
  XOR U2038 ( .A(DB[18]), .B(DB[11]), .Z(n1268) );
  AND U2039 ( .A(n506), .B(n1269), .Z(n1267) );
  XOR U2040 ( .A(DB[4]), .B(DB[11]), .Z(n1269) );
  XOR U2041 ( .A(DB[892]), .B(n1270), .Z(min_val_out[3]) );
  AND U2042 ( .A(n2), .B(n1271), .Z(n1270) );
  XOR U2043 ( .A(n1272), .B(n1273), .Z(n1271) );
  XOR U2044 ( .A(n1274), .B(n1275), .Z(n1273) );
  IV U2045 ( .A(DB[892]), .Z(n1274) );
  AND U2046 ( .A(n6), .B(n1276), .Z(n1272) );
  XOR U2047 ( .A(n1277), .B(n1278), .Z(n1276) );
  XOR U2048 ( .A(DB[885]), .B(DB[878]), .Z(n1278) );
  AND U2049 ( .A(n10), .B(n1279), .Z(n1277) );
  XOR U2050 ( .A(n1280), .B(n1281), .Z(n1279) );
  XOR U2051 ( .A(DB[878]), .B(DB[871]), .Z(n1281) );
  AND U2052 ( .A(n14), .B(n1282), .Z(n1280) );
  XOR U2053 ( .A(n1283), .B(n1284), .Z(n1282) );
  XOR U2054 ( .A(DB[871]), .B(DB[864]), .Z(n1284) );
  AND U2055 ( .A(n18), .B(n1285), .Z(n1283) );
  XOR U2056 ( .A(n1286), .B(n1287), .Z(n1285) );
  XOR U2057 ( .A(DB[864]), .B(DB[857]), .Z(n1287) );
  AND U2058 ( .A(n22), .B(n1288), .Z(n1286) );
  XOR U2059 ( .A(n1289), .B(n1290), .Z(n1288) );
  XOR U2060 ( .A(DB[857]), .B(DB[850]), .Z(n1290) );
  AND U2061 ( .A(n26), .B(n1291), .Z(n1289) );
  XOR U2062 ( .A(n1292), .B(n1293), .Z(n1291) );
  XOR U2063 ( .A(DB[850]), .B(DB[843]), .Z(n1293) );
  AND U2064 ( .A(n30), .B(n1294), .Z(n1292) );
  XOR U2065 ( .A(n1295), .B(n1296), .Z(n1294) );
  XOR U2066 ( .A(DB[843]), .B(DB[836]), .Z(n1296) );
  AND U2067 ( .A(n34), .B(n1297), .Z(n1295) );
  XOR U2068 ( .A(n1298), .B(n1299), .Z(n1297) );
  XOR U2069 ( .A(DB[836]), .B(DB[829]), .Z(n1299) );
  AND U2070 ( .A(n38), .B(n1300), .Z(n1298) );
  XOR U2071 ( .A(n1301), .B(n1302), .Z(n1300) );
  XOR U2072 ( .A(DB[829]), .B(DB[822]), .Z(n1302) );
  AND U2073 ( .A(n42), .B(n1303), .Z(n1301) );
  XOR U2074 ( .A(n1304), .B(n1305), .Z(n1303) );
  XOR U2075 ( .A(DB[822]), .B(DB[815]), .Z(n1305) );
  AND U2076 ( .A(n46), .B(n1306), .Z(n1304) );
  XOR U2077 ( .A(n1307), .B(n1308), .Z(n1306) );
  XOR U2078 ( .A(DB[815]), .B(DB[808]), .Z(n1308) );
  AND U2079 ( .A(n50), .B(n1309), .Z(n1307) );
  XOR U2080 ( .A(n1310), .B(n1311), .Z(n1309) );
  XOR U2081 ( .A(DB[808]), .B(DB[801]), .Z(n1311) );
  AND U2082 ( .A(n54), .B(n1312), .Z(n1310) );
  XOR U2083 ( .A(n1313), .B(n1314), .Z(n1312) );
  XOR U2084 ( .A(DB[801]), .B(DB[794]), .Z(n1314) );
  AND U2085 ( .A(n58), .B(n1315), .Z(n1313) );
  XOR U2086 ( .A(n1316), .B(n1317), .Z(n1315) );
  XOR U2087 ( .A(DB[794]), .B(DB[787]), .Z(n1317) );
  AND U2088 ( .A(n62), .B(n1318), .Z(n1316) );
  XOR U2089 ( .A(n1319), .B(n1320), .Z(n1318) );
  XOR U2090 ( .A(DB[787]), .B(DB[780]), .Z(n1320) );
  AND U2091 ( .A(n66), .B(n1321), .Z(n1319) );
  XOR U2092 ( .A(n1322), .B(n1323), .Z(n1321) );
  XOR U2093 ( .A(DB[780]), .B(DB[773]), .Z(n1323) );
  AND U2094 ( .A(n70), .B(n1324), .Z(n1322) );
  XOR U2095 ( .A(n1325), .B(n1326), .Z(n1324) );
  XOR U2096 ( .A(DB[773]), .B(DB[766]), .Z(n1326) );
  AND U2097 ( .A(n74), .B(n1327), .Z(n1325) );
  XOR U2098 ( .A(n1328), .B(n1329), .Z(n1327) );
  XOR U2099 ( .A(DB[766]), .B(DB[759]), .Z(n1329) );
  AND U2100 ( .A(n78), .B(n1330), .Z(n1328) );
  XOR U2101 ( .A(n1331), .B(n1332), .Z(n1330) );
  XOR U2102 ( .A(DB[759]), .B(DB[752]), .Z(n1332) );
  AND U2103 ( .A(n82), .B(n1333), .Z(n1331) );
  XOR U2104 ( .A(n1334), .B(n1335), .Z(n1333) );
  XOR U2105 ( .A(DB[752]), .B(DB[745]), .Z(n1335) );
  AND U2106 ( .A(n86), .B(n1336), .Z(n1334) );
  XOR U2107 ( .A(n1337), .B(n1338), .Z(n1336) );
  XOR U2108 ( .A(DB[745]), .B(DB[738]), .Z(n1338) );
  AND U2109 ( .A(n90), .B(n1339), .Z(n1337) );
  XOR U2110 ( .A(n1340), .B(n1341), .Z(n1339) );
  XOR U2111 ( .A(DB[738]), .B(DB[731]), .Z(n1341) );
  AND U2112 ( .A(n94), .B(n1342), .Z(n1340) );
  XOR U2113 ( .A(n1343), .B(n1344), .Z(n1342) );
  XOR U2114 ( .A(DB[731]), .B(DB[724]), .Z(n1344) );
  AND U2115 ( .A(n98), .B(n1345), .Z(n1343) );
  XOR U2116 ( .A(n1346), .B(n1347), .Z(n1345) );
  XOR U2117 ( .A(DB[724]), .B(DB[717]), .Z(n1347) );
  AND U2118 ( .A(n102), .B(n1348), .Z(n1346) );
  XOR U2119 ( .A(n1349), .B(n1350), .Z(n1348) );
  XOR U2120 ( .A(DB[717]), .B(DB[710]), .Z(n1350) );
  AND U2121 ( .A(n106), .B(n1351), .Z(n1349) );
  XOR U2122 ( .A(n1352), .B(n1353), .Z(n1351) );
  XOR U2123 ( .A(DB[710]), .B(DB[703]), .Z(n1353) );
  AND U2124 ( .A(n110), .B(n1354), .Z(n1352) );
  XOR U2125 ( .A(n1355), .B(n1356), .Z(n1354) );
  XOR U2126 ( .A(DB[703]), .B(DB[696]), .Z(n1356) );
  AND U2127 ( .A(n114), .B(n1357), .Z(n1355) );
  XOR U2128 ( .A(n1358), .B(n1359), .Z(n1357) );
  XOR U2129 ( .A(DB[696]), .B(DB[689]), .Z(n1359) );
  AND U2130 ( .A(n118), .B(n1360), .Z(n1358) );
  XOR U2131 ( .A(n1361), .B(n1362), .Z(n1360) );
  XOR U2132 ( .A(DB[689]), .B(DB[682]), .Z(n1362) );
  AND U2133 ( .A(n122), .B(n1363), .Z(n1361) );
  XOR U2134 ( .A(n1364), .B(n1365), .Z(n1363) );
  XOR U2135 ( .A(DB[682]), .B(DB[675]), .Z(n1365) );
  AND U2136 ( .A(n126), .B(n1366), .Z(n1364) );
  XOR U2137 ( .A(n1367), .B(n1368), .Z(n1366) );
  XOR U2138 ( .A(DB[675]), .B(DB[668]), .Z(n1368) );
  AND U2139 ( .A(n130), .B(n1369), .Z(n1367) );
  XOR U2140 ( .A(n1370), .B(n1371), .Z(n1369) );
  XOR U2141 ( .A(DB[668]), .B(DB[661]), .Z(n1371) );
  AND U2142 ( .A(n134), .B(n1372), .Z(n1370) );
  XOR U2143 ( .A(n1373), .B(n1374), .Z(n1372) );
  XOR U2144 ( .A(DB[661]), .B(DB[654]), .Z(n1374) );
  AND U2145 ( .A(n138), .B(n1375), .Z(n1373) );
  XOR U2146 ( .A(n1376), .B(n1377), .Z(n1375) );
  XOR U2147 ( .A(DB[654]), .B(DB[647]), .Z(n1377) );
  AND U2148 ( .A(n142), .B(n1378), .Z(n1376) );
  XOR U2149 ( .A(n1379), .B(n1380), .Z(n1378) );
  XOR U2150 ( .A(DB[647]), .B(DB[640]), .Z(n1380) );
  AND U2151 ( .A(n146), .B(n1381), .Z(n1379) );
  XOR U2152 ( .A(n1382), .B(n1383), .Z(n1381) );
  XOR U2153 ( .A(DB[640]), .B(DB[633]), .Z(n1383) );
  AND U2154 ( .A(n150), .B(n1384), .Z(n1382) );
  XOR U2155 ( .A(n1385), .B(n1386), .Z(n1384) );
  XOR U2156 ( .A(DB[633]), .B(DB[626]), .Z(n1386) );
  AND U2157 ( .A(n154), .B(n1387), .Z(n1385) );
  XOR U2158 ( .A(n1388), .B(n1389), .Z(n1387) );
  XOR U2159 ( .A(DB[626]), .B(DB[619]), .Z(n1389) );
  AND U2160 ( .A(n158), .B(n1390), .Z(n1388) );
  XOR U2161 ( .A(n1391), .B(n1392), .Z(n1390) );
  XOR U2162 ( .A(DB[619]), .B(DB[612]), .Z(n1392) );
  AND U2163 ( .A(n162), .B(n1393), .Z(n1391) );
  XOR U2164 ( .A(n1394), .B(n1395), .Z(n1393) );
  XOR U2165 ( .A(DB[612]), .B(DB[605]), .Z(n1395) );
  AND U2166 ( .A(n166), .B(n1396), .Z(n1394) );
  XOR U2167 ( .A(n1397), .B(n1398), .Z(n1396) );
  XOR U2168 ( .A(DB[605]), .B(DB[598]), .Z(n1398) );
  AND U2169 ( .A(n170), .B(n1399), .Z(n1397) );
  XOR U2170 ( .A(n1400), .B(n1401), .Z(n1399) );
  XOR U2171 ( .A(DB[598]), .B(DB[591]), .Z(n1401) );
  AND U2172 ( .A(n174), .B(n1402), .Z(n1400) );
  XOR U2173 ( .A(n1403), .B(n1404), .Z(n1402) );
  XOR U2174 ( .A(DB[591]), .B(DB[584]), .Z(n1404) );
  AND U2175 ( .A(n178), .B(n1405), .Z(n1403) );
  XOR U2176 ( .A(n1406), .B(n1407), .Z(n1405) );
  XOR U2177 ( .A(DB[584]), .B(DB[577]), .Z(n1407) );
  AND U2178 ( .A(n182), .B(n1408), .Z(n1406) );
  XOR U2179 ( .A(n1409), .B(n1410), .Z(n1408) );
  XOR U2180 ( .A(DB[577]), .B(DB[570]), .Z(n1410) );
  AND U2181 ( .A(n186), .B(n1411), .Z(n1409) );
  XOR U2182 ( .A(n1412), .B(n1413), .Z(n1411) );
  XOR U2183 ( .A(DB[570]), .B(DB[563]), .Z(n1413) );
  AND U2184 ( .A(n190), .B(n1414), .Z(n1412) );
  XOR U2185 ( .A(n1415), .B(n1416), .Z(n1414) );
  XOR U2186 ( .A(DB[563]), .B(DB[556]), .Z(n1416) );
  AND U2187 ( .A(n194), .B(n1417), .Z(n1415) );
  XOR U2188 ( .A(n1418), .B(n1419), .Z(n1417) );
  XOR U2189 ( .A(DB[556]), .B(DB[549]), .Z(n1419) );
  AND U2190 ( .A(n198), .B(n1420), .Z(n1418) );
  XOR U2191 ( .A(n1421), .B(n1422), .Z(n1420) );
  XOR U2192 ( .A(DB[549]), .B(DB[542]), .Z(n1422) );
  AND U2193 ( .A(n202), .B(n1423), .Z(n1421) );
  XOR U2194 ( .A(n1424), .B(n1425), .Z(n1423) );
  XOR U2195 ( .A(DB[542]), .B(DB[535]), .Z(n1425) );
  AND U2196 ( .A(n206), .B(n1426), .Z(n1424) );
  XOR U2197 ( .A(n1427), .B(n1428), .Z(n1426) );
  XOR U2198 ( .A(DB[535]), .B(DB[528]), .Z(n1428) );
  AND U2199 ( .A(n210), .B(n1429), .Z(n1427) );
  XOR U2200 ( .A(n1430), .B(n1431), .Z(n1429) );
  XOR U2201 ( .A(DB[528]), .B(DB[521]), .Z(n1431) );
  AND U2202 ( .A(n214), .B(n1432), .Z(n1430) );
  XOR U2203 ( .A(n1433), .B(n1434), .Z(n1432) );
  XOR U2204 ( .A(DB[521]), .B(DB[514]), .Z(n1434) );
  AND U2205 ( .A(n218), .B(n1435), .Z(n1433) );
  XOR U2206 ( .A(n1436), .B(n1437), .Z(n1435) );
  XOR U2207 ( .A(DB[514]), .B(DB[507]), .Z(n1437) );
  AND U2208 ( .A(n222), .B(n1438), .Z(n1436) );
  XOR U2209 ( .A(n1439), .B(n1440), .Z(n1438) );
  XOR U2210 ( .A(DB[507]), .B(DB[500]), .Z(n1440) );
  AND U2211 ( .A(n226), .B(n1441), .Z(n1439) );
  XOR U2212 ( .A(n1442), .B(n1443), .Z(n1441) );
  XOR U2213 ( .A(DB[500]), .B(DB[493]), .Z(n1443) );
  AND U2214 ( .A(n230), .B(n1444), .Z(n1442) );
  XOR U2215 ( .A(n1445), .B(n1446), .Z(n1444) );
  XOR U2216 ( .A(DB[493]), .B(DB[486]), .Z(n1446) );
  AND U2217 ( .A(n234), .B(n1447), .Z(n1445) );
  XOR U2218 ( .A(n1448), .B(n1449), .Z(n1447) );
  XOR U2219 ( .A(DB[486]), .B(DB[479]), .Z(n1449) );
  AND U2220 ( .A(n238), .B(n1450), .Z(n1448) );
  XOR U2221 ( .A(n1451), .B(n1452), .Z(n1450) );
  XOR U2222 ( .A(DB[479]), .B(DB[472]), .Z(n1452) );
  AND U2223 ( .A(n242), .B(n1453), .Z(n1451) );
  XOR U2224 ( .A(n1454), .B(n1455), .Z(n1453) );
  XOR U2225 ( .A(DB[472]), .B(DB[465]), .Z(n1455) );
  AND U2226 ( .A(n246), .B(n1456), .Z(n1454) );
  XOR U2227 ( .A(n1457), .B(n1458), .Z(n1456) );
  XOR U2228 ( .A(DB[465]), .B(DB[458]), .Z(n1458) );
  AND U2229 ( .A(n250), .B(n1459), .Z(n1457) );
  XOR U2230 ( .A(n1460), .B(n1461), .Z(n1459) );
  XOR U2231 ( .A(DB[458]), .B(DB[451]), .Z(n1461) );
  AND U2232 ( .A(n254), .B(n1462), .Z(n1460) );
  XOR U2233 ( .A(n1463), .B(n1464), .Z(n1462) );
  XOR U2234 ( .A(DB[451]), .B(DB[444]), .Z(n1464) );
  AND U2235 ( .A(n258), .B(n1465), .Z(n1463) );
  XOR U2236 ( .A(n1466), .B(n1467), .Z(n1465) );
  XOR U2237 ( .A(DB[444]), .B(DB[437]), .Z(n1467) );
  AND U2238 ( .A(n262), .B(n1468), .Z(n1466) );
  XOR U2239 ( .A(n1469), .B(n1470), .Z(n1468) );
  XOR U2240 ( .A(DB[437]), .B(DB[430]), .Z(n1470) );
  AND U2241 ( .A(n266), .B(n1471), .Z(n1469) );
  XOR U2242 ( .A(n1472), .B(n1473), .Z(n1471) );
  XOR U2243 ( .A(DB[430]), .B(DB[423]), .Z(n1473) );
  AND U2244 ( .A(n270), .B(n1474), .Z(n1472) );
  XOR U2245 ( .A(n1475), .B(n1476), .Z(n1474) );
  XOR U2246 ( .A(DB[423]), .B(DB[416]), .Z(n1476) );
  AND U2247 ( .A(n274), .B(n1477), .Z(n1475) );
  XOR U2248 ( .A(n1478), .B(n1479), .Z(n1477) );
  XOR U2249 ( .A(DB[416]), .B(DB[409]), .Z(n1479) );
  AND U2250 ( .A(n278), .B(n1480), .Z(n1478) );
  XOR U2251 ( .A(n1481), .B(n1482), .Z(n1480) );
  XOR U2252 ( .A(DB[409]), .B(DB[402]), .Z(n1482) );
  AND U2253 ( .A(n282), .B(n1483), .Z(n1481) );
  XOR U2254 ( .A(n1484), .B(n1485), .Z(n1483) );
  XOR U2255 ( .A(DB[402]), .B(DB[395]), .Z(n1485) );
  AND U2256 ( .A(n286), .B(n1486), .Z(n1484) );
  XOR U2257 ( .A(n1487), .B(n1488), .Z(n1486) );
  XOR U2258 ( .A(DB[395]), .B(DB[388]), .Z(n1488) );
  AND U2259 ( .A(n290), .B(n1489), .Z(n1487) );
  XOR U2260 ( .A(n1490), .B(n1491), .Z(n1489) );
  XOR U2261 ( .A(DB[388]), .B(DB[381]), .Z(n1491) );
  AND U2262 ( .A(n294), .B(n1492), .Z(n1490) );
  XOR U2263 ( .A(n1493), .B(n1494), .Z(n1492) );
  XOR U2264 ( .A(DB[381]), .B(DB[374]), .Z(n1494) );
  AND U2265 ( .A(n298), .B(n1495), .Z(n1493) );
  XOR U2266 ( .A(n1496), .B(n1497), .Z(n1495) );
  XOR U2267 ( .A(DB[374]), .B(DB[367]), .Z(n1497) );
  AND U2268 ( .A(n302), .B(n1498), .Z(n1496) );
  XOR U2269 ( .A(n1499), .B(n1500), .Z(n1498) );
  XOR U2270 ( .A(DB[367]), .B(DB[360]), .Z(n1500) );
  AND U2271 ( .A(n306), .B(n1501), .Z(n1499) );
  XOR U2272 ( .A(n1502), .B(n1503), .Z(n1501) );
  XOR U2273 ( .A(DB[360]), .B(DB[353]), .Z(n1503) );
  AND U2274 ( .A(n310), .B(n1504), .Z(n1502) );
  XOR U2275 ( .A(n1505), .B(n1506), .Z(n1504) );
  XOR U2276 ( .A(DB[353]), .B(DB[346]), .Z(n1506) );
  AND U2277 ( .A(n314), .B(n1507), .Z(n1505) );
  XOR U2278 ( .A(n1508), .B(n1509), .Z(n1507) );
  XOR U2279 ( .A(DB[346]), .B(DB[339]), .Z(n1509) );
  AND U2280 ( .A(n318), .B(n1510), .Z(n1508) );
  XOR U2281 ( .A(n1511), .B(n1512), .Z(n1510) );
  XOR U2282 ( .A(DB[339]), .B(DB[332]), .Z(n1512) );
  AND U2283 ( .A(n322), .B(n1513), .Z(n1511) );
  XOR U2284 ( .A(n1514), .B(n1515), .Z(n1513) );
  XOR U2285 ( .A(DB[332]), .B(DB[325]), .Z(n1515) );
  AND U2286 ( .A(n326), .B(n1516), .Z(n1514) );
  XOR U2287 ( .A(n1517), .B(n1518), .Z(n1516) );
  XOR U2288 ( .A(DB[325]), .B(DB[318]), .Z(n1518) );
  AND U2289 ( .A(n330), .B(n1519), .Z(n1517) );
  XOR U2290 ( .A(n1520), .B(n1521), .Z(n1519) );
  XOR U2291 ( .A(DB[318]), .B(DB[311]), .Z(n1521) );
  AND U2292 ( .A(n334), .B(n1522), .Z(n1520) );
  XOR U2293 ( .A(n1523), .B(n1524), .Z(n1522) );
  XOR U2294 ( .A(DB[311]), .B(DB[304]), .Z(n1524) );
  AND U2295 ( .A(n338), .B(n1525), .Z(n1523) );
  XOR U2296 ( .A(n1526), .B(n1527), .Z(n1525) );
  XOR U2297 ( .A(DB[304]), .B(DB[297]), .Z(n1527) );
  AND U2298 ( .A(n342), .B(n1528), .Z(n1526) );
  XOR U2299 ( .A(n1529), .B(n1530), .Z(n1528) );
  XOR U2300 ( .A(DB[297]), .B(DB[290]), .Z(n1530) );
  AND U2301 ( .A(n346), .B(n1531), .Z(n1529) );
  XOR U2302 ( .A(n1532), .B(n1533), .Z(n1531) );
  XOR U2303 ( .A(DB[290]), .B(DB[283]), .Z(n1533) );
  AND U2304 ( .A(n350), .B(n1534), .Z(n1532) );
  XOR U2305 ( .A(n1535), .B(n1536), .Z(n1534) );
  XOR U2306 ( .A(DB[283]), .B(DB[276]), .Z(n1536) );
  AND U2307 ( .A(n354), .B(n1537), .Z(n1535) );
  XOR U2308 ( .A(n1538), .B(n1539), .Z(n1537) );
  XOR U2309 ( .A(DB[276]), .B(DB[269]), .Z(n1539) );
  AND U2310 ( .A(n358), .B(n1540), .Z(n1538) );
  XOR U2311 ( .A(n1541), .B(n1542), .Z(n1540) );
  XOR U2312 ( .A(DB[269]), .B(DB[262]), .Z(n1542) );
  AND U2313 ( .A(n362), .B(n1543), .Z(n1541) );
  XOR U2314 ( .A(n1544), .B(n1545), .Z(n1543) );
  XOR U2315 ( .A(DB[262]), .B(DB[255]), .Z(n1545) );
  AND U2316 ( .A(n366), .B(n1546), .Z(n1544) );
  XOR U2317 ( .A(n1547), .B(n1548), .Z(n1546) );
  XOR U2318 ( .A(DB[255]), .B(DB[248]), .Z(n1548) );
  AND U2319 ( .A(n370), .B(n1549), .Z(n1547) );
  XOR U2320 ( .A(n1550), .B(n1551), .Z(n1549) );
  XOR U2321 ( .A(DB[248]), .B(DB[241]), .Z(n1551) );
  AND U2322 ( .A(n374), .B(n1552), .Z(n1550) );
  XOR U2323 ( .A(n1553), .B(n1554), .Z(n1552) );
  XOR U2324 ( .A(DB[241]), .B(DB[234]), .Z(n1554) );
  AND U2325 ( .A(n378), .B(n1555), .Z(n1553) );
  XOR U2326 ( .A(n1556), .B(n1557), .Z(n1555) );
  XOR U2327 ( .A(DB[234]), .B(DB[227]), .Z(n1557) );
  AND U2328 ( .A(n382), .B(n1558), .Z(n1556) );
  XOR U2329 ( .A(n1559), .B(n1560), .Z(n1558) );
  XOR U2330 ( .A(DB[227]), .B(DB[220]), .Z(n1560) );
  AND U2331 ( .A(n386), .B(n1561), .Z(n1559) );
  XOR U2332 ( .A(n1562), .B(n1563), .Z(n1561) );
  XOR U2333 ( .A(DB[220]), .B(DB[213]), .Z(n1563) );
  AND U2334 ( .A(n390), .B(n1564), .Z(n1562) );
  XOR U2335 ( .A(n1565), .B(n1566), .Z(n1564) );
  XOR U2336 ( .A(DB[213]), .B(DB[206]), .Z(n1566) );
  AND U2337 ( .A(n394), .B(n1567), .Z(n1565) );
  XOR U2338 ( .A(n1568), .B(n1569), .Z(n1567) );
  XOR U2339 ( .A(DB[206]), .B(DB[199]), .Z(n1569) );
  AND U2340 ( .A(n398), .B(n1570), .Z(n1568) );
  XOR U2341 ( .A(n1571), .B(n1572), .Z(n1570) );
  XOR U2342 ( .A(DB[199]), .B(DB[192]), .Z(n1572) );
  AND U2343 ( .A(n402), .B(n1573), .Z(n1571) );
  XOR U2344 ( .A(n1574), .B(n1575), .Z(n1573) );
  XOR U2345 ( .A(DB[192]), .B(DB[185]), .Z(n1575) );
  AND U2346 ( .A(n406), .B(n1576), .Z(n1574) );
  XOR U2347 ( .A(n1577), .B(n1578), .Z(n1576) );
  XOR U2348 ( .A(DB[185]), .B(DB[178]), .Z(n1578) );
  AND U2349 ( .A(n410), .B(n1579), .Z(n1577) );
  XOR U2350 ( .A(n1580), .B(n1581), .Z(n1579) );
  XOR U2351 ( .A(DB[178]), .B(DB[171]), .Z(n1581) );
  AND U2352 ( .A(n414), .B(n1582), .Z(n1580) );
  XOR U2353 ( .A(n1583), .B(n1584), .Z(n1582) );
  XOR U2354 ( .A(DB[171]), .B(DB[164]), .Z(n1584) );
  AND U2355 ( .A(n418), .B(n1585), .Z(n1583) );
  XOR U2356 ( .A(n1586), .B(n1587), .Z(n1585) );
  XOR U2357 ( .A(DB[164]), .B(DB[157]), .Z(n1587) );
  AND U2358 ( .A(n422), .B(n1588), .Z(n1586) );
  XOR U2359 ( .A(n1589), .B(n1590), .Z(n1588) );
  XOR U2360 ( .A(DB[157]), .B(DB[150]), .Z(n1590) );
  AND U2361 ( .A(n426), .B(n1591), .Z(n1589) );
  XOR U2362 ( .A(n1592), .B(n1593), .Z(n1591) );
  XOR U2363 ( .A(DB[150]), .B(DB[143]), .Z(n1593) );
  AND U2364 ( .A(n430), .B(n1594), .Z(n1592) );
  XOR U2365 ( .A(n1595), .B(n1596), .Z(n1594) );
  XOR U2366 ( .A(DB[143]), .B(DB[136]), .Z(n1596) );
  AND U2367 ( .A(n434), .B(n1597), .Z(n1595) );
  XOR U2368 ( .A(n1598), .B(n1599), .Z(n1597) );
  XOR U2369 ( .A(DB[136]), .B(DB[129]), .Z(n1599) );
  AND U2370 ( .A(n438), .B(n1600), .Z(n1598) );
  XOR U2371 ( .A(n1601), .B(n1602), .Z(n1600) );
  XOR U2372 ( .A(DB[129]), .B(DB[122]), .Z(n1602) );
  AND U2373 ( .A(n442), .B(n1603), .Z(n1601) );
  XOR U2374 ( .A(n1604), .B(n1605), .Z(n1603) );
  XOR U2375 ( .A(DB[122]), .B(DB[115]), .Z(n1605) );
  AND U2376 ( .A(n446), .B(n1606), .Z(n1604) );
  XOR U2377 ( .A(n1607), .B(n1608), .Z(n1606) );
  XOR U2378 ( .A(DB[115]), .B(DB[108]), .Z(n1608) );
  AND U2379 ( .A(n450), .B(n1609), .Z(n1607) );
  XOR U2380 ( .A(n1610), .B(n1611), .Z(n1609) );
  XOR U2381 ( .A(DB[108]), .B(DB[101]), .Z(n1611) );
  AND U2382 ( .A(n454), .B(n1612), .Z(n1610) );
  XOR U2383 ( .A(n1613), .B(n1614), .Z(n1612) );
  XOR U2384 ( .A(DB[94]), .B(DB[101]), .Z(n1614) );
  AND U2385 ( .A(n458), .B(n1615), .Z(n1613) );
  XOR U2386 ( .A(n1616), .B(n1617), .Z(n1615) );
  XOR U2387 ( .A(DB[94]), .B(DB[87]), .Z(n1617) );
  AND U2388 ( .A(n462), .B(n1618), .Z(n1616) );
  XOR U2389 ( .A(n1619), .B(n1620), .Z(n1618) );
  XOR U2390 ( .A(DB[87]), .B(DB[80]), .Z(n1620) );
  AND U2391 ( .A(n466), .B(n1621), .Z(n1619) );
  XOR U2392 ( .A(n1622), .B(n1623), .Z(n1621) );
  XOR U2393 ( .A(DB[80]), .B(DB[73]), .Z(n1623) );
  AND U2394 ( .A(n470), .B(n1624), .Z(n1622) );
  XOR U2395 ( .A(n1625), .B(n1626), .Z(n1624) );
  XOR U2396 ( .A(DB[73]), .B(DB[66]), .Z(n1626) );
  AND U2397 ( .A(n474), .B(n1627), .Z(n1625) );
  XOR U2398 ( .A(n1628), .B(n1629), .Z(n1627) );
  XOR U2399 ( .A(DB[66]), .B(DB[59]), .Z(n1629) );
  AND U2400 ( .A(n478), .B(n1630), .Z(n1628) );
  XOR U2401 ( .A(n1631), .B(n1632), .Z(n1630) );
  XOR U2402 ( .A(DB[59]), .B(DB[52]), .Z(n1632) );
  AND U2403 ( .A(n482), .B(n1633), .Z(n1631) );
  XOR U2404 ( .A(n1634), .B(n1635), .Z(n1633) );
  XOR U2405 ( .A(DB[52]), .B(DB[45]), .Z(n1635) );
  AND U2406 ( .A(n486), .B(n1636), .Z(n1634) );
  XOR U2407 ( .A(n1637), .B(n1638), .Z(n1636) );
  XOR U2408 ( .A(DB[45]), .B(DB[38]), .Z(n1638) );
  AND U2409 ( .A(n490), .B(n1639), .Z(n1637) );
  XOR U2410 ( .A(n1640), .B(n1641), .Z(n1639) );
  XOR U2411 ( .A(DB[38]), .B(DB[31]), .Z(n1641) );
  AND U2412 ( .A(n494), .B(n1642), .Z(n1640) );
  XOR U2413 ( .A(n1643), .B(n1644), .Z(n1642) );
  XOR U2414 ( .A(DB[31]), .B(DB[24]), .Z(n1644) );
  AND U2415 ( .A(n498), .B(n1645), .Z(n1643) );
  XOR U2416 ( .A(n1646), .B(n1647), .Z(n1645) );
  XOR U2417 ( .A(DB[24]), .B(DB[17]), .Z(n1647) );
  AND U2418 ( .A(n502), .B(n1648), .Z(n1646) );
  XOR U2419 ( .A(n1649), .B(n1650), .Z(n1648) );
  XOR U2420 ( .A(DB[17]), .B(DB[10]), .Z(n1650) );
  AND U2421 ( .A(n506), .B(n1651), .Z(n1649) );
  XOR U2422 ( .A(DB[3]), .B(DB[10]), .Z(n1651) );
  XOR U2423 ( .A(DB[891]), .B(n1652), .Z(min_val_out[2]) );
  AND U2424 ( .A(n2), .B(n1653), .Z(n1652) );
  XOR U2425 ( .A(n1654), .B(n1655), .Z(n1653) );
  XOR U2426 ( .A(DB[891]), .B(DB[884]), .Z(n1655) );
  AND U2427 ( .A(n6), .B(n1656), .Z(n1654) );
  XOR U2428 ( .A(n1657), .B(n1658), .Z(n1656) );
  XOR U2429 ( .A(DB[884]), .B(DB[877]), .Z(n1658) );
  AND U2430 ( .A(n10), .B(n1659), .Z(n1657) );
  XOR U2431 ( .A(n1660), .B(n1661), .Z(n1659) );
  XOR U2432 ( .A(DB[877]), .B(DB[870]), .Z(n1661) );
  AND U2433 ( .A(n14), .B(n1662), .Z(n1660) );
  XOR U2434 ( .A(n1663), .B(n1664), .Z(n1662) );
  XOR U2435 ( .A(DB[870]), .B(DB[863]), .Z(n1664) );
  AND U2436 ( .A(n18), .B(n1665), .Z(n1663) );
  XOR U2437 ( .A(n1666), .B(n1667), .Z(n1665) );
  XOR U2438 ( .A(DB[863]), .B(DB[856]), .Z(n1667) );
  AND U2439 ( .A(n22), .B(n1668), .Z(n1666) );
  XOR U2440 ( .A(n1669), .B(n1670), .Z(n1668) );
  XOR U2441 ( .A(DB[856]), .B(DB[849]), .Z(n1670) );
  AND U2442 ( .A(n26), .B(n1671), .Z(n1669) );
  XOR U2443 ( .A(n1672), .B(n1673), .Z(n1671) );
  XOR U2444 ( .A(DB[849]), .B(DB[842]), .Z(n1673) );
  AND U2445 ( .A(n30), .B(n1674), .Z(n1672) );
  XOR U2446 ( .A(n1675), .B(n1676), .Z(n1674) );
  XOR U2447 ( .A(DB[842]), .B(DB[835]), .Z(n1676) );
  AND U2448 ( .A(n34), .B(n1677), .Z(n1675) );
  XOR U2449 ( .A(n1678), .B(n1679), .Z(n1677) );
  XOR U2450 ( .A(DB[835]), .B(DB[828]), .Z(n1679) );
  AND U2451 ( .A(n38), .B(n1680), .Z(n1678) );
  XOR U2452 ( .A(n1681), .B(n1682), .Z(n1680) );
  XOR U2453 ( .A(DB[828]), .B(DB[821]), .Z(n1682) );
  AND U2454 ( .A(n42), .B(n1683), .Z(n1681) );
  XOR U2455 ( .A(n1684), .B(n1685), .Z(n1683) );
  XOR U2456 ( .A(DB[821]), .B(DB[814]), .Z(n1685) );
  AND U2457 ( .A(n46), .B(n1686), .Z(n1684) );
  XOR U2458 ( .A(n1687), .B(n1688), .Z(n1686) );
  XOR U2459 ( .A(DB[814]), .B(DB[807]), .Z(n1688) );
  AND U2460 ( .A(n50), .B(n1689), .Z(n1687) );
  XOR U2461 ( .A(n1690), .B(n1691), .Z(n1689) );
  XOR U2462 ( .A(DB[807]), .B(DB[800]), .Z(n1691) );
  AND U2463 ( .A(n54), .B(n1692), .Z(n1690) );
  XOR U2464 ( .A(n1693), .B(n1694), .Z(n1692) );
  XOR U2465 ( .A(DB[800]), .B(DB[793]), .Z(n1694) );
  AND U2466 ( .A(n58), .B(n1695), .Z(n1693) );
  XOR U2467 ( .A(n1696), .B(n1697), .Z(n1695) );
  XOR U2468 ( .A(DB[793]), .B(DB[786]), .Z(n1697) );
  AND U2469 ( .A(n62), .B(n1698), .Z(n1696) );
  XOR U2470 ( .A(n1699), .B(n1700), .Z(n1698) );
  XOR U2471 ( .A(DB[786]), .B(DB[779]), .Z(n1700) );
  AND U2472 ( .A(n66), .B(n1701), .Z(n1699) );
  XOR U2473 ( .A(n1702), .B(n1703), .Z(n1701) );
  XOR U2474 ( .A(DB[779]), .B(DB[772]), .Z(n1703) );
  AND U2475 ( .A(n70), .B(n1704), .Z(n1702) );
  XOR U2476 ( .A(n1705), .B(n1706), .Z(n1704) );
  XOR U2477 ( .A(DB[772]), .B(DB[765]), .Z(n1706) );
  AND U2478 ( .A(n74), .B(n1707), .Z(n1705) );
  XOR U2479 ( .A(n1708), .B(n1709), .Z(n1707) );
  XOR U2480 ( .A(DB[765]), .B(DB[758]), .Z(n1709) );
  AND U2481 ( .A(n78), .B(n1710), .Z(n1708) );
  XOR U2482 ( .A(n1711), .B(n1712), .Z(n1710) );
  XOR U2483 ( .A(DB[758]), .B(DB[751]), .Z(n1712) );
  AND U2484 ( .A(n82), .B(n1713), .Z(n1711) );
  XOR U2485 ( .A(n1714), .B(n1715), .Z(n1713) );
  XOR U2486 ( .A(DB[751]), .B(DB[744]), .Z(n1715) );
  AND U2487 ( .A(n86), .B(n1716), .Z(n1714) );
  XOR U2488 ( .A(n1717), .B(n1718), .Z(n1716) );
  XOR U2489 ( .A(DB[744]), .B(DB[737]), .Z(n1718) );
  AND U2490 ( .A(n90), .B(n1719), .Z(n1717) );
  XOR U2491 ( .A(n1720), .B(n1721), .Z(n1719) );
  XOR U2492 ( .A(DB[737]), .B(DB[730]), .Z(n1721) );
  AND U2493 ( .A(n94), .B(n1722), .Z(n1720) );
  XOR U2494 ( .A(n1723), .B(n1724), .Z(n1722) );
  XOR U2495 ( .A(DB[730]), .B(DB[723]), .Z(n1724) );
  AND U2496 ( .A(n98), .B(n1725), .Z(n1723) );
  XOR U2497 ( .A(n1726), .B(n1727), .Z(n1725) );
  XOR U2498 ( .A(DB[723]), .B(DB[716]), .Z(n1727) );
  AND U2499 ( .A(n102), .B(n1728), .Z(n1726) );
  XOR U2500 ( .A(n1729), .B(n1730), .Z(n1728) );
  XOR U2501 ( .A(DB[716]), .B(DB[709]), .Z(n1730) );
  AND U2502 ( .A(n106), .B(n1731), .Z(n1729) );
  XOR U2503 ( .A(n1732), .B(n1733), .Z(n1731) );
  XOR U2504 ( .A(DB[709]), .B(DB[702]), .Z(n1733) );
  AND U2505 ( .A(n110), .B(n1734), .Z(n1732) );
  XOR U2506 ( .A(n1735), .B(n1736), .Z(n1734) );
  XOR U2507 ( .A(DB[702]), .B(DB[695]), .Z(n1736) );
  AND U2508 ( .A(n114), .B(n1737), .Z(n1735) );
  XOR U2509 ( .A(n1738), .B(n1739), .Z(n1737) );
  XOR U2510 ( .A(DB[695]), .B(DB[688]), .Z(n1739) );
  AND U2511 ( .A(n118), .B(n1740), .Z(n1738) );
  XOR U2512 ( .A(n1741), .B(n1742), .Z(n1740) );
  XOR U2513 ( .A(DB[688]), .B(DB[681]), .Z(n1742) );
  AND U2514 ( .A(n122), .B(n1743), .Z(n1741) );
  XOR U2515 ( .A(n1744), .B(n1745), .Z(n1743) );
  XOR U2516 ( .A(DB[681]), .B(DB[674]), .Z(n1745) );
  AND U2517 ( .A(n126), .B(n1746), .Z(n1744) );
  XOR U2518 ( .A(n1747), .B(n1748), .Z(n1746) );
  XOR U2519 ( .A(DB[674]), .B(DB[667]), .Z(n1748) );
  AND U2520 ( .A(n130), .B(n1749), .Z(n1747) );
  XOR U2521 ( .A(n1750), .B(n1751), .Z(n1749) );
  XOR U2522 ( .A(DB[667]), .B(DB[660]), .Z(n1751) );
  AND U2523 ( .A(n134), .B(n1752), .Z(n1750) );
  XOR U2524 ( .A(n1753), .B(n1754), .Z(n1752) );
  XOR U2525 ( .A(DB[660]), .B(DB[653]), .Z(n1754) );
  AND U2526 ( .A(n138), .B(n1755), .Z(n1753) );
  XOR U2527 ( .A(n1756), .B(n1757), .Z(n1755) );
  XOR U2528 ( .A(DB[653]), .B(DB[646]), .Z(n1757) );
  AND U2529 ( .A(n142), .B(n1758), .Z(n1756) );
  XOR U2530 ( .A(n1759), .B(n1760), .Z(n1758) );
  XOR U2531 ( .A(DB[646]), .B(DB[639]), .Z(n1760) );
  AND U2532 ( .A(n146), .B(n1761), .Z(n1759) );
  XOR U2533 ( .A(n1762), .B(n1763), .Z(n1761) );
  XOR U2534 ( .A(DB[639]), .B(DB[632]), .Z(n1763) );
  AND U2535 ( .A(n150), .B(n1764), .Z(n1762) );
  XOR U2536 ( .A(n1765), .B(n1766), .Z(n1764) );
  XOR U2537 ( .A(DB[632]), .B(DB[625]), .Z(n1766) );
  AND U2538 ( .A(n154), .B(n1767), .Z(n1765) );
  XOR U2539 ( .A(n1768), .B(n1769), .Z(n1767) );
  XOR U2540 ( .A(DB[625]), .B(DB[618]), .Z(n1769) );
  AND U2541 ( .A(n158), .B(n1770), .Z(n1768) );
  XOR U2542 ( .A(n1771), .B(n1772), .Z(n1770) );
  XOR U2543 ( .A(DB[618]), .B(DB[611]), .Z(n1772) );
  AND U2544 ( .A(n162), .B(n1773), .Z(n1771) );
  XOR U2545 ( .A(n1774), .B(n1775), .Z(n1773) );
  XOR U2546 ( .A(DB[611]), .B(DB[604]), .Z(n1775) );
  AND U2547 ( .A(n166), .B(n1776), .Z(n1774) );
  XOR U2548 ( .A(n1777), .B(n1778), .Z(n1776) );
  XOR U2549 ( .A(DB[604]), .B(DB[597]), .Z(n1778) );
  AND U2550 ( .A(n170), .B(n1779), .Z(n1777) );
  XOR U2551 ( .A(n1780), .B(n1781), .Z(n1779) );
  XOR U2552 ( .A(DB[597]), .B(DB[590]), .Z(n1781) );
  AND U2553 ( .A(n174), .B(n1782), .Z(n1780) );
  XOR U2554 ( .A(n1783), .B(n1784), .Z(n1782) );
  XOR U2555 ( .A(DB[590]), .B(DB[583]), .Z(n1784) );
  AND U2556 ( .A(n178), .B(n1785), .Z(n1783) );
  XOR U2557 ( .A(n1786), .B(n1787), .Z(n1785) );
  XOR U2558 ( .A(DB[583]), .B(DB[576]), .Z(n1787) );
  AND U2559 ( .A(n182), .B(n1788), .Z(n1786) );
  XOR U2560 ( .A(n1789), .B(n1790), .Z(n1788) );
  XOR U2561 ( .A(DB[576]), .B(DB[569]), .Z(n1790) );
  AND U2562 ( .A(n186), .B(n1791), .Z(n1789) );
  XOR U2563 ( .A(n1792), .B(n1793), .Z(n1791) );
  XOR U2564 ( .A(DB[569]), .B(DB[562]), .Z(n1793) );
  AND U2565 ( .A(n190), .B(n1794), .Z(n1792) );
  XOR U2566 ( .A(n1795), .B(n1796), .Z(n1794) );
  XOR U2567 ( .A(DB[562]), .B(DB[555]), .Z(n1796) );
  AND U2568 ( .A(n194), .B(n1797), .Z(n1795) );
  XOR U2569 ( .A(n1798), .B(n1799), .Z(n1797) );
  XOR U2570 ( .A(DB[555]), .B(DB[548]), .Z(n1799) );
  AND U2571 ( .A(n198), .B(n1800), .Z(n1798) );
  XOR U2572 ( .A(n1801), .B(n1802), .Z(n1800) );
  XOR U2573 ( .A(DB[548]), .B(DB[541]), .Z(n1802) );
  AND U2574 ( .A(n202), .B(n1803), .Z(n1801) );
  XOR U2575 ( .A(n1804), .B(n1805), .Z(n1803) );
  XOR U2576 ( .A(DB[541]), .B(DB[534]), .Z(n1805) );
  AND U2577 ( .A(n206), .B(n1806), .Z(n1804) );
  XOR U2578 ( .A(n1807), .B(n1808), .Z(n1806) );
  XOR U2579 ( .A(DB[534]), .B(DB[527]), .Z(n1808) );
  AND U2580 ( .A(n210), .B(n1809), .Z(n1807) );
  XOR U2581 ( .A(n1810), .B(n1811), .Z(n1809) );
  XOR U2582 ( .A(DB[527]), .B(DB[520]), .Z(n1811) );
  AND U2583 ( .A(n214), .B(n1812), .Z(n1810) );
  XOR U2584 ( .A(n1813), .B(n1814), .Z(n1812) );
  XOR U2585 ( .A(DB[520]), .B(DB[513]), .Z(n1814) );
  AND U2586 ( .A(n218), .B(n1815), .Z(n1813) );
  XOR U2587 ( .A(n1816), .B(n1817), .Z(n1815) );
  XOR U2588 ( .A(DB[513]), .B(DB[506]), .Z(n1817) );
  AND U2589 ( .A(n222), .B(n1818), .Z(n1816) );
  XOR U2590 ( .A(n1819), .B(n1820), .Z(n1818) );
  XOR U2591 ( .A(DB[506]), .B(DB[499]), .Z(n1820) );
  AND U2592 ( .A(n226), .B(n1821), .Z(n1819) );
  XOR U2593 ( .A(n1822), .B(n1823), .Z(n1821) );
  XOR U2594 ( .A(DB[499]), .B(DB[492]), .Z(n1823) );
  AND U2595 ( .A(n230), .B(n1824), .Z(n1822) );
  XOR U2596 ( .A(n1825), .B(n1826), .Z(n1824) );
  XOR U2597 ( .A(DB[492]), .B(DB[485]), .Z(n1826) );
  AND U2598 ( .A(n234), .B(n1827), .Z(n1825) );
  XOR U2599 ( .A(n1828), .B(n1829), .Z(n1827) );
  XOR U2600 ( .A(DB[485]), .B(DB[478]), .Z(n1829) );
  AND U2601 ( .A(n238), .B(n1830), .Z(n1828) );
  XOR U2602 ( .A(n1831), .B(n1832), .Z(n1830) );
  XOR U2603 ( .A(DB[478]), .B(DB[471]), .Z(n1832) );
  AND U2604 ( .A(n242), .B(n1833), .Z(n1831) );
  XOR U2605 ( .A(n1834), .B(n1835), .Z(n1833) );
  XOR U2606 ( .A(DB[471]), .B(DB[464]), .Z(n1835) );
  AND U2607 ( .A(n246), .B(n1836), .Z(n1834) );
  XOR U2608 ( .A(n1837), .B(n1838), .Z(n1836) );
  XOR U2609 ( .A(DB[464]), .B(DB[457]), .Z(n1838) );
  AND U2610 ( .A(n250), .B(n1839), .Z(n1837) );
  XOR U2611 ( .A(n1840), .B(n1841), .Z(n1839) );
  XOR U2612 ( .A(DB[457]), .B(DB[450]), .Z(n1841) );
  AND U2613 ( .A(n254), .B(n1842), .Z(n1840) );
  XOR U2614 ( .A(n1843), .B(n1844), .Z(n1842) );
  XOR U2615 ( .A(DB[450]), .B(DB[443]), .Z(n1844) );
  AND U2616 ( .A(n258), .B(n1845), .Z(n1843) );
  XOR U2617 ( .A(n1846), .B(n1847), .Z(n1845) );
  XOR U2618 ( .A(DB[443]), .B(DB[436]), .Z(n1847) );
  AND U2619 ( .A(n262), .B(n1848), .Z(n1846) );
  XOR U2620 ( .A(n1849), .B(n1850), .Z(n1848) );
  XOR U2621 ( .A(DB[436]), .B(DB[429]), .Z(n1850) );
  AND U2622 ( .A(n266), .B(n1851), .Z(n1849) );
  XOR U2623 ( .A(n1852), .B(n1853), .Z(n1851) );
  XOR U2624 ( .A(DB[429]), .B(DB[422]), .Z(n1853) );
  AND U2625 ( .A(n270), .B(n1854), .Z(n1852) );
  XOR U2626 ( .A(n1855), .B(n1856), .Z(n1854) );
  XOR U2627 ( .A(DB[422]), .B(DB[415]), .Z(n1856) );
  AND U2628 ( .A(n274), .B(n1857), .Z(n1855) );
  XOR U2629 ( .A(n1858), .B(n1859), .Z(n1857) );
  XOR U2630 ( .A(DB[415]), .B(DB[408]), .Z(n1859) );
  AND U2631 ( .A(n278), .B(n1860), .Z(n1858) );
  XOR U2632 ( .A(n1861), .B(n1862), .Z(n1860) );
  XOR U2633 ( .A(DB[408]), .B(DB[401]), .Z(n1862) );
  AND U2634 ( .A(n282), .B(n1863), .Z(n1861) );
  XOR U2635 ( .A(n1864), .B(n1865), .Z(n1863) );
  XOR U2636 ( .A(DB[401]), .B(DB[394]), .Z(n1865) );
  AND U2637 ( .A(n286), .B(n1866), .Z(n1864) );
  XOR U2638 ( .A(n1867), .B(n1868), .Z(n1866) );
  XOR U2639 ( .A(DB[394]), .B(DB[387]), .Z(n1868) );
  AND U2640 ( .A(n290), .B(n1869), .Z(n1867) );
  XOR U2641 ( .A(n1870), .B(n1871), .Z(n1869) );
  XOR U2642 ( .A(DB[387]), .B(DB[380]), .Z(n1871) );
  AND U2643 ( .A(n294), .B(n1872), .Z(n1870) );
  XOR U2644 ( .A(n1873), .B(n1874), .Z(n1872) );
  XOR U2645 ( .A(DB[380]), .B(DB[373]), .Z(n1874) );
  AND U2646 ( .A(n298), .B(n1875), .Z(n1873) );
  XOR U2647 ( .A(n1876), .B(n1877), .Z(n1875) );
  XOR U2648 ( .A(DB[373]), .B(DB[366]), .Z(n1877) );
  AND U2649 ( .A(n302), .B(n1878), .Z(n1876) );
  XOR U2650 ( .A(n1879), .B(n1880), .Z(n1878) );
  XOR U2651 ( .A(DB[366]), .B(DB[359]), .Z(n1880) );
  AND U2652 ( .A(n306), .B(n1881), .Z(n1879) );
  XOR U2653 ( .A(n1882), .B(n1883), .Z(n1881) );
  XOR U2654 ( .A(DB[359]), .B(DB[352]), .Z(n1883) );
  AND U2655 ( .A(n310), .B(n1884), .Z(n1882) );
  XOR U2656 ( .A(n1885), .B(n1886), .Z(n1884) );
  XOR U2657 ( .A(DB[352]), .B(DB[345]), .Z(n1886) );
  AND U2658 ( .A(n314), .B(n1887), .Z(n1885) );
  XOR U2659 ( .A(n1888), .B(n1889), .Z(n1887) );
  XOR U2660 ( .A(DB[345]), .B(DB[338]), .Z(n1889) );
  AND U2661 ( .A(n318), .B(n1890), .Z(n1888) );
  XOR U2662 ( .A(n1891), .B(n1892), .Z(n1890) );
  XOR U2663 ( .A(DB[338]), .B(DB[331]), .Z(n1892) );
  AND U2664 ( .A(n322), .B(n1893), .Z(n1891) );
  XOR U2665 ( .A(n1894), .B(n1895), .Z(n1893) );
  XOR U2666 ( .A(DB[331]), .B(DB[324]), .Z(n1895) );
  AND U2667 ( .A(n326), .B(n1896), .Z(n1894) );
  XOR U2668 ( .A(n1897), .B(n1898), .Z(n1896) );
  XOR U2669 ( .A(DB[324]), .B(DB[317]), .Z(n1898) );
  AND U2670 ( .A(n330), .B(n1899), .Z(n1897) );
  XOR U2671 ( .A(n1900), .B(n1901), .Z(n1899) );
  XOR U2672 ( .A(DB[317]), .B(DB[310]), .Z(n1901) );
  AND U2673 ( .A(n334), .B(n1902), .Z(n1900) );
  XOR U2674 ( .A(n1903), .B(n1904), .Z(n1902) );
  XOR U2675 ( .A(DB[310]), .B(DB[303]), .Z(n1904) );
  AND U2676 ( .A(n338), .B(n1905), .Z(n1903) );
  XOR U2677 ( .A(n1906), .B(n1907), .Z(n1905) );
  XOR U2678 ( .A(DB[303]), .B(DB[296]), .Z(n1907) );
  AND U2679 ( .A(n342), .B(n1908), .Z(n1906) );
  XOR U2680 ( .A(n1909), .B(n1910), .Z(n1908) );
  XOR U2681 ( .A(DB[296]), .B(DB[289]), .Z(n1910) );
  AND U2682 ( .A(n346), .B(n1911), .Z(n1909) );
  XOR U2683 ( .A(n1912), .B(n1913), .Z(n1911) );
  XOR U2684 ( .A(DB[289]), .B(DB[282]), .Z(n1913) );
  AND U2685 ( .A(n350), .B(n1914), .Z(n1912) );
  XOR U2686 ( .A(n1915), .B(n1916), .Z(n1914) );
  XOR U2687 ( .A(DB[282]), .B(DB[275]), .Z(n1916) );
  AND U2688 ( .A(n354), .B(n1917), .Z(n1915) );
  XOR U2689 ( .A(n1918), .B(n1919), .Z(n1917) );
  XOR U2690 ( .A(DB[275]), .B(DB[268]), .Z(n1919) );
  AND U2691 ( .A(n358), .B(n1920), .Z(n1918) );
  XOR U2692 ( .A(n1921), .B(n1922), .Z(n1920) );
  XOR U2693 ( .A(DB[268]), .B(DB[261]), .Z(n1922) );
  AND U2694 ( .A(n362), .B(n1923), .Z(n1921) );
  XOR U2695 ( .A(n1924), .B(n1925), .Z(n1923) );
  XOR U2696 ( .A(DB[261]), .B(DB[254]), .Z(n1925) );
  AND U2697 ( .A(n366), .B(n1926), .Z(n1924) );
  XOR U2698 ( .A(n1927), .B(n1928), .Z(n1926) );
  XOR U2699 ( .A(DB[254]), .B(DB[247]), .Z(n1928) );
  AND U2700 ( .A(n370), .B(n1929), .Z(n1927) );
  XOR U2701 ( .A(n1930), .B(n1931), .Z(n1929) );
  XOR U2702 ( .A(DB[247]), .B(DB[240]), .Z(n1931) );
  AND U2703 ( .A(n374), .B(n1932), .Z(n1930) );
  XOR U2704 ( .A(n1933), .B(n1934), .Z(n1932) );
  XOR U2705 ( .A(DB[240]), .B(DB[233]), .Z(n1934) );
  AND U2706 ( .A(n378), .B(n1935), .Z(n1933) );
  XOR U2707 ( .A(n1936), .B(n1937), .Z(n1935) );
  XOR U2708 ( .A(DB[233]), .B(DB[226]), .Z(n1937) );
  AND U2709 ( .A(n382), .B(n1938), .Z(n1936) );
  XOR U2710 ( .A(n1939), .B(n1940), .Z(n1938) );
  XOR U2711 ( .A(DB[226]), .B(DB[219]), .Z(n1940) );
  AND U2712 ( .A(n386), .B(n1941), .Z(n1939) );
  XOR U2713 ( .A(n1942), .B(n1943), .Z(n1941) );
  XOR U2714 ( .A(DB[219]), .B(DB[212]), .Z(n1943) );
  AND U2715 ( .A(n390), .B(n1944), .Z(n1942) );
  XOR U2716 ( .A(n1945), .B(n1946), .Z(n1944) );
  XOR U2717 ( .A(DB[212]), .B(DB[205]), .Z(n1946) );
  AND U2718 ( .A(n394), .B(n1947), .Z(n1945) );
  XOR U2719 ( .A(n1948), .B(n1949), .Z(n1947) );
  XOR U2720 ( .A(DB[205]), .B(DB[198]), .Z(n1949) );
  AND U2721 ( .A(n398), .B(n1950), .Z(n1948) );
  XOR U2722 ( .A(n1951), .B(n1952), .Z(n1950) );
  XOR U2723 ( .A(DB[198]), .B(DB[191]), .Z(n1952) );
  AND U2724 ( .A(n402), .B(n1953), .Z(n1951) );
  XOR U2725 ( .A(n1954), .B(n1955), .Z(n1953) );
  XOR U2726 ( .A(DB[191]), .B(DB[184]), .Z(n1955) );
  AND U2727 ( .A(n406), .B(n1956), .Z(n1954) );
  XOR U2728 ( .A(n1957), .B(n1958), .Z(n1956) );
  XOR U2729 ( .A(DB[184]), .B(DB[177]), .Z(n1958) );
  AND U2730 ( .A(n410), .B(n1959), .Z(n1957) );
  XOR U2731 ( .A(n1960), .B(n1961), .Z(n1959) );
  XOR U2732 ( .A(DB[177]), .B(DB[170]), .Z(n1961) );
  AND U2733 ( .A(n414), .B(n1962), .Z(n1960) );
  XOR U2734 ( .A(n1963), .B(n1964), .Z(n1962) );
  XOR U2735 ( .A(DB[170]), .B(DB[163]), .Z(n1964) );
  AND U2736 ( .A(n418), .B(n1965), .Z(n1963) );
  XOR U2737 ( .A(n1966), .B(n1967), .Z(n1965) );
  XOR U2738 ( .A(DB[163]), .B(DB[156]), .Z(n1967) );
  AND U2739 ( .A(n422), .B(n1968), .Z(n1966) );
  XOR U2740 ( .A(n1969), .B(n1970), .Z(n1968) );
  XOR U2741 ( .A(DB[156]), .B(DB[149]), .Z(n1970) );
  AND U2742 ( .A(n426), .B(n1971), .Z(n1969) );
  XOR U2743 ( .A(n1972), .B(n1973), .Z(n1971) );
  XOR U2744 ( .A(DB[149]), .B(DB[142]), .Z(n1973) );
  AND U2745 ( .A(n430), .B(n1974), .Z(n1972) );
  XOR U2746 ( .A(n1975), .B(n1976), .Z(n1974) );
  XOR U2747 ( .A(DB[142]), .B(DB[135]), .Z(n1976) );
  AND U2748 ( .A(n434), .B(n1977), .Z(n1975) );
  XOR U2749 ( .A(n1978), .B(n1979), .Z(n1977) );
  XOR U2750 ( .A(DB[135]), .B(DB[128]), .Z(n1979) );
  AND U2751 ( .A(n438), .B(n1980), .Z(n1978) );
  XOR U2752 ( .A(n1981), .B(n1982), .Z(n1980) );
  XOR U2753 ( .A(DB[128]), .B(DB[121]), .Z(n1982) );
  AND U2754 ( .A(n442), .B(n1983), .Z(n1981) );
  XOR U2755 ( .A(n1984), .B(n1985), .Z(n1983) );
  XOR U2756 ( .A(DB[121]), .B(DB[114]), .Z(n1985) );
  AND U2757 ( .A(n446), .B(n1986), .Z(n1984) );
  XOR U2758 ( .A(n1987), .B(n1988), .Z(n1986) );
  XOR U2759 ( .A(DB[114]), .B(DB[107]), .Z(n1988) );
  AND U2760 ( .A(n450), .B(n1989), .Z(n1987) );
  XOR U2761 ( .A(n1990), .B(n1991), .Z(n1989) );
  XOR U2762 ( .A(DB[107]), .B(DB[100]), .Z(n1991) );
  AND U2763 ( .A(n454), .B(n1992), .Z(n1990) );
  XOR U2764 ( .A(n1993), .B(n1994), .Z(n1992) );
  XOR U2765 ( .A(DB[93]), .B(DB[100]), .Z(n1994) );
  AND U2766 ( .A(n458), .B(n1995), .Z(n1993) );
  XOR U2767 ( .A(n1996), .B(n1997), .Z(n1995) );
  XOR U2768 ( .A(DB[93]), .B(DB[86]), .Z(n1997) );
  AND U2769 ( .A(n462), .B(n1998), .Z(n1996) );
  XOR U2770 ( .A(n1999), .B(n2000), .Z(n1998) );
  XOR U2771 ( .A(DB[86]), .B(DB[79]), .Z(n2000) );
  AND U2772 ( .A(n466), .B(n2001), .Z(n1999) );
  XOR U2773 ( .A(n2002), .B(n2003), .Z(n2001) );
  XOR U2774 ( .A(DB[79]), .B(DB[72]), .Z(n2003) );
  AND U2775 ( .A(n470), .B(n2004), .Z(n2002) );
  XOR U2776 ( .A(n2005), .B(n2006), .Z(n2004) );
  XOR U2777 ( .A(DB[72]), .B(DB[65]), .Z(n2006) );
  AND U2778 ( .A(n474), .B(n2007), .Z(n2005) );
  XOR U2779 ( .A(n2008), .B(n2009), .Z(n2007) );
  XOR U2780 ( .A(DB[65]), .B(DB[58]), .Z(n2009) );
  AND U2781 ( .A(n478), .B(n2010), .Z(n2008) );
  XOR U2782 ( .A(n2011), .B(n2012), .Z(n2010) );
  XOR U2783 ( .A(DB[58]), .B(DB[51]), .Z(n2012) );
  AND U2784 ( .A(n482), .B(n2013), .Z(n2011) );
  XOR U2785 ( .A(n2014), .B(n2015), .Z(n2013) );
  XOR U2786 ( .A(DB[51]), .B(DB[44]), .Z(n2015) );
  AND U2787 ( .A(n486), .B(n2016), .Z(n2014) );
  XOR U2788 ( .A(n2017), .B(n2018), .Z(n2016) );
  XOR U2789 ( .A(DB[44]), .B(DB[37]), .Z(n2018) );
  AND U2790 ( .A(n490), .B(n2019), .Z(n2017) );
  XOR U2791 ( .A(n2020), .B(n2021), .Z(n2019) );
  XOR U2792 ( .A(DB[37]), .B(DB[30]), .Z(n2021) );
  AND U2793 ( .A(n494), .B(n2022), .Z(n2020) );
  XOR U2794 ( .A(n2023), .B(n2024), .Z(n2022) );
  XOR U2795 ( .A(DB[30]), .B(DB[23]), .Z(n2024) );
  AND U2796 ( .A(n498), .B(n2025), .Z(n2023) );
  XOR U2797 ( .A(n2026), .B(n2027), .Z(n2025) );
  XOR U2798 ( .A(DB[23]), .B(DB[16]), .Z(n2027) );
  AND U2799 ( .A(n502), .B(n2028), .Z(n2026) );
  XOR U2800 ( .A(n2029), .B(n2030), .Z(n2028) );
  XOR U2801 ( .A(DB[9]), .B(DB[16]), .Z(n2030) );
  AND U2802 ( .A(n506), .B(n2031), .Z(n2029) );
  XOR U2803 ( .A(DB[9]), .B(DB[2]), .Z(n2031) );
  XOR U2804 ( .A(DB[890]), .B(n2032), .Z(min_val_out[1]) );
  AND U2805 ( .A(n2), .B(n2033), .Z(n2032) );
  XOR U2806 ( .A(n2034), .B(n2035), .Z(n2033) );
  XOR U2807 ( .A(DB[890]), .B(DB[883]), .Z(n2035) );
  AND U2808 ( .A(n6), .B(n2036), .Z(n2034) );
  XOR U2809 ( .A(n2037), .B(n2038), .Z(n2036) );
  XOR U2810 ( .A(DB[883]), .B(DB[876]), .Z(n2038) );
  AND U2811 ( .A(n10), .B(n2039), .Z(n2037) );
  XOR U2812 ( .A(n2040), .B(n2041), .Z(n2039) );
  XOR U2813 ( .A(DB[876]), .B(DB[869]), .Z(n2041) );
  AND U2814 ( .A(n14), .B(n2042), .Z(n2040) );
  XOR U2815 ( .A(n2043), .B(n2044), .Z(n2042) );
  XOR U2816 ( .A(DB[869]), .B(DB[862]), .Z(n2044) );
  AND U2817 ( .A(n18), .B(n2045), .Z(n2043) );
  XOR U2818 ( .A(n2046), .B(n2047), .Z(n2045) );
  XOR U2819 ( .A(DB[862]), .B(DB[855]), .Z(n2047) );
  AND U2820 ( .A(n22), .B(n2048), .Z(n2046) );
  XOR U2821 ( .A(n2049), .B(n2050), .Z(n2048) );
  XOR U2822 ( .A(DB[855]), .B(DB[848]), .Z(n2050) );
  AND U2823 ( .A(n26), .B(n2051), .Z(n2049) );
  XOR U2824 ( .A(n2052), .B(n2053), .Z(n2051) );
  XOR U2825 ( .A(DB[848]), .B(DB[841]), .Z(n2053) );
  AND U2826 ( .A(n30), .B(n2054), .Z(n2052) );
  XOR U2827 ( .A(n2055), .B(n2056), .Z(n2054) );
  XOR U2828 ( .A(DB[841]), .B(DB[834]), .Z(n2056) );
  AND U2829 ( .A(n34), .B(n2057), .Z(n2055) );
  XOR U2830 ( .A(n2058), .B(n2059), .Z(n2057) );
  XOR U2831 ( .A(DB[834]), .B(DB[827]), .Z(n2059) );
  AND U2832 ( .A(n38), .B(n2060), .Z(n2058) );
  XOR U2833 ( .A(n2061), .B(n2062), .Z(n2060) );
  XOR U2834 ( .A(DB[827]), .B(DB[820]), .Z(n2062) );
  AND U2835 ( .A(n42), .B(n2063), .Z(n2061) );
  XOR U2836 ( .A(n2064), .B(n2065), .Z(n2063) );
  XOR U2837 ( .A(DB[820]), .B(DB[813]), .Z(n2065) );
  AND U2838 ( .A(n46), .B(n2066), .Z(n2064) );
  XOR U2839 ( .A(n2067), .B(n2068), .Z(n2066) );
  XOR U2840 ( .A(DB[813]), .B(DB[806]), .Z(n2068) );
  AND U2841 ( .A(n50), .B(n2069), .Z(n2067) );
  XOR U2842 ( .A(n2070), .B(n2071), .Z(n2069) );
  XOR U2843 ( .A(DB[806]), .B(DB[799]), .Z(n2071) );
  AND U2844 ( .A(n54), .B(n2072), .Z(n2070) );
  XOR U2845 ( .A(n2073), .B(n2074), .Z(n2072) );
  XOR U2846 ( .A(DB[799]), .B(DB[792]), .Z(n2074) );
  AND U2847 ( .A(n58), .B(n2075), .Z(n2073) );
  XOR U2848 ( .A(n2076), .B(n2077), .Z(n2075) );
  XOR U2849 ( .A(DB[792]), .B(DB[785]), .Z(n2077) );
  AND U2850 ( .A(n62), .B(n2078), .Z(n2076) );
  XOR U2851 ( .A(n2079), .B(n2080), .Z(n2078) );
  XOR U2852 ( .A(DB[785]), .B(DB[778]), .Z(n2080) );
  AND U2853 ( .A(n66), .B(n2081), .Z(n2079) );
  XOR U2854 ( .A(n2082), .B(n2083), .Z(n2081) );
  XOR U2855 ( .A(DB[778]), .B(DB[771]), .Z(n2083) );
  AND U2856 ( .A(n70), .B(n2084), .Z(n2082) );
  XOR U2857 ( .A(n2085), .B(n2086), .Z(n2084) );
  XOR U2858 ( .A(DB[771]), .B(DB[764]), .Z(n2086) );
  AND U2859 ( .A(n74), .B(n2087), .Z(n2085) );
  XOR U2860 ( .A(n2088), .B(n2089), .Z(n2087) );
  XOR U2861 ( .A(DB[764]), .B(DB[757]), .Z(n2089) );
  AND U2862 ( .A(n78), .B(n2090), .Z(n2088) );
  XOR U2863 ( .A(n2091), .B(n2092), .Z(n2090) );
  XOR U2864 ( .A(DB[757]), .B(DB[750]), .Z(n2092) );
  AND U2865 ( .A(n82), .B(n2093), .Z(n2091) );
  XOR U2866 ( .A(n2094), .B(n2095), .Z(n2093) );
  XOR U2867 ( .A(DB[750]), .B(DB[743]), .Z(n2095) );
  AND U2868 ( .A(n86), .B(n2096), .Z(n2094) );
  XOR U2869 ( .A(n2097), .B(n2098), .Z(n2096) );
  XOR U2870 ( .A(DB[743]), .B(DB[736]), .Z(n2098) );
  AND U2871 ( .A(n90), .B(n2099), .Z(n2097) );
  XOR U2872 ( .A(n2100), .B(n2101), .Z(n2099) );
  XOR U2873 ( .A(DB[736]), .B(DB[729]), .Z(n2101) );
  AND U2874 ( .A(n94), .B(n2102), .Z(n2100) );
  XOR U2875 ( .A(n2103), .B(n2104), .Z(n2102) );
  XOR U2876 ( .A(DB[729]), .B(DB[722]), .Z(n2104) );
  AND U2877 ( .A(n98), .B(n2105), .Z(n2103) );
  XOR U2878 ( .A(n2106), .B(n2107), .Z(n2105) );
  XOR U2879 ( .A(DB[722]), .B(DB[715]), .Z(n2107) );
  AND U2880 ( .A(n102), .B(n2108), .Z(n2106) );
  XOR U2881 ( .A(n2109), .B(n2110), .Z(n2108) );
  XOR U2882 ( .A(DB[715]), .B(DB[708]), .Z(n2110) );
  AND U2883 ( .A(n106), .B(n2111), .Z(n2109) );
  XOR U2884 ( .A(n2112), .B(n2113), .Z(n2111) );
  XOR U2885 ( .A(DB[708]), .B(DB[701]), .Z(n2113) );
  AND U2886 ( .A(n110), .B(n2114), .Z(n2112) );
  XOR U2887 ( .A(n2115), .B(n2116), .Z(n2114) );
  XOR U2888 ( .A(DB[701]), .B(DB[694]), .Z(n2116) );
  AND U2889 ( .A(n114), .B(n2117), .Z(n2115) );
  XOR U2890 ( .A(n2118), .B(n2119), .Z(n2117) );
  XOR U2891 ( .A(DB[694]), .B(DB[687]), .Z(n2119) );
  AND U2892 ( .A(n118), .B(n2120), .Z(n2118) );
  XOR U2893 ( .A(n2121), .B(n2122), .Z(n2120) );
  XOR U2894 ( .A(DB[687]), .B(DB[680]), .Z(n2122) );
  AND U2895 ( .A(n122), .B(n2123), .Z(n2121) );
  XOR U2896 ( .A(n2124), .B(n2125), .Z(n2123) );
  XOR U2897 ( .A(DB[680]), .B(DB[673]), .Z(n2125) );
  AND U2898 ( .A(n126), .B(n2126), .Z(n2124) );
  XOR U2899 ( .A(n2127), .B(n2128), .Z(n2126) );
  XOR U2900 ( .A(DB[673]), .B(DB[666]), .Z(n2128) );
  AND U2901 ( .A(n130), .B(n2129), .Z(n2127) );
  XOR U2902 ( .A(n2130), .B(n2131), .Z(n2129) );
  XOR U2903 ( .A(DB[666]), .B(DB[659]), .Z(n2131) );
  AND U2904 ( .A(n134), .B(n2132), .Z(n2130) );
  XOR U2905 ( .A(n2133), .B(n2134), .Z(n2132) );
  XOR U2906 ( .A(DB[659]), .B(DB[652]), .Z(n2134) );
  AND U2907 ( .A(n138), .B(n2135), .Z(n2133) );
  XOR U2908 ( .A(n2136), .B(n2137), .Z(n2135) );
  XOR U2909 ( .A(DB[652]), .B(DB[645]), .Z(n2137) );
  AND U2910 ( .A(n142), .B(n2138), .Z(n2136) );
  XOR U2911 ( .A(n2139), .B(n2140), .Z(n2138) );
  XOR U2912 ( .A(DB[645]), .B(DB[638]), .Z(n2140) );
  AND U2913 ( .A(n146), .B(n2141), .Z(n2139) );
  XOR U2914 ( .A(n2142), .B(n2143), .Z(n2141) );
  XOR U2915 ( .A(DB[638]), .B(DB[631]), .Z(n2143) );
  AND U2916 ( .A(n150), .B(n2144), .Z(n2142) );
  XOR U2917 ( .A(n2145), .B(n2146), .Z(n2144) );
  XOR U2918 ( .A(DB[631]), .B(DB[624]), .Z(n2146) );
  AND U2919 ( .A(n154), .B(n2147), .Z(n2145) );
  XOR U2920 ( .A(n2148), .B(n2149), .Z(n2147) );
  XOR U2921 ( .A(DB[624]), .B(DB[617]), .Z(n2149) );
  AND U2922 ( .A(n158), .B(n2150), .Z(n2148) );
  XOR U2923 ( .A(n2151), .B(n2152), .Z(n2150) );
  XOR U2924 ( .A(DB[617]), .B(DB[610]), .Z(n2152) );
  AND U2925 ( .A(n162), .B(n2153), .Z(n2151) );
  XOR U2926 ( .A(n2154), .B(n2155), .Z(n2153) );
  XOR U2927 ( .A(DB[610]), .B(DB[603]), .Z(n2155) );
  AND U2928 ( .A(n166), .B(n2156), .Z(n2154) );
  XOR U2929 ( .A(n2157), .B(n2158), .Z(n2156) );
  XOR U2930 ( .A(DB[603]), .B(DB[596]), .Z(n2158) );
  AND U2931 ( .A(n170), .B(n2159), .Z(n2157) );
  XOR U2932 ( .A(n2160), .B(n2161), .Z(n2159) );
  XOR U2933 ( .A(DB[596]), .B(DB[589]), .Z(n2161) );
  AND U2934 ( .A(n174), .B(n2162), .Z(n2160) );
  XOR U2935 ( .A(n2163), .B(n2164), .Z(n2162) );
  XOR U2936 ( .A(DB[589]), .B(DB[582]), .Z(n2164) );
  AND U2937 ( .A(n178), .B(n2165), .Z(n2163) );
  XOR U2938 ( .A(n2166), .B(n2167), .Z(n2165) );
  XOR U2939 ( .A(DB[582]), .B(DB[575]), .Z(n2167) );
  AND U2940 ( .A(n182), .B(n2168), .Z(n2166) );
  XOR U2941 ( .A(n2169), .B(n2170), .Z(n2168) );
  XOR U2942 ( .A(DB[575]), .B(DB[568]), .Z(n2170) );
  AND U2943 ( .A(n186), .B(n2171), .Z(n2169) );
  XOR U2944 ( .A(n2172), .B(n2173), .Z(n2171) );
  XOR U2945 ( .A(DB[568]), .B(DB[561]), .Z(n2173) );
  AND U2946 ( .A(n190), .B(n2174), .Z(n2172) );
  XOR U2947 ( .A(n2175), .B(n2176), .Z(n2174) );
  XOR U2948 ( .A(DB[561]), .B(DB[554]), .Z(n2176) );
  AND U2949 ( .A(n194), .B(n2177), .Z(n2175) );
  XOR U2950 ( .A(n2178), .B(n2179), .Z(n2177) );
  XOR U2951 ( .A(DB[554]), .B(DB[547]), .Z(n2179) );
  AND U2952 ( .A(n198), .B(n2180), .Z(n2178) );
  XOR U2953 ( .A(n2181), .B(n2182), .Z(n2180) );
  XOR U2954 ( .A(DB[547]), .B(DB[540]), .Z(n2182) );
  AND U2955 ( .A(n202), .B(n2183), .Z(n2181) );
  XOR U2956 ( .A(n2184), .B(n2185), .Z(n2183) );
  XOR U2957 ( .A(DB[540]), .B(DB[533]), .Z(n2185) );
  AND U2958 ( .A(n206), .B(n2186), .Z(n2184) );
  XOR U2959 ( .A(n2187), .B(n2188), .Z(n2186) );
  XOR U2960 ( .A(DB[533]), .B(DB[526]), .Z(n2188) );
  AND U2961 ( .A(n210), .B(n2189), .Z(n2187) );
  XOR U2962 ( .A(n2190), .B(n2191), .Z(n2189) );
  XOR U2963 ( .A(DB[526]), .B(DB[519]), .Z(n2191) );
  AND U2964 ( .A(n214), .B(n2192), .Z(n2190) );
  XOR U2965 ( .A(n2193), .B(n2194), .Z(n2192) );
  XOR U2966 ( .A(DB[519]), .B(DB[512]), .Z(n2194) );
  AND U2967 ( .A(n218), .B(n2195), .Z(n2193) );
  XOR U2968 ( .A(n2196), .B(n2197), .Z(n2195) );
  XOR U2969 ( .A(DB[512]), .B(DB[505]), .Z(n2197) );
  AND U2970 ( .A(n222), .B(n2198), .Z(n2196) );
  XOR U2971 ( .A(n2199), .B(n2200), .Z(n2198) );
  XOR U2972 ( .A(DB[505]), .B(DB[498]), .Z(n2200) );
  AND U2973 ( .A(n226), .B(n2201), .Z(n2199) );
  XOR U2974 ( .A(n2202), .B(n2203), .Z(n2201) );
  XOR U2975 ( .A(DB[498]), .B(DB[491]), .Z(n2203) );
  AND U2976 ( .A(n230), .B(n2204), .Z(n2202) );
  XOR U2977 ( .A(n2205), .B(n2206), .Z(n2204) );
  XOR U2978 ( .A(DB[491]), .B(DB[484]), .Z(n2206) );
  AND U2979 ( .A(n234), .B(n2207), .Z(n2205) );
  XOR U2980 ( .A(n2208), .B(n2209), .Z(n2207) );
  XOR U2981 ( .A(DB[484]), .B(DB[477]), .Z(n2209) );
  AND U2982 ( .A(n238), .B(n2210), .Z(n2208) );
  XOR U2983 ( .A(n2211), .B(n2212), .Z(n2210) );
  XOR U2984 ( .A(DB[477]), .B(DB[470]), .Z(n2212) );
  AND U2985 ( .A(n242), .B(n2213), .Z(n2211) );
  XOR U2986 ( .A(n2214), .B(n2215), .Z(n2213) );
  XOR U2987 ( .A(DB[470]), .B(DB[463]), .Z(n2215) );
  AND U2988 ( .A(n246), .B(n2216), .Z(n2214) );
  XOR U2989 ( .A(n2217), .B(n2218), .Z(n2216) );
  XOR U2990 ( .A(DB[463]), .B(DB[456]), .Z(n2218) );
  AND U2991 ( .A(n250), .B(n2219), .Z(n2217) );
  XOR U2992 ( .A(n2220), .B(n2221), .Z(n2219) );
  XOR U2993 ( .A(DB[456]), .B(DB[449]), .Z(n2221) );
  AND U2994 ( .A(n254), .B(n2222), .Z(n2220) );
  XOR U2995 ( .A(n2223), .B(n2224), .Z(n2222) );
  XOR U2996 ( .A(DB[449]), .B(DB[442]), .Z(n2224) );
  AND U2997 ( .A(n258), .B(n2225), .Z(n2223) );
  XOR U2998 ( .A(n2226), .B(n2227), .Z(n2225) );
  XOR U2999 ( .A(DB[442]), .B(DB[435]), .Z(n2227) );
  AND U3000 ( .A(n262), .B(n2228), .Z(n2226) );
  XOR U3001 ( .A(n2229), .B(n2230), .Z(n2228) );
  XOR U3002 ( .A(DB[435]), .B(DB[428]), .Z(n2230) );
  AND U3003 ( .A(n266), .B(n2231), .Z(n2229) );
  XOR U3004 ( .A(n2232), .B(n2233), .Z(n2231) );
  XOR U3005 ( .A(DB[428]), .B(DB[421]), .Z(n2233) );
  AND U3006 ( .A(n270), .B(n2234), .Z(n2232) );
  XOR U3007 ( .A(n2235), .B(n2236), .Z(n2234) );
  XOR U3008 ( .A(DB[421]), .B(DB[414]), .Z(n2236) );
  AND U3009 ( .A(n274), .B(n2237), .Z(n2235) );
  XOR U3010 ( .A(n2238), .B(n2239), .Z(n2237) );
  XOR U3011 ( .A(DB[414]), .B(DB[407]), .Z(n2239) );
  AND U3012 ( .A(n278), .B(n2240), .Z(n2238) );
  XOR U3013 ( .A(n2241), .B(n2242), .Z(n2240) );
  XOR U3014 ( .A(DB[407]), .B(DB[400]), .Z(n2242) );
  AND U3015 ( .A(n282), .B(n2243), .Z(n2241) );
  XOR U3016 ( .A(n2244), .B(n2245), .Z(n2243) );
  XOR U3017 ( .A(DB[400]), .B(DB[393]), .Z(n2245) );
  AND U3018 ( .A(n286), .B(n2246), .Z(n2244) );
  XOR U3019 ( .A(n2247), .B(n2248), .Z(n2246) );
  XOR U3020 ( .A(DB[393]), .B(DB[386]), .Z(n2248) );
  AND U3021 ( .A(n290), .B(n2249), .Z(n2247) );
  XOR U3022 ( .A(n2250), .B(n2251), .Z(n2249) );
  XOR U3023 ( .A(DB[386]), .B(DB[379]), .Z(n2251) );
  AND U3024 ( .A(n294), .B(n2252), .Z(n2250) );
  XOR U3025 ( .A(n2253), .B(n2254), .Z(n2252) );
  XOR U3026 ( .A(DB[379]), .B(DB[372]), .Z(n2254) );
  AND U3027 ( .A(n298), .B(n2255), .Z(n2253) );
  XOR U3028 ( .A(n2256), .B(n2257), .Z(n2255) );
  XOR U3029 ( .A(DB[372]), .B(DB[365]), .Z(n2257) );
  AND U3030 ( .A(n302), .B(n2258), .Z(n2256) );
  XOR U3031 ( .A(n2259), .B(n2260), .Z(n2258) );
  XOR U3032 ( .A(DB[365]), .B(DB[358]), .Z(n2260) );
  AND U3033 ( .A(n306), .B(n2261), .Z(n2259) );
  XOR U3034 ( .A(n2262), .B(n2263), .Z(n2261) );
  XOR U3035 ( .A(DB[358]), .B(DB[351]), .Z(n2263) );
  AND U3036 ( .A(n310), .B(n2264), .Z(n2262) );
  XOR U3037 ( .A(n2265), .B(n2266), .Z(n2264) );
  XOR U3038 ( .A(DB[351]), .B(DB[344]), .Z(n2266) );
  AND U3039 ( .A(n314), .B(n2267), .Z(n2265) );
  XOR U3040 ( .A(n2268), .B(n2269), .Z(n2267) );
  XOR U3041 ( .A(DB[344]), .B(DB[337]), .Z(n2269) );
  AND U3042 ( .A(n318), .B(n2270), .Z(n2268) );
  XOR U3043 ( .A(n2271), .B(n2272), .Z(n2270) );
  XOR U3044 ( .A(DB[337]), .B(DB[330]), .Z(n2272) );
  AND U3045 ( .A(n322), .B(n2273), .Z(n2271) );
  XOR U3046 ( .A(n2274), .B(n2275), .Z(n2273) );
  XOR U3047 ( .A(DB[330]), .B(DB[323]), .Z(n2275) );
  AND U3048 ( .A(n326), .B(n2276), .Z(n2274) );
  XOR U3049 ( .A(n2277), .B(n2278), .Z(n2276) );
  XOR U3050 ( .A(DB[323]), .B(DB[316]), .Z(n2278) );
  AND U3051 ( .A(n330), .B(n2279), .Z(n2277) );
  XOR U3052 ( .A(n2280), .B(n2281), .Z(n2279) );
  XOR U3053 ( .A(DB[316]), .B(DB[309]), .Z(n2281) );
  AND U3054 ( .A(n334), .B(n2282), .Z(n2280) );
  XOR U3055 ( .A(n2283), .B(n2284), .Z(n2282) );
  XOR U3056 ( .A(DB[309]), .B(DB[302]), .Z(n2284) );
  AND U3057 ( .A(n338), .B(n2285), .Z(n2283) );
  XOR U3058 ( .A(n2286), .B(n2287), .Z(n2285) );
  XOR U3059 ( .A(DB[302]), .B(DB[295]), .Z(n2287) );
  AND U3060 ( .A(n342), .B(n2288), .Z(n2286) );
  XOR U3061 ( .A(n2289), .B(n2290), .Z(n2288) );
  XOR U3062 ( .A(DB[295]), .B(DB[288]), .Z(n2290) );
  AND U3063 ( .A(n346), .B(n2291), .Z(n2289) );
  XOR U3064 ( .A(n2292), .B(n2293), .Z(n2291) );
  XOR U3065 ( .A(DB[288]), .B(DB[281]), .Z(n2293) );
  AND U3066 ( .A(n350), .B(n2294), .Z(n2292) );
  XOR U3067 ( .A(n2295), .B(n2296), .Z(n2294) );
  XOR U3068 ( .A(DB[281]), .B(DB[274]), .Z(n2296) );
  AND U3069 ( .A(n354), .B(n2297), .Z(n2295) );
  XOR U3070 ( .A(n2298), .B(n2299), .Z(n2297) );
  XOR U3071 ( .A(DB[274]), .B(DB[267]), .Z(n2299) );
  AND U3072 ( .A(n358), .B(n2300), .Z(n2298) );
  XOR U3073 ( .A(n2301), .B(n2302), .Z(n2300) );
  XOR U3074 ( .A(DB[267]), .B(DB[260]), .Z(n2302) );
  AND U3075 ( .A(n362), .B(n2303), .Z(n2301) );
  XOR U3076 ( .A(n2304), .B(n2305), .Z(n2303) );
  XOR U3077 ( .A(DB[260]), .B(DB[253]), .Z(n2305) );
  AND U3078 ( .A(n366), .B(n2306), .Z(n2304) );
  XOR U3079 ( .A(n2307), .B(n2308), .Z(n2306) );
  XOR U3080 ( .A(DB[253]), .B(DB[246]), .Z(n2308) );
  AND U3081 ( .A(n370), .B(n2309), .Z(n2307) );
  XOR U3082 ( .A(n2310), .B(n2311), .Z(n2309) );
  XOR U3083 ( .A(DB[246]), .B(DB[239]), .Z(n2311) );
  AND U3084 ( .A(n374), .B(n2312), .Z(n2310) );
  XOR U3085 ( .A(n2313), .B(n2314), .Z(n2312) );
  XOR U3086 ( .A(DB[239]), .B(DB[232]), .Z(n2314) );
  AND U3087 ( .A(n378), .B(n2315), .Z(n2313) );
  XOR U3088 ( .A(n2316), .B(n2317), .Z(n2315) );
  XOR U3089 ( .A(DB[232]), .B(DB[225]), .Z(n2317) );
  AND U3090 ( .A(n382), .B(n2318), .Z(n2316) );
  XOR U3091 ( .A(n2319), .B(n2320), .Z(n2318) );
  XOR U3092 ( .A(DB[225]), .B(DB[218]), .Z(n2320) );
  AND U3093 ( .A(n386), .B(n2321), .Z(n2319) );
  XOR U3094 ( .A(n2322), .B(n2323), .Z(n2321) );
  XOR U3095 ( .A(DB[218]), .B(DB[211]), .Z(n2323) );
  AND U3096 ( .A(n390), .B(n2324), .Z(n2322) );
  XOR U3097 ( .A(n2325), .B(n2326), .Z(n2324) );
  XOR U3098 ( .A(DB[211]), .B(DB[204]), .Z(n2326) );
  AND U3099 ( .A(n394), .B(n2327), .Z(n2325) );
  XOR U3100 ( .A(n2328), .B(n2329), .Z(n2327) );
  XOR U3101 ( .A(DB[204]), .B(DB[197]), .Z(n2329) );
  AND U3102 ( .A(n398), .B(n2330), .Z(n2328) );
  XOR U3103 ( .A(n2331), .B(n2332), .Z(n2330) );
  XOR U3104 ( .A(DB[197]), .B(DB[190]), .Z(n2332) );
  AND U3105 ( .A(n402), .B(n2333), .Z(n2331) );
  XOR U3106 ( .A(n2334), .B(n2335), .Z(n2333) );
  XOR U3107 ( .A(DB[190]), .B(DB[183]), .Z(n2335) );
  AND U3108 ( .A(n406), .B(n2336), .Z(n2334) );
  XOR U3109 ( .A(n2337), .B(n2338), .Z(n2336) );
  XOR U3110 ( .A(DB[183]), .B(DB[176]), .Z(n2338) );
  AND U3111 ( .A(n410), .B(n2339), .Z(n2337) );
  XOR U3112 ( .A(n2340), .B(n2341), .Z(n2339) );
  XOR U3113 ( .A(DB[176]), .B(DB[169]), .Z(n2341) );
  AND U3114 ( .A(n414), .B(n2342), .Z(n2340) );
  XOR U3115 ( .A(n2343), .B(n2344), .Z(n2342) );
  XOR U3116 ( .A(DB[169]), .B(DB[162]), .Z(n2344) );
  AND U3117 ( .A(n418), .B(n2345), .Z(n2343) );
  XOR U3118 ( .A(n2346), .B(n2347), .Z(n2345) );
  XOR U3119 ( .A(DB[162]), .B(DB[155]), .Z(n2347) );
  AND U3120 ( .A(n422), .B(n2348), .Z(n2346) );
  XOR U3121 ( .A(n2349), .B(n2350), .Z(n2348) );
  XOR U3122 ( .A(DB[155]), .B(DB[148]), .Z(n2350) );
  AND U3123 ( .A(n426), .B(n2351), .Z(n2349) );
  XOR U3124 ( .A(n2352), .B(n2353), .Z(n2351) );
  XOR U3125 ( .A(DB[148]), .B(DB[141]), .Z(n2353) );
  AND U3126 ( .A(n430), .B(n2354), .Z(n2352) );
  XOR U3127 ( .A(n2355), .B(n2356), .Z(n2354) );
  XOR U3128 ( .A(DB[141]), .B(DB[134]), .Z(n2356) );
  AND U3129 ( .A(n434), .B(n2357), .Z(n2355) );
  XOR U3130 ( .A(n2358), .B(n2359), .Z(n2357) );
  XOR U3131 ( .A(DB[134]), .B(DB[127]), .Z(n2359) );
  AND U3132 ( .A(n438), .B(n2360), .Z(n2358) );
  XOR U3133 ( .A(n2361), .B(n2362), .Z(n2360) );
  XOR U3134 ( .A(DB[127]), .B(DB[120]), .Z(n2362) );
  AND U3135 ( .A(n442), .B(n2363), .Z(n2361) );
  XOR U3136 ( .A(n2364), .B(n2365), .Z(n2363) );
  XOR U3137 ( .A(DB[120]), .B(DB[113]), .Z(n2365) );
  AND U3138 ( .A(n446), .B(n2366), .Z(n2364) );
  XOR U3139 ( .A(n2367), .B(n2368), .Z(n2366) );
  XOR U3140 ( .A(DB[113]), .B(DB[106]), .Z(n2368) );
  AND U3141 ( .A(n450), .B(n2369), .Z(n2367) );
  XOR U3142 ( .A(n2370), .B(n2371), .Z(n2369) );
  XOR U3143 ( .A(DB[99]), .B(DB[106]), .Z(n2371) );
  AND U3144 ( .A(n454), .B(n2372), .Z(n2370) );
  XOR U3145 ( .A(n2373), .B(n2374), .Z(n2372) );
  XOR U3146 ( .A(DB[99]), .B(DB[92]), .Z(n2374) );
  AND U3147 ( .A(n458), .B(n2375), .Z(n2373) );
  XOR U3148 ( .A(n2376), .B(n2377), .Z(n2375) );
  XOR U3149 ( .A(DB[92]), .B(DB[85]), .Z(n2377) );
  AND U3150 ( .A(n462), .B(n2378), .Z(n2376) );
  XOR U3151 ( .A(n2379), .B(n2380), .Z(n2378) );
  XOR U3152 ( .A(DB[85]), .B(DB[78]), .Z(n2380) );
  AND U3153 ( .A(n466), .B(n2381), .Z(n2379) );
  XOR U3154 ( .A(n2382), .B(n2383), .Z(n2381) );
  XOR U3155 ( .A(DB[78]), .B(DB[71]), .Z(n2383) );
  AND U3156 ( .A(n470), .B(n2384), .Z(n2382) );
  XOR U3157 ( .A(n2385), .B(n2386), .Z(n2384) );
  XOR U3158 ( .A(DB[71]), .B(DB[64]), .Z(n2386) );
  AND U3159 ( .A(n474), .B(n2387), .Z(n2385) );
  XOR U3160 ( .A(n2388), .B(n2389), .Z(n2387) );
  XOR U3161 ( .A(DB[64]), .B(DB[57]), .Z(n2389) );
  AND U3162 ( .A(n478), .B(n2390), .Z(n2388) );
  XOR U3163 ( .A(n2391), .B(n2392), .Z(n2390) );
  XOR U3164 ( .A(DB[57]), .B(DB[50]), .Z(n2392) );
  AND U3165 ( .A(n482), .B(n2393), .Z(n2391) );
  XOR U3166 ( .A(n2394), .B(n2395), .Z(n2393) );
  XOR U3167 ( .A(DB[50]), .B(DB[43]), .Z(n2395) );
  AND U3168 ( .A(n486), .B(n2396), .Z(n2394) );
  XOR U3169 ( .A(n2397), .B(n2398), .Z(n2396) );
  XOR U3170 ( .A(DB[43]), .B(DB[36]), .Z(n2398) );
  AND U3171 ( .A(n490), .B(n2399), .Z(n2397) );
  XOR U3172 ( .A(n2400), .B(n2401), .Z(n2399) );
  XOR U3173 ( .A(DB[36]), .B(DB[29]), .Z(n2401) );
  AND U3174 ( .A(n494), .B(n2402), .Z(n2400) );
  XOR U3175 ( .A(n2403), .B(n2404), .Z(n2402) );
  XOR U3176 ( .A(DB[29]), .B(DB[22]), .Z(n2404) );
  AND U3177 ( .A(n498), .B(n2405), .Z(n2403) );
  XOR U3178 ( .A(n2406), .B(n2407), .Z(n2405) );
  XOR U3179 ( .A(DB[22]), .B(DB[15]), .Z(n2407) );
  AND U3180 ( .A(n502), .B(n2408), .Z(n2406) );
  XOR U3181 ( .A(n2409), .B(n2410), .Z(n2408) );
  XOR U3182 ( .A(DB[8]), .B(DB[15]), .Z(n2410) );
  AND U3183 ( .A(n506), .B(n2411), .Z(n2409) );
  XOR U3184 ( .A(DB[8]), .B(DB[1]), .Z(n2411) );
  XOR U3185 ( .A(DB[889]), .B(n2412), .Z(min_val_out[0]) );
  AND U3186 ( .A(n2), .B(n2413), .Z(n2412) );
  XOR U3187 ( .A(n2414), .B(n2415), .Z(n2413) );
  XOR U3188 ( .A(DB[889]), .B(DB[882]), .Z(n2415) );
  AND U3189 ( .A(n6), .B(n2416), .Z(n2414) );
  XOR U3190 ( .A(n2417), .B(n2418), .Z(n2416) );
  XOR U3191 ( .A(DB[882]), .B(DB[875]), .Z(n2418) );
  AND U3192 ( .A(n10), .B(n2419), .Z(n2417) );
  XOR U3193 ( .A(n2420), .B(n2421), .Z(n2419) );
  XOR U3194 ( .A(DB[875]), .B(DB[868]), .Z(n2421) );
  AND U3195 ( .A(n14), .B(n2422), .Z(n2420) );
  XOR U3196 ( .A(n2423), .B(n2424), .Z(n2422) );
  XOR U3197 ( .A(DB[868]), .B(DB[861]), .Z(n2424) );
  AND U3198 ( .A(n18), .B(n2425), .Z(n2423) );
  XOR U3199 ( .A(n2426), .B(n2427), .Z(n2425) );
  XOR U3200 ( .A(DB[861]), .B(DB[854]), .Z(n2427) );
  AND U3201 ( .A(n22), .B(n2428), .Z(n2426) );
  XOR U3202 ( .A(n2429), .B(n2430), .Z(n2428) );
  XOR U3203 ( .A(DB[854]), .B(DB[847]), .Z(n2430) );
  AND U3204 ( .A(n26), .B(n2431), .Z(n2429) );
  XOR U3205 ( .A(n2432), .B(n2433), .Z(n2431) );
  XOR U3206 ( .A(DB[847]), .B(DB[840]), .Z(n2433) );
  AND U3207 ( .A(n30), .B(n2434), .Z(n2432) );
  XOR U3208 ( .A(n2435), .B(n2436), .Z(n2434) );
  XOR U3209 ( .A(DB[840]), .B(DB[833]), .Z(n2436) );
  AND U3210 ( .A(n34), .B(n2437), .Z(n2435) );
  XOR U3211 ( .A(n2438), .B(n2439), .Z(n2437) );
  XOR U3212 ( .A(DB[833]), .B(DB[826]), .Z(n2439) );
  AND U3213 ( .A(n38), .B(n2440), .Z(n2438) );
  XOR U3214 ( .A(n2441), .B(n2442), .Z(n2440) );
  XOR U3215 ( .A(DB[826]), .B(DB[819]), .Z(n2442) );
  AND U3216 ( .A(n42), .B(n2443), .Z(n2441) );
  XOR U3217 ( .A(n2444), .B(n2445), .Z(n2443) );
  XOR U3218 ( .A(DB[819]), .B(DB[812]), .Z(n2445) );
  AND U3219 ( .A(n46), .B(n2446), .Z(n2444) );
  XOR U3220 ( .A(n2447), .B(n2448), .Z(n2446) );
  XOR U3221 ( .A(DB[812]), .B(DB[805]), .Z(n2448) );
  AND U3222 ( .A(n50), .B(n2449), .Z(n2447) );
  XOR U3223 ( .A(n2450), .B(n2451), .Z(n2449) );
  XOR U3224 ( .A(DB[805]), .B(DB[798]), .Z(n2451) );
  AND U3225 ( .A(n54), .B(n2452), .Z(n2450) );
  XOR U3226 ( .A(n2453), .B(n2454), .Z(n2452) );
  XOR U3227 ( .A(DB[798]), .B(DB[791]), .Z(n2454) );
  AND U3228 ( .A(n58), .B(n2455), .Z(n2453) );
  XOR U3229 ( .A(n2456), .B(n2457), .Z(n2455) );
  XOR U3230 ( .A(DB[791]), .B(DB[784]), .Z(n2457) );
  AND U3231 ( .A(n62), .B(n2458), .Z(n2456) );
  XOR U3232 ( .A(n2459), .B(n2460), .Z(n2458) );
  XOR U3233 ( .A(DB[784]), .B(DB[777]), .Z(n2460) );
  AND U3234 ( .A(n66), .B(n2461), .Z(n2459) );
  XOR U3235 ( .A(n2462), .B(n2463), .Z(n2461) );
  XOR U3236 ( .A(DB[777]), .B(DB[770]), .Z(n2463) );
  AND U3237 ( .A(n70), .B(n2464), .Z(n2462) );
  XOR U3238 ( .A(n2465), .B(n2466), .Z(n2464) );
  XOR U3239 ( .A(DB[770]), .B(DB[763]), .Z(n2466) );
  AND U3240 ( .A(n74), .B(n2467), .Z(n2465) );
  XOR U3241 ( .A(n2468), .B(n2469), .Z(n2467) );
  XOR U3242 ( .A(DB[763]), .B(DB[756]), .Z(n2469) );
  AND U3243 ( .A(n78), .B(n2470), .Z(n2468) );
  XOR U3244 ( .A(n2471), .B(n2472), .Z(n2470) );
  XOR U3245 ( .A(DB[756]), .B(DB[749]), .Z(n2472) );
  AND U3246 ( .A(n82), .B(n2473), .Z(n2471) );
  XOR U3247 ( .A(n2474), .B(n2475), .Z(n2473) );
  XOR U3248 ( .A(DB[749]), .B(DB[742]), .Z(n2475) );
  AND U3249 ( .A(n86), .B(n2476), .Z(n2474) );
  XOR U3250 ( .A(n2477), .B(n2478), .Z(n2476) );
  XOR U3251 ( .A(DB[742]), .B(DB[735]), .Z(n2478) );
  AND U3252 ( .A(n90), .B(n2479), .Z(n2477) );
  XOR U3253 ( .A(n2480), .B(n2481), .Z(n2479) );
  XOR U3254 ( .A(DB[735]), .B(DB[728]), .Z(n2481) );
  AND U3255 ( .A(n94), .B(n2482), .Z(n2480) );
  XOR U3256 ( .A(n2483), .B(n2484), .Z(n2482) );
  XOR U3257 ( .A(DB[728]), .B(DB[721]), .Z(n2484) );
  AND U3258 ( .A(n98), .B(n2485), .Z(n2483) );
  XOR U3259 ( .A(n2486), .B(n2487), .Z(n2485) );
  XOR U3260 ( .A(DB[721]), .B(DB[714]), .Z(n2487) );
  AND U3261 ( .A(n102), .B(n2488), .Z(n2486) );
  XOR U3262 ( .A(n2489), .B(n2490), .Z(n2488) );
  XOR U3263 ( .A(DB[714]), .B(DB[707]), .Z(n2490) );
  AND U3264 ( .A(n106), .B(n2491), .Z(n2489) );
  XOR U3265 ( .A(n2492), .B(n2493), .Z(n2491) );
  XOR U3266 ( .A(DB[707]), .B(DB[700]), .Z(n2493) );
  AND U3267 ( .A(n110), .B(n2494), .Z(n2492) );
  XOR U3268 ( .A(n2495), .B(n2496), .Z(n2494) );
  XOR U3269 ( .A(DB[700]), .B(DB[693]), .Z(n2496) );
  AND U3270 ( .A(n114), .B(n2497), .Z(n2495) );
  XOR U3271 ( .A(n2498), .B(n2499), .Z(n2497) );
  XOR U3272 ( .A(DB[693]), .B(DB[686]), .Z(n2499) );
  AND U3273 ( .A(n118), .B(n2500), .Z(n2498) );
  XOR U3274 ( .A(n2501), .B(n2502), .Z(n2500) );
  XOR U3275 ( .A(DB[686]), .B(DB[679]), .Z(n2502) );
  AND U3276 ( .A(n122), .B(n2503), .Z(n2501) );
  XOR U3277 ( .A(n2504), .B(n2505), .Z(n2503) );
  XOR U3278 ( .A(DB[679]), .B(DB[672]), .Z(n2505) );
  AND U3279 ( .A(n126), .B(n2506), .Z(n2504) );
  XOR U3280 ( .A(n2507), .B(n2508), .Z(n2506) );
  XOR U3281 ( .A(DB[672]), .B(DB[665]), .Z(n2508) );
  AND U3282 ( .A(n130), .B(n2509), .Z(n2507) );
  XOR U3283 ( .A(n2510), .B(n2511), .Z(n2509) );
  XOR U3284 ( .A(DB[665]), .B(DB[658]), .Z(n2511) );
  AND U3285 ( .A(n134), .B(n2512), .Z(n2510) );
  XOR U3286 ( .A(n2513), .B(n2514), .Z(n2512) );
  XOR U3287 ( .A(DB[658]), .B(DB[651]), .Z(n2514) );
  AND U3288 ( .A(n138), .B(n2515), .Z(n2513) );
  XOR U3289 ( .A(n2516), .B(n2517), .Z(n2515) );
  XOR U3290 ( .A(DB[651]), .B(DB[644]), .Z(n2517) );
  AND U3291 ( .A(n142), .B(n2518), .Z(n2516) );
  XOR U3292 ( .A(n2519), .B(n2520), .Z(n2518) );
  XOR U3293 ( .A(DB[644]), .B(DB[637]), .Z(n2520) );
  AND U3294 ( .A(n146), .B(n2521), .Z(n2519) );
  XOR U3295 ( .A(n2522), .B(n2523), .Z(n2521) );
  XOR U3296 ( .A(DB[637]), .B(DB[630]), .Z(n2523) );
  AND U3297 ( .A(n150), .B(n2524), .Z(n2522) );
  XOR U3298 ( .A(n2525), .B(n2526), .Z(n2524) );
  XOR U3299 ( .A(DB[630]), .B(DB[623]), .Z(n2526) );
  AND U3300 ( .A(n154), .B(n2527), .Z(n2525) );
  XOR U3301 ( .A(n2528), .B(n2529), .Z(n2527) );
  XOR U3302 ( .A(DB[623]), .B(DB[616]), .Z(n2529) );
  AND U3303 ( .A(n158), .B(n2530), .Z(n2528) );
  XOR U3304 ( .A(n2531), .B(n2532), .Z(n2530) );
  XOR U3305 ( .A(DB[616]), .B(DB[609]), .Z(n2532) );
  AND U3306 ( .A(n162), .B(n2533), .Z(n2531) );
  XOR U3307 ( .A(n2534), .B(n2535), .Z(n2533) );
  XOR U3308 ( .A(DB[609]), .B(DB[602]), .Z(n2535) );
  AND U3309 ( .A(n166), .B(n2536), .Z(n2534) );
  XOR U3310 ( .A(n2537), .B(n2538), .Z(n2536) );
  XOR U3311 ( .A(DB[602]), .B(DB[595]), .Z(n2538) );
  AND U3312 ( .A(n170), .B(n2539), .Z(n2537) );
  XOR U3313 ( .A(n2540), .B(n2541), .Z(n2539) );
  XOR U3314 ( .A(DB[595]), .B(DB[588]), .Z(n2541) );
  AND U3315 ( .A(n174), .B(n2542), .Z(n2540) );
  XOR U3316 ( .A(n2543), .B(n2544), .Z(n2542) );
  XOR U3317 ( .A(DB[588]), .B(DB[581]), .Z(n2544) );
  AND U3318 ( .A(n178), .B(n2545), .Z(n2543) );
  XOR U3319 ( .A(n2546), .B(n2547), .Z(n2545) );
  XOR U3320 ( .A(DB[581]), .B(DB[574]), .Z(n2547) );
  AND U3321 ( .A(n182), .B(n2548), .Z(n2546) );
  XOR U3322 ( .A(n2549), .B(n2550), .Z(n2548) );
  XOR U3323 ( .A(DB[574]), .B(DB[567]), .Z(n2550) );
  AND U3324 ( .A(n186), .B(n2551), .Z(n2549) );
  XOR U3325 ( .A(n2552), .B(n2553), .Z(n2551) );
  XOR U3326 ( .A(DB[567]), .B(DB[560]), .Z(n2553) );
  AND U3327 ( .A(n190), .B(n2554), .Z(n2552) );
  XOR U3328 ( .A(n2555), .B(n2556), .Z(n2554) );
  XOR U3329 ( .A(DB[560]), .B(DB[553]), .Z(n2556) );
  AND U3330 ( .A(n194), .B(n2557), .Z(n2555) );
  XOR U3331 ( .A(n2558), .B(n2559), .Z(n2557) );
  XOR U3332 ( .A(DB[553]), .B(DB[546]), .Z(n2559) );
  AND U3333 ( .A(n198), .B(n2560), .Z(n2558) );
  XOR U3334 ( .A(n2561), .B(n2562), .Z(n2560) );
  XOR U3335 ( .A(DB[546]), .B(DB[539]), .Z(n2562) );
  AND U3336 ( .A(n202), .B(n2563), .Z(n2561) );
  XOR U3337 ( .A(n2564), .B(n2565), .Z(n2563) );
  XOR U3338 ( .A(DB[539]), .B(DB[532]), .Z(n2565) );
  AND U3339 ( .A(n206), .B(n2566), .Z(n2564) );
  XOR U3340 ( .A(n2567), .B(n2568), .Z(n2566) );
  XOR U3341 ( .A(DB[532]), .B(DB[525]), .Z(n2568) );
  AND U3342 ( .A(n210), .B(n2569), .Z(n2567) );
  XOR U3343 ( .A(n2570), .B(n2571), .Z(n2569) );
  XOR U3344 ( .A(DB[525]), .B(DB[518]), .Z(n2571) );
  AND U3345 ( .A(n214), .B(n2572), .Z(n2570) );
  XOR U3346 ( .A(n2573), .B(n2574), .Z(n2572) );
  XOR U3347 ( .A(DB[518]), .B(DB[511]), .Z(n2574) );
  AND U3348 ( .A(n218), .B(n2575), .Z(n2573) );
  XOR U3349 ( .A(n2576), .B(n2577), .Z(n2575) );
  XOR U3350 ( .A(DB[511]), .B(DB[504]), .Z(n2577) );
  AND U3351 ( .A(n222), .B(n2578), .Z(n2576) );
  XOR U3352 ( .A(n2579), .B(n2580), .Z(n2578) );
  XOR U3353 ( .A(DB[504]), .B(DB[497]), .Z(n2580) );
  AND U3354 ( .A(n226), .B(n2581), .Z(n2579) );
  XOR U3355 ( .A(n2582), .B(n2583), .Z(n2581) );
  XOR U3356 ( .A(DB[497]), .B(DB[490]), .Z(n2583) );
  AND U3357 ( .A(n230), .B(n2584), .Z(n2582) );
  XOR U3358 ( .A(n2585), .B(n2586), .Z(n2584) );
  XOR U3359 ( .A(DB[490]), .B(DB[483]), .Z(n2586) );
  AND U3360 ( .A(n234), .B(n2587), .Z(n2585) );
  XOR U3361 ( .A(n2588), .B(n2589), .Z(n2587) );
  XOR U3362 ( .A(DB[483]), .B(DB[476]), .Z(n2589) );
  AND U3363 ( .A(n238), .B(n2590), .Z(n2588) );
  XOR U3364 ( .A(n2591), .B(n2592), .Z(n2590) );
  XOR U3365 ( .A(DB[476]), .B(DB[469]), .Z(n2592) );
  AND U3366 ( .A(n242), .B(n2593), .Z(n2591) );
  XOR U3367 ( .A(n2594), .B(n2595), .Z(n2593) );
  XOR U3368 ( .A(DB[469]), .B(DB[462]), .Z(n2595) );
  AND U3369 ( .A(n246), .B(n2596), .Z(n2594) );
  XOR U3370 ( .A(n2597), .B(n2598), .Z(n2596) );
  XOR U3371 ( .A(DB[462]), .B(DB[455]), .Z(n2598) );
  AND U3372 ( .A(n250), .B(n2599), .Z(n2597) );
  XOR U3373 ( .A(n2600), .B(n2601), .Z(n2599) );
  XOR U3374 ( .A(DB[455]), .B(DB[448]), .Z(n2601) );
  AND U3375 ( .A(n254), .B(n2602), .Z(n2600) );
  XOR U3376 ( .A(n2603), .B(n2604), .Z(n2602) );
  XOR U3377 ( .A(DB[448]), .B(DB[441]), .Z(n2604) );
  AND U3378 ( .A(n258), .B(n2605), .Z(n2603) );
  XOR U3379 ( .A(n2606), .B(n2607), .Z(n2605) );
  XOR U3380 ( .A(DB[441]), .B(DB[434]), .Z(n2607) );
  AND U3381 ( .A(n262), .B(n2608), .Z(n2606) );
  XOR U3382 ( .A(n2609), .B(n2610), .Z(n2608) );
  XOR U3383 ( .A(DB[434]), .B(DB[427]), .Z(n2610) );
  AND U3384 ( .A(n266), .B(n2611), .Z(n2609) );
  XOR U3385 ( .A(n2612), .B(n2613), .Z(n2611) );
  XOR U3386 ( .A(DB[427]), .B(DB[420]), .Z(n2613) );
  AND U3387 ( .A(n270), .B(n2614), .Z(n2612) );
  XOR U3388 ( .A(n2615), .B(n2616), .Z(n2614) );
  XOR U3389 ( .A(DB[420]), .B(DB[413]), .Z(n2616) );
  AND U3390 ( .A(n274), .B(n2617), .Z(n2615) );
  XOR U3391 ( .A(n2618), .B(n2619), .Z(n2617) );
  XOR U3392 ( .A(DB[413]), .B(DB[406]), .Z(n2619) );
  AND U3393 ( .A(n278), .B(n2620), .Z(n2618) );
  XOR U3394 ( .A(n2621), .B(n2622), .Z(n2620) );
  XOR U3395 ( .A(DB[406]), .B(DB[399]), .Z(n2622) );
  AND U3396 ( .A(n282), .B(n2623), .Z(n2621) );
  XOR U3397 ( .A(n2624), .B(n2625), .Z(n2623) );
  XOR U3398 ( .A(DB[399]), .B(DB[392]), .Z(n2625) );
  AND U3399 ( .A(n286), .B(n2626), .Z(n2624) );
  XOR U3400 ( .A(n2627), .B(n2628), .Z(n2626) );
  XOR U3401 ( .A(DB[392]), .B(DB[385]), .Z(n2628) );
  AND U3402 ( .A(n290), .B(n2629), .Z(n2627) );
  XOR U3403 ( .A(n2630), .B(n2631), .Z(n2629) );
  XOR U3404 ( .A(DB[385]), .B(DB[378]), .Z(n2631) );
  AND U3405 ( .A(n294), .B(n2632), .Z(n2630) );
  XOR U3406 ( .A(n2633), .B(n2634), .Z(n2632) );
  XOR U3407 ( .A(DB[378]), .B(DB[371]), .Z(n2634) );
  AND U3408 ( .A(n298), .B(n2635), .Z(n2633) );
  XOR U3409 ( .A(n2636), .B(n2637), .Z(n2635) );
  XOR U3410 ( .A(DB[371]), .B(DB[364]), .Z(n2637) );
  AND U3411 ( .A(n302), .B(n2638), .Z(n2636) );
  XOR U3412 ( .A(n2639), .B(n2640), .Z(n2638) );
  XOR U3413 ( .A(DB[364]), .B(DB[357]), .Z(n2640) );
  AND U3414 ( .A(n306), .B(n2641), .Z(n2639) );
  XOR U3415 ( .A(n2642), .B(n2643), .Z(n2641) );
  XOR U3416 ( .A(DB[357]), .B(DB[350]), .Z(n2643) );
  AND U3417 ( .A(n310), .B(n2644), .Z(n2642) );
  XOR U3418 ( .A(n2645), .B(n2646), .Z(n2644) );
  XOR U3419 ( .A(DB[350]), .B(DB[343]), .Z(n2646) );
  AND U3420 ( .A(n314), .B(n2647), .Z(n2645) );
  XOR U3421 ( .A(n2648), .B(n2649), .Z(n2647) );
  XOR U3422 ( .A(DB[343]), .B(DB[336]), .Z(n2649) );
  AND U3423 ( .A(n318), .B(n2650), .Z(n2648) );
  XOR U3424 ( .A(n2651), .B(n2652), .Z(n2650) );
  XOR U3425 ( .A(DB[336]), .B(DB[329]), .Z(n2652) );
  AND U3426 ( .A(n322), .B(n2653), .Z(n2651) );
  XOR U3427 ( .A(n2654), .B(n2655), .Z(n2653) );
  XOR U3428 ( .A(DB[329]), .B(DB[322]), .Z(n2655) );
  AND U3429 ( .A(n326), .B(n2656), .Z(n2654) );
  XOR U3430 ( .A(n2657), .B(n2658), .Z(n2656) );
  XOR U3431 ( .A(DB[322]), .B(DB[315]), .Z(n2658) );
  AND U3432 ( .A(n330), .B(n2659), .Z(n2657) );
  XOR U3433 ( .A(n2660), .B(n2661), .Z(n2659) );
  XOR U3434 ( .A(DB[315]), .B(DB[308]), .Z(n2661) );
  AND U3435 ( .A(n334), .B(n2662), .Z(n2660) );
  XOR U3436 ( .A(n2663), .B(n2664), .Z(n2662) );
  XOR U3437 ( .A(DB[308]), .B(DB[301]), .Z(n2664) );
  AND U3438 ( .A(n338), .B(n2665), .Z(n2663) );
  XOR U3439 ( .A(n2666), .B(n2667), .Z(n2665) );
  XOR U3440 ( .A(DB[301]), .B(DB[294]), .Z(n2667) );
  AND U3441 ( .A(n342), .B(n2668), .Z(n2666) );
  XOR U3442 ( .A(n2669), .B(n2670), .Z(n2668) );
  XOR U3443 ( .A(DB[294]), .B(DB[287]), .Z(n2670) );
  AND U3444 ( .A(n346), .B(n2671), .Z(n2669) );
  XOR U3445 ( .A(n2672), .B(n2673), .Z(n2671) );
  XOR U3446 ( .A(DB[287]), .B(DB[280]), .Z(n2673) );
  AND U3447 ( .A(n350), .B(n2674), .Z(n2672) );
  XOR U3448 ( .A(n2675), .B(n2676), .Z(n2674) );
  XOR U3449 ( .A(DB[280]), .B(DB[273]), .Z(n2676) );
  AND U3450 ( .A(n354), .B(n2677), .Z(n2675) );
  XOR U3451 ( .A(n2678), .B(n2679), .Z(n2677) );
  XOR U3452 ( .A(DB[273]), .B(DB[266]), .Z(n2679) );
  AND U3453 ( .A(n358), .B(n2680), .Z(n2678) );
  XOR U3454 ( .A(n2681), .B(n2682), .Z(n2680) );
  XOR U3455 ( .A(DB[266]), .B(DB[259]), .Z(n2682) );
  AND U3456 ( .A(n362), .B(n2683), .Z(n2681) );
  XOR U3457 ( .A(n2684), .B(n2685), .Z(n2683) );
  XOR U3458 ( .A(DB[259]), .B(DB[252]), .Z(n2685) );
  AND U3459 ( .A(n366), .B(n2686), .Z(n2684) );
  XOR U3460 ( .A(n2687), .B(n2688), .Z(n2686) );
  XOR U3461 ( .A(DB[252]), .B(DB[245]), .Z(n2688) );
  AND U3462 ( .A(n370), .B(n2689), .Z(n2687) );
  XOR U3463 ( .A(n2690), .B(n2691), .Z(n2689) );
  XOR U3464 ( .A(DB[245]), .B(DB[238]), .Z(n2691) );
  AND U3465 ( .A(n374), .B(n2692), .Z(n2690) );
  XOR U3466 ( .A(n2693), .B(n2694), .Z(n2692) );
  XOR U3467 ( .A(DB[238]), .B(DB[231]), .Z(n2694) );
  AND U3468 ( .A(n378), .B(n2695), .Z(n2693) );
  XOR U3469 ( .A(n2696), .B(n2697), .Z(n2695) );
  XOR U3470 ( .A(DB[231]), .B(DB[224]), .Z(n2697) );
  AND U3471 ( .A(n382), .B(n2698), .Z(n2696) );
  XOR U3472 ( .A(n2699), .B(n2700), .Z(n2698) );
  XOR U3473 ( .A(DB[224]), .B(DB[217]), .Z(n2700) );
  AND U3474 ( .A(n386), .B(n2701), .Z(n2699) );
  XOR U3475 ( .A(n2702), .B(n2703), .Z(n2701) );
  XOR U3476 ( .A(DB[217]), .B(DB[210]), .Z(n2703) );
  AND U3477 ( .A(n390), .B(n2704), .Z(n2702) );
  XOR U3478 ( .A(n2705), .B(n2706), .Z(n2704) );
  XOR U3479 ( .A(DB[210]), .B(DB[203]), .Z(n2706) );
  AND U3480 ( .A(n394), .B(n2707), .Z(n2705) );
  XOR U3481 ( .A(n2708), .B(n2709), .Z(n2707) );
  XOR U3482 ( .A(DB[203]), .B(DB[196]), .Z(n2709) );
  AND U3483 ( .A(n398), .B(n2710), .Z(n2708) );
  XOR U3484 ( .A(n2711), .B(n2712), .Z(n2710) );
  XOR U3485 ( .A(DB[196]), .B(DB[189]), .Z(n2712) );
  AND U3486 ( .A(n402), .B(n2713), .Z(n2711) );
  XOR U3487 ( .A(n2714), .B(n2715), .Z(n2713) );
  XOR U3488 ( .A(DB[189]), .B(DB[182]), .Z(n2715) );
  AND U3489 ( .A(n406), .B(n2716), .Z(n2714) );
  XOR U3490 ( .A(n2717), .B(n2718), .Z(n2716) );
  XOR U3491 ( .A(DB[182]), .B(DB[175]), .Z(n2718) );
  AND U3492 ( .A(n410), .B(n2719), .Z(n2717) );
  XOR U3493 ( .A(n2720), .B(n2721), .Z(n2719) );
  XOR U3494 ( .A(DB[175]), .B(DB[168]), .Z(n2721) );
  AND U3495 ( .A(n414), .B(n2722), .Z(n2720) );
  XOR U3496 ( .A(n2723), .B(n2724), .Z(n2722) );
  XOR U3497 ( .A(DB[168]), .B(DB[161]), .Z(n2724) );
  AND U3498 ( .A(n418), .B(n2725), .Z(n2723) );
  XOR U3499 ( .A(n2726), .B(n2727), .Z(n2725) );
  XOR U3500 ( .A(DB[161]), .B(DB[154]), .Z(n2727) );
  AND U3501 ( .A(n422), .B(n2728), .Z(n2726) );
  XOR U3502 ( .A(n2729), .B(n2730), .Z(n2728) );
  XOR U3503 ( .A(DB[154]), .B(DB[147]), .Z(n2730) );
  AND U3504 ( .A(n426), .B(n2731), .Z(n2729) );
  XOR U3505 ( .A(n2732), .B(n2733), .Z(n2731) );
  XOR U3506 ( .A(DB[147]), .B(DB[140]), .Z(n2733) );
  AND U3507 ( .A(n430), .B(n2734), .Z(n2732) );
  XOR U3508 ( .A(n2735), .B(n2736), .Z(n2734) );
  XOR U3509 ( .A(DB[140]), .B(DB[133]), .Z(n2736) );
  AND U3510 ( .A(n434), .B(n2737), .Z(n2735) );
  XOR U3511 ( .A(n2738), .B(n2739), .Z(n2737) );
  XOR U3512 ( .A(DB[133]), .B(DB[126]), .Z(n2739) );
  AND U3513 ( .A(n438), .B(n2740), .Z(n2738) );
  XOR U3514 ( .A(n2741), .B(n2742), .Z(n2740) );
  XOR U3515 ( .A(DB[126]), .B(DB[119]), .Z(n2742) );
  AND U3516 ( .A(n442), .B(n2743), .Z(n2741) );
  XOR U3517 ( .A(n2744), .B(n2745), .Z(n2743) );
  XOR U3518 ( .A(DB[119]), .B(DB[112]), .Z(n2745) );
  AND U3519 ( .A(n446), .B(n2746), .Z(n2744) );
  XOR U3520 ( .A(n2747), .B(n2748), .Z(n2746) );
  XOR U3521 ( .A(DB[112]), .B(DB[105]), .Z(n2748) );
  AND U3522 ( .A(n450), .B(n2749), .Z(n2747) );
  XOR U3523 ( .A(n2750), .B(n2751), .Z(n2749) );
  XOR U3524 ( .A(DB[98]), .B(DB[105]), .Z(n2751) );
  AND U3525 ( .A(n454), .B(n2752), .Z(n2750) );
  XOR U3526 ( .A(n2753), .B(n2754), .Z(n2752) );
  XOR U3527 ( .A(DB[98]), .B(DB[91]), .Z(n2754) );
  AND U3528 ( .A(n458), .B(n2755), .Z(n2753) );
  XOR U3529 ( .A(n2756), .B(n2757), .Z(n2755) );
  XOR U3530 ( .A(DB[91]), .B(DB[84]), .Z(n2757) );
  AND U3531 ( .A(n462), .B(n2758), .Z(n2756) );
  XOR U3532 ( .A(n2759), .B(n2760), .Z(n2758) );
  XOR U3533 ( .A(DB[84]), .B(DB[77]), .Z(n2760) );
  AND U3534 ( .A(n466), .B(n2761), .Z(n2759) );
  XOR U3535 ( .A(n2762), .B(n2763), .Z(n2761) );
  XOR U3536 ( .A(DB[77]), .B(DB[70]), .Z(n2763) );
  AND U3537 ( .A(n470), .B(n2764), .Z(n2762) );
  XOR U3538 ( .A(n2765), .B(n2766), .Z(n2764) );
  XOR U3539 ( .A(DB[70]), .B(DB[63]), .Z(n2766) );
  AND U3540 ( .A(n474), .B(n2767), .Z(n2765) );
  XOR U3541 ( .A(n2768), .B(n2769), .Z(n2767) );
  XOR U3542 ( .A(DB[63]), .B(DB[56]), .Z(n2769) );
  AND U3543 ( .A(n478), .B(n2770), .Z(n2768) );
  XOR U3544 ( .A(n2771), .B(n2772), .Z(n2770) );
  XOR U3545 ( .A(DB[56]), .B(DB[49]), .Z(n2772) );
  AND U3546 ( .A(n482), .B(n2773), .Z(n2771) );
  XOR U3547 ( .A(n2774), .B(n2775), .Z(n2773) );
  XOR U3548 ( .A(DB[49]), .B(DB[42]), .Z(n2775) );
  AND U3549 ( .A(n486), .B(n2776), .Z(n2774) );
  XOR U3550 ( .A(n2777), .B(n2778), .Z(n2776) );
  XOR U3551 ( .A(DB[42]), .B(DB[35]), .Z(n2778) );
  AND U3552 ( .A(n490), .B(n2779), .Z(n2777) );
  XOR U3553 ( .A(n2780), .B(n2781), .Z(n2779) );
  XOR U3554 ( .A(DB[35]), .B(DB[28]), .Z(n2781) );
  AND U3555 ( .A(n494), .B(n2782), .Z(n2780) );
  XOR U3556 ( .A(n2783), .B(n2784), .Z(n2782) );
  XOR U3557 ( .A(DB[28]), .B(DB[21]), .Z(n2784) );
  AND U3558 ( .A(n498), .B(n2785), .Z(n2783) );
  XOR U3559 ( .A(n2786), .B(n2787), .Z(n2785) );
  XOR U3560 ( .A(DB[21]), .B(DB[14]), .Z(n2787) );
  AND U3561 ( .A(n502), .B(n2788), .Z(n2786) );
  XOR U3562 ( .A(n2789), .B(n2790), .Z(n2788) );
  XOR U3563 ( .A(DB[7]), .B(DB[14]), .Z(n2790) );
  AND U3564 ( .A(n506), .B(n2791), .Z(n2789) );
  XOR U3565 ( .A(DB[7]), .B(DB[0]), .Z(n2791) );
  XOR U3566 ( .A(n2792), .B(n2793), .Z(n2) );
  AND U3567 ( .A(n2794), .B(n2795), .Z(n2792) );
  XNOR U3568 ( .A(n2793), .B(n2796), .Z(n2795) );
  XOR U3569 ( .A(n2797), .B(n2798), .Z(n2796) );
  AND U3570 ( .A(n2799), .B(n2800), .Z(n2797) );
  XNOR U3571 ( .A(n2801), .B(n2802), .Z(n2800) );
  XNOR U3572 ( .A(n2793), .B(n2803), .Z(n2794) );
  XNOR U3573 ( .A(n2804), .B(n2805), .Z(n2803) );
  AND U3574 ( .A(n6), .B(n2806), .Z(n2804) );
  XOR U3575 ( .A(n2807), .B(n2805), .Z(n2806) );
  XNOR U3576 ( .A(n2808), .B(n2809), .Z(n2793) );
  NAND U3577 ( .A(n2810), .B(n2811), .Z(n2809) );
  XOR U3578 ( .A(n2799), .B(n2812), .Z(n2811) );
  XNOR U3579 ( .A(n2808), .B(n2801), .Z(n2812) );
  XOR U3580 ( .A(n2813), .B(n2814), .Z(n2801) );
  ANDN U3581 ( .B(n2815), .A(n2816), .Z(n2813) );
  XNOR U3582 ( .A(n2814), .B(n2817), .Z(n2815) );
  XNOR U3583 ( .A(n2798), .B(n2818), .Z(n2799) );
  XNOR U3584 ( .A(n2819), .B(n2820), .Z(n2818) );
  ANDN U3585 ( .B(n2821), .A(n2822), .Z(n2819) );
  XNOR U3586 ( .A(n2823), .B(n2824), .Z(n2821) );
  IV U3587 ( .A(n2820), .Z(n2824) );
  IV U3588 ( .A(n2802), .Z(n2798) );
  XNOR U3589 ( .A(n2825), .B(n2826), .Z(n2802) );
  AND U3590 ( .A(n2827), .B(n2828), .Z(n2825) );
  XNOR U3591 ( .A(n2826), .B(n2829), .Z(n2828) );
  XOR U3592 ( .A(n2830), .B(n2831), .Z(n2810) );
  XNOR U3593 ( .A(n2808), .B(n2832), .Z(n2831) );
  NAND U3594 ( .A(n2833), .B(n6), .Z(n2832) );
  XOR U3595 ( .A(n2834), .B(n2830), .Z(n2833) );
  NAND U3596 ( .A(n2835), .B(n2836), .Z(n2808) );
  XNOR U3597 ( .A(n2827), .B(n2829), .Z(n2836) );
  XOR U3598 ( .A(n2837), .B(n2817), .Z(n2829) );
  XNOR U3599 ( .A(q[6]), .B(DB[895]), .Z(n2817) );
  IV U3600 ( .A(n2816), .Z(n2837) );
  XOR U3601 ( .A(n2814), .B(n2838), .Z(n2816) );
  XNOR U3602 ( .A(q[5]), .B(DB[894]), .Z(n2838) );
  XOR U3603 ( .A(q[4]), .B(DB[893]), .Z(n2814) );
  XNOR U3604 ( .A(n2839), .B(n2840), .Z(n2827) );
  XNOR U3605 ( .A(n2823), .B(n2826), .Z(n2840) );
  XOR U3606 ( .A(q[0]), .B(DB[889]), .Z(n2826) );
  XOR U3607 ( .A(q[3]), .B(DB[892]), .Z(n2823) );
  IV U3608 ( .A(n2822), .Z(n2839) );
  XOR U3609 ( .A(n2820), .B(n2841), .Z(n2822) );
  XNOR U3610 ( .A(q[2]), .B(DB[891]), .Z(n2841) );
  XOR U3611 ( .A(q[1]), .B(DB[890]), .Z(n2820) );
  XOR U3612 ( .A(n2842), .B(n2843), .Z(n2835) );
  AND U3613 ( .A(n6), .B(n2844), .Z(n2842) );
  XOR U3614 ( .A(n2843), .B(n2845), .Z(n2844) );
  XOR U3615 ( .A(n2846), .B(n2847), .Z(n6) );
  AND U3616 ( .A(n2848), .B(n2849), .Z(n2846) );
  XNOR U3617 ( .A(n2847), .B(n2805), .Z(n2849) );
  XNOR U3618 ( .A(n2850), .B(n2851), .Z(n2805) );
  ANDN U3619 ( .B(n2852), .A(n2853), .Z(n2850) );
  XOR U3620 ( .A(n2851), .B(n2854), .Z(n2852) );
  XOR U3621 ( .A(n2847), .B(n2807), .Z(n2848) );
  XOR U3622 ( .A(n2855), .B(n2856), .Z(n2807) );
  AND U3623 ( .A(n10), .B(n2857), .Z(n2855) );
  XOR U3624 ( .A(n2858), .B(n2856), .Z(n2857) );
  XNOR U3625 ( .A(n2859), .B(n2860), .Z(n2847) );
  NAND U3626 ( .A(n2861), .B(n2862), .Z(n2860) );
  XOR U3627 ( .A(n2863), .B(n2830), .Z(n2862) );
  XNOR U3628 ( .A(n2864), .B(n2854), .Z(n2830) );
  XOR U3629 ( .A(n2865), .B(n2866), .Z(n2854) );
  ANDN U3630 ( .B(n2867), .A(n2868), .Z(n2865) );
  XOR U3631 ( .A(n2866), .B(n2869), .Z(n2867) );
  IV U3632 ( .A(n2853), .Z(n2864) );
  XOR U3633 ( .A(n2870), .B(n2871), .Z(n2853) );
  XOR U3634 ( .A(n2872), .B(n2873), .Z(n2871) );
  ANDN U3635 ( .B(n2874), .A(n2875), .Z(n2872) );
  XOR U3636 ( .A(n2876), .B(n2873), .Z(n2874) );
  IV U3637 ( .A(n2851), .Z(n2870) );
  XOR U3638 ( .A(n2877), .B(n2878), .Z(n2851) );
  ANDN U3639 ( .B(n2879), .A(n2880), .Z(n2877) );
  XOR U3640 ( .A(n2878), .B(n2881), .Z(n2879) );
  IV U3641 ( .A(n2859), .Z(n2863) );
  XOR U3642 ( .A(n2859), .B(n2834), .Z(n2861) );
  XOR U3643 ( .A(n2882), .B(n2883), .Z(n2834) );
  AND U3644 ( .A(n10), .B(n2884), .Z(n2882) );
  XOR U3645 ( .A(n2885), .B(n2883), .Z(n2884) );
  NANDN U3646 ( .A(n2843), .B(n2845), .Z(n2859) );
  XOR U3647 ( .A(n2886), .B(n2887), .Z(n2845) );
  AND U3648 ( .A(n10), .B(n2888), .Z(n2886) );
  XOR U3649 ( .A(n2887), .B(n2889), .Z(n2888) );
  XOR U3650 ( .A(n2890), .B(n2891), .Z(n10) );
  AND U3651 ( .A(n2892), .B(n2893), .Z(n2890) );
  XNOR U3652 ( .A(n2891), .B(n2856), .Z(n2893) );
  XNOR U3653 ( .A(n2894), .B(n2895), .Z(n2856) );
  ANDN U3654 ( .B(n2896), .A(n2897), .Z(n2894) );
  XOR U3655 ( .A(n2895), .B(n2898), .Z(n2896) );
  XOR U3656 ( .A(n2891), .B(n2858), .Z(n2892) );
  XOR U3657 ( .A(n2899), .B(n2900), .Z(n2858) );
  AND U3658 ( .A(n14), .B(n2901), .Z(n2899) );
  XOR U3659 ( .A(n2902), .B(n2900), .Z(n2901) );
  XNOR U3660 ( .A(n2903), .B(n2904), .Z(n2891) );
  NAND U3661 ( .A(n2905), .B(n2906), .Z(n2904) );
  XOR U3662 ( .A(n2907), .B(n2883), .Z(n2906) );
  XOR U3663 ( .A(n2897), .B(n2898), .Z(n2883) );
  XOR U3664 ( .A(n2908), .B(n2909), .Z(n2898) );
  ANDN U3665 ( .B(n2910), .A(n2911), .Z(n2908) );
  XOR U3666 ( .A(n2909), .B(n2912), .Z(n2910) );
  XOR U3667 ( .A(n2913), .B(n2914), .Z(n2897) );
  XOR U3668 ( .A(n2915), .B(n2916), .Z(n2914) );
  ANDN U3669 ( .B(n2917), .A(n2918), .Z(n2915) );
  XOR U3670 ( .A(n2919), .B(n2916), .Z(n2917) );
  IV U3671 ( .A(n2895), .Z(n2913) );
  XOR U3672 ( .A(n2920), .B(n2921), .Z(n2895) );
  ANDN U3673 ( .B(n2922), .A(n2923), .Z(n2920) );
  XOR U3674 ( .A(n2921), .B(n2924), .Z(n2922) );
  IV U3675 ( .A(n2903), .Z(n2907) );
  XOR U3676 ( .A(n2903), .B(n2885), .Z(n2905) );
  XOR U3677 ( .A(n2925), .B(n2926), .Z(n2885) );
  AND U3678 ( .A(n14), .B(n2927), .Z(n2925) );
  XOR U3679 ( .A(n2928), .B(n2926), .Z(n2927) );
  NANDN U3680 ( .A(n2887), .B(n2889), .Z(n2903) );
  XOR U3681 ( .A(n2929), .B(n2930), .Z(n2889) );
  AND U3682 ( .A(n14), .B(n2931), .Z(n2929) );
  XOR U3683 ( .A(n2930), .B(n2932), .Z(n2931) );
  XOR U3684 ( .A(n2933), .B(n2934), .Z(n14) );
  AND U3685 ( .A(n2935), .B(n2936), .Z(n2933) );
  XNOR U3686 ( .A(n2934), .B(n2900), .Z(n2936) );
  XNOR U3687 ( .A(n2937), .B(n2938), .Z(n2900) );
  ANDN U3688 ( .B(n2939), .A(n2940), .Z(n2937) );
  XOR U3689 ( .A(n2938), .B(n2941), .Z(n2939) );
  XOR U3690 ( .A(n2934), .B(n2902), .Z(n2935) );
  XOR U3691 ( .A(n2942), .B(n2943), .Z(n2902) );
  AND U3692 ( .A(n18), .B(n2944), .Z(n2942) );
  XOR U3693 ( .A(n2945), .B(n2943), .Z(n2944) );
  XNOR U3694 ( .A(n2946), .B(n2947), .Z(n2934) );
  NAND U3695 ( .A(n2948), .B(n2949), .Z(n2947) );
  XOR U3696 ( .A(n2950), .B(n2926), .Z(n2949) );
  XOR U3697 ( .A(n2940), .B(n2941), .Z(n2926) );
  XOR U3698 ( .A(n2951), .B(n2952), .Z(n2941) );
  ANDN U3699 ( .B(n2953), .A(n2954), .Z(n2951) );
  XOR U3700 ( .A(n2952), .B(n2955), .Z(n2953) );
  XOR U3701 ( .A(n2956), .B(n2957), .Z(n2940) );
  XOR U3702 ( .A(n2958), .B(n2959), .Z(n2957) );
  ANDN U3703 ( .B(n2960), .A(n2961), .Z(n2958) );
  XOR U3704 ( .A(n2962), .B(n2959), .Z(n2960) );
  IV U3705 ( .A(n2938), .Z(n2956) );
  XOR U3706 ( .A(n2963), .B(n2964), .Z(n2938) );
  ANDN U3707 ( .B(n2965), .A(n2966), .Z(n2963) );
  XOR U3708 ( .A(n2964), .B(n2967), .Z(n2965) );
  IV U3709 ( .A(n2946), .Z(n2950) );
  XOR U3710 ( .A(n2946), .B(n2928), .Z(n2948) );
  XOR U3711 ( .A(n2968), .B(n2969), .Z(n2928) );
  AND U3712 ( .A(n18), .B(n2970), .Z(n2968) );
  XOR U3713 ( .A(n2971), .B(n2969), .Z(n2970) );
  NANDN U3714 ( .A(n2930), .B(n2932), .Z(n2946) );
  XOR U3715 ( .A(n2972), .B(n2973), .Z(n2932) );
  AND U3716 ( .A(n18), .B(n2974), .Z(n2972) );
  XOR U3717 ( .A(n2973), .B(n2975), .Z(n2974) );
  XOR U3718 ( .A(n2976), .B(n2977), .Z(n18) );
  AND U3719 ( .A(n2978), .B(n2979), .Z(n2976) );
  XNOR U3720 ( .A(n2977), .B(n2943), .Z(n2979) );
  XNOR U3721 ( .A(n2980), .B(n2981), .Z(n2943) );
  ANDN U3722 ( .B(n2982), .A(n2983), .Z(n2980) );
  XOR U3723 ( .A(n2981), .B(n2984), .Z(n2982) );
  XOR U3724 ( .A(n2977), .B(n2945), .Z(n2978) );
  XOR U3725 ( .A(n2985), .B(n2986), .Z(n2945) );
  AND U3726 ( .A(n22), .B(n2987), .Z(n2985) );
  XOR U3727 ( .A(n2988), .B(n2986), .Z(n2987) );
  XNOR U3728 ( .A(n2989), .B(n2990), .Z(n2977) );
  NAND U3729 ( .A(n2991), .B(n2992), .Z(n2990) );
  XOR U3730 ( .A(n2993), .B(n2969), .Z(n2992) );
  XOR U3731 ( .A(n2983), .B(n2984), .Z(n2969) );
  XOR U3732 ( .A(n2994), .B(n2995), .Z(n2984) );
  ANDN U3733 ( .B(n2996), .A(n2997), .Z(n2994) );
  XOR U3734 ( .A(n2995), .B(n2998), .Z(n2996) );
  XOR U3735 ( .A(n2999), .B(n3000), .Z(n2983) );
  XOR U3736 ( .A(n3001), .B(n3002), .Z(n3000) );
  ANDN U3737 ( .B(n3003), .A(n3004), .Z(n3001) );
  XOR U3738 ( .A(n3005), .B(n3002), .Z(n3003) );
  IV U3739 ( .A(n2981), .Z(n2999) );
  XOR U3740 ( .A(n3006), .B(n3007), .Z(n2981) );
  ANDN U3741 ( .B(n3008), .A(n3009), .Z(n3006) );
  XOR U3742 ( .A(n3007), .B(n3010), .Z(n3008) );
  IV U3743 ( .A(n2989), .Z(n2993) );
  XOR U3744 ( .A(n2989), .B(n2971), .Z(n2991) );
  XOR U3745 ( .A(n3011), .B(n3012), .Z(n2971) );
  AND U3746 ( .A(n22), .B(n3013), .Z(n3011) );
  XOR U3747 ( .A(n3014), .B(n3012), .Z(n3013) );
  NANDN U3748 ( .A(n2973), .B(n2975), .Z(n2989) );
  XOR U3749 ( .A(n3015), .B(n3016), .Z(n2975) );
  AND U3750 ( .A(n22), .B(n3017), .Z(n3015) );
  XOR U3751 ( .A(n3016), .B(n3018), .Z(n3017) );
  XOR U3752 ( .A(n3019), .B(n3020), .Z(n22) );
  AND U3753 ( .A(n3021), .B(n3022), .Z(n3019) );
  XNOR U3754 ( .A(n3020), .B(n2986), .Z(n3022) );
  XNOR U3755 ( .A(n3023), .B(n3024), .Z(n2986) );
  ANDN U3756 ( .B(n3025), .A(n3026), .Z(n3023) );
  XOR U3757 ( .A(n3024), .B(n3027), .Z(n3025) );
  XOR U3758 ( .A(n3020), .B(n2988), .Z(n3021) );
  XOR U3759 ( .A(n3028), .B(n3029), .Z(n2988) );
  AND U3760 ( .A(n26), .B(n3030), .Z(n3028) );
  XOR U3761 ( .A(n3031), .B(n3029), .Z(n3030) );
  XNOR U3762 ( .A(n3032), .B(n3033), .Z(n3020) );
  NAND U3763 ( .A(n3034), .B(n3035), .Z(n3033) );
  XOR U3764 ( .A(n3036), .B(n3012), .Z(n3035) );
  XOR U3765 ( .A(n3026), .B(n3027), .Z(n3012) );
  XOR U3766 ( .A(n3037), .B(n3038), .Z(n3027) );
  ANDN U3767 ( .B(n3039), .A(n3040), .Z(n3037) );
  XOR U3768 ( .A(n3038), .B(n3041), .Z(n3039) );
  XOR U3769 ( .A(n3042), .B(n3043), .Z(n3026) );
  XOR U3770 ( .A(n3044), .B(n3045), .Z(n3043) );
  ANDN U3771 ( .B(n3046), .A(n3047), .Z(n3044) );
  XOR U3772 ( .A(n3048), .B(n3045), .Z(n3046) );
  IV U3773 ( .A(n3024), .Z(n3042) );
  XOR U3774 ( .A(n3049), .B(n3050), .Z(n3024) );
  ANDN U3775 ( .B(n3051), .A(n3052), .Z(n3049) );
  XOR U3776 ( .A(n3050), .B(n3053), .Z(n3051) );
  IV U3777 ( .A(n3032), .Z(n3036) );
  XOR U3778 ( .A(n3032), .B(n3014), .Z(n3034) );
  XOR U3779 ( .A(n3054), .B(n3055), .Z(n3014) );
  AND U3780 ( .A(n26), .B(n3056), .Z(n3054) );
  XOR U3781 ( .A(n3057), .B(n3055), .Z(n3056) );
  NANDN U3782 ( .A(n3016), .B(n3018), .Z(n3032) );
  XOR U3783 ( .A(n3058), .B(n3059), .Z(n3018) );
  AND U3784 ( .A(n26), .B(n3060), .Z(n3058) );
  XOR U3785 ( .A(n3059), .B(n3061), .Z(n3060) );
  XOR U3786 ( .A(n3062), .B(n3063), .Z(n26) );
  AND U3787 ( .A(n3064), .B(n3065), .Z(n3062) );
  XNOR U3788 ( .A(n3063), .B(n3029), .Z(n3065) );
  XNOR U3789 ( .A(n3066), .B(n3067), .Z(n3029) );
  ANDN U3790 ( .B(n3068), .A(n3069), .Z(n3066) );
  XOR U3791 ( .A(n3067), .B(n3070), .Z(n3068) );
  XOR U3792 ( .A(n3063), .B(n3031), .Z(n3064) );
  XOR U3793 ( .A(n3071), .B(n3072), .Z(n3031) );
  AND U3794 ( .A(n30), .B(n3073), .Z(n3071) );
  XOR U3795 ( .A(n3074), .B(n3072), .Z(n3073) );
  XNOR U3796 ( .A(n3075), .B(n3076), .Z(n3063) );
  NAND U3797 ( .A(n3077), .B(n3078), .Z(n3076) );
  XOR U3798 ( .A(n3079), .B(n3055), .Z(n3078) );
  XOR U3799 ( .A(n3069), .B(n3070), .Z(n3055) );
  XOR U3800 ( .A(n3080), .B(n3081), .Z(n3070) );
  ANDN U3801 ( .B(n3082), .A(n3083), .Z(n3080) );
  XOR U3802 ( .A(n3081), .B(n3084), .Z(n3082) );
  XOR U3803 ( .A(n3085), .B(n3086), .Z(n3069) );
  XOR U3804 ( .A(n3087), .B(n3088), .Z(n3086) );
  ANDN U3805 ( .B(n3089), .A(n3090), .Z(n3087) );
  XOR U3806 ( .A(n3091), .B(n3088), .Z(n3089) );
  IV U3807 ( .A(n3067), .Z(n3085) );
  XOR U3808 ( .A(n3092), .B(n3093), .Z(n3067) );
  ANDN U3809 ( .B(n3094), .A(n3095), .Z(n3092) );
  XOR U3810 ( .A(n3093), .B(n3096), .Z(n3094) );
  IV U3811 ( .A(n3075), .Z(n3079) );
  XOR U3812 ( .A(n3075), .B(n3057), .Z(n3077) );
  XOR U3813 ( .A(n3097), .B(n3098), .Z(n3057) );
  AND U3814 ( .A(n30), .B(n3099), .Z(n3097) );
  XOR U3815 ( .A(n3100), .B(n3098), .Z(n3099) );
  NANDN U3816 ( .A(n3059), .B(n3061), .Z(n3075) );
  XOR U3817 ( .A(n3101), .B(n3102), .Z(n3061) );
  AND U3818 ( .A(n30), .B(n3103), .Z(n3101) );
  XOR U3819 ( .A(n3102), .B(n3104), .Z(n3103) );
  XOR U3820 ( .A(n3105), .B(n3106), .Z(n30) );
  AND U3821 ( .A(n3107), .B(n3108), .Z(n3105) );
  XNOR U3822 ( .A(n3106), .B(n3072), .Z(n3108) );
  XNOR U3823 ( .A(n3109), .B(n3110), .Z(n3072) );
  ANDN U3824 ( .B(n3111), .A(n3112), .Z(n3109) );
  XOR U3825 ( .A(n3110), .B(n3113), .Z(n3111) );
  XOR U3826 ( .A(n3106), .B(n3074), .Z(n3107) );
  XOR U3827 ( .A(n3114), .B(n3115), .Z(n3074) );
  AND U3828 ( .A(n34), .B(n3116), .Z(n3114) );
  XOR U3829 ( .A(n3117), .B(n3115), .Z(n3116) );
  XNOR U3830 ( .A(n3118), .B(n3119), .Z(n3106) );
  NAND U3831 ( .A(n3120), .B(n3121), .Z(n3119) );
  XOR U3832 ( .A(n3122), .B(n3098), .Z(n3121) );
  XOR U3833 ( .A(n3112), .B(n3113), .Z(n3098) );
  XOR U3834 ( .A(n3123), .B(n3124), .Z(n3113) );
  ANDN U3835 ( .B(n3125), .A(n3126), .Z(n3123) );
  XOR U3836 ( .A(n3124), .B(n3127), .Z(n3125) );
  XOR U3837 ( .A(n3128), .B(n3129), .Z(n3112) );
  XOR U3838 ( .A(n3130), .B(n3131), .Z(n3129) );
  ANDN U3839 ( .B(n3132), .A(n3133), .Z(n3130) );
  XOR U3840 ( .A(n3134), .B(n3131), .Z(n3132) );
  IV U3841 ( .A(n3110), .Z(n3128) );
  XOR U3842 ( .A(n3135), .B(n3136), .Z(n3110) );
  ANDN U3843 ( .B(n3137), .A(n3138), .Z(n3135) );
  XOR U3844 ( .A(n3136), .B(n3139), .Z(n3137) );
  IV U3845 ( .A(n3118), .Z(n3122) );
  XOR U3846 ( .A(n3118), .B(n3100), .Z(n3120) );
  XOR U3847 ( .A(n3140), .B(n3141), .Z(n3100) );
  AND U3848 ( .A(n34), .B(n3142), .Z(n3140) );
  XOR U3849 ( .A(n3143), .B(n3141), .Z(n3142) );
  NANDN U3850 ( .A(n3102), .B(n3104), .Z(n3118) );
  XOR U3851 ( .A(n3144), .B(n3145), .Z(n3104) );
  AND U3852 ( .A(n34), .B(n3146), .Z(n3144) );
  XOR U3853 ( .A(n3145), .B(n3147), .Z(n3146) );
  XOR U3854 ( .A(n3148), .B(n3149), .Z(n34) );
  AND U3855 ( .A(n3150), .B(n3151), .Z(n3148) );
  XNOR U3856 ( .A(n3149), .B(n3115), .Z(n3151) );
  XNOR U3857 ( .A(n3152), .B(n3153), .Z(n3115) );
  ANDN U3858 ( .B(n3154), .A(n3155), .Z(n3152) );
  XOR U3859 ( .A(n3153), .B(n3156), .Z(n3154) );
  XOR U3860 ( .A(n3149), .B(n3117), .Z(n3150) );
  XOR U3861 ( .A(n3157), .B(n3158), .Z(n3117) );
  AND U3862 ( .A(n38), .B(n3159), .Z(n3157) );
  XOR U3863 ( .A(n3160), .B(n3158), .Z(n3159) );
  XNOR U3864 ( .A(n3161), .B(n3162), .Z(n3149) );
  NAND U3865 ( .A(n3163), .B(n3164), .Z(n3162) );
  XOR U3866 ( .A(n3165), .B(n3141), .Z(n3164) );
  XOR U3867 ( .A(n3155), .B(n3156), .Z(n3141) );
  XOR U3868 ( .A(n3166), .B(n3167), .Z(n3156) );
  ANDN U3869 ( .B(n3168), .A(n3169), .Z(n3166) );
  XOR U3870 ( .A(n3167), .B(n3170), .Z(n3168) );
  XOR U3871 ( .A(n3171), .B(n3172), .Z(n3155) );
  XOR U3872 ( .A(n3173), .B(n3174), .Z(n3172) );
  ANDN U3873 ( .B(n3175), .A(n3176), .Z(n3173) );
  XOR U3874 ( .A(n3177), .B(n3174), .Z(n3175) );
  IV U3875 ( .A(n3153), .Z(n3171) );
  XOR U3876 ( .A(n3178), .B(n3179), .Z(n3153) );
  ANDN U3877 ( .B(n3180), .A(n3181), .Z(n3178) );
  XOR U3878 ( .A(n3179), .B(n3182), .Z(n3180) );
  IV U3879 ( .A(n3161), .Z(n3165) );
  XOR U3880 ( .A(n3161), .B(n3143), .Z(n3163) );
  XOR U3881 ( .A(n3183), .B(n3184), .Z(n3143) );
  AND U3882 ( .A(n38), .B(n3185), .Z(n3183) );
  XOR U3883 ( .A(n3186), .B(n3184), .Z(n3185) );
  NANDN U3884 ( .A(n3145), .B(n3147), .Z(n3161) );
  XOR U3885 ( .A(n3187), .B(n3188), .Z(n3147) );
  AND U3886 ( .A(n38), .B(n3189), .Z(n3187) );
  XOR U3887 ( .A(n3188), .B(n3190), .Z(n3189) );
  XOR U3888 ( .A(n3191), .B(n3192), .Z(n38) );
  AND U3889 ( .A(n3193), .B(n3194), .Z(n3191) );
  XNOR U3890 ( .A(n3192), .B(n3158), .Z(n3194) );
  XNOR U3891 ( .A(n3195), .B(n3196), .Z(n3158) );
  ANDN U3892 ( .B(n3197), .A(n3198), .Z(n3195) );
  XOR U3893 ( .A(n3196), .B(n3199), .Z(n3197) );
  XOR U3894 ( .A(n3192), .B(n3160), .Z(n3193) );
  XOR U3895 ( .A(n3200), .B(n3201), .Z(n3160) );
  AND U3896 ( .A(n42), .B(n3202), .Z(n3200) );
  XOR U3897 ( .A(n3203), .B(n3201), .Z(n3202) );
  XNOR U3898 ( .A(n3204), .B(n3205), .Z(n3192) );
  NAND U3899 ( .A(n3206), .B(n3207), .Z(n3205) );
  XOR U3900 ( .A(n3208), .B(n3184), .Z(n3207) );
  XOR U3901 ( .A(n3198), .B(n3199), .Z(n3184) );
  XOR U3902 ( .A(n3209), .B(n3210), .Z(n3199) );
  ANDN U3903 ( .B(n3211), .A(n3212), .Z(n3209) );
  XOR U3904 ( .A(n3210), .B(n3213), .Z(n3211) );
  XOR U3905 ( .A(n3214), .B(n3215), .Z(n3198) );
  XOR U3906 ( .A(n3216), .B(n3217), .Z(n3215) );
  ANDN U3907 ( .B(n3218), .A(n3219), .Z(n3216) );
  XOR U3908 ( .A(n3220), .B(n3217), .Z(n3218) );
  IV U3909 ( .A(n3196), .Z(n3214) );
  XOR U3910 ( .A(n3221), .B(n3222), .Z(n3196) );
  ANDN U3911 ( .B(n3223), .A(n3224), .Z(n3221) );
  XOR U3912 ( .A(n3222), .B(n3225), .Z(n3223) );
  IV U3913 ( .A(n3204), .Z(n3208) );
  XOR U3914 ( .A(n3204), .B(n3186), .Z(n3206) );
  XOR U3915 ( .A(n3226), .B(n3227), .Z(n3186) );
  AND U3916 ( .A(n42), .B(n3228), .Z(n3226) );
  XOR U3917 ( .A(n3229), .B(n3227), .Z(n3228) );
  NANDN U3918 ( .A(n3188), .B(n3190), .Z(n3204) );
  XOR U3919 ( .A(n3230), .B(n3231), .Z(n3190) );
  AND U3920 ( .A(n42), .B(n3232), .Z(n3230) );
  XOR U3921 ( .A(n3231), .B(n3233), .Z(n3232) );
  XOR U3922 ( .A(n3234), .B(n3235), .Z(n42) );
  AND U3923 ( .A(n3236), .B(n3237), .Z(n3234) );
  XNOR U3924 ( .A(n3235), .B(n3201), .Z(n3237) );
  XNOR U3925 ( .A(n3238), .B(n3239), .Z(n3201) );
  ANDN U3926 ( .B(n3240), .A(n3241), .Z(n3238) );
  XOR U3927 ( .A(n3239), .B(n3242), .Z(n3240) );
  XOR U3928 ( .A(n3235), .B(n3203), .Z(n3236) );
  XOR U3929 ( .A(n3243), .B(n3244), .Z(n3203) );
  AND U3930 ( .A(n46), .B(n3245), .Z(n3243) );
  XOR U3931 ( .A(n3246), .B(n3244), .Z(n3245) );
  XNOR U3932 ( .A(n3247), .B(n3248), .Z(n3235) );
  NAND U3933 ( .A(n3249), .B(n3250), .Z(n3248) );
  XOR U3934 ( .A(n3251), .B(n3227), .Z(n3250) );
  XOR U3935 ( .A(n3241), .B(n3242), .Z(n3227) );
  XOR U3936 ( .A(n3252), .B(n3253), .Z(n3242) );
  ANDN U3937 ( .B(n3254), .A(n3255), .Z(n3252) );
  XOR U3938 ( .A(n3253), .B(n3256), .Z(n3254) );
  XOR U3939 ( .A(n3257), .B(n3258), .Z(n3241) );
  XOR U3940 ( .A(n3259), .B(n3260), .Z(n3258) );
  ANDN U3941 ( .B(n3261), .A(n3262), .Z(n3259) );
  XOR U3942 ( .A(n3263), .B(n3260), .Z(n3261) );
  IV U3943 ( .A(n3239), .Z(n3257) );
  XOR U3944 ( .A(n3264), .B(n3265), .Z(n3239) );
  ANDN U3945 ( .B(n3266), .A(n3267), .Z(n3264) );
  XOR U3946 ( .A(n3265), .B(n3268), .Z(n3266) );
  IV U3947 ( .A(n3247), .Z(n3251) );
  XOR U3948 ( .A(n3247), .B(n3229), .Z(n3249) );
  XOR U3949 ( .A(n3269), .B(n3270), .Z(n3229) );
  AND U3950 ( .A(n46), .B(n3271), .Z(n3269) );
  XOR U3951 ( .A(n3272), .B(n3270), .Z(n3271) );
  NANDN U3952 ( .A(n3231), .B(n3233), .Z(n3247) );
  XOR U3953 ( .A(n3273), .B(n3274), .Z(n3233) );
  AND U3954 ( .A(n46), .B(n3275), .Z(n3273) );
  XOR U3955 ( .A(n3274), .B(n3276), .Z(n3275) );
  XOR U3956 ( .A(n3277), .B(n3278), .Z(n46) );
  AND U3957 ( .A(n3279), .B(n3280), .Z(n3277) );
  XNOR U3958 ( .A(n3278), .B(n3244), .Z(n3280) );
  XNOR U3959 ( .A(n3281), .B(n3282), .Z(n3244) );
  ANDN U3960 ( .B(n3283), .A(n3284), .Z(n3281) );
  XOR U3961 ( .A(n3282), .B(n3285), .Z(n3283) );
  XOR U3962 ( .A(n3278), .B(n3246), .Z(n3279) );
  XOR U3963 ( .A(n3286), .B(n3287), .Z(n3246) );
  AND U3964 ( .A(n50), .B(n3288), .Z(n3286) );
  XOR U3965 ( .A(n3289), .B(n3287), .Z(n3288) );
  XNOR U3966 ( .A(n3290), .B(n3291), .Z(n3278) );
  NAND U3967 ( .A(n3292), .B(n3293), .Z(n3291) );
  XOR U3968 ( .A(n3294), .B(n3270), .Z(n3293) );
  XOR U3969 ( .A(n3284), .B(n3285), .Z(n3270) );
  XOR U3970 ( .A(n3295), .B(n3296), .Z(n3285) );
  ANDN U3971 ( .B(n3297), .A(n3298), .Z(n3295) );
  XOR U3972 ( .A(n3296), .B(n3299), .Z(n3297) );
  XOR U3973 ( .A(n3300), .B(n3301), .Z(n3284) );
  XOR U3974 ( .A(n3302), .B(n3303), .Z(n3301) );
  ANDN U3975 ( .B(n3304), .A(n3305), .Z(n3302) );
  XOR U3976 ( .A(n3306), .B(n3303), .Z(n3304) );
  IV U3977 ( .A(n3282), .Z(n3300) );
  XOR U3978 ( .A(n3307), .B(n3308), .Z(n3282) );
  ANDN U3979 ( .B(n3309), .A(n3310), .Z(n3307) );
  XOR U3980 ( .A(n3308), .B(n3311), .Z(n3309) );
  IV U3981 ( .A(n3290), .Z(n3294) );
  XOR U3982 ( .A(n3290), .B(n3272), .Z(n3292) );
  XOR U3983 ( .A(n3312), .B(n3313), .Z(n3272) );
  AND U3984 ( .A(n50), .B(n3314), .Z(n3312) );
  XOR U3985 ( .A(n3315), .B(n3313), .Z(n3314) );
  NANDN U3986 ( .A(n3274), .B(n3276), .Z(n3290) );
  XOR U3987 ( .A(n3316), .B(n3317), .Z(n3276) );
  AND U3988 ( .A(n50), .B(n3318), .Z(n3316) );
  XOR U3989 ( .A(n3317), .B(n3319), .Z(n3318) );
  XOR U3990 ( .A(n3320), .B(n3321), .Z(n50) );
  AND U3991 ( .A(n3322), .B(n3323), .Z(n3320) );
  XNOR U3992 ( .A(n3321), .B(n3287), .Z(n3323) );
  XNOR U3993 ( .A(n3324), .B(n3325), .Z(n3287) );
  ANDN U3994 ( .B(n3326), .A(n3327), .Z(n3324) );
  XOR U3995 ( .A(n3325), .B(n3328), .Z(n3326) );
  XOR U3996 ( .A(n3321), .B(n3289), .Z(n3322) );
  XOR U3997 ( .A(n3329), .B(n3330), .Z(n3289) );
  AND U3998 ( .A(n54), .B(n3331), .Z(n3329) );
  XOR U3999 ( .A(n3332), .B(n3330), .Z(n3331) );
  XNOR U4000 ( .A(n3333), .B(n3334), .Z(n3321) );
  NAND U4001 ( .A(n3335), .B(n3336), .Z(n3334) );
  XOR U4002 ( .A(n3337), .B(n3313), .Z(n3336) );
  XOR U4003 ( .A(n3327), .B(n3328), .Z(n3313) );
  XOR U4004 ( .A(n3338), .B(n3339), .Z(n3328) );
  ANDN U4005 ( .B(n3340), .A(n3341), .Z(n3338) );
  XOR U4006 ( .A(n3339), .B(n3342), .Z(n3340) );
  XOR U4007 ( .A(n3343), .B(n3344), .Z(n3327) );
  XOR U4008 ( .A(n3345), .B(n3346), .Z(n3344) );
  ANDN U4009 ( .B(n3347), .A(n3348), .Z(n3345) );
  XOR U4010 ( .A(n3349), .B(n3346), .Z(n3347) );
  IV U4011 ( .A(n3325), .Z(n3343) );
  XOR U4012 ( .A(n3350), .B(n3351), .Z(n3325) );
  ANDN U4013 ( .B(n3352), .A(n3353), .Z(n3350) );
  XOR U4014 ( .A(n3351), .B(n3354), .Z(n3352) );
  IV U4015 ( .A(n3333), .Z(n3337) );
  XOR U4016 ( .A(n3333), .B(n3315), .Z(n3335) );
  XOR U4017 ( .A(n3355), .B(n3356), .Z(n3315) );
  AND U4018 ( .A(n54), .B(n3357), .Z(n3355) );
  XOR U4019 ( .A(n3358), .B(n3356), .Z(n3357) );
  NANDN U4020 ( .A(n3317), .B(n3319), .Z(n3333) );
  XOR U4021 ( .A(n3359), .B(n3360), .Z(n3319) );
  AND U4022 ( .A(n54), .B(n3361), .Z(n3359) );
  XOR U4023 ( .A(n3360), .B(n3362), .Z(n3361) );
  XOR U4024 ( .A(n3363), .B(n3364), .Z(n54) );
  AND U4025 ( .A(n3365), .B(n3366), .Z(n3363) );
  XNOR U4026 ( .A(n3364), .B(n3330), .Z(n3366) );
  XNOR U4027 ( .A(n3367), .B(n3368), .Z(n3330) );
  ANDN U4028 ( .B(n3369), .A(n3370), .Z(n3367) );
  XOR U4029 ( .A(n3368), .B(n3371), .Z(n3369) );
  XOR U4030 ( .A(n3364), .B(n3332), .Z(n3365) );
  XOR U4031 ( .A(n3372), .B(n3373), .Z(n3332) );
  AND U4032 ( .A(n58), .B(n3374), .Z(n3372) );
  XOR U4033 ( .A(n3375), .B(n3373), .Z(n3374) );
  XNOR U4034 ( .A(n3376), .B(n3377), .Z(n3364) );
  NAND U4035 ( .A(n3378), .B(n3379), .Z(n3377) );
  XOR U4036 ( .A(n3380), .B(n3356), .Z(n3379) );
  XOR U4037 ( .A(n3370), .B(n3371), .Z(n3356) );
  XOR U4038 ( .A(n3381), .B(n3382), .Z(n3371) );
  ANDN U4039 ( .B(n3383), .A(n3384), .Z(n3381) );
  XOR U4040 ( .A(n3382), .B(n3385), .Z(n3383) );
  XOR U4041 ( .A(n3386), .B(n3387), .Z(n3370) );
  XOR U4042 ( .A(n3388), .B(n3389), .Z(n3387) );
  ANDN U4043 ( .B(n3390), .A(n3391), .Z(n3388) );
  XOR U4044 ( .A(n3392), .B(n3389), .Z(n3390) );
  IV U4045 ( .A(n3368), .Z(n3386) );
  XOR U4046 ( .A(n3393), .B(n3394), .Z(n3368) );
  ANDN U4047 ( .B(n3395), .A(n3396), .Z(n3393) );
  XOR U4048 ( .A(n3394), .B(n3397), .Z(n3395) );
  IV U4049 ( .A(n3376), .Z(n3380) );
  XOR U4050 ( .A(n3376), .B(n3358), .Z(n3378) );
  XOR U4051 ( .A(n3398), .B(n3399), .Z(n3358) );
  AND U4052 ( .A(n58), .B(n3400), .Z(n3398) );
  XOR U4053 ( .A(n3401), .B(n3399), .Z(n3400) );
  NANDN U4054 ( .A(n3360), .B(n3362), .Z(n3376) );
  XOR U4055 ( .A(n3402), .B(n3403), .Z(n3362) );
  AND U4056 ( .A(n58), .B(n3404), .Z(n3402) );
  XOR U4057 ( .A(n3403), .B(n3405), .Z(n3404) );
  XOR U4058 ( .A(n3406), .B(n3407), .Z(n58) );
  AND U4059 ( .A(n3408), .B(n3409), .Z(n3406) );
  XNOR U4060 ( .A(n3407), .B(n3373), .Z(n3409) );
  XNOR U4061 ( .A(n3410), .B(n3411), .Z(n3373) );
  ANDN U4062 ( .B(n3412), .A(n3413), .Z(n3410) );
  XOR U4063 ( .A(n3411), .B(n3414), .Z(n3412) );
  XOR U4064 ( .A(n3407), .B(n3375), .Z(n3408) );
  XOR U4065 ( .A(n3415), .B(n3416), .Z(n3375) );
  AND U4066 ( .A(n62), .B(n3417), .Z(n3415) );
  XOR U4067 ( .A(n3418), .B(n3416), .Z(n3417) );
  XNOR U4068 ( .A(n3419), .B(n3420), .Z(n3407) );
  NAND U4069 ( .A(n3421), .B(n3422), .Z(n3420) );
  XOR U4070 ( .A(n3423), .B(n3399), .Z(n3422) );
  XOR U4071 ( .A(n3413), .B(n3414), .Z(n3399) );
  XOR U4072 ( .A(n3424), .B(n3425), .Z(n3414) );
  ANDN U4073 ( .B(n3426), .A(n3427), .Z(n3424) );
  XOR U4074 ( .A(n3425), .B(n3428), .Z(n3426) );
  XOR U4075 ( .A(n3429), .B(n3430), .Z(n3413) );
  XOR U4076 ( .A(n3431), .B(n3432), .Z(n3430) );
  ANDN U4077 ( .B(n3433), .A(n3434), .Z(n3431) );
  XOR U4078 ( .A(n3435), .B(n3432), .Z(n3433) );
  IV U4079 ( .A(n3411), .Z(n3429) );
  XOR U4080 ( .A(n3436), .B(n3437), .Z(n3411) );
  ANDN U4081 ( .B(n3438), .A(n3439), .Z(n3436) );
  XOR U4082 ( .A(n3437), .B(n3440), .Z(n3438) );
  IV U4083 ( .A(n3419), .Z(n3423) );
  XOR U4084 ( .A(n3419), .B(n3401), .Z(n3421) );
  XOR U4085 ( .A(n3441), .B(n3442), .Z(n3401) );
  AND U4086 ( .A(n62), .B(n3443), .Z(n3441) );
  XOR U4087 ( .A(n3444), .B(n3442), .Z(n3443) );
  NANDN U4088 ( .A(n3403), .B(n3405), .Z(n3419) );
  XOR U4089 ( .A(n3445), .B(n3446), .Z(n3405) );
  AND U4090 ( .A(n62), .B(n3447), .Z(n3445) );
  XOR U4091 ( .A(n3446), .B(n3448), .Z(n3447) );
  XOR U4092 ( .A(n3449), .B(n3450), .Z(n62) );
  AND U4093 ( .A(n3451), .B(n3452), .Z(n3449) );
  XNOR U4094 ( .A(n3450), .B(n3416), .Z(n3452) );
  XNOR U4095 ( .A(n3453), .B(n3454), .Z(n3416) );
  ANDN U4096 ( .B(n3455), .A(n3456), .Z(n3453) );
  XOR U4097 ( .A(n3454), .B(n3457), .Z(n3455) );
  XOR U4098 ( .A(n3450), .B(n3418), .Z(n3451) );
  XOR U4099 ( .A(n3458), .B(n3459), .Z(n3418) );
  AND U4100 ( .A(n66), .B(n3460), .Z(n3458) );
  XOR U4101 ( .A(n3461), .B(n3459), .Z(n3460) );
  XNOR U4102 ( .A(n3462), .B(n3463), .Z(n3450) );
  NAND U4103 ( .A(n3464), .B(n3465), .Z(n3463) );
  XOR U4104 ( .A(n3466), .B(n3442), .Z(n3465) );
  XOR U4105 ( .A(n3456), .B(n3457), .Z(n3442) );
  XOR U4106 ( .A(n3467), .B(n3468), .Z(n3457) );
  ANDN U4107 ( .B(n3469), .A(n3470), .Z(n3467) );
  XOR U4108 ( .A(n3468), .B(n3471), .Z(n3469) );
  XOR U4109 ( .A(n3472), .B(n3473), .Z(n3456) );
  XOR U4110 ( .A(n3474), .B(n3475), .Z(n3473) );
  ANDN U4111 ( .B(n3476), .A(n3477), .Z(n3474) );
  XOR U4112 ( .A(n3478), .B(n3475), .Z(n3476) );
  IV U4113 ( .A(n3454), .Z(n3472) );
  XOR U4114 ( .A(n3479), .B(n3480), .Z(n3454) );
  ANDN U4115 ( .B(n3481), .A(n3482), .Z(n3479) );
  XOR U4116 ( .A(n3480), .B(n3483), .Z(n3481) );
  IV U4117 ( .A(n3462), .Z(n3466) );
  XOR U4118 ( .A(n3462), .B(n3444), .Z(n3464) );
  XOR U4119 ( .A(n3484), .B(n3485), .Z(n3444) );
  AND U4120 ( .A(n66), .B(n3486), .Z(n3484) );
  XOR U4121 ( .A(n3487), .B(n3485), .Z(n3486) );
  NANDN U4122 ( .A(n3446), .B(n3448), .Z(n3462) );
  XOR U4123 ( .A(n3488), .B(n3489), .Z(n3448) );
  AND U4124 ( .A(n66), .B(n3490), .Z(n3488) );
  XOR U4125 ( .A(n3489), .B(n3491), .Z(n3490) );
  XOR U4126 ( .A(n3492), .B(n3493), .Z(n66) );
  AND U4127 ( .A(n3494), .B(n3495), .Z(n3492) );
  XNOR U4128 ( .A(n3493), .B(n3459), .Z(n3495) );
  XNOR U4129 ( .A(n3496), .B(n3497), .Z(n3459) );
  ANDN U4130 ( .B(n3498), .A(n3499), .Z(n3496) );
  XOR U4131 ( .A(n3497), .B(n3500), .Z(n3498) );
  XOR U4132 ( .A(n3493), .B(n3461), .Z(n3494) );
  XOR U4133 ( .A(n3501), .B(n3502), .Z(n3461) );
  AND U4134 ( .A(n70), .B(n3503), .Z(n3501) );
  XOR U4135 ( .A(n3504), .B(n3502), .Z(n3503) );
  XNOR U4136 ( .A(n3505), .B(n3506), .Z(n3493) );
  NAND U4137 ( .A(n3507), .B(n3508), .Z(n3506) );
  XOR U4138 ( .A(n3509), .B(n3485), .Z(n3508) );
  XOR U4139 ( .A(n3499), .B(n3500), .Z(n3485) );
  XOR U4140 ( .A(n3510), .B(n3511), .Z(n3500) );
  ANDN U4141 ( .B(n3512), .A(n3513), .Z(n3510) );
  XOR U4142 ( .A(n3511), .B(n3514), .Z(n3512) );
  XOR U4143 ( .A(n3515), .B(n3516), .Z(n3499) );
  XOR U4144 ( .A(n3517), .B(n3518), .Z(n3516) );
  ANDN U4145 ( .B(n3519), .A(n3520), .Z(n3517) );
  XOR U4146 ( .A(n3521), .B(n3518), .Z(n3519) );
  IV U4147 ( .A(n3497), .Z(n3515) );
  XOR U4148 ( .A(n3522), .B(n3523), .Z(n3497) );
  ANDN U4149 ( .B(n3524), .A(n3525), .Z(n3522) );
  XOR U4150 ( .A(n3523), .B(n3526), .Z(n3524) );
  IV U4151 ( .A(n3505), .Z(n3509) );
  XOR U4152 ( .A(n3505), .B(n3487), .Z(n3507) );
  XOR U4153 ( .A(n3527), .B(n3528), .Z(n3487) );
  AND U4154 ( .A(n70), .B(n3529), .Z(n3527) );
  XOR U4155 ( .A(n3530), .B(n3528), .Z(n3529) );
  NANDN U4156 ( .A(n3489), .B(n3491), .Z(n3505) );
  XOR U4157 ( .A(n3531), .B(n3532), .Z(n3491) );
  AND U4158 ( .A(n70), .B(n3533), .Z(n3531) );
  XOR U4159 ( .A(n3532), .B(n3534), .Z(n3533) );
  XOR U4160 ( .A(n3535), .B(n3536), .Z(n70) );
  AND U4161 ( .A(n3537), .B(n3538), .Z(n3535) );
  XNOR U4162 ( .A(n3536), .B(n3502), .Z(n3538) );
  XNOR U4163 ( .A(n3539), .B(n3540), .Z(n3502) );
  ANDN U4164 ( .B(n3541), .A(n3542), .Z(n3539) );
  XOR U4165 ( .A(n3540), .B(n3543), .Z(n3541) );
  XOR U4166 ( .A(n3536), .B(n3504), .Z(n3537) );
  XOR U4167 ( .A(n3544), .B(n3545), .Z(n3504) );
  AND U4168 ( .A(n74), .B(n3546), .Z(n3544) );
  XOR U4169 ( .A(n3547), .B(n3545), .Z(n3546) );
  XNOR U4170 ( .A(n3548), .B(n3549), .Z(n3536) );
  NAND U4171 ( .A(n3550), .B(n3551), .Z(n3549) );
  XOR U4172 ( .A(n3552), .B(n3528), .Z(n3551) );
  XOR U4173 ( .A(n3542), .B(n3543), .Z(n3528) );
  XOR U4174 ( .A(n3553), .B(n3554), .Z(n3543) );
  ANDN U4175 ( .B(n3555), .A(n3556), .Z(n3553) );
  XOR U4176 ( .A(n3554), .B(n3557), .Z(n3555) );
  XOR U4177 ( .A(n3558), .B(n3559), .Z(n3542) );
  XOR U4178 ( .A(n3560), .B(n3561), .Z(n3559) );
  ANDN U4179 ( .B(n3562), .A(n3563), .Z(n3560) );
  XOR U4180 ( .A(n3564), .B(n3561), .Z(n3562) );
  IV U4181 ( .A(n3540), .Z(n3558) );
  XOR U4182 ( .A(n3565), .B(n3566), .Z(n3540) );
  ANDN U4183 ( .B(n3567), .A(n3568), .Z(n3565) );
  XOR U4184 ( .A(n3566), .B(n3569), .Z(n3567) );
  IV U4185 ( .A(n3548), .Z(n3552) );
  XOR U4186 ( .A(n3548), .B(n3530), .Z(n3550) );
  XOR U4187 ( .A(n3570), .B(n3571), .Z(n3530) );
  AND U4188 ( .A(n74), .B(n3572), .Z(n3570) );
  XOR U4189 ( .A(n3573), .B(n3571), .Z(n3572) );
  NANDN U4190 ( .A(n3532), .B(n3534), .Z(n3548) );
  XOR U4191 ( .A(n3574), .B(n3575), .Z(n3534) );
  AND U4192 ( .A(n74), .B(n3576), .Z(n3574) );
  XOR U4193 ( .A(n3575), .B(n3577), .Z(n3576) );
  XOR U4194 ( .A(n3578), .B(n3579), .Z(n74) );
  AND U4195 ( .A(n3580), .B(n3581), .Z(n3578) );
  XNOR U4196 ( .A(n3579), .B(n3545), .Z(n3581) );
  XNOR U4197 ( .A(n3582), .B(n3583), .Z(n3545) );
  ANDN U4198 ( .B(n3584), .A(n3585), .Z(n3582) );
  XOR U4199 ( .A(n3583), .B(n3586), .Z(n3584) );
  XOR U4200 ( .A(n3579), .B(n3547), .Z(n3580) );
  XOR U4201 ( .A(n3587), .B(n3588), .Z(n3547) );
  AND U4202 ( .A(n78), .B(n3589), .Z(n3587) );
  XOR U4203 ( .A(n3590), .B(n3588), .Z(n3589) );
  XNOR U4204 ( .A(n3591), .B(n3592), .Z(n3579) );
  NAND U4205 ( .A(n3593), .B(n3594), .Z(n3592) );
  XOR U4206 ( .A(n3595), .B(n3571), .Z(n3594) );
  XOR U4207 ( .A(n3585), .B(n3586), .Z(n3571) );
  XOR U4208 ( .A(n3596), .B(n3597), .Z(n3586) );
  ANDN U4209 ( .B(n3598), .A(n3599), .Z(n3596) );
  XOR U4210 ( .A(n3597), .B(n3600), .Z(n3598) );
  XOR U4211 ( .A(n3601), .B(n3602), .Z(n3585) );
  XOR U4212 ( .A(n3603), .B(n3604), .Z(n3602) );
  ANDN U4213 ( .B(n3605), .A(n3606), .Z(n3603) );
  XOR U4214 ( .A(n3607), .B(n3604), .Z(n3605) );
  IV U4215 ( .A(n3583), .Z(n3601) );
  XOR U4216 ( .A(n3608), .B(n3609), .Z(n3583) );
  ANDN U4217 ( .B(n3610), .A(n3611), .Z(n3608) );
  XOR U4218 ( .A(n3609), .B(n3612), .Z(n3610) );
  IV U4219 ( .A(n3591), .Z(n3595) );
  XOR U4220 ( .A(n3591), .B(n3573), .Z(n3593) );
  XOR U4221 ( .A(n3613), .B(n3614), .Z(n3573) );
  AND U4222 ( .A(n78), .B(n3615), .Z(n3613) );
  XOR U4223 ( .A(n3616), .B(n3614), .Z(n3615) );
  NANDN U4224 ( .A(n3575), .B(n3577), .Z(n3591) );
  XOR U4225 ( .A(n3617), .B(n3618), .Z(n3577) );
  AND U4226 ( .A(n78), .B(n3619), .Z(n3617) );
  XOR U4227 ( .A(n3618), .B(n3620), .Z(n3619) );
  XOR U4228 ( .A(n3621), .B(n3622), .Z(n78) );
  AND U4229 ( .A(n3623), .B(n3624), .Z(n3621) );
  XNOR U4230 ( .A(n3622), .B(n3588), .Z(n3624) );
  XNOR U4231 ( .A(n3625), .B(n3626), .Z(n3588) );
  ANDN U4232 ( .B(n3627), .A(n3628), .Z(n3625) );
  XOR U4233 ( .A(n3626), .B(n3629), .Z(n3627) );
  XOR U4234 ( .A(n3622), .B(n3590), .Z(n3623) );
  XOR U4235 ( .A(n3630), .B(n3631), .Z(n3590) );
  AND U4236 ( .A(n82), .B(n3632), .Z(n3630) );
  XOR U4237 ( .A(n3633), .B(n3631), .Z(n3632) );
  XNOR U4238 ( .A(n3634), .B(n3635), .Z(n3622) );
  NAND U4239 ( .A(n3636), .B(n3637), .Z(n3635) );
  XOR U4240 ( .A(n3638), .B(n3614), .Z(n3637) );
  XOR U4241 ( .A(n3628), .B(n3629), .Z(n3614) );
  XOR U4242 ( .A(n3639), .B(n3640), .Z(n3629) );
  ANDN U4243 ( .B(n3641), .A(n3642), .Z(n3639) );
  XOR U4244 ( .A(n3640), .B(n3643), .Z(n3641) );
  XOR U4245 ( .A(n3644), .B(n3645), .Z(n3628) );
  XOR U4246 ( .A(n3646), .B(n3647), .Z(n3645) );
  ANDN U4247 ( .B(n3648), .A(n3649), .Z(n3646) );
  XOR U4248 ( .A(n3650), .B(n3647), .Z(n3648) );
  IV U4249 ( .A(n3626), .Z(n3644) );
  XOR U4250 ( .A(n3651), .B(n3652), .Z(n3626) );
  ANDN U4251 ( .B(n3653), .A(n3654), .Z(n3651) );
  XOR U4252 ( .A(n3652), .B(n3655), .Z(n3653) );
  IV U4253 ( .A(n3634), .Z(n3638) );
  XOR U4254 ( .A(n3634), .B(n3616), .Z(n3636) );
  XOR U4255 ( .A(n3656), .B(n3657), .Z(n3616) );
  AND U4256 ( .A(n82), .B(n3658), .Z(n3656) );
  XOR U4257 ( .A(n3659), .B(n3657), .Z(n3658) );
  NANDN U4258 ( .A(n3618), .B(n3620), .Z(n3634) );
  XOR U4259 ( .A(n3660), .B(n3661), .Z(n3620) );
  AND U4260 ( .A(n82), .B(n3662), .Z(n3660) );
  XOR U4261 ( .A(n3661), .B(n3663), .Z(n3662) );
  XOR U4262 ( .A(n3664), .B(n3665), .Z(n82) );
  AND U4263 ( .A(n3666), .B(n3667), .Z(n3664) );
  XNOR U4264 ( .A(n3665), .B(n3631), .Z(n3667) );
  XNOR U4265 ( .A(n3668), .B(n3669), .Z(n3631) );
  ANDN U4266 ( .B(n3670), .A(n3671), .Z(n3668) );
  XOR U4267 ( .A(n3669), .B(n3672), .Z(n3670) );
  XOR U4268 ( .A(n3665), .B(n3633), .Z(n3666) );
  XOR U4269 ( .A(n3673), .B(n3674), .Z(n3633) );
  AND U4270 ( .A(n86), .B(n3675), .Z(n3673) );
  XOR U4271 ( .A(n3676), .B(n3674), .Z(n3675) );
  XNOR U4272 ( .A(n3677), .B(n3678), .Z(n3665) );
  NAND U4273 ( .A(n3679), .B(n3680), .Z(n3678) );
  XOR U4274 ( .A(n3681), .B(n3657), .Z(n3680) );
  XOR U4275 ( .A(n3671), .B(n3672), .Z(n3657) );
  XOR U4276 ( .A(n3682), .B(n3683), .Z(n3672) );
  ANDN U4277 ( .B(n3684), .A(n3685), .Z(n3682) );
  XOR U4278 ( .A(n3683), .B(n3686), .Z(n3684) );
  XOR U4279 ( .A(n3687), .B(n3688), .Z(n3671) );
  XOR U4280 ( .A(n3689), .B(n3690), .Z(n3688) );
  ANDN U4281 ( .B(n3691), .A(n3692), .Z(n3689) );
  XOR U4282 ( .A(n3693), .B(n3690), .Z(n3691) );
  IV U4283 ( .A(n3669), .Z(n3687) );
  XOR U4284 ( .A(n3694), .B(n3695), .Z(n3669) );
  ANDN U4285 ( .B(n3696), .A(n3697), .Z(n3694) );
  XOR U4286 ( .A(n3695), .B(n3698), .Z(n3696) );
  IV U4287 ( .A(n3677), .Z(n3681) );
  XOR U4288 ( .A(n3677), .B(n3659), .Z(n3679) );
  XOR U4289 ( .A(n3699), .B(n3700), .Z(n3659) );
  AND U4290 ( .A(n86), .B(n3701), .Z(n3699) );
  XOR U4291 ( .A(n3702), .B(n3700), .Z(n3701) );
  NANDN U4292 ( .A(n3661), .B(n3663), .Z(n3677) );
  XOR U4293 ( .A(n3703), .B(n3704), .Z(n3663) );
  AND U4294 ( .A(n86), .B(n3705), .Z(n3703) );
  XOR U4295 ( .A(n3704), .B(n3706), .Z(n3705) );
  XOR U4296 ( .A(n3707), .B(n3708), .Z(n86) );
  AND U4297 ( .A(n3709), .B(n3710), .Z(n3707) );
  XNOR U4298 ( .A(n3708), .B(n3674), .Z(n3710) );
  XNOR U4299 ( .A(n3711), .B(n3712), .Z(n3674) );
  ANDN U4300 ( .B(n3713), .A(n3714), .Z(n3711) );
  XOR U4301 ( .A(n3712), .B(n3715), .Z(n3713) );
  XOR U4302 ( .A(n3708), .B(n3676), .Z(n3709) );
  XOR U4303 ( .A(n3716), .B(n3717), .Z(n3676) );
  AND U4304 ( .A(n90), .B(n3718), .Z(n3716) );
  XOR U4305 ( .A(n3719), .B(n3717), .Z(n3718) );
  XNOR U4306 ( .A(n3720), .B(n3721), .Z(n3708) );
  NAND U4307 ( .A(n3722), .B(n3723), .Z(n3721) );
  XOR U4308 ( .A(n3724), .B(n3700), .Z(n3723) );
  XOR U4309 ( .A(n3714), .B(n3715), .Z(n3700) );
  XOR U4310 ( .A(n3725), .B(n3726), .Z(n3715) );
  ANDN U4311 ( .B(n3727), .A(n3728), .Z(n3725) );
  XOR U4312 ( .A(n3726), .B(n3729), .Z(n3727) );
  XOR U4313 ( .A(n3730), .B(n3731), .Z(n3714) );
  XOR U4314 ( .A(n3732), .B(n3733), .Z(n3731) );
  ANDN U4315 ( .B(n3734), .A(n3735), .Z(n3732) );
  XOR U4316 ( .A(n3736), .B(n3733), .Z(n3734) );
  IV U4317 ( .A(n3712), .Z(n3730) );
  XOR U4318 ( .A(n3737), .B(n3738), .Z(n3712) );
  ANDN U4319 ( .B(n3739), .A(n3740), .Z(n3737) );
  XOR U4320 ( .A(n3738), .B(n3741), .Z(n3739) );
  IV U4321 ( .A(n3720), .Z(n3724) );
  XOR U4322 ( .A(n3720), .B(n3702), .Z(n3722) );
  XOR U4323 ( .A(n3742), .B(n3743), .Z(n3702) );
  AND U4324 ( .A(n90), .B(n3744), .Z(n3742) );
  XOR U4325 ( .A(n3745), .B(n3743), .Z(n3744) );
  NANDN U4326 ( .A(n3704), .B(n3706), .Z(n3720) );
  XOR U4327 ( .A(n3746), .B(n3747), .Z(n3706) );
  AND U4328 ( .A(n90), .B(n3748), .Z(n3746) );
  XOR U4329 ( .A(n3747), .B(n3749), .Z(n3748) );
  XOR U4330 ( .A(n3750), .B(n3751), .Z(n90) );
  AND U4331 ( .A(n3752), .B(n3753), .Z(n3750) );
  XNOR U4332 ( .A(n3751), .B(n3717), .Z(n3753) );
  XNOR U4333 ( .A(n3754), .B(n3755), .Z(n3717) );
  ANDN U4334 ( .B(n3756), .A(n3757), .Z(n3754) );
  XOR U4335 ( .A(n3755), .B(n3758), .Z(n3756) );
  XOR U4336 ( .A(n3751), .B(n3719), .Z(n3752) );
  XOR U4337 ( .A(n3759), .B(n3760), .Z(n3719) );
  AND U4338 ( .A(n94), .B(n3761), .Z(n3759) );
  XOR U4339 ( .A(n3762), .B(n3760), .Z(n3761) );
  XNOR U4340 ( .A(n3763), .B(n3764), .Z(n3751) );
  NAND U4341 ( .A(n3765), .B(n3766), .Z(n3764) );
  XOR U4342 ( .A(n3767), .B(n3743), .Z(n3766) );
  XOR U4343 ( .A(n3757), .B(n3758), .Z(n3743) );
  XOR U4344 ( .A(n3768), .B(n3769), .Z(n3758) );
  ANDN U4345 ( .B(n3770), .A(n3771), .Z(n3768) );
  XOR U4346 ( .A(n3769), .B(n3772), .Z(n3770) );
  XOR U4347 ( .A(n3773), .B(n3774), .Z(n3757) );
  XOR U4348 ( .A(n3775), .B(n3776), .Z(n3774) );
  ANDN U4349 ( .B(n3777), .A(n3778), .Z(n3775) );
  XOR U4350 ( .A(n3779), .B(n3776), .Z(n3777) );
  IV U4351 ( .A(n3755), .Z(n3773) );
  XOR U4352 ( .A(n3780), .B(n3781), .Z(n3755) );
  ANDN U4353 ( .B(n3782), .A(n3783), .Z(n3780) );
  XOR U4354 ( .A(n3781), .B(n3784), .Z(n3782) );
  IV U4355 ( .A(n3763), .Z(n3767) );
  XOR U4356 ( .A(n3763), .B(n3745), .Z(n3765) );
  XOR U4357 ( .A(n3785), .B(n3786), .Z(n3745) );
  AND U4358 ( .A(n94), .B(n3787), .Z(n3785) );
  XOR U4359 ( .A(n3788), .B(n3786), .Z(n3787) );
  NANDN U4360 ( .A(n3747), .B(n3749), .Z(n3763) );
  XOR U4361 ( .A(n3789), .B(n3790), .Z(n3749) );
  AND U4362 ( .A(n94), .B(n3791), .Z(n3789) );
  XOR U4363 ( .A(n3790), .B(n3792), .Z(n3791) );
  XOR U4364 ( .A(n3793), .B(n3794), .Z(n94) );
  AND U4365 ( .A(n3795), .B(n3796), .Z(n3793) );
  XNOR U4366 ( .A(n3794), .B(n3760), .Z(n3796) );
  XNOR U4367 ( .A(n3797), .B(n3798), .Z(n3760) );
  ANDN U4368 ( .B(n3799), .A(n3800), .Z(n3797) );
  XOR U4369 ( .A(n3798), .B(n3801), .Z(n3799) );
  XOR U4370 ( .A(n3794), .B(n3762), .Z(n3795) );
  XOR U4371 ( .A(n3802), .B(n3803), .Z(n3762) );
  AND U4372 ( .A(n98), .B(n3804), .Z(n3802) );
  XOR U4373 ( .A(n3805), .B(n3803), .Z(n3804) );
  XNOR U4374 ( .A(n3806), .B(n3807), .Z(n3794) );
  NAND U4375 ( .A(n3808), .B(n3809), .Z(n3807) );
  XOR U4376 ( .A(n3810), .B(n3786), .Z(n3809) );
  XOR U4377 ( .A(n3800), .B(n3801), .Z(n3786) );
  XOR U4378 ( .A(n3811), .B(n3812), .Z(n3801) );
  ANDN U4379 ( .B(n3813), .A(n3814), .Z(n3811) );
  XOR U4380 ( .A(n3812), .B(n3815), .Z(n3813) );
  XOR U4381 ( .A(n3816), .B(n3817), .Z(n3800) );
  XOR U4382 ( .A(n3818), .B(n3819), .Z(n3817) );
  ANDN U4383 ( .B(n3820), .A(n3821), .Z(n3818) );
  XOR U4384 ( .A(n3822), .B(n3819), .Z(n3820) );
  IV U4385 ( .A(n3798), .Z(n3816) );
  XOR U4386 ( .A(n3823), .B(n3824), .Z(n3798) );
  ANDN U4387 ( .B(n3825), .A(n3826), .Z(n3823) );
  XOR U4388 ( .A(n3824), .B(n3827), .Z(n3825) );
  IV U4389 ( .A(n3806), .Z(n3810) );
  XOR U4390 ( .A(n3806), .B(n3788), .Z(n3808) );
  XOR U4391 ( .A(n3828), .B(n3829), .Z(n3788) );
  AND U4392 ( .A(n98), .B(n3830), .Z(n3828) );
  XOR U4393 ( .A(n3831), .B(n3829), .Z(n3830) );
  NANDN U4394 ( .A(n3790), .B(n3792), .Z(n3806) );
  XOR U4395 ( .A(n3832), .B(n3833), .Z(n3792) );
  AND U4396 ( .A(n98), .B(n3834), .Z(n3832) );
  XOR U4397 ( .A(n3833), .B(n3835), .Z(n3834) );
  XOR U4398 ( .A(n3836), .B(n3837), .Z(n98) );
  AND U4399 ( .A(n3838), .B(n3839), .Z(n3836) );
  XNOR U4400 ( .A(n3837), .B(n3803), .Z(n3839) );
  XNOR U4401 ( .A(n3840), .B(n3841), .Z(n3803) );
  ANDN U4402 ( .B(n3842), .A(n3843), .Z(n3840) );
  XOR U4403 ( .A(n3841), .B(n3844), .Z(n3842) );
  XOR U4404 ( .A(n3837), .B(n3805), .Z(n3838) );
  XOR U4405 ( .A(n3845), .B(n3846), .Z(n3805) );
  AND U4406 ( .A(n102), .B(n3847), .Z(n3845) );
  XOR U4407 ( .A(n3848), .B(n3846), .Z(n3847) );
  XNOR U4408 ( .A(n3849), .B(n3850), .Z(n3837) );
  NAND U4409 ( .A(n3851), .B(n3852), .Z(n3850) );
  XOR U4410 ( .A(n3853), .B(n3829), .Z(n3852) );
  XOR U4411 ( .A(n3843), .B(n3844), .Z(n3829) );
  XOR U4412 ( .A(n3854), .B(n3855), .Z(n3844) );
  ANDN U4413 ( .B(n3856), .A(n3857), .Z(n3854) );
  XOR U4414 ( .A(n3855), .B(n3858), .Z(n3856) );
  XOR U4415 ( .A(n3859), .B(n3860), .Z(n3843) );
  XOR U4416 ( .A(n3861), .B(n3862), .Z(n3860) );
  ANDN U4417 ( .B(n3863), .A(n3864), .Z(n3861) );
  XOR U4418 ( .A(n3865), .B(n3862), .Z(n3863) );
  IV U4419 ( .A(n3841), .Z(n3859) );
  XOR U4420 ( .A(n3866), .B(n3867), .Z(n3841) );
  ANDN U4421 ( .B(n3868), .A(n3869), .Z(n3866) );
  XOR U4422 ( .A(n3867), .B(n3870), .Z(n3868) );
  IV U4423 ( .A(n3849), .Z(n3853) );
  XOR U4424 ( .A(n3849), .B(n3831), .Z(n3851) );
  XOR U4425 ( .A(n3871), .B(n3872), .Z(n3831) );
  AND U4426 ( .A(n102), .B(n3873), .Z(n3871) );
  XOR U4427 ( .A(n3874), .B(n3872), .Z(n3873) );
  NANDN U4428 ( .A(n3833), .B(n3835), .Z(n3849) );
  XOR U4429 ( .A(n3875), .B(n3876), .Z(n3835) );
  AND U4430 ( .A(n102), .B(n3877), .Z(n3875) );
  XOR U4431 ( .A(n3876), .B(n3878), .Z(n3877) );
  XOR U4432 ( .A(n3879), .B(n3880), .Z(n102) );
  AND U4433 ( .A(n3881), .B(n3882), .Z(n3879) );
  XNOR U4434 ( .A(n3880), .B(n3846), .Z(n3882) );
  XNOR U4435 ( .A(n3883), .B(n3884), .Z(n3846) );
  ANDN U4436 ( .B(n3885), .A(n3886), .Z(n3883) );
  XOR U4437 ( .A(n3884), .B(n3887), .Z(n3885) );
  XOR U4438 ( .A(n3880), .B(n3848), .Z(n3881) );
  XOR U4439 ( .A(n3888), .B(n3889), .Z(n3848) );
  AND U4440 ( .A(n106), .B(n3890), .Z(n3888) );
  XOR U4441 ( .A(n3891), .B(n3889), .Z(n3890) );
  XNOR U4442 ( .A(n3892), .B(n3893), .Z(n3880) );
  NAND U4443 ( .A(n3894), .B(n3895), .Z(n3893) );
  XOR U4444 ( .A(n3896), .B(n3872), .Z(n3895) );
  XOR U4445 ( .A(n3886), .B(n3887), .Z(n3872) );
  XOR U4446 ( .A(n3897), .B(n3898), .Z(n3887) );
  ANDN U4447 ( .B(n3899), .A(n3900), .Z(n3897) );
  XOR U4448 ( .A(n3898), .B(n3901), .Z(n3899) );
  XOR U4449 ( .A(n3902), .B(n3903), .Z(n3886) );
  XOR U4450 ( .A(n3904), .B(n3905), .Z(n3903) );
  ANDN U4451 ( .B(n3906), .A(n3907), .Z(n3904) );
  XOR U4452 ( .A(n3908), .B(n3905), .Z(n3906) );
  IV U4453 ( .A(n3884), .Z(n3902) );
  XOR U4454 ( .A(n3909), .B(n3910), .Z(n3884) );
  ANDN U4455 ( .B(n3911), .A(n3912), .Z(n3909) );
  XOR U4456 ( .A(n3910), .B(n3913), .Z(n3911) );
  IV U4457 ( .A(n3892), .Z(n3896) );
  XOR U4458 ( .A(n3892), .B(n3874), .Z(n3894) );
  XOR U4459 ( .A(n3914), .B(n3915), .Z(n3874) );
  AND U4460 ( .A(n106), .B(n3916), .Z(n3914) );
  XOR U4461 ( .A(n3917), .B(n3915), .Z(n3916) );
  NANDN U4462 ( .A(n3876), .B(n3878), .Z(n3892) );
  XOR U4463 ( .A(n3918), .B(n3919), .Z(n3878) );
  AND U4464 ( .A(n106), .B(n3920), .Z(n3918) );
  XOR U4465 ( .A(n3919), .B(n3921), .Z(n3920) );
  XOR U4466 ( .A(n3922), .B(n3923), .Z(n106) );
  AND U4467 ( .A(n3924), .B(n3925), .Z(n3922) );
  XNOR U4468 ( .A(n3923), .B(n3889), .Z(n3925) );
  XNOR U4469 ( .A(n3926), .B(n3927), .Z(n3889) );
  ANDN U4470 ( .B(n3928), .A(n3929), .Z(n3926) );
  XOR U4471 ( .A(n3927), .B(n3930), .Z(n3928) );
  XOR U4472 ( .A(n3923), .B(n3891), .Z(n3924) );
  XOR U4473 ( .A(n3931), .B(n3932), .Z(n3891) );
  AND U4474 ( .A(n110), .B(n3933), .Z(n3931) );
  XOR U4475 ( .A(n3934), .B(n3932), .Z(n3933) );
  XNOR U4476 ( .A(n3935), .B(n3936), .Z(n3923) );
  NAND U4477 ( .A(n3937), .B(n3938), .Z(n3936) );
  XOR U4478 ( .A(n3939), .B(n3915), .Z(n3938) );
  XOR U4479 ( .A(n3929), .B(n3930), .Z(n3915) );
  XOR U4480 ( .A(n3940), .B(n3941), .Z(n3930) );
  ANDN U4481 ( .B(n3942), .A(n3943), .Z(n3940) );
  XOR U4482 ( .A(n3941), .B(n3944), .Z(n3942) );
  XOR U4483 ( .A(n3945), .B(n3946), .Z(n3929) );
  XOR U4484 ( .A(n3947), .B(n3948), .Z(n3946) );
  ANDN U4485 ( .B(n3949), .A(n3950), .Z(n3947) );
  XOR U4486 ( .A(n3951), .B(n3948), .Z(n3949) );
  IV U4487 ( .A(n3927), .Z(n3945) );
  XOR U4488 ( .A(n3952), .B(n3953), .Z(n3927) );
  ANDN U4489 ( .B(n3954), .A(n3955), .Z(n3952) );
  XOR U4490 ( .A(n3953), .B(n3956), .Z(n3954) );
  IV U4491 ( .A(n3935), .Z(n3939) );
  XOR U4492 ( .A(n3935), .B(n3917), .Z(n3937) );
  XOR U4493 ( .A(n3957), .B(n3958), .Z(n3917) );
  AND U4494 ( .A(n110), .B(n3959), .Z(n3957) );
  XOR U4495 ( .A(n3960), .B(n3958), .Z(n3959) );
  NANDN U4496 ( .A(n3919), .B(n3921), .Z(n3935) );
  XOR U4497 ( .A(n3961), .B(n3962), .Z(n3921) );
  AND U4498 ( .A(n110), .B(n3963), .Z(n3961) );
  XOR U4499 ( .A(n3962), .B(n3964), .Z(n3963) );
  XOR U4500 ( .A(n3965), .B(n3966), .Z(n110) );
  AND U4501 ( .A(n3967), .B(n3968), .Z(n3965) );
  XNOR U4502 ( .A(n3966), .B(n3932), .Z(n3968) );
  XNOR U4503 ( .A(n3969), .B(n3970), .Z(n3932) );
  ANDN U4504 ( .B(n3971), .A(n3972), .Z(n3969) );
  XOR U4505 ( .A(n3970), .B(n3973), .Z(n3971) );
  XOR U4506 ( .A(n3966), .B(n3934), .Z(n3967) );
  XOR U4507 ( .A(n3974), .B(n3975), .Z(n3934) );
  AND U4508 ( .A(n114), .B(n3976), .Z(n3974) );
  XOR U4509 ( .A(n3977), .B(n3975), .Z(n3976) );
  XNOR U4510 ( .A(n3978), .B(n3979), .Z(n3966) );
  NAND U4511 ( .A(n3980), .B(n3981), .Z(n3979) );
  XOR U4512 ( .A(n3982), .B(n3958), .Z(n3981) );
  XOR U4513 ( .A(n3972), .B(n3973), .Z(n3958) );
  XOR U4514 ( .A(n3983), .B(n3984), .Z(n3973) );
  ANDN U4515 ( .B(n3985), .A(n3986), .Z(n3983) );
  XOR U4516 ( .A(n3984), .B(n3987), .Z(n3985) );
  XOR U4517 ( .A(n3988), .B(n3989), .Z(n3972) );
  XOR U4518 ( .A(n3990), .B(n3991), .Z(n3989) );
  ANDN U4519 ( .B(n3992), .A(n3993), .Z(n3990) );
  XOR U4520 ( .A(n3994), .B(n3991), .Z(n3992) );
  IV U4521 ( .A(n3970), .Z(n3988) );
  XOR U4522 ( .A(n3995), .B(n3996), .Z(n3970) );
  ANDN U4523 ( .B(n3997), .A(n3998), .Z(n3995) );
  XOR U4524 ( .A(n3996), .B(n3999), .Z(n3997) );
  IV U4525 ( .A(n3978), .Z(n3982) );
  XOR U4526 ( .A(n3978), .B(n3960), .Z(n3980) );
  XOR U4527 ( .A(n4000), .B(n4001), .Z(n3960) );
  AND U4528 ( .A(n114), .B(n4002), .Z(n4000) );
  XOR U4529 ( .A(n4003), .B(n4001), .Z(n4002) );
  NANDN U4530 ( .A(n3962), .B(n3964), .Z(n3978) );
  XOR U4531 ( .A(n4004), .B(n4005), .Z(n3964) );
  AND U4532 ( .A(n114), .B(n4006), .Z(n4004) );
  XOR U4533 ( .A(n4005), .B(n4007), .Z(n4006) );
  XOR U4534 ( .A(n4008), .B(n4009), .Z(n114) );
  AND U4535 ( .A(n4010), .B(n4011), .Z(n4008) );
  XNOR U4536 ( .A(n4009), .B(n3975), .Z(n4011) );
  XNOR U4537 ( .A(n4012), .B(n4013), .Z(n3975) );
  ANDN U4538 ( .B(n4014), .A(n4015), .Z(n4012) );
  XOR U4539 ( .A(n4013), .B(n4016), .Z(n4014) );
  XOR U4540 ( .A(n4009), .B(n3977), .Z(n4010) );
  XOR U4541 ( .A(n4017), .B(n4018), .Z(n3977) );
  AND U4542 ( .A(n118), .B(n4019), .Z(n4017) );
  XOR U4543 ( .A(n4020), .B(n4018), .Z(n4019) );
  XNOR U4544 ( .A(n4021), .B(n4022), .Z(n4009) );
  NAND U4545 ( .A(n4023), .B(n4024), .Z(n4022) );
  XOR U4546 ( .A(n4025), .B(n4001), .Z(n4024) );
  XOR U4547 ( .A(n4015), .B(n4016), .Z(n4001) );
  XOR U4548 ( .A(n4026), .B(n4027), .Z(n4016) );
  ANDN U4549 ( .B(n4028), .A(n4029), .Z(n4026) );
  XOR U4550 ( .A(n4027), .B(n4030), .Z(n4028) );
  XOR U4551 ( .A(n4031), .B(n4032), .Z(n4015) );
  XOR U4552 ( .A(n4033), .B(n4034), .Z(n4032) );
  ANDN U4553 ( .B(n4035), .A(n4036), .Z(n4033) );
  XOR U4554 ( .A(n4037), .B(n4034), .Z(n4035) );
  IV U4555 ( .A(n4013), .Z(n4031) );
  XOR U4556 ( .A(n4038), .B(n4039), .Z(n4013) );
  ANDN U4557 ( .B(n4040), .A(n4041), .Z(n4038) );
  XOR U4558 ( .A(n4039), .B(n4042), .Z(n4040) );
  IV U4559 ( .A(n4021), .Z(n4025) );
  XOR U4560 ( .A(n4021), .B(n4003), .Z(n4023) );
  XOR U4561 ( .A(n4043), .B(n4044), .Z(n4003) );
  AND U4562 ( .A(n118), .B(n4045), .Z(n4043) );
  XOR U4563 ( .A(n4046), .B(n4044), .Z(n4045) );
  NANDN U4564 ( .A(n4005), .B(n4007), .Z(n4021) );
  XOR U4565 ( .A(n4047), .B(n4048), .Z(n4007) );
  AND U4566 ( .A(n118), .B(n4049), .Z(n4047) );
  XOR U4567 ( .A(n4048), .B(n4050), .Z(n4049) );
  XOR U4568 ( .A(n4051), .B(n4052), .Z(n118) );
  AND U4569 ( .A(n4053), .B(n4054), .Z(n4051) );
  XNOR U4570 ( .A(n4052), .B(n4018), .Z(n4054) );
  XNOR U4571 ( .A(n4055), .B(n4056), .Z(n4018) );
  ANDN U4572 ( .B(n4057), .A(n4058), .Z(n4055) );
  XOR U4573 ( .A(n4056), .B(n4059), .Z(n4057) );
  XOR U4574 ( .A(n4052), .B(n4020), .Z(n4053) );
  XOR U4575 ( .A(n4060), .B(n4061), .Z(n4020) );
  AND U4576 ( .A(n122), .B(n4062), .Z(n4060) );
  XOR U4577 ( .A(n4063), .B(n4061), .Z(n4062) );
  XNOR U4578 ( .A(n4064), .B(n4065), .Z(n4052) );
  NAND U4579 ( .A(n4066), .B(n4067), .Z(n4065) );
  XOR U4580 ( .A(n4068), .B(n4044), .Z(n4067) );
  XOR U4581 ( .A(n4058), .B(n4059), .Z(n4044) );
  XOR U4582 ( .A(n4069), .B(n4070), .Z(n4059) );
  ANDN U4583 ( .B(n4071), .A(n4072), .Z(n4069) );
  XOR U4584 ( .A(n4070), .B(n4073), .Z(n4071) );
  XOR U4585 ( .A(n4074), .B(n4075), .Z(n4058) );
  XOR U4586 ( .A(n4076), .B(n4077), .Z(n4075) );
  ANDN U4587 ( .B(n4078), .A(n4079), .Z(n4076) );
  XOR U4588 ( .A(n4080), .B(n4077), .Z(n4078) );
  IV U4589 ( .A(n4056), .Z(n4074) );
  XOR U4590 ( .A(n4081), .B(n4082), .Z(n4056) );
  ANDN U4591 ( .B(n4083), .A(n4084), .Z(n4081) );
  XOR U4592 ( .A(n4082), .B(n4085), .Z(n4083) );
  IV U4593 ( .A(n4064), .Z(n4068) );
  XOR U4594 ( .A(n4064), .B(n4046), .Z(n4066) );
  XOR U4595 ( .A(n4086), .B(n4087), .Z(n4046) );
  AND U4596 ( .A(n122), .B(n4088), .Z(n4086) );
  XOR U4597 ( .A(n4089), .B(n4087), .Z(n4088) );
  NANDN U4598 ( .A(n4048), .B(n4050), .Z(n4064) );
  XOR U4599 ( .A(n4090), .B(n4091), .Z(n4050) );
  AND U4600 ( .A(n122), .B(n4092), .Z(n4090) );
  XOR U4601 ( .A(n4091), .B(n4093), .Z(n4092) );
  XOR U4602 ( .A(n4094), .B(n4095), .Z(n122) );
  AND U4603 ( .A(n4096), .B(n4097), .Z(n4094) );
  XNOR U4604 ( .A(n4095), .B(n4061), .Z(n4097) );
  XNOR U4605 ( .A(n4098), .B(n4099), .Z(n4061) );
  ANDN U4606 ( .B(n4100), .A(n4101), .Z(n4098) );
  XOR U4607 ( .A(n4099), .B(n4102), .Z(n4100) );
  XOR U4608 ( .A(n4095), .B(n4063), .Z(n4096) );
  XOR U4609 ( .A(n4103), .B(n4104), .Z(n4063) );
  AND U4610 ( .A(n126), .B(n4105), .Z(n4103) );
  XOR U4611 ( .A(n4106), .B(n4104), .Z(n4105) );
  XNOR U4612 ( .A(n4107), .B(n4108), .Z(n4095) );
  NAND U4613 ( .A(n4109), .B(n4110), .Z(n4108) );
  XOR U4614 ( .A(n4111), .B(n4087), .Z(n4110) );
  XOR U4615 ( .A(n4101), .B(n4102), .Z(n4087) );
  XOR U4616 ( .A(n4112), .B(n4113), .Z(n4102) );
  ANDN U4617 ( .B(n4114), .A(n4115), .Z(n4112) );
  XOR U4618 ( .A(n4113), .B(n4116), .Z(n4114) );
  XOR U4619 ( .A(n4117), .B(n4118), .Z(n4101) );
  XOR U4620 ( .A(n4119), .B(n4120), .Z(n4118) );
  ANDN U4621 ( .B(n4121), .A(n4122), .Z(n4119) );
  XOR U4622 ( .A(n4123), .B(n4120), .Z(n4121) );
  IV U4623 ( .A(n4099), .Z(n4117) );
  XOR U4624 ( .A(n4124), .B(n4125), .Z(n4099) );
  ANDN U4625 ( .B(n4126), .A(n4127), .Z(n4124) );
  XOR U4626 ( .A(n4125), .B(n4128), .Z(n4126) );
  IV U4627 ( .A(n4107), .Z(n4111) );
  XOR U4628 ( .A(n4107), .B(n4089), .Z(n4109) );
  XOR U4629 ( .A(n4129), .B(n4130), .Z(n4089) );
  AND U4630 ( .A(n126), .B(n4131), .Z(n4129) );
  XOR U4631 ( .A(n4132), .B(n4130), .Z(n4131) );
  NANDN U4632 ( .A(n4091), .B(n4093), .Z(n4107) );
  XOR U4633 ( .A(n4133), .B(n4134), .Z(n4093) );
  AND U4634 ( .A(n126), .B(n4135), .Z(n4133) );
  XOR U4635 ( .A(n4134), .B(n4136), .Z(n4135) );
  XOR U4636 ( .A(n4137), .B(n4138), .Z(n126) );
  AND U4637 ( .A(n4139), .B(n4140), .Z(n4137) );
  XNOR U4638 ( .A(n4138), .B(n4104), .Z(n4140) );
  XNOR U4639 ( .A(n4141), .B(n4142), .Z(n4104) );
  ANDN U4640 ( .B(n4143), .A(n4144), .Z(n4141) );
  XOR U4641 ( .A(n4142), .B(n4145), .Z(n4143) );
  XOR U4642 ( .A(n4138), .B(n4106), .Z(n4139) );
  XOR U4643 ( .A(n4146), .B(n4147), .Z(n4106) );
  AND U4644 ( .A(n130), .B(n4148), .Z(n4146) );
  XOR U4645 ( .A(n4149), .B(n4147), .Z(n4148) );
  XNOR U4646 ( .A(n4150), .B(n4151), .Z(n4138) );
  NAND U4647 ( .A(n4152), .B(n4153), .Z(n4151) );
  XOR U4648 ( .A(n4154), .B(n4130), .Z(n4153) );
  XOR U4649 ( .A(n4144), .B(n4145), .Z(n4130) );
  XOR U4650 ( .A(n4155), .B(n4156), .Z(n4145) );
  ANDN U4651 ( .B(n4157), .A(n4158), .Z(n4155) );
  XOR U4652 ( .A(n4156), .B(n4159), .Z(n4157) );
  XOR U4653 ( .A(n4160), .B(n4161), .Z(n4144) );
  XOR U4654 ( .A(n4162), .B(n4163), .Z(n4161) );
  ANDN U4655 ( .B(n4164), .A(n4165), .Z(n4162) );
  XOR U4656 ( .A(n4166), .B(n4163), .Z(n4164) );
  IV U4657 ( .A(n4142), .Z(n4160) );
  XOR U4658 ( .A(n4167), .B(n4168), .Z(n4142) );
  ANDN U4659 ( .B(n4169), .A(n4170), .Z(n4167) );
  XOR U4660 ( .A(n4168), .B(n4171), .Z(n4169) );
  IV U4661 ( .A(n4150), .Z(n4154) );
  XOR U4662 ( .A(n4150), .B(n4132), .Z(n4152) );
  XOR U4663 ( .A(n4172), .B(n4173), .Z(n4132) );
  AND U4664 ( .A(n130), .B(n4174), .Z(n4172) );
  XOR U4665 ( .A(n4175), .B(n4173), .Z(n4174) );
  NANDN U4666 ( .A(n4134), .B(n4136), .Z(n4150) );
  XOR U4667 ( .A(n4176), .B(n4177), .Z(n4136) );
  AND U4668 ( .A(n130), .B(n4178), .Z(n4176) );
  XOR U4669 ( .A(n4177), .B(n4179), .Z(n4178) );
  XOR U4670 ( .A(n4180), .B(n4181), .Z(n130) );
  AND U4671 ( .A(n4182), .B(n4183), .Z(n4180) );
  XNOR U4672 ( .A(n4181), .B(n4147), .Z(n4183) );
  XNOR U4673 ( .A(n4184), .B(n4185), .Z(n4147) );
  ANDN U4674 ( .B(n4186), .A(n4187), .Z(n4184) );
  XOR U4675 ( .A(n4185), .B(n4188), .Z(n4186) );
  XOR U4676 ( .A(n4181), .B(n4149), .Z(n4182) );
  XOR U4677 ( .A(n4189), .B(n4190), .Z(n4149) );
  AND U4678 ( .A(n134), .B(n4191), .Z(n4189) );
  XOR U4679 ( .A(n4192), .B(n4190), .Z(n4191) );
  XNOR U4680 ( .A(n4193), .B(n4194), .Z(n4181) );
  NAND U4681 ( .A(n4195), .B(n4196), .Z(n4194) );
  XOR U4682 ( .A(n4197), .B(n4173), .Z(n4196) );
  XOR U4683 ( .A(n4187), .B(n4188), .Z(n4173) );
  XOR U4684 ( .A(n4198), .B(n4199), .Z(n4188) );
  ANDN U4685 ( .B(n4200), .A(n4201), .Z(n4198) );
  XOR U4686 ( .A(n4199), .B(n4202), .Z(n4200) );
  XOR U4687 ( .A(n4203), .B(n4204), .Z(n4187) );
  XOR U4688 ( .A(n4205), .B(n4206), .Z(n4204) );
  ANDN U4689 ( .B(n4207), .A(n4208), .Z(n4205) );
  XOR U4690 ( .A(n4209), .B(n4206), .Z(n4207) );
  IV U4691 ( .A(n4185), .Z(n4203) );
  XOR U4692 ( .A(n4210), .B(n4211), .Z(n4185) );
  ANDN U4693 ( .B(n4212), .A(n4213), .Z(n4210) );
  XOR U4694 ( .A(n4211), .B(n4214), .Z(n4212) );
  IV U4695 ( .A(n4193), .Z(n4197) );
  XOR U4696 ( .A(n4193), .B(n4175), .Z(n4195) );
  XOR U4697 ( .A(n4215), .B(n4216), .Z(n4175) );
  AND U4698 ( .A(n134), .B(n4217), .Z(n4215) );
  XOR U4699 ( .A(n4218), .B(n4216), .Z(n4217) );
  NANDN U4700 ( .A(n4177), .B(n4179), .Z(n4193) );
  XOR U4701 ( .A(n4219), .B(n4220), .Z(n4179) );
  AND U4702 ( .A(n134), .B(n4221), .Z(n4219) );
  XOR U4703 ( .A(n4220), .B(n4222), .Z(n4221) );
  XOR U4704 ( .A(n4223), .B(n4224), .Z(n134) );
  AND U4705 ( .A(n4225), .B(n4226), .Z(n4223) );
  XNOR U4706 ( .A(n4224), .B(n4190), .Z(n4226) );
  XNOR U4707 ( .A(n4227), .B(n4228), .Z(n4190) );
  ANDN U4708 ( .B(n4229), .A(n4230), .Z(n4227) );
  XOR U4709 ( .A(n4228), .B(n4231), .Z(n4229) );
  XOR U4710 ( .A(n4224), .B(n4192), .Z(n4225) );
  XOR U4711 ( .A(n4232), .B(n4233), .Z(n4192) );
  AND U4712 ( .A(n138), .B(n4234), .Z(n4232) );
  XOR U4713 ( .A(n4235), .B(n4233), .Z(n4234) );
  XNOR U4714 ( .A(n4236), .B(n4237), .Z(n4224) );
  NAND U4715 ( .A(n4238), .B(n4239), .Z(n4237) );
  XOR U4716 ( .A(n4240), .B(n4216), .Z(n4239) );
  XOR U4717 ( .A(n4230), .B(n4231), .Z(n4216) );
  XOR U4718 ( .A(n4241), .B(n4242), .Z(n4231) );
  ANDN U4719 ( .B(n4243), .A(n4244), .Z(n4241) );
  XOR U4720 ( .A(n4242), .B(n4245), .Z(n4243) );
  XOR U4721 ( .A(n4246), .B(n4247), .Z(n4230) );
  XOR U4722 ( .A(n4248), .B(n4249), .Z(n4247) );
  ANDN U4723 ( .B(n4250), .A(n4251), .Z(n4248) );
  XOR U4724 ( .A(n4252), .B(n4249), .Z(n4250) );
  IV U4725 ( .A(n4228), .Z(n4246) );
  XOR U4726 ( .A(n4253), .B(n4254), .Z(n4228) );
  ANDN U4727 ( .B(n4255), .A(n4256), .Z(n4253) );
  XOR U4728 ( .A(n4254), .B(n4257), .Z(n4255) );
  IV U4729 ( .A(n4236), .Z(n4240) );
  XOR U4730 ( .A(n4236), .B(n4218), .Z(n4238) );
  XOR U4731 ( .A(n4258), .B(n4259), .Z(n4218) );
  AND U4732 ( .A(n138), .B(n4260), .Z(n4258) );
  XOR U4733 ( .A(n4261), .B(n4259), .Z(n4260) );
  NANDN U4734 ( .A(n4220), .B(n4222), .Z(n4236) );
  XOR U4735 ( .A(n4262), .B(n4263), .Z(n4222) );
  AND U4736 ( .A(n138), .B(n4264), .Z(n4262) );
  XOR U4737 ( .A(n4263), .B(n4265), .Z(n4264) );
  XOR U4738 ( .A(n4266), .B(n4267), .Z(n138) );
  AND U4739 ( .A(n4268), .B(n4269), .Z(n4266) );
  XNOR U4740 ( .A(n4267), .B(n4233), .Z(n4269) );
  XNOR U4741 ( .A(n4270), .B(n4271), .Z(n4233) );
  ANDN U4742 ( .B(n4272), .A(n4273), .Z(n4270) );
  XOR U4743 ( .A(n4271), .B(n4274), .Z(n4272) );
  XOR U4744 ( .A(n4267), .B(n4235), .Z(n4268) );
  XOR U4745 ( .A(n4275), .B(n4276), .Z(n4235) );
  AND U4746 ( .A(n142), .B(n4277), .Z(n4275) );
  XOR U4747 ( .A(n4278), .B(n4276), .Z(n4277) );
  XNOR U4748 ( .A(n4279), .B(n4280), .Z(n4267) );
  NAND U4749 ( .A(n4281), .B(n4282), .Z(n4280) );
  XOR U4750 ( .A(n4283), .B(n4259), .Z(n4282) );
  XOR U4751 ( .A(n4273), .B(n4274), .Z(n4259) );
  XOR U4752 ( .A(n4284), .B(n4285), .Z(n4274) );
  ANDN U4753 ( .B(n4286), .A(n4287), .Z(n4284) );
  XOR U4754 ( .A(n4285), .B(n4288), .Z(n4286) );
  XOR U4755 ( .A(n4289), .B(n4290), .Z(n4273) );
  XOR U4756 ( .A(n4291), .B(n4292), .Z(n4290) );
  ANDN U4757 ( .B(n4293), .A(n4294), .Z(n4291) );
  XOR U4758 ( .A(n4295), .B(n4292), .Z(n4293) );
  IV U4759 ( .A(n4271), .Z(n4289) );
  XOR U4760 ( .A(n4296), .B(n4297), .Z(n4271) );
  ANDN U4761 ( .B(n4298), .A(n4299), .Z(n4296) );
  XOR U4762 ( .A(n4297), .B(n4300), .Z(n4298) );
  IV U4763 ( .A(n4279), .Z(n4283) );
  XOR U4764 ( .A(n4279), .B(n4261), .Z(n4281) );
  XOR U4765 ( .A(n4301), .B(n4302), .Z(n4261) );
  AND U4766 ( .A(n142), .B(n4303), .Z(n4301) );
  XOR U4767 ( .A(n4304), .B(n4302), .Z(n4303) );
  NANDN U4768 ( .A(n4263), .B(n4265), .Z(n4279) );
  XOR U4769 ( .A(n4305), .B(n4306), .Z(n4265) );
  AND U4770 ( .A(n142), .B(n4307), .Z(n4305) );
  XOR U4771 ( .A(n4306), .B(n4308), .Z(n4307) );
  XOR U4772 ( .A(n4309), .B(n4310), .Z(n142) );
  AND U4773 ( .A(n4311), .B(n4312), .Z(n4309) );
  XNOR U4774 ( .A(n4310), .B(n4276), .Z(n4312) );
  XNOR U4775 ( .A(n4313), .B(n4314), .Z(n4276) );
  ANDN U4776 ( .B(n4315), .A(n4316), .Z(n4313) );
  XOR U4777 ( .A(n4314), .B(n4317), .Z(n4315) );
  XOR U4778 ( .A(n4310), .B(n4278), .Z(n4311) );
  XOR U4779 ( .A(n4318), .B(n4319), .Z(n4278) );
  AND U4780 ( .A(n146), .B(n4320), .Z(n4318) );
  XOR U4781 ( .A(n4321), .B(n4319), .Z(n4320) );
  XNOR U4782 ( .A(n4322), .B(n4323), .Z(n4310) );
  NAND U4783 ( .A(n4324), .B(n4325), .Z(n4323) );
  XOR U4784 ( .A(n4326), .B(n4302), .Z(n4325) );
  XOR U4785 ( .A(n4316), .B(n4317), .Z(n4302) );
  XOR U4786 ( .A(n4327), .B(n4328), .Z(n4317) );
  ANDN U4787 ( .B(n4329), .A(n4330), .Z(n4327) );
  XOR U4788 ( .A(n4328), .B(n4331), .Z(n4329) );
  XOR U4789 ( .A(n4332), .B(n4333), .Z(n4316) );
  XOR U4790 ( .A(n4334), .B(n4335), .Z(n4333) );
  ANDN U4791 ( .B(n4336), .A(n4337), .Z(n4334) );
  XOR U4792 ( .A(n4338), .B(n4335), .Z(n4336) );
  IV U4793 ( .A(n4314), .Z(n4332) );
  XOR U4794 ( .A(n4339), .B(n4340), .Z(n4314) );
  ANDN U4795 ( .B(n4341), .A(n4342), .Z(n4339) );
  XOR U4796 ( .A(n4340), .B(n4343), .Z(n4341) );
  IV U4797 ( .A(n4322), .Z(n4326) );
  XOR U4798 ( .A(n4322), .B(n4304), .Z(n4324) );
  XOR U4799 ( .A(n4344), .B(n4345), .Z(n4304) );
  AND U4800 ( .A(n146), .B(n4346), .Z(n4344) );
  XOR U4801 ( .A(n4347), .B(n4345), .Z(n4346) );
  NANDN U4802 ( .A(n4306), .B(n4308), .Z(n4322) );
  XOR U4803 ( .A(n4348), .B(n4349), .Z(n4308) );
  AND U4804 ( .A(n146), .B(n4350), .Z(n4348) );
  XOR U4805 ( .A(n4349), .B(n4351), .Z(n4350) );
  XOR U4806 ( .A(n4352), .B(n4353), .Z(n146) );
  AND U4807 ( .A(n4354), .B(n4355), .Z(n4352) );
  XNOR U4808 ( .A(n4353), .B(n4319), .Z(n4355) );
  XNOR U4809 ( .A(n4356), .B(n4357), .Z(n4319) );
  ANDN U4810 ( .B(n4358), .A(n4359), .Z(n4356) );
  XOR U4811 ( .A(n4357), .B(n4360), .Z(n4358) );
  XOR U4812 ( .A(n4353), .B(n4321), .Z(n4354) );
  XOR U4813 ( .A(n4361), .B(n4362), .Z(n4321) );
  AND U4814 ( .A(n150), .B(n4363), .Z(n4361) );
  XOR U4815 ( .A(n4364), .B(n4362), .Z(n4363) );
  XNOR U4816 ( .A(n4365), .B(n4366), .Z(n4353) );
  NAND U4817 ( .A(n4367), .B(n4368), .Z(n4366) );
  XOR U4818 ( .A(n4369), .B(n4345), .Z(n4368) );
  XOR U4819 ( .A(n4359), .B(n4360), .Z(n4345) );
  XOR U4820 ( .A(n4370), .B(n4371), .Z(n4360) );
  ANDN U4821 ( .B(n4372), .A(n4373), .Z(n4370) );
  XOR U4822 ( .A(n4371), .B(n4374), .Z(n4372) );
  XOR U4823 ( .A(n4375), .B(n4376), .Z(n4359) );
  XOR U4824 ( .A(n4377), .B(n4378), .Z(n4376) );
  ANDN U4825 ( .B(n4379), .A(n4380), .Z(n4377) );
  XOR U4826 ( .A(n4381), .B(n4378), .Z(n4379) );
  IV U4827 ( .A(n4357), .Z(n4375) );
  XOR U4828 ( .A(n4382), .B(n4383), .Z(n4357) );
  ANDN U4829 ( .B(n4384), .A(n4385), .Z(n4382) );
  XOR U4830 ( .A(n4383), .B(n4386), .Z(n4384) );
  IV U4831 ( .A(n4365), .Z(n4369) );
  XOR U4832 ( .A(n4365), .B(n4347), .Z(n4367) );
  XOR U4833 ( .A(n4387), .B(n4388), .Z(n4347) );
  AND U4834 ( .A(n150), .B(n4389), .Z(n4387) );
  XOR U4835 ( .A(n4390), .B(n4388), .Z(n4389) );
  NANDN U4836 ( .A(n4349), .B(n4351), .Z(n4365) );
  XOR U4837 ( .A(n4391), .B(n4392), .Z(n4351) );
  AND U4838 ( .A(n150), .B(n4393), .Z(n4391) );
  XOR U4839 ( .A(n4392), .B(n4394), .Z(n4393) );
  XOR U4840 ( .A(n4395), .B(n4396), .Z(n150) );
  AND U4841 ( .A(n4397), .B(n4398), .Z(n4395) );
  XNOR U4842 ( .A(n4396), .B(n4362), .Z(n4398) );
  XNOR U4843 ( .A(n4399), .B(n4400), .Z(n4362) );
  ANDN U4844 ( .B(n4401), .A(n4402), .Z(n4399) );
  XOR U4845 ( .A(n4400), .B(n4403), .Z(n4401) );
  XOR U4846 ( .A(n4396), .B(n4364), .Z(n4397) );
  XOR U4847 ( .A(n4404), .B(n4405), .Z(n4364) );
  AND U4848 ( .A(n154), .B(n4406), .Z(n4404) );
  XOR U4849 ( .A(n4407), .B(n4405), .Z(n4406) );
  XNOR U4850 ( .A(n4408), .B(n4409), .Z(n4396) );
  NAND U4851 ( .A(n4410), .B(n4411), .Z(n4409) );
  XOR U4852 ( .A(n4412), .B(n4388), .Z(n4411) );
  XOR U4853 ( .A(n4402), .B(n4403), .Z(n4388) );
  XOR U4854 ( .A(n4413), .B(n4414), .Z(n4403) );
  ANDN U4855 ( .B(n4415), .A(n4416), .Z(n4413) );
  XOR U4856 ( .A(n4414), .B(n4417), .Z(n4415) );
  XOR U4857 ( .A(n4418), .B(n4419), .Z(n4402) );
  XOR U4858 ( .A(n4420), .B(n4421), .Z(n4419) );
  ANDN U4859 ( .B(n4422), .A(n4423), .Z(n4420) );
  XOR U4860 ( .A(n4424), .B(n4421), .Z(n4422) );
  IV U4861 ( .A(n4400), .Z(n4418) );
  XOR U4862 ( .A(n4425), .B(n4426), .Z(n4400) );
  ANDN U4863 ( .B(n4427), .A(n4428), .Z(n4425) );
  XOR U4864 ( .A(n4426), .B(n4429), .Z(n4427) );
  IV U4865 ( .A(n4408), .Z(n4412) );
  XOR U4866 ( .A(n4408), .B(n4390), .Z(n4410) );
  XOR U4867 ( .A(n4430), .B(n4431), .Z(n4390) );
  AND U4868 ( .A(n154), .B(n4432), .Z(n4430) );
  XOR U4869 ( .A(n4433), .B(n4431), .Z(n4432) );
  NANDN U4870 ( .A(n4392), .B(n4394), .Z(n4408) );
  XOR U4871 ( .A(n4434), .B(n4435), .Z(n4394) );
  AND U4872 ( .A(n154), .B(n4436), .Z(n4434) );
  XOR U4873 ( .A(n4435), .B(n4437), .Z(n4436) );
  XOR U4874 ( .A(n4438), .B(n4439), .Z(n154) );
  AND U4875 ( .A(n4440), .B(n4441), .Z(n4438) );
  XNOR U4876 ( .A(n4439), .B(n4405), .Z(n4441) );
  XNOR U4877 ( .A(n4442), .B(n4443), .Z(n4405) );
  ANDN U4878 ( .B(n4444), .A(n4445), .Z(n4442) );
  XOR U4879 ( .A(n4443), .B(n4446), .Z(n4444) );
  XOR U4880 ( .A(n4439), .B(n4407), .Z(n4440) );
  XOR U4881 ( .A(n4447), .B(n4448), .Z(n4407) );
  AND U4882 ( .A(n158), .B(n4449), .Z(n4447) );
  XOR U4883 ( .A(n4450), .B(n4448), .Z(n4449) );
  XNOR U4884 ( .A(n4451), .B(n4452), .Z(n4439) );
  NAND U4885 ( .A(n4453), .B(n4454), .Z(n4452) );
  XOR U4886 ( .A(n4455), .B(n4431), .Z(n4454) );
  XOR U4887 ( .A(n4445), .B(n4446), .Z(n4431) );
  XOR U4888 ( .A(n4456), .B(n4457), .Z(n4446) );
  ANDN U4889 ( .B(n4458), .A(n4459), .Z(n4456) );
  XOR U4890 ( .A(n4457), .B(n4460), .Z(n4458) );
  XOR U4891 ( .A(n4461), .B(n4462), .Z(n4445) );
  XOR U4892 ( .A(n4463), .B(n4464), .Z(n4462) );
  ANDN U4893 ( .B(n4465), .A(n4466), .Z(n4463) );
  XOR U4894 ( .A(n4467), .B(n4464), .Z(n4465) );
  IV U4895 ( .A(n4443), .Z(n4461) );
  XOR U4896 ( .A(n4468), .B(n4469), .Z(n4443) );
  ANDN U4897 ( .B(n4470), .A(n4471), .Z(n4468) );
  XOR U4898 ( .A(n4469), .B(n4472), .Z(n4470) );
  IV U4899 ( .A(n4451), .Z(n4455) );
  XOR U4900 ( .A(n4451), .B(n4433), .Z(n4453) );
  XOR U4901 ( .A(n4473), .B(n4474), .Z(n4433) );
  AND U4902 ( .A(n158), .B(n4475), .Z(n4473) );
  XOR U4903 ( .A(n4476), .B(n4474), .Z(n4475) );
  NANDN U4904 ( .A(n4435), .B(n4437), .Z(n4451) );
  XOR U4905 ( .A(n4477), .B(n4478), .Z(n4437) );
  AND U4906 ( .A(n158), .B(n4479), .Z(n4477) );
  XOR U4907 ( .A(n4478), .B(n4480), .Z(n4479) );
  XOR U4908 ( .A(n4481), .B(n4482), .Z(n158) );
  AND U4909 ( .A(n4483), .B(n4484), .Z(n4481) );
  XNOR U4910 ( .A(n4482), .B(n4448), .Z(n4484) );
  XNOR U4911 ( .A(n4485), .B(n4486), .Z(n4448) );
  ANDN U4912 ( .B(n4487), .A(n4488), .Z(n4485) );
  XOR U4913 ( .A(n4486), .B(n4489), .Z(n4487) );
  XOR U4914 ( .A(n4482), .B(n4450), .Z(n4483) );
  XOR U4915 ( .A(n4490), .B(n4491), .Z(n4450) );
  AND U4916 ( .A(n162), .B(n4492), .Z(n4490) );
  XOR U4917 ( .A(n4493), .B(n4491), .Z(n4492) );
  XNOR U4918 ( .A(n4494), .B(n4495), .Z(n4482) );
  NAND U4919 ( .A(n4496), .B(n4497), .Z(n4495) );
  XOR U4920 ( .A(n4498), .B(n4474), .Z(n4497) );
  XOR U4921 ( .A(n4488), .B(n4489), .Z(n4474) );
  XOR U4922 ( .A(n4499), .B(n4500), .Z(n4489) );
  ANDN U4923 ( .B(n4501), .A(n4502), .Z(n4499) );
  XOR U4924 ( .A(n4500), .B(n4503), .Z(n4501) );
  XOR U4925 ( .A(n4504), .B(n4505), .Z(n4488) );
  XOR U4926 ( .A(n4506), .B(n4507), .Z(n4505) );
  ANDN U4927 ( .B(n4508), .A(n4509), .Z(n4506) );
  XOR U4928 ( .A(n4510), .B(n4507), .Z(n4508) );
  IV U4929 ( .A(n4486), .Z(n4504) );
  XOR U4930 ( .A(n4511), .B(n4512), .Z(n4486) );
  ANDN U4931 ( .B(n4513), .A(n4514), .Z(n4511) );
  XOR U4932 ( .A(n4512), .B(n4515), .Z(n4513) );
  IV U4933 ( .A(n4494), .Z(n4498) );
  XOR U4934 ( .A(n4494), .B(n4476), .Z(n4496) );
  XOR U4935 ( .A(n4516), .B(n4517), .Z(n4476) );
  AND U4936 ( .A(n162), .B(n4518), .Z(n4516) );
  XOR U4937 ( .A(n4519), .B(n4517), .Z(n4518) );
  NANDN U4938 ( .A(n4478), .B(n4480), .Z(n4494) );
  XOR U4939 ( .A(n4520), .B(n4521), .Z(n4480) );
  AND U4940 ( .A(n162), .B(n4522), .Z(n4520) );
  XOR U4941 ( .A(n4521), .B(n4523), .Z(n4522) );
  XOR U4942 ( .A(n4524), .B(n4525), .Z(n162) );
  AND U4943 ( .A(n4526), .B(n4527), .Z(n4524) );
  XNOR U4944 ( .A(n4525), .B(n4491), .Z(n4527) );
  XNOR U4945 ( .A(n4528), .B(n4529), .Z(n4491) );
  ANDN U4946 ( .B(n4530), .A(n4531), .Z(n4528) );
  XOR U4947 ( .A(n4529), .B(n4532), .Z(n4530) );
  XOR U4948 ( .A(n4525), .B(n4493), .Z(n4526) );
  XOR U4949 ( .A(n4533), .B(n4534), .Z(n4493) );
  AND U4950 ( .A(n166), .B(n4535), .Z(n4533) );
  XOR U4951 ( .A(n4536), .B(n4534), .Z(n4535) );
  XNOR U4952 ( .A(n4537), .B(n4538), .Z(n4525) );
  NAND U4953 ( .A(n4539), .B(n4540), .Z(n4538) );
  XOR U4954 ( .A(n4541), .B(n4517), .Z(n4540) );
  XOR U4955 ( .A(n4531), .B(n4532), .Z(n4517) );
  XOR U4956 ( .A(n4542), .B(n4543), .Z(n4532) );
  ANDN U4957 ( .B(n4544), .A(n4545), .Z(n4542) );
  XOR U4958 ( .A(n4543), .B(n4546), .Z(n4544) );
  XOR U4959 ( .A(n4547), .B(n4548), .Z(n4531) );
  XOR U4960 ( .A(n4549), .B(n4550), .Z(n4548) );
  ANDN U4961 ( .B(n4551), .A(n4552), .Z(n4549) );
  XOR U4962 ( .A(n4553), .B(n4550), .Z(n4551) );
  IV U4963 ( .A(n4529), .Z(n4547) );
  XOR U4964 ( .A(n4554), .B(n4555), .Z(n4529) );
  ANDN U4965 ( .B(n4556), .A(n4557), .Z(n4554) );
  XOR U4966 ( .A(n4555), .B(n4558), .Z(n4556) );
  IV U4967 ( .A(n4537), .Z(n4541) );
  XOR U4968 ( .A(n4537), .B(n4519), .Z(n4539) );
  XOR U4969 ( .A(n4559), .B(n4560), .Z(n4519) );
  AND U4970 ( .A(n166), .B(n4561), .Z(n4559) );
  XOR U4971 ( .A(n4562), .B(n4560), .Z(n4561) );
  NANDN U4972 ( .A(n4521), .B(n4523), .Z(n4537) );
  XOR U4973 ( .A(n4563), .B(n4564), .Z(n4523) );
  AND U4974 ( .A(n166), .B(n4565), .Z(n4563) );
  XOR U4975 ( .A(n4564), .B(n4566), .Z(n4565) );
  XOR U4976 ( .A(n4567), .B(n4568), .Z(n166) );
  AND U4977 ( .A(n4569), .B(n4570), .Z(n4567) );
  XNOR U4978 ( .A(n4568), .B(n4534), .Z(n4570) );
  XNOR U4979 ( .A(n4571), .B(n4572), .Z(n4534) );
  ANDN U4980 ( .B(n4573), .A(n4574), .Z(n4571) );
  XOR U4981 ( .A(n4572), .B(n4575), .Z(n4573) );
  XOR U4982 ( .A(n4568), .B(n4536), .Z(n4569) );
  XOR U4983 ( .A(n4576), .B(n4577), .Z(n4536) );
  AND U4984 ( .A(n170), .B(n4578), .Z(n4576) );
  XOR U4985 ( .A(n4579), .B(n4577), .Z(n4578) );
  XNOR U4986 ( .A(n4580), .B(n4581), .Z(n4568) );
  NAND U4987 ( .A(n4582), .B(n4583), .Z(n4581) );
  XOR U4988 ( .A(n4584), .B(n4560), .Z(n4583) );
  XOR U4989 ( .A(n4574), .B(n4575), .Z(n4560) );
  XOR U4990 ( .A(n4585), .B(n4586), .Z(n4575) );
  ANDN U4991 ( .B(n4587), .A(n4588), .Z(n4585) );
  XOR U4992 ( .A(n4586), .B(n4589), .Z(n4587) );
  XOR U4993 ( .A(n4590), .B(n4591), .Z(n4574) );
  XOR U4994 ( .A(n4592), .B(n4593), .Z(n4591) );
  ANDN U4995 ( .B(n4594), .A(n4595), .Z(n4592) );
  XOR U4996 ( .A(n4596), .B(n4593), .Z(n4594) );
  IV U4997 ( .A(n4572), .Z(n4590) );
  XOR U4998 ( .A(n4597), .B(n4598), .Z(n4572) );
  ANDN U4999 ( .B(n4599), .A(n4600), .Z(n4597) );
  XOR U5000 ( .A(n4598), .B(n4601), .Z(n4599) );
  IV U5001 ( .A(n4580), .Z(n4584) );
  XOR U5002 ( .A(n4580), .B(n4562), .Z(n4582) );
  XOR U5003 ( .A(n4602), .B(n4603), .Z(n4562) );
  AND U5004 ( .A(n170), .B(n4604), .Z(n4602) );
  XOR U5005 ( .A(n4605), .B(n4603), .Z(n4604) );
  NANDN U5006 ( .A(n4564), .B(n4566), .Z(n4580) );
  XOR U5007 ( .A(n4606), .B(n4607), .Z(n4566) );
  AND U5008 ( .A(n170), .B(n4608), .Z(n4606) );
  XOR U5009 ( .A(n4607), .B(n4609), .Z(n4608) );
  XOR U5010 ( .A(n4610), .B(n4611), .Z(n170) );
  AND U5011 ( .A(n4612), .B(n4613), .Z(n4610) );
  XNOR U5012 ( .A(n4611), .B(n4577), .Z(n4613) );
  XNOR U5013 ( .A(n4614), .B(n4615), .Z(n4577) );
  ANDN U5014 ( .B(n4616), .A(n4617), .Z(n4614) );
  XOR U5015 ( .A(n4615), .B(n4618), .Z(n4616) );
  XOR U5016 ( .A(n4611), .B(n4579), .Z(n4612) );
  XOR U5017 ( .A(n4619), .B(n4620), .Z(n4579) );
  AND U5018 ( .A(n174), .B(n4621), .Z(n4619) );
  XOR U5019 ( .A(n4622), .B(n4620), .Z(n4621) );
  XNOR U5020 ( .A(n4623), .B(n4624), .Z(n4611) );
  NAND U5021 ( .A(n4625), .B(n4626), .Z(n4624) );
  XOR U5022 ( .A(n4627), .B(n4603), .Z(n4626) );
  XOR U5023 ( .A(n4617), .B(n4618), .Z(n4603) );
  XOR U5024 ( .A(n4628), .B(n4629), .Z(n4618) );
  ANDN U5025 ( .B(n4630), .A(n4631), .Z(n4628) );
  XOR U5026 ( .A(n4629), .B(n4632), .Z(n4630) );
  XOR U5027 ( .A(n4633), .B(n4634), .Z(n4617) );
  XOR U5028 ( .A(n4635), .B(n4636), .Z(n4634) );
  ANDN U5029 ( .B(n4637), .A(n4638), .Z(n4635) );
  XOR U5030 ( .A(n4639), .B(n4636), .Z(n4637) );
  IV U5031 ( .A(n4615), .Z(n4633) );
  XOR U5032 ( .A(n4640), .B(n4641), .Z(n4615) );
  ANDN U5033 ( .B(n4642), .A(n4643), .Z(n4640) );
  XOR U5034 ( .A(n4641), .B(n4644), .Z(n4642) );
  IV U5035 ( .A(n4623), .Z(n4627) );
  XOR U5036 ( .A(n4623), .B(n4605), .Z(n4625) );
  XOR U5037 ( .A(n4645), .B(n4646), .Z(n4605) );
  AND U5038 ( .A(n174), .B(n4647), .Z(n4645) );
  XOR U5039 ( .A(n4648), .B(n4646), .Z(n4647) );
  NANDN U5040 ( .A(n4607), .B(n4609), .Z(n4623) );
  XOR U5041 ( .A(n4649), .B(n4650), .Z(n4609) );
  AND U5042 ( .A(n174), .B(n4651), .Z(n4649) );
  XOR U5043 ( .A(n4650), .B(n4652), .Z(n4651) );
  XOR U5044 ( .A(n4653), .B(n4654), .Z(n174) );
  AND U5045 ( .A(n4655), .B(n4656), .Z(n4653) );
  XNOR U5046 ( .A(n4654), .B(n4620), .Z(n4656) );
  XNOR U5047 ( .A(n4657), .B(n4658), .Z(n4620) );
  ANDN U5048 ( .B(n4659), .A(n4660), .Z(n4657) );
  XOR U5049 ( .A(n4658), .B(n4661), .Z(n4659) );
  XOR U5050 ( .A(n4654), .B(n4622), .Z(n4655) );
  XOR U5051 ( .A(n4662), .B(n4663), .Z(n4622) );
  AND U5052 ( .A(n178), .B(n4664), .Z(n4662) );
  XOR U5053 ( .A(n4665), .B(n4663), .Z(n4664) );
  XNOR U5054 ( .A(n4666), .B(n4667), .Z(n4654) );
  NAND U5055 ( .A(n4668), .B(n4669), .Z(n4667) );
  XOR U5056 ( .A(n4670), .B(n4646), .Z(n4669) );
  XOR U5057 ( .A(n4660), .B(n4661), .Z(n4646) );
  XOR U5058 ( .A(n4671), .B(n4672), .Z(n4661) );
  ANDN U5059 ( .B(n4673), .A(n4674), .Z(n4671) );
  XOR U5060 ( .A(n4672), .B(n4675), .Z(n4673) );
  XOR U5061 ( .A(n4676), .B(n4677), .Z(n4660) );
  XOR U5062 ( .A(n4678), .B(n4679), .Z(n4677) );
  ANDN U5063 ( .B(n4680), .A(n4681), .Z(n4678) );
  XOR U5064 ( .A(n4682), .B(n4679), .Z(n4680) );
  IV U5065 ( .A(n4658), .Z(n4676) );
  XOR U5066 ( .A(n4683), .B(n4684), .Z(n4658) );
  ANDN U5067 ( .B(n4685), .A(n4686), .Z(n4683) );
  XOR U5068 ( .A(n4684), .B(n4687), .Z(n4685) );
  IV U5069 ( .A(n4666), .Z(n4670) );
  XOR U5070 ( .A(n4666), .B(n4648), .Z(n4668) );
  XOR U5071 ( .A(n4688), .B(n4689), .Z(n4648) );
  AND U5072 ( .A(n178), .B(n4690), .Z(n4688) );
  XOR U5073 ( .A(n4691), .B(n4689), .Z(n4690) );
  NANDN U5074 ( .A(n4650), .B(n4652), .Z(n4666) );
  XOR U5075 ( .A(n4692), .B(n4693), .Z(n4652) );
  AND U5076 ( .A(n178), .B(n4694), .Z(n4692) );
  XOR U5077 ( .A(n4693), .B(n4695), .Z(n4694) );
  XOR U5078 ( .A(n4696), .B(n4697), .Z(n178) );
  AND U5079 ( .A(n4698), .B(n4699), .Z(n4696) );
  XNOR U5080 ( .A(n4697), .B(n4663), .Z(n4699) );
  XNOR U5081 ( .A(n4700), .B(n4701), .Z(n4663) );
  ANDN U5082 ( .B(n4702), .A(n4703), .Z(n4700) );
  XOR U5083 ( .A(n4701), .B(n4704), .Z(n4702) );
  XOR U5084 ( .A(n4697), .B(n4665), .Z(n4698) );
  XOR U5085 ( .A(n4705), .B(n4706), .Z(n4665) );
  AND U5086 ( .A(n182), .B(n4707), .Z(n4705) );
  XOR U5087 ( .A(n4708), .B(n4706), .Z(n4707) );
  XNOR U5088 ( .A(n4709), .B(n4710), .Z(n4697) );
  NAND U5089 ( .A(n4711), .B(n4712), .Z(n4710) );
  XOR U5090 ( .A(n4713), .B(n4689), .Z(n4712) );
  XOR U5091 ( .A(n4703), .B(n4704), .Z(n4689) );
  XOR U5092 ( .A(n4714), .B(n4715), .Z(n4704) );
  ANDN U5093 ( .B(n4716), .A(n4717), .Z(n4714) );
  XOR U5094 ( .A(n4715), .B(n4718), .Z(n4716) );
  XOR U5095 ( .A(n4719), .B(n4720), .Z(n4703) );
  XOR U5096 ( .A(n4721), .B(n4722), .Z(n4720) );
  ANDN U5097 ( .B(n4723), .A(n4724), .Z(n4721) );
  XOR U5098 ( .A(n4725), .B(n4722), .Z(n4723) );
  IV U5099 ( .A(n4701), .Z(n4719) );
  XOR U5100 ( .A(n4726), .B(n4727), .Z(n4701) );
  ANDN U5101 ( .B(n4728), .A(n4729), .Z(n4726) );
  XOR U5102 ( .A(n4727), .B(n4730), .Z(n4728) );
  IV U5103 ( .A(n4709), .Z(n4713) );
  XOR U5104 ( .A(n4709), .B(n4691), .Z(n4711) );
  XOR U5105 ( .A(n4731), .B(n4732), .Z(n4691) );
  AND U5106 ( .A(n182), .B(n4733), .Z(n4731) );
  XOR U5107 ( .A(n4734), .B(n4732), .Z(n4733) );
  NANDN U5108 ( .A(n4693), .B(n4695), .Z(n4709) );
  XOR U5109 ( .A(n4735), .B(n4736), .Z(n4695) );
  AND U5110 ( .A(n182), .B(n4737), .Z(n4735) );
  XOR U5111 ( .A(n4736), .B(n4738), .Z(n4737) );
  XOR U5112 ( .A(n4739), .B(n4740), .Z(n182) );
  AND U5113 ( .A(n4741), .B(n4742), .Z(n4739) );
  XNOR U5114 ( .A(n4740), .B(n4706), .Z(n4742) );
  XNOR U5115 ( .A(n4743), .B(n4744), .Z(n4706) );
  ANDN U5116 ( .B(n4745), .A(n4746), .Z(n4743) );
  XOR U5117 ( .A(n4744), .B(n4747), .Z(n4745) );
  XOR U5118 ( .A(n4740), .B(n4708), .Z(n4741) );
  XOR U5119 ( .A(n4748), .B(n4749), .Z(n4708) );
  AND U5120 ( .A(n186), .B(n4750), .Z(n4748) );
  XOR U5121 ( .A(n4751), .B(n4749), .Z(n4750) );
  XNOR U5122 ( .A(n4752), .B(n4753), .Z(n4740) );
  NAND U5123 ( .A(n4754), .B(n4755), .Z(n4753) );
  XOR U5124 ( .A(n4756), .B(n4732), .Z(n4755) );
  XOR U5125 ( .A(n4746), .B(n4747), .Z(n4732) );
  XOR U5126 ( .A(n4757), .B(n4758), .Z(n4747) );
  ANDN U5127 ( .B(n4759), .A(n4760), .Z(n4757) );
  XOR U5128 ( .A(n4758), .B(n4761), .Z(n4759) );
  XOR U5129 ( .A(n4762), .B(n4763), .Z(n4746) );
  XOR U5130 ( .A(n4764), .B(n4765), .Z(n4763) );
  ANDN U5131 ( .B(n4766), .A(n4767), .Z(n4764) );
  XOR U5132 ( .A(n4768), .B(n4765), .Z(n4766) );
  IV U5133 ( .A(n4744), .Z(n4762) );
  XOR U5134 ( .A(n4769), .B(n4770), .Z(n4744) );
  ANDN U5135 ( .B(n4771), .A(n4772), .Z(n4769) );
  XOR U5136 ( .A(n4770), .B(n4773), .Z(n4771) );
  IV U5137 ( .A(n4752), .Z(n4756) );
  XOR U5138 ( .A(n4752), .B(n4734), .Z(n4754) );
  XOR U5139 ( .A(n4774), .B(n4775), .Z(n4734) );
  AND U5140 ( .A(n186), .B(n4776), .Z(n4774) );
  XOR U5141 ( .A(n4777), .B(n4775), .Z(n4776) );
  NANDN U5142 ( .A(n4736), .B(n4738), .Z(n4752) );
  XOR U5143 ( .A(n4778), .B(n4779), .Z(n4738) );
  AND U5144 ( .A(n186), .B(n4780), .Z(n4778) );
  XOR U5145 ( .A(n4779), .B(n4781), .Z(n4780) );
  XOR U5146 ( .A(n4782), .B(n4783), .Z(n186) );
  AND U5147 ( .A(n4784), .B(n4785), .Z(n4782) );
  XNOR U5148 ( .A(n4783), .B(n4749), .Z(n4785) );
  XNOR U5149 ( .A(n4786), .B(n4787), .Z(n4749) );
  ANDN U5150 ( .B(n4788), .A(n4789), .Z(n4786) );
  XOR U5151 ( .A(n4787), .B(n4790), .Z(n4788) );
  XOR U5152 ( .A(n4783), .B(n4751), .Z(n4784) );
  XOR U5153 ( .A(n4791), .B(n4792), .Z(n4751) );
  AND U5154 ( .A(n190), .B(n4793), .Z(n4791) );
  XOR U5155 ( .A(n4794), .B(n4792), .Z(n4793) );
  XNOR U5156 ( .A(n4795), .B(n4796), .Z(n4783) );
  NAND U5157 ( .A(n4797), .B(n4798), .Z(n4796) );
  XOR U5158 ( .A(n4799), .B(n4775), .Z(n4798) );
  XOR U5159 ( .A(n4789), .B(n4790), .Z(n4775) );
  XOR U5160 ( .A(n4800), .B(n4801), .Z(n4790) );
  ANDN U5161 ( .B(n4802), .A(n4803), .Z(n4800) );
  XOR U5162 ( .A(n4801), .B(n4804), .Z(n4802) );
  XOR U5163 ( .A(n4805), .B(n4806), .Z(n4789) );
  XOR U5164 ( .A(n4807), .B(n4808), .Z(n4806) );
  ANDN U5165 ( .B(n4809), .A(n4810), .Z(n4807) );
  XOR U5166 ( .A(n4811), .B(n4808), .Z(n4809) );
  IV U5167 ( .A(n4787), .Z(n4805) );
  XOR U5168 ( .A(n4812), .B(n4813), .Z(n4787) );
  ANDN U5169 ( .B(n4814), .A(n4815), .Z(n4812) );
  XOR U5170 ( .A(n4813), .B(n4816), .Z(n4814) );
  IV U5171 ( .A(n4795), .Z(n4799) );
  XOR U5172 ( .A(n4795), .B(n4777), .Z(n4797) );
  XOR U5173 ( .A(n4817), .B(n4818), .Z(n4777) );
  AND U5174 ( .A(n190), .B(n4819), .Z(n4817) );
  XOR U5175 ( .A(n4820), .B(n4818), .Z(n4819) );
  NANDN U5176 ( .A(n4779), .B(n4781), .Z(n4795) );
  XOR U5177 ( .A(n4821), .B(n4822), .Z(n4781) );
  AND U5178 ( .A(n190), .B(n4823), .Z(n4821) );
  XOR U5179 ( .A(n4822), .B(n4824), .Z(n4823) );
  XOR U5180 ( .A(n4825), .B(n4826), .Z(n190) );
  AND U5181 ( .A(n4827), .B(n4828), .Z(n4825) );
  XNOR U5182 ( .A(n4826), .B(n4792), .Z(n4828) );
  XNOR U5183 ( .A(n4829), .B(n4830), .Z(n4792) );
  ANDN U5184 ( .B(n4831), .A(n4832), .Z(n4829) );
  XOR U5185 ( .A(n4830), .B(n4833), .Z(n4831) );
  XOR U5186 ( .A(n4826), .B(n4794), .Z(n4827) );
  XOR U5187 ( .A(n4834), .B(n4835), .Z(n4794) );
  AND U5188 ( .A(n194), .B(n4836), .Z(n4834) );
  XOR U5189 ( .A(n4837), .B(n4835), .Z(n4836) );
  XNOR U5190 ( .A(n4838), .B(n4839), .Z(n4826) );
  NAND U5191 ( .A(n4840), .B(n4841), .Z(n4839) );
  XOR U5192 ( .A(n4842), .B(n4818), .Z(n4841) );
  XOR U5193 ( .A(n4832), .B(n4833), .Z(n4818) );
  XOR U5194 ( .A(n4843), .B(n4844), .Z(n4833) );
  ANDN U5195 ( .B(n4845), .A(n4846), .Z(n4843) );
  XOR U5196 ( .A(n4844), .B(n4847), .Z(n4845) );
  XOR U5197 ( .A(n4848), .B(n4849), .Z(n4832) );
  XOR U5198 ( .A(n4850), .B(n4851), .Z(n4849) );
  ANDN U5199 ( .B(n4852), .A(n4853), .Z(n4850) );
  XOR U5200 ( .A(n4854), .B(n4851), .Z(n4852) );
  IV U5201 ( .A(n4830), .Z(n4848) );
  XOR U5202 ( .A(n4855), .B(n4856), .Z(n4830) );
  ANDN U5203 ( .B(n4857), .A(n4858), .Z(n4855) );
  XOR U5204 ( .A(n4856), .B(n4859), .Z(n4857) );
  IV U5205 ( .A(n4838), .Z(n4842) );
  XOR U5206 ( .A(n4838), .B(n4820), .Z(n4840) );
  XOR U5207 ( .A(n4860), .B(n4861), .Z(n4820) );
  AND U5208 ( .A(n194), .B(n4862), .Z(n4860) );
  XOR U5209 ( .A(n4863), .B(n4861), .Z(n4862) );
  NANDN U5210 ( .A(n4822), .B(n4824), .Z(n4838) );
  XOR U5211 ( .A(n4864), .B(n4865), .Z(n4824) );
  AND U5212 ( .A(n194), .B(n4866), .Z(n4864) );
  XOR U5213 ( .A(n4865), .B(n4867), .Z(n4866) );
  XOR U5214 ( .A(n4868), .B(n4869), .Z(n194) );
  AND U5215 ( .A(n4870), .B(n4871), .Z(n4868) );
  XNOR U5216 ( .A(n4869), .B(n4835), .Z(n4871) );
  XNOR U5217 ( .A(n4872), .B(n4873), .Z(n4835) );
  ANDN U5218 ( .B(n4874), .A(n4875), .Z(n4872) );
  XOR U5219 ( .A(n4873), .B(n4876), .Z(n4874) );
  XOR U5220 ( .A(n4869), .B(n4837), .Z(n4870) );
  XOR U5221 ( .A(n4877), .B(n4878), .Z(n4837) );
  AND U5222 ( .A(n198), .B(n4879), .Z(n4877) );
  XOR U5223 ( .A(n4880), .B(n4878), .Z(n4879) );
  XNOR U5224 ( .A(n4881), .B(n4882), .Z(n4869) );
  NAND U5225 ( .A(n4883), .B(n4884), .Z(n4882) );
  XOR U5226 ( .A(n4885), .B(n4861), .Z(n4884) );
  XOR U5227 ( .A(n4875), .B(n4876), .Z(n4861) );
  XOR U5228 ( .A(n4886), .B(n4887), .Z(n4876) );
  ANDN U5229 ( .B(n4888), .A(n4889), .Z(n4886) );
  XOR U5230 ( .A(n4887), .B(n4890), .Z(n4888) );
  XOR U5231 ( .A(n4891), .B(n4892), .Z(n4875) );
  XOR U5232 ( .A(n4893), .B(n4894), .Z(n4892) );
  ANDN U5233 ( .B(n4895), .A(n4896), .Z(n4893) );
  XOR U5234 ( .A(n4897), .B(n4894), .Z(n4895) );
  IV U5235 ( .A(n4873), .Z(n4891) );
  XOR U5236 ( .A(n4898), .B(n4899), .Z(n4873) );
  ANDN U5237 ( .B(n4900), .A(n4901), .Z(n4898) );
  XOR U5238 ( .A(n4899), .B(n4902), .Z(n4900) );
  IV U5239 ( .A(n4881), .Z(n4885) );
  XOR U5240 ( .A(n4881), .B(n4863), .Z(n4883) );
  XOR U5241 ( .A(n4903), .B(n4904), .Z(n4863) );
  AND U5242 ( .A(n198), .B(n4905), .Z(n4903) );
  XOR U5243 ( .A(n4906), .B(n4904), .Z(n4905) );
  NANDN U5244 ( .A(n4865), .B(n4867), .Z(n4881) );
  XOR U5245 ( .A(n4907), .B(n4908), .Z(n4867) );
  AND U5246 ( .A(n198), .B(n4909), .Z(n4907) );
  XOR U5247 ( .A(n4908), .B(n4910), .Z(n4909) );
  XOR U5248 ( .A(n4911), .B(n4912), .Z(n198) );
  AND U5249 ( .A(n4913), .B(n4914), .Z(n4911) );
  XNOR U5250 ( .A(n4912), .B(n4878), .Z(n4914) );
  XNOR U5251 ( .A(n4915), .B(n4916), .Z(n4878) );
  ANDN U5252 ( .B(n4917), .A(n4918), .Z(n4915) );
  XOR U5253 ( .A(n4916), .B(n4919), .Z(n4917) );
  XOR U5254 ( .A(n4912), .B(n4880), .Z(n4913) );
  XOR U5255 ( .A(n4920), .B(n4921), .Z(n4880) );
  AND U5256 ( .A(n202), .B(n4922), .Z(n4920) );
  XOR U5257 ( .A(n4923), .B(n4921), .Z(n4922) );
  XNOR U5258 ( .A(n4924), .B(n4925), .Z(n4912) );
  NAND U5259 ( .A(n4926), .B(n4927), .Z(n4925) );
  XOR U5260 ( .A(n4928), .B(n4904), .Z(n4927) );
  XOR U5261 ( .A(n4918), .B(n4919), .Z(n4904) );
  XOR U5262 ( .A(n4929), .B(n4930), .Z(n4919) );
  ANDN U5263 ( .B(n4931), .A(n4932), .Z(n4929) );
  XOR U5264 ( .A(n4930), .B(n4933), .Z(n4931) );
  XOR U5265 ( .A(n4934), .B(n4935), .Z(n4918) );
  XOR U5266 ( .A(n4936), .B(n4937), .Z(n4935) );
  ANDN U5267 ( .B(n4938), .A(n4939), .Z(n4936) );
  XOR U5268 ( .A(n4940), .B(n4937), .Z(n4938) );
  IV U5269 ( .A(n4916), .Z(n4934) );
  XOR U5270 ( .A(n4941), .B(n4942), .Z(n4916) );
  ANDN U5271 ( .B(n4943), .A(n4944), .Z(n4941) );
  XOR U5272 ( .A(n4942), .B(n4945), .Z(n4943) );
  IV U5273 ( .A(n4924), .Z(n4928) );
  XOR U5274 ( .A(n4924), .B(n4906), .Z(n4926) );
  XOR U5275 ( .A(n4946), .B(n4947), .Z(n4906) );
  AND U5276 ( .A(n202), .B(n4948), .Z(n4946) );
  XOR U5277 ( .A(n4949), .B(n4947), .Z(n4948) );
  NANDN U5278 ( .A(n4908), .B(n4910), .Z(n4924) );
  XOR U5279 ( .A(n4950), .B(n4951), .Z(n4910) );
  AND U5280 ( .A(n202), .B(n4952), .Z(n4950) );
  XOR U5281 ( .A(n4951), .B(n4953), .Z(n4952) );
  XOR U5282 ( .A(n4954), .B(n4955), .Z(n202) );
  AND U5283 ( .A(n4956), .B(n4957), .Z(n4954) );
  XNOR U5284 ( .A(n4955), .B(n4921), .Z(n4957) );
  XNOR U5285 ( .A(n4958), .B(n4959), .Z(n4921) );
  ANDN U5286 ( .B(n4960), .A(n4961), .Z(n4958) );
  XOR U5287 ( .A(n4959), .B(n4962), .Z(n4960) );
  XOR U5288 ( .A(n4955), .B(n4923), .Z(n4956) );
  XOR U5289 ( .A(n4963), .B(n4964), .Z(n4923) );
  AND U5290 ( .A(n206), .B(n4965), .Z(n4963) );
  XOR U5291 ( .A(n4966), .B(n4964), .Z(n4965) );
  XNOR U5292 ( .A(n4967), .B(n4968), .Z(n4955) );
  NAND U5293 ( .A(n4969), .B(n4970), .Z(n4968) );
  XOR U5294 ( .A(n4971), .B(n4947), .Z(n4970) );
  XOR U5295 ( .A(n4961), .B(n4962), .Z(n4947) );
  XOR U5296 ( .A(n4972), .B(n4973), .Z(n4962) );
  ANDN U5297 ( .B(n4974), .A(n4975), .Z(n4972) );
  XOR U5298 ( .A(n4973), .B(n4976), .Z(n4974) );
  XOR U5299 ( .A(n4977), .B(n4978), .Z(n4961) );
  XOR U5300 ( .A(n4979), .B(n4980), .Z(n4978) );
  ANDN U5301 ( .B(n4981), .A(n4982), .Z(n4979) );
  XOR U5302 ( .A(n4983), .B(n4980), .Z(n4981) );
  IV U5303 ( .A(n4959), .Z(n4977) );
  XOR U5304 ( .A(n4984), .B(n4985), .Z(n4959) );
  ANDN U5305 ( .B(n4986), .A(n4987), .Z(n4984) );
  XOR U5306 ( .A(n4985), .B(n4988), .Z(n4986) );
  IV U5307 ( .A(n4967), .Z(n4971) );
  XOR U5308 ( .A(n4967), .B(n4949), .Z(n4969) );
  XOR U5309 ( .A(n4989), .B(n4990), .Z(n4949) );
  AND U5310 ( .A(n206), .B(n4991), .Z(n4989) );
  XOR U5311 ( .A(n4992), .B(n4990), .Z(n4991) );
  NANDN U5312 ( .A(n4951), .B(n4953), .Z(n4967) );
  XOR U5313 ( .A(n4993), .B(n4994), .Z(n4953) );
  AND U5314 ( .A(n206), .B(n4995), .Z(n4993) );
  XOR U5315 ( .A(n4994), .B(n4996), .Z(n4995) );
  XOR U5316 ( .A(n4997), .B(n4998), .Z(n206) );
  AND U5317 ( .A(n4999), .B(n5000), .Z(n4997) );
  XNOR U5318 ( .A(n4998), .B(n4964), .Z(n5000) );
  XNOR U5319 ( .A(n5001), .B(n5002), .Z(n4964) );
  ANDN U5320 ( .B(n5003), .A(n5004), .Z(n5001) );
  XOR U5321 ( .A(n5002), .B(n5005), .Z(n5003) );
  XOR U5322 ( .A(n4998), .B(n4966), .Z(n4999) );
  XOR U5323 ( .A(n5006), .B(n5007), .Z(n4966) );
  AND U5324 ( .A(n210), .B(n5008), .Z(n5006) );
  XOR U5325 ( .A(n5009), .B(n5007), .Z(n5008) );
  XNOR U5326 ( .A(n5010), .B(n5011), .Z(n4998) );
  NAND U5327 ( .A(n5012), .B(n5013), .Z(n5011) );
  XOR U5328 ( .A(n5014), .B(n4990), .Z(n5013) );
  XOR U5329 ( .A(n5004), .B(n5005), .Z(n4990) );
  XOR U5330 ( .A(n5015), .B(n5016), .Z(n5005) );
  ANDN U5331 ( .B(n5017), .A(n5018), .Z(n5015) );
  XOR U5332 ( .A(n5016), .B(n5019), .Z(n5017) );
  XOR U5333 ( .A(n5020), .B(n5021), .Z(n5004) );
  XOR U5334 ( .A(n5022), .B(n5023), .Z(n5021) );
  ANDN U5335 ( .B(n5024), .A(n5025), .Z(n5022) );
  XOR U5336 ( .A(n5026), .B(n5023), .Z(n5024) );
  IV U5337 ( .A(n5002), .Z(n5020) );
  XOR U5338 ( .A(n5027), .B(n5028), .Z(n5002) );
  ANDN U5339 ( .B(n5029), .A(n5030), .Z(n5027) );
  XOR U5340 ( .A(n5028), .B(n5031), .Z(n5029) );
  IV U5341 ( .A(n5010), .Z(n5014) );
  XOR U5342 ( .A(n5010), .B(n4992), .Z(n5012) );
  XOR U5343 ( .A(n5032), .B(n5033), .Z(n4992) );
  AND U5344 ( .A(n210), .B(n5034), .Z(n5032) );
  XOR U5345 ( .A(n5035), .B(n5033), .Z(n5034) );
  NANDN U5346 ( .A(n4994), .B(n4996), .Z(n5010) );
  XOR U5347 ( .A(n5036), .B(n5037), .Z(n4996) );
  AND U5348 ( .A(n210), .B(n5038), .Z(n5036) );
  XOR U5349 ( .A(n5037), .B(n5039), .Z(n5038) );
  XOR U5350 ( .A(n5040), .B(n5041), .Z(n210) );
  AND U5351 ( .A(n5042), .B(n5043), .Z(n5040) );
  XNOR U5352 ( .A(n5041), .B(n5007), .Z(n5043) );
  XNOR U5353 ( .A(n5044), .B(n5045), .Z(n5007) );
  ANDN U5354 ( .B(n5046), .A(n5047), .Z(n5044) );
  XOR U5355 ( .A(n5045), .B(n5048), .Z(n5046) );
  XOR U5356 ( .A(n5041), .B(n5009), .Z(n5042) );
  XOR U5357 ( .A(n5049), .B(n5050), .Z(n5009) );
  AND U5358 ( .A(n214), .B(n5051), .Z(n5049) );
  XOR U5359 ( .A(n5052), .B(n5050), .Z(n5051) );
  XNOR U5360 ( .A(n5053), .B(n5054), .Z(n5041) );
  NAND U5361 ( .A(n5055), .B(n5056), .Z(n5054) );
  XOR U5362 ( .A(n5057), .B(n5033), .Z(n5056) );
  XOR U5363 ( .A(n5047), .B(n5048), .Z(n5033) );
  XOR U5364 ( .A(n5058), .B(n5059), .Z(n5048) );
  ANDN U5365 ( .B(n5060), .A(n5061), .Z(n5058) );
  XOR U5366 ( .A(n5059), .B(n5062), .Z(n5060) );
  XOR U5367 ( .A(n5063), .B(n5064), .Z(n5047) );
  XOR U5368 ( .A(n5065), .B(n5066), .Z(n5064) );
  ANDN U5369 ( .B(n5067), .A(n5068), .Z(n5065) );
  XOR U5370 ( .A(n5069), .B(n5066), .Z(n5067) );
  IV U5371 ( .A(n5045), .Z(n5063) );
  XOR U5372 ( .A(n5070), .B(n5071), .Z(n5045) );
  ANDN U5373 ( .B(n5072), .A(n5073), .Z(n5070) );
  XOR U5374 ( .A(n5071), .B(n5074), .Z(n5072) );
  IV U5375 ( .A(n5053), .Z(n5057) );
  XOR U5376 ( .A(n5053), .B(n5035), .Z(n5055) );
  XOR U5377 ( .A(n5075), .B(n5076), .Z(n5035) );
  AND U5378 ( .A(n214), .B(n5077), .Z(n5075) );
  XOR U5379 ( .A(n5078), .B(n5076), .Z(n5077) );
  NANDN U5380 ( .A(n5037), .B(n5039), .Z(n5053) );
  XOR U5381 ( .A(n5079), .B(n5080), .Z(n5039) );
  AND U5382 ( .A(n214), .B(n5081), .Z(n5079) );
  XOR U5383 ( .A(n5080), .B(n5082), .Z(n5081) );
  XOR U5384 ( .A(n5083), .B(n5084), .Z(n214) );
  AND U5385 ( .A(n5085), .B(n5086), .Z(n5083) );
  XNOR U5386 ( .A(n5084), .B(n5050), .Z(n5086) );
  XNOR U5387 ( .A(n5087), .B(n5088), .Z(n5050) );
  ANDN U5388 ( .B(n5089), .A(n5090), .Z(n5087) );
  XOR U5389 ( .A(n5088), .B(n5091), .Z(n5089) );
  XOR U5390 ( .A(n5084), .B(n5052), .Z(n5085) );
  XOR U5391 ( .A(n5092), .B(n5093), .Z(n5052) );
  AND U5392 ( .A(n218), .B(n5094), .Z(n5092) );
  XOR U5393 ( .A(n5095), .B(n5093), .Z(n5094) );
  XNOR U5394 ( .A(n5096), .B(n5097), .Z(n5084) );
  NAND U5395 ( .A(n5098), .B(n5099), .Z(n5097) );
  XOR U5396 ( .A(n5100), .B(n5076), .Z(n5099) );
  XOR U5397 ( .A(n5090), .B(n5091), .Z(n5076) );
  XOR U5398 ( .A(n5101), .B(n5102), .Z(n5091) );
  ANDN U5399 ( .B(n5103), .A(n5104), .Z(n5101) );
  XOR U5400 ( .A(n5102), .B(n5105), .Z(n5103) );
  XOR U5401 ( .A(n5106), .B(n5107), .Z(n5090) );
  XOR U5402 ( .A(n5108), .B(n5109), .Z(n5107) );
  ANDN U5403 ( .B(n5110), .A(n5111), .Z(n5108) );
  XOR U5404 ( .A(n5112), .B(n5109), .Z(n5110) );
  IV U5405 ( .A(n5088), .Z(n5106) );
  XOR U5406 ( .A(n5113), .B(n5114), .Z(n5088) );
  ANDN U5407 ( .B(n5115), .A(n5116), .Z(n5113) );
  XOR U5408 ( .A(n5114), .B(n5117), .Z(n5115) );
  IV U5409 ( .A(n5096), .Z(n5100) );
  XOR U5410 ( .A(n5096), .B(n5078), .Z(n5098) );
  XOR U5411 ( .A(n5118), .B(n5119), .Z(n5078) );
  AND U5412 ( .A(n218), .B(n5120), .Z(n5118) );
  XOR U5413 ( .A(n5121), .B(n5119), .Z(n5120) );
  NANDN U5414 ( .A(n5080), .B(n5082), .Z(n5096) );
  XOR U5415 ( .A(n5122), .B(n5123), .Z(n5082) );
  AND U5416 ( .A(n218), .B(n5124), .Z(n5122) );
  XOR U5417 ( .A(n5123), .B(n5125), .Z(n5124) );
  XOR U5418 ( .A(n5126), .B(n5127), .Z(n218) );
  AND U5419 ( .A(n5128), .B(n5129), .Z(n5126) );
  XNOR U5420 ( .A(n5127), .B(n5093), .Z(n5129) );
  XNOR U5421 ( .A(n5130), .B(n5131), .Z(n5093) );
  ANDN U5422 ( .B(n5132), .A(n5133), .Z(n5130) );
  XOR U5423 ( .A(n5131), .B(n5134), .Z(n5132) );
  XOR U5424 ( .A(n5127), .B(n5095), .Z(n5128) );
  XOR U5425 ( .A(n5135), .B(n5136), .Z(n5095) );
  AND U5426 ( .A(n222), .B(n5137), .Z(n5135) );
  XOR U5427 ( .A(n5138), .B(n5136), .Z(n5137) );
  XNOR U5428 ( .A(n5139), .B(n5140), .Z(n5127) );
  NAND U5429 ( .A(n5141), .B(n5142), .Z(n5140) );
  XOR U5430 ( .A(n5143), .B(n5119), .Z(n5142) );
  XOR U5431 ( .A(n5133), .B(n5134), .Z(n5119) );
  XOR U5432 ( .A(n5144), .B(n5145), .Z(n5134) );
  ANDN U5433 ( .B(n5146), .A(n5147), .Z(n5144) );
  XOR U5434 ( .A(n5145), .B(n5148), .Z(n5146) );
  XOR U5435 ( .A(n5149), .B(n5150), .Z(n5133) );
  XOR U5436 ( .A(n5151), .B(n5152), .Z(n5150) );
  ANDN U5437 ( .B(n5153), .A(n5154), .Z(n5151) );
  XOR U5438 ( .A(n5155), .B(n5152), .Z(n5153) );
  IV U5439 ( .A(n5131), .Z(n5149) );
  XOR U5440 ( .A(n5156), .B(n5157), .Z(n5131) );
  ANDN U5441 ( .B(n5158), .A(n5159), .Z(n5156) );
  XOR U5442 ( .A(n5157), .B(n5160), .Z(n5158) );
  IV U5443 ( .A(n5139), .Z(n5143) );
  XOR U5444 ( .A(n5139), .B(n5121), .Z(n5141) );
  XOR U5445 ( .A(n5161), .B(n5162), .Z(n5121) );
  AND U5446 ( .A(n222), .B(n5163), .Z(n5161) );
  XOR U5447 ( .A(n5164), .B(n5162), .Z(n5163) );
  NANDN U5448 ( .A(n5123), .B(n5125), .Z(n5139) );
  XOR U5449 ( .A(n5165), .B(n5166), .Z(n5125) );
  AND U5450 ( .A(n222), .B(n5167), .Z(n5165) );
  XOR U5451 ( .A(n5166), .B(n5168), .Z(n5167) );
  XOR U5452 ( .A(n5169), .B(n5170), .Z(n222) );
  AND U5453 ( .A(n5171), .B(n5172), .Z(n5169) );
  XNOR U5454 ( .A(n5170), .B(n5136), .Z(n5172) );
  XNOR U5455 ( .A(n5173), .B(n5174), .Z(n5136) );
  ANDN U5456 ( .B(n5175), .A(n5176), .Z(n5173) );
  XOR U5457 ( .A(n5174), .B(n5177), .Z(n5175) );
  XOR U5458 ( .A(n5170), .B(n5138), .Z(n5171) );
  XOR U5459 ( .A(n5178), .B(n5179), .Z(n5138) );
  AND U5460 ( .A(n226), .B(n5180), .Z(n5178) );
  XOR U5461 ( .A(n5181), .B(n5179), .Z(n5180) );
  XNOR U5462 ( .A(n5182), .B(n5183), .Z(n5170) );
  NAND U5463 ( .A(n5184), .B(n5185), .Z(n5183) );
  XOR U5464 ( .A(n5186), .B(n5162), .Z(n5185) );
  XOR U5465 ( .A(n5176), .B(n5177), .Z(n5162) );
  XOR U5466 ( .A(n5187), .B(n5188), .Z(n5177) );
  ANDN U5467 ( .B(n5189), .A(n5190), .Z(n5187) );
  XOR U5468 ( .A(n5188), .B(n5191), .Z(n5189) );
  XOR U5469 ( .A(n5192), .B(n5193), .Z(n5176) );
  XOR U5470 ( .A(n5194), .B(n5195), .Z(n5193) );
  ANDN U5471 ( .B(n5196), .A(n5197), .Z(n5194) );
  XOR U5472 ( .A(n5198), .B(n5195), .Z(n5196) );
  IV U5473 ( .A(n5174), .Z(n5192) );
  XOR U5474 ( .A(n5199), .B(n5200), .Z(n5174) );
  ANDN U5475 ( .B(n5201), .A(n5202), .Z(n5199) );
  XOR U5476 ( .A(n5200), .B(n5203), .Z(n5201) );
  IV U5477 ( .A(n5182), .Z(n5186) );
  XOR U5478 ( .A(n5182), .B(n5164), .Z(n5184) );
  XOR U5479 ( .A(n5204), .B(n5205), .Z(n5164) );
  AND U5480 ( .A(n226), .B(n5206), .Z(n5204) );
  XOR U5481 ( .A(n5207), .B(n5205), .Z(n5206) );
  NANDN U5482 ( .A(n5166), .B(n5168), .Z(n5182) );
  XOR U5483 ( .A(n5208), .B(n5209), .Z(n5168) );
  AND U5484 ( .A(n226), .B(n5210), .Z(n5208) );
  XOR U5485 ( .A(n5209), .B(n5211), .Z(n5210) );
  XOR U5486 ( .A(n5212), .B(n5213), .Z(n226) );
  AND U5487 ( .A(n5214), .B(n5215), .Z(n5212) );
  XNOR U5488 ( .A(n5213), .B(n5179), .Z(n5215) );
  XNOR U5489 ( .A(n5216), .B(n5217), .Z(n5179) );
  ANDN U5490 ( .B(n5218), .A(n5219), .Z(n5216) );
  XOR U5491 ( .A(n5217), .B(n5220), .Z(n5218) );
  XOR U5492 ( .A(n5213), .B(n5181), .Z(n5214) );
  XOR U5493 ( .A(n5221), .B(n5222), .Z(n5181) );
  AND U5494 ( .A(n230), .B(n5223), .Z(n5221) );
  XOR U5495 ( .A(n5224), .B(n5222), .Z(n5223) );
  XNOR U5496 ( .A(n5225), .B(n5226), .Z(n5213) );
  NAND U5497 ( .A(n5227), .B(n5228), .Z(n5226) );
  XOR U5498 ( .A(n5229), .B(n5205), .Z(n5228) );
  XOR U5499 ( .A(n5219), .B(n5220), .Z(n5205) );
  XOR U5500 ( .A(n5230), .B(n5231), .Z(n5220) );
  ANDN U5501 ( .B(n5232), .A(n5233), .Z(n5230) );
  XOR U5502 ( .A(n5231), .B(n5234), .Z(n5232) );
  XOR U5503 ( .A(n5235), .B(n5236), .Z(n5219) );
  XOR U5504 ( .A(n5237), .B(n5238), .Z(n5236) );
  ANDN U5505 ( .B(n5239), .A(n5240), .Z(n5237) );
  XOR U5506 ( .A(n5241), .B(n5238), .Z(n5239) );
  IV U5507 ( .A(n5217), .Z(n5235) );
  XOR U5508 ( .A(n5242), .B(n5243), .Z(n5217) );
  ANDN U5509 ( .B(n5244), .A(n5245), .Z(n5242) );
  XOR U5510 ( .A(n5243), .B(n5246), .Z(n5244) );
  IV U5511 ( .A(n5225), .Z(n5229) );
  XOR U5512 ( .A(n5225), .B(n5207), .Z(n5227) );
  XOR U5513 ( .A(n5247), .B(n5248), .Z(n5207) );
  AND U5514 ( .A(n230), .B(n5249), .Z(n5247) );
  XOR U5515 ( .A(n5250), .B(n5248), .Z(n5249) );
  NANDN U5516 ( .A(n5209), .B(n5211), .Z(n5225) );
  XOR U5517 ( .A(n5251), .B(n5252), .Z(n5211) );
  AND U5518 ( .A(n230), .B(n5253), .Z(n5251) );
  XOR U5519 ( .A(n5252), .B(n5254), .Z(n5253) );
  XOR U5520 ( .A(n5255), .B(n5256), .Z(n230) );
  AND U5521 ( .A(n5257), .B(n5258), .Z(n5255) );
  XNOR U5522 ( .A(n5256), .B(n5222), .Z(n5258) );
  XNOR U5523 ( .A(n5259), .B(n5260), .Z(n5222) );
  ANDN U5524 ( .B(n5261), .A(n5262), .Z(n5259) );
  XOR U5525 ( .A(n5260), .B(n5263), .Z(n5261) );
  XOR U5526 ( .A(n5256), .B(n5224), .Z(n5257) );
  XOR U5527 ( .A(n5264), .B(n5265), .Z(n5224) );
  AND U5528 ( .A(n234), .B(n5266), .Z(n5264) );
  XOR U5529 ( .A(n5267), .B(n5265), .Z(n5266) );
  XNOR U5530 ( .A(n5268), .B(n5269), .Z(n5256) );
  NAND U5531 ( .A(n5270), .B(n5271), .Z(n5269) );
  XOR U5532 ( .A(n5272), .B(n5248), .Z(n5271) );
  XOR U5533 ( .A(n5262), .B(n5263), .Z(n5248) );
  XOR U5534 ( .A(n5273), .B(n5274), .Z(n5263) );
  ANDN U5535 ( .B(n5275), .A(n5276), .Z(n5273) );
  XOR U5536 ( .A(n5274), .B(n5277), .Z(n5275) );
  XOR U5537 ( .A(n5278), .B(n5279), .Z(n5262) );
  XOR U5538 ( .A(n5280), .B(n5281), .Z(n5279) );
  ANDN U5539 ( .B(n5282), .A(n5283), .Z(n5280) );
  XOR U5540 ( .A(n5284), .B(n5281), .Z(n5282) );
  IV U5541 ( .A(n5260), .Z(n5278) );
  XOR U5542 ( .A(n5285), .B(n5286), .Z(n5260) );
  ANDN U5543 ( .B(n5287), .A(n5288), .Z(n5285) );
  XOR U5544 ( .A(n5286), .B(n5289), .Z(n5287) );
  IV U5545 ( .A(n5268), .Z(n5272) );
  XOR U5546 ( .A(n5268), .B(n5250), .Z(n5270) );
  XOR U5547 ( .A(n5290), .B(n5291), .Z(n5250) );
  AND U5548 ( .A(n234), .B(n5292), .Z(n5290) );
  XOR U5549 ( .A(n5293), .B(n5291), .Z(n5292) );
  NANDN U5550 ( .A(n5252), .B(n5254), .Z(n5268) );
  XOR U5551 ( .A(n5294), .B(n5295), .Z(n5254) );
  AND U5552 ( .A(n234), .B(n5296), .Z(n5294) );
  XOR U5553 ( .A(n5295), .B(n5297), .Z(n5296) );
  XOR U5554 ( .A(n5298), .B(n5299), .Z(n234) );
  AND U5555 ( .A(n5300), .B(n5301), .Z(n5298) );
  XNOR U5556 ( .A(n5299), .B(n5265), .Z(n5301) );
  XNOR U5557 ( .A(n5302), .B(n5303), .Z(n5265) );
  ANDN U5558 ( .B(n5304), .A(n5305), .Z(n5302) );
  XOR U5559 ( .A(n5303), .B(n5306), .Z(n5304) );
  XOR U5560 ( .A(n5299), .B(n5267), .Z(n5300) );
  XOR U5561 ( .A(n5307), .B(n5308), .Z(n5267) );
  AND U5562 ( .A(n238), .B(n5309), .Z(n5307) );
  XOR U5563 ( .A(n5310), .B(n5308), .Z(n5309) );
  XNOR U5564 ( .A(n5311), .B(n5312), .Z(n5299) );
  NAND U5565 ( .A(n5313), .B(n5314), .Z(n5312) );
  XOR U5566 ( .A(n5315), .B(n5291), .Z(n5314) );
  XOR U5567 ( .A(n5305), .B(n5306), .Z(n5291) );
  XOR U5568 ( .A(n5316), .B(n5317), .Z(n5306) );
  ANDN U5569 ( .B(n5318), .A(n5319), .Z(n5316) );
  XOR U5570 ( .A(n5317), .B(n5320), .Z(n5318) );
  XOR U5571 ( .A(n5321), .B(n5322), .Z(n5305) );
  XOR U5572 ( .A(n5323), .B(n5324), .Z(n5322) );
  ANDN U5573 ( .B(n5325), .A(n5326), .Z(n5323) );
  XOR U5574 ( .A(n5327), .B(n5324), .Z(n5325) );
  IV U5575 ( .A(n5303), .Z(n5321) );
  XOR U5576 ( .A(n5328), .B(n5329), .Z(n5303) );
  ANDN U5577 ( .B(n5330), .A(n5331), .Z(n5328) );
  XOR U5578 ( .A(n5329), .B(n5332), .Z(n5330) );
  IV U5579 ( .A(n5311), .Z(n5315) );
  XOR U5580 ( .A(n5311), .B(n5293), .Z(n5313) );
  XOR U5581 ( .A(n5333), .B(n5334), .Z(n5293) );
  AND U5582 ( .A(n238), .B(n5335), .Z(n5333) );
  XOR U5583 ( .A(n5336), .B(n5334), .Z(n5335) );
  NANDN U5584 ( .A(n5295), .B(n5297), .Z(n5311) );
  XOR U5585 ( .A(n5337), .B(n5338), .Z(n5297) );
  AND U5586 ( .A(n238), .B(n5339), .Z(n5337) );
  XOR U5587 ( .A(n5338), .B(n5340), .Z(n5339) );
  XOR U5588 ( .A(n5341), .B(n5342), .Z(n238) );
  AND U5589 ( .A(n5343), .B(n5344), .Z(n5341) );
  XNOR U5590 ( .A(n5342), .B(n5308), .Z(n5344) );
  XNOR U5591 ( .A(n5345), .B(n5346), .Z(n5308) );
  ANDN U5592 ( .B(n5347), .A(n5348), .Z(n5345) );
  XOR U5593 ( .A(n5346), .B(n5349), .Z(n5347) );
  XOR U5594 ( .A(n5342), .B(n5310), .Z(n5343) );
  XOR U5595 ( .A(n5350), .B(n5351), .Z(n5310) );
  AND U5596 ( .A(n242), .B(n5352), .Z(n5350) );
  XOR U5597 ( .A(n5353), .B(n5351), .Z(n5352) );
  XNOR U5598 ( .A(n5354), .B(n5355), .Z(n5342) );
  NAND U5599 ( .A(n5356), .B(n5357), .Z(n5355) );
  XOR U5600 ( .A(n5358), .B(n5334), .Z(n5357) );
  XOR U5601 ( .A(n5348), .B(n5349), .Z(n5334) );
  XOR U5602 ( .A(n5359), .B(n5360), .Z(n5349) );
  ANDN U5603 ( .B(n5361), .A(n5362), .Z(n5359) );
  XOR U5604 ( .A(n5360), .B(n5363), .Z(n5361) );
  XOR U5605 ( .A(n5364), .B(n5365), .Z(n5348) );
  XOR U5606 ( .A(n5366), .B(n5367), .Z(n5365) );
  ANDN U5607 ( .B(n5368), .A(n5369), .Z(n5366) );
  XOR U5608 ( .A(n5370), .B(n5367), .Z(n5368) );
  IV U5609 ( .A(n5346), .Z(n5364) );
  XOR U5610 ( .A(n5371), .B(n5372), .Z(n5346) );
  ANDN U5611 ( .B(n5373), .A(n5374), .Z(n5371) );
  XOR U5612 ( .A(n5372), .B(n5375), .Z(n5373) );
  IV U5613 ( .A(n5354), .Z(n5358) );
  XOR U5614 ( .A(n5354), .B(n5336), .Z(n5356) );
  XOR U5615 ( .A(n5376), .B(n5377), .Z(n5336) );
  AND U5616 ( .A(n242), .B(n5378), .Z(n5376) );
  XOR U5617 ( .A(n5379), .B(n5377), .Z(n5378) );
  NANDN U5618 ( .A(n5338), .B(n5340), .Z(n5354) );
  XOR U5619 ( .A(n5380), .B(n5381), .Z(n5340) );
  AND U5620 ( .A(n242), .B(n5382), .Z(n5380) );
  XOR U5621 ( .A(n5381), .B(n5383), .Z(n5382) );
  XOR U5622 ( .A(n5384), .B(n5385), .Z(n242) );
  AND U5623 ( .A(n5386), .B(n5387), .Z(n5384) );
  XNOR U5624 ( .A(n5385), .B(n5351), .Z(n5387) );
  XNOR U5625 ( .A(n5388), .B(n5389), .Z(n5351) );
  ANDN U5626 ( .B(n5390), .A(n5391), .Z(n5388) );
  XOR U5627 ( .A(n5389), .B(n5392), .Z(n5390) );
  XOR U5628 ( .A(n5385), .B(n5353), .Z(n5386) );
  XOR U5629 ( .A(n5393), .B(n5394), .Z(n5353) );
  AND U5630 ( .A(n246), .B(n5395), .Z(n5393) );
  XOR U5631 ( .A(n5396), .B(n5394), .Z(n5395) );
  XNOR U5632 ( .A(n5397), .B(n5398), .Z(n5385) );
  NAND U5633 ( .A(n5399), .B(n5400), .Z(n5398) );
  XOR U5634 ( .A(n5401), .B(n5377), .Z(n5400) );
  XOR U5635 ( .A(n5391), .B(n5392), .Z(n5377) );
  XOR U5636 ( .A(n5402), .B(n5403), .Z(n5392) );
  ANDN U5637 ( .B(n5404), .A(n5405), .Z(n5402) );
  XOR U5638 ( .A(n5403), .B(n5406), .Z(n5404) );
  XOR U5639 ( .A(n5407), .B(n5408), .Z(n5391) );
  XOR U5640 ( .A(n5409), .B(n5410), .Z(n5408) );
  ANDN U5641 ( .B(n5411), .A(n5412), .Z(n5409) );
  XOR U5642 ( .A(n5413), .B(n5410), .Z(n5411) );
  IV U5643 ( .A(n5389), .Z(n5407) );
  XOR U5644 ( .A(n5414), .B(n5415), .Z(n5389) );
  ANDN U5645 ( .B(n5416), .A(n5417), .Z(n5414) );
  XOR U5646 ( .A(n5415), .B(n5418), .Z(n5416) );
  IV U5647 ( .A(n5397), .Z(n5401) );
  XOR U5648 ( .A(n5397), .B(n5379), .Z(n5399) );
  XOR U5649 ( .A(n5419), .B(n5420), .Z(n5379) );
  AND U5650 ( .A(n246), .B(n5421), .Z(n5419) );
  XOR U5651 ( .A(n5422), .B(n5420), .Z(n5421) );
  NANDN U5652 ( .A(n5381), .B(n5383), .Z(n5397) );
  XOR U5653 ( .A(n5423), .B(n5424), .Z(n5383) );
  AND U5654 ( .A(n246), .B(n5425), .Z(n5423) );
  XOR U5655 ( .A(n5424), .B(n5426), .Z(n5425) );
  XOR U5656 ( .A(n5427), .B(n5428), .Z(n246) );
  AND U5657 ( .A(n5429), .B(n5430), .Z(n5427) );
  XNOR U5658 ( .A(n5428), .B(n5394), .Z(n5430) );
  XNOR U5659 ( .A(n5431), .B(n5432), .Z(n5394) );
  ANDN U5660 ( .B(n5433), .A(n5434), .Z(n5431) );
  XOR U5661 ( .A(n5432), .B(n5435), .Z(n5433) );
  XOR U5662 ( .A(n5428), .B(n5396), .Z(n5429) );
  XOR U5663 ( .A(n5436), .B(n5437), .Z(n5396) );
  AND U5664 ( .A(n250), .B(n5438), .Z(n5436) );
  XOR U5665 ( .A(n5439), .B(n5437), .Z(n5438) );
  XNOR U5666 ( .A(n5440), .B(n5441), .Z(n5428) );
  NAND U5667 ( .A(n5442), .B(n5443), .Z(n5441) );
  XOR U5668 ( .A(n5444), .B(n5420), .Z(n5443) );
  XOR U5669 ( .A(n5434), .B(n5435), .Z(n5420) );
  XOR U5670 ( .A(n5445), .B(n5446), .Z(n5435) );
  ANDN U5671 ( .B(n5447), .A(n5448), .Z(n5445) );
  XOR U5672 ( .A(n5446), .B(n5449), .Z(n5447) );
  XOR U5673 ( .A(n5450), .B(n5451), .Z(n5434) );
  XOR U5674 ( .A(n5452), .B(n5453), .Z(n5451) );
  ANDN U5675 ( .B(n5454), .A(n5455), .Z(n5452) );
  XOR U5676 ( .A(n5456), .B(n5453), .Z(n5454) );
  IV U5677 ( .A(n5432), .Z(n5450) );
  XOR U5678 ( .A(n5457), .B(n5458), .Z(n5432) );
  ANDN U5679 ( .B(n5459), .A(n5460), .Z(n5457) );
  XOR U5680 ( .A(n5458), .B(n5461), .Z(n5459) );
  IV U5681 ( .A(n5440), .Z(n5444) );
  XOR U5682 ( .A(n5440), .B(n5422), .Z(n5442) );
  XOR U5683 ( .A(n5462), .B(n5463), .Z(n5422) );
  AND U5684 ( .A(n250), .B(n5464), .Z(n5462) );
  XOR U5685 ( .A(n5465), .B(n5463), .Z(n5464) );
  NANDN U5686 ( .A(n5424), .B(n5426), .Z(n5440) );
  XOR U5687 ( .A(n5466), .B(n5467), .Z(n5426) );
  AND U5688 ( .A(n250), .B(n5468), .Z(n5466) );
  XOR U5689 ( .A(n5467), .B(n5469), .Z(n5468) );
  XOR U5690 ( .A(n5470), .B(n5471), .Z(n250) );
  AND U5691 ( .A(n5472), .B(n5473), .Z(n5470) );
  XNOR U5692 ( .A(n5471), .B(n5437), .Z(n5473) );
  XNOR U5693 ( .A(n5474), .B(n5475), .Z(n5437) );
  ANDN U5694 ( .B(n5476), .A(n5477), .Z(n5474) );
  XOR U5695 ( .A(n5475), .B(n5478), .Z(n5476) );
  XOR U5696 ( .A(n5471), .B(n5439), .Z(n5472) );
  XOR U5697 ( .A(n5479), .B(n5480), .Z(n5439) );
  AND U5698 ( .A(n254), .B(n5481), .Z(n5479) );
  XOR U5699 ( .A(n5482), .B(n5480), .Z(n5481) );
  XNOR U5700 ( .A(n5483), .B(n5484), .Z(n5471) );
  NAND U5701 ( .A(n5485), .B(n5486), .Z(n5484) );
  XOR U5702 ( .A(n5487), .B(n5463), .Z(n5486) );
  XOR U5703 ( .A(n5477), .B(n5478), .Z(n5463) );
  XOR U5704 ( .A(n5488), .B(n5489), .Z(n5478) );
  ANDN U5705 ( .B(n5490), .A(n5491), .Z(n5488) );
  XOR U5706 ( .A(n5489), .B(n5492), .Z(n5490) );
  XOR U5707 ( .A(n5493), .B(n5494), .Z(n5477) );
  XOR U5708 ( .A(n5495), .B(n5496), .Z(n5494) );
  ANDN U5709 ( .B(n5497), .A(n5498), .Z(n5495) );
  XOR U5710 ( .A(n5499), .B(n5496), .Z(n5497) );
  IV U5711 ( .A(n5475), .Z(n5493) );
  XOR U5712 ( .A(n5500), .B(n5501), .Z(n5475) );
  ANDN U5713 ( .B(n5502), .A(n5503), .Z(n5500) );
  XOR U5714 ( .A(n5501), .B(n5504), .Z(n5502) );
  IV U5715 ( .A(n5483), .Z(n5487) );
  XOR U5716 ( .A(n5483), .B(n5465), .Z(n5485) );
  XOR U5717 ( .A(n5505), .B(n5506), .Z(n5465) );
  AND U5718 ( .A(n254), .B(n5507), .Z(n5505) );
  XOR U5719 ( .A(n5508), .B(n5506), .Z(n5507) );
  NANDN U5720 ( .A(n5467), .B(n5469), .Z(n5483) );
  XOR U5721 ( .A(n5509), .B(n5510), .Z(n5469) );
  AND U5722 ( .A(n254), .B(n5511), .Z(n5509) );
  XOR U5723 ( .A(n5510), .B(n5512), .Z(n5511) );
  XOR U5724 ( .A(n5513), .B(n5514), .Z(n254) );
  AND U5725 ( .A(n5515), .B(n5516), .Z(n5513) );
  XNOR U5726 ( .A(n5514), .B(n5480), .Z(n5516) );
  XNOR U5727 ( .A(n5517), .B(n5518), .Z(n5480) );
  ANDN U5728 ( .B(n5519), .A(n5520), .Z(n5517) );
  XOR U5729 ( .A(n5518), .B(n5521), .Z(n5519) );
  XOR U5730 ( .A(n5514), .B(n5482), .Z(n5515) );
  XOR U5731 ( .A(n5522), .B(n5523), .Z(n5482) );
  AND U5732 ( .A(n258), .B(n5524), .Z(n5522) );
  XOR U5733 ( .A(n5525), .B(n5523), .Z(n5524) );
  XNOR U5734 ( .A(n5526), .B(n5527), .Z(n5514) );
  NAND U5735 ( .A(n5528), .B(n5529), .Z(n5527) );
  XOR U5736 ( .A(n5530), .B(n5506), .Z(n5529) );
  XOR U5737 ( .A(n5520), .B(n5521), .Z(n5506) );
  XOR U5738 ( .A(n5531), .B(n5532), .Z(n5521) );
  ANDN U5739 ( .B(n5533), .A(n5534), .Z(n5531) );
  XOR U5740 ( .A(n5532), .B(n5535), .Z(n5533) );
  XOR U5741 ( .A(n5536), .B(n5537), .Z(n5520) );
  XOR U5742 ( .A(n5538), .B(n5539), .Z(n5537) );
  ANDN U5743 ( .B(n5540), .A(n5541), .Z(n5538) );
  XOR U5744 ( .A(n5542), .B(n5539), .Z(n5540) );
  IV U5745 ( .A(n5518), .Z(n5536) );
  XOR U5746 ( .A(n5543), .B(n5544), .Z(n5518) );
  ANDN U5747 ( .B(n5545), .A(n5546), .Z(n5543) );
  XOR U5748 ( .A(n5544), .B(n5547), .Z(n5545) );
  IV U5749 ( .A(n5526), .Z(n5530) );
  XOR U5750 ( .A(n5526), .B(n5508), .Z(n5528) );
  XOR U5751 ( .A(n5548), .B(n5549), .Z(n5508) );
  AND U5752 ( .A(n258), .B(n5550), .Z(n5548) );
  XOR U5753 ( .A(n5551), .B(n5549), .Z(n5550) );
  NANDN U5754 ( .A(n5510), .B(n5512), .Z(n5526) );
  XOR U5755 ( .A(n5552), .B(n5553), .Z(n5512) );
  AND U5756 ( .A(n258), .B(n5554), .Z(n5552) );
  XOR U5757 ( .A(n5553), .B(n5555), .Z(n5554) );
  XOR U5758 ( .A(n5556), .B(n5557), .Z(n258) );
  AND U5759 ( .A(n5558), .B(n5559), .Z(n5556) );
  XNOR U5760 ( .A(n5557), .B(n5523), .Z(n5559) );
  XNOR U5761 ( .A(n5560), .B(n5561), .Z(n5523) );
  ANDN U5762 ( .B(n5562), .A(n5563), .Z(n5560) );
  XOR U5763 ( .A(n5561), .B(n5564), .Z(n5562) );
  XOR U5764 ( .A(n5557), .B(n5525), .Z(n5558) );
  XOR U5765 ( .A(n5565), .B(n5566), .Z(n5525) );
  AND U5766 ( .A(n262), .B(n5567), .Z(n5565) );
  XOR U5767 ( .A(n5568), .B(n5566), .Z(n5567) );
  XNOR U5768 ( .A(n5569), .B(n5570), .Z(n5557) );
  NAND U5769 ( .A(n5571), .B(n5572), .Z(n5570) );
  XOR U5770 ( .A(n5573), .B(n5549), .Z(n5572) );
  XOR U5771 ( .A(n5563), .B(n5564), .Z(n5549) );
  XOR U5772 ( .A(n5574), .B(n5575), .Z(n5564) );
  ANDN U5773 ( .B(n5576), .A(n5577), .Z(n5574) );
  XOR U5774 ( .A(n5575), .B(n5578), .Z(n5576) );
  XOR U5775 ( .A(n5579), .B(n5580), .Z(n5563) );
  XOR U5776 ( .A(n5581), .B(n5582), .Z(n5580) );
  ANDN U5777 ( .B(n5583), .A(n5584), .Z(n5581) );
  XOR U5778 ( .A(n5585), .B(n5582), .Z(n5583) );
  IV U5779 ( .A(n5561), .Z(n5579) );
  XOR U5780 ( .A(n5586), .B(n5587), .Z(n5561) );
  ANDN U5781 ( .B(n5588), .A(n5589), .Z(n5586) );
  XOR U5782 ( .A(n5587), .B(n5590), .Z(n5588) );
  IV U5783 ( .A(n5569), .Z(n5573) );
  XOR U5784 ( .A(n5569), .B(n5551), .Z(n5571) );
  XOR U5785 ( .A(n5591), .B(n5592), .Z(n5551) );
  AND U5786 ( .A(n262), .B(n5593), .Z(n5591) );
  XOR U5787 ( .A(n5594), .B(n5592), .Z(n5593) );
  NANDN U5788 ( .A(n5553), .B(n5555), .Z(n5569) );
  XOR U5789 ( .A(n5595), .B(n5596), .Z(n5555) );
  AND U5790 ( .A(n262), .B(n5597), .Z(n5595) );
  XOR U5791 ( .A(n5596), .B(n5598), .Z(n5597) );
  XOR U5792 ( .A(n5599), .B(n5600), .Z(n262) );
  AND U5793 ( .A(n5601), .B(n5602), .Z(n5599) );
  XNOR U5794 ( .A(n5600), .B(n5566), .Z(n5602) );
  XNOR U5795 ( .A(n5603), .B(n5604), .Z(n5566) );
  ANDN U5796 ( .B(n5605), .A(n5606), .Z(n5603) );
  XOR U5797 ( .A(n5604), .B(n5607), .Z(n5605) );
  XOR U5798 ( .A(n5600), .B(n5568), .Z(n5601) );
  XOR U5799 ( .A(n5608), .B(n5609), .Z(n5568) );
  AND U5800 ( .A(n266), .B(n5610), .Z(n5608) );
  XOR U5801 ( .A(n5611), .B(n5609), .Z(n5610) );
  XNOR U5802 ( .A(n5612), .B(n5613), .Z(n5600) );
  NAND U5803 ( .A(n5614), .B(n5615), .Z(n5613) );
  XOR U5804 ( .A(n5616), .B(n5592), .Z(n5615) );
  XOR U5805 ( .A(n5606), .B(n5607), .Z(n5592) );
  XOR U5806 ( .A(n5617), .B(n5618), .Z(n5607) );
  ANDN U5807 ( .B(n5619), .A(n5620), .Z(n5617) );
  XOR U5808 ( .A(n5618), .B(n5621), .Z(n5619) );
  XOR U5809 ( .A(n5622), .B(n5623), .Z(n5606) );
  XOR U5810 ( .A(n5624), .B(n5625), .Z(n5623) );
  ANDN U5811 ( .B(n5626), .A(n5627), .Z(n5624) );
  XOR U5812 ( .A(n5628), .B(n5625), .Z(n5626) );
  IV U5813 ( .A(n5604), .Z(n5622) );
  XOR U5814 ( .A(n5629), .B(n5630), .Z(n5604) );
  ANDN U5815 ( .B(n5631), .A(n5632), .Z(n5629) );
  XOR U5816 ( .A(n5630), .B(n5633), .Z(n5631) );
  IV U5817 ( .A(n5612), .Z(n5616) );
  XOR U5818 ( .A(n5612), .B(n5594), .Z(n5614) );
  XOR U5819 ( .A(n5634), .B(n5635), .Z(n5594) );
  AND U5820 ( .A(n266), .B(n5636), .Z(n5634) );
  XOR U5821 ( .A(n5637), .B(n5635), .Z(n5636) );
  NANDN U5822 ( .A(n5596), .B(n5598), .Z(n5612) );
  XOR U5823 ( .A(n5638), .B(n5639), .Z(n5598) );
  AND U5824 ( .A(n266), .B(n5640), .Z(n5638) );
  XOR U5825 ( .A(n5639), .B(n5641), .Z(n5640) );
  XOR U5826 ( .A(n5642), .B(n5643), .Z(n266) );
  AND U5827 ( .A(n5644), .B(n5645), .Z(n5642) );
  XNOR U5828 ( .A(n5643), .B(n5609), .Z(n5645) );
  XNOR U5829 ( .A(n5646), .B(n5647), .Z(n5609) );
  ANDN U5830 ( .B(n5648), .A(n5649), .Z(n5646) );
  XOR U5831 ( .A(n5647), .B(n5650), .Z(n5648) );
  XOR U5832 ( .A(n5643), .B(n5611), .Z(n5644) );
  XOR U5833 ( .A(n5651), .B(n5652), .Z(n5611) );
  AND U5834 ( .A(n270), .B(n5653), .Z(n5651) );
  XOR U5835 ( .A(n5654), .B(n5652), .Z(n5653) );
  XNOR U5836 ( .A(n5655), .B(n5656), .Z(n5643) );
  NAND U5837 ( .A(n5657), .B(n5658), .Z(n5656) );
  XOR U5838 ( .A(n5659), .B(n5635), .Z(n5658) );
  XOR U5839 ( .A(n5649), .B(n5650), .Z(n5635) );
  XOR U5840 ( .A(n5660), .B(n5661), .Z(n5650) );
  ANDN U5841 ( .B(n5662), .A(n5663), .Z(n5660) );
  XOR U5842 ( .A(n5661), .B(n5664), .Z(n5662) );
  XOR U5843 ( .A(n5665), .B(n5666), .Z(n5649) );
  XOR U5844 ( .A(n5667), .B(n5668), .Z(n5666) );
  ANDN U5845 ( .B(n5669), .A(n5670), .Z(n5667) );
  XOR U5846 ( .A(n5671), .B(n5668), .Z(n5669) );
  IV U5847 ( .A(n5647), .Z(n5665) );
  XOR U5848 ( .A(n5672), .B(n5673), .Z(n5647) );
  ANDN U5849 ( .B(n5674), .A(n5675), .Z(n5672) );
  XOR U5850 ( .A(n5673), .B(n5676), .Z(n5674) );
  IV U5851 ( .A(n5655), .Z(n5659) );
  XOR U5852 ( .A(n5655), .B(n5637), .Z(n5657) );
  XOR U5853 ( .A(n5677), .B(n5678), .Z(n5637) );
  AND U5854 ( .A(n270), .B(n5679), .Z(n5677) );
  XOR U5855 ( .A(n5680), .B(n5678), .Z(n5679) );
  NANDN U5856 ( .A(n5639), .B(n5641), .Z(n5655) );
  XOR U5857 ( .A(n5681), .B(n5682), .Z(n5641) );
  AND U5858 ( .A(n270), .B(n5683), .Z(n5681) );
  XOR U5859 ( .A(n5682), .B(n5684), .Z(n5683) );
  XOR U5860 ( .A(n5685), .B(n5686), .Z(n270) );
  AND U5861 ( .A(n5687), .B(n5688), .Z(n5685) );
  XNOR U5862 ( .A(n5686), .B(n5652), .Z(n5688) );
  XNOR U5863 ( .A(n5689), .B(n5690), .Z(n5652) );
  ANDN U5864 ( .B(n5691), .A(n5692), .Z(n5689) );
  XOR U5865 ( .A(n5690), .B(n5693), .Z(n5691) );
  XOR U5866 ( .A(n5686), .B(n5654), .Z(n5687) );
  XOR U5867 ( .A(n5694), .B(n5695), .Z(n5654) );
  AND U5868 ( .A(n274), .B(n5696), .Z(n5694) );
  XOR U5869 ( .A(n5697), .B(n5695), .Z(n5696) );
  XNOR U5870 ( .A(n5698), .B(n5699), .Z(n5686) );
  NAND U5871 ( .A(n5700), .B(n5701), .Z(n5699) );
  XOR U5872 ( .A(n5702), .B(n5678), .Z(n5701) );
  XOR U5873 ( .A(n5692), .B(n5693), .Z(n5678) );
  XOR U5874 ( .A(n5703), .B(n5704), .Z(n5693) );
  ANDN U5875 ( .B(n5705), .A(n5706), .Z(n5703) );
  XOR U5876 ( .A(n5704), .B(n5707), .Z(n5705) );
  XOR U5877 ( .A(n5708), .B(n5709), .Z(n5692) );
  XOR U5878 ( .A(n5710), .B(n5711), .Z(n5709) );
  ANDN U5879 ( .B(n5712), .A(n5713), .Z(n5710) );
  XOR U5880 ( .A(n5714), .B(n5711), .Z(n5712) );
  IV U5881 ( .A(n5690), .Z(n5708) );
  XOR U5882 ( .A(n5715), .B(n5716), .Z(n5690) );
  ANDN U5883 ( .B(n5717), .A(n5718), .Z(n5715) );
  XOR U5884 ( .A(n5716), .B(n5719), .Z(n5717) );
  IV U5885 ( .A(n5698), .Z(n5702) );
  XOR U5886 ( .A(n5698), .B(n5680), .Z(n5700) );
  XOR U5887 ( .A(n5720), .B(n5721), .Z(n5680) );
  AND U5888 ( .A(n274), .B(n5722), .Z(n5720) );
  XOR U5889 ( .A(n5723), .B(n5721), .Z(n5722) );
  NANDN U5890 ( .A(n5682), .B(n5684), .Z(n5698) );
  XOR U5891 ( .A(n5724), .B(n5725), .Z(n5684) );
  AND U5892 ( .A(n274), .B(n5726), .Z(n5724) );
  XOR U5893 ( .A(n5725), .B(n5727), .Z(n5726) );
  XOR U5894 ( .A(n5728), .B(n5729), .Z(n274) );
  AND U5895 ( .A(n5730), .B(n5731), .Z(n5728) );
  XNOR U5896 ( .A(n5729), .B(n5695), .Z(n5731) );
  XNOR U5897 ( .A(n5732), .B(n5733), .Z(n5695) );
  ANDN U5898 ( .B(n5734), .A(n5735), .Z(n5732) );
  XOR U5899 ( .A(n5733), .B(n5736), .Z(n5734) );
  XOR U5900 ( .A(n5729), .B(n5697), .Z(n5730) );
  XOR U5901 ( .A(n5737), .B(n5738), .Z(n5697) );
  AND U5902 ( .A(n278), .B(n5739), .Z(n5737) );
  XOR U5903 ( .A(n5740), .B(n5738), .Z(n5739) );
  XNOR U5904 ( .A(n5741), .B(n5742), .Z(n5729) );
  NAND U5905 ( .A(n5743), .B(n5744), .Z(n5742) );
  XOR U5906 ( .A(n5745), .B(n5721), .Z(n5744) );
  XOR U5907 ( .A(n5735), .B(n5736), .Z(n5721) );
  XOR U5908 ( .A(n5746), .B(n5747), .Z(n5736) );
  ANDN U5909 ( .B(n5748), .A(n5749), .Z(n5746) );
  XOR U5910 ( .A(n5747), .B(n5750), .Z(n5748) );
  XOR U5911 ( .A(n5751), .B(n5752), .Z(n5735) );
  XOR U5912 ( .A(n5753), .B(n5754), .Z(n5752) );
  ANDN U5913 ( .B(n5755), .A(n5756), .Z(n5753) );
  XOR U5914 ( .A(n5757), .B(n5754), .Z(n5755) );
  IV U5915 ( .A(n5733), .Z(n5751) );
  XOR U5916 ( .A(n5758), .B(n5759), .Z(n5733) );
  ANDN U5917 ( .B(n5760), .A(n5761), .Z(n5758) );
  XOR U5918 ( .A(n5759), .B(n5762), .Z(n5760) );
  IV U5919 ( .A(n5741), .Z(n5745) );
  XOR U5920 ( .A(n5741), .B(n5723), .Z(n5743) );
  XOR U5921 ( .A(n5763), .B(n5764), .Z(n5723) );
  AND U5922 ( .A(n278), .B(n5765), .Z(n5763) );
  XOR U5923 ( .A(n5766), .B(n5764), .Z(n5765) );
  NANDN U5924 ( .A(n5725), .B(n5727), .Z(n5741) );
  XOR U5925 ( .A(n5767), .B(n5768), .Z(n5727) );
  AND U5926 ( .A(n278), .B(n5769), .Z(n5767) );
  XOR U5927 ( .A(n5768), .B(n5770), .Z(n5769) );
  XOR U5928 ( .A(n5771), .B(n5772), .Z(n278) );
  AND U5929 ( .A(n5773), .B(n5774), .Z(n5771) );
  XNOR U5930 ( .A(n5772), .B(n5738), .Z(n5774) );
  XNOR U5931 ( .A(n5775), .B(n5776), .Z(n5738) );
  ANDN U5932 ( .B(n5777), .A(n5778), .Z(n5775) );
  XOR U5933 ( .A(n5776), .B(n5779), .Z(n5777) );
  XOR U5934 ( .A(n5772), .B(n5740), .Z(n5773) );
  XOR U5935 ( .A(n5780), .B(n5781), .Z(n5740) );
  AND U5936 ( .A(n282), .B(n5782), .Z(n5780) );
  XOR U5937 ( .A(n5783), .B(n5781), .Z(n5782) );
  XNOR U5938 ( .A(n5784), .B(n5785), .Z(n5772) );
  NAND U5939 ( .A(n5786), .B(n5787), .Z(n5785) );
  XOR U5940 ( .A(n5788), .B(n5764), .Z(n5787) );
  XOR U5941 ( .A(n5778), .B(n5779), .Z(n5764) );
  XOR U5942 ( .A(n5789), .B(n5790), .Z(n5779) );
  ANDN U5943 ( .B(n5791), .A(n5792), .Z(n5789) );
  XOR U5944 ( .A(n5790), .B(n5793), .Z(n5791) );
  XOR U5945 ( .A(n5794), .B(n5795), .Z(n5778) );
  XOR U5946 ( .A(n5796), .B(n5797), .Z(n5795) );
  ANDN U5947 ( .B(n5798), .A(n5799), .Z(n5796) );
  XOR U5948 ( .A(n5800), .B(n5797), .Z(n5798) );
  IV U5949 ( .A(n5776), .Z(n5794) );
  XOR U5950 ( .A(n5801), .B(n5802), .Z(n5776) );
  ANDN U5951 ( .B(n5803), .A(n5804), .Z(n5801) );
  XOR U5952 ( .A(n5802), .B(n5805), .Z(n5803) );
  IV U5953 ( .A(n5784), .Z(n5788) );
  XOR U5954 ( .A(n5784), .B(n5766), .Z(n5786) );
  XOR U5955 ( .A(n5806), .B(n5807), .Z(n5766) );
  AND U5956 ( .A(n282), .B(n5808), .Z(n5806) );
  XOR U5957 ( .A(n5809), .B(n5807), .Z(n5808) );
  NANDN U5958 ( .A(n5768), .B(n5770), .Z(n5784) );
  XOR U5959 ( .A(n5810), .B(n5811), .Z(n5770) );
  AND U5960 ( .A(n282), .B(n5812), .Z(n5810) );
  XOR U5961 ( .A(n5811), .B(n5813), .Z(n5812) );
  XOR U5962 ( .A(n5814), .B(n5815), .Z(n282) );
  AND U5963 ( .A(n5816), .B(n5817), .Z(n5814) );
  XNOR U5964 ( .A(n5815), .B(n5781), .Z(n5817) );
  XNOR U5965 ( .A(n5818), .B(n5819), .Z(n5781) );
  ANDN U5966 ( .B(n5820), .A(n5821), .Z(n5818) );
  XOR U5967 ( .A(n5819), .B(n5822), .Z(n5820) );
  XOR U5968 ( .A(n5815), .B(n5783), .Z(n5816) );
  XOR U5969 ( .A(n5823), .B(n5824), .Z(n5783) );
  AND U5970 ( .A(n286), .B(n5825), .Z(n5823) );
  XOR U5971 ( .A(n5826), .B(n5824), .Z(n5825) );
  XNOR U5972 ( .A(n5827), .B(n5828), .Z(n5815) );
  NAND U5973 ( .A(n5829), .B(n5830), .Z(n5828) );
  XOR U5974 ( .A(n5831), .B(n5807), .Z(n5830) );
  XOR U5975 ( .A(n5821), .B(n5822), .Z(n5807) );
  XOR U5976 ( .A(n5832), .B(n5833), .Z(n5822) );
  ANDN U5977 ( .B(n5834), .A(n5835), .Z(n5832) );
  XOR U5978 ( .A(n5833), .B(n5836), .Z(n5834) );
  XOR U5979 ( .A(n5837), .B(n5838), .Z(n5821) );
  XOR U5980 ( .A(n5839), .B(n5840), .Z(n5838) );
  ANDN U5981 ( .B(n5841), .A(n5842), .Z(n5839) );
  XOR U5982 ( .A(n5843), .B(n5840), .Z(n5841) );
  IV U5983 ( .A(n5819), .Z(n5837) );
  XOR U5984 ( .A(n5844), .B(n5845), .Z(n5819) );
  ANDN U5985 ( .B(n5846), .A(n5847), .Z(n5844) );
  XOR U5986 ( .A(n5845), .B(n5848), .Z(n5846) );
  IV U5987 ( .A(n5827), .Z(n5831) );
  XOR U5988 ( .A(n5827), .B(n5809), .Z(n5829) );
  XOR U5989 ( .A(n5849), .B(n5850), .Z(n5809) );
  AND U5990 ( .A(n286), .B(n5851), .Z(n5849) );
  XOR U5991 ( .A(n5852), .B(n5850), .Z(n5851) );
  NANDN U5992 ( .A(n5811), .B(n5813), .Z(n5827) );
  XOR U5993 ( .A(n5853), .B(n5854), .Z(n5813) );
  AND U5994 ( .A(n286), .B(n5855), .Z(n5853) );
  XOR U5995 ( .A(n5854), .B(n5856), .Z(n5855) );
  XOR U5996 ( .A(n5857), .B(n5858), .Z(n286) );
  AND U5997 ( .A(n5859), .B(n5860), .Z(n5857) );
  XNOR U5998 ( .A(n5858), .B(n5824), .Z(n5860) );
  XNOR U5999 ( .A(n5861), .B(n5862), .Z(n5824) );
  ANDN U6000 ( .B(n5863), .A(n5864), .Z(n5861) );
  XOR U6001 ( .A(n5862), .B(n5865), .Z(n5863) );
  XOR U6002 ( .A(n5858), .B(n5826), .Z(n5859) );
  XOR U6003 ( .A(n5866), .B(n5867), .Z(n5826) );
  AND U6004 ( .A(n290), .B(n5868), .Z(n5866) );
  XOR U6005 ( .A(n5869), .B(n5867), .Z(n5868) );
  XNOR U6006 ( .A(n5870), .B(n5871), .Z(n5858) );
  NAND U6007 ( .A(n5872), .B(n5873), .Z(n5871) );
  XOR U6008 ( .A(n5874), .B(n5850), .Z(n5873) );
  XOR U6009 ( .A(n5864), .B(n5865), .Z(n5850) );
  XOR U6010 ( .A(n5875), .B(n5876), .Z(n5865) );
  ANDN U6011 ( .B(n5877), .A(n5878), .Z(n5875) );
  XOR U6012 ( .A(n5876), .B(n5879), .Z(n5877) );
  XOR U6013 ( .A(n5880), .B(n5881), .Z(n5864) );
  XOR U6014 ( .A(n5882), .B(n5883), .Z(n5881) );
  ANDN U6015 ( .B(n5884), .A(n5885), .Z(n5882) );
  XOR U6016 ( .A(n5886), .B(n5883), .Z(n5884) );
  IV U6017 ( .A(n5862), .Z(n5880) );
  XOR U6018 ( .A(n5887), .B(n5888), .Z(n5862) );
  ANDN U6019 ( .B(n5889), .A(n5890), .Z(n5887) );
  XOR U6020 ( .A(n5888), .B(n5891), .Z(n5889) );
  IV U6021 ( .A(n5870), .Z(n5874) );
  XOR U6022 ( .A(n5870), .B(n5852), .Z(n5872) );
  XOR U6023 ( .A(n5892), .B(n5893), .Z(n5852) );
  AND U6024 ( .A(n290), .B(n5894), .Z(n5892) );
  XOR U6025 ( .A(n5895), .B(n5893), .Z(n5894) );
  NANDN U6026 ( .A(n5854), .B(n5856), .Z(n5870) );
  XOR U6027 ( .A(n5896), .B(n5897), .Z(n5856) );
  AND U6028 ( .A(n290), .B(n5898), .Z(n5896) );
  XOR U6029 ( .A(n5897), .B(n5899), .Z(n5898) );
  XOR U6030 ( .A(n5900), .B(n5901), .Z(n290) );
  AND U6031 ( .A(n5902), .B(n5903), .Z(n5900) );
  XNOR U6032 ( .A(n5901), .B(n5867), .Z(n5903) );
  XNOR U6033 ( .A(n5904), .B(n5905), .Z(n5867) );
  ANDN U6034 ( .B(n5906), .A(n5907), .Z(n5904) );
  XOR U6035 ( .A(n5905), .B(n5908), .Z(n5906) );
  XOR U6036 ( .A(n5901), .B(n5869), .Z(n5902) );
  XOR U6037 ( .A(n5909), .B(n5910), .Z(n5869) );
  AND U6038 ( .A(n294), .B(n5911), .Z(n5909) );
  XOR U6039 ( .A(n5912), .B(n5910), .Z(n5911) );
  XNOR U6040 ( .A(n5913), .B(n5914), .Z(n5901) );
  NAND U6041 ( .A(n5915), .B(n5916), .Z(n5914) );
  XOR U6042 ( .A(n5917), .B(n5893), .Z(n5916) );
  XOR U6043 ( .A(n5907), .B(n5908), .Z(n5893) );
  XOR U6044 ( .A(n5918), .B(n5919), .Z(n5908) );
  ANDN U6045 ( .B(n5920), .A(n5921), .Z(n5918) );
  XOR U6046 ( .A(n5919), .B(n5922), .Z(n5920) );
  XOR U6047 ( .A(n5923), .B(n5924), .Z(n5907) );
  XOR U6048 ( .A(n5925), .B(n5926), .Z(n5924) );
  ANDN U6049 ( .B(n5927), .A(n5928), .Z(n5925) );
  XOR U6050 ( .A(n5929), .B(n5926), .Z(n5927) );
  IV U6051 ( .A(n5905), .Z(n5923) );
  XOR U6052 ( .A(n5930), .B(n5931), .Z(n5905) );
  ANDN U6053 ( .B(n5932), .A(n5933), .Z(n5930) );
  XOR U6054 ( .A(n5931), .B(n5934), .Z(n5932) );
  IV U6055 ( .A(n5913), .Z(n5917) );
  XOR U6056 ( .A(n5913), .B(n5895), .Z(n5915) );
  XOR U6057 ( .A(n5935), .B(n5936), .Z(n5895) );
  AND U6058 ( .A(n294), .B(n5937), .Z(n5935) );
  XOR U6059 ( .A(n5938), .B(n5936), .Z(n5937) );
  NANDN U6060 ( .A(n5897), .B(n5899), .Z(n5913) );
  XOR U6061 ( .A(n5939), .B(n5940), .Z(n5899) );
  AND U6062 ( .A(n294), .B(n5941), .Z(n5939) );
  XOR U6063 ( .A(n5940), .B(n5942), .Z(n5941) );
  XOR U6064 ( .A(n5943), .B(n5944), .Z(n294) );
  AND U6065 ( .A(n5945), .B(n5946), .Z(n5943) );
  XNOR U6066 ( .A(n5944), .B(n5910), .Z(n5946) );
  XNOR U6067 ( .A(n5947), .B(n5948), .Z(n5910) );
  ANDN U6068 ( .B(n5949), .A(n5950), .Z(n5947) );
  XOR U6069 ( .A(n5948), .B(n5951), .Z(n5949) );
  XOR U6070 ( .A(n5944), .B(n5912), .Z(n5945) );
  XOR U6071 ( .A(n5952), .B(n5953), .Z(n5912) );
  AND U6072 ( .A(n298), .B(n5954), .Z(n5952) );
  XOR U6073 ( .A(n5955), .B(n5953), .Z(n5954) );
  XNOR U6074 ( .A(n5956), .B(n5957), .Z(n5944) );
  NAND U6075 ( .A(n5958), .B(n5959), .Z(n5957) );
  XOR U6076 ( .A(n5960), .B(n5936), .Z(n5959) );
  XOR U6077 ( .A(n5950), .B(n5951), .Z(n5936) );
  XOR U6078 ( .A(n5961), .B(n5962), .Z(n5951) );
  ANDN U6079 ( .B(n5963), .A(n5964), .Z(n5961) );
  XOR U6080 ( .A(n5962), .B(n5965), .Z(n5963) );
  XOR U6081 ( .A(n5966), .B(n5967), .Z(n5950) );
  XOR U6082 ( .A(n5968), .B(n5969), .Z(n5967) );
  ANDN U6083 ( .B(n5970), .A(n5971), .Z(n5968) );
  XOR U6084 ( .A(n5972), .B(n5969), .Z(n5970) );
  IV U6085 ( .A(n5948), .Z(n5966) );
  XOR U6086 ( .A(n5973), .B(n5974), .Z(n5948) );
  ANDN U6087 ( .B(n5975), .A(n5976), .Z(n5973) );
  XOR U6088 ( .A(n5974), .B(n5977), .Z(n5975) );
  IV U6089 ( .A(n5956), .Z(n5960) );
  XOR U6090 ( .A(n5956), .B(n5938), .Z(n5958) );
  XOR U6091 ( .A(n5978), .B(n5979), .Z(n5938) );
  AND U6092 ( .A(n298), .B(n5980), .Z(n5978) );
  XOR U6093 ( .A(n5981), .B(n5979), .Z(n5980) );
  NANDN U6094 ( .A(n5940), .B(n5942), .Z(n5956) );
  XOR U6095 ( .A(n5982), .B(n5983), .Z(n5942) );
  AND U6096 ( .A(n298), .B(n5984), .Z(n5982) );
  XOR U6097 ( .A(n5983), .B(n5985), .Z(n5984) );
  XOR U6098 ( .A(n5986), .B(n5987), .Z(n298) );
  AND U6099 ( .A(n5988), .B(n5989), .Z(n5986) );
  XNOR U6100 ( .A(n5987), .B(n5953), .Z(n5989) );
  XNOR U6101 ( .A(n5990), .B(n5991), .Z(n5953) );
  ANDN U6102 ( .B(n5992), .A(n5993), .Z(n5990) );
  XOR U6103 ( .A(n5991), .B(n5994), .Z(n5992) );
  XOR U6104 ( .A(n5987), .B(n5955), .Z(n5988) );
  XOR U6105 ( .A(n5995), .B(n5996), .Z(n5955) );
  AND U6106 ( .A(n302), .B(n5997), .Z(n5995) );
  XOR U6107 ( .A(n5998), .B(n5996), .Z(n5997) );
  XNOR U6108 ( .A(n5999), .B(n6000), .Z(n5987) );
  NAND U6109 ( .A(n6001), .B(n6002), .Z(n6000) );
  XOR U6110 ( .A(n6003), .B(n5979), .Z(n6002) );
  XOR U6111 ( .A(n5993), .B(n5994), .Z(n5979) );
  XOR U6112 ( .A(n6004), .B(n6005), .Z(n5994) );
  ANDN U6113 ( .B(n6006), .A(n6007), .Z(n6004) );
  XOR U6114 ( .A(n6005), .B(n6008), .Z(n6006) );
  XOR U6115 ( .A(n6009), .B(n6010), .Z(n5993) );
  XOR U6116 ( .A(n6011), .B(n6012), .Z(n6010) );
  ANDN U6117 ( .B(n6013), .A(n6014), .Z(n6011) );
  XOR U6118 ( .A(n6015), .B(n6012), .Z(n6013) );
  IV U6119 ( .A(n5991), .Z(n6009) );
  XOR U6120 ( .A(n6016), .B(n6017), .Z(n5991) );
  ANDN U6121 ( .B(n6018), .A(n6019), .Z(n6016) );
  XOR U6122 ( .A(n6017), .B(n6020), .Z(n6018) );
  IV U6123 ( .A(n5999), .Z(n6003) );
  XOR U6124 ( .A(n5999), .B(n5981), .Z(n6001) );
  XOR U6125 ( .A(n6021), .B(n6022), .Z(n5981) );
  AND U6126 ( .A(n302), .B(n6023), .Z(n6021) );
  XOR U6127 ( .A(n6024), .B(n6022), .Z(n6023) );
  NANDN U6128 ( .A(n5983), .B(n5985), .Z(n5999) );
  XOR U6129 ( .A(n6025), .B(n6026), .Z(n5985) );
  AND U6130 ( .A(n302), .B(n6027), .Z(n6025) );
  XOR U6131 ( .A(n6026), .B(n6028), .Z(n6027) );
  XOR U6132 ( .A(n6029), .B(n6030), .Z(n302) );
  AND U6133 ( .A(n6031), .B(n6032), .Z(n6029) );
  XNOR U6134 ( .A(n6030), .B(n5996), .Z(n6032) );
  XNOR U6135 ( .A(n6033), .B(n6034), .Z(n5996) );
  ANDN U6136 ( .B(n6035), .A(n6036), .Z(n6033) );
  XOR U6137 ( .A(n6034), .B(n6037), .Z(n6035) );
  XOR U6138 ( .A(n6030), .B(n5998), .Z(n6031) );
  XOR U6139 ( .A(n6038), .B(n6039), .Z(n5998) );
  AND U6140 ( .A(n306), .B(n6040), .Z(n6038) );
  XOR U6141 ( .A(n6041), .B(n6039), .Z(n6040) );
  XNOR U6142 ( .A(n6042), .B(n6043), .Z(n6030) );
  NAND U6143 ( .A(n6044), .B(n6045), .Z(n6043) );
  XOR U6144 ( .A(n6046), .B(n6022), .Z(n6045) );
  XOR U6145 ( .A(n6036), .B(n6037), .Z(n6022) );
  XOR U6146 ( .A(n6047), .B(n6048), .Z(n6037) );
  ANDN U6147 ( .B(n6049), .A(n6050), .Z(n6047) );
  XOR U6148 ( .A(n6048), .B(n6051), .Z(n6049) );
  XOR U6149 ( .A(n6052), .B(n6053), .Z(n6036) );
  XOR U6150 ( .A(n6054), .B(n6055), .Z(n6053) );
  ANDN U6151 ( .B(n6056), .A(n6057), .Z(n6054) );
  XOR U6152 ( .A(n6058), .B(n6055), .Z(n6056) );
  IV U6153 ( .A(n6034), .Z(n6052) );
  XOR U6154 ( .A(n6059), .B(n6060), .Z(n6034) );
  ANDN U6155 ( .B(n6061), .A(n6062), .Z(n6059) );
  XOR U6156 ( .A(n6060), .B(n6063), .Z(n6061) );
  IV U6157 ( .A(n6042), .Z(n6046) );
  XOR U6158 ( .A(n6042), .B(n6024), .Z(n6044) );
  XOR U6159 ( .A(n6064), .B(n6065), .Z(n6024) );
  AND U6160 ( .A(n306), .B(n6066), .Z(n6064) );
  XOR U6161 ( .A(n6067), .B(n6065), .Z(n6066) );
  NANDN U6162 ( .A(n6026), .B(n6028), .Z(n6042) );
  XOR U6163 ( .A(n6068), .B(n6069), .Z(n6028) );
  AND U6164 ( .A(n306), .B(n6070), .Z(n6068) );
  XOR U6165 ( .A(n6069), .B(n6071), .Z(n6070) );
  XOR U6166 ( .A(n6072), .B(n6073), .Z(n306) );
  AND U6167 ( .A(n6074), .B(n6075), .Z(n6072) );
  XNOR U6168 ( .A(n6073), .B(n6039), .Z(n6075) );
  XNOR U6169 ( .A(n6076), .B(n6077), .Z(n6039) );
  ANDN U6170 ( .B(n6078), .A(n6079), .Z(n6076) );
  XOR U6171 ( .A(n6077), .B(n6080), .Z(n6078) );
  XOR U6172 ( .A(n6073), .B(n6041), .Z(n6074) );
  XOR U6173 ( .A(n6081), .B(n6082), .Z(n6041) );
  AND U6174 ( .A(n310), .B(n6083), .Z(n6081) );
  XOR U6175 ( .A(n6084), .B(n6082), .Z(n6083) );
  XNOR U6176 ( .A(n6085), .B(n6086), .Z(n6073) );
  NAND U6177 ( .A(n6087), .B(n6088), .Z(n6086) );
  XOR U6178 ( .A(n6089), .B(n6065), .Z(n6088) );
  XOR U6179 ( .A(n6079), .B(n6080), .Z(n6065) );
  XOR U6180 ( .A(n6090), .B(n6091), .Z(n6080) );
  ANDN U6181 ( .B(n6092), .A(n6093), .Z(n6090) );
  XOR U6182 ( .A(n6091), .B(n6094), .Z(n6092) );
  XOR U6183 ( .A(n6095), .B(n6096), .Z(n6079) );
  XOR U6184 ( .A(n6097), .B(n6098), .Z(n6096) );
  ANDN U6185 ( .B(n6099), .A(n6100), .Z(n6097) );
  XOR U6186 ( .A(n6101), .B(n6098), .Z(n6099) );
  IV U6187 ( .A(n6077), .Z(n6095) );
  XOR U6188 ( .A(n6102), .B(n6103), .Z(n6077) );
  ANDN U6189 ( .B(n6104), .A(n6105), .Z(n6102) );
  XOR U6190 ( .A(n6103), .B(n6106), .Z(n6104) );
  IV U6191 ( .A(n6085), .Z(n6089) );
  XOR U6192 ( .A(n6085), .B(n6067), .Z(n6087) );
  XOR U6193 ( .A(n6107), .B(n6108), .Z(n6067) );
  AND U6194 ( .A(n310), .B(n6109), .Z(n6107) );
  XOR U6195 ( .A(n6110), .B(n6108), .Z(n6109) );
  NANDN U6196 ( .A(n6069), .B(n6071), .Z(n6085) );
  XOR U6197 ( .A(n6111), .B(n6112), .Z(n6071) );
  AND U6198 ( .A(n310), .B(n6113), .Z(n6111) );
  XOR U6199 ( .A(n6112), .B(n6114), .Z(n6113) );
  XOR U6200 ( .A(n6115), .B(n6116), .Z(n310) );
  AND U6201 ( .A(n6117), .B(n6118), .Z(n6115) );
  XNOR U6202 ( .A(n6116), .B(n6082), .Z(n6118) );
  XNOR U6203 ( .A(n6119), .B(n6120), .Z(n6082) );
  ANDN U6204 ( .B(n6121), .A(n6122), .Z(n6119) );
  XOR U6205 ( .A(n6120), .B(n6123), .Z(n6121) );
  XOR U6206 ( .A(n6116), .B(n6084), .Z(n6117) );
  XOR U6207 ( .A(n6124), .B(n6125), .Z(n6084) );
  AND U6208 ( .A(n314), .B(n6126), .Z(n6124) );
  XOR U6209 ( .A(n6127), .B(n6125), .Z(n6126) );
  XNOR U6210 ( .A(n6128), .B(n6129), .Z(n6116) );
  NAND U6211 ( .A(n6130), .B(n6131), .Z(n6129) );
  XOR U6212 ( .A(n6132), .B(n6108), .Z(n6131) );
  XOR U6213 ( .A(n6122), .B(n6123), .Z(n6108) );
  XOR U6214 ( .A(n6133), .B(n6134), .Z(n6123) );
  ANDN U6215 ( .B(n6135), .A(n6136), .Z(n6133) );
  XOR U6216 ( .A(n6134), .B(n6137), .Z(n6135) );
  XOR U6217 ( .A(n6138), .B(n6139), .Z(n6122) );
  XOR U6218 ( .A(n6140), .B(n6141), .Z(n6139) );
  ANDN U6219 ( .B(n6142), .A(n6143), .Z(n6140) );
  XOR U6220 ( .A(n6144), .B(n6141), .Z(n6142) );
  IV U6221 ( .A(n6120), .Z(n6138) );
  XOR U6222 ( .A(n6145), .B(n6146), .Z(n6120) );
  ANDN U6223 ( .B(n6147), .A(n6148), .Z(n6145) );
  XOR U6224 ( .A(n6146), .B(n6149), .Z(n6147) );
  IV U6225 ( .A(n6128), .Z(n6132) );
  XOR U6226 ( .A(n6128), .B(n6110), .Z(n6130) );
  XOR U6227 ( .A(n6150), .B(n6151), .Z(n6110) );
  AND U6228 ( .A(n314), .B(n6152), .Z(n6150) );
  XOR U6229 ( .A(n6153), .B(n6151), .Z(n6152) );
  NANDN U6230 ( .A(n6112), .B(n6114), .Z(n6128) );
  XOR U6231 ( .A(n6154), .B(n6155), .Z(n6114) );
  AND U6232 ( .A(n314), .B(n6156), .Z(n6154) );
  XOR U6233 ( .A(n6155), .B(n6157), .Z(n6156) );
  XOR U6234 ( .A(n6158), .B(n6159), .Z(n314) );
  AND U6235 ( .A(n6160), .B(n6161), .Z(n6158) );
  XNOR U6236 ( .A(n6159), .B(n6125), .Z(n6161) );
  XNOR U6237 ( .A(n6162), .B(n6163), .Z(n6125) );
  ANDN U6238 ( .B(n6164), .A(n6165), .Z(n6162) );
  XOR U6239 ( .A(n6163), .B(n6166), .Z(n6164) );
  XOR U6240 ( .A(n6159), .B(n6127), .Z(n6160) );
  XOR U6241 ( .A(n6167), .B(n6168), .Z(n6127) );
  AND U6242 ( .A(n318), .B(n6169), .Z(n6167) );
  XOR U6243 ( .A(n6170), .B(n6168), .Z(n6169) );
  XNOR U6244 ( .A(n6171), .B(n6172), .Z(n6159) );
  NAND U6245 ( .A(n6173), .B(n6174), .Z(n6172) );
  XOR U6246 ( .A(n6175), .B(n6151), .Z(n6174) );
  XOR U6247 ( .A(n6165), .B(n6166), .Z(n6151) );
  XOR U6248 ( .A(n6176), .B(n6177), .Z(n6166) );
  ANDN U6249 ( .B(n6178), .A(n6179), .Z(n6176) );
  XOR U6250 ( .A(n6177), .B(n6180), .Z(n6178) );
  XOR U6251 ( .A(n6181), .B(n6182), .Z(n6165) );
  XOR U6252 ( .A(n6183), .B(n6184), .Z(n6182) );
  ANDN U6253 ( .B(n6185), .A(n6186), .Z(n6183) );
  XOR U6254 ( .A(n6187), .B(n6184), .Z(n6185) );
  IV U6255 ( .A(n6163), .Z(n6181) );
  XOR U6256 ( .A(n6188), .B(n6189), .Z(n6163) );
  ANDN U6257 ( .B(n6190), .A(n6191), .Z(n6188) );
  XOR U6258 ( .A(n6189), .B(n6192), .Z(n6190) );
  IV U6259 ( .A(n6171), .Z(n6175) );
  XOR U6260 ( .A(n6171), .B(n6153), .Z(n6173) );
  XOR U6261 ( .A(n6193), .B(n6194), .Z(n6153) );
  AND U6262 ( .A(n318), .B(n6195), .Z(n6193) );
  XOR U6263 ( .A(n6196), .B(n6194), .Z(n6195) );
  NANDN U6264 ( .A(n6155), .B(n6157), .Z(n6171) );
  XOR U6265 ( .A(n6197), .B(n6198), .Z(n6157) );
  AND U6266 ( .A(n318), .B(n6199), .Z(n6197) );
  XOR U6267 ( .A(n6198), .B(n6200), .Z(n6199) );
  XOR U6268 ( .A(n6201), .B(n6202), .Z(n318) );
  AND U6269 ( .A(n6203), .B(n6204), .Z(n6201) );
  XNOR U6270 ( .A(n6202), .B(n6168), .Z(n6204) );
  XNOR U6271 ( .A(n6205), .B(n6206), .Z(n6168) );
  ANDN U6272 ( .B(n6207), .A(n6208), .Z(n6205) );
  XOR U6273 ( .A(n6206), .B(n6209), .Z(n6207) );
  XOR U6274 ( .A(n6202), .B(n6170), .Z(n6203) );
  XOR U6275 ( .A(n6210), .B(n6211), .Z(n6170) );
  AND U6276 ( .A(n322), .B(n6212), .Z(n6210) );
  XOR U6277 ( .A(n6213), .B(n6211), .Z(n6212) );
  XNOR U6278 ( .A(n6214), .B(n6215), .Z(n6202) );
  NAND U6279 ( .A(n6216), .B(n6217), .Z(n6215) );
  XOR U6280 ( .A(n6218), .B(n6194), .Z(n6217) );
  XOR U6281 ( .A(n6208), .B(n6209), .Z(n6194) );
  XOR U6282 ( .A(n6219), .B(n6220), .Z(n6209) );
  ANDN U6283 ( .B(n6221), .A(n6222), .Z(n6219) );
  XOR U6284 ( .A(n6220), .B(n6223), .Z(n6221) );
  XOR U6285 ( .A(n6224), .B(n6225), .Z(n6208) );
  XOR U6286 ( .A(n6226), .B(n6227), .Z(n6225) );
  ANDN U6287 ( .B(n6228), .A(n6229), .Z(n6226) );
  XOR U6288 ( .A(n6230), .B(n6227), .Z(n6228) );
  IV U6289 ( .A(n6206), .Z(n6224) );
  XOR U6290 ( .A(n6231), .B(n6232), .Z(n6206) );
  ANDN U6291 ( .B(n6233), .A(n6234), .Z(n6231) );
  XOR U6292 ( .A(n6232), .B(n6235), .Z(n6233) );
  IV U6293 ( .A(n6214), .Z(n6218) );
  XOR U6294 ( .A(n6214), .B(n6196), .Z(n6216) );
  XOR U6295 ( .A(n6236), .B(n6237), .Z(n6196) );
  AND U6296 ( .A(n322), .B(n6238), .Z(n6236) );
  XOR U6297 ( .A(n6239), .B(n6237), .Z(n6238) );
  NANDN U6298 ( .A(n6198), .B(n6200), .Z(n6214) );
  XOR U6299 ( .A(n6240), .B(n6241), .Z(n6200) );
  AND U6300 ( .A(n322), .B(n6242), .Z(n6240) );
  XOR U6301 ( .A(n6241), .B(n6243), .Z(n6242) );
  XOR U6302 ( .A(n6244), .B(n6245), .Z(n322) );
  AND U6303 ( .A(n6246), .B(n6247), .Z(n6244) );
  XNOR U6304 ( .A(n6245), .B(n6211), .Z(n6247) );
  XNOR U6305 ( .A(n6248), .B(n6249), .Z(n6211) );
  ANDN U6306 ( .B(n6250), .A(n6251), .Z(n6248) );
  XOR U6307 ( .A(n6249), .B(n6252), .Z(n6250) );
  XOR U6308 ( .A(n6245), .B(n6213), .Z(n6246) );
  XOR U6309 ( .A(n6253), .B(n6254), .Z(n6213) );
  AND U6310 ( .A(n326), .B(n6255), .Z(n6253) );
  XOR U6311 ( .A(n6256), .B(n6254), .Z(n6255) );
  XNOR U6312 ( .A(n6257), .B(n6258), .Z(n6245) );
  NAND U6313 ( .A(n6259), .B(n6260), .Z(n6258) );
  XOR U6314 ( .A(n6261), .B(n6237), .Z(n6260) );
  XOR U6315 ( .A(n6251), .B(n6252), .Z(n6237) );
  XOR U6316 ( .A(n6262), .B(n6263), .Z(n6252) );
  ANDN U6317 ( .B(n6264), .A(n6265), .Z(n6262) );
  XOR U6318 ( .A(n6263), .B(n6266), .Z(n6264) );
  XOR U6319 ( .A(n6267), .B(n6268), .Z(n6251) );
  XOR U6320 ( .A(n6269), .B(n6270), .Z(n6268) );
  ANDN U6321 ( .B(n6271), .A(n6272), .Z(n6269) );
  XOR U6322 ( .A(n6273), .B(n6270), .Z(n6271) );
  IV U6323 ( .A(n6249), .Z(n6267) );
  XOR U6324 ( .A(n6274), .B(n6275), .Z(n6249) );
  ANDN U6325 ( .B(n6276), .A(n6277), .Z(n6274) );
  XOR U6326 ( .A(n6275), .B(n6278), .Z(n6276) );
  IV U6327 ( .A(n6257), .Z(n6261) );
  XOR U6328 ( .A(n6257), .B(n6239), .Z(n6259) );
  XOR U6329 ( .A(n6279), .B(n6280), .Z(n6239) );
  AND U6330 ( .A(n326), .B(n6281), .Z(n6279) );
  XOR U6331 ( .A(n6282), .B(n6280), .Z(n6281) );
  NANDN U6332 ( .A(n6241), .B(n6243), .Z(n6257) );
  XOR U6333 ( .A(n6283), .B(n6284), .Z(n6243) );
  AND U6334 ( .A(n326), .B(n6285), .Z(n6283) );
  XOR U6335 ( .A(n6284), .B(n6286), .Z(n6285) );
  XOR U6336 ( .A(n6287), .B(n6288), .Z(n326) );
  AND U6337 ( .A(n6289), .B(n6290), .Z(n6287) );
  XNOR U6338 ( .A(n6288), .B(n6254), .Z(n6290) );
  XNOR U6339 ( .A(n6291), .B(n6292), .Z(n6254) );
  ANDN U6340 ( .B(n6293), .A(n6294), .Z(n6291) );
  XOR U6341 ( .A(n6292), .B(n6295), .Z(n6293) );
  XOR U6342 ( .A(n6288), .B(n6256), .Z(n6289) );
  XOR U6343 ( .A(n6296), .B(n6297), .Z(n6256) );
  AND U6344 ( .A(n330), .B(n6298), .Z(n6296) );
  XOR U6345 ( .A(n6299), .B(n6297), .Z(n6298) );
  XNOR U6346 ( .A(n6300), .B(n6301), .Z(n6288) );
  NAND U6347 ( .A(n6302), .B(n6303), .Z(n6301) );
  XOR U6348 ( .A(n6304), .B(n6280), .Z(n6303) );
  XOR U6349 ( .A(n6294), .B(n6295), .Z(n6280) );
  XOR U6350 ( .A(n6305), .B(n6306), .Z(n6295) );
  ANDN U6351 ( .B(n6307), .A(n6308), .Z(n6305) );
  XOR U6352 ( .A(n6306), .B(n6309), .Z(n6307) );
  XOR U6353 ( .A(n6310), .B(n6311), .Z(n6294) );
  XOR U6354 ( .A(n6312), .B(n6313), .Z(n6311) );
  ANDN U6355 ( .B(n6314), .A(n6315), .Z(n6312) );
  XOR U6356 ( .A(n6316), .B(n6313), .Z(n6314) );
  IV U6357 ( .A(n6292), .Z(n6310) );
  XOR U6358 ( .A(n6317), .B(n6318), .Z(n6292) );
  ANDN U6359 ( .B(n6319), .A(n6320), .Z(n6317) );
  XOR U6360 ( .A(n6318), .B(n6321), .Z(n6319) );
  IV U6361 ( .A(n6300), .Z(n6304) );
  XOR U6362 ( .A(n6300), .B(n6282), .Z(n6302) );
  XOR U6363 ( .A(n6322), .B(n6323), .Z(n6282) );
  AND U6364 ( .A(n330), .B(n6324), .Z(n6322) );
  XOR U6365 ( .A(n6325), .B(n6323), .Z(n6324) );
  NANDN U6366 ( .A(n6284), .B(n6286), .Z(n6300) );
  XOR U6367 ( .A(n6326), .B(n6327), .Z(n6286) );
  AND U6368 ( .A(n330), .B(n6328), .Z(n6326) );
  XOR U6369 ( .A(n6327), .B(n6329), .Z(n6328) );
  XOR U6370 ( .A(n6330), .B(n6331), .Z(n330) );
  AND U6371 ( .A(n6332), .B(n6333), .Z(n6330) );
  XNOR U6372 ( .A(n6331), .B(n6297), .Z(n6333) );
  XNOR U6373 ( .A(n6334), .B(n6335), .Z(n6297) );
  ANDN U6374 ( .B(n6336), .A(n6337), .Z(n6334) );
  XOR U6375 ( .A(n6335), .B(n6338), .Z(n6336) );
  XOR U6376 ( .A(n6331), .B(n6299), .Z(n6332) );
  XOR U6377 ( .A(n6339), .B(n6340), .Z(n6299) );
  AND U6378 ( .A(n334), .B(n6341), .Z(n6339) );
  XOR U6379 ( .A(n6342), .B(n6340), .Z(n6341) );
  XNOR U6380 ( .A(n6343), .B(n6344), .Z(n6331) );
  NAND U6381 ( .A(n6345), .B(n6346), .Z(n6344) );
  XOR U6382 ( .A(n6347), .B(n6323), .Z(n6346) );
  XOR U6383 ( .A(n6337), .B(n6338), .Z(n6323) );
  XOR U6384 ( .A(n6348), .B(n6349), .Z(n6338) );
  ANDN U6385 ( .B(n6350), .A(n6351), .Z(n6348) );
  XOR U6386 ( .A(n6349), .B(n6352), .Z(n6350) );
  XOR U6387 ( .A(n6353), .B(n6354), .Z(n6337) );
  XOR U6388 ( .A(n6355), .B(n6356), .Z(n6354) );
  ANDN U6389 ( .B(n6357), .A(n6358), .Z(n6355) );
  XOR U6390 ( .A(n6359), .B(n6356), .Z(n6357) );
  IV U6391 ( .A(n6335), .Z(n6353) );
  XOR U6392 ( .A(n6360), .B(n6361), .Z(n6335) );
  ANDN U6393 ( .B(n6362), .A(n6363), .Z(n6360) );
  XOR U6394 ( .A(n6361), .B(n6364), .Z(n6362) );
  IV U6395 ( .A(n6343), .Z(n6347) );
  XOR U6396 ( .A(n6343), .B(n6325), .Z(n6345) );
  XOR U6397 ( .A(n6365), .B(n6366), .Z(n6325) );
  AND U6398 ( .A(n334), .B(n6367), .Z(n6365) );
  XOR U6399 ( .A(n6368), .B(n6366), .Z(n6367) );
  NANDN U6400 ( .A(n6327), .B(n6329), .Z(n6343) );
  XOR U6401 ( .A(n6369), .B(n6370), .Z(n6329) );
  AND U6402 ( .A(n334), .B(n6371), .Z(n6369) );
  XOR U6403 ( .A(n6370), .B(n6372), .Z(n6371) );
  XOR U6404 ( .A(n6373), .B(n6374), .Z(n334) );
  AND U6405 ( .A(n6375), .B(n6376), .Z(n6373) );
  XNOR U6406 ( .A(n6374), .B(n6340), .Z(n6376) );
  XNOR U6407 ( .A(n6377), .B(n6378), .Z(n6340) );
  ANDN U6408 ( .B(n6379), .A(n6380), .Z(n6377) );
  XOR U6409 ( .A(n6378), .B(n6381), .Z(n6379) );
  XOR U6410 ( .A(n6374), .B(n6342), .Z(n6375) );
  XOR U6411 ( .A(n6382), .B(n6383), .Z(n6342) );
  AND U6412 ( .A(n338), .B(n6384), .Z(n6382) );
  XOR U6413 ( .A(n6385), .B(n6383), .Z(n6384) );
  XNOR U6414 ( .A(n6386), .B(n6387), .Z(n6374) );
  NAND U6415 ( .A(n6388), .B(n6389), .Z(n6387) );
  XOR U6416 ( .A(n6390), .B(n6366), .Z(n6389) );
  XOR U6417 ( .A(n6380), .B(n6381), .Z(n6366) );
  XOR U6418 ( .A(n6391), .B(n6392), .Z(n6381) );
  ANDN U6419 ( .B(n6393), .A(n6394), .Z(n6391) );
  XOR U6420 ( .A(n6392), .B(n6395), .Z(n6393) );
  XOR U6421 ( .A(n6396), .B(n6397), .Z(n6380) );
  XOR U6422 ( .A(n6398), .B(n6399), .Z(n6397) );
  ANDN U6423 ( .B(n6400), .A(n6401), .Z(n6398) );
  XOR U6424 ( .A(n6402), .B(n6399), .Z(n6400) );
  IV U6425 ( .A(n6378), .Z(n6396) );
  XOR U6426 ( .A(n6403), .B(n6404), .Z(n6378) );
  ANDN U6427 ( .B(n6405), .A(n6406), .Z(n6403) );
  XOR U6428 ( .A(n6404), .B(n6407), .Z(n6405) );
  IV U6429 ( .A(n6386), .Z(n6390) );
  XOR U6430 ( .A(n6386), .B(n6368), .Z(n6388) );
  XOR U6431 ( .A(n6408), .B(n6409), .Z(n6368) );
  AND U6432 ( .A(n338), .B(n6410), .Z(n6408) );
  XOR U6433 ( .A(n6411), .B(n6409), .Z(n6410) );
  NANDN U6434 ( .A(n6370), .B(n6372), .Z(n6386) );
  XOR U6435 ( .A(n6412), .B(n6413), .Z(n6372) );
  AND U6436 ( .A(n338), .B(n6414), .Z(n6412) );
  XOR U6437 ( .A(n6413), .B(n6415), .Z(n6414) );
  XOR U6438 ( .A(n6416), .B(n6417), .Z(n338) );
  AND U6439 ( .A(n6418), .B(n6419), .Z(n6416) );
  XNOR U6440 ( .A(n6417), .B(n6383), .Z(n6419) );
  XNOR U6441 ( .A(n6420), .B(n6421), .Z(n6383) );
  ANDN U6442 ( .B(n6422), .A(n6423), .Z(n6420) );
  XOR U6443 ( .A(n6421), .B(n6424), .Z(n6422) );
  XOR U6444 ( .A(n6417), .B(n6385), .Z(n6418) );
  XOR U6445 ( .A(n6425), .B(n6426), .Z(n6385) );
  AND U6446 ( .A(n342), .B(n6427), .Z(n6425) );
  XOR U6447 ( .A(n6428), .B(n6426), .Z(n6427) );
  XNOR U6448 ( .A(n6429), .B(n6430), .Z(n6417) );
  NAND U6449 ( .A(n6431), .B(n6432), .Z(n6430) );
  XOR U6450 ( .A(n6433), .B(n6409), .Z(n6432) );
  XOR U6451 ( .A(n6423), .B(n6424), .Z(n6409) );
  XOR U6452 ( .A(n6434), .B(n6435), .Z(n6424) );
  ANDN U6453 ( .B(n6436), .A(n6437), .Z(n6434) );
  XOR U6454 ( .A(n6435), .B(n6438), .Z(n6436) );
  XOR U6455 ( .A(n6439), .B(n6440), .Z(n6423) );
  XOR U6456 ( .A(n6441), .B(n6442), .Z(n6440) );
  ANDN U6457 ( .B(n6443), .A(n6444), .Z(n6441) );
  XOR U6458 ( .A(n6445), .B(n6442), .Z(n6443) );
  IV U6459 ( .A(n6421), .Z(n6439) );
  XOR U6460 ( .A(n6446), .B(n6447), .Z(n6421) );
  ANDN U6461 ( .B(n6448), .A(n6449), .Z(n6446) );
  XOR U6462 ( .A(n6447), .B(n6450), .Z(n6448) );
  IV U6463 ( .A(n6429), .Z(n6433) );
  XOR U6464 ( .A(n6429), .B(n6411), .Z(n6431) );
  XOR U6465 ( .A(n6451), .B(n6452), .Z(n6411) );
  AND U6466 ( .A(n342), .B(n6453), .Z(n6451) );
  XOR U6467 ( .A(n6454), .B(n6452), .Z(n6453) );
  NANDN U6468 ( .A(n6413), .B(n6415), .Z(n6429) );
  XOR U6469 ( .A(n6455), .B(n6456), .Z(n6415) );
  AND U6470 ( .A(n342), .B(n6457), .Z(n6455) );
  XOR U6471 ( .A(n6456), .B(n6458), .Z(n6457) );
  XOR U6472 ( .A(n6459), .B(n6460), .Z(n342) );
  AND U6473 ( .A(n6461), .B(n6462), .Z(n6459) );
  XNOR U6474 ( .A(n6460), .B(n6426), .Z(n6462) );
  XNOR U6475 ( .A(n6463), .B(n6464), .Z(n6426) );
  ANDN U6476 ( .B(n6465), .A(n6466), .Z(n6463) );
  XOR U6477 ( .A(n6464), .B(n6467), .Z(n6465) );
  XOR U6478 ( .A(n6460), .B(n6428), .Z(n6461) );
  XOR U6479 ( .A(n6468), .B(n6469), .Z(n6428) );
  AND U6480 ( .A(n346), .B(n6470), .Z(n6468) );
  XOR U6481 ( .A(n6471), .B(n6469), .Z(n6470) );
  XNOR U6482 ( .A(n6472), .B(n6473), .Z(n6460) );
  NAND U6483 ( .A(n6474), .B(n6475), .Z(n6473) );
  XOR U6484 ( .A(n6476), .B(n6452), .Z(n6475) );
  XOR U6485 ( .A(n6466), .B(n6467), .Z(n6452) );
  XOR U6486 ( .A(n6477), .B(n6478), .Z(n6467) );
  ANDN U6487 ( .B(n6479), .A(n6480), .Z(n6477) );
  XOR U6488 ( .A(n6478), .B(n6481), .Z(n6479) );
  XOR U6489 ( .A(n6482), .B(n6483), .Z(n6466) );
  XOR U6490 ( .A(n6484), .B(n6485), .Z(n6483) );
  ANDN U6491 ( .B(n6486), .A(n6487), .Z(n6484) );
  XOR U6492 ( .A(n6488), .B(n6485), .Z(n6486) );
  IV U6493 ( .A(n6464), .Z(n6482) );
  XOR U6494 ( .A(n6489), .B(n6490), .Z(n6464) );
  ANDN U6495 ( .B(n6491), .A(n6492), .Z(n6489) );
  XOR U6496 ( .A(n6490), .B(n6493), .Z(n6491) );
  IV U6497 ( .A(n6472), .Z(n6476) );
  XOR U6498 ( .A(n6472), .B(n6454), .Z(n6474) );
  XOR U6499 ( .A(n6494), .B(n6495), .Z(n6454) );
  AND U6500 ( .A(n346), .B(n6496), .Z(n6494) );
  XOR U6501 ( .A(n6497), .B(n6495), .Z(n6496) );
  NANDN U6502 ( .A(n6456), .B(n6458), .Z(n6472) );
  XOR U6503 ( .A(n6498), .B(n6499), .Z(n6458) );
  AND U6504 ( .A(n346), .B(n6500), .Z(n6498) );
  XOR U6505 ( .A(n6499), .B(n6501), .Z(n6500) );
  XOR U6506 ( .A(n6502), .B(n6503), .Z(n346) );
  AND U6507 ( .A(n6504), .B(n6505), .Z(n6502) );
  XNOR U6508 ( .A(n6503), .B(n6469), .Z(n6505) );
  XNOR U6509 ( .A(n6506), .B(n6507), .Z(n6469) );
  ANDN U6510 ( .B(n6508), .A(n6509), .Z(n6506) );
  XOR U6511 ( .A(n6507), .B(n6510), .Z(n6508) );
  XOR U6512 ( .A(n6503), .B(n6471), .Z(n6504) );
  XOR U6513 ( .A(n6511), .B(n6512), .Z(n6471) );
  AND U6514 ( .A(n350), .B(n6513), .Z(n6511) );
  XOR U6515 ( .A(n6514), .B(n6512), .Z(n6513) );
  XNOR U6516 ( .A(n6515), .B(n6516), .Z(n6503) );
  NAND U6517 ( .A(n6517), .B(n6518), .Z(n6516) );
  XOR U6518 ( .A(n6519), .B(n6495), .Z(n6518) );
  XOR U6519 ( .A(n6509), .B(n6510), .Z(n6495) );
  XOR U6520 ( .A(n6520), .B(n6521), .Z(n6510) );
  ANDN U6521 ( .B(n6522), .A(n6523), .Z(n6520) );
  XOR U6522 ( .A(n6521), .B(n6524), .Z(n6522) );
  XOR U6523 ( .A(n6525), .B(n6526), .Z(n6509) );
  XOR U6524 ( .A(n6527), .B(n6528), .Z(n6526) );
  ANDN U6525 ( .B(n6529), .A(n6530), .Z(n6527) );
  XOR U6526 ( .A(n6531), .B(n6528), .Z(n6529) );
  IV U6527 ( .A(n6507), .Z(n6525) );
  XOR U6528 ( .A(n6532), .B(n6533), .Z(n6507) );
  ANDN U6529 ( .B(n6534), .A(n6535), .Z(n6532) );
  XOR U6530 ( .A(n6533), .B(n6536), .Z(n6534) );
  IV U6531 ( .A(n6515), .Z(n6519) );
  XOR U6532 ( .A(n6515), .B(n6497), .Z(n6517) );
  XOR U6533 ( .A(n6537), .B(n6538), .Z(n6497) );
  AND U6534 ( .A(n350), .B(n6539), .Z(n6537) );
  XOR U6535 ( .A(n6540), .B(n6538), .Z(n6539) );
  NANDN U6536 ( .A(n6499), .B(n6501), .Z(n6515) );
  XOR U6537 ( .A(n6541), .B(n6542), .Z(n6501) );
  AND U6538 ( .A(n350), .B(n6543), .Z(n6541) );
  XOR U6539 ( .A(n6542), .B(n6544), .Z(n6543) );
  XOR U6540 ( .A(n6545), .B(n6546), .Z(n350) );
  AND U6541 ( .A(n6547), .B(n6548), .Z(n6545) );
  XNOR U6542 ( .A(n6546), .B(n6512), .Z(n6548) );
  XNOR U6543 ( .A(n6549), .B(n6550), .Z(n6512) );
  ANDN U6544 ( .B(n6551), .A(n6552), .Z(n6549) );
  XOR U6545 ( .A(n6550), .B(n6553), .Z(n6551) );
  XOR U6546 ( .A(n6546), .B(n6514), .Z(n6547) );
  XOR U6547 ( .A(n6554), .B(n6555), .Z(n6514) );
  AND U6548 ( .A(n354), .B(n6556), .Z(n6554) );
  XOR U6549 ( .A(n6557), .B(n6555), .Z(n6556) );
  XNOR U6550 ( .A(n6558), .B(n6559), .Z(n6546) );
  NAND U6551 ( .A(n6560), .B(n6561), .Z(n6559) );
  XOR U6552 ( .A(n6562), .B(n6538), .Z(n6561) );
  XOR U6553 ( .A(n6552), .B(n6553), .Z(n6538) );
  XOR U6554 ( .A(n6563), .B(n6564), .Z(n6553) );
  ANDN U6555 ( .B(n6565), .A(n6566), .Z(n6563) );
  XOR U6556 ( .A(n6564), .B(n6567), .Z(n6565) );
  XOR U6557 ( .A(n6568), .B(n6569), .Z(n6552) );
  XOR U6558 ( .A(n6570), .B(n6571), .Z(n6569) );
  ANDN U6559 ( .B(n6572), .A(n6573), .Z(n6570) );
  XOR U6560 ( .A(n6574), .B(n6571), .Z(n6572) );
  IV U6561 ( .A(n6550), .Z(n6568) );
  XOR U6562 ( .A(n6575), .B(n6576), .Z(n6550) );
  ANDN U6563 ( .B(n6577), .A(n6578), .Z(n6575) );
  XOR U6564 ( .A(n6576), .B(n6579), .Z(n6577) );
  IV U6565 ( .A(n6558), .Z(n6562) );
  XOR U6566 ( .A(n6558), .B(n6540), .Z(n6560) );
  XOR U6567 ( .A(n6580), .B(n6581), .Z(n6540) );
  AND U6568 ( .A(n354), .B(n6582), .Z(n6580) );
  XOR U6569 ( .A(n6583), .B(n6581), .Z(n6582) );
  NANDN U6570 ( .A(n6542), .B(n6544), .Z(n6558) );
  XOR U6571 ( .A(n6584), .B(n6585), .Z(n6544) );
  AND U6572 ( .A(n354), .B(n6586), .Z(n6584) );
  XOR U6573 ( .A(n6585), .B(n6587), .Z(n6586) );
  XOR U6574 ( .A(n6588), .B(n6589), .Z(n354) );
  AND U6575 ( .A(n6590), .B(n6591), .Z(n6588) );
  XNOR U6576 ( .A(n6589), .B(n6555), .Z(n6591) );
  XNOR U6577 ( .A(n6592), .B(n6593), .Z(n6555) );
  ANDN U6578 ( .B(n6594), .A(n6595), .Z(n6592) );
  XOR U6579 ( .A(n6593), .B(n6596), .Z(n6594) );
  XOR U6580 ( .A(n6589), .B(n6557), .Z(n6590) );
  XOR U6581 ( .A(n6597), .B(n6598), .Z(n6557) );
  AND U6582 ( .A(n358), .B(n6599), .Z(n6597) );
  XOR U6583 ( .A(n6600), .B(n6598), .Z(n6599) );
  XNOR U6584 ( .A(n6601), .B(n6602), .Z(n6589) );
  NAND U6585 ( .A(n6603), .B(n6604), .Z(n6602) );
  XOR U6586 ( .A(n6605), .B(n6581), .Z(n6604) );
  XOR U6587 ( .A(n6595), .B(n6596), .Z(n6581) );
  XOR U6588 ( .A(n6606), .B(n6607), .Z(n6596) );
  ANDN U6589 ( .B(n6608), .A(n6609), .Z(n6606) );
  XOR U6590 ( .A(n6607), .B(n6610), .Z(n6608) );
  XOR U6591 ( .A(n6611), .B(n6612), .Z(n6595) );
  XOR U6592 ( .A(n6613), .B(n6614), .Z(n6612) );
  ANDN U6593 ( .B(n6615), .A(n6616), .Z(n6613) );
  XOR U6594 ( .A(n6617), .B(n6614), .Z(n6615) );
  IV U6595 ( .A(n6593), .Z(n6611) );
  XOR U6596 ( .A(n6618), .B(n6619), .Z(n6593) );
  ANDN U6597 ( .B(n6620), .A(n6621), .Z(n6618) );
  XOR U6598 ( .A(n6619), .B(n6622), .Z(n6620) );
  IV U6599 ( .A(n6601), .Z(n6605) );
  XOR U6600 ( .A(n6601), .B(n6583), .Z(n6603) );
  XOR U6601 ( .A(n6623), .B(n6624), .Z(n6583) );
  AND U6602 ( .A(n358), .B(n6625), .Z(n6623) );
  XOR U6603 ( .A(n6626), .B(n6624), .Z(n6625) );
  NANDN U6604 ( .A(n6585), .B(n6587), .Z(n6601) );
  XOR U6605 ( .A(n6627), .B(n6628), .Z(n6587) );
  AND U6606 ( .A(n358), .B(n6629), .Z(n6627) );
  XOR U6607 ( .A(n6628), .B(n6630), .Z(n6629) );
  XOR U6608 ( .A(n6631), .B(n6632), .Z(n358) );
  AND U6609 ( .A(n6633), .B(n6634), .Z(n6631) );
  XNOR U6610 ( .A(n6632), .B(n6598), .Z(n6634) );
  XNOR U6611 ( .A(n6635), .B(n6636), .Z(n6598) );
  ANDN U6612 ( .B(n6637), .A(n6638), .Z(n6635) );
  XOR U6613 ( .A(n6636), .B(n6639), .Z(n6637) );
  XOR U6614 ( .A(n6632), .B(n6600), .Z(n6633) );
  XOR U6615 ( .A(n6640), .B(n6641), .Z(n6600) );
  AND U6616 ( .A(n362), .B(n6642), .Z(n6640) );
  XOR U6617 ( .A(n6643), .B(n6641), .Z(n6642) );
  XNOR U6618 ( .A(n6644), .B(n6645), .Z(n6632) );
  NAND U6619 ( .A(n6646), .B(n6647), .Z(n6645) );
  XOR U6620 ( .A(n6648), .B(n6624), .Z(n6647) );
  XOR U6621 ( .A(n6638), .B(n6639), .Z(n6624) );
  XOR U6622 ( .A(n6649), .B(n6650), .Z(n6639) );
  ANDN U6623 ( .B(n6651), .A(n6652), .Z(n6649) );
  XOR U6624 ( .A(n6650), .B(n6653), .Z(n6651) );
  XOR U6625 ( .A(n6654), .B(n6655), .Z(n6638) );
  XOR U6626 ( .A(n6656), .B(n6657), .Z(n6655) );
  ANDN U6627 ( .B(n6658), .A(n6659), .Z(n6656) );
  XOR U6628 ( .A(n6660), .B(n6657), .Z(n6658) );
  IV U6629 ( .A(n6636), .Z(n6654) );
  XOR U6630 ( .A(n6661), .B(n6662), .Z(n6636) );
  ANDN U6631 ( .B(n6663), .A(n6664), .Z(n6661) );
  XOR U6632 ( .A(n6662), .B(n6665), .Z(n6663) );
  IV U6633 ( .A(n6644), .Z(n6648) );
  XOR U6634 ( .A(n6644), .B(n6626), .Z(n6646) );
  XOR U6635 ( .A(n6666), .B(n6667), .Z(n6626) );
  AND U6636 ( .A(n362), .B(n6668), .Z(n6666) );
  XOR U6637 ( .A(n6669), .B(n6667), .Z(n6668) );
  NANDN U6638 ( .A(n6628), .B(n6630), .Z(n6644) );
  XOR U6639 ( .A(n6670), .B(n6671), .Z(n6630) );
  AND U6640 ( .A(n362), .B(n6672), .Z(n6670) );
  XOR U6641 ( .A(n6671), .B(n6673), .Z(n6672) );
  XOR U6642 ( .A(n6674), .B(n6675), .Z(n362) );
  AND U6643 ( .A(n6676), .B(n6677), .Z(n6674) );
  XNOR U6644 ( .A(n6675), .B(n6641), .Z(n6677) );
  XNOR U6645 ( .A(n6678), .B(n6679), .Z(n6641) );
  ANDN U6646 ( .B(n6680), .A(n6681), .Z(n6678) );
  XOR U6647 ( .A(n6679), .B(n6682), .Z(n6680) );
  XOR U6648 ( .A(n6675), .B(n6643), .Z(n6676) );
  XOR U6649 ( .A(n6683), .B(n6684), .Z(n6643) );
  AND U6650 ( .A(n366), .B(n6685), .Z(n6683) );
  XOR U6651 ( .A(n6686), .B(n6684), .Z(n6685) );
  XNOR U6652 ( .A(n6687), .B(n6688), .Z(n6675) );
  NAND U6653 ( .A(n6689), .B(n6690), .Z(n6688) );
  XOR U6654 ( .A(n6691), .B(n6667), .Z(n6690) );
  XOR U6655 ( .A(n6681), .B(n6682), .Z(n6667) );
  XOR U6656 ( .A(n6692), .B(n6693), .Z(n6682) );
  ANDN U6657 ( .B(n6694), .A(n6695), .Z(n6692) );
  XOR U6658 ( .A(n6693), .B(n6696), .Z(n6694) );
  XOR U6659 ( .A(n6697), .B(n6698), .Z(n6681) );
  XOR U6660 ( .A(n6699), .B(n6700), .Z(n6698) );
  ANDN U6661 ( .B(n6701), .A(n6702), .Z(n6699) );
  XOR U6662 ( .A(n6703), .B(n6700), .Z(n6701) );
  IV U6663 ( .A(n6679), .Z(n6697) );
  XOR U6664 ( .A(n6704), .B(n6705), .Z(n6679) );
  ANDN U6665 ( .B(n6706), .A(n6707), .Z(n6704) );
  XOR U6666 ( .A(n6705), .B(n6708), .Z(n6706) );
  IV U6667 ( .A(n6687), .Z(n6691) );
  XOR U6668 ( .A(n6687), .B(n6669), .Z(n6689) );
  XOR U6669 ( .A(n6709), .B(n6710), .Z(n6669) );
  AND U6670 ( .A(n366), .B(n6711), .Z(n6709) );
  XOR U6671 ( .A(n6712), .B(n6710), .Z(n6711) );
  NANDN U6672 ( .A(n6671), .B(n6673), .Z(n6687) );
  XOR U6673 ( .A(n6713), .B(n6714), .Z(n6673) );
  AND U6674 ( .A(n366), .B(n6715), .Z(n6713) );
  XOR U6675 ( .A(n6714), .B(n6716), .Z(n6715) );
  XOR U6676 ( .A(n6717), .B(n6718), .Z(n366) );
  AND U6677 ( .A(n6719), .B(n6720), .Z(n6717) );
  XNOR U6678 ( .A(n6718), .B(n6684), .Z(n6720) );
  XNOR U6679 ( .A(n6721), .B(n6722), .Z(n6684) );
  ANDN U6680 ( .B(n6723), .A(n6724), .Z(n6721) );
  XOR U6681 ( .A(n6722), .B(n6725), .Z(n6723) );
  XOR U6682 ( .A(n6718), .B(n6686), .Z(n6719) );
  XOR U6683 ( .A(n6726), .B(n6727), .Z(n6686) );
  AND U6684 ( .A(n370), .B(n6728), .Z(n6726) );
  XOR U6685 ( .A(n6729), .B(n6727), .Z(n6728) );
  XNOR U6686 ( .A(n6730), .B(n6731), .Z(n6718) );
  NAND U6687 ( .A(n6732), .B(n6733), .Z(n6731) );
  XOR U6688 ( .A(n6734), .B(n6710), .Z(n6733) );
  XOR U6689 ( .A(n6724), .B(n6725), .Z(n6710) );
  XOR U6690 ( .A(n6735), .B(n6736), .Z(n6725) );
  ANDN U6691 ( .B(n6737), .A(n6738), .Z(n6735) );
  XOR U6692 ( .A(n6736), .B(n6739), .Z(n6737) );
  XOR U6693 ( .A(n6740), .B(n6741), .Z(n6724) );
  XOR U6694 ( .A(n6742), .B(n6743), .Z(n6741) );
  ANDN U6695 ( .B(n6744), .A(n6745), .Z(n6742) );
  XOR U6696 ( .A(n6746), .B(n6743), .Z(n6744) );
  IV U6697 ( .A(n6722), .Z(n6740) );
  XOR U6698 ( .A(n6747), .B(n6748), .Z(n6722) );
  ANDN U6699 ( .B(n6749), .A(n6750), .Z(n6747) );
  XOR U6700 ( .A(n6748), .B(n6751), .Z(n6749) );
  IV U6701 ( .A(n6730), .Z(n6734) );
  XOR U6702 ( .A(n6730), .B(n6712), .Z(n6732) );
  XOR U6703 ( .A(n6752), .B(n6753), .Z(n6712) );
  AND U6704 ( .A(n370), .B(n6754), .Z(n6752) );
  XOR U6705 ( .A(n6755), .B(n6753), .Z(n6754) );
  NANDN U6706 ( .A(n6714), .B(n6716), .Z(n6730) );
  XOR U6707 ( .A(n6756), .B(n6757), .Z(n6716) );
  AND U6708 ( .A(n370), .B(n6758), .Z(n6756) );
  XOR U6709 ( .A(n6757), .B(n6759), .Z(n6758) );
  XOR U6710 ( .A(n6760), .B(n6761), .Z(n370) );
  AND U6711 ( .A(n6762), .B(n6763), .Z(n6760) );
  XNOR U6712 ( .A(n6761), .B(n6727), .Z(n6763) );
  XNOR U6713 ( .A(n6764), .B(n6765), .Z(n6727) );
  ANDN U6714 ( .B(n6766), .A(n6767), .Z(n6764) );
  XOR U6715 ( .A(n6765), .B(n6768), .Z(n6766) );
  XOR U6716 ( .A(n6761), .B(n6729), .Z(n6762) );
  XOR U6717 ( .A(n6769), .B(n6770), .Z(n6729) );
  AND U6718 ( .A(n374), .B(n6771), .Z(n6769) );
  XOR U6719 ( .A(n6772), .B(n6770), .Z(n6771) );
  XNOR U6720 ( .A(n6773), .B(n6774), .Z(n6761) );
  NAND U6721 ( .A(n6775), .B(n6776), .Z(n6774) );
  XOR U6722 ( .A(n6777), .B(n6753), .Z(n6776) );
  XOR U6723 ( .A(n6767), .B(n6768), .Z(n6753) );
  XOR U6724 ( .A(n6778), .B(n6779), .Z(n6768) );
  ANDN U6725 ( .B(n6780), .A(n6781), .Z(n6778) );
  XOR U6726 ( .A(n6779), .B(n6782), .Z(n6780) );
  XOR U6727 ( .A(n6783), .B(n6784), .Z(n6767) );
  XOR U6728 ( .A(n6785), .B(n6786), .Z(n6784) );
  ANDN U6729 ( .B(n6787), .A(n6788), .Z(n6785) );
  XOR U6730 ( .A(n6789), .B(n6786), .Z(n6787) );
  IV U6731 ( .A(n6765), .Z(n6783) );
  XOR U6732 ( .A(n6790), .B(n6791), .Z(n6765) );
  ANDN U6733 ( .B(n6792), .A(n6793), .Z(n6790) );
  XOR U6734 ( .A(n6791), .B(n6794), .Z(n6792) );
  IV U6735 ( .A(n6773), .Z(n6777) );
  XOR U6736 ( .A(n6773), .B(n6755), .Z(n6775) );
  XOR U6737 ( .A(n6795), .B(n6796), .Z(n6755) );
  AND U6738 ( .A(n374), .B(n6797), .Z(n6795) );
  XOR U6739 ( .A(n6798), .B(n6796), .Z(n6797) );
  NANDN U6740 ( .A(n6757), .B(n6759), .Z(n6773) );
  XOR U6741 ( .A(n6799), .B(n6800), .Z(n6759) );
  AND U6742 ( .A(n374), .B(n6801), .Z(n6799) );
  XOR U6743 ( .A(n6800), .B(n6802), .Z(n6801) );
  XOR U6744 ( .A(n6803), .B(n6804), .Z(n374) );
  AND U6745 ( .A(n6805), .B(n6806), .Z(n6803) );
  XNOR U6746 ( .A(n6804), .B(n6770), .Z(n6806) );
  XNOR U6747 ( .A(n6807), .B(n6808), .Z(n6770) );
  ANDN U6748 ( .B(n6809), .A(n6810), .Z(n6807) );
  XOR U6749 ( .A(n6808), .B(n6811), .Z(n6809) );
  XOR U6750 ( .A(n6804), .B(n6772), .Z(n6805) );
  XOR U6751 ( .A(n6812), .B(n6813), .Z(n6772) );
  AND U6752 ( .A(n378), .B(n6814), .Z(n6812) );
  XOR U6753 ( .A(n6815), .B(n6813), .Z(n6814) );
  XNOR U6754 ( .A(n6816), .B(n6817), .Z(n6804) );
  NAND U6755 ( .A(n6818), .B(n6819), .Z(n6817) );
  XOR U6756 ( .A(n6820), .B(n6796), .Z(n6819) );
  XOR U6757 ( .A(n6810), .B(n6811), .Z(n6796) );
  XOR U6758 ( .A(n6821), .B(n6822), .Z(n6811) );
  ANDN U6759 ( .B(n6823), .A(n6824), .Z(n6821) );
  XOR U6760 ( .A(n6822), .B(n6825), .Z(n6823) );
  XOR U6761 ( .A(n6826), .B(n6827), .Z(n6810) );
  XOR U6762 ( .A(n6828), .B(n6829), .Z(n6827) );
  ANDN U6763 ( .B(n6830), .A(n6831), .Z(n6828) );
  XOR U6764 ( .A(n6832), .B(n6829), .Z(n6830) );
  IV U6765 ( .A(n6808), .Z(n6826) );
  XOR U6766 ( .A(n6833), .B(n6834), .Z(n6808) );
  ANDN U6767 ( .B(n6835), .A(n6836), .Z(n6833) );
  XOR U6768 ( .A(n6834), .B(n6837), .Z(n6835) );
  IV U6769 ( .A(n6816), .Z(n6820) );
  XOR U6770 ( .A(n6816), .B(n6798), .Z(n6818) );
  XOR U6771 ( .A(n6838), .B(n6839), .Z(n6798) );
  AND U6772 ( .A(n378), .B(n6840), .Z(n6838) );
  XOR U6773 ( .A(n6841), .B(n6839), .Z(n6840) );
  NANDN U6774 ( .A(n6800), .B(n6802), .Z(n6816) );
  XOR U6775 ( .A(n6842), .B(n6843), .Z(n6802) );
  AND U6776 ( .A(n378), .B(n6844), .Z(n6842) );
  XOR U6777 ( .A(n6843), .B(n6845), .Z(n6844) );
  XOR U6778 ( .A(n6846), .B(n6847), .Z(n378) );
  AND U6779 ( .A(n6848), .B(n6849), .Z(n6846) );
  XNOR U6780 ( .A(n6847), .B(n6813), .Z(n6849) );
  XNOR U6781 ( .A(n6850), .B(n6851), .Z(n6813) );
  ANDN U6782 ( .B(n6852), .A(n6853), .Z(n6850) );
  XOR U6783 ( .A(n6851), .B(n6854), .Z(n6852) );
  XOR U6784 ( .A(n6847), .B(n6815), .Z(n6848) );
  XOR U6785 ( .A(n6855), .B(n6856), .Z(n6815) );
  AND U6786 ( .A(n382), .B(n6857), .Z(n6855) );
  XOR U6787 ( .A(n6858), .B(n6856), .Z(n6857) );
  XNOR U6788 ( .A(n6859), .B(n6860), .Z(n6847) );
  NAND U6789 ( .A(n6861), .B(n6862), .Z(n6860) );
  XOR U6790 ( .A(n6863), .B(n6839), .Z(n6862) );
  XOR U6791 ( .A(n6853), .B(n6854), .Z(n6839) );
  XOR U6792 ( .A(n6864), .B(n6865), .Z(n6854) );
  ANDN U6793 ( .B(n6866), .A(n6867), .Z(n6864) );
  XOR U6794 ( .A(n6865), .B(n6868), .Z(n6866) );
  XOR U6795 ( .A(n6869), .B(n6870), .Z(n6853) );
  XOR U6796 ( .A(n6871), .B(n6872), .Z(n6870) );
  ANDN U6797 ( .B(n6873), .A(n6874), .Z(n6871) );
  XOR U6798 ( .A(n6875), .B(n6872), .Z(n6873) );
  IV U6799 ( .A(n6851), .Z(n6869) );
  XOR U6800 ( .A(n6876), .B(n6877), .Z(n6851) );
  ANDN U6801 ( .B(n6878), .A(n6879), .Z(n6876) );
  XOR U6802 ( .A(n6877), .B(n6880), .Z(n6878) );
  IV U6803 ( .A(n6859), .Z(n6863) );
  XOR U6804 ( .A(n6859), .B(n6841), .Z(n6861) );
  XOR U6805 ( .A(n6881), .B(n6882), .Z(n6841) );
  AND U6806 ( .A(n382), .B(n6883), .Z(n6881) );
  XOR U6807 ( .A(n6884), .B(n6882), .Z(n6883) );
  NANDN U6808 ( .A(n6843), .B(n6845), .Z(n6859) );
  XOR U6809 ( .A(n6885), .B(n6886), .Z(n6845) );
  AND U6810 ( .A(n382), .B(n6887), .Z(n6885) );
  XOR U6811 ( .A(n6886), .B(n6888), .Z(n6887) );
  XOR U6812 ( .A(n6889), .B(n6890), .Z(n382) );
  AND U6813 ( .A(n6891), .B(n6892), .Z(n6889) );
  XNOR U6814 ( .A(n6890), .B(n6856), .Z(n6892) );
  XNOR U6815 ( .A(n6893), .B(n6894), .Z(n6856) );
  ANDN U6816 ( .B(n6895), .A(n6896), .Z(n6893) );
  XOR U6817 ( .A(n6894), .B(n6897), .Z(n6895) );
  XOR U6818 ( .A(n6890), .B(n6858), .Z(n6891) );
  XOR U6819 ( .A(n6898), .B(n6899), .Z(n6858) );
  AND U6820 ( .A(n386), .B(n6900), .Z(n6898) );
  XOR U6821 ( .A(n6901), .B(n6899), .Z(n6900) );
  XNOR U6822 ( .A(n6902), .B(n6903), .Z(n6890) );
  NAND U6823 ( .A(n6904), .B(n6905), .Z(n6903) );
  XOR U6824 ( .A(n6906), .B(n6882), .Z(n6905) );
  XOR U6825 ( .A(n6896), .B(n6897), .Z(n6882) );
  XOR U6826 ( .A(n6907), .B(n6908), .Z(n6897) );
  ANDN U6827 ( .B(n6909), .A(n6910), .Z(n6907) );
  XOR U6828 ( .A(n6908), .B(n6911), .Z(n6909) );
  XOR U6829 ( .A(n6912), .B(n6913), .Z(n6896) );
  XOR U6830 ( .A(n6914), .B(n6915), .Z(n6913) );
  ANDN U6831 ( .B(n6916), .A(n6917), .Z(n6914) );
  XOR U6832 ( .A(n6918), .B(n6915), .Z(n6916) );
  IV U6833 ( .A(n6894), .Z(n6912) );
  XOR U6834 ( .A(n6919), .B(n6920), .Z(n6894) );
  ANDN U6835 ( .B(n6921), .A(n6922), .Z(n6919) );
  XOR U6836 ( .A(n6920), .B(n6923), .Z(n6921) );
  IV U6837 ( .A(n6902), .Z(n6906) );
  XOR U6838 ( .A(n6902), .B(n6884), .Z(n6904) );
  XOR U6839 ( .A(n6924), .B(n6925), .Z(n6884) );
  AND U6840 ( .A(n386), .B(n6926), .Z(n6924) );
  XOR U6841 ( .A(n6927), .B(n6925), .Z(n6926) );
  NANDN U6842 ( .A(n6886), .B(n6888), .Z(n6902) );
  XOR U6843 ( .A(n6928), .B(n6929), .Z(n6888) );
  AND U6844 ( .A(n386), .B(n6930), .Z(n6928) );
  XOR U6845 ( .A(n6929), .B(n6931), .Z(n6930) );
  XOR U6846 ( .A(n6932), .B(n6933), .Z(n386) );
  AND U6847 ( .A(n6934), .B(n6935), .Z(n6932) );
  XNOR U6848 ( .A(n6933), .B(n6899), .Z(n6935) );
  XNOR U6849 ( .A(n6936), .B(n6937), .Z(n6899) );
  ANDN U6850 ( .B(n6938), .A(n6939), .Z(n6936) );
  XOR U6851 ( .A(n6937), .B(n6940), .Z(n6938) );
  XOR U6852 ( .A(n6933), .B(n6901), .Z(n6934) );
  XOR U6853 ( .A(n6941), .B(n6942), .Z(n6901) );
  AND U6854 ( .A(n390), .B(n6943), .Z(n6941) );
  XOR U6855 ( .A(n6944), .B(n6942), .Z(n6943) );
  XNOR U6856 ( .A(n6945), .B(n6946), .Z(n6933) );
  NAND U6857 ( .A(n6947), .B(n6948), .Z(n6946) );
  XOR U6858 ( .A(n6949), .B(n6925), .Z(n6948) );
  XOR U6859 ( .A(n6939), .B(n6940), .Z(n6925) );
  XOR U6860 ( .A(n6950), .B(n6951), .Z(n6940) );
  ANDN U6861 ( .B(n6952), .A(n6953), .Z(n6950) );
  XOR U6862 ( .A(n6951), .B(n6954), .Z(n6952) );
  XOR U6863 ( .A(n6955), .B(n6956), .Z(n6939) );
  XOR U6864 ( .A(n6957), .B(n6958), .Z(n6956) );
  ANDN U6865 ( .B(n6959), .A(n6960), .Z(n6957) );
  XOR U6866 ( .A(n6961), .B(n6958), .Z(n6959) );
  IV U6867 ( .A(n6937), .Z(n6955) );
  XOR U6868 ( .A(n6962), .B(n6963), .Z(n6937) );
  ANDN U6869 ( .B(n6964), .A(n6965), .Z(n6962) );
  XOR U6870 ( .A(n6963), .B(n6966), .Z(n6964) );
  IV U6871 ( .A(n6945), .Z(n6949) );
  XOR U6872 ( .A(n6945), .B(n6927), .Z(n6947) );
  XOR U6873 ( .A(n6967), .B(n6968), .Z(n6927) );
  AND U6874 ( .A(n390), .B(n6969), .Z(n6967) );
  XOR U6875 ( .A(n6970), .B(n6968), .Z(n6969) );
  NANDN U6876 ( .A(n6929), .B(n6931), .Z(n6945) );
  XOR U6877 ( .A(n6971), .B(n6972), .Z(n6931) );
  AND U6878 ( .A(n390), .B(n6973), .Z(n6971) );
  XOR U6879 ( .A(n6972), .B(n6974), .Z(n6973) );
  XOR U6880 ( .A(n6975), .B(n6976), .Z(n390) );
  AND U6881 ( .A(n6977), .B(n6978), .Z(n6975) );
  XNOR U6882 ( .A(n6976), .B(n6942), .Z(n6978) );
  XNOR U6883 ( .A(n6979), .B(n6980), .Z(n6942) );
  ANDN U6884 ( .B(n6981), .A(n6982), .Z(n6979) );
  XOR U6885 ( .A(n6980), .B(n6983), .Z(n6981) );
  XOR U6886 ( .A(n6976), .B(n6944), .Z(n6977) );
  XOR U6887 ( .A(n6984), .B(n6985), .Z(n6944) );
  AND U6888 ( .A(n394), .B(n6986), .Z(n6984) );
  XOR U6889 ( .A(n6987), .B(n6985), .Z(n6986) );
  XNOR U6890 ( .A(n6988), .B(n6989), .Z(n6976) );
  NAND U6891 ( .A(n6990), .B(n6991), .Z(n6989) );
  XOR U6892 ( .A(n6992), .B(n6968), .Z(n6991) );
  XOR U6893 ( .A(n6982), .B(n6983), .Z(n6968) );
  XOR U6894 ( .A(n6993), .B(n6994), .Z(n6983) );
  ANDN U6895 ( .B(n6995), .A(n6996), .Z(n6993) );
  XOR U6896 ( .A(n6994), .B(n6997), .Z(n6995) );
  XOR U6897 ( .A(n6998), .B(n6999), .Z(n6982) );
  XOR U6898 ( .A(n7000), .B(n7001), .Z(n6999) );
  ANDN U6899 ( .B(n7002), .A(n7003), .Z(n7000) );
  XOR U6900 ( .A(n7004), .B(n7001), .Z(n7002) );
  IV U6901 ( .A(n6980), .Z(n6998) );
  XOR U6902 ( .A(n7005), .B(n7006), .Z(n6980) );
  ANDN U6903 ( .B(n7007), .A(n7008), .Z(n7005) );
  XOR U6904 ( .A(n7006), .B(n7009), .Z(n7007) );
  IV U6905 ( .A(n6988), .Z(n6992) );
  XOR U6906 ( .A(n6988), .B(n6970), .Z(n6990) );
  XOR U6907 ( .A(n7010), .B(n7011), .Z(n6970) );
  AND U6908 ( .A(n394), .B(n7012), .Z(n7010) );
  XOR U6909 ( .A(n7013), .B(n7011), .Z(n7012) );
  NANDN U6910 ( .A(n6972), .B(n6974), .Z(n6988) );
  XOR U6911 ( .A(n7014), .B(n7015), .Z(n6974) );
  AND U6912 ( .A(n394), .B(n7016), .Z(n7014) );
  XOR U6913 ( .A(n7015), .B(n7017), .Z(n7016) );
  XOR U6914 ( .A(n7018), .B(n7019), .Z(n394) );
  AND U6915 ( .A(n7020), .B(n7021), .Z(n7018) );
  XNOR U6916 ( .A(n7019), .B(n6985), .Z(n7021) );
  XNOR U6917 ( .A(n7022), .B(n7023), .Z(n6985) );
  ANDN U6918 ( .B(n7024), .A(n7025), .Z(n7022) );
  XOR U6919 ( .A(n7023), .B(n7026), .Z(n7024) );
  XOR U6920 ( .A(n7019), .B(n6987), .Z(n7020) );
  XOR U6921 ( .A(n7027), .B(n7028), .Z(n6987) );
  AND U6922 ( .A(n398), .B(n7029), .Z(n7027) );
  XOR U6923 ( .A(n7030), .B(n7028), .Z(n7029) );
  XNOR U6924 ( .A(n7031), .B(n7032), .Z(n7019) );
  NAND U6925 ( .A(n7033), .B(n7034), .Z(n7032) );
  XOR U6926 ( .A(n7035), .B(n7011), .Z(n7034) );
  XOR U6927 ( .A(n7025), .B(n7026), .Z(n7011) );
  XOR U6928 ( .A(n7036), .B(n7037), .Z(n7026) );
  ANDN U6929 ( .B(n7038), .A(n7039), .Z(n7036) );
  XOR U6930 ( .A(n7037), .B(n7040), .Z(n7038) );
  XOR U6931 ( .A(n7041), .B(n7042), .Z(n7025) );
  XOR U6932 ( .A(n7043), .B(n7044), .Z(n7042) );
  ANDN U6933 ( .B(n7045), .A(n7046), .Z(n7043) );
  XOR U6934 ( .A(n7047), .B(n7044), .Z(n7045) );
  IV U6935 ( .A(n7023), .Z(n7041) );
  XOR U6936 ( .A(n7048), .B(n7049), .Z(n7023) );
  ANDN U6937 ( .B(n7050), .A(n7051), .Z(n7048) );
  XOR U6938 ( .A(n7049), .B(n7052), .Z(n7050) );
  IV U6939 ( .A(n7031), .Z(n7035) );
  XOR U6940 ( .A(n7031), .B(n7013), .Z(n7033) );
  XOR U6941 ( .A(n7053), .B(n7054), .Z(n7013) );
  AND U6942 ( .A(n398), .B(n7055), .Z(n7053) );
  XOR U6943 ( .A(n7056), .B(n7054), .Z(n7055) );
  NANDN U6944 ( .A(n7015), .B(n7017), .Z(n7031) );
  XOR U6945 ( .A(n7057), .B(n7058), .Z(n7017) );
  AND U6946 ( .A(n398), .B(n7059), .Z(n7057) );
  XOR U6947 ( .A(n7058), .B(n7060), .Z(n7059) );
  XOR U6948 ( .A(n7061), .B(n7062), .Z(n398) );
  AND U6949 ( .A(n7063), .B(n7064), .Z(n7061) );
  XNOR U6950 ( .A(n7062), .B(n7028), .Z(n7064) );
  XNOR U6951 ( .A(n7065), .B(n7066), .Z(n7028) );
  ANDN U6952 ( .B(n7067), .A(n7068), .Z(n7065) );
  XOR U6953 ( .A(n7066), .B(n7069), .Z(n7067) );
  XOR U6954 ( .A(n7062), .B(n7030), .Z(n7063) );
  XOR U6955 ( .A(n7070), .B(n7071), .Z(n7030) );
  AND U6956 ( .A(n402), .B(n7072), .Z(n7070) );
  XOR U6957 ( .A(n7073), .B(n7071), .Z(n7072) );
  XNOR U6958 ( .A(n7074), .B(n7075), .Z(n7062) );
  NAND U6959 ( .A(n7076), .B(n7077), .Z(n7075) );
  XOR U6960 ( .A(n7078), .B(n7054), .Z(n7077) );
  XOR U6961 ( .A(n7068), .B(n7069), .Z(n7054) );
  XOR U6962 ( .A(n7079), .B(n7080), .Z(n7069) );
  ANDN U6963 ( .B(n7081), .A(n7082), .Z(n7079) );
  XOR U6964 ( .A(n7080), .B(n7083), .Z(n7081) );
  XOR U6965 ( .A(n7084), .B(n7085), .Z(n7068) );
  XOR U6966 ( .A(n7086), .B(n7087), .Z(n7085) );
  ANDN U6967 ( .B(n7088), .A(n7089), .Z(n7086) );
  XOR U6968 ( .A(n7090), .B(n7087), .Z(n7088) );
  IV U6969 ( .A(n7066), .Z(n7084) );
  XOR U6970 ( .A(n7091), .B(n7092), .Z(n7066) );
  ANDN U6971 ( .B(n7093), .A(n7094), .Z(n7091) );
  XOR U6972 ( .A(n7092), .B(n7095), .Z(n7093) );
  IV U6973 ( .A(n7074), .Z(n7078) );
  XOR U6974 ( .A(n7074), .B(n7056), .Z(n7076) );
  XOR U6975 ( .A(n7096), .B(n7097), .Z(n7056) );
  AND U6976 ( .A(n402), .B(n7098), .Z(n7096) );
  XOR U6977 ( .A(n7099), .B(n7097), .Z(n7098) );
  NANDN U6978 ( .A(n7058), .B(n7060), .Z(n7074) );
  XOR U6979 ( .A(n7100), .B(n7101), .Z(n7060) );
  AND U6980 ( .A(n402), .B(n7102), .Z(n7100) );
  XOR U6981 ( .A(n7101), .B(n7103), .Z(n7102) );
  XOR U6982 ( .A(n7104), .B(n7105), .Z(n402) );
  AND U6983 ( .A(n7106), .B(n7107), .Z(n7104) );
  XNOR U6984 ( .A(n7105), .B(n7071), .Z(n7107) );
  XNOR U6985 ( .A(n7108), .B(n7109), .Z(n7071) );
  ANDN U6986 ( .B(n7110), .A(n7111), .Z(n7108) );
  XOR U6987 ( .A(n7109), .B(n7112), .Z(n7110) );
  XOR U6988 ( .A(n7105), .B(n7073), .Z(n7106) );
  XOR U6989 ( .A(n7113), .B(n7114), .Z(n7073) );
  AND U6990 ( .A(n406), .B(n7115), .Z(n7113) );
  XOR U6991 ( .A(n7116), .B(n7114), .Z(n7115) );
  XNOR U6992 ( .A(n7117), .B(n7118), .Z(n7105) );
  NAND U6993 ( .A(n7119), .B(n7120), .Z(n7118) );
  XOR U6994 ( .A(n7121), .B(n7097), .Z(n7120) );
  XOR U6995 ( .A(n7111), .B(n7112), .Z(n7097) );
  XOR U6996 ( .A(n7122), .B(n7123), .Z(n7112) );
  ANDN U6997 ( .B(n7124), .A(n7125), .Z(n7122) );
  XOR U6998 ( .A(n7123), .B(n7126), .Z(n7124) );
  XOR U6999 ( .A(n7127), .B(n7128), .Z(n7111) );
  XOR U7000 ( .A(n7129), .B(n7130), .Z(n7128) );
  ANDN U7001 ( .B(n7131), .A(n7132), .Z(n7129) );
  XOR U7002 ( .A(n7133), .B(n7130), .Z(n7131) );
  IV U7003 ( .A(n7109), .Z(n7127) );
  XOR U7004 ( .A(n7134), .B(n7135), .Z(n7109) );
  ANDN U7005 ( .B(n7136), .A(n7137), .Z(n7134) );
  XOR U7006 ( .A(n7135), .B(n7138), .Z(n7136) );
  IV U7007 ( .A(n7117), .Z(n7121) );
  XOR U7008 ( .A(n7117), .B(n7099), .Z(n7119) );
  XOR U7009 ( .A(n7139), .B(n7140), .Z(n7099) );
  AND U7010 ( .A(n406), .B(n7141), .Z(n7139) );
  XOR U7011 ( .A(n7142), .B(n7140), .Z(n7141) );
  NANDN U7012 ( .A(n7101), .B(n7103), .Z(n7117) );
  XOR U7013 ( .A(n7143), .B(n7144), .Z(n7103) );
  AND U7014 ( .A(n406), .B(n7145), .Z(n7143) );
  XOR U7015 ( .A(n7144), .B(n7146), .Z(n7145) );
  XOR U7016 ( .A(n7147), .B(n7148), .Z(n406) );
  AND U7017 ( .A(n7149), .B(n7150), .Z(n7147) );
  XNOR U7018 ( .A(n7148), .B(n7114), .Z(n7150) );
  XNOR U7019 ( .A(n7151), .B(n7152), .Z(n7114) );
  ANDN U7020 ( .B(n7153), .A(n7154), .Z(n7151) );
  XOR U7021 ( .A(n7152), .B(n7155), .Z(n7153) );
  XOR U7022 ( .A(n7148), .B(n7116), .Z(n7149) );
  XOR U7023 ( .A(n7156), .B(n7157), .Z(n7116) );
  AND U7024 ( .A(n410), .B(n7158), .Z(n7156) );
  XOR U7025 ( .A(n7159), .B(n7157), .Z(n7158) );
  XNOR U7026 ( .A(n7160), .B(n7161), .Z(n7148) );
  NAND U7027 ( .A(n7162), .B(n7163), .Z(n7161) );
  XOR U7028 ( .A(n7164), .B(n7140), .Z(n7163) );
  XOR U7029 ( .A(n7154), .B(n7155), .Z(n7140) );
  XOR U7030 ( .A(n7165), .B(n7166), .Z(n7155) );
  ANDN U7031 ( .B(n7167), .A(n7168), .Z(n7165) );
  XOR U7032 ( .A(n7166), .B(n7169), .Z(n7167) );
  XOR U7033 ( .A(n7170), .B(n7171), .Z(n7154) );
  XOR U7034 ( .A(n7172), .B(n7173), .Z(n7171) );
  ANDN U7035 ( .B(n7174), .A(n7175), .Z(n7172) );
  XOR U7036 ( .A(n7176), .B(n7173), .Z(n7174) );
  IV U7037 ( .A(n7152), .Z(n7170) );
  XOR U7038 ( .A(n7177), .B(n7178), .Z(n7152) );
  ANDN U7039 ( .B(n7179), .A(n7180), .Z(n7177) );
  XOR U7040 ( .A(n7178), .B(n7181), .Z(n7179) );
  IV U7041 ( .A(n7160), .Z(n7164) );
  XOR U7042 ( .A(n7160), .B(n7142), .Z(n7162) );
  XOR U7043 ( .A(n7182), .B(n7183), .Z(n7142) );
  AND U7044 ( .A(n410), .B(n7184), .Z(n7182) );
  XOR U7045 ( .A(n7185), .B(n7183), .Z(n7184) );
  NANDN U7046 ( .A(n7144), .B(n7146), .Z(n7160) );
  XOR U7047 ( .A(n7186), .B(n7187), .Z(n7146) );
  AND U7048 ( .A(n410), .B(n7188), .Z(n7186) );
  XOR U7049 ( .A(n7187), .B(n7189), .Z(n7188) );
  XOR U7050 ( .A(n7190), .B(n7191), .Z(n410) );
  AND U7051 ( .A(n7192), .B(n7193), .Z(n7190) );
  XNOR U7052 ( .A(n7191), .B(n7157), .Z(n7193) );
  XNOR U7053 ( .A(n7194), .B(n7195), .Z(n7157) );
  ANDN U7054 ( .B(n7196), .A(n7197), .Z(n7194) );
  XOR U7055 ( .A(n7195), .B(n7198), .Z(n7196) );
  XOR U7056 ( .A(n7191), .B(n7159), .Z(n7192) );
  XOR U7057 ( .A(n7199), .B(n7200), .Z(n7159) );
  AND U7058 ( .A(n414), .B(n7201), .Z(n7199) );
  XOR U7059 ( .A(n7202), .B(n7200), .Z(n7201) );
  XNOR U7060 ( .A(n7203), .B(n7204), .Z(n7191) );
  NAND U7061 ( .A(n7205), .B(n7206), .Z(n7204) );
  XOR U7062 ( .A(n7207), .B(n7183), .Z(n7206) );
  XOR U7063 ( .A(n7197), .B(n7198), .Z(n7183) );
  XOR U7064 ( .A(n7208), .B(n7209), .Z(n7198) );
  ANDN U7065 ( .B(n7210), .A(n7211), .Z(n7208) );
  XOR U7066 ( .A(n7209), .B(n7212), .Z(n7210) );
  XOR U7067 ( .A(n7213), .B(n7214), .Z(n7197) );
  XOR U7068 ( .A(n7215), .B(n7216), .Z(n7214) );
  ANDN U7069 ( .B(n7217), .A(n7218), .Z(n7215) );
  XOR U7070 ( .A(n7219), .B(n7216), .Z(n7217) );
  IV U7071 ( .A(n7195), .Z(n7213) );
  XOR U7072 ( .A(n7220), .B(n7221), .Z(n7195) );
  ANDN U7073 ( .B(n7222), .A(n7223), .Z(n7220) );
  XOR U7074 ( .A(n7221), .B(n7224), .Z(n7222) );
  IV U7075 ( .A(n7203), .Z(n7207) );
  XOR U7076 ( .A(n7203), .B(n7185), .Z(n7205) );
  XOR U7077 ( .A(n7225), .B(n7226), .Z(n7185) );
  AND U7078 ( .A(n414), .B(n7227), .Z(n7225) );
  XOR U7079 ( .A(n7228), .B(n7226), .Z(n7227) );
  NANDN U7080 ( .A(n7187), .B(n7189), .Z(n7203) );
  XOR U7081 ( .A(n7229), .B(n7230), .Z(n7189) );
  AND U7082 ( .A(n414), .B(n7231), .Z(n7229) );
  XOR U7083 ( .A(n7230), .B(n7232), .Z(n7231) );
  XOR U7084 ( .A(n7233), .B(n7234), .Z(n414) );
  AND U7085 ( .A(n7235), .B(n7236), .Z(n7233) );
  XNOR U7086 ( .A(n7234), .B(n7200), .Z(n7236) );
  XNOR U7087 ( .A(n7237), .B(n7238), .Z(n7200) );
  ANDN U7088 ( .B(n7239), .A(n7240), .Z(n7237) );
  XOR U7089 ( .A(n7238), .B(n7241), .Z(n7239) );
  XOR U7090 ( .A(n7234), .B(n7202), .Z(n7235) );
  XOR U7091 ( .A(n7242), .B(n7243), .Z(n7202) );
  AND U7092 ( .A(n418), .B(n7244), .Z(n7242) );
  XOR U7093 ( .A(n7245), .B(n7243), .Z(n7244) );
  XNOR U7094 ( .A(n7246), .B(n7247), .Z(n7234) );
  NAND U7095 ( .A(n7248), .B(n7249), .Z(n7247) );
  XOR U7096 ( .A(n7250), .B(n7226), .Z(n7249) );
  XOR U7097 ( .A(n7240), .B(n7241), .Z(n7226) );
  XOR U7098 ( .A(n7251), .B(n7252), .Z(n7241) );
  ANDN U7099 ( .B(n7253), .A(n7254), .Z(n7251) );
  XOR U7100 ( .A(n7252), .B(n7255), .Z(n7253) );
  XOR U7101 ( .A(n7256), .B(n7257), .Z(n7240) );
  XOR U7102 ( .A(n7258), .B(n7259), .Z(n7257) );
  ANDN U7103 ( .B(n7260), .A(n7261), .Z(n7258) );
  XOR U7104 ( .A(n7262), .B(n7259), .Z(n7260) );
  IV U7105 ( .A(n7238), .Z(n7256) );
  XOR U7106 ( .A(n7263), .B(n7264), .Z(n7238) );
  ANDN U7107 ( .B(n7265), .A(n7266), .Z(n7263) );
  XOR U7108 ( .A(n7264), .B(n7267), .Z(n7265) );
  IV U7109 ( .A(n7246), .Z(n7250) );
  XOR U7110 ( .A(n7246), .B(n7228), .Z(n7248) );
  XOR U7111 ( .A(n7268), .B(n7269), .Z(n7228) );
  AND U7112 ( .A(n418), .B(n7270), .Z(n7268) );
  XOR U7113 ( .A(n7271), .B(n7269), .Z(n7270) );
  NANDN U7114 ( .A(n7230), .B(n7232), .Z(n7246) );
  XOR U7115 ( .A(n7272), .B(n7273), .Z(n7232) );
  AND U7116 ( .A(n418), .B(n7274), .Z(n7272) );
  XOR U7117 ( .A(n7273), .B(n7275), .Z(n7274) );
  XOR U7118 ( .A(n7276), .B(n7277), .Z(n418) );
  AND U7119 ( .A(n7278), .B(n7279), .Z(n7276) );
  XNOR U7120 ( .A(n7277), .B(n7243), .Z(n7279) );
  XNOR U7121 ( .A(n7280), .B(n7281), .Z(n7243) );
  ANDN U7122 ( .B(n7282), .A(n7283), .Z(n7280) );
  XOR U7123 ( .A(n7281), .B(n7284), .Z(n7282) );
  XOR U7124 ( .A(n7277), .B(n7245), .Z(n7278) );
  XOR U7125 ( .A(n7285), .B(n7286), .Z(n7245) );
  AND U7126 ( .A(n422), .B(n7287), .Z(n7285) );
  XOR U7127 ( .A(n7288), .B(n7286), .Z(n7287) );
  XNOR U7128 ( .A(n7289), .B(n7290), .Z(n7277) );
  NAND U7129 ( .A(n7291), .B(n7292), .Z(n7290) );
  XOR U7130 ( .A(n7293), .B(n7269), .Z(n7292) );
  XOR U7131 ( .A(n7283), .B(n7284), .Z(n7269) );
  XOR U7132 ( .A(n7294), .B(n7295), .Z(n7284) );
  ANDN U7133 ( .B(n7296), .A(n7297), .Z(n7294) );
  XOR U7134 ( .A(n7295), .B(n7298), .Z(n7296) );
  XOR U7135 ( .A(n7299), .B(n7300), .Z(n7283) );
  XOR U7136 ( .A(n7301), .B(n7302), .Z(n7300) );
  ANDN U7137 ( .B(n7303), .A(n7304), .Z(n7301) );
  XOR U7138 ( .A(n7305), .B(n7302), .Z(n7303) );
  IV U7139 ( .A(n7281), .Z(n7299) );
  XOR U7140 ( .A(n7306), .B(n7307), .Z(n7281) );
  ANDN U7141 ( .B(n7308), .A(n7309), .Z(n7306) );
  XOR U7142 ( .A(n7307), .B(n7310), .Z(n7308) );
  IV U7143 ( .A(n7289), .Z(n7293) );
  XOR U7144 ( .A(n7289), .B(n7271), .Z(n7291) );
  XOR U7145 ( .A(n7311), .B(n7312), .Z(n7271) );
  AND U7146 ( .A(n422), .B(n7313), .Z(n7311) );
  XOR U7147 ( .A(n7314), .B(n7312), .Z(n7313) );
  NANDN U7148 ( .A(n7273), .B(n7275), .Z(n7289) );
  XOR U7149 ( .A(n7315), .B(n7316), .Z(n7275) );
  AND U7150 ( .A(n422), .B(n7317), .Z(n7315) );
  XOR U7151 ( .A(n7316), .B(n7318), .Z(n7317) );
  XOR U7152 ( .A(n7319), .B(n7320), .Z(n422) );
  AND U7153 ( .A(n7321), .B(n7322), .Z(n7319) );
  XNOR U7154 ( .A(n7320), .B(n7286), .Z(n7322) );
  XNOR U7155 ( .A(n7323), .B(n7324), .Z(n7286) );
  ANDN U7156 ( .B(n7325), .A(n7326), .Z(n7323) );
  XOR U7157 ( .A(n7324), .B(n7327), .Z(n7325) );
  XOR U7158 ( .A(n7320), .B(n7288), .Z(n7321) );
  XOR U7159 ( .A(n7328), .B(n7329), .Z(n7288) );
  AND U7160 ( .A(n426), .B(n7330), .Z(n7328) );
  XOR U7161 ( .A(n7331), .B(n7329), .Z(n7330) );
  XNOR U7162 ( .A(n7332), .B(n7333), .Z(n7320) );
  NAND U7163 ( .A(n7334), .B(n7335), .Z(n7333) );
  XOR U7164 ( .A(n7336), .B(n7312), .Z(n7335) );
  XOR U7165 ( .A(n7326), .B(n7327), .Z(n7312) );
  XOR U7166 ( .A(n7337), .B(n7338), .Z(n7327) );
  ANDN U7167 ( .B(n7339), .A(n7340), .Z(n7337) );
  XOR U7168 ( .A(n7338), .B(n7341), .Z(n7339) );
  XOR U7169 ( .A(n7342), .B(n7343), .Z(n7326) );
  XOR U7170 ( .A(n7344), .B(n7345), .Z(n7343) );
  ANDN U7171 ( .B(n7346), .A(n7347), .Z(n7344) );
  XOR U7172 ( .A(n7348), .B(n7345), .Z(n7346) );
  IV U7173 ( .A(n7324), .Z(n7342) );
  XOR U7174 ( .A(n7349), .B(n7350), .Z(n7324) );
  ANDN U7175 ( .B(n7351), .A(n7352), .Z(n7349) );
  XOR U7176 ( .A(n7350), .B(n7353), .Z(n7351) );
  IV U7177 ( .A(n7332), .Z(n7336) );
  XOR U7178 ( .A(n7332), .B(n7314), .Z(n7334) );
  XOR U7179 ( .A(n7354), .B(n7355), .Z(n7314) );
  AND U7180 ( .A(n426), .B(n7356), .Z(n7354) );
  XOR U7181 ( .A(n7357), .B(n7355), .Z(n7356) );
  NANDN U7182 ( .A(n7316), .B(n7318), .Z(n7332) );
  XOR U7183 ( .A(n7358), .B(n7359), .Z(n7318) );
  AND U7184 ( .A(n426), .B(n7360), .Z(n7358) );
  XOR U7185 ( .A(n7359), .B(n7361), .Z(n7360) );
  XOR U7186 ( .A(n7362), .B(n7363), .Z(n426) );
  AND U7187 ( .A(n7364), .B(n7365), .Z(n7362) );
  XNOR U7188 ( .A(n7363), .B(n7329), .Z(n7365) );
  XNOR U7189 ( .A(n7366), .B(n7367), .Z(n7329) );
  ANDN U7190 ( .B(n7368), .A(n7369), .Z(n7366) );
  XOR U7191 ( .A(n7367), .B(n7370), .Z(n7368) );
  XOR U7192 ( .A(n7363), .B(n7331), .Z(n7364) );
  XOR U7193 ( .A(n7371), .B(n7372), .Z(n7331) );
  AND U7194 ( .A(n430), .B(n7373), .Z(n7371) );
  XOR U7195 ( .A(n7374), .B(n7372), .Z(n7373) );
  XNOR U7196 ( .A(n7375), .B(n7376), .Z(n7363) );
  NAND U7197 ( .A(n7377), .B(n7378), .Z(n7376) );
  XOR U7198 ( .A(n7379), .B(n7355), .Z(n7378) );
  XOR U7199 ( .A(n7369), .B(n7370), .Z(n7355) );
  XOR U7200 ( .A(n7380), .B(n7381), .Z(n7370) );
  ANDN U7201 ( .B(n7382), .A(n7383), .Z(n7380) );
  XOR U7202 ( .A(n7381), .B(n7384), .Z(n7382) );
  XOR U7203 ( .A(n7385), .B(n7386), .Z(n7369) );
  XOR U7204 ( .A(n7387), .B(n7388), .Z(n7386) );
  ANDN U7205 ( .B(n7389), .A(n7390), .Z(n7387) );
  XOR U7206 ( .A(n7391), .B(n7388), .Z(n7389) );
  IV U7207 ( .A(n7367), .Z(n7385) );
  XOR U7208 ( .A(n7392), .B(n7393), .Z(n7367) );
  ANDN U7209 ( .B(n7394), .A(n7395), .Z(n7392) );
  XOR U7210 ( .A(n7393), .B(n7396), .Z(n7394) );
  IV U7211 ( .A(n7375), .Z(n7379) );
  XOR U7212 ( .A(n7375), .B(n7357), .Z(n7377) );
  XOR U7213 ( .A(n7397), .B(n7398), .Z(n7357) );
  AND U7214 ( .A(n430), .B(n7399), .Z(n7397) );
  XOR U7215 ( .A(n7400), .B(n7398), .Z(n7399) );
  NANDN U7216 ( .A(n7359), .B(n7361), .Z(n7375) );
  XOR U7217 ( .A(n7401), .B(n7402), .Z(n7361) );
  AND U7218 ( .A(n430), .B(n7403), .Z(n7401) );
  XOR U7219 ( .A(n7402), .B(n7404), .Z(n7403) );
  XOR U7220 ( .A(n7405), .B(n7406), .Z(n430) );
  AND U7221 ( .A(n7407), .B(n7408), .Z(n7405) );
  XNOR U7222 ( .A(n7406), .B(n7372), .Z(n7408) );
  XNOR U7223 ( .A(n7409), .B(n7410), .Z(n7372) );
  ANDN U7224 ( .B(n7411), .A(n7412), .Z(n7409) );
  XOR U7225 ( .A(n7410), .B(n7413), .Z(n7411) );
  XOR U7226 ( .A(n7406), .B(n7374), .Z(n7407) );
  XOR U7227 ( .A(n7414), .B(n7415), .Z(n7374) );
  AND U7228 ( .A(n434), .B(n7416), .Z(n7414) );
  XOR U7229 ( .A(n7417), .B(n7415), .Z(n7416) );
  XNOR U7230 ( .A(n7418), .B(n7419), .Z(n7406) );
  NAND U7231 ( .A(n7420), .B(n7421), .Z(n7419) );
  XOR U7232 ( .A(n7422), .B(n7398), .Z(n7421) );
  XOR U7233 ( .A(n7412), .B(n7413), .Z(n7398) );
  XOR U7234 ( .A(n7423), .B(n7424), .Z(n7413) );
  ANDN U7235 ( .B(n7425), .A(n7426), .Z(n7423) );
  XOR U7236 ( .A(n7424), .B(n7427), .Z(n7425) );
  XOR U7237 ( .A(n7428), .B(n7429), .Z(n7412) );
  XOR U7238 ( .A(n7430), .B(n7431), .Z(n7429) );
  ANDN U7239 ( .B(n7432), .A(n7433), .Z(n7430) );
  XOR U7240 ( .A(n7434), .B(n7431), .Z(n7432) );
  IV U7241 ( .A(n7410), .Z(n7428) );
  XOR U7242 ( .A(n7435), .B(n7436), .Z(n7410) );
  ANDN U7243 ( .B(n7437), .A(n7438), .Z(n7435) );
  XOR U7244 ( .A(n7436), .B(n7439), .Z(n7437) );
  IV U7245 ( .A(n7418), .Z(n7422) );
  XOR U7246 ( .A(n7418), .B(n7400), .Z(n7420) );
  XOR U7247 ( .A(n7440), .B(n7441), .Z(n7400) );
  AND U7248 ( .A(n434), .B(n7442), .Z(n7440) );
  XOR U7249 ( .A(n7443), .B(n7441), .Z(n7442) );
  NANDN U7250 ( .A(n7402), .B(n7404), .Z(n7418) );
  XOR U7251 ( .A(n7444), .B(n7445), .Z(n7404) );
  AND U7252 ( .A(n434), .B(n7446), .Z(n7444) );
  XOR U7253 ( .A(n7445), .B(n7447), .Z(n7446) );
  XOR U7254 ( .A(n7448), .B(n7449), .Z(n434) );
  AND U7255 ( .A(n7450), .B(n7451), .Z(n7448) );
  XNOR U7256 ( .A(n7449), .B(n7415), .Z(n7451) );
  XNOR U7257 ( .A(n7452), .B(n7453), .Z(n7415) );
  ANDN U7258 ( .B(n7454), .A(n7455), .Z(n7452) );
  XOR U7259 ( .A(n7453), .B(n7456), .Z(n7454) );
  XOR U7260 ( .A(n7449), .B(n7417), .Z(n7450) );
  XOR U7261 ( .A(n7457), .B(n7458), .Z(n7417) );
  AND U7262 ( .A(n438), .B(n7459), .Z(n7457) );
  XOR U7263 ( .A(n7460), .B(n7458), .Z(n7459) );
  XNOR U7264 ( .A(n7461), .B(n7462), .Z(n7449) );
  NAND U7265 ( .A(n7463), .B(n7464), .Z(n7462) );
  XOR U7266 ( .A(n7465), .B(n7441), .Z(n7464) );
  XOR U7267 ( .A(n7455), .B(n7456), .Z(n7441) );
  XOR U7268 ( .A(n7466), .B(n7467), .Z(n7456) );
  ANDN U7269 ( .B(n7468), .A(n7469), .Z(n7466) );
  XOR U7270 ( .A(n7467), .B(n7470), .Z(n7468) );
  XOR U7271 ( .A(n7471), .B(n7472), .Z(n7455) );
  XOR U7272 ( .A(n7473), .B(n7474), .Z(n7472) );
  ANDN U7273 ( .B(n7475), .A(n7476), .Z(n7473) );
  XOR U7274 ( .A(n7477), .B(n7474), .Z(n7475) );
  IV U7275 ( .A(n7453), .Z(n7471) );
  XOR U7276 ( .A(n7478), .B(n7479), .Z(n7453) );
  ANDN U7277 ( .B(n7480), .A(n7481), .Z(n7478) );
  XOR U7278 ( .A(n7479), .B(n7482), .Z(n7480) );
  IV U7279 ( .A(n7461), .Z(n7465) );
  XOR U7280 ( .A(n7461), .B(n7443), .Z(n7463) );
  XOR U7281 ( .A(n7483), .B(n7484), .Z(n7443) );
  AND U7282 ( .A(n438), .B(n7485), .Z(n7483) );
  XOR U7283 ( .A(n7486), .B(n7484), .Z(n7485) );
  NANDN U7284 ( .A(n7445), .B(n7447), .Z(n7461) );
  XOR U7285 ( .A(n7487), .B(n7488), .Z(n7447) );
  AND U7286 ( .A(n438), .B(n7489), .Z(n7487) );
  XOR U7287 ( .A(n7488), .B(n7490), .Z(n7489) );
  XOR U7288 ( .A(n7491), .B(n7492), .Z(n438) );
  AND U7289 ( .A(n7493), .B(n7494), .Z(n7491) );
  XNOR U7290 ( .A(n7492), .B(n7458), .Z(n7494) );
  XNOR U7291 ( .A(n7495), .B(n7496), .Z(n7458) );
  ANDN U7292 ( .B(n7497), .A(n7498), .Z(n7495) );
  XOR U7293 ( .A(n7496), .B(n7499), .Z(n7497) );
  XOR U7294 ( .A(n7492), .B(n7460), .Z(n7493) );
  XOR U7295 ( .A(n7500), .B(n7501), .Z(n7460) );
  AND U7296 ( .A(n442), .B(n7502), .Z(n7500) );
  XOR U7297 ( .A(n7503), .B(n7501), .Z(n7502) );
  XNOR U7298 ( .A(n7504), .B(n7505), .Z(n7492) );
  NAND U7299 ( .A(n7506), .B(n7507), .Z(n7505) );
  XOR U7300 ( .A(n7508), .B(n7484), .Z(n7507) );
  XOR U7301 ( .A(n7498), .B(n7499), .Z(n7484) );
  XOR U7302 ( .A(n7509), .B(n7510), .Z(n7499) );
  ANDN U7303 ( .B(n7511), .A(n7512), .Z(n7509) );
  XOR U7304 ( .A(n7510), .B(n7513), .Z(n7511) );
  XOR U7305 ( .A(n7514), .B(n7515), .Z(n7498) );
  XOR U7306 ( .A(n7516), .B(n7517), .Z(n7515) );
  ANDN U7307 ( .B(n7518), .A(n7519), .Z(n7516) );
  XOR U7308 ( .A(n7520), .B(n7517), .Z(n7518) );
  IV U7309 ( .A(n7496), .Z(n7514) );
  XOR U7310 ( .A(n7521), .B(n7522), .Z(n7496) );
  ANDN U7311 ( .B(n7523), .A(n7524), .Z(n7521) );
  XOR U7312 ( .A(n7522), .B(n7525), .Z(n7523) );
  IV U7313 ( .A(n7504), .Z(n7508) );
  XOR U7314 ( .A(n7504), .B(n7486), .Z(n7506) );
  XOR U7315 ( .A(n7526), .B(n7527), .Z(n7486) );
  AND U7316 ( .A(n442), .B(n7528), .Z(n7526) );
  XOR U7317 ( .A(n7529), .B(n7527), .Z(n7528) );
  NANDN U7318 ( .A(n7488), .B(n7490), .Z(n7504) );
  XOR U7319 ( .A(n7530), .B(n7531), .Z(n7490) );
  AND U7320 ( .A(n442), .B(n7532), .Z(n7530) );
  XOR U7321 ( .A(n7531), .B(n7533), .Z(n7532) );
  XOR U7322 ( .A(n7534), .B(n7535), .Z(n442) );
  AND U7323 ( .A(n7536), .B(n7537), .Z(n7534) );
  XNOR U7324 ( .A(n7535), .B(n7501), .Z(n7537) );
  XNOR U7325 ( .A(n7538), .B(n7539), .Z(n7501) );
  ANDN U7326 ( .B(n7540), .A(n7541), .Z(n7538) );
  XOR U7327 ( .A(n7539), .B(n7542), .Z(n7540) );
  XOR U7328 ( .A(n7535), .B(n7503), .Z(n7536) );
  XOR U7329 ( .A(n7543), .B(n7544), .Z(n7503) );
  AND U7330 ( .A(n446), .B(n7545), .Z(n7543) );
  XOR U7331 ( .A(n7546), .B(n7544), .Z(n7545) );
  XNOR U7332 ( .A(n7547), .B(n7548), .Z(n7535) );
  NAND U7333 ( .A(n7549), .B(n7550), .Z(n7548) );
  XOR U7334 ( .A(n7551), .B(n7527), .Z(n7550) );
  XOR U7335 ( .A(n7541), .B(n7542), .Z(n7527) );
  XOR U7336 ( .A(n7552), .B(n7553), .Z(n7542) );
  ANDN U7337 ( .B(n7554), .A(n7555), .Z(n7552) );
  XOR U7338 ( .A(n7553), .B(n7556), .Z(n7554) );
  XOR U7339 ( .A(n7557), .B(n7558), .Z(n7541) );
  XOR U7340 ( .A(n7559), .B(n7560), .Z(n7558) );
  ANDN U7341 ( .B(n7561), .A(n7562), .Z(n7559) );
  XOR U7342 ( .A(n7563), .B(n7560), .Z(n7561) );
  IV U7343 ( .A(n7539), .Z(n7557) );
  XOR U7344 ( .A(n7564), .B(n7565), .Z(n7539) );
  ANDN U7345 ( .B(n7566), .A(n7567), .Z(n7564) );
  XOR U7346 ( .A(n7565), .B(n7568), .Z(n7566) );
  IV U7347 ( .A(n7547), .Z(n7551) );
  XOR U7348 ( .A(n7547), .B(n7529), .Z(n7549) );
  XOR U7349 ( .A(n7569), .B(n7570), .Z(n7529) );
  AND U7350 ( .A(n446), .B(n7571), .Z(n7569) );
  XOR U7351 ( .A(n7572), .B(n7570), .Z(n7571) );
  NANDN U7352 ( .A(n7531), .B(n7533), .Z(n7547) );
  XOR U7353 ( .A(n7573), .B(n7574), .Z(n7533) );
  AND U7354 ( .A(n446), .B(n7575), .Z(n7573) );
  XOR U7355 ( .A(n7574), .B(n7576), .Z(n7575) );
  XOR U7356 ( .A(n7577), .B(n7578), .Z(n446) );
  AND U7357 ( .A(n7579), .B(n7580), .Z(n7577) );
  XNOR U7358 ( .A(n7578), .B(n7544), .Z(n7580) );
  XNOR U7359 ( .A(n7581), .B(n7582), .Z(n7544) );
  ANDN U7360 ( .B(n7583), .A(n7584), .Z(n7581) );
  XOR U7361 ( .A(n7582), .B(n7585), .Z(n7583) );
  XOR U7362 ( .A(n7578), .B(n7546), .Z(n7579) );
  XOR U7363 ( .A(n7586), .B(n7587), .Z(n7546) );
  AND U7364 ( .A(n450), .B(n7588), .Z(n7586) );
  XOR U7365 ( .A(n7589), .B(n7587), .Z(n7588) );
  XNOR U7366 ( .A(n7590), .B(n7591), .Z(n7578) );
  NAND U7367 ( .A(n7592), .B(n7593), .Z(n7591) );
  XOR U7368 ( .A(n7594), .B(n7570), .Z(n7593) );
  XOR U7369 ( .A(n7584), .B(n7585), .Z(n7570) );
  XOR U7370 ( .A(n7595), .B(n7596), .Z(n7585) );
  ANDN U7371 ( .B(n7597), .A(n7598), .Z(n7595) );
  XOR U7372 ( .A(n7596), .B(n7599), .Z(n7597) );
  XOR U7373 ( .A(n7600), .B(n7601), .Z(n7584) );
  XOR U7374 ( .A(n7602), .B(n7603), .Z(n7601) );
  ANDN U7375 ( .B(n7604), .A(n7605), .Z(n7602) );
  XOR U7376 ( .A(n7606), .B(n7603), .Z(n7604) );
  IV U7377 ( .A(n7582), .Z(n7600) );
  XOR U7378 ( .A(n7607), .B(n7608), .Z(n7582) );
  ANDN U7379 ( .B(n7609), .A(n7610), .Z(n7607) );
  XOR U7380 ( .A(n7608), .B(n7611), .Z(n7609) );
  IV U7381 ( .A(n7590), .Z(n7594) );
  XOR U7382 ( .A(n7590), .B(n7572), .Z(n7592) );
  XOR U7383 ( .A(n7612), .B(n7613), .Z(n7572) );
  AND U7384 ( .A(n450), .B(n7614), .Z(n7612) );
  XOR U7385 ( .A(n7615), .B(n7613), .Z(n7614) );
  NANDN U7386 ( .A(n7574), .B(n7576), .Z(n7590) );
  XOR U7387 ( .A(n7616), .B(n7617), .Z(n7576) );
  AND U7388 ( .A(n450), .B(n7618), .Z(n7616) );
  XOR U7389 ( .A(n7617), .B(n7619), .Z(n7618) );
  XOR U7390 ( .A(n7620), .B(n7621), .Z(n450) );
  AND U7391 ( .A(n7622), .B(n7623), .Z(n7620) );
  XNOR U7392 ( .A(n7621), .B(n7587), .Z(n7623) );
  XNOR U7393 ( .A(n7624), .B(n7625), .Z(n7587) );
  ANDN U7394 ( .B(n7626), .A(n7627), .Z(n7624) );
  XOR U7395 ( .A(n7625), .B(n7628), .Z(n7626) );
  XOR U7396 ( .A(n7621), .B(n7589), .Z(n7622) );
  XOR U7397 ( .A(n7629), .B(n7630), .Z(n7589) );
  AND U7398 ( .A(n454), .B(n7631), .Z(n7629) );
  XOR U7399 ( .A(n7632), .B(n7630), .Z(n7631) );
  XNOR U7400 ( .A(n7633), .B(n7634), .Z(n7621) );
  NAND U7401 ( .A(n7635), .B(n7636), .Z(n7634) );
  XOR U7402 ( .A(n7637), .B(n7613), .Z(n7636) );
  XOR U7403 ( .A(n7627), .B(n7628), .Z(n7613) );
  XOR U7404 ( .A(n7638), .B(n7639), .Z(n7628) );
  ANDN U7405 ( .B(n7640), .A(n7641), .Z(n7638) );
  XOR U7406 ( .A(n7639), .B(n7642), .Z(n7640) );
  XOR U7407 ( .A(n7643), .B(n7644), .Z(n7627) );
  XOR U7408 ( .A(n7645), .B(n7646), .Z(n7644) );
  ANDN U7409 ( .B(n7647), .A(n7648), .Z(n7645) );
  XOR U7410 ( .A(n7649), .B(n7646), .Z(n7647) );
  IV U7411 ( .A(n7625), .Z(n7643) );
  XOR U7412 ( .A(n7650), .B(n7651), .Z(n7625) );
  ANDN U7413 ( .B(n7652), .A(n7653), .Z(n7650) );
  XOR U7414 ( .A(n7651), .B(n7654), .Z(n7652) );
  IV U7415 ( .A(n7633), .Z(n7637) );
  XOR U7416 ( .A(n7633), .B(n7615), .Z(n7635) );
  XOR U7417 ( .A(n7655), .B(n7656), .Z(n7615) );
  AND U7418 ( .A(n454), .B(n7657), .Z(n7655) );
  XOR U7419 ( .A(n7658), .B(n7656), .Z(n7657) );
  NANDN U7420 ( .A(n7617), .B(n7619), .Z(n7633) );
  XOR U7421 ( .A(n7659), .B(n7660), .Z(n7619) );
  AND U7422 ( .A(n454), .B(n7661), .Z(n7659) );
  XOR U7423 ( .A(n7660), .B(n7662), .Z(n7661) );
  XOR U7424 ( .A(n7663), .B(n7664), .Z(n454) );
  AND U7425 ( .A(n7665), .B(n7666), .Z(n7663) );
  XNOR U7426 ( .A(n7664), .B(n7630), .Z(n7666) );
  XNOR U7427 ( .A(n7667), .B(n7668), .Z(n7630) );
  ANDN U7428 ( .B(n7669), .A(n7670), .Z(n7667) );
  XOR U7429 ( .A(n7668), .B(n7671), .Z(n7669) );
  XOR U7430 ( .A(n7664), .B(n7632), .Z(n7665) );
  XOR U7431 ( .A(n7672), .B(n7673), .Z(n7632) );
  AND U7432 ( .A(n458), .B(n7674), .Z(n7672) );
  XOR U7433 ( .A(n7675), .B(n7673), .Z(n7674) );
  XNOR U7434 ( .A(n7676), .B(n7677), .Z(n7664) );
  NAND U7435 ( .A(n7678), .B(n7679), .Z(n7677) );
  XOR U7436 ( .A(n7680), .B(n7656), .Z(n7679) );
  XOR U7437 ( .A(n7670), .B(n7671), .Z(n7656) );
  XOR U7438 ( .A(n7681), .B(n7682), .Z(n7671) );
  ANDN U7439 ( .B(n7683), .A(n7684), .Z(n7681) );
  XOR U7440 ( .A(n7682), .B(n7685), .Z(n7683) );
  XOR U7441 ( .A(n7686), .B(n7687), .Z(n7670) );
  XOR U7442 ( .A(n7688), .B(n7689), .Z(n7687) );
  ANDN U7443 ( .B(n7690), .A(n7691), .Z(n7688) );
  XOR U7444 ( .A(n7692), .B(n7689), .Z(n7690) );
  IV U7445 ( .A(n7668), .Z(n7686) );
  XOR U7446 ( .A(n7693), .B(n7694), .Z(n7668) );
  ANDN U7447 ( .B(n7695), .A(n7696), .Z(n7693) );
  XOR U7448 ( .A(n7694), .B(n7697), .Z(n7695) );
  IV U7449 ( .A(n7676), .Z(n7680) );
  XOR U7450 ( .A(n7676), .B(n7658), .Z(n7678) );
  XOR U7451 ( .A(n7698), .B(n7699), .Z(n7658) );
  AND U7452 ( .A(n458), .B(n7700), .Z(n7698) );
  XOR U7453 ( .A(n7701), .B(n7699), .Z(n7700) );
  NANDN U7454 ( .A(n7660), .B(n7662), .Z(n7676) );
  XOR U7455 ( .A(n7702), .B(n7703), .Z(n7662) );
  AND U7456 ( .A(n458), .B(n7704), .Z(n7702) );
  XOR U7457 ( .A(n7703), .B(n7705), .Z(n7704) );
  XOR U7458 ( .A(n7706), .B(n7707), .Z(n458) );
  AND U7459 ( .A(n7708), .B(n7709), .Z(n7706) );
  XNOR U7460 ( .A(n7707), .B(n7673), .Z(n7709) );
  XNOR U7461 ( .A(n7710), .B(n7711), .Z(n7673) );
  ANDN U7462 ( .B(n7712), .A(n7713), .Z(n7710) );
  XOR U7463 ( .A(n7711), .B(n7714), .Z(n7712) );
  XOR U7464 ( .A(n7707), .B(n7675), .Z(n7708) );
  XOR U7465 ( .A(n7715), .B(n7716), .Z(n7675) );
  AND U7466 ( .A(n462), .B(n7717), .Z(n7715) );
  XOR U7467 ( .A(n7718), .B(n7716), .Z(n7717) );
  XNOR U7468 ( .A(n7719), .B(n7720), .Z(n7707) );
  NAND U7469 ( .A(n7721), .B(n7722), .Z(n7720) );
  XOR U7470 ( .A(n7723), .B(n7699), .Z(n7722) );
  XOR U7471 ( .A(n7713), .B(n7714), .Z(n7699) );
  XOR U7472 ( .A(n7724), .B(n7725), .Z(n7714) );
  ANDN U7473 ( .B(n7726), .A(n7727), .Z(n7724) );
  XOR U7474 ( .A(n7725), .B(n7728), .Z(n7726) );
  XOR U7475 ( .A(n7729), .B(n7730), .Z(n7713) );
  XOR U7476 ( .A(n7731), .B(n7732), .Z(n7730) );
  ANDN U7477 ( .B(n7733), .A(n7734), .Z(n7731) );
  XOR U7478 ( .A(n7735), .B(n7732), .Z(n7733) );
  IV U7479 ( .A(n7711), .Z(n7729) );
  XOR U7480 ( .A(n7736), .B(n7737), .Z(n7711) );
  ANDN U7481 ( .B(n7738), .A(n7739), .Z(n7736) );
  XOR U7482 ( .A(n7737), .B(n7740), .Z(n7738) );
  IV U7483 ( .A(n7719), .Z(n7723) );
  XOR U7484 ( .A(n7719), .B(n7701), .Z(n7721) );
  XOR U7485 ( .A(n7741), .B(n7742), .Z(n7701) );
  AND U7486 ( .A(n462), .B(n7743), .Z(n7741) );
  XOR U7487 ( .A(n7744), .B(n7742), .Z(n7743) );
  NANDN U7488 ( .A(n7703), .B(n7705), .Z(n7719) );
  XOR U7489 ( .A(n7745), .B(n7746), .Z(n7705) );
  AND U7490 ( .A(n462), .B(n7747), .Z(n7745) );
  XOR U7491 ( .A(n7746), .B(n7748), .Z(n7747) );
  XOR U7492 ( .A(n7749), .B(n7750), .Z(n462) );
  AND U7493 ( .A(n7751), .B(n7752), .Z(n7749) );
  XNOR U7494 ( .A(n7750), .B(n7716), .Z(n7752) );
  XNOR U7495 ( .A(n7753), .B(n7754), .Z(n7716) );
  ANDN U7496 ( .B(n7755), .A(n7756), .Z(n7753) );
  XOR U7497 ( .A(n7754), .B(n7757), .Z(n7755) );
  XOR U7498 ( .A(n7750), .B(n7718), .Z(n7751) );
  XOR U7499 ( .A(n7758), .B(n7759), .Z(n7718) );
  AND U7500 ( .A(n466), .B(n7760), .Z(n7758) );
  XOR U7501 ( .A(n7761), .B(n7759), .Z(n7760) );
  XNOR U7502 ( .A(n7762), .B(n7763), .Z(n7750) );
  NAND U7503 ( .A(n7764), .B(n7765), .Z(n7763) );
  XOR U7504 ( .A(n7766), .B(n7742), .Z(n7765) );
  XOR U7505 ( .A(n7756), .B(n7757), .Z(n7742) );
  XOR U7506 ( .A(n7767), .B(n7768), .Z(n7757) );
  ANDN U7507 ( .B(n7769), .A(n7770), .Z(n7767) );
  XOR U7508 ( .A(n7768), .B(n7771), .Z(n7769) );
  XOR U7509 ( .A(n7772), .B(n7773), .Z(n7756) );
  XOR U7510 ( .A(n7774), .B(n7775), .Z(n7773) );
  ANDN U7511 ( .B(n7776), .A(n7777), .Z(n7774) );
  XOR U7512 ( .A(n7778), .B(n7775), .Z(n7776) );
  IV U7513 ( .A(n7754), .Z(n7772) );
  XOR U7514 ( .A(n7779), .B(n7780), .Z(n7754) );
  ANDN U7515 ( .B(n7781), .A(n7782), .Z(n7779) );
  XOR U7516 ( .A(n7780), .B(n7783), .Z(n7781) );
  IV U7517 ( .A(n7762), .Z(n7766) );
  XOR U7518 ( .A(n7762), .B(n7744), .Z(n7764) );
  XOR U7519 ( .A(n7784), .B(n7785), .Z(n7744) );
  AND U7520 ( .A(n466), .B(n7786), .Z(n7784) );
  XOR U7521 ( .A(n7787), .B(n7785), .Z(n7786) );
  NANDN U7522 ( .A(n7746), .B(n7748), .Z(n7762) );
  XOR U7523 ( .A(n7788), .B(n7789), .Z(n7748) );
  AND U7524 ( .A(n466), .B(n7790), .Z(n7788) );
  XOR U7525 ( .A(n7789), .B(n7791), .Z(n7790) );
  XOR U7526 ( .A(n7792), .B(n7793), .Z(n466) );
  AND U7527 ( .A(n7794), .B(n7795), .Z(n7792) );
  XNOR U7528 ( .A(n7793), .B(n7759), .Z(n7795) );
  XNOR U7529 ( .A(n7796), .B(n7797), .Z(n7759) );
  ANDN U7530 ( .B(n7798), .A(n7799), .Z(n7796) );
  XOR U7531 ( .A(n7797), .B(n7800), .Z(n7798) );
  XOR U7532 ( .A(n7793), .B(n7761), .Z(n7794) );
  XOR U7533 ( .A(n7801), .B(n7802), .Z(n7761) );
  AND U7534 ( .A(n470), .B(n7803), .Z(n7801) );
  XOR U7535 ( .A(n7804), .B(n7802), .Z(n7803) );
  XNOR U7536 ( .A(n7805), .B(n7806), .Z(n7793) );
  NAND U7537 ( .A(n7807), .B(n7808), .Z(n7806) );
  XOR U7538 ( .A(n7809), .B(n7785), .Z(n7808) );
  XOR U7539 ( .A(n7799), .B(n7800), .Z(n7785) );
  XOR U7540 ( .A(n7810), .B(n7811), .Z(n7800) );
  ANDN U7541 ( .B(n7812), .A(n7813), .Z(n7810) );
  XOR U7542 ( .A(n7811), .B(n7814), .Z(n7812) );
  XOR U7543 ( .A(n7815), .B(n7816), .Z(n7799) );
  XOR U7544 ( .A(n7817), .B(n7818), .Z(n7816) );
  ANDN U7545 ( .B(n7819), .A(n7820), .Z(n7817) );
  XOR U7546 ( .A(n7821), .B(n7818), .Z(n7819) );
  IV U7547 ( .A(n7797), .Z(n7815) );
  XOR U7548 ( .A(n7822), .B(n7823), .Z(n7797) );
  ANDN U7549 ( .B(n7824), .A(n7825), .Z(n7822) );
  XOR U7550 ( .A(n7823), .B(n7826), .Z(n7824) );
  IV U7551 ( .A(n7805), .Z(n7809) );
  XOR U7552 ( .A(n7805), .B(n7787), .Z(n7807) );
  XOR U7553 ( .A(n7827), .B(n7828), .Z(n7787) );
  AND U7554 ( .A(n470), .B(n7829), .Z(n7827) );
  XOR U7555 ( .A(n7830), .B(n7828), .Z(n7829) );
  NANDN U7556 ( .A(n7789), .B(n7791), .Z(n7805) );
  XOR U7557 ( .A(n7831), .B(n7832), .Z(n7791) );
  AND U7558 ( .A(n470), .B(n7833), .Z(n7831) );
  XOR U7559 ( .A(n7832), .B(n7834), .Z(n7833) );
  XOR U7560 ( .A(n7835), .B(n7836), .Z(n470) );
  AND U7561 ( .A(n7837), .B(n7838), .Z(n7835) );
  XNOR U7562 ( .A(n7836), .B(n7802), .Z(n7838) );
  XNOR U7563 ( .A(n7839), .B(n7840), .Z(n7802) );
  ANDN U7564 ( .B(n7841), .A(n7842), .Z(n7839) );
  XOR U7565 ( .A(n7840), .B(n7843), .Z(n7841) );
  XOR U7566 ( .A(n7836), .B(n7804), .Z(n7837) );
  XOR U7567 ( .A(n7844), .B(n7845), .Z(n7804) );
  AND U7568 ( .A(n474), .B(n7846), .Z(n7844) );
  XOR U7569 ( .A(n7847), .B(n7845), .Z(n7846) );
  XNOR U7570 ( .A(n7848), .B(n7849), .Z(n7836) );
  NAND U7571 ( .A(n7850), .B(n7851), .Z(n7849) );
  XOR U7572 ( .A(n7852), .B(n7828), .Z(n7851) );
  XOR U7573 ( .A(n7842), .B(n7843), .Z(n7828) );
  XOR U7574 ( .A(n7853), .B(n7854), .Z(n7843) );
  ANDN U7575 ( .B(n7855), .A(n7856), .Z(n7853) );
  XOR U7576 ( .A(n7854), .B(n7857), .Z(n7855) );
  XOR U7577 ( .A(n7858), .B(n7859), .Z(n7842) );
  XOR U7578 ( .A(n7860), .B(n7861), .Z(n7859) );
  ANDN U7579 ( .B(n7862), .A(n7863), .Z(n7860) );
  XOR U7580 ( .A(n7864), .B(n7861), .Z(n7862) );
  IV U7581 ( .A(n7840), .Z(n7858) );
  XOR U7582 ( .A(n7865), .B(n7866), .Z(n7840) );
  ANDN U7583 ( .B(n7867), .A(n7868), .Z(n7865) );
  XOR U7584 ( .A(n7866), .B(n7869), .Z(n7867) );
  IV U7585 ( .A(n7848), .Z(n7852) );
  XOR U7586 ( .A(n7848), .B(n7830), .Z(n7850) );
  XOR U7587 ( .A(n7870), .B(n7871), .Z(n7830) );
  AND U7588 ( .A(n474), .B(n7872), .Z(n7870) );
  XOR U7589 ( .A(n7873), .B(n7871), .Z(n7872) );
  NANDN U7590 ( .A(n7832), .B(n7834), .Z(n7848) );
  XOR U7591 ( .A(n7874), .B(n7875), .Z(n7834) );
  AND U7592 ( .A(n474), .B(n7876), .Z(n7874) );
  XOR U7593 ( .A(n7875), .B(n7877), .Z(n7876) );
  XOR U7594 ( .A(n7878), .B(n7879), .Z(n474) );
  AND U7595 ( .A(n7880), .B(n7881), .Z(n7878) );
  XNOR U7596 ( .A(n7879), .B(n7845), .Z(n7881) );
  XNOR U7597 ( .A(n7882), .B(n7883), .Z(n7845) );
  ANDN U7598 ( .B(n7884), .A(n7885), .Z(n7882) );
  XOR U7599 ( .A(n7883), .B(n7886), .Z(n7884) );
  XOR U7600 ( .A(n7879), .B(n7847), .Z(n7880) );
  XOR U7601 ( .A(n7887), .B(n7888), .Z(n7847) );
  AND U7602 ( .A(n478), .B(n7889), .Z(n7887) );
  XOR U7603 ( .A(n7890), .B(n7888), .Z(n7889) );
  XNOR U7604 ( .A(n7891), .B(n7892), .Z(n7879) );
  NAND U7605 ( .A(n7893), .B(n7894), .Z(n7892) );
  XOR U7606 ( .A(n7895), .B(n7871), .Z(n7894) );
  XOR U7607 ( .A(n7885), .B(n7886), .Z(n7871) );
  XOR U7608 ( .A(n7896), .B(n7897), .Z(n7886) );
  ANDN U7609 ( .B(n7898), .A(n7899), .Z(n7896) );
  XOR U7610 ( .A(n7897), .B(n7900), .Z(n7898) );
  XOR U7611 ( .A(n7901), .B(n7902), .Z(n7885) );
  XOR U7612 ( .A(n7903), .B(n7904), .Z(n7902) );
  ANDN U7613 ( .B(n7905), .A(n7906), .Z(n7903) );
  XOR U7614 ( .A(n7907), .B(n7904), .Z(n7905) );
  IV U7615 ( .A(n7883), .Z(n7901) );
  XOR U7616 ( .A(n7908), .B(n7909), .Z(n7883) );
  ANDN U7617 ( .B(n7910), .A(n7911), .Z(n7908) );
  XOR U7618 ( .A(n7909), .B(n7912), .Z(n7910) );
  IV U7619 ( .A(n7891), .Z(n7895) );
  XOR U7620 ( .A(n7891), .B(n7873), .Z(n7893) );
  XOR U7621 ( .A(n7913), .B(n7914), .Z(n7873) );
  AND U7622 ( .A(n478), .B(n7915), .Z(n7913) );
  XOR U7623 ( .A(n7916), .B(n7914), .Z(n7915) );
  NANDN U7624 ( .A(n7875), .B(n7877), .Z(n7891) );
  XOR U7625 ( .A(n7917), .B(n7918), .Z(n7877) );
  AND U7626 ( .A(n478), .B(n7919), .Z(n7917) );
  XOR U7627 ( .A(n7918), .B(n7920), .Z(n7919) );
  XOR U7628 ( .A(n7921), .B(n7922), .Z(n478) );
  AND U7629 ( .A(n7923), .B(n7924), .Z(n7921) );
  XNOR U7630 ( .A(n7922), .B(n7888), .Z(n7924) );
  XNOR U7631 ( .A(n7925), .B(n7926), .Z(n7888) );
  ANDN U7632 ( .B(n7927), .A(n7928), .Z(n7925) );
  XOR U7633 ( .A(n7926), .B(n7929), .Z(n7927) );
  XOR U7634 ( .A(n7922), .B(n7890), .Z(n7923) );
  XOR U7635 ( .A(n7930), .B(n7931), .Z(n7890) );
  AND U7636 ( .A(n482), .B(n7932), .Z(n7930) );
  XOR U7637 ( .A(n7933), .B(n7931), .Z(n7932) );
  XNOR U7638 ( .A(n7934), .B(n7935), .Z(n7922) );
  NAND U7639 ( .A(n7936), .B(n7937), .Z(n7935) );
  XOR U7640 ( .A(n7938), .B(n7914), .Z(n7937) );
  XOR U7641 ( .A(n7928), .B(n7929), .Z(n7914) );
  XOR U7642 ( .A(n7939), .B(n7940), .Z(n7929) );
  ANDN U7643 ( .B(n7941), .A(n7942), .Z(n7939) );
  XOR U7644 ( .A(n7940), .B(n7943), .Z(n7941) );
  XOR U7645 ( .A(n7944), .B(n7945), .Z(n7928) );
  XOR U7646 ( .A(n7946), .B(n7947), .Z(n7945) );
  ANDN U7647 ( .B(n7948), .A(n7949), .Z(n7946) );
  XOR U7648 ( .A(n7950), .B(n7947), .Z(n7948) );
  IV U7649 ( .A(n7926), .Z(n7944) );
  XOR U7650 ( .A(n7951), .B(n7952), .Z(n7926) );
  ANDN U7651 ( .B(n7953), .A(n7954), .Z(n7951) );
  XOR U7652 ( .A(n7952), .B(n7955), .Z(n7953) );
  IV U7653 ( .A(n7934), .Z(n7938) );
  XOR U7654 ( .A(n7934), .B(n7916), .Z(n7936) );
  XOR U7655 ( .A(n7956), .B(n7957), .Z(n7916) );
  AND U7656 ( .A(n482), .B(n7958), .Z(n7956) );
  XOR U7657 ( .A(n7959), .B(n7957), .Z(n7958) );
  NANDN U7658 ( .A(n7918), .B(n7920), .Z(n7934) );
  XOR U7659 ( .A(n7960), .B(n7961), .Z(n7920) );
  AND U7660 ( .A(n482), .B(n7962), .Z(n7960) );
  XOR U7661 ( .A(n7961), .B(n7963), .Z(n7962) );
  XOR U7662 ( .A(n7964), .B(n7965), .Z(n482) );
  AND U7663 ( .A(n7966), .B(n7967), .Z(n7964) );
  XNOR U7664 ( .A(n7965), .B(n7931), .Z(n7967) );
  XNOR U7665 ( .A(n7968), .B(n7969), .Z(n7931) );
  ANDN U7666 ( .B(n7970), .A(n7971), .Z(n7968) );
  XOR U7667 ( .A(n7969), .B(n7972), .Z(n7970) );
  XOR U7668 ( .A(n7965), .B(n7933), .Z(n7966) );
  XOR U7669 ( .A(n7973), .B(n7974), .Z(n7933) );
  AND U7670 ( .A(n486), .B(n7975), .Z(n7973) );
  XOR U7671 ( .A(n7976), .B(n7974), .Z(n7975) );
  XNOR U7672 ( .A(n7977), .B(n7978), .Z(n7965) );
  NAND U7673 ( .A(n7979), .B(n7980), .Z(n7978) );
  XOR U7674 ( .A(n7981), .B(n7957), .Z(n7980) );
  XOR U7675 ( .A(n7971), .B(n7972), .Z(n7957) );
  XOR U7676 ( .A(n7982), .B(n7983), .Z(n7972) );
  ANDN U7677 ( .B(n7984), .A(n7985), .Z(n7982) );
  XOR U7678 ( .A(n7983), .B(n7986), .Z(n7984) );
  XOR U7679 ( .A(n7987), .B(n7988), .Z(n7971) );
  XOR U7680 ( .A(n7989), .B(n7990), .Z(n7988) );
  ANDN U7681 ( .B(n7991), .A(n7992), .Z(n7989) );
  XOR U7682 ( .A(n7993), .B(n7990), .Z(n7991) );
  IV U7683 ( .A(n7969), .Z(n7987) );
  XOR U7684 ( .A(n7994), .B(n7995), .Z(n7969) );
  ANDN U7685 ( .B(n7996), .A(n7997), .Z(n7994) );
  XOR U7686 ( .A(n7995), .B(n7998), .Z(n7996) );
  IV U7687 ( .A(n7977), .Z(n7981) );
  XOR U7688 ( .A(n7977), .B(n7959), .Z(n7979) );
  XOR U7689 ( .A(n7999), .B(n8000), .Z(n7959) );
  AND U7690 ( .A(n486), .B(n8001), .Z(n7999) );
  XOR U7691 ( .A(n8002), .B(n8000), .Z(n8001) );
  NANDN U7692 ( .A(n7961), .B(n7963), .Z(n7977) );
  XOR U7693 ( .A(n8003), .B(n8004), .Z(n7963) );
  AND U7694 ( .A(n486), .B(n8005), .Z(n8003) );
  XOR U7695 ( .A(n8004), .B(n8006), .Z(n8005) );
  XOR U7696 ( .A(n8007), .B(n8008), .Z(n486) );
  AND U7697 ( .A(n8009), .B(n8010), .Z(n8007) );
  XNOR U7698 ( .A(n8008), .B(n7974), .Z(n8010) );
  XNOR U7699 ( .A(n8011), .B(n8012), .Z(n7974) );
  ANDN U7700 ( .B(n8013), .A(n8014), .Z(n8011) );
  XOR U7701 ( .A(n8012), .B(n8015), .Z(n8013) );
  XOR U7702 ( .A(n8008), .B(n7976), .Z(n8009) );
  XOR U7703 ( .A(n8016), .B(n8017), .Z(n7976) );
  AND U7704 ( .A(n490), .B(n8018), .Z(n8016) );
  XOR U7705 ( .A(n8019), .B(n8017), .Z(n8018) );
  XNOR U7706 ( .A(n8020), .B(n8021), .Z(n8008) );
  NAND U7707 ( .A(n8022), .B(n8023), .Z(n8021) );
  XOR U7708 ( .A(n8024), .B(n8000), .Z(n8023) );
  XOR U7709 ( .A(n8014), .B(n8015), .Z(n8000) );
  XOR U7710 ( .A(n8025), .B(n8026), .Z(n8015) );
  ANDN U7711 ( .B(n8027), .A(n8028), .Z(n8025) );
  XOR U7712 ( .A(n8026), .B(n8029), .Z(n8027) );
  XOR U7713 ( .A(n8030), .B(n8031), .Z(n8014) );
  XOR U7714 ( .A(n8032), .B(n8033), .Z(n8031) );
  ANDN U7715 ( .B(n8034), .A(n8035), .Z(n8032) );
  XOR U7716 ( .A(n8036), .B(n8033), .Z(n8034) );
  IV U7717 ( .A(n8012), .Z(n8030) );
  XOR U7718 ( .A(n8037), .B(n8038), .Z(n8012) );
  ANDN U7719 ( .B(n8039), .A(n8040), .Z(n8037) );
  XOR U7720 ( .A(n8038), .B(n8041), .Z(n8039) );
  IV U7721 ( .A(n8020), .Z(n8024) );
  XOR U7722 ( .A(n8020), .B(n8002), .Z(n8022) );
  XOR U7723 ( .A(n8042), .B(n8043), .Z(n8002) );
  AND U7724 ( .A(n490), .B(n8044), .Z(n8042) );
  XOR U7725 ( .A(n8045), .B(n8043), .Z(n8044) );
  NANDN U7726 ( .A(n8004), .B(n8006), .Z(n8020) );
  XOR U7727 ( .A(n8046), .B(n8047), .Z(n8006) );
  AND U7728 ( .A(n490), .B(n8048), .Z(n8046) );
  XOR U7729 ( .A(n8047), .B(n8049), .Z(n8048) );
  XOR U7730 ( .A(n8050), .B(n8051), .Z(n490) );
  AND U7731 ( .A(n8052), .B(n8053), .Z(n8050) );
  XNOR U7732 ( .A(n8051), .B(n8017), .Z(n8053) );
  XNOR U7733 ( .A(n8054), .B(n8055), .Z(n8017) );
  ANDN U7734 ( .B(n8056), .A(n8057), .Z(n8054) );
  XOR U7735 ( .A(n8055), .B(n8058), .Z(n8056) );
  XOR U7736 ( .A(n8051), .B(n8019), .Z(n8052) );
  XOR U7737 ( .A(n8059), .B(n8060), .Z(n8019) );
  AND U7738 ( .A(n494), .B(n8061), .Z(n8059) );
  XOR U7739 ( .A(n8062), .B(n8060), .Z(n8061) );
  XNOR U7740 ( .A(n8063), .B(n8064), .Z(n8051) );
  NAND U7741 ( .A(n8065), .B(n8066), .Z(n8064) );
  XOR U7742 ( .A(n8067), .B(n8043), .Z(n8066) );
  XOR U7743 ( .A(n8057), .B(n8058), .Z(n8043) );
  XOR U7744 ( .A(n8068), .B(n8069), .Z(n8058) );
  ANDN U7745 ( .B(n8070), .A(n8071), .Z(n8068) );
  XOR U7746 ( .A(n8069), .B(n8072), .Z(n8070) );
  XOR U7747 ( .A(n8073), .B(n8074), .Z(n8057) );
  XOR U7748 ( .A(n8075), .B(n8076), .Z(n8074) );
  ANDN U7749 ( .B(n8077), .A(n8078), .Z(n8075) );
  XOR U7750 ( .A(n8079), .B(n8076), .Z(n8077) );
  IV U7751 ( .A(n8055), .Z(n8073) );
  XOR U7752 ( .A(n8080), .B(n8081), .Z(n8055) );
  ANDN U7753 ( .B(n8082), .A(n8083), .Z(n8080) );
  XOR U7754 ( .A(n8081), .B(n8084), .Z(n8082) );
  IV U7755 ( .A(n8063), .Z(n8067) );
  XOR U7756 ( .A(n8063), .B(n8045), .Z(n8065) );
  XOR U7757 ( .A(n8085), .B(n8086), .Z(n8045) );
  AND U7758 ( .A(n494), .B(n8087), .Z(n8085) );
  XOR U7759 ( .A(n8088), .B(n8086), .Z(n8087) );
  NANDN U7760 ( .A(n8047), .B(n8049), .Z(n8063) );
  XOR U7761 ( .A(n8089), .B(n8090), .Z(n8049) );
  AND U7762 ( .A(n494), .B(n8091), .Z(n8089) );
  XOR U7763 ( .A(n8090), .B(n8092), .Z(n8091) );
  XOR U7764 ( .A(n8093), .B(n8094), .Z(n494) );
  AND U7765 ( .A(n8095), .B(n8096), .Z(n8093) );
  XNOR U7766 ( .A(n8094), .B(n8060), .Z(n8096) );
  XNOR U7767 ( .A(n8097), .B(n8098), .Z(n8060) );
  ANDN U7768 ( .B(n8099), .A(n8100), .Z(n8097) );
  XOR U7769 ( .A(n8098), .B(n8101), .Z(n8099) );
  XOR U7770 ( .A(n8094), .B(n8062), .Z(n8095) );
  XOR U7771 ( .A(n8102), .B(n8103), .Z(n8062) );
  AND U7772 ( .A(n498), .B(n8104), .Z(n8102) );
  XOR U7773 ( .A(n8105), .B(n8103), .Z(n8104) );
  XNOR U7774 ( .A(n8106), .B(n8107), .Z(n8094) );
  NAND U7775 ( .A(n8108), .B(n8109), .Z(n8107) );
  XOR U7776 ( .A(n8110), .B(n8086), .Z(n8109) );
  XOR U7777 ( .A(n8100), .B(n8101), .Z(n8086) );
  XOR U7778 ( .A(n8111), .B(n8112), .Z(n8101) );
  ANDN U7779 ( .B(n8113), .A(n8114), .Z(n8111) );
  XOR U7780 ( .A(n8112), .B(n8115), .Z(n8113) );
  XOR U7781 ( .A(n8116), .B(n8117), .Z(n8100) );
  XOR U7782 ( .A(n8118), .B(n8119), .Z(n8117) );
  ANDN U7783 ( .B(n8120), .A(n8121), .Z(n8118) );
  XOR U7784 ( .A(n8122), .B(n8119), .Z(n8120) );
  IV U7785 ( .A(n8098), .Z(n8116) );
  XOR U7786 ( .A(n8123), .B(n8124), .Z(n8098) );
  ANDN U7787 ( .B(n8125), .A(n8126), .Z(n8123) );
  XOR U7788 ( .A(n8124), .B(n8127), .Z(n8125) );
  IV U7789 ( .A(n8106), .Z(n8110) );
  XOR U7790 ( .A(n8106), .B(n8088), .Z(n8108) );
  XOR U7791 ( .A(n8128), .B(n8129), .Z(n8088) );
  AND U7792 ( .A(n498), .B(n8130), .Z(n8128) );
  XOR U7793 ( .A(n8131), .B(n8129), .Z(n8130) );
  NANDN U7794 ( .A(n8090), .B(n8092), .Z(n8106) );
  XOR U7795 ( .A(n8132), .B(n8133), .Z(n8092) );
  AND U7796 ( .A(n498), .B(n8134), .Z(n8132) );
  XOR U7797 ( .A(n8133), .B(n8135), .Z(n8134) );
  XOR U7798 ( .A(n8136), .B(n8137), .Z(n498) );
  AND U7799 ( .A(n8138), .B(n8139), .Z(n8136) );
  XNOR U7800 ( .A(n8137), .B(n8103), .Z(n8139) );
  XNOR U7801 ( .A(n8140), .B(n8141), .Z(n8103) );
  ANDN U7802 ( .B(n8142), .A(n8143), .Z(n8140) );
  XOR U7803 ( .A(n8141), .B(n8144), .Z(n8142) );
  XOR U7804 ( .A(n8137), .B(n8105), .Z(n8138) );
  XOR U7805 ( .A(n8145), .B(n8146), .Z(n8105) );
  AND U7806 ( .A(n502), .B(n8147), .Z(n8145) );
  XOR U7807 ( .A(n8148), .B(n8146), .Z(n8147) );
  XNOR U7808 ( .A(n8149), .B(n8150), .Z(n8137) );
  NAND U7809 ( .A(n8151), .B(n8152), .Z(n8150) );
  XOR U7810 ( .A(n8153), .B(n8129), .Z(n8152) );
  XOR U7811 ( .A(n8143), .B(n8144), .Z(n8129) );
  XOR U7812 ( .A(n8154), .B(n8155), .Z(n8144) );
  ANDN U7813 ( .B(n8156), .A(n8157), .Z(n8154) );
  XOR U7814 ( .A(n8155), .B(n8158), .Z(n8156) );
  XOR U7815 ( .A(n8159), .B(n8160), .Z(n8143) );
  XOR U7816 ( .A(n8161), .B(n8162), .Z(n8160) );
  ANDN U7817 ( .B(n8163), .A(n8164), .Z(n8161) );
  XOR U7818 ( .A(n8165), .B(n8162), .Z(n8163) );
  IV U7819 ( .A(n8141), .Z(n8159) );
  XOR U7820 ( .A(n8166), .B(n8167), .Z(n8141) );
  ANDN U7821 ( .B(n8168), .A(n8169), .Z(n8166) );
  XOR U7822 ( .A(n8167), .B(n8170), .Z(n8168) );
  IV U7823 ( .A(n8149), .Z(n8153) );
  XOR U7824 ( .A(n8149), .B(n8131), .Z(n8151) );
  XOR U7825 ( .A(n8171), .B(n8172), .Z(n8131) );
  AND U7826 ( .A(n502), .B(n8173), .Z(n8171) );
  XOR U7827 ( .A(n8174), .B(n8172), .Z(n8173) );
  NANDN U7828 ( .A(n8133), .B(n8135), .Z(n8149) );
  XOR U7829 ( .A(n8175), .B(n8176), .Z(n8135) );
  AND U7830 ( .A(n502), .B(n8177), .Z(n8175) );
  XOR U7831 ( .A(n8176), .B(n8178), .Z(n8177) );
  XOR U7832 ( .A(n8179), .B(n8180), .Z(n502) );
  AND U7833 ( .A(n8181), .B(n8182), .Z(n8179) );
  XNOR U7834 ( .A(n8180), .B(n8146), .Z(n8182) );
  XNOR U7835 ( .A(n8183), .B(n8184), .Z(n8146) );
  ANDN U7836 ( .B(n8185), .A(n8186), .Z(n8183) );
  XOR U7837 ( .A(n8184), .B(n8187), .Z(n8185) );
  XOR U7838 ( .A(n8180), .B(n8148), .Z(n8181) );
  XOR U7839 ( .A(n8188), .B(n8189), .Z(n8148) );
  AND U7840 ( .A(n506), .B(n8190), .Z(n8188) );
  XOR U7841 ( .A(n8191), .B(n8189), .Z(n8190) );
  XNOR U7842 ( .A(n8192), .B(n8193), .Z(n8180) );
  NAND U7843 ( .A(n8194), .B(n8195), .Z(n8193) );
  XOR U7844 ( .A(n8196), .B(n8172), .Z(n8195) );
  XOR U7845 ( .A(n8186), .B(n8187), .Z(n8172) );
  XOR U7846 ( .A(n8197), .B(n8198), .Z(n8187) );
  ANDN U7847 ( .B(n8199), .A(n8200), .Z(n8197) );
  XOR U7848 ( .A(n8198), .B(n8201), .Z(n8199) );
  XOR U7849 ( .A(n8202), .B(n8203), .Z(n8186) );
  XOR U7850 ( .A(n8204), .B(n8205), .Z(n8203) );
  ANDN U7851 ( .B(n8206), .A(n8207), .Z(n8204) );
  XOR U7852 ( .A(n8208), .B(n8205), .Z(n8206) );
  IV U7853 ( .A(n8184), .Z(n8202) );
  XOR U7854 ( .A(n8209), .B(n8210), .Z(n8184) );
  ANDN U7855 ( .B(n8211), .A(n8212), .Z(n8209) );
  XOR U7856 ( .A(n8210), .B(n8213), .Z(n8211) );
  IV U7857 ( .A(n8192), .Z(n8196) );
  XOR U7858 ( .A(n8192), .B(n8174), .Z(n8194) );
  XOR U7859 ( .A(n8214), .B(n8215), .Z(n8174) );
  AND U7860 ( .A(n506), .B(n8216), .Z(n8214) );
  XNOR U7861 ( .A(n8217), .B(n8215), .Z(n8216) );
  NANDN U7862 ( .A(n8176), .B(n8178), .Z(n8192) );
  XOR U7863 ( .A(n8218), .B(n8219), .Z(n8178) );
  AND U7864 ( .A(n506), .B(n8220), .Z(n8218) );
  XOR U7865 ( .A(n8219), .B(n8221), .Z(n8220) );
  XOR U7866 ( .A(n8222), .B(n8223), .Z(n506) );
  AND U7867 ( .A(n8224), .B(n8225), .Z(n8222) );
  XNOR U7868 ( .A(n8223), .B(n8189), .Z(n8225) );
  XNOR U7869 ( .A(n8226), .B(n8227), .Z(n8189) );
  ANDN U7870 ( .B(n8228), .A(n8229), .Z(n8226) );
  XOR U7871 ( .A(n8227), .B(n8230), .Z(n8228) );
  XOR U7872 ( .A(n8223), .B(n8191), .Z(n8224) );
  XNOR U7873 ( .A(n8231), .B(n8232), .Z(n8191) );
  ANDN U7874 ( .B(n8233), .A(n8234), .Z(n8231) );
  XOR U7875 ( .A(n8232), .B(n8235), .Z(n8233) );
  XNOR U7876 ( .A(n8236), .B(n8237), .Z(n8223) );
  NAND U7877 ( .A(n8238), .B(n8239), .Z(n8237) );
  XOR U7878 ( .A(n8240), .B(n8215), .Z(n8239) );
  XOR U7879 ( .A(n8229), .B(n8230), .Z(n8215) );
  XOR U7880 ( .A(n8241), .B(n8242), .Z(n8230) );
  ANDN U7881 ( .B(n8243), .A(n8244), .Z(n8241) );
  XOR U7882 ( .A(n8242), .B(n8245), .Z(n8243) );
  XOR U7883 ( .A(n8246), .B(n8247), .Z(n8229) );
  XOR U7884 ( .A(n8248), .B(n8249), .Z(n8247) );
  ANDN U7885 ( .B(n8250), .A(n8251), .Z(n8248) );
  XOR U7886 ( .A(n8252), .B(n8249), .Z(n8250) );
  IV U7887 ( .A(n8227), .Z(n8246) );
  XOR U7888 ( .A(n8253), .B(n8254), .Z(n8227) );
  ANDN U7889 ( .B(n8255), .A(n8256), .Z(n8253) );
  XOR U7890 ( .A(n8254), .B(n8257), .Z(n8255) );
  IV U7891 ( .A(n8236), .Z(n8240) );
  XNOR U7892 ( .A(n8236), .B(n8217), .Z(n8238) );
  XOR U7893 ( .A(n8258), .B(n8235), .Z(n8217) );
  XOR U7894 ( .A(n8259), .B(n8260), .Z(n8235) );
  ANDN U7895 ( .B(n8261), .A(n8262), .Z(n8259) );
  XOR U7896 ( .A(n8260), .B(n8263), .Z(n8261) );
  IV U7897 ( .A(n8234), .Z(n8258) );
  XOR U7898 ( .A(n8264), .B(n8265), .Z(n8234) );
  XOR U7899 ( .A(n8266), .B(n8267), .Z(n8265) );
  ANDN U7900 ( .B(n8268), .A(n8269), .Z(n8266) );
  XOR U7901 ( .A(n8270), .B(n8267), .Z(n8268) );
  IV U7902 ( .A(n8232), .Z(n8264) );
  XNOR U7903 ( .A(n8271), .B(n8272), .Z(n8232) );
  ANDN U7904 ( .B(n8273), .A(n8274), .Z(n8271) );
  XNOR U7905 ( .A(n8272), .B(n8275), .Z(n8273) );
  NANDN U7906 ( .A(n8219), .B(n8221), .Z(n8236) );
  XOR U7907 ( .A(n8276), .B(n8275), .Z(n8221) );
  XOR U7908 ( .A(n8277), .B(n8263), .Z(n8275) );
  XNOR U7909 ( .A(q[6]), .B(DB[6]), .Z(n8263) );
  IV U7910 ( .A(n8262), .Z(n8277) );
  XNOR U7911 ( .A(n8260), .B(n8278), .Z(n8262) );
  XNOR U7912 ( .A(q[5]), .B(DB[5]), .Z(n8278) );
  XNOR U7913 ( .A(q[4]), .B(DB[4]), .Z(n8260) );
  IV U7914 ( .A(n8274), .Z(n8276) );
  XOR U7915 ( .A(n8279), .B(n8280), .Z(n8274) );
  XOR U7916 ( .A(n8272), .B(n8270), .Z(n8280) );
  XNOR U7917 ( .A(q[3]), .B(DB[3]), .Z(n8270) );
  XOR U7918 ( .A(q[0]), .B(DB[0]), .Z(n8272) );
  IV U7919 ( .A(n8269), .Z(n8279) );
  XNOR U7920 ( .A(n8267), .B(n8281), .Z(n8269) );
  XNOR U7921 ( .A(q[2]), .B(DB[2]), .Z(n8281) );
  XNOR U7922 ( .A(q[1]), .B(DB[1]), .Z(n8267) );
  XOR U7923 ( .A(n8282), .B(n8257), .Z(n8219) );
  XOR U7924 ( .A(n8283), .B(n8245), .Z(n8257) );
  XNOR U7925 ( .A(q[6]), .B(DB[13]), .Z(n8245) );
  IV U7926 ( .A(n8244), .Z(n8283) );
  XNOR U7927 ( .A(n8242), .B(n8284), .Z(n8244) );
  XNOR U7928 ( .A(q[5]), .B(DB[12]), .Z(n8284) );
  XNOR U7929 ( .A(q[4]), .B(DB[11]), .Z(n8242) );
  IV U7930 ( .A(n8256), .Z(n8282) );
  XOR U7931 ( .A(n8285), .B(n8286), .Z(n8256) );
  XNOR U7932 ( .A(n8252), .B(n8254), .Z(n8286) );
  XNOR U7933 ( .A(q[0]), .B(DB[7]), .Z(n8254) );
  XNOR U7934 ( .A(q[3]), .B(DB[10]), .Z(n8252) );
  IV U7935 ( .A(n8251), .Z(n8285) );
  XNOR U7936 ( .A(n8249), .B(n8287), .Z(n8251) );
  XNOR U7937 ( .A(q[2]), .B(DB[9]), .Z(n8287) );
  XNOR U7938 ( .A(q[1]), .B(DB[8]), .Z(n8249) );
  XOR U7939 ( .A(n8288), .B(n8213), .Z(n8176) );
  XOR U7940 ( .A(n8289), .B(n8201), .Z(n8213) );
  XNOR U7941 ( .A(q[6]), .B(DB[20]), .Z(n8201) );
  IV U7942 ( .A(n8200), .Z(n8289) );
  XNOR U7943 ( .A(n8198), .B(n8290), .Z(n8200) );
  XNOR U7944 ( .A(q[5]), .B(DB[19]), .Z(n8290) );
  XNOR U7945 ( .A(q[4]), .B(DB[18]), .Z(n8198) );
  IV U7946 ( .A(n8212), .Z(n8288) );
  XOR U7947 ( .A(n8291), .B(n8292), .Z(n8212) );
  XNOR U7948 ( .A(n8208), .B(n8210), .Z(n8292) );
  XNOR U7949 ( .A(q[0]), .B(DB[14]), .Z(n8210) );
  XNOR U7950 ( .A(q[3]), .B(DB[17]), .Z(n8208) );
  IV U7951 ( .A(n8207), .Z(n8291) );
  XNOR U7952 ( .A(n8205), .B(n8293), .Z(n8207) );
  XNOR U7953 ( .A(q[2]), .B(DB[16]), .Z(n8293) );
  XNOR U7954 ( .A(q[1]), .B(DB[15]), .Z(n8205) );
  XOR U7955 ( .A(n8294), .B(n8170), .Z(n8133) );
  XOR U7956 ( .A(n8295), .B(n8158), .Z(n8170) );
  XNOR U7957 ( .A(q[6]), .B(DB[27]), .Z(n8158) );
  IV U7958 ( .A(n8157), .Z(n8295) );
  XNOR U7959 ( .A(n8155), .B(n8296), .Z(n8157) );
  XNOR U7960 ( .A(q[5]), .B(DB[26]), .Z(n8296) );
  XNOR U7961 ( .A(q[4]), .B(DB[25]), .Z(n8155) );
  IV U7962 ( .A(n8169), .Z(n8294) );
  XOR U7963 ( .A(n8297), .B(n8298), .Z(n8169) );
  XNOR U7964 ( .A(n8165), .B(n8167), .Z(n8298) );
  XNOR U7965 ( .A(q[0]), .B(DB[21]), .Z(n8167) );
  XNOR U7966 ( .A(q[3]), .B(DB[24]), .Z(n8165) );
  IV U7967 ( .A(n8164), .Z(n8297) );
  XNOR U7968 ( .A(n8162), .B(n8299), .Z(n8164) );
  XNOR U7969 ( .A(q[2]), .B(DB[23]), .Z(n8299) );
  XNOR U7970 ( .A(q[1]), .B(DB[22]), .Z(n8162) );
  XOR U7971 ( .A(n8300), .B(n8127), .Z(n8090) );
  XOR U7972 ( .A(n8301), .B(n8115), .Z(n8127) );
  XNOR U7973 ( .A(q[6]), .B(DB[34]), .Z(n8115) );
  IV U7974 ( .A(n8114), .Z(n8301) );
  XNOR U7975 ( .A(n8112), .B(n8302), .Z(n8114) );
  XNOR U7976 ( .A(q[5]), .B(DB[33]), .Z(n8302) );
  XNOR U7977 ( .A(q[4]), .B(DB[32]), .Z(n8112) );
  IV U7978 ( .A(n8126), .Z(n8300) );
  XOR U7979 ( .A(n8303), .B(n8304), .Z(n8126) );
  XNOR U7980 ( .A(n8122), .B(n8124), .Z(n8304) );
  XNOR U7981 ( .A(q[0]), .B(DB[28]), .Z(n8124) );
  XNOR U7982 ( .A(q[3]), .B(DB[31]), .Z(n8122) );
  IV U7983 ( .A(n8121), .Z(n8303) );
  XNOR U7984 ( .A(n8119), .B(n8305), .Z(n8121) );
  XNOR U7985 ( .A(q[2]), .B(DB[30]), .Z(n8305) );
  XNOR U7986 ( .A(q[1]), .B(DB[29]), .Z(n8119) );
  XOR U7987 ( .A(n8306), .B(n8084), .Z(n8047) );
  XOR U7988 ( .A(n8307), .B(n8072), .Z(n8084) );
  XNOR U7989 ( .A(q[6]), .B(DB[41]), .Z(n8072) );
  IV U7990 ( .A(n8071), .Z(n8307) );
  XNOR U7991 ( .A(n8069), .B(n8308), .Z(n8071) );
  XNOR U7992 ( .A(q[5]), .B(DB[40]), .Z(n8308) );
  XNOR U7993 ( .A(q[4]), .B(DB[39]), .Z(n8069) );
  IV U7994 ( .A(n8083), .Z(n8306) );
  XOR U7995 ( .A(n8309), .B(n8310), .Z(n8083) );
  XNOR U7996 ( .A(n8079), .B(n8081), .Z(n8310) );
  XNOR U7997 ( .A(q[0]), .B(DB[35]), .Z(n8081) );
  XNOR U7998 ( .A(q[3]), .B(DB[38]), .Z(n8079) );
  IV U7999 ( .A(n8078), .Z(n8309) );
  XNOR U8000 ( .A(n8076), .B(n8311), .Z(n8078) );
  XNOR U8001 ( .A(q[2]), .B(DB[37]), .Z(n8311) );
  XNOR U8002 ( .A(q[1]), .B(DB[36]), .Z(n8076) );
  XOR U8003 ( .A(n8312), .B(n8041), .Z(n8004) );
  XOR U8004 ( .A(n8313), .B(n8029), .Z(n8041) );
  XNOR U8005 ( .A(q[6]), .B(DB[48]), .Z(n8029) );
  IV U8006 ( .A(n8028), .Z(n8313) );
  XNOR U8007 ( .A(n8026), .B(n8314), .Z(n8028) );
  XNOR U8008 ( .A(q[5]), .B(DB[47]), .Z(n8314) );
  XNOR U8009 ( .A(q[4]), .B(DB[46]), .Z(n8026) );
  IV U8010 ( .A(n8040), .Z(n8312) );
  XOR U8011 ( .A(n8315), .B(n8316), .Z(n8040) );
  XNOR U8012 ( .A(n8036), .B(n8038), .Z(n8316) );
  XNOR U8013 ( .A(q[0]), .B(DB[42]), .Z(n8038) );
  XNOR U8014 ( .A(q[3]), .B(DB[45]), .Z(n8036) );
  IV U8015 ( .A(n8035), .Z(n8315) );
  XNOR U8016 ( .A(n8033), .B(n8317), .Z(n8035) );
  XNOR U8017 ( .A(q[2]), .B(DB[44]), .Z(n8317) );
  XNOR U8018 ( .A(q[1]), .B(DB[43]), .Z(n8033) );
  XOR U8019 ( .A(n8318), .B(n7998), .Z(n7961) );
  XOR U8020 ( .A(n8319), .B(n7986), .Z(n7998) );
  XNOR U8021 ( .A(q[6]), .B(DB[55]), .Z(n7986) );
  IV U8022 ( .A(n7985), .Z(n8319) );
  XNOR U8023 ( .A(n7983), .B(n8320), .Z(n7985) );
  XNOR U8024 ( .A(q[5]), .B(DB[54]), .Z(n8320) );
  XNOR U8025 ( .A(q[4]), .B(DB[53]), .Z(n7983) );
  IV U8026 ( .A(n7997), .Z(n8318) );
  XOR U8027 ( .A(n8321), .B(n8322), .Z(n7997) );
  XNOR U8028 ( .A(n7993), .B(n7995), .Z(n8322) );
  XNOR U8029 ( .A(q[0]), .B(DB[49]), .Z(n7995) );
  XNOR U8030 ( .A(q[3]), .B(DB[52]), .Z(n7993) );
  IV U8031 ( .A(n7992), .Z(n8321) );
  XNOR U8032 ( .A(n7990), .B(n8323), .Z(n7992) );
  XNOR U8033 ( .A(q[2]), .B(DB[51]), .Z(n8323) );
  XNOR U8034 ( .A(q[1]), .B(DB[50]), .Z(n7990) );
  XOR U8035 ( .A(n8324), .B(n7955), .Z(n7918) );
  XOR U8036 ( .A(n8325), .B(n7943), .Z(n7955) );
  XNOR U8037 ( .A(q[6]), .B(DB[62]), .Z(n7943) );
  IV U8038 ( .A(n7942), .Z(n8325) );
  XNOR U8039 ( .A(n7940), .B(n8326), .Z(n7942) );
  XNOR U8040 ( .A(q[5]), .B(DB[61]), .Z(n8326) );
  XNOR U8041 ( .A(q[4]), .B(DB[60]), .Z(n7940) );
  IV U8042 ( .A(n7954), .Z(n8324) );
  XOR U8043 ( .A(n8327), .B(n8328), .Z(n7954) );
  XNOR U8044 ( .A(n7950), .B(n7952), .Z(n8328) );
  XNOR U8045 ( .A(q[0]), .B(DB[56]), .Z(n7952) );
  XNOR U8046 ( .A(q[3]), .B(DB[59]), .Z(n7950) );
  IV U8047 ( .A(n7949), .Z(n8327) );
  XNOR U8048 ( .A(n7947), .B(n8329), .Z(n7949) );
  XNOR U8049 ( .A(q[2]), .B(DB[58]), .Z(n8329) );
  XNOR U8050 ( .A(q[1]), .B(DB[57]), .Z(n7947) );
  XOR U8051 ( .A(n8330), .B(n7912), .Z(n7875) );
  XOR U8052 ( .A(n8331), .B(n7900), .Z(n7912) );
  XNOR U8053 ( .A(q[6]), .B(DB[69]), .Z(n7900) );
  IV U8054 ( .A(n7899), .Z(n8331) );
  XNOR U8055 ( .A(n7897), .B(n8332), .Z(n7899) );
  XNOR U8056 ( .A(q[5]), .B(DB[68]), .Z(n8332) );
  XNOR U8057 ( .A(q[4]), .B(DB[67]), .Z(n7897) );
  IV U8058 ( .A(n7911), .Z(n8330) );
  XOR U8059 ( .A(n8333), .B(n8334), .Z(n7911) );
  XNOR U8060 ( .A(n7907), .B(n7909), .Z(n8334) );
  XNOR U8061 ( .A(q[0]), .B(DB[63]), .Z(n7909) );
  XNOR U8062 ( .A(q[3]), .B(DB[66]), .Z(n7907) );
  IV U8063 ( .A(n7906), .Z(n8333) );
  XNOR U8064 ( .A(n7904), .B(n8335), .Z(n7906) );
  XNOR U8065 ( .A(q[2]), .B(DB[65]), .Z(n8335) );
  XNOR U8066 ( .A(q[1]), .B(DB[64]), .Z(n7904) );
  XOR U8067 ( .A(n8336), .B(n7869), .Z(n7832) );
  XOR U8068 ( .A(n8337), .B(n7857), .Z(n7869) );
  XNOR U8069 ( .A(q[6]), .B(DB[76]), .Z(n7857) );
  IV U8070 ( .A(n7856), .Z(n8337) );
  XNOR U8071 ( .A(n7854), .B(n8338), .Z(n7856) );
  XNOR U8072 ( .A(q[5]), .B(DB[75]), .Z(n8338) );
  XNOR U8073 ( .A(q[4]), .B(DB[74]), .Z(n7854) );
  IV U8074 ( .A(n7868), .Z(n8336) );
  XOR U8075 ( .A(n8339), .B(n8340), .Z(n7868) );
  XNOR U8076 ( .A(n7864), .B(n7866), .Z(n8340) );
  XNOR U8077 ( .A(q[0]), .B(DB[70]), .Z(n7866) );
  XNOR U8078 ( .A(q[3]), .B(DB[73]), .Z(n7864) );
  IV U8079 ( .A(n7863), .Z(n8339) );
  XNOR U8080 ( .A(n7861), .B(n8341), .Z(n7863) );
  XNOR U8081 ( .A(q[2]), .B(DB[72]), .Z(n8341) );
  XNOR U8082 ( .A(q[1]), .B(DB[71]), .Z(n7861) );
  XOR U8083 ( .A(n8342), .B(n7826), .Z(n7789) );
  XOR U8084 ( .A(n8343), .B(n7814), .Z(n7826) );
  XNOR U8085 ( .A(q[6]), .B(DB[83]), .Z(n7814) );
  IV U8086 ( .A(n7813), .Z(n8343) );
  XNOR U8087 ( .A(n7811), .B(n8344), .Z(n7813) );
  XNOR U8088 ( .A(q[5]), .B(DB[82]), .Z(n8344) );
  XNOR U8089 ( .A(q[4]), .B(DB[81]), .Z(n7811) );
  IV U8090 ( .A(n7825), .Z(n8342) );
  XOR U8091 ( .A(n8345), .B(n8346), .Z(n7825) );
  XNOR U8092 ( .A(n7821), .B(n7823), .Z(n8346) );
  XNOR U8093 ( .A(q[0]), .B(DB[77]), .Z(n7823) );
  XNOR U8094 ( .A(q[3]), .B(DB[80]), .Z(n7821) );
  IV U8095 ( .A(n7820), .Z(n8345) );
  XNOR U8096 ( .A(n7818), .B(n8347), .Z(n7820) );
  XNOR U8097 ( .A(q[2]), .B(DB[79]), .Z(n8347) );
  XNOR U8098 ( .A(q[1]), .B(DB[78]), .Z(n7818) );
  XOR U8099 ( .A(n8348), .B(n7783), .Z(n7746) );
  XOR U8100 ( .A(n8349), .B(n7771), .Z(n7783) );
  XNOR U8101 ( .A(q[6]), .B(DB[90]), .Z(n7771) );
  IV U8102 ( .A(n7770), .Z(n8349) );
  XNOR U8103 ( .A(n7768), .B(n8350), .Z(n7770) );
  XNOR U8104 ( .A(q[5]), .B(DB[89]), .Z(n8350) );
  XNOR U8105 ( .A(q[4]), .B(DB[88]), .Z(n7768) );
  IV U8106 ( .A(n7782), .Z(n8348) );
  XOR U8107 ( .A(n8351), .B(n8352), .Z(n7782) );
  XNOR U8108 ( .A(n7778), .B(n7780), .Z(n8352) );
  XNOR U8109 ( .A(q[0]), .B(DB[84]), .Z(n7780) );
  XNOR U8110 ( .A(q[3]), .B(DB[87]), .Z(n7778) );
  IV U8111 ( .A(n7777), .Z(n8351) );
  XNOR U8112 ( .A(n7775), .B(n8353), .Z(n7777) );
  XNOR U8113 ( .A(q[2]), .B(DB[86]), .Z(n8353) );
  XNOR U8114 ( .A(q[1]), .B(DB[85]), .Z(n7775) );
  XOR U8115 ( .A(n8354), .B(n7740), .Z(n7703) );
  XOR U8116 ( .A(n8355), .B(n7728), .Z(n7740) );
  XNOR U8117 ( .A(q[6]), .B(DB[97]), .Z(n7728) );
  IV U8118 ( .A(n7727), .Z(n8355) );
  XNOR U8119 ( .A(n7725), .B(n8356), .Z(n7727) );
  XNOR U8120 ( .A(q[5]), .B(DB[96]), .Z(n8356) );
  XNOR U8121 ( .A(q[4]), .B(DB[95]), .Z(n7725) );
  IV U8122 ( .A(n7739), .Z(n8354) );
  XOR U8123 ( .A(n8357), .B(n8358), .Z(n7739) );
  XNOR U8124 ( .A(n7735), .B(n7737), .Z(n8358) );
  XNOR U8125 ( .A(q[0]), .B(DB[91]), .Z(n7737) );
  XNOR U8126 ( .A(q[3]), .B(DB[94]), .Z(n7735) );
  IV U8127 ( .A(n7734), .Z(n8357) );
  XNOR U8128 ( .A(n7732), .B(n8359), .Z(n7734) );
  XNOR U8129 ( .A(q[2]), .B(DB[93]), .Z(n8359) );
  XNOR U8130 ( .A(q[1]), .B(DB[92]), .Z(n7732) );
  XOR U8131 ( .A(n8360), .B(n7697), .Z(n7660) );
  XOR U8132 ( .A(n8361), .B(n7685), .Z(n7697) );
  XNOR U8133 ( .A(q[6]), .B(DB[104]), .Z(n7685) );
  IV U8134 ( .A(n7684), .Z(n8361) );
  XNOR U8135 ( .A(n7682), .B(n8362), .Z(n7684) );
  XNOR U8136 ( .A(q[5]), .B(DB[103]), .Z(n8362) );
  XNOR U8137 ( .A(q[4]), .B(DB[102]), .Z(n7682) );
  IV U8138 ( .A(n7696), .Z(n8360) );
  XOR U8139 ( .A(n8363), .B(n8364), .Z(n7696) );
  XNOR U8140 ( .A(n7692), .B(n7694), .Z(n8364) );
  XNOR U8141 ( .A(q[0]), .B(DB[98]), .Z(n7694) );
  XNOR U8142 ( .A(q[3]), .B(DB[101]), .Z(n7692) );
  IV U8143 ( .A(n7691), .Z(n8363) );
  XNOR U8144 ( .A(n7689), .B(n8365), .Z(n7691) );
  XNOR U8145 ( .A(q[2]), .B(DB[100]), .Z(n8365) );
  XNOR U8146 ( .A(q[1]), .B(DB[99]), .Z(n7689) );
  XOR U8147 ( .A(n8366), .B(n7654), .Z(n7617) );
  XOR U8148 ( .A(n8367), .B(n7642), .Z(n7654) );
  XNOR U8149 ( .A(q[6]), .B(DB[111]), .Z(n7642) );
  IV U8150 ( .A(n7641), .Z(n8367) );
  XNOR U8151 ( .A(n7639), .B(n8368), .Z(n7641) );
  XNOR U8152 ( .A(q[5]), .B(DB[110]), .Z(n8368) );
  XNOR U8153 ( .A(q[4]), .B(DB[109]), .Z(n7639) );
  IV U8154 ( .A(n7653), .Z(n8366) );
  XOR U8155 ( .A(n8369), .B(n8370), .Z(n7653) );
  XNOR U8156 ( .A(n7649), .B(n7651), .Z(n8370) );
  XNOR U8157 ( .A(q[0]), .B(DB[105]), .Z(n7651) );
  XNOR U8158 ( .A(q[3]), .B(DB[108]), .Z(n7649) );
  IV U8159 ( .A(n7648), .Z(n8369) );
  XNOR U8160 ( .A(n7646), .B(n8371), .Z(n7648) );
  XNOR U8161 ( .A(q[2]), .B(DB[107]), .Z(n8371) );
  XNOR U8162 ( .A(q[1]), .B(DB[106]), .Z(n7646) );
  XOR U8163 ( .A(n8372), .B(n7611), .Z(n7574) );
  XOR U8164 ( .A(n8373), .B(n7599), .Z(n7611) );
  XNOR U8165 ( .A(q[6]), .B(DB[118]), .Z(n7599) );
  IV U8166 ( .A(n7598), .Z(n8373) );
  XNOR U8167 ( .A(n7596), .B(n8374), .Z(n7598) );
  XNOR U8168 ( .A(q[5]), .B(DB[117]), .Z(n8374) );
  XNOR U8169 ( .A(q[4]), .B(DB[116]), .Z(n7596) );
  IV U8170 ( .A(n7610), .Z(n8372) );
  XOR U8171 ( .A(n8375), .B(n8376), .Z(n7610) );
  XNOR U8172 ( .A(n7606), .B(n7608), .Z(n8376) );
  XNOR U8173 ( .A(q[0]), .B(DB[112]), .Z(n7608) );
  XNOR U8174 ( .A(q[3]), .B(DB[115]), .Z(n7606) );
  IV U8175 ( .A(n7605), .Z(n8375) );
  XNOR U8176 ( .A(n7603), .B(n8377), .Z(n7605) );
  XNOR U8177 ( .A(q[2]), .B(DB[114]), .Z(n8377) );
  XNOR U8178 ( .A(q[1]), .B(DB[113]), .Z(n7603) );
  XOR U8179 ( .A(n8378), .B(n7568), .Z(n7531) );
  XOR U8180 ( .A(n8379), .B(n7556), .Z(n7568) );
  XNOR U8181 ( .A(q[6]), .B(DB[125]), .Z(n7556) );
  IV U8182 ( .A(n7555), .Z(n8379) );
  XNOR U8183 ( .A(n7553), .B(n8380), .Z(n7555) );
  XNOR U8184 ( .A(q[5]), .B(DB[124]), .Z(n8380) );
  XNOR U8185 ( .A(q[4]), .B(DB[123]), .Z(n7553) );
  IV U8186 ( .A(n7567), .Z(n8378) );
  XOR U8187 ( .A(n8381), .B(n8382), .Z(n7567) );
  XNOR U8188 ( .A(n7563), .B(n7565), .Z(n8382) );
  XNOR U8189 ( .A(q[0]), .B(DB[119]), .Z(n7565) );
  XNOR U8190 ( .A(q[3]), .B(DB[122]), .Z(n7563) );
  IV U8191 ( .A(n7562), .Z(n8381) );
  XNOR U8192 ( .A(n7560), .B(n8383), .Z(n7562) );
  XNOR U8193 ( .A(q[2]), .B(DB[121]), .Z(n8383) );
  XNOR U8194 ( .A(q[1]), .B(DB[120]), .Z(n7560) );
  XOR U8195 ( .A(n8384), .B(n7525), .Z(n7488) );
  XOR U8196 ( .A(n8385), .B(n7513), .Z(n7525) );
  XNOR U8197 ( .A(q[6]), .B(DB[132]), .Z(n7513) );
  IV U8198 ( .A(n7512), .Z(n8385) );
  XNOR U8199 ( .A(n7510), .B(n8386), .Z(n7512) );
  XNOR U8200 ( .A(q[5]), .B(DB[131]), .Z(n8386) );
  XNOR U8201 ( .A(q[4]), .B(DB[130]), .Z(n7510) );
  IV U8202 ( .A(n7524), .Z(n8384) );
  XOR U8203 ( .A(n8387), .B(n8388), .Z(n7524) );
  XNOR U8204 ( .A(n7520), .B(n7522), .Z(n8388) );
  XNOR U8205 ( .A(q[0]), .B(DB[126]), .Z(n7522) );
  XNOR U8206 ( .A(q[3]), .B(DB[129]), .Z(n7520) );
  IV U8207 ( .A(n7519), .Z(n8387) );
  XNOR U8208 ( .A(n7517), .B(n8389), .Z(n7519) );
  XNOR U8209 ( .A(q[2]), .B(DB[128]), .Z(n8389) );
  XNOR U8210 ( .A(q[1]), .B(DB[127]), .Z(n7517) );
  XOR U8211 ( .A(n8390), .B(n7482), .Z(n7445) );
  XOR U8212 ( .A(n8391), .B(n7470), .Z(n7482) );
  XNOR U8213 ( .A(q[6]), .B(DB[139]), .Z(n7470) );
  IV U8214 ( .A(n7469), .Z(n8391) );
  XNOR U8215 ( .A(n7467), .B(n8392), .Z(n7469) );
  XNOR U8216 ( .A(q[5]), .B(DB[138]), .Z(n8392) );
  XNOR U8217 ( .A(q[4]), .B(DB[137]), .Z(n7467) );
  IV U8218 ( .A(n7481), .Z(n8390) );
  XOR U8219 ( .A(n8393), .B(n8394), .Z(n7481) );
  XNOR U8220 ( .A(n7477), .B(n7479), .Z(n8394) );
  XNOR U8221 ( .A(q[0]), .B(DB[133]), .Z(n7479) );
  XNOR U8222 ( .A(q[3]), .B(DB[136]), .Z(n7477) );
  IV U8223 ( .A(n7476), .Z(n8393) );
  XNOR U8224 ( .A(n7474), .B(n8395), .Z(n7476) );
  XNOR U8225 ( .A(q[2]), .B(DB[135]), .Z(n8395) );
  XNOR U8226 ( .A(q[1]), .B(DB[134]), .Z(n7474) );
  XOR U8227 ( .A(n8396), .B(n7439), .Z(n7402) );
  XOR U8228 ( .A(n8397), .B(n7427), .Z(n7439) );
  XNOR U8229 ( .A(q[6]), .B(DB[146]), .Z(n7427) );
  IV U8230 ( .A(n7426), .Z(n8397) );
  XNOR U8231 ( .A(n7424), .B(n8398), .Z(n7426) );
  XNOR U8232 ( .A(q[5]), .B(DB[145]), .Z(n8398) );
  XNOR U8233 ( .A(q[4]), .B(DB[144]), .Z(n7424) );
  IV U8234 ( .A(n7438), .Z(n8396) );
  XOR U8235 ( .A(n8399), .B(n8400), .Z(n7438) );
  XNOR U8236 ( .A(n7434), .B(n7436), .Z(n8400) );
  XNOR U8237 ( .A(q[0]), .B(DB[140]), .Z(n7436) );
  XNOR U8238 ( .A(q[3]), .B(DB[143]), .Z(n7434) );
  IV U8239 ( .A(n7433), .Z(n8399) );
  XNOR U8240 ( .A(n7431), .B(n8401), .Z(n7433) );
  XNOR U8241 ( .A(q[2]), .B(DB[142]), .Z(n8401) );
  XNOR U8242 ( .A(q[1]), .B(DB[141]), .Z(n7431) );
  XOR U8243 ( .A(n8402), .B(n7396), .Z(n7359) );
  XOR U8244 ( .A(n8403), .B(n7384), .Z(n7396) );
  XNOR U8245 ( .A(q[6]), .B(DB[153]), .Z(n7384) );
  IV U8246 ( .A(n7383), .Z(n8403) );
  XNOR U8247 ( .A(n7381), .B(n8404), .Z(n7383) );
  XNOR U8248 ( .A(q[5]), .B(DB[152]), .Z(n8404) );
  XNOR U8249 ( .A(q[4]), .B(DB[151]), .Z(n7381) );
  IV U8250 ( .A(n7395), .Z(n8402) );
  XOR U8251 ( .A(n8405), .B(n8406), .Z(n7395) );
  XNOR U8252 ( .A(n7391), .B(n7393), .Z(n8406) );
  XNOR U8253 ( .A(q[0]), .B(DB[147]), .Z(n7393) );
  XNOR U8254 ( .A(q[3]), .B(DB[150]), .Z(n7391) );
  IV U8255 ( .A(n7390), .Z(n8405) );
  XNOR U8256 ( .A(n7388), .B(n8407), .Z(n7390) );
  XNOR U8257 ( .A(q[2]), .B(DB[149]), .Z(n8407) );
  XNOR U8258 ( .A(q[1]), .B(DB[148]), .Z(n7388) );
  XOR U8259 ( .A(n8408), .B(n7353), .Z(n7316) );
  XOR U8260 ( .A(n8409), .B(n7341), .Z(n7353) );
  XNOR U8261 ( .A(q[6]), .B(DB[160]), .Z(n7341) );
  IV U8262 ( .A(n7340), .Z(n8409) );
  XNOR U8263 ( .A(n7338), .B(n8410), .Z(n7340) );
  XNOR U8264 ( .A(q[5]), .B(DB[159]), .Z(n8410) );
  XNOR U8265 ( .A(q[4]), .B(DB[158]), .Z(n7338) );
  IV U8266 ( .A(n7352), .Z(n8408) );
  XOR U8267 ( .A(n8411), .B(n8412), .Z(n7352) );
  XNOR U8268 ( .A(n7348), .B(n7350), .Z(n8412) );
  XNOR U8269 ( .A(q[0]), .B(DB[154]), .Z(n7350) );
  XNOR U8270 ( .A(q[3]), .B(DB[157]), .Z(n7348) );
  IV U8271 ( .A(n7347), .Z(n8411) );
  XNOR U8272 ( .A(n7345), .B(n8413), .Z(n7347) );
  XNOR U8273 ( .A(q[2]), .B(DB[156]), .Z(n8413) );
  XNOR U8274 ( .A(q[1]), .B(DB[155]), .Z(n7345) );
  XOR U8275 ( .A(n8414), .B(n7310), .Z(n7273) );
  XOR U8276 ( .A(n8415), .B(n7298), .Z(n7310) );
  XNOR U8277 ( .A(q[6]), .B(DB[167]), .Z(n7298) );
  IV U8278 ( .A(n7297), .Z(n8415) );
  XNOR U8279 ( .A(n7295), .B(n8416), .Z(n7297) );
  XNOR U8280 ( .A(q[5]), .B(DB[166]), .Z(n8416) );
  XNOR U8281 ( .A(q[4]), .B(DB[165]), .Z(n7295) );
  IV U8282 ( .A(n7309), .Z(n8414) );
  XOR U8283 ( .A(n8417), .B(n8418), .Z(n7309) );
  XNOR U8284 ( .A(n7305), .B(n7307), .Z(n8418) );
  XNOR U8285 ( .A(q[0]), .B(DB[161]), .Z(n7307) );
  XNOR U8286 ( .A(q[3]), .B(DB[164]), .Z(n7305) );
  IV U8287 ( .A(n7304), .Z(n8417) );
  XNOR U8288 ( .A(n7302), .B(n8419), .Z(n7304) );
  XNOR U8289 ( .A(q[2]), .B(DB[163]), .Z(n8419) );
  XNOR U8290 ( .A(q[1]), .B(DB[162]), .Z(n7302) );
  XOR U8291 ( .A(n8420), .B(n7267), .Z(n7230) );
  XOR U8292 ( .A(n8421), .B(n7255), .Z(n7267) );
  XNOR U8293 ( .A(q[6]), .B(DB[174]), .Z(n7255) );
  IV U8294 ( .A(n7254), .Z(n8421) );
  XNOR U8295 ( .A(n7252), .B(n8422), .Z(n7254) );
  XNOR U8296 ( .A(q[5]), .B(DB[173]), .Z(n8422) );
  XNOR U8297 ( .A(q[4]), .B(DB[172]), .Z(n7252) );
  IV U8298 ( .A(n7266), .Z(n8420) );
  XOR U8299 ( .A(n8423), .B(n8424), .Z(n7266) );
  XNOR U8300 ( .A(n7262), .B(n7264), .Z(n8424) );
  XNOR U8301 ( .A(q[0]), .B(DB[168]), .Z(n7264) );
  XNOR U8302 ( .A(q[3]), .B(DB[171]), .Z(n7262) );
  IV U8303 ( .A(n7261), .Z(n8423) );
  XNOR U8304 ( .A(n7259), .B(n8425), .Z(n7261) );
  XNOR U8305 ( .A(q[2]), .B(DB[170]), .Z(n8425) );
  XNOR U8306 ( .A(q[1]), .B(DB[169]), .Z(n7259) );
  XOR U8307 ( .A(n8426), .B(n7224), .Z(n7187) );
  XOR U8308 ( .A(n8427), .B(n7212), .Z(n7224) );
  XNOR U8309 ( .A(q[6]), .B(DB[181]), .Z(n7212) );
  IV U8310 ( .A(n7211), .Z(n8427) );
  XNOR U8311 ( .A(n7209), .B(n8428), .Z(n7211) );
  XNOR U8312 ( .A(q[5]), .B(DB[180]), .Z(n8428) );
  XNOR U8313 ( .A(q[4]), .B(DB[179]), .Z(n7209) );
  IV U8314 ( .A(n7223), .Z(n8426) );
  XOR U8315 ( .A(n8429), .B(n8430), .Z(n7223) );
  XNOR U8316 ( .A(n7219), .B(n7221), .Z(n8430) );
  XNOR U8317 ( .A(q[0]), .B(DB[175]), .Z(n7221) );
  XNOR U8318 ( .A(q[3]), .B(DB[178]), .Z(n7219) );
  IV U8319 ( .A(n7218), .Z(n8429) );
  XNOR U8320 ( .A(n7216), .B(n8431), .Z(n7218) );
  XNOR U8321 ( .A(q[2]), .B(DB[177]), .Z(n8431) );
  XNOR U8322 ( .A(q[1]), .B(DB[176]), .Z(n7216) );
  XOR U8323 ( .A(n8432), .B(n7181), .Z(n7144) );
  XOR U8324 ( .A(n8433), .B(n7169), .Z(n7181) );
  XNOR U8325 ( .A(q[6]), .B(DB[188]), .Z(n7169) );
  IV U8326 ( .A(n7168), .Z(n8433) );
  XNOR U8327 ( .A(n7166), .B(n8434), .Z(n7168) );
  XNOR U8328 ( .A(q[5]), .B(DB[187]), .Z(n8434) );
  XNOR U8329 ( .A(q[4]), .B(DB[186]), .Z(n7166) );
  IV U8330 ( .A(n7180), .Z(n8432) );
  XOR U8331 ( .A(n8435), .B(n8436), .Z(n7180) );
  XNOR U8332 ( .A(n7176), .B(n7178), .Z(n8436) );
  XNOR U8333 ( .A(q[0]), .B(DB[182]), .Z(n7178) );
  XNOR U8334 ( .A(q[3]), .B(DB[185]), .Z(n7176) );
  IV U8335 ( .A(n7175), .Z(n8435) );
  XNOR U8336 ( .A(n7173), .B(n8437), .Z(n7175) );
  XNOR U8337 ( .A(q[2]), .B(DB[184]), .Z(n8437) );
  XNOR U8338 ( .A(q[1]), .B(DB[183]), .Z(n7173) );
  XOR U8339 ( .A(n8438), .B(n7138), .Z(n7101) );
  XOR U8340 ( .A(n8439), .B(n7126), .Z(n7138) );
  XNOR U8341 ( .A(q[6]), .B(DB[195]), .Z(n7126) );
  IV U8342 ( .A(n7125), .Z(n8439) );
  XNOR U8343 ( .A(n7123), .B(n8440), .Z(n7125) );
  XNOR U8344 ( .A(q[5]), .B(DB[194]), .Z(n8440) );
  XNOR U8345 ( .A(q[4]), .B(DB[193]), .Z(n7123) );
  IV U8346 ( .A(n7137), .Z(n8438) );
  XOR U8347 ( .A(n8441), .B(n8442), .Z(n7137) );
  XNOR U8348 ( .A(n7133), .B(n7135), .Z(n8442) );
  XNOR U8349 ( .A(q[0]), .B(DB[189]), .Z(n7135) );
  XNOR U8350 ( .A(q[3]), .B(DB[192]), .Z(n7133) );
  IV U8351 ( .A(n7132), .Z(n8441) );
  XNOR U8352 ( .A(n7130), .B(n8443), .Z(n7132) );
  XNOR U8353 ( .A(q[2]), .B(DB[191]), .Z(n8443) );
  XNOR U8354 ( .A(q[1]), .B(DB[190]), .Z(n7130) );
  XOR U8355 ( .A(n8444), .B(n7095), .Z(n7058) );
  XOR U8356 ( .A(n8445), .B(n7083), .Z(n7095) );
  XNOR U8357 ( .A(q[6]), .B(DB[202]), .Z(n7083) );
  IV U8358 ( .A(n7082), .Z(n8445) );
  XNOR U8359 ( .A(n7080), .B(n8446), .Z(n7082) );
  XNOR U8360 ( .A(q[5]), .B(DB[201]), .Z(n8446) );
  XNOR U8361 ( .A(q[4]), .B(DB[200]), .Z(n7080) );
  IV U8362 ( .A(n7094), .Z(n8444) );
  XOR U8363 ( .A(n8447), .B(n8448), .Z(n7094) );
  XNOR U8364 ( .A(n7090), .B(n7092), .Z(n8448) );
  XNOR U8365 ( .A(q[0]), .B(DB[196]), .Z(n7092) );
  XNOR U8366 ( .A(q[3]), .B(DB[199]), .Z(n7090) );
  IV U8367 ( .A(n7089), .Z(n8447) );
  XNOR U8368 ( .A(n7087), .B(n8449), .Z(n7089) );
  XNOR U8369 ( .A(q[2]), .B(DB[198]), .Z(n8449) );
  XNOR U8370 ( .A(q[1]), .B(DB[197]), .Z(n7087) );
  XOR U8371 ( .A(n8450), .B(n7052), .Z(n7015) );
  XOR U8372 ( .A(n8451), .B(n7040), .Z(n7052) );
  XNOR U8373 ( .A(q[6]), .B(DB[209]), .Z(n7040) );
  IV U8374 ( .A(n7039), .Z(n8451) );
  XNOR U8375 ( .A(n7037), .B(n8452), .Z(n7039) );
  XNOR U8376 ( .A(q[5]), .B(DB[208]), .Z(n8452) );
  XNOR U8377 ( .A(q[4]), .B(DB[207]), .Z(n7037) );
  IV U8378 ( .A(n7051), .Z(n8450) );
  XOR U8379 ( .A(n8453), .B(n8454), .Z(n7051) );
  XNOR U8380 ( .A(n7047), .B(n7049), .Z(n8454) );
  XNOR U8381 ( .A(q[0]), .B(DB[203]), .Z(n7049) );
  XNOR U8382 ( .A(q[3]), .B(DB[206]), .Z(n7047) );
  IV U8383 ( .A(n7046), .Z(n8453) );
  XNOR U8384 ( .A(n7044), .B(n8455), .Z(n7046) );
  XNOR U8385 ( .A(q[2]), .B(DB[205]), .Z(n8455) );
  XNOR U8386 ( .A(q[1]), .B(DB[204]), .Z(n7044) );
  XOR U8387 ( .A(n8456), .B(n7009), .Z(n6972) );
  XOR U8388 ( .A(n8457), .B(n6997), .Z(n7009) );
  XNOR U8389 ( .A(q[6]), .B(DB[216]), .Z(n6997) );
  IV U8390 ( .A(n6996), .Z(n8457) );
  XNOR U8391 ( .A(n6994), .B(n8458), .Z(n6996) );
  XNOR U8392 ( .A(q[5]), .B(DB[215]), .Z(n8458) );
  XNOR U8393 ( .A(q[4]), .B(DB[214]), .Z(n6994) );
  IV U8394 ( .A(n7008), .Z(n8456) );
  XOR U8395 ( .A(n8459), .B(n8460), .Z(n7008) );
  XNOR U8396 ( .A(n7004), .B(n7006), .Z(n8460) );
  XNOR U8397 ( .A(q[0]), .B(DB[210]), .Z(n7006) );
  XNOR U8398 ( .A(q[3]), .B(DB[213]), .Z(n7004) );
  IV U8399 ( .A(n7003), .Z(n8459) );
  XNOR U8400 ( .A(n7001), .B(n8461), .Z(n7003) );
  XNOR U8401 ( .A(q[2]), .B(DB[212]), .Z(n8461) );
  XNOR U8402 ( .A(q[1]), .B(DB[211]), .Z(n7001) );
  XOR U8403 ( .A(n8462), .B(n6966), .Z(n6929) );
  XOR U8404 ( .A(n8463), .B(n6954), .Z(n6966) );
  XNOR U8405 ( .A(q[6]), .B(DB[223]), .Z(n6954) );
  IV U8406 ( .A(n6953), .Z(n8463) );
  XNOR U8407 ( .A(n6951), .B(n8464), .Z(n6953) );
  XNOR U8408 ( .A(q[5]), .B(DB[222]), .Z(n8464) );
  XNOR U8409 ( .A(q[4]), .B(DB[221]), .Z(n6951) );
  IV U8410 ( .A(n6965), .Z(n8462) );
  XOR U8411 ( .A(n8465), .B(n8466), .Z(n6965) );
  XNOR U8412 ( .A(n6961), .B(n6963), .Z(n8466) );
  XNOR U8413 ( .A(q[0]), .B(DB[217]), .Z(n6963) );
  XNOR U8414 ( .A(q[3]), .B(DB[220]), .Z(n6961) );
  IV U8415 ( .A(n6960), .Z(n8465) );
  XNOR U8416 ( .A(n6958), .B(n8467), .Z(n6960) );
  XNOR U8417 ( .A(q[2]), .B(DB[219]), .Z(n8467) );
  XNOR U8418 ( .A(q[1]), .B(DB[218]), .Z(n6958) );
  XOR U8419 ( .A(n8468), .B(n6923), .Z(n6886) );
  XOR U8420 ( .A(n8469), .B(n6911), .Z(n6923) );
  XNOR U8421 ( .A(q[6]), .B(DB[230]), .Z(n6911) );
  IV U8422 ( .A(n6910), .Z(n8469) );
  XNOR U8423 ( .A(n6908), .B(n8470), .Z(n6910) );
  XNOR U8424 ( .A(q[5]), .B(DB[229]), .Z(n8470) );
  XNOR U8425 ( .A(q[4]), .B(DB[228]), .Z(n6908) );
  IV U8426 ( .A(n6922), .Z(n8468) );
  XOR U8427 ( .A(n8471), .B(n8472), .Z(n6922) );
  XNOR U8428 ( .A(n6918), .B(n6920), .Z(n8472) );
  XNOR U8429 ( .A(q[0]), .B(DB[224]), .Z(n6920) );
  XNOR U8430 ( .A(q[3]), .B(DB[227]), .Z(n6918) );
  IV U8431 ( .A(n6917), .Z(n8471) );
  XNOR U8432 ( .A(n6915), .B(n8473), .Z(n6917) );
  XNOR U8433 ( .A(q[2]), .B(DB[226]), .Z(n8473) );
  XNOR U8434 ( .A(q[1]), .B(DB[225]), .Z(n6915) );
  XOR U8435 ( .A(n8474), .B(n6880), .Z(n6843) );
  XOR U8436 ( .A(n8475), .B(n6868), .Z(n6880) );
  XNOR U8437 ( .A(q[6]), .B(DB[237]), .Z(n6868) );
  IV U8438 ( .A(n6867), .Z(n8475) );
  XNOR U8439 ( .A(n6865), .B(n8476), .Z(n6867) );
  XNOR U8440 ( .A(q[5]), .B(DB[236]), .Z(n8476) );
  XNOR U8441 ( .A(q[4]), .B(DB[235]), .Z(n6865) );
  IV U8442 ( .A(n6879), .Z(n8474) );
  XOR U8443 ( .A(n8477), .B(n8478), .Z(n6879) );
  XNOR U8444 ( .A(n6875), .B(n6877), .Z(n8478) );
  XNOR U8445 ( .A(q[0]), .B(DB[231]), .Z(n6877) );
  XNOR U8446 ( .A(q[3]), .B(DB[234]), .Z(n6875) );
  IV U8447 ( .A(n6874), .Z(n8477) );
  XNOR U8448 ( .A(n6872), .B(n8479), .Z(n6874) );
  XNOR U8449 ( .A(q[2]), .B(DB[233]), .Z(n8479) );
  XNOR U8450 ( .A(q[1]), .B(DB[232]), .Z(n6872) );
  XOR U8451 ( .A(n8480), .B(n6837), .Z(n6800) );
  XOR U8452 ( .A(n8481), .B(n6825), .Z(n6837) );
  XNOR U8453 ( .A(q[6]), .B(DB[244]), .Z(n6825) );
  IV U8454 ( .A(n6824), .Z(n8481) );
  XNOR U8455 ( .A(n6822), .B(n8482), .Z(n6824) );
  XNOR U8456 ( .A(q[5]), .B(DB[243]), .Z(n8482) );
  XNOR U8457 ( .A(q[4]), .B(DB[242]), .Z(n6822) );
  IV U8458 ( .A(n6836), .Z(n8480) );
  XOR U8459 ( .A(n8483), .B(n8484), .Z(n6836) );
  XNOR U8460 ( .A(n6832), .B(n6834), .Z(n8484) );
  XNOR U8461 ( .A(q[0]), .B(DB[238]), .Z(n6834) );
  XNOR U8462 ( .A(q[3]), .B(DB[241]), .Z(n6832) );
  IV U8463 ( .A(n6831), .Z(n8483) );
  XNOR U8464 ( .A(n6829), .B(n8485), .Z(n6831) );
  XNOR U8465 ( .A(q[2]), .B(DB[240]), .Z(n8485) );
  XNOR U8466 ( .A(q[1]), .B(DB[239]), .Z(n6829) );
  XOR U8467 ( .A(n8486), .B(n6794), .Z(n6757) );
  XOR U8468 ( .A(n8487), .B(n6782), .Z(n6794) );
  XNOR U8469 ( .A(q[6]), .B(DB[251]), .Z(n6782) );
  IV U8470 ( .A(n6781), .Z(n8487) );
  XNOR U8471 ( .A(n6779), .B(n8488), .Z(n6781) );
  XNOR U8472 ( .A(q[5]), .B(DB[250]), .Z(n8488) );
  XNOR U8473 ( .A(q[4]), .B(DB[249]), .Z(n6779) );
  IV U8474 ( .A(n6793), .Z(n8486) );
  XOR U8475 ( .A(n8489), .B(n8490), .Z(n6793) );
  XNOR U8476 ( .A(n6789), .B(n6791), .Z(n8490) );
  XNOR U8477 ( .A(q[0]), .B(DB[245]), .Z(n6791) );
  XNOR U8478 ( .A(q[3]), .B(DB[248]), .Z(n6789) );
  IV U8479 ( .A(n6788), .Z(n8489) );
  XNOR U8480 ( .A(n6786), .B(n8491), .Z(n6788) );
  XNOR U8481 ( .A(q[2]), .B(DB[247]), .Z(n8491) );
  XNOR U8482 ( .A(q[1]), .B(DB[246]), .Z(n6786) );
  XOR U8483 ( .A(n8492), .B(n6751), .Z(n6714) );
  XOR U8484 ( .A(n8493), .B(n6739), .Z(n6751) );
  XNOR U8485 ( .A(q[6]), .B(DB[258]), .Z(n6739) );
  IV U8486 ( .A(n6738), .Z(n8493) );
  XNOR U8487 ( .A(n6736), .B(n8494), .Z(n6738) );
  XNOR U8488 ( .A(q[5]), .B(DB[257]), .Z(n8494) );
  XNOR U8489 ( .A(q[4]), .B(DB[256]), .Z(n6736) );
  IV U8490 ( .A(n6750), .Z(n8492) );
  XOR U8491 ( .A(n8495), .B(n8496), .Z(n6750) );
  XNOR U8492 ( .A(n6746), .B(n6748), .Z(n8496) );
  XNOR U8493 ( .A(q[0]), .B(DB[252]), .Z(n6748) );
  XNOR U8494 ( .A(q[3]), .B(DB[255]), .Z(n6746) );
  IV U8495 ( .A(n6745), .Z(n8495) );
  XNOR U8496 ( .A(n6743), .B(n8497), .Z(n6745) );
  XNOR U8497 ( .A(q[2]), .B(DB[254]), .Z(n8497) );
  XNOR U8498 ( .A(q[1]), .B(DB[253]), .Z(n6743) );
  XOR U8499 ( .A(n8498), .B(n6708), .Z(n6671) );
  XOR U8500 ( .A(n8499), .B(n6696), .Z(n6708) );
  XNOR U8501 ( .A(q[6]), .B(DB[265]), .Z(n6696) );
  IV U8502 ( .A(n6695), .Z(n8499) );
  XNOR U8503 ( .A(n6693), .B(n8500), .Z(n6695) );
  XNOR U8504 ( .A(q[5]), .B(DB[264]), .Z(n8500) );
  XNOR U8505 ( .A(q[4]), .B(DB[263]), .Z(n6693) );
  IV U8506 ( .A(n6707), .Z(n8498) );
  XOR U8507 ( .A(n8501), .B(n8502), .Z(n6707) );
  XNOR U8508 ( .A(n6703), .B(n6705), .Z(n8502) );
  XNOR U8509 ( .A(q[0]), .B(DB[259]), .Z(n6705) );
  XNOR U8510 ( .A(q[3]), .B(DB[262]), .Z(n6703) );
  IV U8511 ( .A(n6702), .Z(n8501) );
  XNOR U8512 ( .A(n6700), .B(n8503), .Z(n6702) );
  XNOR U8513 ( .A(q[2]), .B(DB[261]), .Z(n8503) );
  XNOR U8514 ( .A(q[1]), .B(DB[260]), .Z(n6700) );
  XOR U8515 ( .A(n8504), .B(n6665), .Z(n6628) );
  XOR U8516 ( .A(n8505), .B(n6653), .Z(n6665) );
  XNOR U8517 ( .A(q[6]), .B(DB[272]), .Z(n6653) );
  IV U8518 ( .A(n6652), .Z(n8505) );
  XNOR U8519 ( .A(n6650), .B(n8506), .Z(n6652) );
  XNOR U8520 ( .A(q[5]), .B(DB[271]), .Z(n8506) );
  XNOR U8521 ( .A(q[4]), .B(DB[270]), .Z(n6650) );
  IV U8522 ( .A(n6664), .Z(n8504) );
  XOR U8523 ( .A(n8507), .B(n8508), .Z(n6664) );
  XNOR U8524 ( .A(n6660), .B(n6662), .Z(n8508) );
  XNOR U8525 ( .A(q[0]), .B(DB[266]), .Z(n6662) );
  XNOR U8526 ( .A(q[3]), .B(DB[269]), .Z(n6660) );
  IV U8527 ( .A(n6659), .Z(n8507) );
  XNOR U8528 ( .A(n6657), .B(n8509), .Z(n6659) );
  XNOR U8529 ( .A(q[2]), .B(DB[268]), .Z(n8509) );
  XNOR U8530 ( .A(q[1]), .B(DB[267]), .Z(n6657) );
  XOR U8531 ( .A(n8510), .B(n6622), .Z(n6585) );
  XOR U8532 ( .A(n8511), .B(n6610), .Z(n6622) );
  XNOR U8533 ( .A(q[6]), .B(DB[279]), .Z(n6610) );
  IV U8534 ( .A(n6609), .Z(n8511) );
  XNOR U8535 ( .A(n6607), .B(n8512), .Z(n6609) );
  XNOR U8536 ( .A(q[5]), .B(DB[278]), .Z(n8512) );
  XNOR U8537 ( .A(q[4]), .B(DB[277]), .Z(n6607) );
  IV U8538 ( .A(n6621), .Z(n8510) );
  XOR U8539 ( .A(n8513), .B(n8514), .Z(n6621) );
  XNOR U8540 ( .A(n6617), .B(n6619), .Z(n8514) );
  XNOR U8541 ( .A(q[0]), .B(DB[273]), .Z(n6619) );
  XNOR U8542 ( .A(q[3]), .B(DB[276]), .Z(n6617) );
  IV U8543 ( .A(n6616), .Z(n8513) );
  XNOR U8544 ( .A(n6614), .B(n8515), .Z(n6616) );
  XNOR U8545 ( .A(q[2]), .B(DB[275]), .Z(n8515) );
  XNOR U8546 ( .A(q[1]), .B(DB[274]), .Z(n6614) );
  XOR U8547 ( .A(n8516), .B(n6579), .Z(n6542) );
  XOR U8548 ( .A(n8517), .B(n6567), .Z(n6579) );
  XNOR U8549 ( .A(q[6]), .B(DB[286]), .Z(n6567) );
  IV U8550 ( .A(n6566), .Z(n8517) );
  XNOR U8551 ( .A(n6564), .B(n8518), .Z(n6566) );
  XNOR U8552 ( .A(q[5]), .B(DB[285]), .Z(n8518) );
  XNOR U8553 ( .A(q[4]), .B(DB[284]), .Z(n6564) );
  IV U8554 ( .A(n6578), .Z(n8516) );
  XOR U8555 ( .A(n8519), .B(n8520), .Z(n6578) );
  XNOR U8556 ( .A(n6574), .B(n6576), .Z(n8520) );
  XNOR U8557 ( .A(q[0]), .B(DB[280]), .Z(n6576) );
  XNOR U8558 ( .A(q[3]), .B(DB[283]), .Z(n6574) );
  IV U8559 ( .A(n6573), .Z(n8519) );
  XNOR U8560 ( .A(n6571), .B(n8521), .Z(n6573) );
  XNOR U8561 ( .A(q[2]), .B(DB[282]), .Z(n8521) );
  XNOR U8562 ( .A(q[1]), .B(DB[281]), .Z(n6571) );
  XOR U8563 ( .A(n8522), .B(n6536), .Z(n6499) );
  XOR U8564 ( .A(n8523), .B(n6524), .Z(n6536) );
  XNOR U8565 ( .A(q[6]), .B(DB[293]), .Z(n6524) );
  IV U8566 ( .A(n6523), .Z(n8523) );
  XNOR U8567 ( .A(n6521), .B(n8524), .Z(n6523) );
  XNOR U8568 ( .A(q[5]), .B(DB[292]), .Z(n8524) );
  XNOR U8569 ( .A(q[4]), .B(DB[291]), .Z(n6521) );
  IV U8570 ( .A(n6535), .Z(n8522) );
  XOR U8571 ( .A(n8525), .B(n8526), .Z(n6535) );
  XNOR U8572 ( .A(n6531), .B(n6533), .Z(n8526) );
  XNOR U8573 ( .A(q[0]), .B(DB[287]), .Z(n6533) );
  XNOR U8574 ( .A(q[3]), .B(DB[290]), .Z(n6531) );
  IV U8575 ( .A(n6530), .Z(n8525) );
  XNOR U8576 ( .A(n6528), .B(n8527), .Z(n6530) );
  XNOR U8577 ( .A(q[2]), .B(DB[289]), .Z(n8527) );
  XNOR U8578 ( .A(q[1]), .B(DB[288]), .Z(n6528) );
  XOR U8579 ( .A(n8528), .B(n6493), .Z(n6456) );
  XOR U8580 ( .A(n8529), .B(n6481), .Z(n6493) );
  XNOR U8581 ( .A(q[6]), .B(DB[300]), .Z(n6481) );
  IV U8582 ( .A(n6480), .Z(n8529) );
  XNOR U8583 ( .A(n6478), .B(n8530), .Z(n6480) );
  XNOR U8584 ( .A(q[5]), .B(DB[299]), .Z(n8530) );
  XNOR U8585 ( .A(q[4]), .B(DB[298]), .Z(n6478) );
  IV U8586 ( .A(n6492), .Z(n8528) );
  XOR U8587 ( .A(n8531), .B(n8532), .Z(n6492) );
  XNOR U8588 ( .A(n6488), .B(n6490), .Z(n8532) );
  XNOR U8589 ( .A(q[0]), .B(DB[294]), .Z(n6490) );
  XNOR U8590 ( .A(q[3]), .B(DB[297]), .Z(n6488) );
  IV U8591 ( .A(n6487), .Z(n8531) );
  XNOR U8592 ( .A(n6485), .B(n8533), .Z(n6487) );
  XNOR U8593 ( .A(q[2]), .B(DB[296]), .Z(n8533) );
  XNOR U8594 ( .A(q[1]), .B(DB[295]), .Z(n6485) );
  XOR U8595 ( .A(n8534), .B(n6450), .Z(n6413) );
  XOR U8596 ( .A(n8535), .B(n6438), .Z(n6450) );
  XNOR U8597 ( .A(q[6]), .B(DB[307]), .Z(n6438) );
  IV U8598 ( .A(n6437), .Z(n8535) );
  XNOR U8599 ( .A(n6435), .B(n8536), .Z(n6437) );
  XNOR U8600 ( .A(q[5]), .B(DB[306]), .Z(n8536) );
  XNOR U8601 ( .A(q[4]), .B(DB[305]), .Z(n6435) );
  IV U8602 ( .A(n6449), .Z(n8534) );
  XOR U8603 ( .A(n8537), .B(n8538), .Z(n6449) );
  XNOR U8604 ( .A(n6445), .B(n6447), .Z(n8538) );
  XNOR U8605 ( .A(q[0]), .B(DB[301]), .Z(n6447) );
  XNOR U8606 ( .A(q[3]), .B(DB[304]), .Z(n6445) );
  IV U8607 ( .A(n6444), .Z(n8537) );
  XNOR U8608 ( .A(n6442), .B(n8539), .Z(n6444) );
  XNOR U8609 ( .A(q[2]), .B(DB[303]), .Z(n8539) );
  XNOR U8610 ( .A(q[1]), .B(DB[302]), .Z(n6442) );
  XOR U8611 ( .A(n8540), .B(n6407), .Z(n6370) );
  XOR U8612 ( .A(n8541), .B(n6395), .Z(n6407) );
  XNOR U8613 ( .A(q[6]), .B(DB[314]), .Z(n6395) );
  IV U8614 ( .A(n6394), .Z(n8541) );
  XNOR U8615 ( .A(n6392), .B(n8542), .Z(n6394) );
  XNOR U8616 ( .A(q[5]), .B(DB[313]), .Z(n8542) );
  XNOR U8617 ( .A(q[4]), .B(DB[312]), .Z(n6392) );
  IV U8618 ( .A(n6406), .Z(n8540) );
  XOR U8619 ( .A(n8543), .B(n8544), .Z(n6406) );
  XNOR U8620 ( .A(n6402), .B(n6404), .Z(n8544) );
  XNOR U8621 ( .A(q[0]), .B(DB[308]), .Z(n6404) );
  XNOR U8622 ( .A(q[3]), .B(DB[311]), .Z(n6402) );
  IV U8623 ( .A(n6401), .Z(n8543) );
  XNOR U8624 ( .A(n6399), .B(n8545), .Z(n6401) );
  XNOR U8625 ( .A(q[2]), .B(DB[310]), .Z(n8545) );
  XNOR U8626 ( .A(q[1]), .B(DB[309]), .Z(n6399) );
  XOR U8627 ( .A(n8546), .B(n6364), .Z(n6327) );
  XOR U8628 ( .A(n8547), .B(n6352), .Z(n6364) );
  XNOR U8629 ( .A(q[6]), .B(DB[321]), .Z(n6352) );
  IV U8630 ( .A(n6351), .Z(n8547) );
  XNOR U8631 ( .A(n6349), .B(n8548), .Z(n6351) );
  XNOR U8632 ( .A(q[5]), .B(DB[320]), .Z(n8548) );
  XNOR U8633 ( .A(q[4]), .B(DB[319]), .Z(n6349) );
  IV U8634 ( .A(n6363), .Z(n8546) );
  XOR U8635 ( .A(n8549), .B(n8550), .Z(n6363) );
  XNOR U8636 ( .A(n6359), .B(n6361), .Z(n8550) );
  XNOR U8637 ( .A(q[0]), .B(DB[315]), .Z(n6361) );
  XNOR U8638 ( .A(q[3]), .B(DB[318]), .Z(n6359) );
  IV U8639 ( .A(n6358), .Z(n8549) );
  XNOR U8640 ( .A(n6356), .B(n8551), .Z(n6358) );
  XNOR U8641 ( .A(q[2]), .B(DB[317]), .Z(n8551) );
  XNOR U8642 ( .A(q[1]), .B(DB[316]), .Z(n6356) );
  XOR U8643 ( .A(n8552), .B(n6321), .Z(n6284) );
  XOR U8644 ( .A(n8553), .B(n6309), .Z(n6321) );
  XNOR U8645 ( .A(q[6]), .B(DB[328]), .Z(n6309) );
  IV U8646 ( .A(n6308), .Z(n8553) );
  XNOR U8647 ( .A(n6306), .B(n8554), .Z(n6308) );
  XNOR U8648 ( .A(q[5]), .B(DB[327]), .Z(n8554) );
  XNOR U8649 ( .A(q[4]), .B(DB[326]), .Z(n6306) );
  IV U8650 ( .A(n6320), .Z(n8552) );
  XOR U8651 ( .A(n8555), .B(n8556), .Z(n6320) );
  XNOR U8652 ( .A(n6316), .B(n6318), .Z(n8556) );
  XNOR U8653 ( .A(q[0]), .B(DB[322]), .Z(n6318) );
  XNOR U8654 ( .A(q[3]), .B(DB[325]), .Z(n6316) );
  IV U8655 ( .A(n6315), .Z(n8555) );
  XNOR U8656 ( .A(n6313), .B(n8557), .Z(n6315) );
  XNOR U8657 ( .A(q[2]), .B(DB[324]), .Z(n8557) );
  XNOR U8658 ( .A(q[1]), .B(DB[323]), .Z(n6313) );
  XOR U8659 ( .A(n8558), .B(n6278), .Z(n6241) );
  XOR U8660 ( .A(n8559), .B(n6266), .Z(n6278) );
  XNOR U8661 ( .A(q[6]), .B(DB[335]), .Z(n6266) );
  IV U8662 ( .A(n6265), .Z(n8559) );
  XNOR U8663 ( .A(n6263), .B(n8560), .Z(n6265) );
  XNOR U8664 ( .A(q[5]), .B(DB[334]), .Z(n8560) );
  XNOR U8665 ( .A(q[4]), .B(DB[333]), .Z(n6263) );
  IV U8666 ( .A(n6277), .Z(n8558) );
  XOR U8667 ( .A(n8561), .B(n8562), .Z(n6277) );
  XNOR U8668 ( .A(n6273), .B(n6275), .Z(n8562) );
  XNOR U8669 ( .A(q[0]), .B(DB[329]), .Z(n6275) );
  XNOR U8670 ( .A(q[3]), .B(DB[332]), .Z(n6273) );
  IV U8671 ( .A(n6272), .Z(n8561) );
  XNOR U8672 ( .A(n6270), .B(n8563), .Z(n6272) );
  XNOR U8673 ( .A(q[2]), .B(DB[331]), .Z(n8563) );
  XNOR U8674 ( .A(q[1]), .B(DB[330]), .Z(n6270) );
  XOR U8675 ( .A(n8564), .B(n6235), .Z(n6198) );
  XOR U8676 ( .A(n8565), .B(n6223), .Z(n6235) );
  XNOR U8677 ( .A(q[6]), .B(DB[342]), .Z(n6223) );
  IV U8678 ( .A(n6222), .Z(n8565) );
  XNOR U8679 ( .A(n6220), .B(n8566), .Z(n6222) );
  XNOR U8680 ( .A(q[5]), .B(DB[341]), .Z(n8566) );
  XNOR U8681 ( .A(q[4]), .B(DB[340]), .Z(n6220) );
  IV U8682 ( .A(n6234), .Z(n8564) );
  XOR U8683 ( .A(n8567), .B(n8568), .Z(n6234) );
  XNOR U8684 ( .A(n6230), .B(n6232), .Z(n8568) );
  XNOR U8685 ( .A(q[0]), .B(DB[336]), .Z(n6232) );
  XNOR U8686 ( .A(q[3]), .B(DB[339]), .Z(n6230) );
  IV U8687 ( .A(n6229), .Z(n8567) );
  XNOR U8688 ( .A(n6227), .B(n8569), .Z(n6229) );
  XNOR U8689 ( .A(q[2]), .B(DB[338]), .Z(n8569) );
  XNOR U8690 ( .A(q[1]), .B(DB[337]), .Z(n6227) );
  XOR U8691 ( .A(n8570), .B(n6192), .Z(n6155) );
  XOR U8692 ( .A(n8571), .B(n6180), .Z(n6192) );
  XNOR U8693 ( .A(q[6]), .B(DB[349]), .Z(n6180) );
  IV U8694 ( .A(n6179), .Z(n8571) );
  XNOR U8695 ( .A(n6177), .B(n8572), .Z(n6179) );
  XNOR U8696 ( .A(q[5]), .B(DB[348]), .Z(n8572) );
  XNOR U8697 ( .A(q[4]), .B(DB[347]), .Z(n6177) );
  IV U8698 ( .A(n6191), .Z(n8570) );
  XOR U8699 ( .A(n8573), .B(n8574), .Z(n6191) );
  XNOR U8700 ( .A(n6187), .B(n6189), .Z(n8574) );
  XNOR U8701 ( .A(q[0]), .B(DB[343]), .Z(n6189) );
  XNOR U8702 ( .A(q[3]), .B(DB[346]), .Z(n6187) );
  IV U8703 ( .A(n6186), .Z(n8573) );
  XNOR U8704 ( .A(n6184), .B(n8575), .Z(n6186) );
  XNOR U8705 ( .A(q[2]), .B(DB[345]), .Z(n8575) );
  XNOR U8706 ( .A(q[1]), .B(DB[344]), .Z(n6184) );
  XOR U8707 ( .A(n8576), .B(n6149), .Z(n6112) );
  XOR U8708 ( .A(n8577), .B(n6137), .Z(n6149) );
  XNOR U8709 ( .A(q[6]), .B(DB[356]), .Z(n6137) );
  IV U8710 ( .A(n6136), .Z(n8577) );
  XNOR U8711 ( .A(n6134), .B(n8578), .Z(n6136) );
  XNOR U8712 ( .A(q[5]), .B(DB[355]), .Z(n8578) );
  XNOR U8713 ( .A(q[4]), .B(DB[354]), .Z(n6134) );
  IV U8714 ( .A(n6148), .Z(n8576) );
  XOR U8715 ( .A(n8579), .B(n8580), .Z(n6148) );
  XNOR U8716 ( .A(n6144), .B(n6146), .Z(n8580) );
  XNOR U8717 ( .A(q[0]), .B(DB[350]), .Z(n6146) );
  XNOR U8718 ( .A(q[3]), .B(DB[353]), .Z(n6144) );
  IV U8719 ( .A(n6143), .Z(n8579) );
  XNOR U8720 ( .A(n6141), .B(n8581), .Z(n6143) );
  XNOR U8721 ( .A(q[2]), .B(DB[352]), .Z(n8581) );
  XNOR U8722 ( .A(q[1]), .B(DB[351]), .Z(n6141) );
  XOR U8723 ( .A(n8582), .B(n6106), .Z(n6069) );
  XOR U8724 ( .A(n8583), .B(n6094), .Z(n6106) );
  XNOR U8725 ( .A(q[6]), .B(DB[363]), .Z(n6094) );
  IV U8726 ( .A(n6093), .Z(n8583) );
  XNOR U8727 ( .A(n6091), .B(n8584), .Z(n6093) );
  XNOR U8728 ( .A(q[5]), .B(DB[362]), .Z(n8584) );
  XNOR U8729 ( .A(q[4]), .B(DB[361]), .Z(n6091) );
  IV U8730 ( .A(n6105), .Z(n8582) );
  XOR U8731 ( .A(n8585), .B(n8586), .Z(n6105) );
  XNOR U8732 ( .A(n6101), .B(n6103), .Z(n8586) );
  XNOR U8733 ( .A(q[0]), .B(DB[357]), .Z(n6103) );
  XNOR U8734 ( .A(q[3]), .B(DB[360]), .Z(n6101) );
  IV U8735 ( .A(n6100), .Z(n8585) );
  XNOR U8736 ( .A(n6098), .B(n8587), .Z(n6100) );
  XNOR U8737 ( .A(q[2]), .B(DB[359]), .Z(n8587) );
  XNOR U8738 ( .A(q[1]), .B(DB[358]), .Z(n6098) );
  XOR U8739 ( .A(n8588), .B(n6063), .Z(n6026) );
  XOR U8740 ( .A(n8589), .B(n6051), .Z(n6063) );
  XNOR U8741 ( .A(q[6]), .B(DB[370]), .Z(n6051) );
  IV U8742 ( .A(n6050), .Z(n8589) );
  XNOR U8743 ( .A(n6048), .B(n8590), .Z(n6050) );
  XNOR U8744 ( .A(q[5]), .B(DB[369]), .Z(n8590) );
  XNOR U8745 ( .A(q[4]), .B(DB[368]), .Z(n6048) );
  IV U8746 ( .A(n6062), .Z(n8588) );
  XOR U8747 ( .A(n8591), .B(n8592), .Z(n6062) );
  XNOR U8748 ( .A(n6058), .B(n6060), .Z(n8592) );
  XNOR U8749 ( .A(q[0]), .B(DB[364]), .Z(n6060) );
  XNOR U8750 ( .A(q[3]), .B(DB[367]), .Z(n6058) );
  IV U8751 ( .A(n6057), .Z(n8591) );
  XNOR U8752 ( .A(n6055), .B(n8593), .Z(n6057) );
  XNOR U8753 ( .A(q[2]), .B(DB[366]), .Z(n8593) );
  XNOR U8754 ( .A(q[1]), .B(DB[365]), .Z(n6055) );
  XOR U8755 ( .A(n8594), .B(n6020), .Z(n5983) );
  XOR U8756 ( .A(n8595), .B(n6008), .Z(n6020) );
  XNOR U8757 ( .A(q[6]), .B(DB[377]), .Z(n6008) );
  IV U8758 ( .A(n6007), .Z(n8595) );
  XNOR U8759 ( .A(n6005), .B(n8596), .Z(n6007) );
  XNOR U8760 ( .A(q[5]), .B(DB[376]), .Z(n8596) );
  XNOR U8761 ( .A(q[4]), .B(DB[375]), .Z(n6005) );
  IV U8762 ( .A(n6019), .Z(n8594) );
  XOR U8763 ( .A(n8597), .B(n8598), .Z(n6019) );
  XNOR U8764 ( .A(n6015), .B(n6017), .Z(n8598) );
  XNOR U8765 ( .A(q[0]), .B(DB[371]), .Z(n6017) );
  XNOR U8766 ( .A(q[3]), .B(DB[374]), .Z(n6015) );
  IV U8767 ( .A(n6014), .Z(n8597) );
  XNOR U8768 ( .A(n6012), .B(n8599), .Z(n6014) );
  XNOR U8769 ( .A(q[2]), .B(DB[373]), .Z(n8599) );
  XNOR U8770 ( .A(q[1]), .B(DB[372]), .Z(n6012) );
  XOR U8771 ( .A(n8600), .B(n5977), .Z(n5940) );
  XOR U8772 ( .A(n8601), .B(n5965), .Z(n5977) );
  XNOR U8773 ( .A(q[6]), .B(DB[384]), .Z(n5965) );
  IV U8774 ( .A(n5964), .Z(n8601) );
  XNOR U8775 ( .A(n5962), .B(n8602), .Z(n5964) );
  XNOR U8776 ( .A(q[5]), .B(DB[383]), .Z(n8602) );
  XNOR U8777 ( .A(q[4]), .B(DB[382]), .Z(n5962) );
  IV U8778 ( .A(n5976), .Z(n8600) );
  XOR U8779 ( .A(n8603), .B(n8604), .Z(n5976) );
  XNOR U8780 ( .A(n5972), .B(n5974), .Z(n8604) );
  XNOR U8781 ( .A(q[0]), .B(DB[378]), .Z(n5974) );
  XNOR U8782 ( .A(q[3]), .B(DB[381]), .Z(n5972) );
  IV U8783 ( .A(n5971), .Z(n8603) );
  XNOR U8784 ( .A(n5969), .B(n8605), .Z(n5971) );
  XNOR U8785 ( .A(q[2]), .B(DB[380]), .Z(n8605) );
  XNOR U8786 ( .A(q[1]), .B(DB[379]), .Z(n5969) );
  XOR U8787 ( .A(n8606), .B(n5934), .Z(n5897) );
  XOR U8788 ( .A(n8607), .B(n5922), .Z(n5934) );
  XNOR U8789 ( .A(q[6]), .B(DB[391]), .Z(n5922) );
  IV U8790 ( .A(n5921), .Z(n8607) );
  XNOR U8791 ( .A(n5919), .B(n8608), .Z(n5921) );
  XNOR U8792 ( .A(q[5]), .B(DB[390]), .Z(n8608) );
  XNOR U8793 ( .A(q[4]), .B(DB[389]), .Z(n5919) );
  IV U8794 ( .A(n5933), .Z(n8606) );
  XOR U8795 ( .A(n8609), .B(n8610), .Z(n5933) );
  XNOR U8796 ( .A(n5929), .B(n5931), .Z(n8610) );
  XNOR U8797 ( .A(q[0]), .B(DB[385]), .Z(n5931) );
  XNOR U8798 ( .A(q[3]), .B(DB[388]), .Z(n5929) );
  IV U8799 ( .A(n5928), .Z(n8609) );
  XNOR U8800 ( .A(n5926), .B(n8611), .Z(n5928) );
  XNOR U8801 ( .A(q[2]), .B(DB[387]), .Z(n8611) );
  XNOR U8802 ( .A(q[1]), .B(DB[386]), .Z(n5926) );
  XOR U8803 ( .A(n8612), .B(n5891), .Z(n5854) );
  XOR U8804 ( .A(n8613), .B(n5879), .Z(n5891) );
  XNOR U8805 ( .A(q[6]), .B(DB[398]), .Z(n5879) );
  IV U8806 ( .A(n5878), .Z(n8613) );
  XNOR U8807 ( .A(n5876), .B(n8614), .Z(n5878) );
  XNOR U8808 ( .A(q[5]), .B(DB[397]), .Z(n8614) );
  XNOR U8809 ( .A(q[4]), .B(DB[396]), .Z(n5876) );
  IV U8810 ( .A(n5890), .Z(n8612) );
  XOR U8811 ( .A(n8615), .B(n8616), .Z(n5890) );
  XNOR U8812 ( .A(n5886), .B(n5888), .Z(n8616) );
  XNOR U8813 ( .A(q[0]), .B(DB[392]), .Z(n5888) );
  XNOR U8814 ( .A(q[3]), .B(DB[395]), .Z(n5886) );
  IV U8815 ( .A(n5885), .Z(n8615) );
  XNOR U8816 ( .A(n5883), .B(n8617), .Z(n5885) );
  XNOR U8817 ( .A(q[2]), .B(DB[394]), .Z(n8617) );
  XNOR U8818 ( .A(q[1]), .B(DB[393]), .Z(n5883) );
  XOR U8819 ( .A(n8618), .B(n5848), .Z(n5811) );
  XOR U8820 ( .A(n8619), .B(n5836), .Z(n5848) );
  XNOR U8821 ( .A(q[6]), .B(DB[405]), .Z(n5836) );
  IV U8822 ( .A(n5835), .Z(n8619) );
  XNOR U8823 ( .A(n5833), .B(n8620), .Z(n5835) );
  XNOR U8824 ( .A(q[5]), .B(DB[404]), .Z(n8620) );
  XNOR U8825 ( .A(q[4]), .B(DB[403]), .Z(n5833) );
  IV U8826 ( .A(n5847), .Z(n8618) );
  XOR U8827 ( .A(n8621), .B(n8622), .Z(n5847) );
  XNOR U8828 ( .A(n5843), .B(n5845), .Z(n8622) );
  XNOR U8829 ( .A(q[0]), .B(DB[399]), .Z(n5845) );
  XNOR U8830 ( .A(q[3]), .B(DB[402]), .Z(n5843) );
  IV U8831 ( .A(n5842), .Z(n8621) );
  XNOR U8832 ( .A(n5840), .B(n8623), .Z(n5842) );
  XNOR U8833 ( .A(q[2]), .B(DB[401]), .Z(n8623) );
  XNOR U8834 ( .A(q[1]), .B(DB[400]), .Z(n5840) );
  XOR U8835 ( .A(n8624), .B(n5805), .Z(n5768) );
  XOR U8836 ( .A(n8625), .B(n5793), .Z(n5805) );
  XNOR U8837 ( .A(q[6]), .B(DB[412]), .Z(n5793) );
  IV U8838 ( .A(n5792), .Z(n8625) );
  XNOR U8839 ( .A(n5790), .B(n8626), .Z(n5792) );
  XNOR U8840 ( .A(q[5]), .B(DB[411]), .Z(n8626) );
  XNOR U8841 ( .A(q[4]), .B(DB[410]), .Z(n5790) );
  IV U8842 ( .A(n5804), .Z(n8624) );
  XOR U8843 ( .A(n8627), .B(n8628), .Z(n5804) );
  XNOR U8844 ( .A(n5800), .B(n5802), .Z(n8628) );
  XNOR U8845 ( .A(q[0]), .B(DB[406]), .Z(n5802) );
  XNOR U8846 ( .A(q[3]), .B(DB[409]), .Z(n5800) );
  IV U8847 ( .A(n5799), .Z(n8627) );
  XNOR U8848 ( .A(n5797), .B(n8629), .Z(n5799) );
  XNOR U8849 ( .A(q[2]), .B(DB[408]), .Z(n8629) );
  XNOR U8850 ( .A(q[1]), .B(DB[407]), .Z(n5797) );
  XOR U8851 ( .A(n8630), .B(n5762), .Z(n5725) );
  XOR U8852 ( .A(n8631), .B(n5750), .Z(n5762) );
  XNOR U8853 ( .A(q[6]), .B(DB[419]), .Z(n5750) );
  IV U8854 ( .A(n5749), .Z(n8631) );
  XNOR U8855 ( .A(n5747), .B(n8632), .Z(n5749) );
  XNOR U8856 ( .A(q[5]), .B(DB[418]), .Z(n8632) );
  XNOR U8857 ( .A(q[4]), .B(DB[417]), .Z(n5747) );
  IV U8858 ( .A(n5761), .Z(n8630) );
  XOR U8859 ( .A(n8633), .B(n8634), .Z(n5761) );
  XNOR U8860 ( .A(n5757), .B(n5759), .Z(n8634) );
  XNOR U8861 ( .A(q[0]), .B(DB[413]), .Z(n5759) );
  XNOR U8862 ( .A(q[3]), .B(DB[416]), .Z(n5757) );
  IV U8863 ( .A(n5756), .Z(n8633) );
  XNOR U8864 ( .A(n5754), .B(n8635), .Z(n5756) );
  XNOR U8865 ( .A(q[2]), .B(DB[415]), .Z(n8635) );
  XNOR U8866 ( .A(q[1]), .B(DB[414]), .Z(n5754) );
  XOR U8867 ( .A(n8636), .B(n5719), .Z(n5682) );
  XOR U8868 ( .A(n8637), .B(n5707), .Z(n5719) );
  XNOR U8869 ( .A(q[6]), .B(DB[426]), .Z(n5707) );
  IV U8870 ( .A(n5706), .Z(n8637) );
  XNOR U8871 ( .A(n5704), .B(n8638), .Z(n5706) );
  XNOR U8872 ( .A(q[5]), .B(DB[425]), .Z(n8638) );
  XNOR U8873 ( .A(q[4]), .B(DB[424]), .Z(n5704) );
  IV U8874 ( .A(n5718), .Z(n8636) );
  XOR U8875 ( .A(n8639), .B(n8640), .Z(n5718) );
  XNOR U8876 ( .A(n5714), .B(n5716), .Z(n8640) );
  XNOR U8877 ( .A(q[0]), .B(DB[420]), .Z(n5716) );
  XNOR U8878 ( .A(q[3]), .B(DB[423]), .Z(n5714) );
  IV U8879 ( .A(n5713), .Z(n8639) );
  XNOR U8880 ( .A(n5711), .B(n8641), .Z(n5713) );
  XNOR U8881 ( .A(q[2]), .B(DB[422]), .Z(n8641) );
  XNOR U8882 ( .A(q[1]), .B(DB[421]), .Z(n5711) );
  XOR U8883 ( .A(n8642), .B(n5676), .Z(n5639) );
  XOR U8884 ( .A(n8643), .B(n5664), .Z(n5676) );
  XNOR U8885 ( .A(q[6]), .B(DB[433]), .Z(n5664) );
  IV U8886 ( .A(n5663), .Z(n8643) );
  XNOR U8887 ( .A(n5661), .B(n8644), .Z(n5663) );
  XNOR U8888 ( .A(q[5]), .B(DB[432]), .Z(n8644) );
  XNOR U8889 ( .A(q[4]), .B(DB[431]), .Z(n5661) );
  IV U8890 ( .A(n5675), .Z(n8642) );
  XOR U8891 ( .A(n8645), .B(n8646), .Z(n5675) );
  XNOR U8892 ( .A(n5671), .B(n5673), .Z(n8646) );
  XNOR U8893 ( .A(q[0]), .B(DB[427]), .Z(n5673) );
  XNOR U8894 ( .A(q[3]), .B(DB[430]), .Z(n5671) );
  IV U8895 ( .A(n5670), .Z(n8645) );
  XNOR U8896 ( .A(n5668), .B(n8647), .Z(n5670) );
  XNOR U8897 ( .A(q[2]), .B(DB[429]), .Z(n8647) );
  XNOR U8898 ( .A(q[1]), .B(DB[428]), .Z(n5668) );
  XOR U8899 ( .A(n8648), .B(n5633), .Z(n5596) );
  XOR U8900 ( .A(n8649), .B(n5621), .Z(n5633) );
  XNOR U8901 ( .A(q[6]), .B(DB[440]), .Z(n5621) );
  IV U8902 ( .A(n5620), .Z(n8649) );
  XNOR U8903 ( .A(n5618), .B(n8650), .Z(n5620) );
  XNOR U8904 ( .A(q[5]), .B(DB[439]), .Z(n8650) );
  XNOR U8905 ( .A(q[4]), .B(DB[438]), .Z(n5618) );
  IV U8906 ( .A(n5632), .Z(n8648) );
  XOR U8907 ( .A(n8651), .B(n8652), .Z(n5632) );
  XNOR U8908 ( .A(n5628), .B(n5630), .Z(n8652) );
  XNOR U8909 ( .A(q[0]), .B(DB[434]), .Z(n5630) );
  XNOR U8910 ( .A(q[3]), .B(DB[437]), .Z(n5628) );
  IV U8911 ( .A(n5627), .Z(n8651) );
  XNOR U8912 ( .A(n5625), .B(n8653), .Z(n5627) );
  XNOR U8913 ( .A(q[2]), .B(DB[436]), .Z(n8653) );
  XNOR U8914 ( .A(q[1]), .B(DB[435]), .Z(n5625) );
  XOR U8915 ( .A(n8654), .B(n5590), .Z(n5553) );
  XOR U8916 ( .A(n8655), .B(n5578), .Z(n5590) );
  XNOR U8917 ( .A(q[6]), .B(DB[447]), .Z(n5578) );
  IV U8918 ( .A(n5577), .Z(n8655) );
  XNOR U8919 ( .A(n5575), .B(n8656), .Z(n5577) );
  XNOR U8920 ( .A(q[5]), .B(DB[446]), .Z(n8656) );
  XNOR U8921 ( .A(q[4]), .B(DB[445]), .Z(n5575) );
  IV U8922 ( .A(n5589), .Z(n8654) );
  XOR U8923 ( .A(n8657), .B(n8658), .Z(n5589) );
  XNOR U8924 ( .A(n5585), .B(n5587), .Z(n8658) );
  XNOR U8925 ( .A(q[0]), .B(DB[441]), .Z(n5587) );
  XNOR U8926 ( .A(q[3]), .B(DB[444]), .Z(n5585) );
  IV U8927 ( .A(n5584), .Z(n8657) );
  XNOR U8928 ( .A(n5582), .B(n8659), .Z(n5584) );
  XNOR U8929 ( .A(q[2]), .B(DB[443]), .Z(n8659) );
  XNOR U8930 ( .A(q[1]), .B(DB[442]), .Z(n5582) );
  XOR U8931 ( .A(n8660), .B(n5547), .Z(n5510) );
  XOR U8932 ( .A(n8661), .B(n5535), .Z(n5547) );
  XNOR U8933 ( .A(q[6]), .B(DB[454]), .Z(n5535) );
  IV U8934 ( .A(n5534), .Z(n8661) );
  XNOR U8935 ( .A(n5532), .B(n8662), .Z(n5534) );
  XNOR U8936 ( .A(q[5]), .B(DB[453]), .Z(n8662) );
  XNOR U8937 ( .A(q[4]), .B(DB[452]), .Z(n5532) );
  IV U8938 ( .A(n5546), .Z(n8660) );
  XOR U8939 ( .A(n8663), .B(n8664), .Z(n5546) );
  XNOR U8940 ( .A(n5542), .B(n5544), .Z(n8664) );
  XNOR U8941 ( .A(q[0]), .B(DB[448]), .Z(n5544) );
  XNOR U8942 ( .A(q[3]), .B(DB[451]), .Z(n5542) );
  IV U8943 ( .A(n5541), .Z(n8663) );
  XNOR U8944 ( .A(n5539), .B(n8665), .Z(n5541) );
  XNOR U8945 ( .A(q[2]), .B(DB[450]), .Z(n8665) );
  XNOR U8946 ( .A(q[1]), .B(DB[449]), .Z(n5539) );
  XOR U8947 ( .A(n8666), .B(n5504), .Z(n5467) );
  XOR U8948 ( .A(n8667), .B(n5492), .Z(n5504) );
  XNOR U8949 ( .A(q[6]), .B(DB[461]), .Z(n5492) );
  IV U8950 ( .A(n5491), .Z(n8667) );
  XNOR U8951 ( .A(n5489), .B(n8668), .Z(n5491) );
  XNOR U8952 ( .A(q[5]), .B(DB[460]), .Z(n8668) );
  XNOR U8953 ( .A(q[4]), .B(DB[459]), .Z(n5489) );
  IV U8954 ( .A(n5503), .Z(n8666) );
  XOR U8955 ( .A(n8669), .B(n8670), .Z(n5503) );
  XNOR U8956 ( .A(n5499), .B(n5501), .Z(n8670) );
  XNOR U8957 ( .A(q[0]), .B(DB[455]), .Z(n5501) );
  XNOR U8958 ( .A(q[3]), .B(DB[458]), .Z(n5499) );
  IV U8959 ( .A(n5498), .Z(n8669) );
  XNOR U8960 ( .A(n5496), .B(n8671), .Z(n5498) );
  XNOR U8961 ( .A(q[2]), .B(DB[457]), .Z(n8671) );
  XNOR U8962 ( .A(q[1]), .B(DB[456]), .Z(n5496) );
  XOR U8963 ( .A(n8672), .B(n5461), .Z(n5424) );
  XOR U8964 ( .A(n8673), .B(n5449), .Z(n5461) );
  XNOR U8965 ( .A(q[6]), .B(DB[468]), .Z(n5449) );
  IV U8966 ( .A(n5448), .Z(n8673) );
  XNOR U8967 ( .A(n5446), .B(n8674), .Z(n5448) );
  XNOR U8968 ( .A(q[5]), .B(DB[467]), .Z(n8674) );
  XNOR U8969 ( .A(q[4]), .B(DB[466]), .Z(n5446) );
  IV U8970 ( .A(n5460), .Z(n8672) );
  XOR U8971 ( .A(n8675), .B(n8676), .Z(n5460) );
  XNOR U8972 ( .A(n5456), .B(n5458), .Z(n8676) );
  XNOR U8973 ( .A(q[0]), .B(DB[462]), .Z(n5458) );
  XNOR U8974 ( .A(q[3]), .B(DB[465]), .Z(n5456) );
  IV U8975 ( .A(n5455), .Z(n8675) );
  XNOR U8976 ( .A(n5453), .B(n8677), .Z(n5455) );
  XNOR U8977 ( .A(q[2]), .B(DB[464]), .Z(n8677) );
  XNOR U8978 ( .A(q[1]), .B(DB[463]), .Z(n5453) );
  XOR U8979 ( .A(n8678), .B(n5418), .Z(n5381) );
  XOR U8980 ( .A(n8679), .B(n5406), .Z(n5418) );
  XNOR U8981 ( .A(q[6]), .B(DB[475]), .Z(n5406) );
  IV U8982 ( .A(n5405), .Z(n8679) );
  XNOR U8983 ( .A(n5403), .B(n8680), .Z(n5405) );
  XNOR U8984 ( .A(q[5]), .B(DB[474]), .Z(n8680) );
  XNOR U8985 ( .A(q[4]), .B(DB[473]), .Z(n5403) );
  IV U8986 ( .A(n5417), .Z(n8678) );
  XOR U8987 ( .A(n8681), .B(n8682), .Z(n5417) );
  XNOR U8988 ( .A(n5413), .B(n5415), .Z(n8682) );
  XNOR U8989 ( .A(q[0]), .B(DB[469]), .Z(n5415) );
  XNOR U8990 ( .A(q[3]), .B(DB[472]), .Z(n5413) );
  IV U8991 ( .A(n5412), .Z(n8681) );
  XNOR U8992 ( .A(n5410), .B(n8683), .Z(n5412) );
  XNOR U8993 ( .A(q[2]), .B(DB[471]), .Z(n8683) );
  XNOR U8994 ( .A(q[1]), .B(DB[470]), .Z(n5410) );
  XOR U8995 ( .A(n8684), .B(n5375), .Z(n5338) );
  XOR U8996 ( .A(n8685), .B(n5363), .Z(n5375) );
  XNOR U8997 ( .A(q[6]), .B(DB[482]), .Z(n5363) );
  IV U8998 ( .A(n5362), .Z(n8685) );
  XNOR U8999 ( .A(n5360), .B(n8686), .Z(n5362) );
  XNOR U9000 ( .A(q[5]), .B(DB[481]), .Z(n8686) );
  XNOR U9001 ( .A(q[4]), .B(DB[480]), .Z(n5360) );
  IV U9002 ( .A(n5374), .Z(n8684) );
  XOR U9003 ( .A(n8687), .B(n8688), .Z(n5374) );
  XNOR U9004 ( .A(n5370), .B(n5372), .Z(n8688) );
  XNOR U9005 ( .A(q[0]), .B(DB[476]), .Z(n5372) );
  XNOR U9006 ( .A(q[3]), .B(DB[479]), .Z(n5370) );
  IV U9007 ( .A(n5369), .Z(n8687) );
  XNOR U9008 ( .A(n5367), .B(n8689), .Z(n5369) );
  XNOR U9009 ( .A(q[2]), .B(DB[478]), .Z(n8689) );
  XNOR U9010 ( .A(q[1]), .B(DB[477]), .Z(n5367) );
  XOR U9011 ( .A(n8690), .B(n5332), .Z(n5295) );
  XOR U9012 ( .A(n8691), .B(n5320), .Z(n5332) );
  XNOR U9013 ( .A(q[6]), .B(DB[489]), .Z(n5320) );
  IV U9014 ( .A(n5319), .Z(n8691) );
  XNOR U9015 ( .A(n5317), .B(n8692), .Z(n5319) );
  XNOR U9016 ( .A(q[5]), .B(DB[488]), .Z(n8692) );
  XNOR U9017 ( .A(q[4]), .B(DB[487]), .Z(n5317) );
  IV U9018 ( .A(n5331), .Z(n8690) );
  XOR U9019 ( .A(n8693), .B(n8694), .Z(n5331) );
  XNOR U9020 ( .A(n5327), .B(n5329), .Z(n8694) );
  XNOR U9021 ( .A(q[0]), .B(DB[483]), .Z(n5329) );
  XNOR U9022 ( .A(q[3]), .B(DB[486]), .Z(n5327) );
  IV U9023 ( .A(n5326), .Z(n8693) );
  XNOR U9024 ( .A(n5324), .B(n8695), .Z(n5326) );
  XNOR U9025 ( .A(q[2]), .B(DB[485]), .Z(n8695) );
  XNOR U9026 ( .A(q[1]), .B(DB[484]), .Z(n5324) );
  XOR U9027 ( .A(n8696), .B(n5289), .Z(n5252) );
  XOR U9028 ( .A(n8697), .B(n5277), .Z(n5289) );
  XNOR U9029 ( .A(q[6]), .B(DB[496]), .Z(n5277) );
  IV U9030 ( .A(n5276), .Z(n8697) );
  XNOR U9031 ( .A(n5274), .B(n8698), .Z(n5276) );
  XNOR U9032 ( .A(q[5]), .B(DB[495]), .Z(n8698) );
  XNOR U9033 ( .A(q[4]), .B(DB[494]), .Z(n5274) );
  IV U9034 ( .A(n5288), .Z(n8696) );
  XOR U9035 ( .A(n8699), .B(n8700), .Z(n5288) );
  XNOR U9036 ( .A(n5284), .B(n5286), .Z(n8700) );
  XNOR U9037 ( .A(q[0]), .B(DB[490]), .Z(n5286) );
  XNOR U9038 ( .A(q[3]), .B(DB[493]), .Z(n5284) );
  IV U9039 ( .A(n5283), .Z(n8699) );
  XNOR U9040 ( .A(n5281), .B(n8701), .Z(n5283) );
  XNOR U9041 ( .A(q[2]), .B(DB[492]), .Z(n8701) );
  XNOR U9042 ( .A(q[1]), .B(DB[491]), .Z(n5281) );
  XOR U9043 ( .A(n8702), .B(n5246), .Z(n5209) );
  XOR U9044 ( .A(n8703), .B(n5234), .Z(n5246) );
  XNOR U9045 ( .A(q[6]), .B(DB[503]), .Z(n5234) );
  IV U9046 ( .A(n5233), .Z(n8703) );
  XNOR U9047 ( .A(n5231), .B(n8704), .Z(n5233) );
  XNOR U9048 ( .A(q[5]), .B(DB[502]), .Z(n8704) );
  XNOR U9049 ( .A(q[4]), .B(DB[501]), .Z(n5231) );
  IV U9050 ( .A(n5245), .Z(n8702) );
  XOR U9051 ( .A(n8705), .B(n8706), .Z(n5245) );
  XNOR U9052 ( .A(n5241), .B(n5243), .Z(n8706) );
  XNOR U9053 ( .A(q[0]), .B(DB[497]), .Z(n5243) );
  XNOR U9054 ( .A(q[3]), .B(DB[500]), .Z(n5241) );
  IV U9055 ( .A(n5240), .Z(n8705) );
  XNOR U9056 ( .A(n5238), .B(n8707), .Z(n5240) );
  XNOR U9057 ( .A(q[2]), .B(DB[499]), .Z(n8707) );
  XNOR U9058 ( .A(q[1]), .B(DB[498]), .Z(n5238) );
  XOR U9059 ( .A(n8708), .B(n5203), .Z(n5166) );
  XOR U9060 ( .A(n8709), .B(n5191), .Z(n5203) );
  XNOR U9061 ( .A(q[6]), .B(DB[510]), .Z(n5191) );
  IV U9062 ( .A(n5190), .Z(n8709) );
  XNOR U9063 ( .A(n5188), .B(n8710), .Z(n5190) );
  XNOR U9064 ( .A(q[5]), .B(DB[509]), .Z(n8710) );
  XNOR U9065 ( .A(q[4]), .B(DB[508]), .Z(n5188) );
  IV U9066 ( .A(n5202), .Z(n8708) );
  XOR U9067 ( .A(n8711), .B(n8712), .Z(n5202) );
  XNOR U9068 ( .A(n5198), .B(n5200), .Z(n8712) );
  XNOR U9069 ( .A(q[0]), .B(DB[504]), .Z(n5200) );
  XNOR U9070 ( .A(q[3]), .B(DB[507]), .Z(n5198) );
  IV U9071 ( .A(n5197), .Z(n8711) );
  XNOR U9072 ( .A(n5195), .B(n8713), .Z(n5197) );
  XNOR U9073 ( .A(q[2]), .B(DB[506]), .Z(n8713) );
  XNOR U9074 ( .A(q[1]), .B(DB[505]), .Z(n5195) );
  XOR U9075 ( .A(n8714), .B(n5160), .Z(n5123) );
  XOR U9076 ( .A(n8715), .B(n5148), .Z(n5160) );
  XNOR U9077 ( .A(q[6]), .B(DB[517]), .Z(n5148) );
  IV U9078 ( .A(n5147), .Z(n8715) );
  XNOR U9079 ( .A(n5145), .B(n8716), .Z(n5147) );
  XNOR U9080 ( .A(q[5]), .B(DB[516]), .Z(n8716) );
  XNOR U9081 ( .A(q[4]), .B(DB[515]), .Z(n5145) );
  IV U9082 ( .A(n5159), .Z(n8714) );
  XOR U9083 ( .A(n8717), .B(n8718), .Z(n5159) );
  XNOR U9084 ( .A(n5155), .B(n5157), .Z(n8718) );
  XNOR U9085 ( .A(q[0]), .B(DB[511]), .Z(n5157) );
  XNOR U9086 ( .A(q[3]), .B(DB[514]), .Z(n5155) );
  IV U9087 ( .A(n5154), .Z(n8717) );
  XNOR U9088 ( .A(n5152), .B(n8719), .Z(n5154) );
  XNOR U9089 ( .A(q[2]), .B(DB[513]), .Z(n8719) );
  XNOR U9090 ( .A(q[1]), .B(DB[512]), .Z(n5152) );
  XOR U9091 ( .A(n8720), .B(n5117), .Z(n5080) );
  XOR U9092 ( .A(n8721), .B(n5105), .Z(n5117) );
  XNOR U9093 ( .A(q[6]), .B(DB[524]), .Z(n5105) );
  IV U9094 ( .A(n5104), .Z(n8721) );
  XNOR U9095 ( .A(n5102), .B(n8722), .Z(n5104) );
  XNOR U9096 ( .A(q[5]), .B(DB[523]), .Z(n8722) );
  XNOR U9097 ( .A(q[4]), .B(DB[522]), .Z(n5102) );
  IV U9098 ( .A(n5116), .Z(n8720) );
  XOR U9099 ( .A(n8723), .B(n8724), .Z(n5116) );
  XNOR U9100 ( .A(n5112), .B(n5114), .Z(n8724) );
  XNOR U9101 ( .A(q[0]), .B(DB[518]), .Z(n5114) );
  XNOR U9102 ( .A(q[3]), .B(DB[521]), .Z(n5112) );
  IV U9103 ( .A(n5111), .Z(n8723) );
  XNOR U9104 ( .A(n5109), .B(n8725), .Z(n5111) );
  XNOR U9105 ( .A(q[2]), .B(DB[520]), .Z(n8725) );
  XNOR U9106 ( .A(q[1]), .B(DB[519]), .Z(n5109) );
  XOR U9107 ( .A(n8726), .B(n5074), .Z(n5037) );
  XOR U9108 ( .A(n8727), .B(n5062), .Z(n5074) );
  XNOR U9109 ( .A(q[6]), .B(DB[531]), .Z(n5062) );
  IV U9110 ( .A(n5061), .Z(n8727) );
  XNOR U9111 ( .A(n5059), .B(n8728), .Z(n5061) );
  XNOR U9112 ( .A(q[5]), .B(DB[530]), .Z(n8728) );
  XNOR U9113 ( .A(q[4]), .B(DB[529]), .Z(n5059) );
  IV U9114 ( .A(n5073), .Z(n8726) );
  XOR U9115 ( .A(n8729), .B(n8730), .Z(n5073) );
  XNOR U9116 ( .A(n5069), .B(n5071), .Z(n8730) );
  XNOR U9117 ( .A(q[0]), .B(DB[525]), .Z(n5071) );
  XNOR U9118 ( .A(q[3]), .B(DB[528]), .Z(n5069) );
  IV U9119 ( .A(n5068), .Z(n8729) );
  XNOR U9120 ( .A(n5066), .B(n8731), .Z(n5068) );
  XNOR U9121 ( .A(q[2]), .B(DB[527]), .Z(n8731) );
  XNOR U9122 ( .A(q[1]), .B(DB[526]), .Z(n5066) );
  XOR U9123 ( .A(n8732), .B(n5031), .Z(n4994) );
  XOR U9124 ( .A(n8733), .B(n5019), .Z(n5031) );
  XNOR U9125 ( .A(q[6]), .B(DB[538]), .Z(n5019) );
  IV U9126 ( .A(n5018), .Z(n8733) );
  XNOR U9127 ( .A(n5016), .B(n8734), .Z(n5018) );
  XNOR U9128 ( .A(q[5]), .B(DB[537]), .Z(n8734) );
  XNOR U9129 ( .A(q[4]), .B(DB[536]), .Z(n5016) );
  IV U9130 ( .A(n5030), .Z(n8732) );
  XOR U9131 ( .A(n8735), .B(n8736), .Z(n5030) );
  XNOR U9132 ( .A(n5026), .B(n5028), .Z(n8736) );
  XNOR U9133 ( .A(q[0]), .B(DB[532]), .Z(n5028) );
  XNOR U9134 ( .A(q[3]), .B(DB[535]), .Z(n5026) );
  IV U9135 ( .A(n5025), .Z(n8735) );
  XNOR U9136 ( .A(n5023), .B(n8737), .Z(n5025) );
  XNOR U9137 ( .A(q[2]), .B(DB[534]), .Z(n8737) );
  XNOR U9138 ( .A(q[1]), .B(DB[533]), .Z(n5023) );
  XOR U9139 ( .A(n8738), .B(n4988), .Z(n4951) );
  XOR U9140 ( .A(n8739), .B(n4976), .Z(n4988) );
  XNOR U9141 ( .A(q[6]), .B(DB[545]), .Z(n4976) );
  IV U9142 ( .A(n4975), .Z(n8739) );
  XNOR U9143 ( .A(n4973), .B(n8740), .Z(n4975) );
  XNOR U9144 ( .A(q[5]), .B(DB[544]), .Z(n8740) );
  XNOR U9145 ( .A(q[4]), .B(DB[543]), .Z(n4973) );
  IV U9146 ( .A(n4987), .Z(n8738) );
  XOR U9147 ( .A(n8741), .B(n8742), .Z(n4987) );
  XNOR U9148 ( .A(n4983), .B(n4985), .Z(n8742) );
  XNOR U9149 ( .A(q[0]), .B(DB[539]), .Z(n4985) );
  XNOR U9150 ( .A(q[3]), .B(DB[542]), .Z(n4983) );
  IV U9151 ( .A(n4982), .Z(n8741) );
  XNOR U9152 ( .A(n4980), .B(n8743), .Z(n4982) );
  XNOR U9153 ( .A(q[2]), .B(DB[541]), .Z(n8743) );
  XNOR U9154 ( .A(q[1]), .B(DB[540]), .Z(n4980) );
  XOR U9155 ( .A(n8744), .B(n4945), .Z(n4908) );
  XOR U9156 ( .A(n8745), .B(n4933), .Z(n4945) );
  XNOR U9157 ( .A(q[6]), .B(DB[552]), .Z(n4933) );
  IV U9158 ( .A(n4932), .Z(n8745) );
  XNOR U9159 ( .A(n4930), .B(n8746), .Z(n4932) );
  XNOR U9160 ( .A(q[5]), .B(DB[551]), .Z(n8746) );
  XNOR U9161 ( .A(q[4]), .B(DB[550]), .Z(n4930) );
  IV U9162 ( .A(n4944), .Z(n8744) );
  XOR U9163 ( .A(n8747), .B(n8748), .Z(n4944) );
  XNOR U9164 ( .A(n4940), .B(n4942), .Z(n8748) );
  XNOR U9165 ( .A(q[0]), .B(DB[546]), .Z(n4942) );
  XNOR U9166 ( .A(q[3]), .B(DB[549]), .Z(n4940) );
  IV U9167 ( .A(n4939), .Z(n8747) );
  XNOR U9168 ( .A(n4937), .B(n8749), .Z(n4939) );
  XNOR U9169 ( .A(q[2]), .B(DB[548]), .Z(n8749) );
  XNOR U9170 ( .A(q[1]), .B(DB[547]), .Z(n4937) );
  XOR U9171 ( .A(n8750), .B(n4902), .Z(n4865) );
  XOR U9172 ( .A(n8751), .B(n4890), .Z(n4902) );
  XNOR U9173 ( .A(q[6]), .B(DB[559]), .Z(n4890) );
  IV U9174 ( .A(n4889), .Z(n8751) );
  XNOR U9175 ( .A(n4887), .B(n8752), .Z(n4889) );
  XNOR U9176 ( .A(q[5]), .B(DB[558]), .Z(n8752) );
  XNOR U9177 ( .A(q[4]), .B(DB[557]), .Z(n4887) );
  IV U9178 ( .A(n4901), .Z(n8750) );
  XOR U9179 ( .A(n8753), .B(n8754), .Z(n4901) );
  XNOR U9180 ( .A(n4897), .B(n4899), .Z(n8754) );
  XNOR U9181 ( .A(q[0]), .B(DB[553]), .Z(n4899) );
  XNOR U9182 ( .A(q[3]), .B(DB[556]), .Z(n4897) );
  IV U9183 ( .A(n4896), .Z(n8753) );
  XNOR U9184 ( .A(n4894), .B(n8755), .Z(n4896) );
  XNOR U9185 ( .A(q[2]), .B(DB[555]), .Z(n8755) );
  XNOR U9186 ( .A(q[1]), .B(DB[554]), .Z(n4894) );
  XOR U9187 ( .A(n8756), .B(n4859), .Z(n4822) );
  XOR U9188 ( .A(n8757), .B(n4847), .Z(n4859) );
  XNOR U9189 ( .A(q[6]), .B(DB[566]), .Z(n4847) );
  IV U9190 ( .A(n4846), .Z(n8757) );
  XNOR U9191 ( .A(n4844), .B(n8758), .Z(n4846) );
  XNOR U9192 ( .A(q[5]), .B(DB[565]), .Z(n8758) );
  XNOR U9193 ( .A(q[4]), .B(DB[564]), .Z(n4844) );
  IV U9194 ( .A(n4858), .Z(n8756) );
  XOR U9195 ( .A(n8759), .B(n8760), .Z(n4858) );
  XNOR U9196 ( .A(n4854), .B(n4856), .Z(n8760) );
  XNOR U9197 ( .A(q[0]), .B(DB[560]), .Z(n4856) );
  XNOR U9198 ( .A(q[3]), .B(DB[563]), .Z(n4854) );
  IV U9199 ( .A(n4853), .Z(n8759) );
  XNOR U9200 ( .A(n4851), .B(n8761), .Z(n4853) );
  XNOR U9201 ( .A(q[2]), .B(DB[562]), .Z(n8761) );
  XNOR U9202 ( .A(q[1]), .B(DB[561]), .Z(n4851) );
  XOR U9203 ( .A(n8762), .B(n4816), .Z(n4779) );
  XOR U9204 ( .A(n8763), .B(n4804), .Z(n4816) );
  XNOR U9205 ( .A(q[6]), .B(DB[573]), .Z(n4804) );
  IV U9206 ( .A(n4803), .Z(n8763) );
  XNOR U9207 ( .A(n4801), .B(n8764), .Z(n4803) );
  XNOR U9208 ( .A(q[5]), .B(DB[572]), .Z(n8764) );
  XNOR U9209 ( .A(q[4]), .B(DB[571]), .Z(n4801) );
  IV U9210 ( .A(n4815), .Z(n8762) );
  XOR U9211 ( .A(n8765), .B(n8766), .Z(n4815) );
  XNOR U9212 ( .A(n4811), .B(n4813), .Z(n8766) );
  XNOR U9213 ( .A(q[0]), .B(DB[567]), .Z(n4813) );
  XNOR U9214 ( .A(q[3]), .B(DB[570]), .Z(n4811) );
  IV U9215 ( .A(n4810), .Z(n8765) );
  XNOR U9216 ( .A(n4808), .B(n8767), .Z(n4810) );
  XNOR U9217 ( .A(q[2]), .B(DB[569]), .Z(n8767) );
  XNOR U9218 ( .A(q[1]), .B(DB[568]), .Z(n4808) );
  XOR U9219 ( .A(n8768), .B(n4773), .Z(n4736) );
  XOR U9220 ( .A(n8769), .B(n4761), .Z(n4773) );
  XNOR U9221 ( .A(q[6]), .B(DB[580]), .Z(n4761) );
  IV U9222 ( .A(n4760), .Z(n8769) );
  XNOR U9223 ( .A(n4758), .B(n8770), .Z(n4760) );
  XNOR U9224 ( .A(q[5]), .B(DB[579]), .Z(n8770) );
  XNOR U9225 ( .A(q[4]), .B(DB[578]), .Z(n4758) );
  IV U9226 ( .A(n4772), .Z(n8768) );
  XOR U9227 ( .A(n8771), .B(n8772), .Z(n4772) );
  XNOR U9228 ( .A(n4768), .B(n4770), .Z(n8772) );
  XNOR U9229 ( .A(q[0]), .B(DB[574]), .Z(n4770) );
  XNOR U9230 ( .A(q[3]), .B(DB[577]), .Z(n4768) );
  IV U9231 ( .A(n4767), .Z(n8771) );
  XNOR U9232 ( .A(n4765), .B(n8773), .Z(n4767) );
  XNOR U9233 ( .A(q[2]), .B(DB[576]), .Z(n8773) );
  XNOR U9234 ( .A(q[1]), .B(DB[575]), .Z(n4765) );
  XOR U9235 ( .A(n8774), .B(n4730), .Z(n4693) );
  XOR U9236 ( .A(n8775), .B(n4718), .Z(n4730) );
  XNOR U9237 ( .A(q[6]), .B(DB[587]), .Z(n4718) );
  IV U9238 ( .A(n4717), .Z(n8775) );
  XNOR U9239 ( .A(n4715), .B(n8776), .Z(n4717) );
  XNOR U9240 ( .A(q[5]), .B(DB[586]), .Z(n8776) );
  XNOR U9241 ( .A(q[4]), .B(DB[585]), .Z(n4715) );
  IV U9242 ( .A(n4729), .Z(n8774) );
  XOR U9243 ( .A(n8777), .B(n8778), .Z(n4729) );
  XNOR U9244 ( .A(n4725), .B(n4727), .Z(n8778) );
  XNOR U9245 ( .A(q[0]), .B(DB[581]), .Z(n4727) );
  XNOR U9246 ( .A(q[3]), .B(DB[584]), .Z(n4725) );
  IV U9247 ( .A(n4724), .Z(n8777) );
  XNOR U9248 ( .A(n4722), .B(n8779), .Z(n4724) );
  XNOR U9249 ( .A(q[2]), .B(DB[583]), .Z(n8779) );
  XNOR U9250 ( .A(q[1]), .B(DB[582]), .Z(n4722) );
  XOR U9251 ( .A(n8780), .B(n4687), .Z(n4650) );
  XOR U9252 ( .A(n8781), .B(n4675), .Z(n4687) );
  XNOR U9253 ( .A(q[6]), .B(DB[594]), .Z(n4675) );
  IV U9254 ( .A(n4674), .Z(n8781) );
  XNOR U9255 ( .A(n4672), .B(n8782), .Z(n4674) );
  XNOR U9256 ( .A(q[5]), .B(DB[593]), .Z(n8782) );
  XNOR U9257 ( .A(q[4]), .B(DB[592]), .Z(n4672) );
  IV U9258 ( .A(n4686), .Z(n8780) );
  XOR U9259 ( .A(n8783), .B(n8784), .Z(n4686) );
  XNOR U9260 ( .A(n4682), .B(n4684), .Z(n8784) );
  XNOR U9261 ( .A(q[0]), .B(DB[588]), .Z(n4684) );
  XNOR U9262 ( .A(q[3]), .B(DB[591]), .Z(n4682) );
  IV U9263 ( .A(n4681), .Z(n8783) );
  XNOR U9264 ( .A(n4679), .B(n8785), .Z(n4681) );
  XNOR U9265 ( .A(q[2]), .B(DB[590]), .Z(n8785) );
  XNOR U9266 ( .A(q[1]), .B(DB[589]), .Z(n4679) );
  XOR U9267 ( .A(n8786), .B(n4644), .Z(n4607) );
  XOR U9268 ( .A(n8787), .B(n4632), .Z(n4644) );
  XNOR U9269 ( .A(q[6]), .B(DB[601]), .Z(n4632) );
  IV U9270 ( .A(n4631), .Z(n8787) );
  XNOR U9271 ( .A(n4629), .B(n8788), .Z(n4631) );
  XNOR U9272 ( .A(q[5]), .B(DB[600]), .Z(n8788) );
  XNOR U9273 ( .A(q[4]), .B(DB[599]), .Z(n4629) );
  IV U9274 ( .A(n4643), .Z(n8786) );
  XOR U9275 ( .A(n8789), .B(n8790), .Z(n4643) );
  XNOR U9276 ( .A(n4639), .B(n4641), .Z(n8790) );
  XNOR U9277 ( .A(q[0]), .B(DB[595]), .Z(n4641) );
  XNOR U9278 ( .A(q[3]), .B(DB[598]), .Z(n4639) );
  IV U9279 ( .A(n4638), .Z(n8789) );
  XNOR U9280 ( .A(n4636), .B(n8791), .Z(n4638) );
  XNOR U9281 ( .A(q[2]), .B(DB[597]), .Z(n8791) );
  XNOR U9282 ( .A(q[1]), .B(DB[596]), .Z(n4636) );
  XOR U9283 ( .A(n8792), .B(n4601), .Z(n4564) );
  XOR U9284 ( .A(n8793), .B(n4589), .Z(n4601) );
  XNOR U9285 ( .A(q[6]), .B(DB[608]), .Z(n4589) );
  IV U9286 ( .A(n4588), .Z(n8793) );
  XNOR U9287 ( .A(n4586), .B(n8794), .Z(n4588) );
  XNOR U9288 ( .A(q[5]), .B(DB[607]), .Z(n8794) );
  XNOR U9289 ( .A(q[4]), .B(DB[606]), .Z(n4586) );
  IV U9290 ( .A(n4600), .Z(n8792) );
  XOR U9291 ( .A(n8795), .B(n8796), .Z(n4600) );
  XNOR U9292 ( .A(n4596), .B(n4598), .Z(n8796) );
  XNOR U9293 ( .A(q[0]), .B(DB[602]), .Z(n4598) );
  XNOR U9294 ( .A(q[3]), .B(DB[605]), .Z(n4596) );
  IV U9295 ( .A(n4595), .Z(n8795) );
  XNOR U9296 ( .A(n4593), .B(n8797), .Z(n4595) );
  XNOR U9297 ( .A(q[2]), .B(DB[604]), .Z(n8797) );
  XNOR U9298 ( .A(q[1]), .B(DB[603]), .Z(n4593) );
  XOR U9299 ( .A(n8798), .B(n4558), .Z(n4521) );
  XOR U9300 ( .A(n8799), .B(n4546), .Z(n4558) );
  XNOR U9301 ( .A(q[6]), .B(DB[615]), .Z(n4546) );
  IV U9302 ( .A(n4545), .Z(n8799) );
  XNOR U9303 ( .A(n4543), .B(n8800), .Z(n4545) );
  XNOR U9304 ( .A(q[5]), .B(DB[614]), .Z(n8800) );
  XNOR U9305 ( .A(q[4]), .B(DB[613]), .Z(n4543) );
  IV U9306 ( .A(n4557), .Z(n8798) );
  XOR U9307 ( .A(n8801), .B(n8802), .Z(n4557) );
  XNOR U9308 ( .A(n4553), .B(n4555), .Z(n8802) );
  XNOR U9309 ( .A(q[0]), .B(DB[609]), .Z(n4555) );
  XNOR U9310 ( .A(q[3]), .B(DB[612]), .Z(n4553) );
  IV U9311 ( .A(n4552), .Z(n8801) );
  XNOR U9312 ( .A(n4550), .B(n8803), .Z(n4552) );
  XNOR U9313 ( .A(q[2]), .B(DB[611]), .Z(n8803) );
  XNOR U9314 ( .A(q[1]), .B(DB[610]), .Z(n4550) );
  XOR U9315 ( .A(n8804), .B(n4515), .Z(n4478) );
  XOR U9316 ( .A(n8805), .B(n4503), .Z(n4515) );
  XNOR U9317 ( .A(q[6]), .B(DB[622]), .Z(n4503) );
  IV U9318 ( .A(n4502), .Z(n8805) );
  XNOR U9319 ( .A(n4500), .B(n8806), .Z(n4502) );
  XNOR U9320 ( .A(q[5]), .B(DB[621]), .Z(n8806) );
  XNOR U9321 ( .A(q[4]), .B(DB[620]), .Z(n4500) );
  IV U9322 ( .A(n4514), .Z(n8804) );
  XOR U9323 ( .A(n8807), .B(n8808), .Z(n4514) );
  XNOR U9324 ( .A(n4510), .B(n4512), .Z(n8808) );
  XNOR U9325 ( .A(q[0]), .B(DB[616]), .Z(n4512) );
  XNOR U9326 ( .A(q[3]), .B(DB[619]), .Z(n4510) );
  IV U9327 ( .A(n4509), .Z(n8807) );
  XNOR U9328 ( .A(n4507), .B(n8809), .Z(n4509) );
  XNOR U9329 ( .A(q[2]), .B(DB[618]), .Z(n8809) );
  XNOR U9330 ( .A(q[1]), .B(DB[617]), .Z(n4507) );
  XOR U9331 ( .A(n8810), .B(n4472), .Z(n4435) );
  XOR U9332 ( .A(n8811), .B(n4460), .Z(n4472) );
  XNOR U9333 ( .A(q[6]), .B(DB[629]), .Z(n4460) );
  IV U9334 ( .A(n4459), .Z(n8811) );
  XNOR U9335 ( .A(n4457), .B(n8812), .Z(n4459) );
  XNOR U9336 ( .A(q[5]), .B(DB[628]), .Z(n8812) );
  XNOR U9337 ( .A(q[4]), .B(DB[627]), .Z(n4457) );
  IV U9338 ( .A(n4471), .Z(n8810) );
  XOR U9339 ( .A(n8813), .B(n8814), .Z(n4471) );
  XNOR U9340 ( .A(n4467), .B(n4469), .Z(n8814) );
  XNOR U9341 ( .A(q[0]), .B(DB[623]), .Z(n4469) );
  XNOR U9342 ( .A(q[3]), .B(DB[626]), .Z(n4467) );
  IV U9343 ( .A(n4466), .Z(n8813) );
  XNOR U9344 ( .A(n4464), .B(n8815), .Z(n4466) );
  XNOR U9345 ( .A(q[2]), .B(DB[625]), .Z(n8815) );
  XNOR U9346 ( .A(q[1]), .B(DB[624]), .Z(n4464) );
  XOR U9347 ( .A(n8816), .B(n4429), .Z(n4392) );
  XOR U9348 ( .A(n8817), .B(n4417), .Z(n4429) );
  XNOR U9349 ( .A(q[6]), .B(DB[636]), .Z(n4417) );
  IV U9350 ( .A(n4416), .Z(n8817) );
  XNOR U9351 ( .A(n4414), .B(n8818), .Z(n4416) );
  XNOR U9352 ( .A(q[5]), .B(DB[635]), .Z(n8818) );
  XNOR U9353 ( .A(q[4]), .B(DB[634]), .Z(n4414) );
  IV U9354 ( .A(n4428), .Z(n8816) );
  XOR U9355 ( .A(n8819), .B(n8820), .Z(n4428) );
  XNOR U9356 ( .A(n4424), .B(n4426), .Z(n8820) );
  XNOR U9357 ( .A(q[0]), .B(DB[630]), .Z(n4426) );
  XNOR U9358 ( .A(q[3]), .B(DB[633]), .Z(n4424) );
  IV U9359 ( .A(n4423), .Z(n8819) );
  XNOR U9360 ( .A(n4421), .B(n8821), .Z(n4423) );
  XNOR U9361 ( .A(q[2]), .B(DB[632]), .Z(n8821) );
  XNOR U9362 ( .A(q[1]), .B(DB[631]), .Z(n4421) );
  XOR U9363 ( .A(n8822), .B(n4386), .Z(n4349) );
  XOR U9364 ( .A(n8823), .B(n4374), .Z(n4386) );
  XNOR U9365 ( .A(q[6]), .B(DB[643]), .Z(n4374) );
  IV U9366 ( .A(n4373), .Z(n8823) );
  XNOR U9367 ( .A(n4371), .B(n8824), .Z(n4373) );
  XNOR U9368 ( .A(q[5]), .B(DB[642]), .Z(n8824) );
  XNOR U9369 ( .A(q[4]), .B(DB[641]), .Z(n4371) );
  IV U9370 ( .A(n4385), .Z(n8822) );
  XOR U9371 ( .A(n8825), .B(n8826), .Z(n4385) );
  XNOR U9372 ( .A(n4381), .B(n4383), .Z(n8826) );
  XNOR U9373 ( .A(q[0]), .B(DB[637]), .Z(n4383) );
  XNOR U9374 ( .A(q[3]), .B(DB[640]), .Z(n4381) );
  IV U9375 ( .A(n4380), .Z(n8825) );
  XNOR U9376 ( .A(n4378), .B(n8827), .Z(n4380) );
  XNOR U9377 ( .A(q[2]), .B(DB[639]), .Z(n8827) );
  XNOR U9378 ( .A(q[1]), .B(DB[638]), .Z(n4378) );
  XOR U9379 ( .A(n8828), .B(n4343), .Z(n4306) );
  XOR U9380 ( .A(n8829), .B(n4331), .Z(n4343) );
  XNOR U9381 ( .A(q[6]), .B(DB[650]), .Z(n4331) );
  IV U9382 ( .A(n4330), .Z(n8829) );
  XNOR U9383 ( .A(n4328), .B(n8830), .Z(n4330) );
  XNOR U9384 ( .A(q[5]), .B(DB[649]), .Z(n8830) );
  XNOR U9385 ( .A(q[4]), .B(DB[648]), .Z(n4328) );
  IV U9386 ( .A(n4342), .Z(n8828) );
  XOR U9387 ( .A(n8831), .B(n8832), .Z(n4342) );
  XNOR U9388 ( .A(n4338), .B(n4340), .Z(n8832) );
  XNOR U9389 ( .A(q[0]), .B(DB[644]), .Z(n4340) );
  XNOR U9390 ( .A(q[3]), .B(DB[647]), .Z(n4338) );
  IV U9391 ( .A(n4337), .Z(n8831) );
  XNOR U9392 ( .A(n4335), .B(n8833), .Z(n4337) );
  XNOR U9393 ( .A(q[2]), .B(DB[646]), .Z(n8833) );
  XNOR U9394 ( .A(q[1]), .B(DB[645]), .Z(n4335) );
  XOR U9395 ( .A(n8834), .B(n4300), .Z(n4263) );
  XOR U9396 ( .A(n8835), .B(n4288), .Z(n4300) );
  XNOR U9397 ( .A(q[6]), .B(DB[657]), .Z(n4288) );
  IV U9398 ( .A(n4287), .Z(n8835) );
  XNOR U9399 ( .A(n4285), .B(n8836), .Z(n4287) );
  XNOR U9400 ( .A(q[5]), .B(DB[656]), .Z(n8836) );
  XNOR U9401 ( .A(q[4]), .B(DB[655]), .Z(n4285) );
  IV U9402 ( .A(n4299), .Z(n8834) );
  XOR U9403 ( .A(n8837), .B(n8838), .Z(n4299) );
  XNOR U9404 ( .A(n4295), .B(n4297), .Z(n8838) );
  XNOR U9405 ( .A(q[0]), .B(DB[651]), .Z(n4297) );
  XNOR U9406 ( .A(q[3]), .B(DB[654]), .Z(n4295) );
  IV U9407 ( .A(n4294), .Z(n8837) );
  XNOR U9408 ( .A(n4292), .B(n8839), .Z(n4294) );
  XNOR U9409 ( .A(q[2]), .B(DB[653]), .Z(n8839) );
  XNOR U9410 ( .A(q[1]), .B(DB[652]), .Z(n4292) );
  XOR U9411 ( .A(n8840), .B(n4257), .Z(n4220) );
  XOR U9412 ( .A(n8841), .B(n4245), .Z(n4257) );
  XNOR U9413 ( .A(q[6]), .B(DB[664]), .Z(n4245) );
  IV U9414 ( .A(n4244), .Z(n8841) );
  XNOR U9415 ( .A(n4242), .B(n8842), .Z(n4244) );
  XNOR U9416 ( .A(q[5]), .B(DB[663]), .Z(n8842) );
  XNOR U9417 ( .A(q[4]), .B(DB[662]), .Z(n4242) );
  IV U9418 ( .A(n4256), .Z(n8840) );
  XOR U9419 ( .A(n8843), .B(n8844), .Z(n4256) );
  XNOR U9420 ( .A(n4252), .B(n4254), .Z(n8844) );
  XNOR U9421 ( .A(q[0]), .B(DB[658]), .Z(n4254) );
  XNOR U9422 ( .A(q[3]), .B(DB[661]), .Z(n4252) );
  IV U9423 ( .A(n4251), .Z(n8843) );
  XNOR U9424 ( .A(n4249), .B(n8845), .Z(n4251) );
  XNOR U9425 ( .A(q[2]), .B(DB[660]), .Z(n8845) );
  XNOR U9426 ( .A(q[1]), .B(DB[659]), .Z(n4249) );
  XOR U9427 ( .A(n8846), .B(n4214), .Z(n4177) );
  XOR U9428 ( .A(n8847), .B(n4202), .Z(n4214) );
  XNOR U9429 ( .A(q[6]), .B(DB[671]), .Z(n4202) );
  IV U9430 ( .A(n4201), .Z(n8847) );
  XNOR U9431 ( .A(n4199), .B(n8848), .Z(n4201) );
  XNOR U9432 ( .A(q[5]), .B(DB[670]), .Z(n8848) );
  XNOR U9433 ( .A(q[4]), .B(DB[669]), .Z(n4199) );
  IV U9434 ( .A(n4213), .Z(n8846) );
  XOR U9435 ( .A(n8849), .B(n8850), .Z(n4213) );
  XNOR U9436 ( .A(n4209), .B(n4211), .Z(n8850) );
  XNOR U9437 ( .A(q[0]), .B(DB[665]), .Z(n4211) );
  XNOR U9438 ( .A(q[3]), .B(DB[668]), .Z(n4209) );
  IV U9439 ( .A(n4208), .Z(n8849) );
  XNOR U9440 ( .A(n4206), .B(n8851), .Z(n4208) );
  XNOR U9441 ( .A(q[2]), .B(DB[667]), .Z(n8851) );
  XNOR U9442 ( .A(q[1]), .B(DB[666]), .Z(n4206) );
  XOR U9443 ( .A(n8852), .B(n4171), .Z(n4134) );
  XOR U9444 ( .A(n8853), .B(n4159), .Z(n4171) );
  XNOR U9445 ( .A(q[6]), .B(DB[678]), .Z(n4159) );
  IV U9446 ( .A(n4158), .Z(n8853) );
  XNOR U9447 ( .A(n4156), .B(n8854), .Z(n4158) );
  XNOR U9448 ( .A(q[5]), .B(DB[677]), .Z(n8854) );
  XNOR U9449 ( .A(q[4]), .B(DB[676]), .Z(n4156) );
  IV U9450 ( .A(n4170), .Z(n8852) );
  XOR U9451 ( .A(n8855), .B(n8856), .Z(n4170) );
  XNOR U9452 ( .A(n4166), .B(n4168), .Z(n8856) );
  XNOR U9453 ( .A(q[0]), .B(DB[672]), .Z(n4168) );
  XNOR U9454 ( .A(q[3]), .B(DB[675]), .Z(n4166) );
  IV U9455 ( .A(n4165), .Z(n8855) );
  XNOR U9456 ( .A(n4163), .B(n8857), .Z(n4165) );
  XNOR U9457 ( .A(q[2]), .B(DB[674]), .Z(n8857) );
  XNOR U9458 ( .A(q[1]), .B(DB[673]), .Z(n4163) );
  XOR U9459 ( .A(n8858), .B(n4128), .Z(n4091) );
  XOR U9460 ( .A(n8859), .B(n4116), .Z(n4128) );
  XNOR U9461 ( .A(q[6]), .B(DB[685]), .Z(n4116) );
  IV U9462 ( .A(n4115), .Z(n8859) );
  XNOR U9463 ( .A(n4113), .B(n8860), .Z(n4115) );
  XNOR U9464 ( .A(q[5]), .B(DB[684]), .Z(n8860) );
  XNOR U9465 ( .A(q[4]), .B(DB[683]), .Z(n4113) );
  IV U9466 ( .A(n4127), .Z(n8858) );
  XOR U9467 ( .A(n8861), .B(n8862), .Z(n4127) );
  XNOR U9468 ( .A(n4123), .B(n4125), .Z(n8862) );
  XNOR U9469 ( .A(q[0]), .B(DB[679]), .Z(n4125) );
  XNOR U9470 ( .A(q[3]), .B(DB[682]), .Z(n4123) );
  IV U9471 ( .A(n4122), .Z(n8861) );
  XNOR U9472 ( .A(n4120), .B(n8863), .Z(n4122) );
  XNOR U9473 ( .A(q[2]), .B(DB[681]), .Z(n8863) );
  XNOR U9474 ( .A(q[1]), .B(DB[680]), .Z(n4120) );
  XOR U9475 ( .A(n8864), .B(n4085), .Z(n4048) );
  XOR U9476 ( .A(n8865), .B(n4073), .Z(n4085) );
  XNOR U9477 ( .A(q[6]), .B(DB[692]), .Z(n4073) );
  IV U9478 ( .A(n4072), .Z(n8865) );
  XNOR U9479 ( .A(n4070), .B(n8866), .Z(n4072) );
  XNOR U9480 ( .A(q[5]), .B(DB[691]), .Z(n8866) );
  XNOR U9481 ( .A(q[4]), .B(DB[690]), .Z(n4070) );
  IV U9482 ( .A(n4084), .Z(n8864) );
  XOR U9483 ( .A(n8867), .B(n8868), .Z(n4084) );
  XNOR U9484 ( .A(n4080), .B(n4082), .Z(n8868) );
  XNOR U9485 ( .A(q[0]), .B(DB[686]), .Z(n4082) );
  XNOR U9486 ( .A(q[3]), .B(DB[689]), .Z(n4080) );
  IV U9487 ( .A(n4079), .Z(n8867) );
  XNOR U9488 ( .A(n4077), .B(n8869), .Z(n4079) );
  XNOR U9489 ( .A(q[2]), .B(DB[688]), .Z(n8869) );
  XNOR U9490 ( .A(q[1]), .B(DB[687]), .Z(n4077) );
  XOR U9491 ( .A(n8870), .B(n4042), .Z(n4005) );
  XOR U9492 ( .A(n8871), .B(n4030), .Z(n4042) );
  XNOR U9493 ( .A(q[6]), .B(DB[699]), .Z(n4030) );
  IV U9494 ( .A(n4029), .Z(n8871) );
  XNOR U9495 ( .A(n4027), .B(n8872), .Z(n4029) );
  XNOR U9496 ( .A(q[5]), .B(DB[698]), .Z(n8872) );
  XNOR U9497 ( .A(q[4]), .B(DB[697]), .Z(n4027) );
  IV U9498 ( .A(n4041), .Z(n8870) );
  XOR U9499 ( .A(n8873), .B(n8874), .Z(n4041) );
  XNOR U9500 ( .A(n4037), .B(n4039), .Z(n8874) );
  XNOR U9501 ( .A(q[0]), .B(DB[693]), .Z(n4039) );
  XNOR U9502 ( .A(q[3]), .B(DB[696]), .Z(n4037) );
  IV U9503 ( .A(n4036), .Z(n8873) );
  XNOR U9504 ( .A(n4034), .B(n8875), .Z(n4036) );
  XNOR U9505 ( .A(q[2]), .B(DB[695]), .Z(n8875) );
  XNOR U9506 ( .A(q[1]), .B(DB[694]), .Z(n4034) );
  XOR U9507 ( .A(n8876), .B(n3999), .Z(n3962) );
  XOR U9508 ( .A(n8877), .B(n3987), .Z(n3999) );
  XNOR U9509 ( .A(q[6]), .B(DB[706]), .Z(n3987) );
  IV U9510 ( .A(n3986), .Z(n8877) );
  XNOR U9511 ( .A(n3984), .B(n8878), .Z(n3986) );
  XNOR U9512 ( .A(q[5]), .B(DB[705]), .Z(n8878) );
  XNOR U9513 ( .A(q[4]), .B(DB[704]), .Z(n3984) );
  IV U9514 ( .A(n3998), .Z(n8876) );
  XOR U9515 ( .A(n8879), .B(n8880), .Z(n3998) );
  XNOR U9516 ( .A(n3994), .B(n3996), .Z(n8880) );
  XNOR U9517 ( .A(q[0]), .B(DB[700]), .Z(n3996) );
  XNOR U9518 ( .A(q[3]), .B(DB[703]), .Z(n3994) );
  IV U9519 ( .A(n3993), .Z(n8879) );
  XNOR U9520 ( .A(n3991), .B(n8881), .Z(n3993) );
  XNOR U9521 ( .A(q[2]), .B(DB[702]), .Z(n8881) );
  XNOR U9522 ( .A(q[1]), .B(DB[701]), .Z(n3991) );
  XOR U9523 ( .A(n8882), .B(n3956), .Z(n3919) );
  XOR U9524 ( .A(n8883), .B(n3944), .Z(n3956) );
  XNOR U9525 ( .A(q[6]), .B(DB[713]), .Z(n3944) );
  IV U9526 ( .A(n3943), .Z(n8883) );
  XNOR U9527 ( .A(n3941), .B(n8884), .Z(n3943) );
  XNOR U9528 ( .A(q[5]), .B(DB[712]), .Z(n8884) );
  XNOR U9529 ( .A(q[4]), .B(DB[711]), .Z(n3941) );
  IV U9530 ( .A(n3955), .Z(n8882) );
  XOR U9531 ( .A(n8885), .B(n8886), .Z(n3955) );
  XNOR U9532 ( .A(n3951), .B(n3953), .Z(n8886) );
  XNOR U9533 ( .A(q[0]), .B(DB[707]), .Z(n3953) );
  XNOR U9534 ( .A(q[3]), .B(DB[710]), .Z(n3951) );
  IV U9535 ( .A(n3950), .Z(n8885) );
  XNOR U9536 ( .A(n3948), .B(n8887), .Z(n3950) );
  XNOR U9537 ( .A(q[2]), .B(DB[709]), .Z(n8887) );
  XNOR U9538 ( .A(q[1]), .B(DB[708]), .Z(n3948) );
  XOR U9539 ( .A(n8888), .B(n3913), .Z(n3876) );
  XOR U9540 ( .A(n8889), .B(n3901), .Z(n3913) );
  XNOR U9541 ( .A(q[6]), .B(DB[720]), .Z(n3901) );
  IV U9542 ( .A(n3900), .Z(n8889) );
  XNOR U9543 ( .A(n3898), .B(n8890), .Z(n3900) );
  XNOR U9544 ( .A(q[5]), .B(DB[719]), .Z(n8890) );
  XNOR U9545 ( .A(q[4]), .B(DB[718]), .Z(n3898) );
  IV U9546 ( .A(n3912), .Z(n8888) );
  XOR U9547 ( .A(n8891), .B(n8892), .Z(n3912) );
  XNOR U9548 ( .A(n3908), .B(n3910), .Z(n8892) );
  XNOR U9549 ( .A(q[0]), .B(DB[714]), .Z(n3910) );
  XNOR U9550 ( .A(q[3]), .B(DB[717]), .Z(n3908) );
  IV U9551 ( .A(n3907), .Z(n8891) );
  XNOR U9552 ( .A(n3905), .B(n8893), .Z(n3907) );
  XNOR U9553 ( .A(q[2]), .B(DB[716]), .Z(n8893) );
  XNOR U9554 ( .A(q[1]), .B(DB[715]), .Z(n3905) );
  XOR U9555 ( .A(n8894), .B(n3870), .Z(n3833) );
  XOR U9556 ( .A(n8895), .B(n3858), .Z(n3870) );
  XNOR U9557 ( .A(q[6]), .B(DB[727]), .Z(n3858) );
  IV U9558 ( .A(n3857), .Z(n8895) );
  XNOR U9559 ( .A(n3855), .B(n8896), .Z(n3857) );
  XNOR U9560 ( .A(q[5]), .B(DB[726]), .Z(n8896) );
  XNOR U9561 ( .A(q[4]), .B(DB[725]), .Z(n3855) );
  IV U9562 ( .A(n3869), .Z(n8894) );
  XOR U9563 ( .A(n8897), .B(n8898), .Z(n3869) );
  XNOR U9564 ( .A(n3865), .B(n3867), .Z(n8898) );
  XNOR U9565 ( .A(q[0]), .B(DB[721]), .Z(n3867) );
  XNOR U9566 ( .A(q[3]), .B(DB[724]), .Z(n3865) );
  IV U9567 ( .A(n3864), .Z(n8897) );
  XNOR U9568 ( .A(n3862), .B(n8899), .Z(n3864) );
  XNOR U9569 ( .A(q[2]), .B(DB[723]), .Z(n8899) );
  XNOR U9570 ( .A(q[1]), .B(DB[722]), .Z(n3862) );
  XOR U9571 ( .A(n8900), .B(n3827), .Z(n3790) );
  XOR U9572 ( .A(n8901), .B(n3815), .Z(n3827) );
  XNOR U9573 ( .A(q[6]), .B(DB[734]), .Z(n3815) );
  IV U9574 ( .A(n3814), .Z(n8901) );
  XNOR U9575 ( .A(n3812), .B(n8902), .Z(n3814) );
  XNOR U9576 ( .A(q[5]), .B(DB[733]), .Z(n8902) );
  XNOR U9577 ( .A(q[4]), .B(DB[732]), .Z(n3812) );
  IV U9578 ( .A(n3826), .Z(n8900) );
  XOR U9579 ( .A(n8903), .B(n8904), .Z(n3826) );
  XNOR U9580 ( .A(n3822), .B(n3824), .Z(n8904) );
  XNOR U9581 ( .A(q[0]), .B(DB[728]), .Z(n3824) );
  XNOR U9582 ( .A(q[3]), .B(DB[731]), .Z(n3822) );
  IV U9583 ( .A(n3821), .Z(n8903) );
  XNOR U9584 ( .A(n3819), .B(n8905), .Z(n3821) );
  XNOR U9585 ( .A(q[2]), .B(DB[730]), .Z(n8905) );
  XNOR U9586 ( .A(q[1]), .B(DB[729]), .Z(n3819) );
  XOR U9587 ( .A(n8906), .B(n3784), .Z(n3747) );
  XOR U9588 ( .A(n8907), .B(n3772), .Z(n3784) );
  XNOR U9589 ( .A(q[6]), .B(DB[741]), .Z(n3772) );
  IV U9590 ( .A(n3771), .Z(n8907) );
  XNOR U9591 ( .A(n3769), .B(n8908), .Z(n3771) );
  XNOR U9592 ( .A(q[5]), .B(DB[740]), .Z(n8908) );
  XNOR U9593 ( .A(q[4]), .B(DB[739]), .Z(n3769) );
  IV U9594 ( .A(n3783), .Z(n8906) );
  XOR U9595 ( .A(n8909), .B(n8910), .Z(n3783) );
  XNOR U9596 ( .A(n3779), .B(n3781), .Z(n8910) );
  XNOR U9597 ( .A(q[0]), .B(DB[735]), .Z(n3781) );
  XNOR U9598 ( .A(q[3]), .B(DB[738]), .Z(n3779) );
  IV U9599 ( .A(n3778), .Z(n8909) );
  XNOR U9600 ( .A(n3776), .B(n8911), .Z(n3778) );
  XNOR U9601 ( .A(q[2]), .B(DB[737]), .Z(n8911) );
  XNOR U9602 ( .A(q[1]), .B(DB[736]), .Z(n3776) );
  XOR U9603 ( .A(n8912), .B(n3741), .Z(n3704) );
  XOR U9604 ( .A(n8913), .B(n3729), .Z(n3741) );
  XNOR U9605 ( .A(q[6]), .B(DB[748]), .Z(n3729) );
  IV U9606 ( .A(n3728), .Z(n8913) );
  XNOR U9607 ( .A(n3726), .B(n8914), .Z(n3728) );
  XNOR U9608 ( .A(q[5]), .B(DB[747]), .Z(n8914) );
  XNOR U9609 ( .A(q[4]), .B(DB[746]), .Z(n3726) );
  IV U9610 ( .A(n3740), .Z(n8912) );
  XOR U9611 ( .A(n8915), .B(n8916), .Z(n3740) );
  XNOR U9612 ( .A(n3736), .B(n3738), .Z(n8916) );
  XNOR U9613 ( .A(q[0]), .B(DB[742]), .Z(n3738) );
  XNOR U9614 ( .A(q[3]), .B(DB[745]), .Z(n3736) );
  IV U9615 ( .A(n3735), .Z(n8915) );
  XNOR U9616 ( .A(n3733), .B(n8917), .Z(n3735) );
  XNOR U9617 ( .A(q[2]), .B(DB[744]), .Z(n8917) );
  XNOR U9618 ( .A(q[1]), .B(DB[743]), .Z(n3733) );
  XOR U9619 ( .A(n8918), .B(n3698), .Z(n3661) );
  XOR U9620 ( .A(n8919), .B(n3686), .Z(n3698) );
  XNOR U9621 ( .A(q[6]), .B(DB[755]), .Z(n3686) );
  IV U9622 ( .A(n3685), .Z(n8919) );
  XNOR U9623 ( .A(n3683), .B(n8920), .Z(n3685) );
  XNOR U9624 ( .A(q[5]), .B(DB[754]), .Z(n8920) );
  XNOR U9625 ( .A(q[4]), .B(DB[753]), .Z(n3683) );
  IV U9626 ( .A(n3697), .Z(n8918) );
  XOR U9627 ( .A(n8921), .B(n8922), .Z(n3697) );
  XNOR U9628 ( .A(n3693), .B(n3695), .Z(n8922) );
  XNOR U9629 ( .A(q[0]), .B(DB[749]), .Z(n3695) );
  XNOR U9630 ( .A(q[3]), .B(DB[752]), .Z(n3693) );
  IV U9631 ( .A(n3692), .Z(n8921) );
  XNOR U9632 ( .A(n3690), .B(n8923), .Z(n3692) );
  XNOR U9633 ( .A(q[2]), .B(DB[751]), .Z(n8923) );
  XNOR U9634 ( .A(q[1]), .B(DB[750]), .Z(n3690) );
  XOR U9635 ( .A(n8924), .B(n3655), .Z(n3618) );
  XOR U9636 ( .A(n8925), .B(n3643), .Z(n3655) );
  XNOR U9637 ( .A(q[6]), .B(DB[762]), .Z(n3643) );
  IV U9638 ( .A(n3642), .Z(n8925) );
  XNOR U9639 ( .A(n3640), .B(n8926), .Z(n3642) );
  XNOR U9640 ( .A(q[5]), .B(DB[761]), .Z(n8926) );
  XNOR U9641 ( .A(q[4]), .B(DB[760]), .Z(n3640) );
  IV U9642 ( .A(n3654), .Z(n8924) );
  XOR U9643 ( .A(n8927), .B(n8928), .Z(n3654) );
  XNOR U9644 ( .A(n3650), .B(n3652), .Z(n8928) );
  XNOR U9645 ( .A(q[0]), .B(DB[756]), .Z(n3652) );
  XNOR U9646 ( .A(q[3]), .B(DB[759]), .Z(n3650) );
  IV U9647 ( .A(n3649), .Z(n8927) );
  XNOR U9648 ( .A(n3647), .B(n8929), .Z(n3649) );
  XNOR U9649 ( .A(q[2]), .B(DB[758]), .Z(n8929) );
  XNOR U9650 ( .A(q[1]), .B(DB[757]), .Z(n3647) );
  XOR U9651 ( .A(n8930), .B(n3612), .Z(n3575) );
  XOR U9652 ( .A(n8931), .B(n3600), .Z(n3612) );
  XNOR U9653 ( .A(q[6]), .B(DB[769]), .Z(n3600) );
  IV U9654 ( .A(n3599), .Z(n8931) );
  XNOR U9655 ( .A(n3597), .B(n8932), .Z(n3599) );
  XNOR U9656 ( .A(q[5]), .B(DB[768]), .Z(n8932) );
  XNOR U9657 ( .A(q[4]), .B(DB[767]), .Z(n3597) );
  IV U9658 ( .A(n3611), .Z(n8930) );
  XOR U9659 ( .A(n8933), .B(n8934), .Z(n3611) );
  XNOR U9660 ( .A(n3607), .B(n3609), .Z(n8934) );
  XNOR U9661 ( .A(q[0]), .B(DB[763]), .Z(n3609) );
  XNOR U9662 ( .A(q[3]), .B(DB[766]), .Z(n3607) );
  IV U9663 ( .A(n3606), .Z(n8933) );
  XNOR U9664 ( .A(n3604), .B(n8935), .Z(n3606) );
  XNOR U9665 ( .A(q[2]), .B(DB[765]), .Z(n8935) );
  XNOR U9666 ( .A(q[1]), .B(DB[764]), .Z(n3604) );
  XOR U9667 ( .A(n8936), .B(n3569), .Z(n3532) );
  XOR U9668 ( .A(n8937), .B(n3557), .Z(n3569) );
  XNOR U9669 ( .A(q[6]), .B(DB[776]), .Z(n3557) );
  IV U9670 ( .A(n3556), .Z(n8937) );
  XNOR U9671 ( .A(n3554), .B(n8938), .Z(n3556) );
  XNOR U9672 ( .A(q[5]), .B(DB[775]), .Z(n8938) );
  XNOR U9673 ( .A(q[4]), .B(DB[774]), .Z(n3554) );
  IV U9674 ( .A(n3568), .Z(n8936) );
  XOR U9675 ( .A(n8939), .B(n8940), .Z(n3568) );
  XNOR U9676 ( .A(n3564), .B(n3566), .Z(n8940) );
  XNOR U9677 ( .A(q[0]), .B(DB[770]), .Z(n3566) );
  XNOR U9678 ( .A(q[3]), .B(DB[773]), .Z(n3564) );
  IV U9679 ( .A(n3563), .Z(n8939) );
  XNOR U9680 ( .A(n3561), .B(n8941), .Z(n3563) );
  XNOR U9681 ( .A(q[2]), .B(DB[772]), .Z(n8941) );
  XNOR U9682 ( .A(q[1]), .B(DB[771]), .Z(n3561) );
  XOR U9683 ( .A(n8942), .B(n3526), .Z(n3489) );
  XOR U9684 ( .A(n8943), .B(n3514), .Z(n3526) );
  XNOR U9685 ( .A(q[6]), .B(DB[783]), .Z(n3514) );
  IV U9686 ( .A(n3513), .Z(n8943) );
  XNOR U9687 ( .A(n3511), .B(n8944), .Z(n3513) );
  XNOR U9688 ( .A(q[5]), .B(DB[782]), .Z(n8944) );
  XNOR U9689 ( .A(q[4]), .B(DB[781]), .Z(n3511) );
  IV U9690 ( .A(n3525), .Z(n8942) );
  XOR U9691 ( .A(n8945), .B(n8946), .Z(n3525) );
  XNOR U9692 ( .A(n3521), .B(n3523), .Z(n8946) );
  XNOR U9693 ( .A(q[0]), .B(DB[777]), .Z(n3523) );
  XNOR U9694 ( .A(q[3]), .B(DB[780]), .Z(n3521) );
  IV U9695 ( .A(n3520), .Z(n8945) );
  XNOR U9696 ( .A(n3518), .B(n8947), .Z(n3520) );
  XNOR U9697 ( .A(q[2]), .B(DB[779]), .Z(n8947) );
  XNOR U9698 ( .A(q[1]), .B(DB[778]), .Z(n3518) );
  XOR U9699 ( .A(n8948), .B(n3483), .Z(n3446) );
  XOR U9700 ( .A(n8949), .B(n3471), .Z(n3483) );
  XNOR U9701 ( .A(q[6]), .B(DB[790]), .Z(n3471) );
  IV U9702 ( .A(n3470), .Z(n8949) );
  XNOR U9703 ( .A(n3468), .B(n8950), .Z(n3470) );
  XNOR U9704 ( .A(q[5]), .B(DB[789]), .Z(n8950) );
  XNOR U9705 ( .A(q[4]), .B(DB[788]), .Z(n3468) );
  IV U9706 ( .A(n3482), .Z(n8948) );
  XOR U9707 ( .A(n8951), .B(n8952), .Z(n3482) );
  XNOR U9708 ( .A(n3478), .B(n3480), .Z(n8952) );
  XNOR U9709 ( .A(q[0]), .B(DB[784]), .Z(n3480) );
  XNOR U9710 ( .A(q[3]), .B(DB[787]), .Z(n3478) );
  IV U9711 ( .A(n3477), .Z(n8951) );
  XNOR U9712 ( .A(n3475), .B(n8953), .Z(n3477) );
  XNOR U9713 ( .A(q[2]), .B(DB[786]), .Z(n8953) );
  XNOR U9714 ( .A(q[1]), .B(DB[785]), .Z(n3475) );
  XOR U9715 ( .A(n8954), .B(n3440), .Z(n3403) );
  XOR U9716 ( .A(n8955), .B(n3428), .Z(n3440) );
  XNOR U9717 ( .A(q[6]), .B(DB[797]), .Z(n3428) );
  IV U9718 ( .A(n3427), .Z(n8955) );
  XNOR U9719 ( .A(n3425), .B(n8956), .Z(n3427) );
  XNOR U9720 ( .A(q[5]), .B(DB[796]), .Z(n8956) );
  XNOR U9721 ( .A(q[4]), .B(DB[795]), .Z(n3425) );
  IV U9722 ( .A(n3439), .Z(n8954) );
  XOR U9723 ( .A(n8957), .B(n8958), .Z(n3439) );
  XNOR U9724 ( .A(n3435), .B(n3437), .Z(n8958) );
  XNOR U9725 ( .A(q[0]), .B(DB[791]), .Z(n3437) );
  XNOR U9726 ( .A(q[3]), .B(DB[794]), .Z(n3435) );
  IV U9727 ( .A(n3434), .Z(n8957) );
  XNOR U9728 ( .A(n3432), .B(n8959), .Z(n3434) );
  XNOR U9729 ( .A(q[2]), .B(DB[793]), .Z(n8959) );
  XNOR U9730 ( .A(q[1]), .B(DB[792]), .Z(n3432) );
  XOR U9731 ( .A(n8960), .B(n3397), .Z(n3360) );
  XOR U9732 ( .A(n8961), .B(n3385), .Z(n3397) );
  XNOR U9733 ( .A(q[6]), .B(DB[804]), .Z(n3385) );
  IV U9734 ( .A(n3384), .Z(n8961) );
  XNOR U9735 ( .A(n3382), .B(n8962), .Z(n3384) );
  XNOR U9736 ( .A(q[5]), .B(DB[803]), .Z(n8962) );
  XNOR U9737 ( .A(q[4]), .B(DB[802]), .Z(n3382) );
  IV U9738 ( .A(n3396), .Z(n8960) );
  XOR U9739 ( .A(n8963), .B(n8964), .Z(n3396) );
  XNOR U9740 ( .A(n3392), .B(n3394), .Z(n8964) );
  XNOR U9741 ( .A(q[0]), .B(DB[798]), .Z(n3394) );
  XNOR U9742 ( .A(q[3]), .B(DB[801]), .Z(n3392) );
  IV U9743 ( .A(n3391), .Z(n8963) );
  XNOR U9744 ( .A(n3389), .B(n8965), .Z(n3391) );
  XNOR U9745 ( .A(q[2]), .B(DB[800]), .Z(n8965) );
  XNOR U9746 ( .A(q[1]), .B(DB[799]), .Z(n3389) );
  XOR U9747 ( .A(n8966), .B(n3354), .Z(n3317) );
  XOR U9748 ( .A(n8967), .B(n3342), .Z(n3354) );
  XNOR U9749 ( .A(q[6]), .B(DB[811]), .Z(n3342) );
  IV U9750 ( .A(n3341), .Z(n8967) );
  XNOR U9751 ( .A(n3339), .B(n8968), .Z(n3341) );
  XNOR U9752 ( .A(q[5]), .B(DB[810]), .Z(n8968) );
  XNOR U9753 ( .A(q[4]), .B(DB[809]), .Z(n3339) );
  IV U9754 ( .A(n3353), .Z(n8966) );
  XOR U9755 ( .A(n8969), .B(n8970), .Z(n3353) );
  XNOR U9756 ( .A(n3349), .B(n3351), .Z(n8970) );
  XNOR U9757 ( .A(q[0]), .B(DB[805]), .Z(n3351) );
  XNOR U9758 ( .A(q[3]), .B(DB[808]), .Z(n3349) );
  IV U9759 ( .A(n3348), .Z(n8969) );
  XNOR U9760 ( .A(n3346), .B(n8971), .Z(n3348) );
  XNOR U9761 ( .A(q[2]), .B(DB[807]), .Z(n8971) );
  XNOR U9762 ( .A(q[1]), .B(DB[806]), .Z(n3346) );
  XOR U9763 ( .A(n8972), .B(n3311), .Z(n3274) );
  XOR U9764 ( .A(n8973), .B(n3299), .Z(n3311) );
  XNOR U9765 ( .A(q[6]), .B(DB[818]), .Z(n3299) );
  IV U9766 ( .A(n3298), .Z(n8973) );
  XNOR U9767 ( .A(n3296), .B(n8974), .Z(n3298) );
  XNOR U9768 ( .A(q[5]), .B(DB[817]), .Z(n8974) );
  XNOR U9769 ( .A(q[4]), .B(DB[816]), .Z(n3296) );
  IV U9770 ( .A(n3310), .Z(n8972) );
  XOR U9771 ( .A(n8975), .B(n8976), .Z(n3310) );
  XNOR U9772 ( .A(n3306), .B(n3308), .Z(n8976) );
  XNOR U9773 ( .A(q[0]), .B(DB[812]), .Z(n3308) );
  XNOR U9774 ( .A(q[3]), .B(DB[815]), .Z(n3306) );
  IV U9775 ( .A(n3305), .Z(n8975) );
  XNOR U9776 ( .A(n3303), .B(n8977), .Z(n3305) );
  XNOR U9777 ( .A(q[2]), .B(DB[814]), .Z(n8977) );
  XNOR U9778 ( .A(q[1]), .B(DB[813]), .Z(n3303) );
  XOR U9779 ( .A(n8978), .B(n3268), .Z(n3231) );
  XOR U9780 ( .A(n8979), .B(n3256), .Z(n3268) );
  XNOR U9781 ( .A(q[6]), .B(DB[825]), .Z(n3256) );
  IV U9782 ( .A(n3255), .Z(n8979) );
  XNOR U9783 ( .A(n3253), .B(n8980), .Z(n3255) );
  XNOR U9784 ( .A(q[5]), .B(DB[824]), .Z(n8980) );
  XNOR U9785 ( .A(q[4]), .B(DB[823]), .Z(n3253) );
  IV U9786 ( .A(n3267), .Z(n8978) );
  XOR U9787 ( .A(n8981), .B(n8982), .Z(n3267) );
  XNOR U9788 ( .A(n3263), .B(n3265), .Z(n8982) );
  XNOR U9789 ( .A(q[0]), .B(DB[819]), .Z(n3265) );
  XNOR U9790 ( .A(q[3]), .B(DB[822]), .Z(n3263) );
  IV U9791 ( .A(n3262), .Z(n8981) );
  XNOR U9792 ( .A(n3260), .B(n8983), .Z(n3262) );
  XNOR U9793 ( .A(q[2]), .B(DB[821]), .Z(n8983) );
  XNOR U9794 ( .A(q[1]), .B(DB[820]), .Z(n3260) );
  XOR U9795 ( .A(n8984), .B(n3225), .Z(n3188) );
  XOR U9796 ( .A(n8985), .B(n3213), .Z(n3225) );
  XNOR U9797 ( .A(q[6]), .B(DB[832]), .Z(n3213) );
  IV U9798 ( .A(n3212), .Z(n8985) );
  XNOR U9799 ( .A(n3210), .B(n8986), .Z(n3212) );
  XNOR U9800 ( .A(q[5]), .B(DB[831]), .Z(n8986) );
  XNOR U9801 ( .A(q[4]), .B(DB[830]), .Z(n3210) );
  IV U9802 ( .A(n3224), .Z(n8984) );
  XOR U9803 ( .A(n8987), .B(n8988), .Z(n3224) );
  XNOR U9804 ( .A(n3220), .B(n3222), .Z(n8988) );
  XNOR U9805 ( .A(q[0]), .B(DB[826]), .Z(n3222) );
  XNOR U9806 ( .A(q[3]), .B(DB[829]), .Z(n3220) );
  IV U9807 ( .A(n3219), .Z(n8987) );
  XNOR U9808 ( .A(n3217), .B(n8989), .Z(n3219) );
  XNOR U9809 ( .A(q[2]), .B(DB[828]), .Z(n8989) );
  XNOR U9810 ( .A(q[1]), .B(DB[827]), .Z(n3217) );
  XOR U9811 ( .A(n8990), .B(n3182), .Z(n3145) );
  XOR U9812 ( .A(n8991), .B(n3170), .Z(n3182) );
  XNOR U9813 ( .A(q[6]), .B(DB[839]), .Z(n3170) );
  IV U9814 ( .A(n3169), .Z(n8991) );
  XNOR U9815 ( .A(n3167), .B(n8992), .Z(n3169) );
  XNOR U9816 ( .A(q[5]), .B(DB[838]), .Z(n8992) );
  XNOR U9817 ( .A(q[4]), .B(DB[837]), .Z(n3167) );
  IV U9818 ( .A(n3181), .Z(n8990) );
  XOR U9819 ( .A(n8993), .B(n8994), .Z(n3181) );
  XNOR U9820 ( .A(n3177), .B(n3179), .Z(n8994) );
  XNOR U9821 ( .A(q[0]), .B(DB[833]), .Z(n3179) );
  XNOR U9822 ( .A(q[3]), .B(DB[836]), .Z(n3177) );
  IV U9823 ( .A(n3176), .Z(n8993) );
  XNOR U9824 ( .A(n3174), .B(n8995), .Z(n3176) );
  XNOR U9825 ( .A(q[2]), .B(DB[835]), .Z(n8995) );
  XNOR U9826 ( .A(q[1]), .B(DB[834]), .Z(n3174) );
  XOR U9827 ( .A(n8996), .B(n3139), .Z(n3102) );
  XOR U9828 ( .A(n8997), .B(n3127), .Z(n3139) );
  XNOR U9829 ( .A(q[6]), .B(DB[846]), .Z(n3127) );
  IV U9830 ( .A(n3126), .Z(n8997) );
  XNOR U9831 ( .A(n3124), .B(n8998), .Z(n3126) );
  XNOR U9832 ( .A(q[5]), .B(DB[845]), .Z(n8998) );
  XNOR U9833 ( .A(q[4]), .B(DB[844]), .Z(n3124) );
  IV U9834 ( .A(n3138), .Z(n8996) );
  XOR U9835 ( .A(n8999), .B(n9000), .Z(n3138) );
  XNOR U9836 ( .A(n3134), .B(n3136), .Z(n9000) );
  XNOR U9837 ( .A(q[0]), .B(DB[840]), .Z(n3136) );
  XNOR U9838 ( .A(q[3]), .B(DB[843]), .Z(n3134) );
  IV U9839 ( .A(n3133), .Z(n8999) );
  XNOR U9840 ( .A(n3131), .B(n9001), .Z(n3133) );
  XNOR U9841 ( .A(q[2]), .B(DB[842]), .Z(n9001) );
  XNOR U9842 ( .A(q[1]), .B(DB[841]), .Z(n3131) );
  XOR U9843 ( .A(n9002), .B(n3096), .Z(n3059) );
  XOR U9844 ( .A(n9003), .B(n3084), .Z(n3096) );
  XNOR U9845 ( .A(q[6]), .B(DB[853]), .Z(n3084) );
  IV U9846 ( .A(n3083), .Z(n9003) );
  XNOR U9847 ( .A(n3081), .B(n9004), .Z(n3083) );
  XNOR U9848 ( .A(q[5]), .B(DB[852]), .Z(n9004) );
  XNOR U9849 ( .A(q[4]), .B(DB[851]), .Z(n3081) );
  IV U9850 ( .A(n3095), .Z(n9002) );
  XOR U9851 ( .A(n9005), .B(n9006), .Z(n3095) );
  XNOR U9852 ( .A(n3091), .B(n3093), .Z(n9006) );
  XNOR U9853 ( .A(q[0]), .B(DB[847]), .Z(n3093) );
  XNOR U9854 ( .A(q[3]), .B(DB[850]), .Z(n3091) );
  IV U9855 ( .A(n3090), .Z(n9005) );
  XNOR U9856 ( .A(n3088), .B(n9007), .Z(n3090) );
  XNOR U9857 ( .A(q[2]), .B(DB[849]), .Z(n9007) );
  XNOR U9858 ( .A(q[1]), .B(DB[848]), .Z(n3088) );
  XOR U9859 ( .A(n9008), .B(n3053), .Z(n3016) );
  XOR U9860 ( .A(n9009), .B(n3041), .Z(n3053) );
  XNOR U9861 ( .A(q[6]), .B(DB[860]), .Z(n3041) );
  IV U9862 ( .A(n3040), .Z(n9009) );
  XNOR U9863 ( .A(n3038), .B(n9010), .Z(n3040) );
  XNOR U9864 ( .A(q[5]), .B(DB[859]), .Z(n9010) );
  XNOR U9865 ( .A(q[4]), .B(DB[858]), .Z(n3038) );
  IV U9866 ( .A(n3052), .Z(n9008) );
  XOR U9867 ( .A(n9011), .B(n9012), .Z(n3052) );
  XNOR U9868 ( .A(n3048), .B(n3050), .Z(n9012) );
  XNOR U9869 ( .A(q[0]), .B(DB[854]), .Z(n3050) );
  XNOR U9870 ( .A(q[3]), .B(DB[857]), .Z(n3048) );
  IV U9871 ( .A(n3047), .Z(n9011) );
  XNOR U9872 ( .A(n3045), .B(n9013), .Z(n3047) );
  XNOR U9873 ( .A(q[2]), .B(DB[856]), .Z(n9013) );
  XNOR U9874 ( .A(q[1]), .B(DB[855]), .Z(n3045) );
  XOR U9875 ( .A(n9014), .B(n3010), .Z(n2973) );
  XOR U9876 ( .A(n9015), .B(n2998), .Z(n3010) );
  XNOR U9877 ( .A(q[6]), .B(DB[867]), .Z(n2998) );
  IV U9878 ( .A(n2997), .Z(n9015) );
  XNOR U9879 ( .A(n2995), .B(n9016), .Z(n2997) );
  XNOR U9880 ( .A(q[5]), .B(DB[866]), .Z(n9016) );
  XNOR U9881 ( .A(q[4]), .B(DB[865]), .Z(n2995) );
  IV U9882 ( .A(n3009), .Z(n9014) );
  XOR U9883 ( .A(n9017), .B(n9018), .Z(n3009) );
  XNOR U9884 ( .A(n3005), .B(n3007), .Z(n9018) );
  XNOR U9885 ( .A(q[0]), .B(DB[861]), .Z(n3007) );
  XNOR U9886 ( .A(q[3]), .B(DB[864]), .Z(n3005) );
  IV U9887 ( .A(n3004), .Z(n9017) );
  XNOR U9888 ( .A(n3002), .B(n9019), .Z(n3004) );
  XNOR U9889 ( .A(q[2]), .B(DB[863]), .Z(n9019) );
  XNOR U9890 ( .A(q[1]), .B(DB[862]), .Z(n3002) );
  XOR U9891 ( .A(n9020), .B(n2967), .Z(n2930) );
  XOR U9892 ( .A(n9021), .B(n2955), .Z(n2967) );
  XNOR U9893 ( .A(q[6]), .B(DB[874]), .Z(n2955) );
  IV U9894 ( .A(n2954), .Z(n9021) );
  XNOR U9895 ( .A(n2952), .B(n9022), .Z(n2954) );
  XNOR U9896 ( .A(q[5]), .B(DB[873]), .Z(n9022) );
  XNOR U9897 ( .A(q[4]), .B(DB[872]), .Z(n2952) );
  IV U9898 ( .A(n2966), .Z(n9020) );
  XOR U9899 ( .A(n9023), .B(n9024), .Z(n2966) );
  XNOR U9900 ( .A(n2962), .B(n2964), .Z(n9024) );
  XNOR U9901 ( .A(q[0]), .B(DB[868]), .Z(n2964) );
  XNOR U9902 ( .A(q[3]), .B(DB[871]), .Z(n2962) );
  IV U9903 ( .A(n2961), .Z(n9023) );
  XNOR U9904 ( .A(n2959), .B(n9025), .Z(n2961) );
  XNOR U9905 ( .A(q[2]), .B(DB[870]), .Z(n9025) );
  XNOR U9906 ( .A(q[1]), .B(DB[869]), .Z(n2959) );
  XOR U9907 ( .A(n9026), .B(n2924), .Z(n2887) );
  XOR U9908 ( .A(n9027), .B(n2912), .Z(n2924) );
  XNOR U9909 ( .A(q[6]), .B(DB[881]), .Z(n2912) );
  IV U9910 ( .A(n2911), .Z(n9027) );
  XNOR U9911 ( .A(n2909), .B(n9028), .Z(n2911) );
  XNOR U9912 ( .A(q[5]), .B(DB[880]), .Z(n9028) );
  XNOR U9913 ( .A(q[4]), .B(DB[879]), .Z(n2909) );
  IV U9914 ( .A(n2923), .Z(n9026) );
  XOR U9915 ( .A(n9029), .B(n9030), .Z(n2923) );
  XNOR U9916 ( .A(n2919), .B(n2921), .Z(n9030) );
  XNOR U9917 ( .A(q[0]), .B(DB[875]), .Z(n2921) );
  XNOR U9918 ( .A(q[3]), .B(DB[878]), .Z(n2919) );
  IV U9919 ( .A(n2918), .Z(n9029) );
  XNOR U9920 ( .A(n2916), .B(n9031), .Z(n2918) );
  XNOR U9921 ( .A(q[2]), .B(DB[877]), .Z(n9031) );
  XNOR U9922 ( .A(q[1]), .B(DB[876]), .Z(n2916) );
  XOR U9923 ( .A(n9032), .B(n2881), .Z(n2843) );
  XOR U9924 ( .A(n9033), .B(n2869), .Z(n2881) );
  XNOR U9925 ( .A(q[6]), .B(DB[888]), .Z(n2869) );
  IV U9926 ( .A(n2868), .Z(n9033) );
  XNOR U9927 ( .A(n2866), .B(n9034), .Z(n2868) );
  XNOR U9928 ( .A(q[5]), .B(DB[887]), .Z(n9034) );
  XOR U9929 ( .A(q[4]), .B(n893), .Z(n2866) );
  IV U9930 ( .A(DB[886]), .Z(n893) );
  IV U9931 ( .A(n2880), .Z(n9032) );
  XOR U9932 ( .A(n9035), .B(n9036), .Z(n2880) );
  XNOR U9933 ( .A(n2876), .B(n2878), .Z(n9036) );
  XNOR U9934 ( .A(q[0]), .B(DB[882]), .Z(n2878) );
  XOR U9935 ( .A(q[3]), .B(n1275), .Z(n2876) );
  IV U9936 ( .A(DB[885]), .Z(n1275) );
  IV U9937 ( .A(n2875), .Z(n9035) );
  XNOR U9938 ( .A(n2873), .B(n9037), .Z(n2875) );
  XNOR U9939 ( .A(q[2]), .B(DB[884]), .Z(n9037) );
  XNOR U9940 ( .A(q[1]), .B(DB[883]), .Z(n2873) );
endmodule

