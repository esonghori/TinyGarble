
module hamming_N16000_CC64 ( clk, rst, x, y, o );
  input [249:0] x;
  input [249:0] y;
  output [13:0] o;
  input clk, rst;
  wire   n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035;
  wire   [13:0] oglobal;

  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[0]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[1]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[2]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[3]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[4]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[5]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[6]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[7]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[8]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[9]) );
  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[10]) );
  DFF \oglobal_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[11]) );
  DFF \oglobal_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[12]) );
  DFF \oglobal_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        oglobal[13]) );
  XNOR U267 ( .A(n334), .B(n335), .Z(n347) );
  XNOR U268 ( .A(n315), .B(n566), .Z(n321) );
  XNOR U269 ( .A(n365), .B(n642), .Z(n371) );
  XNOR U270 ( .A(n383), .B(n384), .Z(n396) );
  XNOR U271 ( .A(n224), .B(n225), .Z(n233) );
  XNOR U272 ( .A(n297), .B(n509), .Z(n280) );
  XNOR U273 ( .A(n417), .B(n419), .Z(n438) );
  XNOR U274 ( .A(n154), .B(n251), .Z(n137) );
  XNOR U275 ( .A(n40), .B(n53), .Z(n42) );
  XNOR U276 ( .A(n187), .B(n299), .Z(n161) );
  XNOR U277 ( .A(n267), .B(n490), .Z(n273) );
  XNOR U278 ( .A(n116), .B(n118), .Z(n130) );
  XNOR U279 ( .A(n493), .B(n495), .Z(n514) );
  XNOR U280 ( .A(n645), .B(n647), .Z(n666) );
  XNOR U281 ( .A(n102), .B(n182), .Z(n108) );
  XNOR U282 ( .A(n232), .B(n233), .Z(n257) );
  XNOR U283 ( .A(n436), .B(n438), .Z(n476) );
  XNOR U284 ( .A(n588), .B(n590), .Z(n628) );
  XNOR U285 ( .A(n57), .B(n86), .Z(n63) );
  XNOR U286 ( .A(n354), .B(n547), .Z(n304) );
  XOR U287 ( .A(oglobal[7]), .B(n37), .Z(n15) );
  XOR U288 ( .A(oglobal[4]), .B(n111), .Z(n21) );
  ANDN U289 ( .B(n1015), .A(n686), .Z(n688) );
  XNOR U290 ( .A(n140), .B(n263), .Z(n142) );
  XNOR U291 ( .A(n359), .B(n360), .Z(n372) );
  XNOR U292 ( .A(n1003), .B(n1002), .Z(n1022) );
  XNOR U293 ( .A(n982), .B(n981), .Z(n979) );
  XNOR U294 ( .A(n940), .B(n939), .Z(n937) );
  XNOR U295 ( .A(n898), .B(n897), .Z(n895) );
  XNOR U296 ( .A(n858), .B(n857), .Z(n855) );
  XNOR U297 ( .A(n814), .B(n813), .Z(n811) );
  XNOR U298 ( .A(n774), .B(n773), .Z(n771) );
  XNOR U299 ( .A(n732), .B(n731), .Z(n729) );
  XNOR U300 ( .A(n148), .B(n275), .Z(n154) );
  XNOR U301 ( .A(n249), .B(n433), .Z(n232) );
  XNOR U302 ( .A(n395), .B(n661), .Z(n378) );
  XNOR U303 ( .A(n569), .B(n571), .Z(n590) );
  XNOR U304 ( .A(n71), .B(n73), .Z(n85) );
  XNOR U305 ( .A(n129), .B(n130), .Z(n138) );
  XNOR U306 ( .A(n280), .B(n471), .Z(n256) );
  XNOR U307 ( .A(n329), .B(n330), .Z(n355) );
  XNOR U308 ( .A(n664), .B(n951), .Z(n626) );
  XNOR U309 ( .A(n108), .B(n156), .Z(n91) );
  XNOR U310 ( .A(n474), .B(n476), .Z(n552) );
  XOR U311 ( .A(oglobal[6]), .B(n45), .Z(n17) );
  XOR U312 ( .A(oglobal[3]), .B(n207), .Z(n23) );
  ANDN U313 ( .B(n847), .A(n534), .Z(n536) );
  ANDN U314 ( .B(n929), .A(n610), .Z(n612) );
  XNOR U315 ( .A(n190), .B(n361), .Z(n192) );
  XNOR U316 ( .A(n243), .B(n452), .Z(n249) );
  XNOR U317 ( .A(n261), .B(n262), .Z(n274) );
  XNOR U318 ( .A(n285), .B(n286), .Z(n298) );
  XNOR U319 ( .A(n309), .B(n310), .Z(n322) );
  XNOR U320 ( .A(n1026), .B(n1025), .Z(n1023) );
  XNOR U321 ( .A(n961), .B(n960), .Z(n978) );
  XNOR U322 ( .A(n917), .B(n916), .Z(n936) );
  XNOR U323 ( .A(n877), .B(n876), .Z(n894) );
  XNOR U324 ( .A(n835), .B(n834), .Z(n854) );
  XNOR U325 ( .A(n793), .B(n792), .Z(n810) );
  XNOR U326 ( .A(n198), .B(n373), .Z(n204) );
  XNOR U327 ( .A(n346), .B(n585), .Z(n329) );
  XNOR U328 ( .A(n455), .B(n741), .Z(n436) );
  XNOR U329 ( .A(n96), .B(n97), .Z(n109) );
  XNOR U330 ( .A(n180), .B(n181), .Z(n188) );
  XNOR U331 ( .A(n378), .B(n623), .Z(n354) );
  XNOR U332 ( .A(n512), .B(n783), .Z(n474) );
  XNOR U333 ( .A(n50), .B(n52), .Z(n64) );
  XNOR U334 ( .A(n84), .B(n85), .Z(n92) );
  XNOR U335 ( .A(n137), .B(n138), .Z(n162) );
  XNOR U336 ( .A(n256), .B(n257), .Z(n305) );
  XNOR U337 ( .A(n626), .B(n867), .Z(n550) );
  XOR U338 ( .A(oglobal[5]), .B(n66), .Z(n19) );
  XOR U339 ( .A(oglobal[2]), .B(n398), .Z(n25) );
  ANDN U340 ( .B(n721), .A(n420), .Z(n422) );
  ANDN U341 ( .B(n763), .A(n458), .Z(n460) );
  ANDN U342 ( .B(n803), .A(n496), .Z(n498) );
  ANDN U343 ( .B(n887), .A(n572), .Z(n574) );
  ANDN U344 ( .B(n971), .A(n648), .Z(n650) );
  XNOR U345 ( .A(n212), .B(n213), .Z(n225) );
  XNOR U346 ( .A(n237), .B(n238), .Z(n250) );
  XNOR U347 ( .A(n291), .B(n528), .Z(n297) );
  XNOR U348 ( .A(n340), .B(n604), .Z(n346) );
  XNOR U349 ( .A(n389), .B(n680), .Z(n395) );
  XNOR U350 ( .A(n751), .B(n750), .Z(n770) );
  XNOR U351 ( .A(n711), .B(n710), .Z(n728) );
  XNOR U352 ( .A(n142), .B(n143), .Z(n155) );
  XNOR U353 ( .A(n166), .B(n168), .Z(n181) );
  XNOR U354 ( .A(n192), .B(n193), .Z(n205) );
  XNOR U355 ( .A(n273), .B(n274), .Z(n281) );
  XNOR U356 ( .A(n321), .B(n322), .Z(n330) );
  XNOR U357 ( .A(n371), .B(n372), .Z(n379) );
  XNOR U358 ( .A(n531), .B(n825), .Z(n512) );
  XNOR U359 ( .A(n607), .B(n907), .Z(n588) );
  XNOR U360 ( .A(n683), .B(n993), .Z(n664) );
  XNOR U361 ( .A(n42), .B(n43), .Z(n18) );
  XNOR U362 ( .A(n63), .B(n64), .Z(n20) );
  XNOR U363 ( .A(n91), .B(n92), .Z(n22) );
  XNOR U364 ( .A(n161), .B(n162), .Z(n24) );
  XNOR U365 ( .A(n304), .B(n305), .Z(n26) );
  XNOR U366 ( .A(n550), .B(n552), .Z(n28) );
  XNOR U367 ( .A(n15), .B(n16), .Z(o[7]) );
  XOR U368 ( .A(n17), .B(n18), .Z(o[6]) );
  XOR U369 ( .A(n19), .B(n20), .Z(o[5]) );
  XOR U370 ( .A(n21), .B(n22), .Z(o[4]) );
  XOR U371 ( .A(n23), .B(n24), .Z(o[3]) );
  XOR U372 ( .A(n25), .B(n26), .Z(o[2]) );
  XOR U373 ( .A(n27), .B(n28), .Z(o[1]) );
  XOR U374 ( .A(n29), .B(n30), .Z(o[13]) );
  XOR U375 ( .A(oglobal[13]), .B(n31), .Z(n30) );
  AND U376 ( .A(n29), .B(o[12]), .Z(n31) );
  XOR U377 ( .A(oglobal[12]), .B(n29), .Z(o[12]) );
  ANDN U378 ( .B(n32), .A(o[11]), .Z(n29) );
  XOR U379 ( .A(oglobal[11]), .B(n32), .Z(o[11]) );
  ANDN U380 ( .B(n33), .A(o[10]), .Z(n32) );
  XOR U381 ( .A(oglobal[10]), .B(n33), .Z(o[10]) );
  ANDN U382 ( .B(n34), .A(o[9]), .Z(n33) );
  XOR U383 ( .A(oglobal[9]), .B(n34), .Z(o[9]) );
  ANDN U384 ( .B(n35), .A(o[8]), .Z(n34) );
  XOR U385 ( .A(oglobal[8]), .B(n35), .Z(o[8]) );
  XNOR U386 ( .A(n36), .B(n37), .Z(n35) );
  ANDN U387 ( .B(n38), .A(n15), .Z(n36) );
  XNOR U388 ( .A(n37), .B(n16), .Z(n38) );
  XNOR U389 ( .A(n39), .B(n40), .Z(n16) );
  ANDN U390 ( .B(n41), .A(n42), .Z(n39) );
  XOR U391 ( .A(n40), .B(n43), .Z(n41) );
  XOR U392 ( .A(n44), .B(n45), .Z(n37) );
  ANDN U393 ( .B(n46), .A(n17), .Z(n44) );
  XOR U394 ( .A(n45), .B(n18), .Z(n46) );
  XNOR U395 ( .A(n47), .B(n48), .Z(n43) );
  ANDN U396 ( .B(n49), .A(n50), .Z(n47) );
  XOR U397 ( .A(n51), .B(n52), .Z(n49) );
  XNOR U398 ( .A(n54), .B(n55), .Z(n53) );
  ANDN U399 ( .B(n56), .A(n57), .Z(n54) );
  XNOR U400 ( .A(n58), .B(n59), .Z(n56) );
  XOR U401 ( .A(n60), .B(n61), .Z(n40) );
  ANDN U402 ( .B(n62), .A(n63), .Z(n60) );
  XOR U403 ( .A(n61), .B(n64), .Z(n62) );
  XOR U404 ( .A(n65), .B(n66), .Z(n45) );
  ANDN U405 ( .B(n67), .A(n19), .Z(n65) );
  XOR U406 ( .A(n66), .B(n20), .Z(n67) );
  XNOR U407 ( .A(n68), .B(n69), .Z(n52) );
  ANDN U408 ( .B(n70), .A(n71), .Z(n68) );
  XOR U409 ( .A(n72), .B(n73), .Z(n70) );
  XOR U410 ( .A(n48), .B(n74), .Z(n50) );
  XNOR U411 ( .A(n75), .B(n76), .Z(n74) );
  ANDN U412 ( .B(n77), .A(n78), .Z(n75) );
  XNOR U413 ( .A(n79), .B(n80), .Z(n77) );
  IV U414 ( .A(n51), .Z(n48) );
  XOR U415 ( .A(n81), .B(n82), .Z(n51) );
  ANDN U416 ( .B(n83), .A(n84), .Z(n81) );
  XOR U417 ( .A(n82), .B(n85), .Z(n83) );
  XNOR U418 ( .A(n58), .B(n87), .Z(n86) );
  IV U419 ( .A(n61), .Z(n87) );
  XOR U420 ( .A(n88), .B(n89), .Z(n61) );
  ANDN U421 ( .B(n90), .A(n91), .Z(n88) );
  XOR U422 ( .A(n89), .B(n92), .Z(n90) );
  XNOR U423 ( .A(n93), .B(n94), .Z(n58) );
  ANDN U424 ( .B(n95), .A(n96), .Z(n93) );
  XOR U425 ( .A(n94), .B(n97), .Z(n95) );
  XOR U426 ( .A(n55), .B(n98), .Z(n57) );
  XNOR U427 ( .A(n99), .B(n100), .Z(n98) );
  ANDN U428 ( .B(n101), .A(n102), .Z(n99) );
  XNOR U429 ( .A(n103), .B(n104), .Z(n101) );
  IV U430 ( .A(n59), .Z(n55) );
  XOR U431 ( .A(n105), .B(n106), .Z(n59) );
  ANDN U432 ( .B(n107), .A(n108), .Z(n105) );
  XOR U433 ( .A(n109), .B(n106), .Z(n107) );
  XOR U434 ( .A(n110), .B(n111), .Z(n66) );
  ANDN U435 ( .B(n112), .A(n21), .Z(n110) );
  XOR U436 ( .A(n111), .B(n22), .Z(n112) );
  XNOR U437 ( .A(n113), .B(n114), .Z(n73) );
  ANDN U438 ( .B(n115), .A(n116), .Z(n113) );
  XOR U439 ( .A(n117), .B(n118), .Z(n115) );
  XOR U440 ( .A(n69), .B(n119), .Z(n71) );
  XNOR U441 ( .A(n120), .B(n121), .Z(n119) );
  ANDN U442 ( .B(n122), .A(n123), .Z(n120) );
  XNOR U443 ( .A(n124), .B(n125), .Z(n122) );
  IV U444 ( .A(n72), .Z(n69) );
  XOR U445 ( .A(n126), .B(n127), .Z(n72) );
  ANDN U446 ( .B(n128), .A(n129), .Z(n126) );
  XOR U447 ( .A(n127), .B(n130), .Z(n128) );
  XOR U448 ( .A(n131), .B(n132), .Z(n84) );
  XNOR U449 ( .A(n79), .B(n133), .Z(n132) );
  IV U450 ( .A(n82), .Z(n133) );
  XOR U451 ( .A(n134), .B(n135), .Z(n82) );
  ANDN U452 ( .B(n136), .A(n137), .Z(n134) );
  XOR U453 ( .A(n135), .B(n138), .Z(n136) );
  XNOR U454 ( .A(n139), .B(n140), .Z(n79) );
  ANDN U455 ( .B(n141), .A(n142), .Z(n139) );
  XOR U456 ( .A(n140), .B(n143), .Z(n141) );
  IV U457 ( .A(n78), .Z(n131) );
  XOR U458 ( .A(n76), .B(n144), .Z(n78) );
  XNOR U459 ( .A(n145), .B(n146), .Z(n144) );
  ANDN U460 ( .B(n147), .A(n148), .Z(n145) );
  XNOR U461 ( .A(n149), .B(n150), .Z(n147) );
  IV U462 ( .A(n80), .Z(n76) );
  XOR U463 ( .A(n151), .B(n152), .Z(n80) );
  ANDN U464 ( .B(n153), .A(n154), .Z(n151) );
  XOR U465 ( .A(n155), .B(n152), .Z(n153) );
  XOR U466 ( .A(n109), .B(n157), .Z(n156) );
  IV U467 ( .A(n89), .Z(n157) );
  XOR U468 ( .A(n158), .B(n159), .Z(n89) );
  ANDN U469 ( .B(n160), .A(n161), .Z(n158) );
  XOR U470 ( .A(n159), .B(n162), .Z(n160) );
  XNOR U471 ( .A(n163), .B(n164), .Z(n97) );
  ANDN U472 ( .B(n165), .A(n166), .Z(n163) );
  XOR U473 ( .A(n167), .B(n168), .Z(n165) );
  XOR U474 ( .A(n169), .B(n170), .Z(n96) );
  XNOR U475 ( .A(n171), .B(n172), .Z(n170) );
  ANDN U476 ( .B(n173), .A(n174), .Z(n171) );
  XNOR U477 ( .A(n175), .B(n176), .Z(n173) );
  IV U478 ( .A(n94), .Z(n169) );
  XOR U479 ( .A(n177), .B(n178), .Z(n94) );
  ANDN U480 ( .B(n179), .A(n180), .Z(n177) );
  XOR U481 ( .A(n178), .B(n181), .Z(n179) );
  XNOR U482 ( .A(n103), .B(n183), .Z(n182) );
  IV U483 ( .A(n106), .Z(n183) );
  XOR U484 ( .A(n184), .B(n185), .Z(n106) );
  ANDN U485 ( .B(n186), .A(n187), .Z(n184) );
  XOR U486 ( .A(n188), .B(n185), .Z(n186) );
  XNOR U487 ( .A(n189), .B(n190), .Z(n103) );
  ANDN U488 ( .B(n191), .A(n192), .Z(n189) );
  XOR U489 ( .A(n190), .B(n193), .Z(n191) );
  XOR U490 ( .A(n100), .B(n194), .Z(n102) );
  XNOR U491 ( .A(n195), .B(n196), .Z(n194) );
  ANDN U492 ( .B(n197), .A(n198), .Z(n195) );
  XNOR U493 ( .A(n199), .B(n200), .Z(n197) );
  IV U494 ( .A(n104), .Z(n100) );
  XOR U495 ( .A(n201), .B(n202), .Z(n104) );
  ANDN U496 ( .B(n203), .A(n204), .Z(n201) );
  XOR U497 ( .A(n205), .B(n202), .Z(n203) );
  XOR U498 ( .A(n206), .B(n207), .Z(n111) );
  ANDN U499 ( .B(n208), .A(n23), .Z(n206) );
  XOR U500 ( .A(n207), .B(n24), .Z(n208) );
  XNOR U501 ( .A(n209), .B(n210), .Z(n118) );
  ANDN U502 ( .B(n211), .A(n212), .Z(n209) );
  XNOR U503 ( .A(n210), .B(n213), .Z(n211) );
  XOR U504 ( .A(n114), .B(n214), .Z(n116) );
  XNOR U505 ( .A(n215), .B(n216), .Z(n214) );
  ANDN U506 ( .B(n217), .A(n218), .Z(n215) );
  XNOR U507 ( .A(n219), .B(n220), .Z(n217) );
  IV U508 ( .A(n117), .Z(n114) );
  XOR U509 ( .A(n221), .B(n222), .Z(n117) );
  ANDN U510 ( .B(n223), .A(n224), .Z(n221) );
  XOR U511 ( .A(n222), .B(n225), .Z(n223) );
  XOR U512 ( .A(n226), .B(n227), .Z(n129) );
  XNOR U513 ( .A(n124), .B(n228), .Z(n227) );
  IV U514 ( .A(n127), .Z(n228) );
  XOR U515 ( .A(n229), .B(n230), .Z(n127) );
  ANDN U516 ( .B(n231), .A(n232), .Z(n229) );
  XOR U517 ( .A(n230), .B(n233), .Z(n231) );
  XOR U518 ( .A(n234), .B(n235), .Z(n124) );
  ANDN U519 ( .B(n236), .A(n237), .Z(n234) );
  XNOR U520 ( .A(n235), .B(n238), .Z(n236) );
  IV U521 ( .A(n123), .Z(n226) );
  XOR U522 ( .A(n121), .B(n239), .Z(n123) );
  XNOR U523 ( .A(n240), .B(n241), .Z(n239) );
  ANDN U524 ( .B(n242), .A(n243), .Z(n240) );
  XNOR U525 ( .A(n244), .B(n245), .Z(n242) );
  IV U526 ( .A(n125), .Z(n121) );
  XOR U527 ( .A(n246), .B(n247), .Z(n125) );
  ANDN U528 ( .B(n248), .A(n249), .Z(n246) );
  XOR U529 ( .A(n250), .B(n247), .Z(n248) );
  XOR U530 ( .A(n155), .B(n252), .Z(n251) );
  IV U531 ( .A(n135), .Z(n252) );
  XOR U532 ( .A(n253), .B(n254), .Z(n135) );
  ANDN U533 ( .B(n255), .A(n256), .Z(n253) );
  XOR U534 ( .A(n254), .B(n257), .Z(n255) );
  XNOR U535 ( .A(n258), .B(n259), .Z(n143) );
  ANDN U536 ( .B(n260), .A(n261), .Z(n258) );
  XNOR U537 ( .A(n259), .B(n262), .Z(n260) );
  XNOR U538 ( .A(n264), .B(n265), .Z(n263) );
  ANDN U539 ( .B(n266), .A(n267), .Z(n264) );
  XNOR U540 ( .A(n268), .B(n269), .Z(n266) );
  XOR U541 ( .A(n270), .B(n271), .Z(n140) );
  ANDN U542 ( .B(n272), .A(n273), .Z(n270) );
  XOR U543 ( .A(n271), .B(n274), .Z(n272) );
  XNOR U544 ( .A(n149), .B(n276), .Z(n275) );
  IV U545 ( .A(n152), .Z(n276) );
  XOR U546 ( .A(n277), .B(n278), .Z(n152) );
  ANDN U547 ( .B(n279), .A(n280), .Z(n277) );
  XOR U548 ( .A(n281), .B(n278), .Z(n279) );
  XOR U549 ( .A(n282), .B(n283), .Z(n149) );
  ANDN U550 ( .B(n284), .A(n285), .Z(n282) );
  XNOR U551 ( .A(n283), .B(n286), .Z(n284) );
  XOR U552 ( .A(n146), .B(n287), .Z(n148) );
  XNOR U553 ( .A(n288), .B(n289), .Z(n287) );
  ANDN U554 ( .B(n290), .A(n291), .Z(n288) );
  XNOR U555 ( .A(n292), .B(n293), .Z(n290) );
  IV U556 ( .A(n150), .Z(n146) );
  XOR U557 ( .A(n294), .B(n295), .Z(n150) );
  ANDN U558 ( .B(n296), .A(n297), .Z(n294) );
  XOR U559 ( .A(n298), .B(n295), .Z(n296) );
  XOR U560 ( .A(n188), .B(n300), .Z(n299) );
  IV U561 ( .A(n159), .Z(n300) );
  XOR U562 ( .A(n301), .B(n302), .Z(n159) );
  ANDN U563 ( .B(n303), .A(n304), .Z(n301) );
  XOR U564 ( .A(n302), .B(n305), .Z(n303) );
  XNOR U565 ( .A(n306), .B(n307), .Z(n168) );
  ANDN U566 ( .B(n308), .A(n309), .Z(n306) );
  XNOR U567 ( .A(n307), .B(n310), .Z(n308) );
  XOR U568 ( .A(n164), .B(n311), .Z(n166) );
  XNOR U569 ( .A(n312), .B(n313), .Z(n311) );
  ANDN U570 ( .B(n314), .A(n315), .Z(n312) );
  XNOR U571 ( .A(n316), .B(n317), .Z(n314) );
  IV U572 ( .A(n167), .Z(n164) );
  XOR U573 ( .A(n318), .B(n319), .Z(n167) );
  ANDN U574 ( .B(n320), .A(n321), .Z(n318) );
  XOR U575 ( .A(n319), .B(n322), .Z(n320) );
  XOR U576 ( .A(n323), .B(n324), .Z(n180) );
  XNOR U577 ( .A(n175), .B(n325), .Z(n324) );
  IV U578 ( .A(n178), .Z(n325) );
  XOR U579 ( .A(n326), .B(n327), .Z(n178) );
  ANDN U580 ( .B(n328), .A(n329), .Z(n326) );
  XOR U581 ( .A(n327), .B(n330), .Z(n328) );
  XOR U582 ( .A(n331), .B(n332), .Z(n175) );
  ANDN U583 ( .B(n333), .A(n334), .Z(n331) );
  XNOR U584 ( .A(n332), .B(n335), .Z(n333) );
  IV U585 ( .A(n174), .Z(n323) );
  XOR U586 ( .A(n172), .B(n336), .Z(n174) );
  XNOR U587 ( .A(n337), .B(n338), .Z(n336) );
  ANDN U588 ( .B(n339), .A(n340), .Z(n337) );
  XNOR U589 ( .A(n341), .B(n342), .Z(n339) );
  IV U590 ( .A(n176), .Z(n172) );
  XOR U591 ( .A(n343), .B(n344), .Z(n176) );
  ANDN U592 ( .B(n345), .A(n346), .Z(n343) );
  XOR U593 ( .A(n347), .B(n344), .Z(n345) );
  XOR U594 ( .A(n348), .B(n349), .Z(n187) );
  XOR U595 ( .A(n205), .B(n350), .Z(n349) );
  IV U596 ( .A(n185), .Z(n350) );
  XOR U597 ( .A(n351), .B(n352), .Z(n185) );
  ANDN U598 ( .B(n353), .A(n354), .Z(n351) );
  XOR U599 ( .A(n355), .B(n352), .Z(n353) );
  XNOR U600 ( .A(n356), .B(n357), .Z(n193) );
  ANDN U601 ( .B(n358), .A(n359), .Z(n356) );
  XNOR U602 ( .A(n357), .B(n360), .Z(n358) );
  XNOR U603 ( .A(n362), .B(n363), .Z(n361) );
  ANDN U604 ( .B(n364), .A(n365), .Z(n362) );
  XNOR U605 ( .A(n366), .B(n367), .Z(n364) );
  XOR U606 ( .A(n368), .B(n369), .Z(n190) );
  ANDN U607 ( .B(n370), .A(n371), .Z(n368) );
  XOR U608 ( .A(n369), .B(n372), .Z(n370) );
  IV U609 ( .A(n204), .Z(n348) );
  XNOR U610 ( .A(n199), .B(n374), .Z(n373) );
  IV U611 ( .A(n202), .Z(n374) );
  XOR U612 ( .A(n375), .B(n376), .Z(n202) );
  ANDN U613 ( .B(n377), .A(n378), .Z(n375) );
  XOR U614 ( .A(n379), .B(n376), .Z(n377) );
  XOR U615 ( .A(n380), .B(n381), .Z(n199) );
  ANDN U616 ( .B(n382), .A(n383), .Z(n380) );
  XNOR U617 ( .A(n381), .B(n384), .Z(n382) );
  XOR U618 ( .A(n196), .B(n385), .Z(n198) );
  XNOR U619 ( .A(n386), .B(n387), .Z(n385) );
  ANDN U620 ( .B(n388), .A(n389), .Z(n386) );
  XNOR U621 ( .A(n390), .B(n391), .Z(n388) );
  IV U622 ( .A(n200), .Z(n196) );
  XOR U623 ( .A(n392), .B(n393), .Z(n200) );
  ANDN U624 ( .B(n394), .A(n395), .Z(n392) );
  XOR U625 ( .A(n396), .B(n393), .Z(n394) );
  XOR U626 ( .A(n397), .B(n398), .Z(n207) );
  ANDN U627 ( .B(n399), .A(n25), .Z(n397) );
  XOR U628 ( .A(n398), .B(n26), .Z(n399) );
  XNOR U629 ( .A(n400), .B(n401), .Z(n213) );
  NANDN U630 ( .A(n402), .B(n403), .Z(n401) );
  NANDN U631 ( .A(n404), .B(n400), .Z(n403) );
  XNOR U632 ( .A(n405), .B(n210), .Z(n212) );
  XNOR U633 ( .A(n406), .B(n407), .Z(n210) );
  NAND U634 ( .A(n408), .B(n409), .Z(n407) );
  XNOR U635 ( .A(n406), .B(n410), .Z(n408) );
  NOR U636 ( .A(n411), .B(n412), .Z(n405) );
  XOR U637 ( .A(n413), .B(n414), .Z(n224) );
  XOR U638 ( .A(n219), .B(n222), .Z(n414) );
  XNOR U639 ( .A(n415), .B(n416), .Z(n222) );
  NANDN U640 ( .A(n417), .B(n418), .Z(n416) );
  XOR U641 ( .A(n415), .B(n419), .Z(n418) );
  XNOR U642 ( .A(n420), .B(n421), .Z(n219) );
  NANDN U643 ( .A(n422), .B(n423), .Z(n421) );
  NANDN U644 ( .A(n420), .B(n424), .Z(n423) );
  IV U645 ( .A(n218), .Z(n413) );
  XOR U646 ( .A(n425), .B(n220), .Z(n218) );
  IV U647 ( .A(n216), .Z(n220) );
  XNOR U648 ( .A(n426), .B(n427), .Z(n216) );
  NAND U649 ( .A(n428), .B(n429), .Z(n427) );
  XOR U650 ( .A(n426), .B(n430), .Z(n428) );
  NOR U651 ( .A(n431), .B(n432), .Z(n425) );
  XNOR U652 ( .A(n250), .B(n230), .Z(n433) );
  XNOR U653 ( .A(n434), .B(n435), .Z(n230) );
  NANDN U654 ( .A(n436), .B(n437), .Z(n435) );
  XOR U655 ( .A(n434), .B(n438), .Z(n437) );
  XNOR U656 ( .A(n439), .B(n440), .Z(n238) );
  NANDN U657 ( .A(n441), .B(n442), .Z(n440) );
  NANDN U658 ( .A(n443), .B(n439), .Z(n442) );
  XNOR U659 ( .A(n444), .B(n235), .Z(n237) );
  XNOR U660 ( .A(n445), .B(n446), .Z(n235) );
  NAND U661 ( .A(n447), .B(n448), .Z(n446) );
  XNOR U662 ( .A(n445), .B(n449), .Z(n447) );
  NOR U663 ( .A(n450), .B(n451), .Z(n444) );
  XOR U664 ( .A(n244), .B(n247), .Z(n452) );
  XNOR U665 ( .A(n453), .B(n454), .Z(n247) );
  NANDN U666 ( .A(n455), .B(n456), .Z(n454) );
  XNOR U667 ( .A(n453), .B(n457), .Z(n456) );
  XNOR U668 ( .A(n458), .B(n459), .Z(n244) );
  NANDN U669 ( .A(n460), .B(n461), .Z(n459) );
  NANDN U670 ( .A(n458), .B(n462), .Z(n461) );
  XOR U671 ( .A(n463), .B(n245), .Z(n243) );
  IV U672 ( .A(n241), .Z(n245) );
  XNOR U673 ( .A(n464), .B(n465), .Z(n241) );
  NAND U674 ( .A(n466), .B(n467), .Z(n465) );
  XOR U675 ( .A(n464), .B(n468), .Z(n466) );
  NOR U676 ( .A(n469), .B(n470), .Z(n463) );
  XNOR U677 ( .A(n281), .B(n254), .Z(n471) );
  XNOR U678 ( .A(n472), .B(n473), .Z(n254) );
  NANDN U679 ( .A(n474), .B(n475), .Z(n473) );
  XOR U680 ( .A(n472), .B(n476), .Z(n475) );
  XNOR U681 ( .A(n477), .B(n478), .Z(n262) );
  NANDN U682 ( .A(n479), .B(n480), .Z(n478) );
  NANDN U683 ( .A(n481), .B(n477), .Z(n480) );
  XNOR U684 ( .A(n482), .B(n259), .Z(n261) );
  XNOR U685 ( .A(n483), .B(n484), .Z(n259) );
  NAND U686 ( .A(n485), .B(n486), .Z(n484) );
  XNOR U687 ( .A(n483), .B(n487), .Z(n485) );
  NOR U688 ( .A(n488), .B(n489), .Z(n482) );
  XOR U689 ( .A(n268), .B(n271), .Z(n490) );
  XNOR U690 ( .A(n491), .B(n492), .Z(n271) );
  NANDN U691 ( .A(n493), .B(n494), .Z(n492) );
  XOR U692 ( .A(n491), .B(n495), .Z(n494) );
  XNOR U693 ( .A(n496), .B(n497), .Z(n268) );
  NANDN U694 ( .A(n498), .B(n499), .Z(n497) );
  NANDN U695 ( .A(n496), .B(n500), .Z(n499) );
  XOR U696 ( .A(n501), .B(n269), .Z(n267) );
  IV U697 ( .A(n265), .Z(n269) );
  XNOR U698 ( .A(n502), .B(n503), .Z(n265) );
  NAND U699 ( .A(n504), .B(n505), .Z(n503) );
  XOR U700 ( .A(n502), .B(n506), .Z(n504) );
  NOR U701 ( .A(n507), .B(n508), .Z(n501) );
  XNOR U702 ( .A(n298), .B(n278), .Z(n509) );
  XNOR U703 ( .A(n510), .B(n511), .Z(n278) );
  NANDN U704 ( .A(n512), .B(n513), .Z(n511) );
  XOR U705 ( .A(n510), .B(n514), .Z(n513) );
  XNOR U706 ( .A(n515), .B(n516), .Z(n286) );
  NANDN U707 ( .A(n517), .B(n518), .Z(n516) );
  NANDN U708 ( .A(n519), .B(n515), .Z(n518) );
  XNOR U709 ( .A(n520), .B(n283), .Z(n285) );
  XNOR U710 ( .A(n521), .B(n522), .Z(n283) );
  NAND U711 ( .A(n523), .B(n524), .Z(n522) );
  XNOR U712 ( .A(n521), .B(n525), .Z(n523) );
  NOR U713 ( .A(n526), .B(n527), .Z(n520) );
  XOR U714 ( .A(n292), .B(n295), .Z(n528) );
  XNOR U715 ( .A(n529), .B(n530), .Z(n295) );
  NANDN U716 ( .A(n531), .B(n532), .Z(n530) );
  XNOR U717 ( .A(n529), .B(n533), .Z(n532) );
  XNOR U718 ( .A(n534), .B(n535), .Z(n292) );
  NANDN U719 ( .A(n536), .B(n537), .Z(n535) );
  NANDN U720 ( .A(n534), .B(n538), .Z(n537) );
  XOR U721 ( .A(n539), .B(n293), .Z(n291) );
  IV U722 ( .A(n289), .Z(n293) );
  XNOR U723 ( .A(n540), .B(n541), .Z(n289) );
  NAND U724 ( .A(n542), .B(n543), .Z(n541) );
  XOR U725 ( .A(n540), .B(n544), .Z(n542) );
  NOR U726 ( .A(n545), .B(n546), .Z(n539) );
  XNOR U727 ( .A(n355), .B(n302), .Z(n547) );
  XNOR U728 ( .A(n548), .B(n549), .Z(n302) );
  NANDN U729 ( .A(n550), .B(n551), .Z(n549) );
  XOR U730 ( .A(n548), .B(n552), .Z(n551) );
  XNOR U731 ( .A(n553), .B(n554), .Z(n310) );
  NANDN U732 ( .A(n555), .B(n556), .Z(n554) );
  NANDN U733 ( .A(n557), .B(n553), .Z(n556) );
  XNOR U734 ( .A(n558), .B(n307), .Z(n309) );
  XNOR U735 ( .A(n559), .B(n560), .Z(n307) );
  NAND U736 ( .A(n561), .B(n562), .Z(n560) );
  XNOR U737 ( .A(n559), .B(n563), .Z(n561) );
  NOR U738 ( .A(n564), .B(n565), .Z(n558) );
  XOR U739 ( .A(n316), .B(n319), .Z(n566) );
  XNOR U740 ( .A(n567), .B(n568), .Z(n319) );
  NANDN U741 ( .A(n569), .B(n570), .Z(n568) );
  XOR U742 ( .A(n567), .B(n571), .Z(n570) );
  XNOR U743 ( .A(n572), .B(n573), .Z(n316) );
  NANDN U744 ( .A(n574), .B(n575), .Z(n573) );
  NANDN U745 ( .A(n572), .B(n576), .Z(n575) );
  XOR U746 ( .A(n577), .B(n317), .Z(n315) );
  IV U747 ( .A(n313), .Z(n317) );
  XNOR U748 ( .A(n578), .B(n579), .Z(n313) );
  NAND U749 ( .A(n580), .B(n581), .Z(n579) );
  XOR U750 ( .A(n578), .B(n582), .Z(n580) );
  NOR U751 ( .A(n583), .B(n584), .Z(n577) );
  XNOR U752 ( .A(n347), .B(n327), .Z(n585) );
  XNOR U753 ( .A(n586), .B(n587), .Z(n327) );
  NANDN U754 ( .A(n588), .B(n589), .Z(n587) );
  XOR U755 ( .A(n586), .B(n590), .Z(n589) );
  XNOR U756 ( .A(n591), .B(n592), .Z(n335) );
  NANDN U757 ( .A(n593), .B(n594), .Z(n592) );
  NANDN U758 ( .A(n595), .B(n591), .Z(n594) );
  XNOR U759 ( .A(n596), .B(n332), .Z(n334) );
  XNOR U760 ( .A(n597), .B(n598), .Z(n332) );
  NAND U761 ( .A(n599), .B(n600), .Z(n598) );
  XNOR U762 ( .A(n597), .B(n601), .Z(n599) );
  NOR U763 ( .A(n602), .B(n603), .Z(n596) );
  XOR U764 ( .A(n341), .B(n344), .Z(n604) );
  XNOR U765 ( .A(n605), .B(n606), .Z(n344) );
  NANDN U766 ( .A(n607), .B(n608), .Z(n606) );
  XNOR U767 ( .A(n605), .B(n609), .Z(n608) );
  XNOR U768 ( .A(n610), .B(n611), .Z(n341) );
  NANDN U769 ( .A(n612), .B(n613), .Z(n611) );
  NANDN U770 ( .A(n610), .B(n614), .Z(n613) );
  XOR U771 ( .A(n615), .B(n342), .Z(n340) );
  IV U772 ( .A(n338), .Z(n342) );
  XNOR U773 ( .A(n616), .B(n617), .Z(n338) );
  NAND U774 ( .A(n618), .B(n619), .Z(n617) );
  XOR U775 ( .A(n616), .B(n620), .Z(n618) );
  NOR U776 ( .A(n621), .B(n622), .Z(n615) );
  XNOR U777 ( .A(n379), .B(n352), .Z(n623) );
  XNOR U778 ( .A(n624), .B(n625), .Z(n352) );
  NANDN U779 ( .A(n626), .B(n627), .Z(n625) );
  XOR U780 ( .A(n624), .B(n628), .Z(n627) );
  XNOR U781 ( .A(n629), .B(n630), .Z(n360) );
  NANDN U782 ( .A(n631), .B(n632), .Z(n630) );
  NANDN U783 ( .A(n633), .B(n629), .Z(n632) );
  XNOR U784 ( .A(n634), .B(n357), .Z(n359) );
  XNOR U785 ( .A(n635), .B(n636), .Z(n357) );
  NAND U786 ( .A(n637), .B(n638), .Z(n636) );
  XNOR U787 ( .A(n635), .B(n639), .Z(n637) );
  NOR U788 ( .A(n640), .B(n641), .Z(n634) );
  XOR U789 ( .A(n366), .B(n369), .Z(n642) );
  XNOR U790 ( .A(n643), .B(n644), .Z(n369) );
  NANDN U791 ( .A(n645), .B(n646), .Z(n644) );
  XOR U792 ( .A(n643), .B(n647), .Z(n646) );
  XNOR U793 ( .A(n648), .B(n649), .Z(n366) );
  NANDN U794 ( .A(n650), .B(n651), .Z(n649) );
  NANDN U795 ( .A(n648), .B(n652), .Z(n651) );
  XOR U796 ( .A(n653), .B(n367), .Z(n365) );
  IV U797 ( .A(n363), .Z(n367) );
  XNOR U798 ( .A(n654), .B(n655), .Z(n363) );
  NAND U799 ( .A(n656), .B(n657), .Z(n655) );
  XOR U800 ( .A(n654), .B(n658), .Z(n656) );
  NOR U801 ( .A(n659), .B(n660), .Z(n653) );
  XNOR U802 ( .A(n396), .B(n376), .Z(n661) );
  XNOR U803 ( .A(n662), .B(n663), .Z(n376) );
  NANDN U804 ( .A(n664), .B(n665), .Z(n663) );
  XOR U805 ( .A(n662), .B(n666), .Z(n665) );
  XNOR U806 ( .A(n667), .B(n668), .Z(n384) );
  NANDN U807 ( .A(n669), .B(n670), .Z(n668) );
  NANDN U808 ( .A(n671), .B(n667), .Z(n670) );
  XNOR U809 ( .A(n672), .B(n381), .Z(n383) );
  XNOR U810 ( .A(n673), .B(n674), .Z(n381) );
  NAND U811 ( .A(n675), .B(n676), .Z(n674) );
  XNOR U812 ( .A(n673), .B(n677), .Z(n675) );
  NOR U813 ( .A(n678), .B(n679), .Z(n672) );
  XOR U814 ( .A(n390), .B(n393), .Z(n680) );
  XNOR U815 ( .A(n681), .B(n682), .Z(n393) );
  NANDN U816 ( .A(n683), .B(n684), .Z(n682) );
  XNOR U817 ( .A(n681), .B(n685), .Z(n684) );
  XNOR U818 ( .A(n686), .B(n687), .Z(n390) );
  NANDN U819 ( .A(n688), .B(n689), .Z(n687) );
  NANDN U820 ( .A(n686), .B(n690), .Z(n689) );
  XOR U821 ( .A(n691), .B(n391), .Z(n389) );
  IV U822 ( .A(n387), .Z(n391) );
  XNOR U823 ( .A(n692), .B(n693), .Z(n387) );
  NAND U824 ( .A(n694), .B(n695), .Z(n693) );
  XOR U825 ( .A(n692), .B(n696), .Z(n694) );
  NOR U826 ( .A(n697), .B(n698), .Z(n691) );
  XOR U827 ( .A(n699), .B(n700), .Z(n398) );
  NANDN U828 ( .A(n27), .B(n701), .Z(n700) );
  XNOR U829 ( .A(n699), .B(n28), .Z(n701) );
  XOR U830 ( .A(n409), .B(n410), .Z(n419) );
  XOR U831 ( .A(n404), .B(n402), .Z(n410) );
  AND U832 ( .A(n702), .B(n400), .Z(n402) );
  OR U833 ( .A(n703), .B(n704), .Z(n400) );
  OR U834 ( .A(n705), .B(n706), .Z(n702) );
  NOR U835 ( .A(n707), .B(n708), .Z(n404) );
  XOR U836 ( .A(n411), .B(n709), .Z(n409) );
  XOR U837 ( .A(n412), .B(n406), .Z(n709) );
  NOR U838 ( .A(n710), .B(n711), .Z(n406) );
  OR U839 ( .A(n712), .B(n713), .Z(n412) );
  AND U840 ( .A(n714), .B(n715), .Z(n411) );
  OR U841 ( .A(n716), .B(n717), .Z(n715) );
  OR U842 ( .A(n718), .B(n719), .Z(n714) );
  XNOR U843 ( .A(n429), .B(n720), .Z(n417) );
  XNOR U844 ( .A(n415), .B(n430), .Z(n720) );
  XOR U845 ( .A(n424), .B(n422), .Z(n430) );
  NOR U846 ( .A(n722), .B(n723), .Z(n420) );
  OR U847 ( .A(n724), .B(n725), .Z(n721) );
  OR U848 ( .A(n726), .B(n727), .Z(n424) );
  OR U849 ( .A(n728), .B(n729), .Z(n415) );
  XOR U850 ( .A(n431), .B(n730), .Z(n429) );
  XOR U851 ( .A(n432), .B(n426), .Z(n730) );
  NOR U852 ( .A(n731), .B(n732), .Z(n426) );
  OR U853 ( .A(n733), .B(n734), .Z(n432) );
  AND U854 ( .A(n735), .B(n736), .Z(n431) );
  OR U855 ( .A(n737), .B(n738), .Z(n736) );
  OR U856 ( .A(n739), .B(n740), .Z(n735) );
  XOR U857 ( .A(n434), .B(n457), .Z(n741) );
  XNOR U858 ( .A(n448), .B(n449), .Z(n457) );
  XOR U859 ( .A(n443), .B(n441), .Z(n449) );
  AND U860 ( .A(n742), .B(n439), .Z(n441) );
  OR U861 ( .A(n743), .B(n744), .Z(n439) );
  OR U862 ( .A(n745), .B(n746), .Z(n742) );
  NOR U863 ( .A(n747), .B(n748), .Z(n443) );
  XOR U864 ( .A(n450), .B(n749), .Z(n448) );
  XOR U865 ( .A(n451), .B(n445), .Z(n749) );
  NOR U866 ( .A(n750), .B(n751), .Z(n445) );
  OR U867 ( .A(n752), .B(n753), .Z(n451) );
  AND U868 ( .A(n754), .B(n755), .Z(n450) );
  OR U869 ( .A(n756), .B(n757), .Z(n755) );
  OR U870 ( .A(n758), .B(n759), .Z(n754) );
  OR U871 ( .A(n760), .B(n761), .Z(n434) );
  XNOR U872 ( .A(n467), .B(n762), .Z(n455) );
  XNOR U873 ( .A(n453), .B(n468), .Z(n762) );
  XOR U874 ( .A(n462), .B(n460), .Z(n468) );
  NOR U875 ( .A(n764), .B(n765), .Z(n458) );
  OR U876 ( .A(n766), .B(n767), .Z(n763) );
  OR U877 ( .A(n768), .B(n769), .Z(n462) );
  OR U878 ( .A(n770), .B(n771), .Z(n453) );
  XOR U879 ( .A(n469), .B(n772), .Z(n467) );
  XOR U880 ( .A(n470), .B(n464), .Z(n772) );
  NOR U881 ( .A(n773), .B(n774), .Z(n464) );
  OR U882 ( .A(n775), .B(n776), .Z(n470) );
  AND U883 ( .A(n777), .B(n778), .Z(n469) );
  OR U884 ( .A(n779), .B(n780), .Z(n778) );
  OR U885 ( .A(n781), .B(n782), .Z(n777) );
  XNOR U886 ( .A(n472), .B(n514), .Z(n783) );
  XOR U887 ( .A(n486), .B(n487), .Z(n495) );
  XOR U888 ( .A(n481), .B(n479), .Z(n487) );
  AND U889 ( .A(n784), .B(n477), .Z(n479) );
  OR U890 ( .A(n785), .B(n786), .Z(n477) );
  OR U891 ( .A(n787), .B(n788), .Z(n784) );
  NOR U892 ( .A(n789), .B(n790), .Z(n481) );
  XOR U893 ( .A(n488), .B(n791), .Z(n486) );
  XOR U894 ( .A(n489), .B(n483), .Z(n791) );
  NOR U895 ( .A(n792), .B(n793), .Z(n483) );
  OR U896 ( .A(n794), .B(n795), .Z(n489) );
  AND U897 ( .A(n796), .B(n797), .Z(n488) );
  OR U898 ( .A(n798), .B(n799), .Z(n797) );
  OR U899 ( .A(n800), .B(n801), .Z(n796) );
  XNOR U900 ( .A(n505), .B(n802), .Z(n493) );
  XNOR U901 ( .A(n491), .B(n506), .Z(n802) );
  XOR U902 ( .A(n500), .B(n498), .Z(n506) );
  NOR U903 ( .A(n804), .B(n805), .Z(n496) );
  OR U904 ( .A(n806), .B(n807), .Z(n803) );
  OR U905 ( .A(n808), .B(n809), .Z(n500) );
  OR U906 ( .A(n810), .B(n811), .Z(n491) );
  XOR U907 ( .A(n507), .B(n812), .Z(n505) );
  XOR U908 ( .A(n508), .B(n502), .Z(n812) );
  NOR U909 ( .A(n813), .B(n814), .Z(n502) );
  OR U910 ( .A(n815), .B(n816), .Z(n508) );
  AND U911 ( .A(n817), .B(n818), .Z(n507) );
  OR U912 ( .A(n819), .B(n820), .Z(n818) );
  OR U913 ( .A(n821), .B(n822), .Z(n817) );
  OR U914 ( .A(n823), .B(n824), .Z(n472) );
  XOR U915 ( .A(n510), .B(n533), .Z(n825) );
  XNOR U916 ( .A(n524), .B(n525), .Z(n533) );
  XOR U917 ( .A(n519), .B(n517), .Z(n525) );
  AND U918 ( .A(n826), .B(n515), .Z(n517) );
  OR U919 ( .A(n827), .B(n828), .Z(n515) );
  OR U920 ( .A(n829), .B(n830), .Z(n826) );
  NOR U921 ( .A(n831), .B(n832), .Z(n519) );
  XOR U922 ( .A(n526), .B(n833), .Z(n524) );
  XOR U923 ( .A(n527), .B(n521), .Z(n833) );
  NOR U924 ( .A(n834), .B(n835), .Z(n521) );
  OR U925 ( .A(n836), .B(n837), .Z(n527) );
  AND U926 ( .A(n838), .B(n839), .Z(n526) );
  OR U927 ( .A(n840), .B(n841), .Z(n839) );
  OR U928 ( .A(n842), .B(n843), .Z(n838) );
  OR U929 ( .A(n844), .B(n845), .Z(n510) );
  XNOR U930 ( .A(n543), .B(n846), .Z(n531) );
  XNOR U931 ( .A(n529), .B(n544), .Z(n846) );
  XOR U932 ( .A(n538), .B(n536), .Z(n544) );
  NOR U933 ( .A(n848), .B(n849), .Z(n534) );
  OR U934 ( .A(n850), .B(n851), .Z(n847) );
  OR U935 ( .A(n852), .B(n853), .Z(n538) );
  OR U936 ( .A(n854), .B(n855), .Z(n529) );
  XOR U937 ( .A(n545), .B(n856), .Z(n543) );
  XOR U938 ( .A(n546), .B(n540), .Z(n856) );
  NOR U939 ( .A(n857), .B(n858), .Z(n540) );
  OR U940 ( .A(n859), .B(n860), .Z(n546) );
  AND U941 ( .A(n861), .B(n862), .Z(n545) );
  OR U942 ( .A(n863), .B(n864), .Z(n862) );
  OR U943 ( .A(n865), .B(n866), .Z(n861) );
  XNOR U944 ( .A(n548), .B(n628), .Z(n867) );
  XOR U945 ( .A(n562), .B(n563), .Z(n571) );
  XOR U946 ( .A(n557), .B(n555), .Z(n563) );
  AND U947 ( .A(n868), .B(n553), .Z(n555) );
  OR U948 ( .A(n869), .B(n870), .Z(n553) );
  OR U949 ( .A(n871), .B(n872), .Z(n868) );
  NOR U950 ( .A(n873), .B(n874), .Z(n557) );
  XOR U951 ( .A(n564), .B(n875), .Z(n562) );
  XOR U952 ( .A(n565), .B(n559), .Z(n875) );
  NOR U953 ( .A(n876), .B(n877), .Z(n559) );
  OR U954 ( .A(n878), .B(n879), .Z(n565) );
  AND U955 ( .A(n880), .B(n881), .Z(n564) );
  OR U956 ( .A(n882), .B(n883), .Z(n881) );
  OR U957 ( .A(n884), .B(n885), .Z(n880) );
  XNOR U958 ( .A(n581), .B(n886), .Z(n569) );
  XNOR U959 ( .A(n567), .B(n582), .Z(n886) );
  XOR U960 ( .A(n576), .B(n574), .Z(n582) );
  NOR U961 ( .A(n888), .B(n889), .Z(n572) );
  OR U962 ( .A(n890), .B(n891), .Z(n887) );
  OR U963 ( .A(n892), .B(n893), .Z(n576) );
  OR U964 ( .A(n894), .B(n895), .Z(n567) );
  XOR U965 ( .A(n583), .B(n896), .Z(n581) );
  XOR U966 ( .A(n584), .B(n578), .Z(n896) );
  NOR U967 ( .A(n897), .B(n898), .Z(n578) );
  OR U968 ( .A(n899), .B(n900), .Z(n584) );
  AND U969 ( .A(n901), .B(n902), .Z(n583) );
  OR U970 ( .A(n903), .B(n904), .Z(n902) );
  OR U971 ( .A(n905), .B(n906), .Z(n901) );
  XOR U972 ( .A(n586), .B(n609), .Z(n907) );
  XNOR U973 ( .A(n600), .B(n601), .Z(n609) );
  XOR U974 ( .A(n595), .B(n593), .Z(n601) );
  AND U975 ( .A(n908), .B(n591), .Z(n593) );
  OR U976 ( .A(n909), .B(n910), .Z(n591) );
  OR U977 ( .A(n911), .B(n912), .Z(n908) );
  NOR U978 ( .A(n913), .B(n914), .Z(n595) );
  XOR U979 ( .A(n602), .B(n915), .Z(n600) );
  XOR U980 ( .A(n603), .B(n597), .Z(n915) );
  NOR U981 ( .A(n916), .B(n917), .Z(n597) );
  OR U982 ( .A(n918), .B(n919), .Z(n603) );
  AND U983 ( .A(n920), .B(n921), .Z(n602) );
  OR U984 ( .A(n922), .B(n923), .Z(n921) );
  OR U985 ( .A(n924), .B(n925), .Z(n920) );
  OR U986 ( .A(n926), .B(n927), .Z(n586) );
  XNOR U987 ( .A(n619), .B(n928), .Z(n607) );
  XNOR U988 ( .A(n605), .B(n620), .Z(n928) );
  XOR U989 ( .A(n614), .B(n612), .Z(n620) );
  NOR U990 ( .A(n930), .B(n931), .Z(n610) );
  OR U991 ( .A(n932), .B(n933), .Z(n929) );
  OR U992 ( .A(n934), .B(n935), .Z(n614) );
  OR U993 ( .A(n936), .B(n937), .Z(n605) );
  XOR U994 ( .A(n621), .B(n938), .Z(n619) );
  XOR U995 ( .A(n622), .B(n616), .Z(n938) );
  NOR U996 ( .A(n939), .B(n940), .Z(n616) );
  OR U997 ( .A(n941), .B(n942), .Z(n622) );
  AND U998 ( .A(n943), .B(n944), .Z(n621) );
  OR U999 ( .A(n945), .B(n946), .Z(n944) );
  OR U1000 ( .A(n947), .B(n948), .Z(n943) );
  OR U1001 ( .A(n949), .B(n950), .Z(n548) );
  XNOR U1002 ( .A(n624), .B(n666), .Z(n951) );
  XOR U1003 ( .A(n638), .B(n639), .Z(n647) );
  XOR U1004 ( .A(n633), .B(n631), .Z(n639) );
  AND U1005 ( .A(n952), .B(n629), .Z(n631) );
  OR U1006 ( .A(n953), .B(n954), .Z(n629) );
  OR U1007 ( .A(n955), .B(n956), .Z(n952) );
  NOR U1008 ( .A(n957), .B(n958), .Z(n633) );
  XOR U1009 ( .A(n640), .B(n959), .Z(n638) );
  XOR U1010 ( .A(n641), .B(n635), .Z(n959) );
  NOR U1011 ( .A(n960), .B(n961), .Z(n635) );
  OR U1012 ( .A(n962), .B(n963), .Z(n641) );
  AND U1013 ( .A(n964), .B(n965), .Z(n640) );
  OR U1014 ( .A(n966), .B(n967), .Z(n965) );
  OR U1015 ( .A(n968), .B(n969), .Z(n964) );
  XNOR U1016 ( .A(n657), .B(n970), .Z(n645) );
  XNOR U1017 ( .A(n643), .B(n658), .Z(n970) );
  XOR U1018 ( .A(n652), .B(n650), .Z(n658) );
  NOR U1019 ( .A(n972), .B(n973), .Z(n648) );
  OR U1020 ( .A(n974), .B(n975), .Z(n971) );
  OR U1021 ( .A(n976), .B(n977), .Z(n652) );
  OR U1022 ( .A(n978), .B(n979), .Z(n643) );
  XOR U1023 ( .A(n659), .B(n980), .Z(n657) );
  XOR U1024 ( .A(n660), .B(n654), .Z(n980) );
  NOR U1025 ( .A(n981), .B(n982), .Z(n654) );
  OR U1026 ( .A(n983), .B(n984), .Z(n660) );
  AND U1027 ( .A(n985), .B(n986), .Z(n659) );
  OR U1028 ( .A(n987), .B(n988), .Z(n986) );
  OR U1029 ( .A(n989), .B(n990), .Z(n985) );
  OR U1030 ( .A(n991), .B(n992), .Z(n624) );
  XOR U1031 ( .A(n662), .B(n685), .Z(n993) );
  XNOR U1032 ( .A(n676), .B(n677), .Z(n685) );
  XOR U1033 ( .A(n671), .B(n669), .Z(n677) );
  AND U1034 ( .A(n994), .B(n667), .Z(n669) );
  OR U1035 ( .A(n995), .B(n996), .Z(n667) );
  OR U1036 ( .A(n997), .B(n998), .Z(n994) );
  NOR U1037 ( .A(n999), .B(n1000), .Z(n671) );
  XOR U1038 ( .A(n678), .B(n1001), .Z(n676) );
  XOR U1039 ( .A(n679), .B(n673), .Z(n1001) );
  NOR U1040 ( .A(n1002), .B(n1003), .Z(n673) );
  OR U1041 ( .A(n1004), .B(n1005), .Z(n679) );
  AND U1042 ( .A(n1006), .B(n1007), .Z(n678) );
  OR U1043 ( .A(n1008), .B(n1009), .Z(n1007) );
  OR U1044 ( .A(n1010), .B(n1011), .Z(n1006) );
  OR U1045 ( .A(n1012), .B(n1013), .Z(n662) );
  XNOR U1046 ( .A(n695), .B(n1014), .Z(n683) );
  XNOR U1047 ( .A(n681), .B(n696), .Z(n1014) );
  XOR U1048 ( .A(n690), .B(n688), .Z(n696) );
  NOR U1049 ( .A(n1016), .B(n1017), .Z(n686) );
  OR U1050 ( .A(n1018), .B(n1019), .Z(n1015) );
  OR U1051 ( .A(n1020), .B(n1021), .Z(n690) );
  OR U1052 ( .A(n1022), .B(n1023), .Z(n681) );
  XOR U1053 ( .A(n697), .B(n1024), .Z(n695) );
  XOR U1054 ( .A(n698), .B(n692), .Z(n1024) );
  NOR U1055 ( .A(n1025), .B(n1026), .Z(n692) );
  OR U1056 ( .A(n1027), .B(n1028), .Z(n698) );
  AND U1057 ( .A(n1029), .B(n1030), .Z(n697) );
  OR U1058 ( .A(n1031), .B(n1032), .Z(n1030) );
  OR U1059 ( .A(n1033), .B(n1034), .Z(n1029) );
  XNOR U1060 ( .A(oglobal[1]), .B(n699), .Z(n27) );
  ANDN U1061 ( .B(oglobal[0]), .A(n1035), .Z(n699) );
  XNOR U1062 ( .A(oglobal[0]), .B(n1035), .Z(o[0]) );
  XNOR U1063 ( .A(n950), .B(n949), .Z(n1035) );
  XNOR U1064 ( .A(n824), .B(n823), .Z(n949) );
  XNOR U1065 ( .A(n761), .B(n760), .Z(n823) );
  XNOR U1066 ( .A(n729), .B(n728), .Z(n760) );
  XNOR U1067 ( .A(n703), .B(n704), .Z(n710) );
  XNOR U1068 ( .A(n707), .B(n708), .Z(n704) );
  XNOR U1069 ( .A(y[127]), .B(x[127]), .Z(n708) );
  XNOR U1070 ( .A(y[126]), .B(x[126]), .Z(n707) );
  XNOR U1071 ( .A(n705), .B(n706), .Z(n703) );
  XNOR U1072 ( .A(y[125]), .B(x[125]), .Z(n706) );
  XNOR U1073 ( .A(y[124]), .B(x[124]), .Z(n705) );
  XNOR U1074 ( .A(n718), .B(n719), .Z(n711) );
  XNOR U1075 ( .A(n713), .B(n712), .Z(n719) );
  XNOR U1076 ( .A(y[123]), .B(x[123]), .Z(n712) );
  XNOR U1077 ( .A(y[122]), .B(x[122]), .Z(n713) );
  XNOR U1078 ( .A(n716), .B(n717), .Z(n718) );
  XNOR U1079 ( .A(y[121]), .B(x[121]), .Z(n717) );
  XNOR U1080 ( .A(y[120]), .B(x[120]), .Z(n716) );
  XNOR U1081 ( .A(n722), .B(n723), .Z(n731) );
  XNOR U1082 ( .A(n726), .B(n727), .Z(n723) );
  XNOR U1083 ( .A(y[119]), .B(x[119]), .Z(n727) );
  XNOR U1084 ( .A(y[118]), .B(x[118]), .Z(n726) );
  XNOR U1085 ( .A(n724), .B(n725), .Z(n722) );
  XNOR U1086 ( .A(y[117]), .B(x[117]), .Z(n725) );
  XNOR U1087 ( .A(y[116]), .B(x[116]), .Z(n724) );
  XNOR U1088 ( .A(n739), .B(n740), .Z(n732) );
  XNOR U1089 ( .A(n734), .B(n733), .Z(n740) );
  XNOR U1090 ( .A(y[115]), .B(x[115]), .Z(n733) );
  XNOR U1091 ( .A(y[114]), .B(x[114]), .Z(n734) );
  XNOR U1092 ( .A(n737), .B(n738), .Z(n739) );
  XNOR U1093 ( .A(y[113]), .B(x[113]), .Z(n738) );
  XNOR U1094 ( .A(y[112]), .B(x[112]), .Z(n737) );
  XNOR U1095 ( .A(n771), .B(n770), .Z(n761) );
  XNOR U1096 ( .A(n743), .B(n744), .Z(n750) );
  XNOR U1097 ( .A(n747), .B(n748), .Z(n744) );
  XNOR U1098 ( .A(y[111]), .B(x[111]), .Z(n748) );
  XNOR U1099 ( .A(y[110]), .B(x[110]), .Z(n747) );
  XNOR U1100 ( .A(n745), .B(n746), .Z(n743) );
  XNOR U1101 ( .A(y[109]), .B(x[109]), .Z(n746) );
  XNOR U1102 ( .A(y[108]), .B(x[108]), .Z(n745) );
  XNOR U1103 ( .A(n758), .B(n759), .Z(n751) );
  XNOR U1104 ( .A(n753), .B(n752), .Z(n759) );
  XNOR U1105 ( .A(y[107]), .B(x[107]), .Z(n752) );
  XNOR U1106 ( .A(y[106]), .B(x[106]), .Z(n753) );
  XNOR U1107 ( .A(n756), .B(n757), .Z(n758) );
  XNOR U1108 ( .A(y[105]), .B(x[105]), .Z(n757) );
  XNOR U1109 ( .A(y[104]), .B(x[104]), .Z(n756) );
  XNOR U1110 ( .A(n764), .B(n765), .Z(n773) );
  XNOR U1111 ( .A(n768), .B(n769), .Z(n765) );
  XNOR U1112 ( .A(y[103]), .B(x[103]), .Z(n769) );
  XNOR U1113 ( .A(y[102]), .B(x[102]), .Z(n768) );
  XNOR U1114 ( .A(n766), .B(n767), .Z(n764) );
  XNOR U1115 ( .A(y[101]), .B(x[101]), .Z(n767) );
  XNOR U1116 ( .A(y[100]), .B(x[100]), .Z(n766) );
  XNOR U1117 ( .A(n781), .B(n782), .Z(n774) );
  XNOR U1118 ( .A(n776), .B(n775), .Z(n782) );
  XNOR U1119 ( .A(y[99]), .B(x[99]), .Z(n775) );
  XNOR U1120 ( .A(y[98]), .B(x[98]), .Z(n776) );
  XNOR U1121 ( .A(n779), .B(n780), .Z(n781) );
  XNOR U1122 ( .A(y[97]), .B(x[97]), .Z(n780) );
  XNOR U1123 ( .A(y[96]), .B(x[96]), .Z(n779) );
  XNOR U1124 ( .A(n845), .B(n844), .Z(n824) );
  XNOR U1125 ( .A(n811), .B(n810), .Z(n844) );
  XNOR U1126 ( .A(n785), .B(n786), .Z(n792) );
  XNOR U1127 ( .A(n789), .B(n790), .Z(n786) );
  XNOR U1128 ( .A(y[95]), .B(x[95]), .Z(n790) );
  XNOR U1129 ( .A(y[94]), .B(x[94]), .Z(n789) );
  XNOR U1130 ( .A(n787), .B(n788), .Z(n785) );
  XNOR U1131 ( .A(y[93]), .B(x[93]), .Z(n788) );
  XNOR U1132 ( .A(y[92]), .B(x[92]), .Z(n787) );
  XNOR U1133 ( .A(n800), .B(n801), .Z(n793) );
  XNOR U1134 ( .A(n795), .B(n794), .Z(n801) );
  XNOR U1135 ( .A(y[91]), .B(x[91]), .Z(n794) );
  XNOR U1136 ( .A(y[90]), .B(x[90]), .Z(n795) );
  XNOR U1137 ( .A(n798), .B(n799), .Z(n800) );
  XNOR U1138 ( .A(y[89]), .B(x[89]), .Z(n799) );
  XNOR U1139 ( .A(y[88]), .B(x[88]), .Z(n798) );
  XNOR U1140 ( .A(n804), .B(n805), .Z(n813) );
  XNOR U1141 ( .A(n808), .B(n809), .Z(n805) );
  XNOR U1142 ( .A(y[87]), .B(x[87]), .Z(n809) );
  XNOR U1143 ( .A(y[86]), .B(x[86]), .Z(n808) );
  XNOR U1144 ( .A(n806), .B(n807), .Z(n804) );
  XNOR U1145 ( .A(y[85]), .B(x[85]), .Z(n807) );
  XNOR U1146 ( .A(y[84]), .B(x[84]), .Z(n806) );
  XNOR U1147 ( .A(n821), .B(n822), .Z(n814) );
  XNOR U1148 ( .A(n816), .B(n815), .Z(n822) );
  XNOR U1149 ( .A(y[83]), .B(x[83]), .Z(n815) );
  XNOR U1150 ( .A(y[82]), .B(x[82]), .Z(n816) );
  XNOR U1151 ( .A(n819), .B(n820), .Z(n821) );
  XNOR U1152 ( .A(y[81]), .B(x[81]), .Z(n820) );
  XNOR U1153 ( .A(y[80]), .B(x[80]), .Z(n819) );
  XNOR U1154 ( .A(n855), .B(n854), .Z(n845) );
  XNOR U1155 ( .A(n827), .B(n828), .Z(n834) );
  XNOR U1156 ( .A(n831), .B(n832), .Z(n828) );
  XNOR U1157 ( .A(y[79]), .B(x[79]), .Z(n832) );
  XNOR U1158 ( .A(y[78]), .B(x[78]), .Z(n831) );
  XNOR U1159 ( .A(n829), .B(n830), .Z(n827) );
  XNOR U1160 ( .A(y[77]), .B(x[77]), .Z(n830) );
  XNOR U1161 ( .A(y[76]), .B(x[76]), .Z(n829) );
  XNOR U1162 ( .A(n842), .B(n843), .Z(n835) );
  XNOR U1163 ( .A(n837), .B(n836), .Z(n843) );
  XNOR U1164 ( .A(y[75]), .B(x[75]), .Z(n836) );
  XNOR U1165 ( .A(y[74]), .B(x[74]), .Z(n837) );
  XNOR U1166 ( .A(n840), .B(n841), .Z(n842) );
  XNOR U1167 ( .A(y[73]), .B(x[73]), .Z(n841) );
  XNOR U1168 ( .A(y[72]), .B(x[72]), .Z(n840) );
  XNOR U1169 ( .A(n848), .B(n849), .Z(n857) );
  XNOR U1170 ( .A(n852), .B(n853), .Z(n849) );
  XNOR U1171 ( .A(y[71]), .B(x[71]), .Z(n853) );
  XNOR U1172 ( .A(y[70]), .B(x[70]), .Z(n852) );
  XNOR U1173 ( .A(n850), .B(n851), .Z(n848) );
  XNOR U1174 ( .A(y[69]), .B(x[69]), .Z(n851) );
  XNOR U1175 ( .A(y[68]), .B(x[68]), .Z(n850) );
  XNOR U1176 ( .A(n865), .B(n866), .Z(n858) );
  XNOR U1177 ( .A(n860), .B(n859), .Z(n866) );
  XNOR U1178 ( .A(y[67]), .B(x[67]), .Z(n859) );
  XNOR U1179 ( .A(y[66]), .B(x[66]), .Z(n860) );
  XNOR U1180 ( .A(n863), .B(n864), .Z(n865) );
  XNOR U1181 ( .A(y[65]), .B(x[65]), .Z(n864) );
  XNOR U1182 ( .A(y[64]), .B(x[64]), .Z(n863) );
  XNOR U1183 ( .A(n992), .B(n991), .Z(n950) );
  XNOR U1184 ( .A(n927), .B(n926), .Z(n991) );
  XNOR U1185 ( .A(n895), .B(n894), .Z(n926) );
  XNOR U1186 ( .A(n869), .B(n870), .Z(n876) );
  XNOR U1187 ( .A(n873), .B(n874), .Z(n870) );
  XNOR U1188 ( .A(y[63]), .B(x[63]), .Z(n874) );
  XNOR U1189 ( .A(y[62]), .B(x[62]), .Z(n873) );
  XNOR U1190 ( .A(n871), .B(n872), .Z(n869) );
  XNOR U1191 ( .A(y[61]), .B(x[61]), .Z(n872) );
  XNOR U1192 ( .A(y[60]), .B(x[60]), .Z(n871) );
  XNOR U1193 ( .A(n884), .B(n885), .Z(n877) );
  XNOR U1194 ( .A(n879), .B(n878), .Z(n885) );
  XNOR U1195 ( .A(y[59]), .B(x[59]), .Z(n878) );
  XNOR U1196 ( .A(y[58]), .B(x[58]), .Z(n879) );
  XNOR U1197 ( .A(n882), .B(n883), .Z(n884) );
  XNOR U1198 ( .A(y[57]), .B(x[57]), .Z(n883) );
  XNOR U1199 ( .A(y[56]), .B(x[56]), .Z(n882) );
  XNOR U1200 ( .A(n888), .B(n889), .Z(n897) );
  XNOR U1201 ( .A(n892), .B(n893), .Z(n889) );
  XNOR U1202 ( .A(y[55]), .B(x[55]), .Z(n893) );
  XNOR U1203 ( .A(y[54]), .B(x[54]), .Z(n892) );
  XNOR U1204 ( .A(n890), .B(n891), .Z(n888) );
  XNOR U1205 ( .A(y[53]), .B(x[53]), .Z(n891) );
  XNOR U1206 ( .A(y[52]), .B(x[52]), .Z(n890) );
  XNOR U1207 ( .A(n905), .B(n906), .Z(n898) );
  XNOR U1208 ( .A(n900), .B(n899), .Z(n906) );
  XNOR U1209 ( .A(y[51]), .B(x[51]), .Z(n899) );
  XNOR U1210 ( .A(y[50]), .B(x[50]), .Z(n900) );
  XNOR U1211 ( .A(n903), .B(n904), .Z(n905) );
  XNOR U1212 ( .A(y[49]), .B(x[49]), .Z(n904) );
  XNOR U1213 ( .A(y[48]), .B(x[48]), .Z(n903) );
  XNOR U1214 ( .A(n937), .B(n936), .Z(n927) );
  XNOR U1215 ( .A(n909), .B(n910), .Z(n916) );
  XNOR U1216 ( .A(n913), .B(n914), .Z(n910) );
  XNOR U1217 ( .A(y[47]), .B(x[47]), .Z(n914) );
  XNOR U1218 ( .A(y[46]), .B(x[46]), .Z(n913) );
  XNOR U1219 ( .A(n911), .B(n912), .Z(n909) );
  XNOR U1220 ( .A(y[45]), .B(x[45]), .Z(n912) );
  XNOR U1221 ( .A(y[44]), .B(x[44]), .Z(n911) );
  XNOR U1222 ( .A(n924), .B(n925), .Z(n917) );
  XNOR U1223 ( .A(n919), .B(n918), .Z(n925) );
  XNOR U1224 ( .A(y[43]), .B(x[43]), .Z(n918) );
  XNOR U1225 ( .A(y[42]), .B(x[42]), .Z(n919) );
  XNOR U1226 ( .A(n922), .B(n923), .Z(n924) );
  XNOR U1227 ( .A(y[41]), .B(x[41]), .Z(n923) );
  XNOR U1228 ( .A(y[40]), .B(x[40]), .Z(n922) );
  XNOR U1229 ( .A(n930), .B(n931), .Z(n939) );
  XNOR U1230 ( .A(n934), .B(n935), .Z(n931) );
  XNOR U1231 ( .A(y[39]), .B(x[39]), .Z(n935) );
  XNOR U1232 ( .A(y[38]), .B(x[38]), .Z(n934) );
  XNOR U1233 ( .A(n932), .B(n933), .Z(n930) );
  XNOR U1234 ( .A(y[37]), .B(x[37]), .Z(n933) );
  XNOR U1235 ( .A(y[36]), .B(x[36]), .Z(n932) );
  XNOR U1236 ( .A(n947), .B(n948), .Z(n940) );
  XNOR U1237 ( .A(n942), .B(n941), .Z(n948) );
  XNOR U1238 ( .A(y[35]), .B(x[35]), .Z(n941) );
  XNOR U1239 ( .A(y[34]), .B(x[34]), .Z(n942) );
  XNOR U1240 ( .A(n945), .B(n946), .Z(n947) );
  XNOR U1241 ( .A(y[33]), .B(x[33]), .Z(n946) );
  XNOR U1242 ( .A(y[32]), .B(x[32]), .Z(n945) );
  XNOR U1243 ( .A(n1013), .B(n1012), .Z(n992) );
  XNOR U1244 ( .A(n979), .B(n978), .Z(n1012) );
  XNOR U1245 ( .A(n953), .B(n954), .Z(n960) );
  XNOR U1246 ( .A(n957), .B(n958), .Z(n954) );
  XNOR U1247 ( .A(y[31]), .B(x[31]), .Z(n958) );
  XNOR U1248 ( .A(y[30]), .B(x[30]), .Z(n957) );
  XNOR U1249 ( .A(n955), .B(n956), .Z(n953) );
  XNOR U1250 ( .A(y[29]), .B(x[29]), .Z(n956) );
  XNOR U1251 ( .A(y[28]), .B(x[28]), .Z(n955) );
  XNOR U1252 ( .A(n968), .B(n969), .Z(n961) );
  XNOR U1253 ( .A(n963), .B(n962), .Z(n969) );
  XNOR U1254 ( .A(y[27]), .B(x[27]), .Z(n962) );
  XNOR U1255 ( .A(y[26]), .B(x[26]), .Z(n963) );
  XNOR U1256 ( .A(n966), .B(n967), .Z(n968) );
  XNOR U1257 ( .A(y[25]), .B(x[25]), .Z(n967) );
  XNOR U1258 ( .A(y[24]), .B(x[24]), .Z(n966) );
  XNOR U1259 ( .A(n972), .B(n973), .Z(n981) );
  XNOR U1260 ( .A(n976), .B(n977), .Z(n973) );
  XNOR U1261 ( .A(y[23]), .B(x[23]), .Z(n977) );
  XNOR U1262 ( .A(y[22]), .B(x[22]), .Z(n976) );
  XNOR U1263 ( .A(n974), .B(n975), .Z(n972) );
  XNOR U1264 ( .A(y[21]), .B(x[21]), .Z(n975) );
  XNOR U1265 ( .A(y[20]), .B(x[20]), .Z(n974) );
  XNOR U1266 ( .A(n989), .B(n990), .Z(n982) );
  XNOR U1267 ( .A(n984), .B(n983), .Z(n990) );
  XNOR U1268 ( .A(y[19]), .B(x[19]), .Z(n983) );
  XNOR U1269 ( .A(y[18]), .B(x[18]), .Z(n984) );
  XNOR U1270 ( .A(n987), .B(n988), .Z(n989) );
  XNOR U1271 ( .A(y[17]), .B(x[17]), .Z(n988) );
  XNOR U1272 ( .A(y[16]), .B(x[16]), .Z(n987) );
  XNOR U1273 ( .A(n1023), .B(n1022), .Z(n1013) );
  XNOR U1274 ( .A(n995), .B(n996), .Z(n1002) );
  XNOR U1275 ( .A(n999), .B(n1000), .Z(n996) );
  XNOR U1276 ( .A(y[15]), .B(x[15]), .Z(n1000) );
  XNOR U1277 ( .A(y[14]), .B(x[14]), .Z(n999) );
  XNOR U1278 ( .A(n997), .B(n998), .Z(n995) );
  XNOR U1279 ( .A(y[13]), .B(x[13]), .Z(n998) );
  XNOR U1280 ( .A(y[12]), .B(x[12]), .Z(n997) );
  XNOR U1281 ( .A(n1010), .B(n1011), .Z(n1003) );
  XNOR U1282 ( .A(n1005), .B(n1004), .Z(n1011) );
  XNOR U1283 ( .A(y[11]), .B(x[11]), .Z(n1004) );
  XNOR U1284 ( .A(y[10]), .B(x[10]), .Z(n1005) );
  XNOR U1285 ( .A(n1008), .B(n1009), .Z(n1010) );
  XNOR U1286 ( .A(y[9]), .B(x[9]), .Z(n1009) );
  XNOR U1287 ( .A(y[8]), .B(x[8]), .Z(n1008) );
  XNOR U1288 ( .A(n1016), .B(n1017), .Z(n1025) );
  XNOR U1289 ( .A(n1020), .B(n1021), .Z(n1017) );
  XNOR U1290 ( .A(y[7]), .B(x[7]), .Z(n1021) );
  XNOR U1291 ( .A(y[6]), .B(x[6]), .Z(n1020) );
  XNOR U1292 ( .A(n1018), .B(n1019), .Z(n1016) );
  XNOR U1293 ( .A(y[5]), .B(x[5]), .Z(n1019) );
  XNOR U1294 ( .A(y[4]), .B(x[4]), .Z(n1018) );
  XNOR U1295 ( .A(n1033), .B(n1034), .Z(n1026) );
  XNOR U1296 ( .A(n1028), .B(n1027), .Z(n1034) );
  XNOR U1297 ( .A(y[3]), .B(x[3]), .Z(n1027) );
  XNOR U1298 ( .A(y[2]), .B(x[2]), .Z(n1028) );
  XNOR U1299 ( .A(n1031), .B(n1032), .Z(n1033) );
  XNOR U1300 ( .A(y[1]), .B(x[1]), .Z(n1032) );
  XNOR U1301 ( .A(y[0]), .B(x[0]), .Z(n1031) );
endmodule

