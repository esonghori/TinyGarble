
module compare_N16384_CC512 ( clk, rst, x, y, g );
  input [31:0] x;
  input [31:0] y;
  input clk, rst;
  output g;
  wire   ci, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160;

  DFF ci_reg ( .D(g), .CLK(clk), .RST(rst), .I(1'b1), .Q(ci) );
  XOR U36 ( .A(y[3]), .B(n147), .Z(n148) );
  XOR U37 ( .A(y[7]), .B(n131), .Z(n132) );
  XOR U38 ( .A(y[11]), .B(n115), .Z(n116) );
  XOR U39 ( .A(y[15]), .B(n99), .Z(n100) );
  XOR U40 ( .A(y[19]), .B(n83), .Z(n84) );
  XOR U41 ( .A(y[23]), .B(n67), .Z(n68) );
  XOR U42 ( .A(y[27]), .B(n51), .Z(n52) );
  XOR U43 ( .A(y[4]), .B(n143), .Z(n144) );
  XOR U44 ( .A(y[8]), .B(n127), .Z(n128) );
  XOR U45 ( .A(y[12]), .B(n111), .Z(n112) );
  XOR U46 ( .A(y[16]), .B(n95), .Z(n96) );
  XOR U47 ( .A(y[20]), .B(n79), .Z(n80) );
  XOR U48 ( .A(y[24]), .B(n63), .Z(n64) );
  XOR U49 ( .A(y[28]), .B(n47), .Z(n48) );
  XOR U50 ( .A(y[5]), .B(n139), .Z(n140) );
  XOR U51 ( .A(y[9]), .B(n123), .Z(n124) );
  XOR U52 ( .A(y[13]), .B(n107), .Z(n108) );
  XOR U53 ( .A(y[17]), .B(n91), .Z(n92) );
  XOR U54 ( .A(y[21]), .B(n75), .Z(n76) );
  XOR U55 ( .A(y[25]), .B(n59), .Z(n60) );
  XOR U56 ( .A(y[29]), .B(n43), .Z(n44) );
  XOR U57 ( .A(y[2]), .B(n151), .Z(n152) );
  XOR U58 ( .A(y[6]), .B(n135), .Z(n136) );
  XOR U59 ( .A(y[10]), .B(n119), .Z(n120) );
  XOR U60 ( .A(y[14]), .B(n103), .Z(n104) );
  XOR U61 ( .A(y[18]), .B(n87), .Z(n88) );
  XOR U62 ( .A(y[22]), .B(n71), .Z(n72) );
  XOR U63 ( .A(y[26]), .B(n55), .Z(n56) );
  XOR U64 ( .A(y[30]), .B(n39), .Z(n40) );
  XOR U65 ( .A(n34), .B(n35), .Z(g) );
  AND U66 ( .A(n36), .B(n37), .Z(n34) );
  XOR U67 ( .A(x[31]), .B(n35), .Z(n37) );
  XNOR U68 ( .A(y[31]), .B(n35), .Z(n36) );
  XNOR U69 ( .A(n38), .B(n39), .Z(n35) );
  AND U70 ( .A(n40), .B(n41), .Z(n38) );
  XNOR U71 ( .A(x[30]), .B(n39), .Z(n41) );
  XOR U72 ( .A(n42), .B(n43), .Z(n39) );
  AND U73 ( .A(n44), .B(n45), .Z(n42) );
  XNOR U74 ( .A(x[29]), .B(n43), .Z(n45) );
  XOR U75 ( .A(n46), .B(n47), .Z(n43) );
  AND U76 ( .A(n48), .B(n49), .Z(n46) );
  XNOR U77 ( .A(x[28]), .B(n47), .Z(n49) );
  XOR U78 ( .A(n50), .B(n51), .Z(n47) );
  AND U79 ( .A(n52), .B(n53), .Z(n50) );
  XNOR U80 ( .A(x[27]), .B(n51), .Z(n53) );
  XOR U81 ( .A(n54), .B(n55), .Z(n51) );
  AND U82 ( .A(n56), .B(n57), .Z(n54) );
  XNOR U83 ( .A(x[26]), .B(n55), .Z(n57) );
  XOR U84 ( .A(n58), .B(n59), .Z(n55) );
  AND U85 ( .A(n60), .B(n61), .Z(n58) );
  XNOR U86 ( .A(x[25]), .B(n59), .Z(n61) );
  XOR U87 ( .A(n62), .B(n63), .Z(n59) );
  AND U88 ( .A(n64), .B(n65), .Z(n62) );
  XNOR U89 ( .A(x[24]), .B(n63), .Z(n65) );
  XOR U90 ( .A(n66), .B(n67), .Z(n63) );
  AND U91 ( .A(n68), .B(n69), .Z(n66) );
  XNOR U92 ( .A(x[23]), .B(n67), .Z(n69) );
  XOR U93 ( .A(n70), .B(n71), .Z(n67) );
  AND U94 ( .A(n72), .B(n73), .Z(n70) );
  XNOR U95 ( .A(x[22]), .B(n71), .Z(n73) );
  XOR U96 ( .A(n74), .B(n75), .Z(n71) );
  AND U97 ( .A(n76), .B(n77), .Z(n74) );
  XNOR U98 ( .A(x[21]), .B(n75), .Z(n77) );
  XOR U99 ( .A(n78), .B(n79), .Z(n75) );
  AND U100 ( .A(n80), .B(n81), .Z(n78) );
  XNOR U101 ( .A(x[20]), .B(n79), .Z(n81) );
  XOR U102 ( .A(n82), .B(n83), .Z(n79) );
  AND U103 ( .A(n84), .B(n85), .Z(n82) );
  XNOR U104 ( .A(x[19]), .B(n83), .Z(n85) );
  XOR U105 ( .A(n86), .B(n87), .Z(n83) );
  AND U106 ( .A(n88), .B(n89), .Z(n86) );
  XNOR U107 ( .A(x[18]), .B(n87), .Z(n89) );
  XOR U108 ( .A(n90), .B(n91), .Z(n87) );
  AND U109 ( .A(n92), .B(n93), .Z(n90) );
  XNOR U110 ( .A(x[17]), .B(n91), .Z(n93) );
  XOR U111 ( .A(n94), .B(n95), .Z(n91) );
  AND U112 ( .A(n96), .B(n97), .Z(n94) );
  XNOR U113 ( .A(x[16]), .B(n95), .Z(n97) );
  XOR U114 ( .A(n98), .B(n99), .Z(n95) );
  AND U115 ( .A(n100), .B(n101), .Z(n98) );
  XNOR U116 ( .A(x[15]), .B(n99), .Z(n101) );
  XOR U117 ( .A(n102), .B(n103), .Z(n99) );
  AND U118 ( .A(n104), .B(n105), .Z(n102) );
  XNOR U119 ( .A(x[14]), .B(n103), .Z(n105) );
  XOR U120 ( .A(n106), .B(n107), .Z(n103) );
  AND U121 ( .A(n108), .B(n109), .Z(n106) );
  XNOR U122 ( .A(x[13]), .B(n107), .Z(n109) );
  XOR U123 ( .A(n110), .B(n111), .Z(n107) );
  AND U124 ( .A(n112), .B(n113), .Z(n110) );
  XNOR U125 ( .A(x[12]), .B(n111), .Z(n113) );
  XOR U126 ( .A(n114), .B(n115), .Z(n111) );
  AND U127 ( .A(n116), .B(n117), .Z(n114) );
  XNOR U128 ( .A(x[11]), .B(n115), .Z(n117) );
  XOR U129 ( .A(n118), .B(n119), .Z(n115) );
  AND U130 ( .A(n120), .B(n121), .Z(n118) );
  XNOR U131 ( .A(x[10]), .B(n119), .Z(n121) );
  XOR U132 ( .A(n122), .B(n123), .Z(n119) );
  AND U133 ( .A(n124), .B(n125), .Z(n122) );
  XNOR U134 ( .A(x[9]), .B(n123), .Z(n125) );
  XOR U135 ( .A(n126), .B(n127), .Z(n123) );
  AND U136 ( .A(n128), .B(n129), .Z(n126) );
  XNOR U137 ( .A(x[8]), .B(n127), .Z(n129) );
  XOR U138 ( .A(n130), .B(n131), .Z(n127) );
  AND U139 ( .A(n132), .B(n133), .Z(n130) );
  XNOR U140 ( .A(x[7]), .B(n131), .Z(n133) );
  XOR U141 ( .A(n134), .B(n135), .Z(n131) );
  AND U142 ( .A(n136), .B(n137), .Z(n134) );
  XNOR U143 ( .A(x[6]), .B(n135), .Z(n137) );
  XOR U144 ( .A(n138), .B(n139), .Z(n135) );
  AND U145 ( .A(n140), .B(n141), .Z(n138) );
  XNOR U146 ( .A(x[5]), .B(n139), .Z(n141) );
  XOR U147 ( .A(n142), .B(n143), .Z(n139) );
  AND U148 ( .A(n144), .B(n145), .Z(n142) );
  XNOR U149 ( .A(x[4]), .B(n143), .Z(n145) );
  XOR U150 ( .A(n146), .B(n147), .Z(n143) );
  AND U151 ( .A(n148), .B(n149), .Z(n146) );
  XNOR U152 ( .A(x[3]), .B(n147), .Z(n149) );
  XOR U153 ( .A(n150), .B(n151), .Z(n147) );
  AND U154 ( .A(n152), .B(n153), .Z(n150) );
  XNOR U155 ( .A(x[2]), .B(n151), .Z(n153) );
  XOR U156 ( .A(n154), .B(n155), .Z(n151) );
  AND U157 ( .A(n156), .B(n157), .Z(n154) );
  XNOR U158 ( .A(x[1]), .B(n155), .Z(n157) );
  XOR U159 ( .A(y[1]), .B(n155), .Z(n156) );
  XOR U160 ( .A(ci), .B(n158), .Z(n155) );
  NANDN U161 ( .A(n159), .B(n160), .Z(n158) );
  XOR U162 ( .A(x[0]), .B(ci), .Z(n160) );
  XOR U163 ( .A(y[0]), .B(ci), .Z(n159) );
endmodule

