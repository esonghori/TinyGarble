
module sum_N1024_CC4 ( clk, rst, a, b, c );
  input [255:0] a;
  input [255:0] b;
  output [255:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .Q(carry_on) );
  XOR U3 ( .A(a[0]), .B(b[0]), .Z(n1) );
  XOR U4 ( .A(n1), .B(carry_on), .Z(c[0]) );
  XOR U5 ( .A(a[1]), .B(b[1]), .Z(n4) );
  NAND U6 ( .A(b[0]), .B(a[0]), .Z(n3) );
  NAND U7 ( .A(carry_on), .B(n1), .Z(n2) );
  AND U8 ( .A(n3), .B(n2), .Z(n5) );
  XNOR U9 ( .A(n4), .B(n5), .Z(c[1]) );
  XOR U10 ( .A(a[2]), .B(b[2]), .Z(n8) );
  NAND U11 ( .A(b[1]), .B(a[1]), .Z(n7) );
  NANDN U12 ( .A(n5), .B(n4), .Z(n6) );
  AND U13 ( .A(n7), .B(n6), .Z(n9) );
  XNOR U14 ( .A(n8), .B(n9), .Z(c[2]) );
  XOR U15 ( .A(a[3]), .B(b[3]), .Z(n12) );
  NAND U16 ( .A(b[2]), .B(a[2]), .Z(n11) );
  NANDN U17 ( .A(n9), .B(n8), .Z(n10) );
  AND U18 ( .A(n11), .B(n10), .Z(n13) );
  XNOR U19 ( .A(n12), .B(n13), .Z(c[3]) );
  XOR U20 ( .A(a[4]), .B(b[4]), .Z(n16) );
  NAND U21 ( .A(b[3]), .B(a[3]), .Z(n15) );
  NANDN U22 ( .A(n13), .B(n12), .Z(n14) );
  AND U23 ( .A(n15), .B(n14), .Z(n17) );
  XNOR U24 ( .A(n16), .B(n17), .Z(c[4]) );
  XOR U25 ( .A(a[5]), .B(b[5]), .Z(n20) );
  NAND U26 ( .A(b[4]), .B(a[4]), .Z(n19) );
  NANDN U27 ( .A(n17), .B(n16), .Z(n18) );
  AND U28 ( .A(n19), .B(n18), .Z(n21) );
  XNOR U29 ( .A(n20), .B(n21), .Z(c[5]) );
  XOR U30 ( .A(a[6]), .B(b[6]), .Z(n24) );
  NAND U31 ( .A(b[5]), .B(a[5]), .Z(n23) );
  NANDN U32 ( .A(n21), .B(n20), .Z(n22) );
  AND U33 ( .A(n23), .B(n22), .Z(n25) );
  XNOR U34 ( .A(n24), .B(n25), .Z(c[6]) );
  XOR U35 ( .A(a[7]), .B(b[7]), .Z(n28) );
  NAND U36 ( .A(b[6]), .B(a[6]), .Z(n27) );
  NANDN U37 ( .A(n25), .B(n24), .Z(n26) );
  AND U38 ( .A(n27), .B(n26), .Z(n29) );
  XNOR U39 ( .A(n28), .B(n29), .Z(c[7]) );
  XOR U40 ( .A(a[8]), .B(b[8]), .Z(n32) );
  NAND U41 ( .A(b[7]), .B(a[7]), .Z(n31) );
  NANDN U42 ( .A(n29), .B(n28), .Z(n30) );
  AND U43 ( .A(n31), .B(n30), .Z(n33) );
  XNOR U44 ( .A(n32), .B(n33), .Z(c[8]) );
  XOR U45 ( .A(a[9]), .B(b[9]), .Z(n36) );
  NAND U46 ( .A(b[8]), .B(a[8]), .Z(n35) );
  NANDN U47 ( .A(n33), .B(n32), .Z(n34) );
  AND U48 ( .A(n35), .B(n34), .Z(n37) );
  XNOR U49 ( .A(n36), .B(n37), .Z(c[9]) );
  XOR U50 ( .A(a[10]), .B(b[10]), .Z(n40) );
  NAND U51 ( .A(b[9]), .B(a[9]), .Z(n39) );
  NANDN U52 ( .A(n37), .B(n36), .Z(n38) );
  AND U53 ( .A(n39), .B(n38), .Z(n41) );
  XNOR U54 ( .A(n40), .B(n41), .Z(c[10]) );
  XOR U55 ( .A(a[11]), .B(b[11]), .Z(n44) );
  NAND U56 ( .A(b[10]), .B(a[10]), .Z(n43) );
  NANDN U57 ( .A(n41), .B(n40), .Z(n42) );
  AND U58 ( .A(n43), .B(n42), .Z(n45) );
  XNOR U59 ( .A(n44), .B(n45), .Z(c[11]) );
  XOR U60 ( .A(a[12]), .B(b[12]), .Z(n48) );
  NAND U61 ( .A(b[11]), .B(a[11]), .Z(n47) );
  NANDN U62 ( .A(n45), .B(n44), .Z(n46) );
  AND U63 ( .A(n47), .B(n46), .Z(n49) );
  XNOR U64 ( .A(n48), .B(n49), .Z(c[12]) );
  XOR U65 ( .A(a[13]), .B(b[13]), .Z(n52) );
  NAND U66 ( .A(b[12]), .B(a[12]), .Z(n51) );
  NANDN U67 ( .A(n49), .B(n48), .Z(n50) );
  AND U68 ( .A(n51), .B(n50), .Z(n53) );
  XNOR U69 ( .A(n52), .B(n53), .Z(c[13]) );
  XOR U70 ( .A(a[14]), .B(b[14]), .Z(n56) );
  NAND U71 ( .A(b[13]), .B(a[13]), .Z(n55) );
  NANDN U72 ( .A(n53), .B(n52), .Z(n54) );
  AND U73 ( .A(n55), .B(n54), .Z(n57) );
  XNOR U74 ( .A(n56), .B(n57), .Z(c[14]) );
  XOR U75 ( .A(a[15]), .B(b[15]), .Z(n60) );
  NAND U76 ( .A(b[14]), .B(a[14]), .Z(n59) );
  NANDN U77 ( .A(n57), .B(n56), .Z(n58) );
  AND U78 ( .A(n59), .B(n58), .Z(n61) );
  XNOR U79 ( .A(n60), .B(n61), .Z(c[15]) );
  XOR U80 ( .A(a[16]), .B(b[16]), .Z(n64) );
  NAND U81 ( .A(b[15]), .B(a[15]), .Z(n63) );
  NANDN U82 ( .A(n61), .B(n60), .Z(n62) );
  AND U83 ( .A(n63), .B(n62), .Z(n65) );
  XNOR U84 ( .A(n64), .B(n65), .Z(c[16]) );
  XOR U85 ( .A(a[17]), .B(b[17]), .Z(n68) );
  NAND U86 ( .A(b[16]), .B(a[16]), .Z(n67) );
  NANDN U87 ( .A(n65), .B(n64), .Z(n66) );
  AND U88 ( .A(n67), .B(n66), .Z(n69) );
  XNOR U89 ( .A(n68), .B(n69), .Z(c[17]) );
  XOR U90 ( .A(a[18]), .B(b[18]), .Z(n72) );
  NAND U91 ( .A(b[17]), .B(a[17]), .Z(n71) );
  NANDN U92 ( .A(n69), .B(n68), .Z(n70) );
  AND U93 ( .A(n71), .B(n70), .Z(n73) );
  XNOR U94 ( .A(n72), .B(n73), .Z(c[18]) );
  XOR U95 ( .A(a[19]), .B(b[19]), .Z(n76) );
  NAND U96 ( .A(b[18]), .B(a[18]), .Z(n75) );
  NANDN U97 ( .A(n73), .B(n72), .Z(n74) );
  AND U98 ( .A(n75), .B(n74), .Z(n77) );
  XNOR U99 ( .A(n76), .B(n77), .Z(c[19]) );
  XOR U100 ( .A(a[20]), .B(b[20]), .Z(n80) );
  NAND U101 ( .A(b[19]), .B(a[19]), .Z(n79) );
  NANDN U102 ( .A(n77), .B(n76), .Z(n78) );
  AND U103 ( .A(n79), .B(n78), .Z(n81) );
  XNOR U104 ( .A(n80), .B(n81), .Z(c[20]) );
  XOR U105 ( .A(a[21]), .B(b[21]), .Z(n84) );
  NAND U106 ( .A(b[20]), .B(a[20]), .Z(n83) );
  NANDN U107 ( .A(n81), .B(n80), .Z(n82) );
  AND U108 ( .A(n83), .B(n82), .Z(n85) );
  XNOR U109 ( .A(n84), .B(n85), .Z(c[21]) );
  XOR U110 ( .A(a[22]), .B(b[22]), .Z(n88) );
  NAND U111 ( .A(b[21]), .B(a[21]), .Z(n87) );
  NANDN U112 ( .A(n85), .B(n84), .Z(n86) );
  AND U113 ( .A(n87), .B(n86), .Z(n89) );
  XNOR U114 ( .A(n88), .B(n89), .Z(c[22]) );
  XOR U115 ( .A(a[23]), .B(b[23]), .Z(n92) );
  NAND U116 ( .A(b[22]), .B(a[22]), .Z(n91) );
  NANDN U117 ( .A(n89), .B(n88), .Z(n90) );
  AND U118 ( .A(n91), .B(n90), .Z(n93) );
  XNOR U119 ( .A(n92), .B(n93), .Z(c[23]) );
  XOR U120 ( .A(a[24]), .B(b[24]), .Z(n96) );
  NAND U121 ( .A(b[23]), .B(a[23]), .Z(n95) );
  NANDN U122 ( .A(n93), .B(n92), .Z(n94) );
  AND U123 ( .A(n95), .B(n94), .Z(n97) );
  XNOR U124 ( .A(n96), .B(n97), .Z(c[24]) );
  XOR U125 ( .A(a[25]), .B(b[25]), .Z(n100) );
  NAND U126 ( .A(b[24]), .B(a[24]), .Z(n99) );
  NANDN U127 ( .A(n97), .B(n96), .Z(n98) );
  AND U128 ( .A(n99), .B(n98), .Z(n101) );
  XNOR U129 ( .A(n100), .B(n101), .Z(c[25]) );
  XOR U130 ( .A(a[26]), .B(b[26]), .Z(n104) );
  NAND U131 ( .A(b[25]), .B(a[25]), .Z(n103) );
  NANDN U132 ( .A(n101), .B(n100), .Z(n102) );
  AND U133 ( .A(n103), .B(n102), .Z(n105) );
  XNOR U134 ( .A(n104), .B(n105), .Z(c[26]) );
  XOR U135 ( .A(a[27]), .B(b[27]), .Z(n108) );
  NAND U136 ( .A(b[26]), .B(a[26]), .Z(n107) );
  NANDN U137 ( .A(n105), .B(n104), .Z(n106) );
  AND U138 ( .A(n107), .B(n106), .Z(n109) );
  XNOR U139 ( .A(n108), .B(n109), .Z(c[27]) );
  XOR U140 ( .A(a[28]), .B(b[28]), .Z(n112) );
  NAND U141 ( .A(b[27]), .B(a[27]), .Z(n111) );
  NANDN U142 ( .A(n109), .B(n108), .Z(n110) );
  AND U143 ( .A(n111), .B(n110), .Z(n113) );
  XNOR U144 ( .A(n112), .B(n113), .Z(c[28]) );
  XOR U145 ( .A(a[29]), .B(b[29]), .Z(n116) );
  NAND U146 ( .A(b[28]), .B(a[28]), .Z(n115) );
  NANDN U147 ( .A(n113), .B(n112), .Z(n114) );
  AND U148 ( .A(n115), .B(n114), .Z(n117) );
  XNOR U149 ( .A(n116), .B(n117), .Z(c[29]) );
  XOR U150 ( .A(a[30]), .B(b[30]), .Z(n120) );
  NAND U151 ( .A(b[29]), .B(a[29]), .Z(n119) );
  NANDN U152 ( .A(n117), .B(n116), .Z(n118) );
  AND U153 ( .A(n119), .B(n118), .Z(n121) );
  XNOR U154 ( .A(n120), .B(n121), .Z(c[30]) );
  XOR U155 ( .A(a[31]), .B(b[31]), .Z(n124) );
  NAND U156 ( .A(b[30]), .B(a[30]), .Z(n123) );
  NANDN U157 ( .A(n121), .B(n120), .Z(n122) );
  AND U158 ( .A(n123), .B(n122), .Z(n125) );
  XNOR U159 ( .A(n124), .B(n125), .Z(c[31]) );
  XOR U160 ( .A(a[32]), .B(b[32]), .Z(n128) );
  NAND U161 ( .A(b[31]), .B(a[31]), .Z(n127) );
  NANDN U162 ( .A(n125), .B(n124), .Z(n126) );
  AND U163 ( .A(n127), .B(n126), .Z(n129) );
  XNOR U164 ( .A(n128), .B(n129), .Z(c[32]) );
  XOR U165 ( .A(a[33]), .B(b[33]), .Z(n132) );
  NAND U166 ( .A(b[32]), .B(a[32]), .Z(n131) );
  NANDN U167 ( .A(n129), .B(n128), .Z(n130) );
  AND U168 ( .A(n131), .B(n130), .Z(n133) );
  XNOR U169 ( .A(n132), .B(n133), .Z(c[33]) );
  XOR U170 ( .A(a[34]), .B(b[34]), .Z(n136) );
  NAND U171 ( .A(b[33]), .B(a[33]), .Z(n135) );
  NANDN U172 ( .A(n133), .B(n132), .Z(n134) );
  AND U173 ( .A(n135), .B(n134), .Z(n137) );
  XNOR U174 ( .A(n136), .B(n137), .Z(c[34]) );
  XOR U175 ( .A(a[35]), .B(b[35]), .Z(n140) );
  NAND U176 ( .A(b[34]), .B(a[34]), .Z(n139) );
  NANDN U177 ( .A(n137), .B(n136), .Z(n138) );
  AND U178 ( .A(n139), .B(n138), .Z(n141) );
  XNOR U179 ( .A(n140), .B(n141), .Z(c[35]) );
  XOR U180 ( .A(a[36]), .B(b[36]), .Z(n144) );
  NAND U181 ( .A(b[35]), .B(a[35]), .Z(n143) );
  NANDN U182 ( .A(n141), .B(n140), .Z(n142) );
  AND U183 ( .A(n143), .B(n142), .Z(n145) );
  XNOR U184 ( .A(n144), .B(n145), .Z(c[36]) );
  XOR U185 ( .A(a[37]), .B(b[37]), .Z(n148) );
  NAND U186 ( .A(b[36]), .B(a[36]), .Z(n147) );
  NANDN U187 ( .A(n145), .B(n144), .Z(n146) );
  AND U188 ( .A(n147), .B(n146), .Z(n149) );
  XNOR U189 ( .A(n148), .B(n149), .Z(c[37]) );
  XOR U190 ( .A(a[38]), .B(b[38]), .Z(n152) );
  NAND U191 ( .A(b[37]), .B(a[37]), .Z(n151) );
  NANDN U192 ( .A(n149), .B(n148), .Z(n150) );
  AND U193 ( .A(n151), .B(n150), .Z(n153) );
  XNOR U194 ( .A(n152), .B(n153), .Z(c[38]) );
  XOR U195 ( .A(a[39]), .B(b[39]), .Z(n156) );
  NAND U196 ( .A(b[38]), .B(a[38]), .Z(n155) );
  NANDN U197 ( .A(n153), .B(n152), .Z(n154) );
  AND U198 ( .A(n155), .B(n154), .Z(n157) );
  XNOR U199 ( .A(n156), .B(n157), .Z(c[39]) );
  XOR U200 ( .A(a[40]), .B(b[40]), .Z(n160) );
  NAND U201 ( .A(b[39]), .B(a[39]), .Z(n159) );
  NANDN U202 ( .A(n157), .B(n156), .Z(n158) );
  AND U203 ( .A(n159), .B(n158), .Z(n161) );
  XNOR U204 ( .A(n160), .B(n161), .Z(c[40]) );
  XOR U205 ( .A(a[41]), .B(b[41]), .Z(n164) );
  NAND U206 ( .A(b[40]), .B(a[40]), .Z(n163) );
  NANDN U207 ( .A(n161), .B(n160), .Z(n162) );
  AND U208 ( .A(n163), .B(n162), .Z(n165) );
  XNOR U209 ( .A(n164), .B(n165), .Z(c[41]) );
  XOR U210 ( .A(a[42]), .B(b[42]), .Z(n168) );
  NAND U211 ( .A(b[41]), .B(a[41]), .Z(n167) );
  NANDN U212 ( .A(n165), .B(n164), .Z(n166) );
  AND U213 ( .A(n167), .B(n166), .Z(n169) );
  XNOR U214 ( .A(n168), .B(n169), .Z(c[42]) );
  XOR U215 ( .A(a[43]), .B(b[43]), .Z(n172) );
  NAND U216 ( .A(b[42]), .B(a[42]), .Z(n171) );
  NANDN U217 ( .A(n169), .B(n168), .Z(n170) );
  AND U218 ( .A(n171), .B(n170), .Z(n173) );
  XNOR U219 ( .A(n172), .B(n173), .Z(c[43]) );
  XOR U220 ( .A(a[44]), .B(b[44]), .Z(n176) );
  NAND U221 ( .A(b[43]), .B(a[43]), .Z(n175) );
  NANDN U222 ( .A(n173), .B(n172), .Z(n174) );
  AND U223 ( .A(n175), .B(n174), .Z(n177) );
  XNOR U224 ( .A(n176), .B(n177), .Z(c[44]) );
  XOR U225 ( .A(a[45]), .B(b[45]), .Z(n180) );
  NAND U226 ( .A(b[44]), .B(a[44]), .Z(n179) );
  NANDN U227 ( .A(n177), .B(n176), .Z(n178) );
  AND U228 ( .A(n179), .B(n178), .Z(n181) );
  XNOR U229 ( .A(n180), .B(n181), .Z(c[45]) );
  XOR U230 ( .A(a[46]), .B(b[46]), .Z(n184) );
  NAND U231 ( .A(b[45]), .B(a[45]), .Z(n183) );
  NANDN U232 ( .A(n181), .B(n180), .Z(n182) );
  AND U233 ( .A(n183), .B(n182), .Z(n185) );
  XNOR U234 ( .A(n184), .B(n185), .Z(c[46]) );
  XOR U235 ( .A(a[47]), .B(b[47]), .Z(n188) );
  NAND U236 ( .A(b[46]), .B(a[46]), .Z(n187) );
  NANDN U237 ( .A(n185), .B(n184), .Z(n186) );
  AND U238 ( .A(n187), .B(n186), .Z(n189) );
  XNOR U239 ( .A(n188), .B(n189), .Z(c[47]) );
  XOR U240 ( .A(a[48]), .B(b[48]), .Z(n192) );
  NAND U241 ( .A(b[47]), .B(a[47]), .Z(n191) );
  NANDN U242 ( .A(n189), .B(n188), .Z(n190) );
  AND U243 ( .A(n191), .B(n190), .Z(n193) );
  XNOR U244 ( .A(n192), .B(n193), .Z(c[48]) );
  XOR U245 ( .A(a[49]), .B(b[49]), .Z(n196) );
  NAND U246 ( .A(b[48]), .B(a[48]), .Z(n195) );
  NANDN U247 ( .A(n193), .B(n192), .Z(n194) );
  AND U248 ( .A(n195), .B(n194), .Z(n197) );
  XNOR U249 ( .A(n196), .B(n197), .Z(c[49]) );
  XOR U250 ( .A(a[50]), .B(b[50]), .Z(n200) );
  NAND U251 ( .A(b[49]), .B(a[49]), .Z(n199) );
  NANDN U252 ( .A(n197), .B(n196), .Z(n198) );
  AND U253 ( .A(n199), .B(n198), .Z(n201) );
  XNOR U254 ( .A(n200), .B(n201), .Z(c[50]) );
  XOR U255 ( .A(a[51]), .B(b[51]), .Z(n204) );
  NAND U256 ( .A(b[50]), .B(a[50]), .Z(n203) );
  NANDN U257 ( .A(n201), .B(n200), .Z(n202) );
  AND U258 ( .A(n203), .B(n202), .Z(n205) );
  XNOR U259 ( .A(n204), .B(n205), .Z(c[51]) );
  XOR U260 ( .A(a[52]), .B(b[52]), .Z(n208) );
  NAND U261 ( .A(b[51]), .B(a[51]), .Z(n207) );
  NANDN U262 ( .A(n205), .B(n204), .Z(n206) );
  AND U263 ( .A(n207), .B(n206), .Z(n209) );
  XNOR U264 ( .A(n208), .B(n209), .Z(c[52]) );
  XOR U265 ( .A(a[53]), .B(b[53]), .Z(n212) );
  NAND U266 ( .A(b[52]), .B(a[52]), .Z(n211) );
  NANDN U267 ( .A(n209), .B(n208), .Z(n210) );
  AND U268 ( .A(n211), .B(n210), .Z(n213) );
  XNOR U269 ( .A(n212), .B(n213), .Z(c[53]) );
  XOR U270 ( .A(a[54]), .B(b[54]), .Z(n216) );
  NAND U271 ( .A(b[53]), .B(a[53]), .Z(n215) );
  NANDN U272 ( .A(n213), .B(n212), .Z(n214) );
  AND U273 ( .A(n215), .B(n214), .Z(n217) );
  XNOR U274 ( .A(n216), .B(n217), .Z(c[54]) );
  XOR U275 ( .A(a[55]), .B(b[55]), .Z(n220) );
  NAND U276 ( .A(b[54]), .B(a[54]), .Z(n219) );
  NANDN U277 ( .A(n217), .B(n216), .Z(n218) );
  AND U278 ( .A(n219), .B(n218), .Z(n221) );
  XNOR U279 ( .A(n220), .B(n221), .Z(c[55]) );
  XOR U280 ( .A(a[56]), .B(b[56]), .Z(n224) );
  NAND U281 ( .A(b[55]), .B(a[55]), .Z(n223) );
  NANDN U282 ( .A(n221), .B(n220), .Z(n222) );
  AND U283 ( .A(n223), .B(n222), .Z(n225) );
  XNOR U284 ( .A(n224), .B(n225), .Z(c[56]) );
  XOR U285 ( .A(a[57]), .B(b[57]), .Z(n228) );
  NAND U286 ( .A(b[56]), .B(a[56]), .Z(n227) );
  NANDN U287 ( .A(n225), .B(n224), .Z(n226) );
  AND U288 ( .A(n227), .B(n226), .Z(n229) );
  XNOR U289 ( .A(n228), .B(n229), .Z(c[57]) );
  XOR U290 ( .A(a[58]), .B(b[58]), .Z(n232) );
  NAND U291 ( .A(b[57]), .B(a[57]), .Z(n231) );
  NANDN U292 ( .A(n229), .B(n228), .Z(n230) );
  AND U293 ( .A(n231), .B(n230), .Z(n233) );
  XNOR U294 ( .A(n232), .B(n233), .Z(c[58]) );
  XOR U295 ( .A(a[59]), .B(b[59]), .Z(n236) );
  NAND U296 ( .A(b[58]), .B(a[58]), .Z(n235) );
  NANDN U297 ( .A(n233), .B(n232), .Z(n234) );
  AND U298 ( .A(n235), .B(n234), .Z(n237) );
  XNOR U299 ( .A(n236), .B(n237), .Z(c[59]) );
  XOR U300 ( .A(a[60]), .B(b[60]), .Z(n240) );
  NAND U301 ( .A(b[59]), .B(a[59]), .Z(n239) );
  NANDN U302 ( .A(n237), .B(n236), .Z(n238) );
  AND U303 ( .A(n239), .B(n238), .Z(n241) );
  XNOR U304 ( .A(n240), .B(n241), .Z(c[60]) );
  XOR U305 ( .A(a[61]), .B(b[61]), .Z(n244) );
  NAND U306 ( .A(b[60]), .B(a[60]), .Z(n243) );
  NANDN U307 ( .A(n241), .B(n240), .Z(n242) );
  AND U308 ( .A(n243), .B(n242), .Z(n245) );
  XNOR U309 ( .A(n244), .B(n245), .Z(c[61]) );
  XOR U310 ( .A(a[62]), .B(b[62]), .Z(n248) );
  NAND U311 ( .A(b[61]), .B(a[61]), .Z(n247) );
  NANDN U312 ( .A(n245), .B(n244), .Z(n246) );
  AND U313 ( .A(n247), .B(n246), .Z(n249) );
  XNOR U314 ( .A(n248), .B(n249), .Z(c[62]) );
  XOR U315 ( .A(a[63]), .B(b[63]), .Z(n252) );
  NAND U316 ( .A(b[62]), .B(a[62]), .Z(n251) );
  NANDN U317 ( .A(n249), .B(n248), .Z(n250) );
  AND U318 ( .A(n251), .B(n250), .Z(n253) );
  XNOR U319 ( .A(n252), .B(n253), .Z(c[63]) );
  XOR U320 ( .A(a[64]), .B(b[64]), .Z(n256) );
  NAND U321 ( .A(b[63]), .B(a[63]), .Z(n255) );
  NANDN U322 ( .A(n253), .B(n252), .Z(n254) );
  AND U323 ( .A(n255), .B(n254), .Z(n257) );
  XNOR U324 ( .A(n256), .B(n257), .Z(c[64]) );
  XOR U325 ( .A(a[65]), .B(b[65]), .Z(n260) );
  NAND U326 ( .A(b[64]), .B(a[64]), .Z(n259) );
  NANDN U327 ( .A(n257), .B(n256), .Z(n258) );
  AND U328 ( .A(n259), .B(n258), .Z(n261) );
  XNOR U329 ( .A(n260), .B(n261), .Z(c[65]) );
  XOR U330 ( .A(a[66]), .B(b[66]), .Z(n264) );
  NAND U331 ( .A(b[65]), .B(a[65]), .Z(n263) );
  NANDN U332 ( .A(n261), .B(n260), .Z(n262) );
  AND U333 ( .A(n263), .B(n262), .Z(n265) );
  XNOR U334 ( .A(n264), .B(n265), .Z(c[66]) );
  XOR U335 ( .A(a[67]), .B(b[67]), .Z(n268) );
  NAND U336 ( .A(b[66]), .B(a[66]), .Z(n267) );
  NANDN U337 ( .A(n265), .B(n264), .Z(n266) );
  AND U338 ( .A(n267), .B(n266), .Z(n269) );
  XNOR U339 ( .A(n268), .B(n269), .Z(c[67]) );
  XOR U340 ( .A(a[68]), .B(b[68]), .Z(n272) );
  NAND U341 ( .A(b[67]), .B(a[67]), .Z(n271) );
  NANDN U342 ( .A(n269), .B(n268), .Z(n270) );
  AND U343 ( .A(n271), .B(n270), .Z(n273) );
  XNOR U344 ( .A(n272), .B(n273), .Z(c[68]) );
  XOR U345 ( .A(a[69]), .B(b[69]), .Z(n276) );
  NAND U346 ( .A(b[68]), .B(a[68]), .Z(n275) );
  NANDN U347 ( .A(n273), .B(n272), .Z(n274) );
  AND U348 ( .A(n275), .B(n274), .Z(n277) );
  XNOR U349 ( .A(n276), .B(n277), .Z(c[69]) );
  XOR U350 ( .A(a[70]), .B(b[70]), .Z(n280) );
  NAND U351 ( .A(b[69]), .B(a[69]), .Z(n279) );
  NANDN U352 ( .A(n277), .B(n276), .Z(n278) );
  AND U353 ( .A(n279), .B(n278), .Z(n281) );
  XNOR U354 ( .A(n280), .B(n281), .Z(c[70]) );
  XOR U355 ( .A(a[71]), .B(b[71]), .Z(n284) );
  NAND U356 ( .A(b[70]), .B(a[70]), .Z(n283) );
  NANDN U357 ( .A(n281), .B(n280), .Z(n282) );
  AND U358 ( .A(n283), .B(n282), .Z(n285) );
  XNOR U359 ( .A(n284), .B(n285), .Z(c[71]) );
  XOR U360 ( .A(a[72]), .B(b[72]), .Z(n288) );
  NAND U361 ( .A(b[71]), .B(a[71]), .Z(n287) );
  NANDN U362 ( .A(n285), .B(n284), .Z(n286) );
  AND U363 ( .A(n287), .B(n286), .Z(n289) );
  XNOR U364 ( .A(n288), .B(n289), .Z(c[72]) );
  XOR U365 ( .A(a[73]), .B(b[73]), .Z(n292) );
  NAND U366 ( .A(b[72]), .B(a[72]), .Z(n291) );
  NANDN U367 ( .A(n289), .B(n288), .Z(n290) );
  AND U368 ( .A(n291), .B(n290), .Z(n293) );
  XNOR U369 ( .A(n292), .B(n293), .Z(c[73]) );
  XOR U370 ( .A(a[74]), .B(b[74]), .Z(n296) );
  NAND U371 ( .A(b[73]), .B(a[73]), .Z(n295) );
  NANDN U372 ( .A(n293), .B(n292), .Z(n294) );
  AND U373 ( .A(n295), .B(n294), .Z(n297) );
  XNOR U374 ( .A(n296), .B(n297), .Z(c[74]) );
  XOR U375 ( .A(a[75]), .B(b[75]), .Z(n300) );
  NAND U376 ( .A(b[74]), .B(a[74]), .Z(n299) );
  NANDN U377 ( .A(n297), .B(n296), .Z(n298) );
  AND U378 ( .A(n299), .B(n298), .Z(n301) );
  XNOR U379 ( .A(n300), .B(n301), .Z(c[75]) );
  XOR U380 ( .A(a[76]), .B(b[76]), .Z(n304) );
  NAND U381 ( .A(b[75]), .B(a[75]), .Z(n303) );
  NANDN U382 ( .A(n301), .B(n300), .Z(n302) );
  AND U383 ( .A(n303), .B(n302), .Z(n305) );
  XNOR U384 ( .A(n304), .B(n305), .Z(c[76]) );
  XOR U385 ( .A(a[77]), .B(b[77]), .Z(n308) );
  NAND U386 ( .A(b[76]), .B(a[76]), .Z(n307) );
  NANDN U387 ( .A(n305), .B(n304), .Z(n306) );
  AND U388 ( .A(n307), .B(n306), .Z(n309) );
  XNOR U389 ( .A(n308), .B(n309), .Z(c[77]) );
  XOR U390 ( .A(a[78]), .B(b[78]), .Z(n312) );
  NAND U391 ( .A(b[77]), .B(a[77]), .Z(n311) );
  NANDN U392 ( .A(n309), .B(n308), .Z(n310) );
  AND U393 ( .A(n311), .B(n310), .Z(n313) );
  XNOR U394 ( .A(n312), .B(n313), .Z(c[78]) );
  XOR U395 ( .A(a[79]), .B(b[79]), .Z(n316) );
  NAND U396 ( .A(b[78]), .B(a[78]), .Z(n315) );
  NANDN U397 ( .A(n313), .B(n312), .Z(n314) );
  AND U398 ( .A(n315), .B(n314), .Z(n317) );
  XNOR U399 ( .A(n316), .B(n317), .Z(c[79]) );
  XOR U400 ( .A(a[80]), .B(b[80]), .Z(n320) );
  NAND U401 ( .A(b[79]), .B(a[79]), .Z(n319) );
  NANDN U402 ( .A(n317), .B(n316), .Z(n318) );
  AND U403 ( .A(n319), .B(n318), .Z(n321) );
  XNOR U404 ( .A(n320), .B(n321), .Z(c[80]) );
  XOR U405 ( .A(a[81]), .B(b[81]), .Z(n324) );
  NAND U406 ( .A(b[80]), .B(a[80]), .Z(n323) );
  NANDN U407 ( .A(n321), .B(n320), .Z(n322) );
  AND U408 ( .A(n323), .B(n322), .Z(n325) );
  XNOR U409 ( .A(n324), .B(n325), .Z(c[81]) );
  XOR U410 ( .A(a[82]), .B(b[82]), .Z(n328) );
  NAND U411 ( .A(b[81]), .B(a[81]), .Z(n327) );
  NANDN U412 ( .A(n325), .B(n324), .Z(n326) );
  AND U413 ( .A(n327), .B(n326), .Z(n329) );
  XNOR U414 ( .A(n328), .B(n329), .Z(c[82]) );
  XOR U415 ( .A(a[83]), .B(b[83]), .Z(n332) );
  NAND U416 ( .A(b[82]), .B(a[82]), .Z(n331) );
  NANDN U417 ( .A(n329), .B(n328), .Z(n330) );
  AND U418 ( .A(n331), .B(n330), .Z(n333) );
  XNOR U419 ( .A(n332), .B(n333), .Z(c[83]) );
  XOR U420 ( .A(a[84]), .B(b[84]), .Z(n336) );
  NAND U421 ( .A(b[83]), .B(a[83]), .Z(n335) );
  NANDN U422 ( .A(n333), .B(n332), .Z(n334) );
  AND U423 ( .A(n335), .B(n334), .Z(n337) );
  XNOR U424 ( .A(n336), .B(n337), .Z(c[84]) );
  XOR U425 ( .A(a[85]), .B(b[85]), .Z(n340) );
  NAND U426 ( .A(b[84]), .B(a[84]), .Z(n339) );
  NANDN U427 ( .A(n337), .B(n336), .Z(n338) );
  AND U428 ( .A(n339), .B(n338), .Z(n341) );
  XNOR U429 ( .A(n340), .B(n341), .Z(c[85]) );
  XOR U430 ( .A(a[86]), .B(b[86]), .Z(n344) );
  NAND U431 ( .A(b[85]), .B(a[85]), .Z(n343) );
  NANDN U432 ( .A(n341), .B(n340), .Z(n342) );
  AND U433 ( .A(n343), .B(n342), .Z(n345) );
  XNOR U434 ( .A(n344), .B(n345), .Z(c[86]) );
  XOR U435 ( .A(a[87]), .B(b[87]), .Z(n348) );
  NAND U436 ( .A(b[86]), .B(a[86]), .Z(n347) );
  NANDN U437 ( .A(n345), .B(n344), .Z(n346) );
  AND U438 ( .A(n347), .B(n346), .Z(n349) );
  XNOR U439 ( .A(n348), .B(n349), .Z(c[87]) );
  XOR U440 ( .A(a[88]), .B(b[88]), .Z(n352) );
  NAND U441 ( .A(b[87]), .B(a[87]), .Z(n351) );
  NANDN U442 ( .A(n349), .B(n348), .Z(n350) );
  AND U443 ( .A(n351), .B(n350), .Z(n353) );
  XNOR U444 ( .A(n352), .B(n353), .Z(c[88]) );
  XOR U445 ( .A(a[89]), .B(b[89]), .Z(n356) );
  NAND U446 ( .A(b[88]), .B(a[88]), .Z(n355) );
  NANDN U447 ( .A(n353), .B(n352), .Z(n354) );
  AND U448 ( .A(n355), .B(n354), .Z(n357) );
  XNOR U449 ( .A(n356), .B(n357), .Z(c[89]) );
  XOR U450 ( .A(a[90]), .B(b[90]), .Z(n360) );
  NAND U451 ( .A(b[89]), .B(a[89]), .Z(n359) );
  NANDN U452 ( .A(n357), .B(n356), .Z(n358) );
  AND U453 ( .A(n359), .B(n358), .Z(n361) );
  XNOR U454 ( .A(n360), .B(n361), .Z(c[90]) );
  XOR U455 ( .A(a[91]), .B(b[91]), .Z(n364) );
  NAND U456 ( .A(b[90]), .B(a[90]), .Z(n363) );
  NANDN U457 ( .A(n361), .B(n360), .Z(n362) );
  AND U458 ( .A(n363), .B(n362), .Z(n365) );
  XNOR U459 ( .A(n364), .B(n365), .Z(c[91]) );
  XOR U460 ( .A(a[92]), .B(b[92]), .Z(n368) );
  NAND U461 ( .A(b[91]), .B(a[91]), .Z(n367) );
  NANDN U462 ( .A(n365), .B(n364), .Z(n366) );
  AND U463 ( .A(n367), .B(n366), .Z(n369) );
  XNOR U464 ( .A(n368), .B(n369), .Z(c[92]) );
  XOR U465 ( .A(a[93]), .B(b[93]), .Z(n372) );
  NAND U466 ( .A(b[92]), .B(a[92]), .Z(n371) );
  NANDN U467 ( .A(n369), .B(n368), .Z(n370) );
  AND U468 ( .A(n371), .B(n370), .Z(n373) );
  XNOR U469 ( .A(n372), .B(n373), .Z(c[93]) );
  XOR U470 ( .A(a[94]), .B(b[94]), .Z(n376) );
  NAND U471 ( .A(b[93]), .B(a[93]), .Z(n375) );
  NANDN U472 ( .A(n373), .B(n372), .Z(n374) );
  AND U473 ( .A(n375), .B(n374), .Z(n377) );
  XNOR U474 ( .A(n376), .B(n377), .Z(c[94]) );
  XOR U475 ( .A(a[95]), .B(b[95]), .Z(n380) );
  NAND U476 ( .A(b[94]), .B(a[94]), .Z(n379) );
  NANDN U477 ( .A(n377), .B(n376), .Z(n378) );
  AND U478 ( .A(n379), .B(n378), .Z(n381) );
  XNOR U479 ( .A(n380), .B(n381), .Z(c[95]) );
  XOR U480 ( .A(a[96]), .B(b[96]), .Z(n384) );
  NAND U481 ( .A(b[95]), .B(a[95]), .Z(n383) );
  NANDN U482 ( .A(n381), .B(n380), .Z(n382) );
  AND U483 ( .A(n383), .B(n382), .Z(n385) );
  XNOR U484 ( .A(n384), .B(n385), .Z(c[96]) );
  XOR U485 ( .A(a[97]), .B(b[97]), .Z(n388) );
  NAND U486 ( .A(b[96]), .B(a[96]), .Z(n387) );
  NANDN U487 ( .A(n385), .B(n384), .Z(n386) );
  AND U488 ( .A(n387), .B(n386), .Z(n389) );
  XNOR U489 ( .A(n388), .B(n389), .Z(c[97]) );
  XOR U490 ( .A(a[98]), .B(b[98]), .Z(n392) );
  NAND U491 ( .A(b[97]), .B(a[97]), .Z(n391) );
  NANDN U492 ( .A(n389), .B(n388), .Z(n390) );
  AND U493 ( .A(n391), .B(n390), .Z(n393) );
  XNOR U494 ( .A(n392), .B(n393), .Z(c[98]) );
  XOR U495 ( .A(a[99]), .B(b[99]), .Z(n396) );
  NAND U496 ( .A(b[98]), .B(a[98]), .Z(n395) );
  NANDN U497 ( .A(n393), .B(n392), .Z(n394) );
  AND U498 ( .A(n395), .B(n394), .Z(n397) );
  XNOR U499 ( .A(n396), .B(n397), .Z(c[99]) );
  XOR U500 ( .A(a[100]), .B(b[100]), .Z(n400) );
  NAND U501 ( .A(b[99]), .B(a[99]), .Z(n399) );
  NANDN U502 ( .A(n397), .B(n396), .Z(n398) );
  AND U503 ( .A(n399), .B(n398), .Z(n401) );
  XNOR U504 ( .A(n400), .B(n401), .Z(c[100]) );
  XOR U505 ( .A(a[101]), .B(b[101]), .Z(n404) );
  NAND U506 ( .A(b[100]), .B(a[100]), .Z(n403) );
  NANDN U507 ( .A(n401), .B(n400), .Z(n402) );
  AND U508 ( .A(n403), .B(n402), .Z(n405) );
  XNOR U509 ( .A(n404), .B(n405), .Z(c[101]) );
  XOR U510 ( .A(a[102]), .B(b[102]), .Z(n408) );
  NAND U511 ( .A(b[101]), .B(a[101]), .Z(n407) );
  NANDN U512 ( .A(n405), .B(n404), .Z(n406) );
  AND U513 ( .A(n407), .B(n406), .Z(n409) );
  XNOR U514 ( .A(n408), .B(n409), .Z(c[102]) );
  XOR U515 ( .A(a[103]), .B(b[103]), .Z(n412) );
  NAND U516 ( .A(b[102]), .B(a[102]), .Z(n411) );
  NANDN U517 ( .A(n409), .B(n408), .Z(n410) );
  AND U518 ( .A(n411), .B(n410), .Z(n413) );
  XNOR U519 ( .A(n412), .B(n413), .Z(c[103]) );
  XOR U520 ( .A(a[104]), .B(b[104]), .Z(n416) );
  NAND U521 ( .A(b[103]), .B(a[103]), .Z(n415) );
  NANDN U522 ( .A(n413), .B(n412), .Z(n414) );
  AND U523 ( .A(n415), .B(n414), .Z(n417) );
  XNOR U524 ( .A(n416), .B(n417), .Z(c[104]) );
  XOR U525 ( .A(a[105]), .B(b[105]), .Z(n420) );
  NAND U526 ( .A(b[104]), .B(a[104]), .Z(n419) );
  NANDN U527 ( .A(n417), .B(n416), .Z(n418) );
  AND U528 ( .A(n419), .B(n418), .Z(n421) );
  XNOR U529 ( .A(n420), .B(n421), .Z(c[105]) );
  XOR U530 ( .A(a[106]), .B(b[106]), .Z(n424) );
  NAND U531 ( .A(b[105]), .B(a[105]), .Z(n423) );
  NANDN U532 ( .A(n421), .B(n420), .Z(n422) );
  AND U533 ( .A(n423), .B(n422), .Z(n425) );
  XNOR U534 ( .A(n424), .B(n425), .Z(c[106]) );
  XOR U535 ( .A(a[107]), .B(b[107]), .Z(n428) );
  NAND U536 ( .A(b[106]), .B(a[106]), .Z(n427) );
  NANDN U537 ( .A(n425), .B(n424), .Z(n426) );
  AND U538 ( .A(n427), .B(n426), .Z(n429) );
  XNOR U539 ( .A(n428), .B(n429), .Z(c[107]) );
  XOR U540 ( .A(a[108]), .B(b[108]), .Z(n432) );
  NAND U541 ( .A(b[107]), .B(a[107]), .Z(n431) );
  NANDN U542 ( .A(n429), .B(n428), .Z(n430) );
  AND U543 ( .A(n431), .B(n430), .Z(n433) );
  XNOR U544 ( .A(n432), .B(n433), .Z(c[108]) );
  XOR U545 ( .A(a[109]), .B(b[109]), .Z(n436) );
  NAND U546 ( .A(b[108]), .B(a[108]), .Z(n435) );
  NANDN U547 ( .A(n433), .B(n432), .Z(n434) );
  AND U548 ( .A(n435), .B(n434), .Z(n437) );
  XNOR U549 ( .A(n436), .B(n437), .Z(c[109]) );
  XOR U550 ( .A(a[110]), .B(b[110]), .Z(n440) );
  NAND U551 ( .A(b[109]), .B(a[109]), .Z(n439) );
  NANDN U552 ( .A(n437), .B(n436), .Z(n438) );
  AND U553 ( .A(n439), .B(n438), .Z(n441) );
  XNOR U554 ( .A(n440), .B(n441), .Z(c[110]) );
  XOR U555 ( .A(a[111]), .B(b[111]), .Z(n444) );
  NAND U556 ( .A(b[110]), .B(a[110]), .Z(n443) );
  NANDN U557 ( .A(n441), .B(n440), .Z(n442) );
  AND U558 ( .A(n443), .B(n442), .Z(n445) );
  XNOR U559 ( .A(n444), .B(n445), .Z(c[111]) );
  XOR U560 ( .A(a[112]), .B(b[112]), .Z(n448) );
  NAND U561 ( .A(b[111]), .B(a[111]), .Z(n447) );
  NANDN U562 ( .A(n445), .B(n444), .Z(n446) );
  AND U563 ( .A(n447), .B(n446), .Z(n449) );
  XNOR U564 ( .A(n448), .B(n449), .Z(c[112]) );
  XOR U565 ( .A(a[113]), .B(b[113]), .Z(n452) );
  NAND U566 ( .A(b[112]), .B(a[112]), .Z(n451) );
  NANDN U567 ( .A(n449), .B(n448), .Z(n450) );
  AND U568 ( .A(n451), .B(n450), .Z(n453) );
  XNOR U569 ( .A(n452), .B(n453), .Z(c[113]) );
  XOR U570 ( .A(a[114]), .B(b[114]), .Z(n456) );
  NAND U571 ( .A(b[113]), .B(a[113]), .Z(n455) );
  NANDN U572 ( .A(n453), .B(n452), .Z(n454) );
  AND U573 ( .A(n455), .B(n454), .Z(n457) );
  XNOR U574 ( .A(n456), .B(n457), .Z(c[114]) );
  XOR U575 ( .A(a[115]), .B(b[115]), .Z(n460) );
  NAND U576 ( .A(b[114]), .B(a[114]), .Z(n459) );
  NANDN U577 ( .A(n457), .B(n456), .Z(n458) );
  AND U578 ( .A(n459), .B(n458), .Z(n461) );
  XNOR U579 ( .A(n460), .B(n461), .Z(c[115]) );
  XOR U580 ( .A(a[116]), .B(b[116]), .Z(n464) );
  NAND U581 ( .A(b[115]), .B(a[115]), .Z(n463) );
  NANDN U582 ( .A(n461), .B(n460), .Z(n462) );
  AND U583 ( .A(n463), .B(n462), .Z(n465) );
  XNOR U584 ( .A(n464), .B(n465), .Z(c[116]) );
  XOR U585 ( .A(a[117]), .B(b[117]), .Z(n468) );
  NAND U586 ( .A(b[116]), .B(a[116]), .Z(n467) );
  NANDN U587 ( .A(n465), .B(n464), .Z(n466) );
  AND U588 ( .A(n467), .B(n466), .Z(n469) );
  XNOR U589 ( .A(n468), .B(n469), .Z(c[117]) );
  XOR U590 ( .A(a[118]), .B(b[118]), .Z(n472) );
  NAND U591 ( .A(b[117]), .B(a[117]), .Z(n471) );
  NANDN U592 ( .A(n469), .B(n468), .Z(n470) );
  AND U593 ( .A(n471), .B(n470), .Z(n473) );
  XNOR U594 ( .A(n472), .B(n473), .Z(c[118]) );
  XOR U595 ( .A(a[119]), .B(b[119]), .Z(n476) );
  NAND U596 ( .A(b[118]), .B(a[118]), .Z(n475) );
  NANDN U597 ( .A(n473), .B(n472), .Z(n474) );
  AND U598 ( .A(n475), .B(n474), .Z(n477) );
  XNOR U599 ( .A(n476), .B(n477), .Z(c[119]) );
  XOR U600 ( .A(a[120]), .B(b[120]), .Z(n480) );
  NAND U601 ( .A(b[119]), .B(a[119]), .Z(n479) );
  NANDN U602 ( .A(n477), .B(n476), .Z(n478) );
  AND U603 ( .A(n479), .B(n478), .Z(n481) );
  XNOR U604 ( .A(n480), .B(n481), .Z(c[120]) );
  XOR U605 ( .A(a[121]), .B(b[121]), .Z(n484) );
  NAND U606 ( .A(b[120]), .B(a[120]), .Z(n483) );
  NANDN U607 ( .A(n481), .B(n480), .Z(n482) );
  AND U608 ( .A(n483), .B(n482), .Z(n485) );
  XNOR U609 ( .A(n484), .B(n485), .Z(c[121]) );
  XOR U610 ( .A(a[122]), .B(b[122]), .Z(n488) );
  NAND U611 ( .A(b[121]), .B(a[121]), .Z(n487) );
  NANDN U612 ( .A(n485), .B(n484), .Z(n486) );
  AND U613 ( .A(n487), .B(n486), .Z(n489) );
  XNOR U614 ( .A(n488), .B(n489), .Z(c[122]) );
  XOR U615 ( .A(a[123]), .B(b[123]), .Z(n492) );
  NAND U616 ( .A(b[122]), .B(a[122]), .Z(n491) );
  NANDN U617 ( .A(n489), .B(n488), .Z(n490) );
  AND U618 ( .A(n491), .B(n490), .Z(n493) );
  XNOR U619 ( .A(n492), .B(n493), .Z(c[123]) );
  XOR U620 ( .A(a[124]), .B(b[124]), .Z(n496) );
  NAND U621 ( .A(b[123]), .B(a[123]), .Z(n495) );
  NANDN U622 ( .A(n493), .B(n492), .Z(n494) );
  AND U623 ( .A(n495), .B(n494), .Z(n497) );
  XNOR U624 ( .A(n496), .B(n497), .Z(c[124]) );
  XOR U625 ( .A(a[125]), .B(b[125]), .Z(n500) );
  NAND U626 ( .A(b[124]), .B(a[124]), .Z(n499) );
  NANDN U627 ( .A(n497), .B(n496), .Z(n498) );
  AND U628 ( .A(n499), .B(n498), .Z(n501) );
  XNOR U629 ( .A(n500), .B(n501), .Z(c[125]) );
  XOR U630 ( .A(a[126]), .B(b[126]), .Z(n504) );
  NAND U631 ( .A(b[125]), .B(a[125]), .Z(n503) );
  NANDN U632 ( .A(n501), .B(n500), .Z(n502) );
  AND U633 ( .A(n503), .B(n502), .Z(n505) );
  XNOR U634 ( .A(n504), .B(n505), .Z(c[126]) );
  XOR U635 ( .A(a[127]), .B(b[127]), .Z(n508) );
  NAND U636 ( .A(b[126]), .B(a[126]), .Z(n507) );
  NANDN U637 ( .A(n505), .B(n504), .Z(n506) );
  AND U638 ( .A(n507), .B(n506), .Z(n509) );
  XNOR U639 ( .A(n508), .B(n509), .Z(c[127]) );
  XOR U640 ( .A(a[128]), .B(b[128]), .Z(n512) );
  NAND U641 ( .A(b[127]), .B(a[127]), .Z(n511) );
  NANDN U642 ( .A(n509), .B(n508), .Z(n510) );
  AND U643 ( .A(n511), .B(n510), .Z(n513) );
  XNOR U644 ( .A(n512), .B(n513), .Z(c[128]) );
  XOR U645 ( .A(a[129]), .B(b[129]), .Z(n516) );
  NAND U646 ( .A(b[128]), .B(a[128]), .Z(n515) );
  NANDN U647 ( .A(n513), .B(n512), .Z(n514) );
  AND U648 ( .A(n515), .B(n514), .Z(n517) );
  XNOR U649 ( .A(n516), .B(n517), .Z(c[129]) );
  XOR U650 ( .A(a[130]), .B(b[130]), .Z(n520) );
  NAND U651 ( .A(b[129]), .B(a[129]), .Z(n519) );
  NANDN U652 ( .A(n517), .B(n516), .Z(n518) );
  AND U653 ( .A(n519), .B(n518), .Z(n521) );
  XNOR U654 ( .A(n520), .B(n521), .Z(c[130]) );
  XOR U655 ( .A(a[131]), .B(b[131]), .Z(n524) );
  NAND U656 ( .A(b[130]), .B(a[130]), .Z(n523) );
  NANDN U657 ( .A(n521), .B(n520), .Z(n522) );
  AND U658 ( .A(n523), .B(n522), .Z(n525) );
  XNOR U659 ( .A(n524), .B(n525), .Z(c[131]) );
  XOR U660 ( .A(a[132]), .B(b[132]), .Z(n528) );
  NAND U661 ( .A(b[131]), .B(a[131]), .Z(n527) );
  NANDN U662 ( .A(n525), .B(n524), .Z(n526) );
  AND U663 ( .A(n527), .B(n526), .Z(n529) );
  XNOR U664 ( .A(n528), .B(n529), .Z(c[132]) );
  XOR U665 ( .A(a[133]), .B(b[133]), .Z(n532) );
  NAND U666 ( .A(b[132]), .B(a[132]), .Z(n531) );
  NANDN U667 ( .A(n529), .B(n528), .Z(n530) );
  AND U668 ( .A(n531), .B(n530), .Z(n533) );
  XNOR U669 ( .A(n532), .B(n533), .Z(c[133]) );
  XOR U670 ( .A(a[134]), .B(b[134]), .Z(n536) );
  NAND U671 ( .A(b[133]), .B(a[133]), .Z(n535) );
  NANDN U672 ( .A(n533), .B(n532), .Z(n534) );
  AND U673 ( .A(n535), .B(n534), .Z(n537) );
  XNOR U674 ( .A(n536), .B(n537), .Z(c[134]) );
  XOR U675 ( .A(a[135]), .B(b[135]), .Z(n540) );
  NAND U676 ( .A(b[134]), .B(a[134]), .Z(n539) );
  NANDN U677 ( .A(n537), .B(n536), .Z(n538) );
  AND U678 ( .A(n539), .B(n538), .Z(n541) );
  XNOR U679 ( .A(n540), .B(n541), .Z(c[135]) );
  XOR U680 ( .A(a[136]), .B(b[136]), .Z(n544) );
  NAND U681 ( .A(b[135]), .B(a[135]), .Z(n543) );
  NANDN U682 ( .A(n541), .B(n540), .Z(n542) );
  AND U683 ( .A(n543), .B(n542), .Z(n545) );
  XNOR U684 ( .A(n544), .B(n545), .Z(c[136]) );
  XOR U685 ( .A(a[137]), .B(b[137]), .Z(n548) );
  NAND U686 ( .A(b[136]), .B(a[136]), .Z(n547) );
  NANDN U687 ( .A(n545), .B(n544), .Z(n546) );
  AND U688 ( .A(n547), .B(n546), .Z(n549) );
  XNOR U689 ( .A(n548), .B(n549), .Z(c[137]) );
  XOR U690 ( .A(a[138]), .B(b[138]), .Z(n552) );
  NAND U691 ( .A(b[137]), .B(a[137]), .Z(n551) );
  NANDN U692 ( .A(n549), .B(n548), .Z(n550) );
  AND U693 ( .A(n551), .B(n550), .Z(n553) );
  XNOR U694 ( .A(n552), .B(n553), .Z(c[138]) );
  XOR U695 ( .A(a[139]), .B(b[139]), .Z(n556) );
  NAND U696 ( .A(b[138]), .B(a[138]), .Z(n555) );
  NANDN U697 ( .A(n553), .B(n552), .Z(n554) );
  AND U698 ( .A(n555), .B(n554), .Z(n557) );
  XNOR U699 ( .A(n556), .B(n557), .Z(c[139]) );
  XOR U700 ( .A(a[140]), .B(b[140]), .Z(n560) );
  NAND U701 ( .A(b[139]), .B(a[139]), .Z(n559) );
  NANDN U702 ( .A(n557), .B(n556), .Z(n558) );
  AND U703 ( .A(n559), .B(n558), .Z(n561) );
  XNOR U704 ( .A(n560), .B(n561), .Z(c[140]) );
  XOR U705 ( .A(a[141]), .B(b[141]), .Z(n564) );
  NAND U706 ( .A(b[140]), .B(a[140]), .Z(n563) );
  NANDN U707 ( .A(n561), .B(n560), .Z(n562) );
  AND U708 ( .A(n563), .B(n562), .Z(n565) );
  XNOR U709 ( .A(n564), .B(n565), .Z(c[141]) );
  XOR U710 ( .A(a[142]), .B(b[142]), .Z(n568) );
  NAND U711 ( .A(b[141]), .B(a[141]), .Z(n567) );
  NANDN U712 ( .A(n565), .B(n564), .Z(n566) );
  AND U713 ( .A(n567), .B(n566), .Z(n569) );
  XNOR U714 ( .A(n568), .B(n569), .Z(c[142]) );
  XOR U715 ( .A(a[143]), .B(b[143]), .Z(n572) );
  NAND U716 ( .A(b[142]), .B(a[142]), .Z(n571) );
  NANDN U717 ( .A(n569), .B(n568), .Z(n570) );
  AND U718 ( .A(n571), .B(n570), .Z(n573) );
  XNOR U719 ( .A(n572), .B(n573), .Z(c[143]) );
  XOR U720 ( .A(a[144]), .B(b[144]), .Z(n576) );
  NAND U721 ( .A(b[143]), .B(a[143]), .Z(n575) );
  NANDN U722 ( .A(n573), .B(n572), .Z(n574) );
  AND U723 ( .A(n575), .B(n574), .Z(n577) );
  XNOR U724 ( .A(n576), .B(n577), .Z(c[144]) );
  XOR U725 ( .A(a[145]), .B(b[145]), .Z(n580) );
  NAND U726 ( .A(b[144]), .B(a[144]), .Z(n579) );
  NANDN U727 ( .A(n577), .B(n576), .Z(n578) );
  AND U728 ( .A(n579), .B(n578), .Z(n581) );
  XNOR U729 ( .A(n580), .B(n581), .Z(c[145]) );
  XOR U730 ( .A(a[146]), .B(b[146]), .Z(n584) );
  NAND U731 ( .A(b[145]), .B(a[145]), .Z(n583) );
  NANDN U732 ( .A(n581), .B(n580), .Z(n582) );
  AND U733 ( .A(n583), .B(n582), .Z(n585) );
  XNOR U734 ( .A(n584), .B(n585), .Z(c[146]) );
  XOR U735 ( .A(a[147]), .B(b[147]), .Z(n588) );
  NAND U736 ( .A(b[146]), .B(a[146]), .Z(n587) );
  NANDN U737 ( .A(n585), .B(n584), .Z(n586) );
  AND U738 ( .A(n587), .B(n586), .Z(n589) );
  XNOR U739 ( .A(n588), .B(n589), .Z(c[147]) );
  XOR U740 ( .A(a[148]), .B(b[148]), .Z(n592) );
  NAND U741 ( .A(b[147]), .B(a[147]), .Z(n591) );
  NANDN U742 ( .A(n589), .B(n588), .Z(n590) );
  AND U743 ( .A(n591), .B(n590), .Z(n593) );
  XNOR U744 ( .A(n592), .B(n593), .Z(c[148]) );
  XOR U745 ( .A(a[149]), .B(b[149]), .Z(n596) );
  NAND U746 ( .A(b[148]), .B(a[148]), .Z(n595) );
  NANDN U747 ( .A(n593), .B(n592), .Z(n594) );
  AND U748 ( .A(n595), .B(n594), .Z(n597) );
  XNOR U749 ( .A(n596), .B(n597), .Z(c[149]) );
  XOR U750 ( .A(a[150]), .B(b[150]), .Z(n600) );
  NAND U751 ( .A(b[149]), .B(a[149]), .Z(n599) );
  NANDN U752 ( .A(n597), .B(n596), .Z(n598) );
  AND U753 ( .A(n599), .B(n598), .Z(n601) );
  XNOR U754 ( .A(n600), .B(n601), .Z(c[150]) );
  XOR U755 ( .A(a[151]), .B(b[151]), .Z(n604) );
  NAND U756 ( .A(b[150]), .B(a[150]), .Z(n603) );
  NANDN U757 ( .A(n601), .B(n600), .Z(n602) );
  AND U758 ( .A(n603), .B(n602), .Z(n605) );
  XNOR U759 ( .A(n604), .B(n605), .Z(c[151]) );
  XOR U760 ( .A(a[152]), .B(b[152]), .Z(n608) );
  NAND U761 ( .A(b[151]), .B(a[151]), .Z(n607) );
  NANDN U762 ( .A(n605), .B(n604), .Z(n606) );
  AND U763 ( .A(n607), .B(n606), .Z(n609) );
  XNOR U764 ( .A(n608), .B(n609), .Z(c[152]) );
  XOR U765 ( .A(a[153]), .B(b[153]), .Z(n612) );
  NAND U766 ( .A(b[152]), .B(a[152]), .Z(n611) );
  NANDN U767 ( .A(n609), .B(n608), .Z(n610) );
  AND U768 ( .A(n611), .B(n610), .Z(n613) );
  XNOR U769 ( .A(n612), .B(n613), .Z(c[153]) );
  XOR U770 ( .A(a[154]), .B(b[154]), .Z(n616) );
  NAND U771 ( .A(b[153]), .B(a[153]), .Z(n615) );
  NANDN U772 ( .A(n613), .B(n612), .Z(n614) );
  AND U773 ( .A(n615), .B(n614), .Z(n617) );
  XNOR U774 ( .A(n616), .B(n617), .Z(c[154]) );
  XOR U775 ( .A(a[155]), .B(b[155]), .Z(n620) );
  NAND U776 ( .A(b[154]), .B(a[154]), .Z(n619) );
  NANDN U777 ( .A(n617), .B(n616), .Z(n618) );
  AND U778 ( .A(n619), .B(n618), .Z(n621) );
  XNOR U779 ( .A(n620), .B(n621), .Z(c[155]) );
  XOR U780 ( .A(a[156]), .B(b[156]), .Z(n624) );
  NAND U781 ( .A(b[155]), .B(a[155]), .Z(n623) );
  NANDN U782 ( .A(n621), .B(n620), .Z(n622) );
  AND U783 ( .A(n623), .B(n622), .Z(n625) );
  XNOR U784 ( .A(n624), .B(n625), .Z(c[156]) );
  XOR U785 ( .A(a[157]), .B(b[157]), .Z(n628) );
  NAND U786 ( .A(b[156]), .B(a[156]), .Z(n627) );
  NANDN U787 ( .A(n625), .B(n624), .Z(n626) );
  AND U788 ( .A(n627), .B(n626), .Z(n629) );
  XNOR U789 ( .A(n628), .B(n629), .Z(c[157]) );
  XOR U790 ( .A(a[158]), .B(b[158]), .Z(n632) );
  NAND U791 ( .A(b[157]), .B(a[157]), .Z(n631) );
  NANDN U792 ( .A(n629), .B(n628), .Z(n630) );
  AND U793 ( .A(n631), .B(n630), .Z(n633) );
  XNOR U794 ( .A(n632), .B(n633), .Z(c[158]) );
  XOR U795 ( .A(a[159]), .B(b[159]), .Z(n636) );
  NAND U796 ( .A(b[158]), .B(a[158]), .Z(n635) );
  NANDN U797 ( .A(n633), .B(n632), .Z(n634) );
  AND U798 ( .A(n635), .B(n634), .Z(n637) );
  XNOR U799 ( .A(n636), .B(n637), .Z(c[159]) );
  XOR U800 ( .A(a[160]), .B(b[160]), .Z(n640) );
  NAND U801 ( .A(b[159]), .B(a[159]), .Z(n639) );
  NANDN U802 ( .A(n637), .B(n636), .Z(n638) );
  AND U803 ( .A(n639), .B(n638), .Z(n641) );
  XNOR U804 ( .A(n640), .B(n641), .Z(c[160]) );
  XOR U805 ( .A(a[161]), .B(b[161]), .Z(n644) );
  NAND U806 ( .A(b[160]), .B(a[160]), .Z(n643) );
  NANDN U807 ( .A(n641), .B(n640), .Z(n642) );
  AND U808 ( .A(n643), .B(n642), .Z(n645) );
  XNOR U809 ( .A(n644), .B(n645), .Z(c[161]) );
  XOR U810 ( .A(a[162]), .B(b[162]), .Z(n648) );
  NAND U811 ( .A(b[161]), .B(a[161]), .Z(n647) );
  NANDN U812 ( .A(n645), .B(n644), .Z(n646) );
  AND U813 ( .A(n647), .B(n646), .Z(n649) );
  XNOR U814 ( .A(n648), .B(n649), .Z(c[162]) );
  XOR U815 ( .A(a[163]), .B(b[163]), .Z(n652) );
  NAND U816 ( .A(b[162]), .B(a[162]), .Z(n651) );
  NANDN U817 ( .A(n649), .B(n648), .Z(n650) );
  AND U818 ( .A(n651), .B(n650), .Z(n653) );
  XNOR U819 ( .A(n652), .B(n653), .Z(c[163]) );
  XOR U820 ( .A(a[164]), .B(b[164]), .Z(n656) );
  NAND U821 ( .A(b[163]), .B(a[163]), .Z(n655) );
  NANDN U822 ( .A(n653), .B(n652), .Z(n654) );
  AND U823 ( .A(n655), .B(n654), .Z(n657) );
  XNOR U824 ( .A(n656), .B(n657), .Z(c[164]) );
  XOR U825 ( .A(a[165]), .B(b[165]), .Z(n660) );
  NAND U826 ( .A(b[164]), .B(a[164]), .Z(n659) );
  NANDN U827 ( .A(n657), .B(n656), .Z(n658) );
  AND U828 ( .A(n659), .B(n658), .Z(n661) );
  XNOR U829 ( .A(n660), .B(n661), .Z(c[165]) );
  XOR U830 ( .A(a[166]), .B(b[166]), .Z(n664) );
  NAND U831 ( .A(b[165]), .B(a[165]), .Z(n663) );
  NANDN U832 ( .A(n661), .B(n660), .Z(n662) );
  AND U833 ( .A(n663), .B(n662), .Z(n665) );
  XNOR U834 ( .A(n664), .B(n665), .Z(c[166]) );
  XOR U835 ( .A(a[167]), .B(b[167]), .Z(n668) );
  NAND U836 ( .A(b[166]), .B(a[166]), .Z(n667) );
  NANDN U837 ( .A(n665), .B(n664), .Z(n666) );
  AND U838 ( .A(n667), .B(n666), .Z(n669) );
  XNOR U839 ( .A(n668), .B(n669), .Z(c[167]) );
  XOR U840 ( .A(a[168]), .B(b[168]), .Z(n672) );
  NAND U841 ( .A(b[167]), .B(a[167]), .Z(n671) );
  NANDN U842 ( .A(n669), .B(n668), .Z(n670) );
  AND U843 ( .A(n671), .B(n670), .Z(n673) );
  XNOR U844 ( .A(n672), .B(n673), .Z(c[168]) );
  XOR U845 ( .A(a[169]), .B(b[169]), .Z(n676) );
  NAND U846 ( .A(b[168]), .B(a[168]), .Z(n675) );
  NANDN U847 ( .A(n673), .B(n672), .Z(n674) );
  AND U848 ( .A(n675), .B(n674), .Z(n677) );
  XNOR U849 ( .A(n676), .B(n677), .Z(c[169]) );
  XOR U850 ( .A(a[170]), .B(b[170]), .Z(n680) );
  NAND U851 ( .A(b[169]), .B(a[169]), .Z(n679) );
  NANDN U852 ( .A(n677), .B(n676), .Z(n678) );
  AND U853 ( .A(n679), .B(n678), .Z(n681) );
  XNOR U854 ( .A(n680), .B(n681), .Z(c[170]) );
  XOR U855 ( .A(a[171]), .B(b[171]), .Z(n684) );
  NAND U856 ( .A(b[170]), .B(a[170]), .Z(n683) );
  NANDN U857 ( .A(n681), .B(n680), .Z(n682) );
  AND U858 ( .A(n683), .B(n682), .Z(n685) );
  XNOR U859 ( .A(n684), .B(n685), .Z(c[171]) );
  XOR U860 ( .A(a[172]), .B(b[172]), .Z(n688) );
  NAND U861 ( .A(b[171]), .B(a[171]), .Z(n687) );
  NANDN U862 ( .A(n685), .B(n684), .Z(n686) );
  AND U863 ( .A(n687), .B(n686), .Z(n689) );
  XNOR U864 ( .A(n688), .B(n689), .Z(c[172]) );
  XOR U865 ( .A(a[173]), .B(b[173]), .Z(n692) );
  NAND U866 ( .A(b[172]), .B(a[172]), .Z(n691) );
  NANDN U867 ( .A(n689), .B(n688), .Z(n690) );
  AND U868 ( .A(n691), .B(n690), .Z(n693) );
  XNOR U869 ( .A(n692), .B(n693), .Z(c[173]) );
  XOR U870 ( .A(a[174]), .B(b[174]), .Z(n696) );
  NAND U871 ( .A(b[173]), .B(a[173]), .Z(n695) );
  NANDN U872 ( .A(n693), .B(n692), .Z(n694) );
  AND U873 ( .A(n695), .B(n694), .Z(n697) );
  XNOR U874 ( .A(n696), .B(n697), .Z(c[174]) );
  XOR U875 ( .A(a[175]), .B(b[175]), .Z(n700) );
  NAND U876 ( .A(b[174]), .B(a[174]), .Z(n699) );
  NANDN U877 ( .A(n697), .B(n696), .Z(n698) );
  AND U878 ( .A(n699), .B(n698), .Z(n701) );
  XNOR U879 ( .A(n700), .B(n701), .Z(c[175]) );
  XOR U880 ( .A(a[176]), .B(b[176]), .Z(n704) );
  NAND U881 ( .A(b[175]), .B(a[175]), .Z(n703) );
  NANDN U882 ( .A(n701), .B(n700), .Z(n702) );
  AND U883 ( .A(n703), .B(n702), .Z(n705) );
  XNOR U884 ( .A(n704), .B(n705), .Z(c[176]) );
  XOR U885 ( .A(a[177]), .B(b[177]), .Z(n708) );
  NAND U886 ( .A(b[176]), .B(a[176]), .Z(n707) );
  NANDN U887 ( .A(n705), .B(n704), .Z(n706) );
  AND U888 ( .A(n707), .B(n706), .Z(n709) );
  XNOR U889 ( .A(n708), .B(n709), .Z(c[177]) );
  XOR U890 ( .A(a[178]), .B(b[178]), .Z(n712) );
  NAND U891 ( .A(b[177]), .B(a[177]), .Z(n711) );
  NANDN U892 ( .A(n709), .B(n708), .Z(n710) );
  AND U893 ( .A(n711), .B(n710), .Z(n713) );
  XNOR U894 ( .A(n712), .B(n713), .Z(c[178]) );
  XOR U895 ( .A(a[179]), .B(b[179]), .Z(n716) );
  NAND U896 ( .A(b[178]), .B(a[178]), .Z(n715) );
  NANDN U897 ( .A(n713), .B(n712), .Z(n714) );
  AND U898 ( .A(n715), .B(n714), .Z(n717) );
  XNOR U899 ( .A(n716), .B(n717), .Z(c[179]) );
  XOR U900 ( .A(a[180]), .B(b[180]), .Z(n720) );
  NAND U901 ( .A(b[179]), .B(a[179]), .Z(n719) );
  NANDN U902 ( .A(n717), .B(n716), .Z(n718) );
  AND U903 ( .A(n719), .B(n718), .Z(n721) );
  XNOR U904 ( .A(n720), .B(n721), .Z(c[180]) );
  XOR U905 ( .A(a[181]), .B(b[181]), .Z(n724) );
  NAND U906 ( .A(b[180]), .B(a[180]), .Z(n723) );
  NANDN U907 ( .A(n721), .B(n720), .Z(n722) );
  AND U908 ( .A(n723), .B(n722), .Z(n725) );
  XNOR U909 ( .A(n724), .B(n725), .Z(c[181]) );
  XOR U910 ( .A(a[182]), .B(b[182]), .Z(n728) );
  NAND U911 ( .A(b[181]), .B(a[181]), .Z(n727) );
  NANDN U912 ( .A(n725), .B(n724), .Z(n726) );
  AND U913 ( .A(n727), .B(n726), .Z(n729) );
  XNOR U914 ( .A(n728), .B(n729), .Z(c[182]) );
  XOR U915 ( .A(a[183]), .B(b[183]), .Z(n732) );
  NAND U916 ( .A(b[182]), .B(a[182]), .Z(n731) );
  NANDN U917 ( .A(n729), .B(n728), .Z(n730) );
  AND U918 ( .A(n731), .B(n730), .Z(n733) );
  XNOR U919 ( .A(n732), .B(n733), .Z(c[183]) );
  XOR U920 ( .A(a[184]), .B(b[184]), .Z(n736) );
  NAND U921 ( .A(b[183]), .B(a[183]), .Z(n735) );
  NANDN U922 ( .A(n733), .B(n732), .Z(n734) );
  AND U923 ( .A(n735), .B(n734), .Z(n737) );
  XNOR U924 ( .A(n736), .B(n737), .Z(c[184]) );
  XOR U925 ( .A(a[185]), .B(b[185]), .Z(n740) );
  NAND U926 ( .A(b[184]), .B(a[184]), .Z(n739) );
  NANDN U927 ( .A(n737), .B(n736), .Z(n738) );
  AND U928 ( .A(n739), .B(n738), .Z(n741) );
  XNOR U929 ( .A(n740), .B(n741), .Z(c[185]) );
  XOR U930 ( .A(a[186]), .B(b[186]), .Z(n744) );
  NAND U931 ( .A(b[185]), .B(a[185]), .Z(n743) );
  NANDN U932 ( .A(n741), .B(n740), .Z(n742) );
  AND U933 ( .A(n743), .B(n742), .Z(n745) );
  XNOR U934 ( .A(n744), .B(n745), .Z(c[186]) );
  XOR U935 ( .A(a[187]), .B(b[187]), .Z(n748) );
  NAND U936 ( .A(b[186]), .B(a[186]), .Z(n747) );
  NANDN U937 ( .A(n745), .B(n744), .Z(n746) );
  AND U938 ( .A(n747), .B(n746), .Z(n749) );
  XNOR U939 ( .A(n748), .B(n749), .Z(c[187]) );
  XOR U940 ( .A(a[188]), .B(b[188]), .Z(n752) );
  NAND U941 ( .A(b[187]), .B(a[187]), .Z(n751) );
  NANDN U942 ( .A(n749), .B(n748), .Z(n750) );
  AND U943 ( .A(n751), .B(n750), .Z(n753) );
  XNOR U944 ( .A(n752), .B(n753), .Z(c[188]) );
  XOR U945 ( .A(a[189]), .B(b[189]), .Z(n756) );
  NAND U946 ( .A(b[188]), .B(a[188]), .Z(n755) );
  NANDN U947 ( .A(n753), .B(n752), .Z(n754) );
  AND U948 ( .A(n755), .B(n754), .Z(n757) );
  XNOR U949 ( .A(n756), .B(n757), .Z(c[189]) );
  XOR U950 ( .A(a[190]), .B(b[190]), .Z(n760) );
  NAND U951 ( .A(b[189]), .B(a[189]), .Z(n759) );
  NANDN U952 ( .A(n757), .B(n756), .Z(n758) );
  AND U953 ( .A(n759), .B(n758), .Z(n761) );
  XNOR U954 ( .A(n760), .B(n761), .Z(c[190]) );
  XOR U955 ( .A(a[191]), .B(b[191]), .Z(n764) );
  NAND U956 ( .A(b[190]), .B(a[190]), .Z(n763) );
  NANDN U957 ( .A(n761), .B(n760), .Z(n762) );
  AND U958 ( .A(n763), .B(n762), .Z(n765) );
  XNOR U959 ( .A(n764), .B(n765), .Z(c[191]) );
  XOR U960 ( .A(a[192]), .B(b[192]), .Z(n768) );
  NAND U961 ( .A(b[191]), .B(a[191]), .Z(n767) );
  NANDN U962 ( .A(n765), .B(n764), .Z(n766) );
  AND U963 ( .A(n767), .B(n766), .Z(n769) );
  XNOR U964 ( .A(n768), .B(n769), .Z(c[192]) );
  XOR U965 ( .A(a[193]), .B(b[193]), .Z(n772) );
  NAND U966 ( .A(b[192]), .B(a[192]), .Z(n771) );
  NANDN U967 ( .A(n769), .B(n768), .Z(n770) );
  AND U968 ( .A(n771), .B(n770), .Z(n773) );
  XNOR U969 ( .A(n772), .B(n773), .Z(c[193]) );
  XOR U970 ( .A(a[194]), .B(b[194]), .Z(n776) );
  NAND U971 ( .A(b[193]), .B(a[193]), .Z(n775) );
  NANDN U972 ( .A(n773), .B(n772), .Z(n774) );
  AND U973 ( .A(n775), .B(n774), .Z(n777) );
  XNOR U974 ( .A(n776), .B(n777), .Z(c[194]) );
  XOR U975 ( .A(a[195]), .B(b[195]), .Z(n780) );
  NAND U976 ( .A(b[194]), .B(a[194]), .Z(n779) );
  NANDN U977 ( .A(n777), .B(n776), .Z(n778) );
  AND U978 ( .A(n779), .B(n778), .Z(n781) );
  XNOR U979 ( .A(n780), .B(n781), .Z(c[195]) );
  XOR U980 ( .A(a[196]), .B(b[196]), .Z(n784) );
  NAND U981 ( .A(b[195]), .B(a[195]), .Z(n783) );
  NANDN U982 ( .A(n781), .B(n780), .Z(n782) );
  AND U983 ( .A(n783), .B(n782), .Z(n785) );
  XNOR U984 ( .A(n784), .B(n785), .Z(c[196]) );
  XOR U985 ( .A(a[197]), .B(b[197]), .Z(n788) );
  NAND U986 ( .A(b[196]), .B(a[196]), .Z(n787) );
  NANDN U987 ( .A(n785), .B(n784), .Z(n786) );
  AND U988 ( .A(n787), .B(n786), .Z(n789) );
  XNOR U989 ( .A(n788), .B(n789), .Z(c[197]) );
  XOR U990 ( .A(a[198]), .B(b[198]), .Z(n792) );
  NAND U991 ( .A(b[197]), .B(a[197]), .Z(n791) );
  NANDN U992 ( .A(n789), .B(n788), .Z(n790) );
  AND U993 ( .A(n791), .B(n790), .Z(n793) );
  XNOR U994 ( .A(n792), .B(n793), .Z(c[198]) );
  XOR U995 ( .A(a[199]), .B(b[199]), .Z(n796) );
  NAND U996 ( .A(b[198]), .B(a[198]), .Z(n795) );
  NANDN U997 ( .A(n793), .B(n792), .Z(n794) );
  AND U998 ( .A(n795), .B(n794), .Z(n797) );
  XNOR U999 ( .A(n796), .B(n797), .Z(c[199]) );
  XOR U1000 ( .A(a[200]), .B(b[200]), .Z(n800) );
  NAND U1001 ( .A(b[199]), .B(a[199]), .Z(n799) );
  NANDN U1002 ( .A(n797), .B(n796), .Z(n798) );
  AND U1003 ( .A(n799), .B(n798), .Z(n801) );
  XNOR U1004 ( .A(n800), .B(n801), .Z(c[200]) );
  XOR U1005 ( .A(a[201]), .B(b[201]), .Z(n804) );
  NAND U1006 ( .A(b[200]), .B(a[200]), .Z(n803) );
  NANDN U1007 ( .A(n801), .B(n800), .Z(n802) );
  AND U1008 ( .A(n803), .B(n802), .Z(n805) );
  XNOR U1009 ( .A(n804), .B(n805), .Z(c[201]) );
  XOR U1010 ( .A(a[202]), .B(b[202]), .Z(n808) );
  NAND U1011 ( .A(b[201]), .B(a[201]), .Z(n807) );
  NANDN U1012 ( .A(n805), .B(n804), .Z(n806) );
  AND U1013 ( .A(n807), .B(n806), .Z(n809) );
  XNOR U1014 ( .A(n808), .B(n809), .Z(c[202]) );
  XOR U1015 ( .A(a[203]), .B(b[203]), .Z(n812) );
  NAND U1016 ( .A(b[202]), .B(a[202]), .Z(n811) );
  NANDN U1017 ( .A(n809), .B(n808), .Z(n810) );
  AND U1018 ( .A(n811), .B(n810), .Z(n813) );
  XNOR U1019 ( .A(n812), .B(n813), .Z(c[203]) );
  XOR U1020 ( .A(a[204]), .B(b[204]), .Z(n816) );
  NAND U1021 ( .A(b[203]), .B(a[203]), .Z(n815) );
  NANDN U1022 ( .A(n813), .B(n812), .Z(n814) );
  AND U1023 ( .A(n815), .B(n814), .Z(n817) );
  XNOR U1024 ( .A(n816), .B(n817), .Z(c[204]) );
  XOR U1025 ( .A(a[205]), .B(b[205]), .Z(n820) );
  NAND U1026 ( .A(b[204]), .B(a[204]), .Z(n819) );
  NANDN U1027 ( .A(n817), .B(n816), .Z(n818) );
  AND U1028 ( .A(n819), .B(n818), .Z(n821) );
  XNOR U1029 ( .A(n820), .B(n821), .Z(c[205]) );
  XOR U1030 ( .A(a[206]), .B(b[206]), .Z(n824) );
  NAND U1031 ( .A(b[205]), .B(a[205]), .Z(n823) );
  NANDN U1032 ( .A(n821), .B(n820), .Z(n822) );
  AND U1033 ( .A(n823), .B(n822), .Z(n825) );
  XNOR U1034 ( .A(n824), .B(n825), .Z(c[206]) );
  XOR U1035 ( .A(a[207]), .B(b[207]), .Z(n828) );
  NAND U1036 ( .A(b[206]), .B(a[206]), .Z(n827) );
  NANDN U1037 ( .A(n825), .B(n824), .Z(n826) );
  AND U1038 ( .A(n827), .B(n826), .Z(n829) );
  XNOR U1039 ( .A(n828), .B(n829), .Z(c[207]) );
  XOR U1040 ( .A(a[208]), .B(b[208]), .Z(n832) );
  NAND U1041 ( .A(b[207]), .B(a[207]), .Z(n831) );
  NANDN U1042 ( .A(n829), .B(n828), .Z(n830) );
  AND U1043 ( .A(n831), .B(n830), .Z(n833) );
  XNOR U1044 ( .A(n832), .B(n833), .Z(c[208]) );
  XOR U1045 ( .A(a[209]), .B(b[209]), .Z(n836) );
  NAND U1046 ( .A(b[208]), .B(a[208]), .Z(n835) );
  NANDN U1047 ( .A(n833), .B(n832), .Z(n834) );
  AND U1048 ( .A(n835), .B(n834), .Z(n837) );
  XNOR U1049 ( .A(n836), .B(n837), .Z(c[209]) );
  XOR U1050 ( .A(a[210]), .B(b[210]), .Z(n840) );
  NAND U1051 ( .A(b[209]), .B(a[209]), .Z(n839) );
  NANDN U1052 ( .A(n837), .B(n836), .Z(n838) );
  AND U1053 ( .A(n839), .B(n838), .Z(n841) );
  XNOR U1054 ( .A(n840), .B(n841), .Z(c[210]) );
  XOR U1055 ( .A(a[211]), .B(b[211]), .Z(n844) );
  NAND U1056 ( .A(b[210]), .B(a[210]), .Z(n843) );
  NANDN U1057 ( .A(n841), .B(n840), .Z(n842) );
  AND U1058 ( .A(n843), .B(n842), .Z(n845) );
  XNOR U1059 ( .A(n844), .B(n845), .Z(c[211]) );
  XOR U1060 ( .A(a[212]), .B(b[212]), .Z(n848) );
  NAND U1061 ( .A(b[211]), .B(a[211]), .Z(n847) );
  NANDN U1062 ( .A(n845), .B(n844), .Z(n846) );
  AND U1063 ( .A(n847), .B(n846), .Z(n849) );
  XNOR U1064 ( .A(n848), .B(n849), .Z(c[212]) );
  XOR U1065 ( .A(a[213]), .B(b[213]), .Z(n852) );
  NAND U1066 ( .A(b[212]), .B(a[212]), .Z(n851) );
  NANDN U1067 ( .A(n849), .B(n848), .Z(n850) );
  AND U1068 ( .A(n851), .B(n850), .Z(n853) );
  XNOR U1069 ( .A(n852), .B(n853), .Z(c[213]) );
  XOR U1070 ( .A(a[214]), .B(b[214]), .Z(n856) );
  NAND U1071 ( .A(b[213]), .B(a[213]), .Z(n855) );
  NANDN U1072 ( .A(n853), .B(n852), .Z(n854) );
  AND U1073 ( .A(n855), .B(n854), .Z(n857) );
  XNOR U1074 ( .A(n856), .B(n857), .Z(c[214]) );
  XOR U1075 ( .A(a[215]), .B(b[215]), .Z(n860) );
  NAND U1076 ( .A(b[214]), .B(a[214]), .Z(n859) );
  NANDN U1077 ( .A(n857), .B(n856), .Z(n858) );
  AND U1078 ( .A(n859), .B(n858), .Z(n861) );
  XNOR U1079 ( .A(n860), .B(n861), .Z(c[215]) );
  XOR U1080 ( .A(a[216]), .B(b[216]), .Z(n864) );
  NAND U1081 ( .A(b[215]), .B(a[215]), .Z(n863) );
  NANDN U1082 ( .A(n861), .B(n860), .Z(n862) );
  AND U1083 ( .A(n863), .B(n862), .Z(n865) );
  XNOR U1084 ( .A(n864), .B(n865), .Z(c[216]) );
  XOR U1085 ( .A(a[217]), .B(b[217]), .Z(n868) );
  NAND U1086 ( .A(b[216]), .B(a[216]), .Z(n867) );
  NANDN U1087 ( .A(n865), .B(n864), .Z(n866) );
  AND U1088 ( .A(n867), .B(n866), .Z(n869) );
  XNOR U1089 ( .A(n868), .B(n869), .Z(c[217]) );
  XOR U1090 ( .A(a[218]), .B(b[218]), .Z(n872) );
  NAND U1091 ( .A(b[217]), .B(a[217]), .Z(n871) );
  NANDN U1092 ( .A(n869), .B(n868), .Z(n870) );
  AND U1093 ( .A(n871), .B(n870), .Z(n873) );
  XNOR U1094 ( .A(n872), .B(n873), .Z(c[218]) );
  XOR U1095 ( .A(a[219]), .B(b[219]), .Z(n876) );
  NAND U1096 ( .A(b[218]), .B(a[218]), .Z(n875) );
  NANDN U1097 ( .A(n873), .B(n872), .Z(n874) );
  AND U1098 ( .A(n875), .B(n874), .Z(n877) );
  XNOR U1099 ( .A(n876), .B(n877), .Z(c[219]) );
  XOR U1100 ( .A(a[220]), .B(b[220]), .Z(n880) );
  NAND U1101 ( .A(b[219]), .B(a[219]), .Z(n879) );
  NANDN U1102 ( .A(n877), .B(n876), .Z(n878) );
  AND U1103 ( .A(n879), .B(n878), .Z(n881) );
  XNOR U1104 ( .A(n880), .B(n881), .Z(c[220]) );
  XOR U1105 ( .A(a[221]), .B(b[221]), .Z(n884) );
  NAND U1106 ( .A(b[220]), .B(a[220]), .Z(n883) );
  NANDN U1107 ( .A(n881), .B(n880), .Z(n882) );
  AND U1108 ( .A(n883), .B(n882), .Z(n885) );
  XNOR U1109 ( .A(n884), .B(n885), .Z(c[221]) );
  XOR U1110 ( .A(a[222]), .B(b[222]), .Z(n888) );
  NAND U1111 ( .A(b[221]), .B(a[221]), .Z(n887) );
  NANDN U1112 ( .A(n885), .B(n884), .Z(n886) );
  AND U1113 ( .A(n887), .B(n886), .Z(n889) );
  XNOR U1114 ( .A(n888), .B(n889), .Z(c[222]) );
  XOR U1115 ( .A(a[223]), .B(b[223]), .Z(n892) );
  NAND U1116 ( .A(b[222]), .B(a[222]), .Z(n891) );
  NANDN U1117 ( .A(n889), .B(n888), .Z(n890) );
  AND U1118 ( .A(n891), .B(n890), .Z(n893) );
  XNOR U1119 ( .A(n892), .B(n893), .Z(c[223]) );
  XOR U1120 ( .A(a[224]), .B(b[224]), .Z(n896) );
  NAND U1121 ( .A(b[223]), .B(a[223]), .Z(n895) );
  NANDN U1122 ( .A(n893), .B(n892), .Z(n894) );
  AND U1123 ( .A(n895), .B(n894), .Z(n897) );
  XNOR U1124 ( .A(n896), .B(n897), .Z(c[224]) );
  XOR U1125 ( .A(a[225]), .B(b[225]), .Z(n900) );
  NAND U1126 ( .A(b[224]), .B(a[224]), .Z(n899) );
  NANDN U1127 ( .A(n897), .B(n896), .Z(n898) );
  AND U1128 ( .A(n899), .B(n898), .Z(n901) );
  XNOR U1129 ( .A(n900), .B(n901), .Z(c[225]) );
  XOR U1130 ( .A(a[226]), .B(b[226]), .Z(n904) );
  NAND U1131 ( .A(b[225]), .B(a[225]), .Z(n903) );
  NANDN U1132 ( .A(n901), .B(n900), .Z(n902) );
  AND U1133 ( .A(n903), .B(n902), .Z(n905) );
  XNOR U1134 ( .A(n904), .B(n905), .Z(c[226]) );
  XOR U1135 ( .A(a[227]), .B(b[227]), .Z(n908) );
  NAND U1136 ( .A(b[226]), .B(a[226]), .Z(n907) );
  NANDN U1137 ( .A(n905), .B(n904), .Z(n906) );
  AND U1138 ( .A(n907), .B(n906), .Z(n909) );
  XNOR U1139 ( .A(n908), .B(n909), .Z(c[227]) );
  XOR U1140 ( .A(a[228]), .B(b[228]), .Z(n912) );
  NAND U1141 ( .A(b[227]), .B(a[227]), .Z(n911) );
  NANDN U1142 ( .A(n909), .B(n908), .Z(n910) );
  AND U1143 ( .A(n911), .B(n910), .Z(n913) );
  XNOR U1144 ( .A(n912), .B(n913), .Z(c[228]) );
  XOR U1145 ( .A(a[229]), .B(b[229]), .Z(n916) );
  NAND U1146 ( .A(b[228]), .B(a[228]), .Z(n915) );
  NANDN U1147 ( .A(n913), .B(n912), .Z(n914) );
  AND U1148 ( .A(n915), .B(n914), .Z(n917) );
  XNOR U1149 ( .A(n916), .B(n917), .Z(c[229]) );
  XOR U1150 ( .A(a[230]), .B(b[230]), .Z(n920) );
  NAND U1151 ( .A(b[229]), .B(a[229]), .Z(n919) );
  NANDN U1152 ( .A(n917), .B(n916), .Z(n918) );
  AND U1153 ( .A(n919), .B(n918), .Z(n921) );
  XNOR U1154 ( .A(n920), .B(n921), .Z(c[230]) );
  XOR U1155 ( .A(a[231]), .B(b[231]), .Z(n924) );
  NAND U1156 ( .A(b[230]), .B(a[230]), .Z(n923) );
  NANDN U1157 ( .A(n921), .B(n920), .Z(n922) );
  AND U1158 ( .A(n923), .B(n922), .Z(n925) );
  XNOR U1159 ( .A(n924), .B(n925), .Z(c[231]) );
  XOR U1160 ( .A(a[232]), .B(b[232]), .Z(n928) );
  NAND U1161 ( .A(b[231]), .B(a[231]), .Z(n927) );
  NANDN U1162 ( .A(n925), .B(n924), .Z(n926) );
  AND U1163 ( .A(n927), .B(n926), .Z(n929) );
  XNOR U1164 ( .A(n928), .B(n929), .Z(c[232]) );
  XOR U1165 ( .A(a[233]), .B(b[233]), .Z(n932) );
  NAND U1166 ( .A(b[232]), .B(a[232]), .Z(n931) );
  NANDN U1167 ( .A(n929), .B(n928), .Z(n930) );
  AND U1168 ( .A(n931), .B(n930), .Z(n933) );
  XNOR U1169 ( .A(n932), .B(n933), .Z(c[233]) );
  XOR U1170 ( .A(a[234]), .B(b[234]), .Z(n936) );
  NAND U1171 ( .A(b[233]), .B(a[233]), .Z(n935) );
  NANDN U1172 ( .A(n933), .B(n932), .Z(n934) );
  AND U1173 ( .A(n935), .B(n934), .Z(n937) );
  XNOR U1174 ( .A(n936), .B(n937), .Z(c[234]) );
  XOR U1175 ( .A(a[235]), .B(b[235]), .Z(n940) );
  NAND U1176 ( .A(b[234]), .B(a[234]), .Z(n939) );
  NANDN U1177 ( .A(n937), .B(n936), .Z(n938) );
  AND U1178 ( .A(n939), .B(n938), .Z(n941) );
  XNOR U1179 ( .A(n940), .B(n941), .Z(c[235]) );
  XOR U1180 ( .A(a[236]), .B(b[236]), .Z(n944) );
  NAND U1181 ( .A(b[235]), .B(a[235]), .Z(n943) );
  NANDN U1182 ( .A(n941), .B(n940), .Z(n942) );
  AND U1183 ( .A(n943), .B(n942), .Z(n945) );
  XNOR U1184 ( .A(n944), .B(n945), .Z(c[236]) );
  XOR U1185 ( .A(a[237]), .B(b[237]), .Z(n948) );
  NAND U1186 ( .A(b[236]), .B(a[236]), .Z(n947) );
  NANDN U1187 ( .A(n945), .B(n944), .Z(n946) );
  AND U1188 ( .A(n947), .B(n946), .Z(n949) );
  XNOR U1189 ( .A(n948), .B(n949), .Z(c[237]) );
  XOR U1190 ( .A(a[238]), .B(b[238]), .Z(n952) );
  NAND U1191 ( .A(b[237]), .B(a[237]), .Z(n951) );
  NANDN U1192 ( .A(n949), .B(n948), .Z(n950) );
  AND U1193 ( .A(n951), .B(n950), .Z(n953) );
  XNOR U1194 ( .A(n952), .B(n953), .Z(c[238]) );
  XOR U1195 ( .A(a[239]), .B(b[239]), .Z(n956) );
  NAND U1196 ( .A(b[238]), .B(a[238]), .Z(n955) );
  NANDN U1197 ( .A(n953), .B(n952), .Z(n954) );
  AND U1198 ( .A(n955), .B(n954), .Z(n957) );
  XNOR U1199 ( .A(n956), .B(n957), .Z(c[239]) );
  XOR U1200 ( .A(a[240]), .B(b[240]), .Z(n960) );
  NAND U1201 ( .A(b[239]), .B(a[239]), .Z(n959) );
  NANDN U1202 ( .A(n957), .B(n956), .Z(n958) );
  AND U1203 ( .A(n959), .B(n958), .Z(n961) );
  XNOR U1204 ( .A(n960), .B(n961), .Z(c[240]) );
  XOR U1205 ( .A(a[241]), .B(b[241]), .Z(n964) );
  NAND U1206 ( .A(b[240]), .B(a[240]), .Z(n963) );
  NANDN U1207 ( .A(n961), .B(n960), .Z(n962) );
  AND U1208 ( .A(n963), .B(n962), .Z(n965) );
  XNOR U1209 ( .A(n964), .B(n965), .Z(c[241]) );
  XOR U1210 ( .A(a[242]), .B(b[242]), .Z(n968) );
  NAND U1211 ( .A(b[241]), .B(a[241]), .Z(n967) );
  NANDN U1212 ( .A(n965), .B(n964), .Z(n966) );
  AND U1213 ( .A(n967), .B(n966), .Z(n969) );
  XNOR U1214 ( .A(n968), .B(n969), .Z(c[242]) );
  XOR U1215 ( .A(a[243]), .B(b[243]), .Z(n972) );
  NAND U1216 ( .A(b[242]), .B(a[242]), .Z(n971) );
  NANDN U1217 ( .A(n969), .B(n968), .Z(n970) );
  AND U1218 ( .A(n971), .B(n970), .Z(n973) );
  XNOR U1219 ( .A(n972), .B(n973), .Z(c[243]) );
  XOR U1220 ( .A(a[244]), .B(b[244]), .Z(n976) );
  NAND U1221 ( .A(b[243]), .B(a[243]), .Z(n975) );
  NANDN U1222 ( .A(n973), .B(n972), .Z(n974) );
  AND U1223 ( .A(n975), .B(n974), .Z(n977) );
  XNOR U1224 ( .A(n976), .B(n977), .Z(c[244]) );
  XOR U1225 ( .A(a[245]), .B(b[245]), .Z(n980) );
  NAND U1226 ( .A(b[244]), .B(a[244]), .Z(n979) );
  NANDN U1227 ( .A(n977), .B(n976), .Z(n978) );
  AND U1228 ( .A(n979), .B(n978), .Z(n981) );
  XNOR U1229 ( .A(n980), .B(n981), .Z(c[245]) );
  XOR U1230 ( .A(a[246]), .B(b[246]), .Z(n984) );
  NAND U1231 ( .A(b[245]), .B(a[245]), .Z(n983) );
  NANDN U1232 ( .A(n981), .B(n980), .Z(n982) );
  AND U1233 ( .A(n983), .B(n982), .Z(n985) );
  XNOR U1234 ( .A(n984), .B(n985), .Z(c[246]) );
  XOR U1235 ( .A(a[247]), .B(b[247]), .Z(n988) );
  NAND U1236 ( .A(b[246]), .B(a[246]), .Z(n987) );
  NANDN U1237 ( .A(n985), .B(n984), .Z(n986) );
  AND U1238 ( .A(n987), .B(n986), .Z(n989) );
  XNOR U1239 ( .A(n988), .B(n989), .Z(c[247]) );
  XOR U1240 ( .A(a[248]), .B(b[248]), .Z(n992) );
  NAND U1241 ( .A(b[247]), .B(a[247]), .Z(n991) );
  NANDN U1242 ( .A(n989), .B(n988), .Z(n990) );
  AND U1243 ( .A(n991), .B(n990), .Z(n993) );
  XNOR U1244 ( .A(n992), .B(n993), .Z(c[248]) );
  XOR U1245 ( .A(a[249]), .B(b[249]), .Z(n996) );
  NAND U1246 ( .A(b[248]), .B(a[248]), .Z(n995) );
  NANDN U1247 ( .A(n993), .B(n992), .Z(n994) );
  AND U1248 ( .A(n995), .B(n994), .Z(n997) );
  XNOR U1249 ( .A(n996), .B(n997), .Z(c[249]) );
  XOR U1250 ( .A(a[250]), .B(b[250]), .Z(n1000) );
  NAND U1251 ( .A(b[249]), .B(a[249]), .Z(n999) );
  NANDN U1252 ( .A(n997), .B(n996), .Z(n998) );
  AND U1253 ( .A(n999), .B(n998), .Z(n1001) );
  XNOR U1254 ( .A(n1000), .B(n1001), .Z(c[250]) );
  XOR U1255 ( .A(a[251]), .B(b[251]), .Z(n1004) );
  NAND U1256 ( .A(b[250]), .B(a[250]), .Z(n1003) );
  NANDN U1257 ( .A(n1001), .B(n1000), .Z(n1002) );
  AND U1258 ( .A(n1003), .B(n1002), .Z(n1005) );
  XNOR U1259 ( .A(n1004), .B(n1005), .Z(c[251]) );
  XOR U1260 ( .A(a[252]), .B(b[252]), .Z(n1008) );
  NAND U1261 ( .A(b[251]), .B(a[251]), .Z(n1007) );
  NANDN U1262 ( .A(n1005), .B(n1004), .Z(n1006) );
  AND U1263 ( .A(n1007), .B(n1006), .Z(n1009) );
  XNOR U1264 ( .A(n1008), .B(n1009), .Z(c[252]) );
  XOR U1265 ( .A(a[253]), .B(b[253]), .Z(n1012) );
  NAND U1266 ( .A(b[252]), .B(a[252]), .Z(n1011) );
  NANDN U1267 ( .A(n1009), .B(n1008), .Z(n1010) );
  AND U1268 ( .A(n1011), .B(n1010), .Z(n1013) );
  XNOR U1269 ( .A(n1012), .B(n1013), .Z(c[253]) );
  XOR U1270 ( .A(a[254]), .B(b[254]), .Z(n1016) );
  NAND U1271 ( .A(b[253]), .B(a[253]), .Z(n1015) );
  NANDN U1272 ( .A(n1013), .B(n1012), .Z(n1014) );
  AND U1273 ( .A(n1015), .B(n1014), .Z(n1017) );
  XNOR U1274 ( .A(n1016), .B(n1017), .Z(c[254]) );
  NAND U1275 ( .A(b[254]), .B(a[254]), .Z(n1019) );
  NANDN U1276 ( .A(n1017), .B(n1016), .Z(n1018) );
  NAND U1277 ( .A(n1019), .B(n1018), .Z(n1020) );
  XOR U1278 ( .A(a[255]), .B(b[255]), .Z(n1021) );
  XOR U1279 ( .A(n1020), .B(n1021), .Z(c[255]) );
  NAND U1280 ( .A(b[255]), .B(a[255]), .Z(n1023) );
  NAND U1281 ( .A(n1021), .B(n1020), .Z(n1022) );
  NAND U1282 ( .A(n1023), .B(n1022), .Z(carry_on_d) );
endmodule

