
module mult_N256_CC16 ( clk, rst, a, b, c );
  input [255:0] a;
  input [15:0] b;
  output [511:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883;
  wire   [511:0] sreg;

  DFF \sreg_reg[495]  ( .D(c[511]), .CLK(clk), .RST(rst), .Q(sreg[495]) );
  DFF \sreg_reg[494]  ( .D(c[510]), .CLK(clk), .RST(rst), .Q(sreg[494]) );
  DFF \sreg_reg[493]  ( .D(c[509]), .CLK(clk), .RST(rst), .Q(sreg[493]) );
  DFF \sreg_reg[492]  ( .D(c[508]), .CLK(clk), .RST(rst), .Q(sreg[492]) );
  DFF \sreg_reg[491]  ( .D(c[507]), .CLK(clk), .RST(rst), .Q(sreg[491]) );
  DFF \sreg_reg[490]  ( .D(c[506]), .CLK(clk), .RST(rst), .Q(sreg[490]) );
  DFF \sreg_reg[489]  ( .D(c[505]), .CLK(clk), .RST(rst), .Q(sreg[489]) );
  DFF \sreg_reg[488]  ( .D(c[504]), .CLK(clk), .RST(rst), .Q(sreg[488]) );
  DFF \sreg_reg[487]  ( .D(c[503]), .CLK(clk), .RST(rst), .Q(sreg[487]) );
  DFF \sreg_reg[486]  ( .D(c[502]), .CLK(clk), .RST(rst), .Q(sreg[486]) );
  DFF \sreg_reg[485]  ( .D(c[501]), .CLK(clk), .RST(rst), .Q(sreg[485]) );
  DFF \sreg_reg[484]  ( .D(c[500]), .CLK(clk), .RST(rst), .Q(sreg[484]) );
  DFF \sreg_reg[483]  ( .D(c[499]), .CLK(clk), .RST(rst), .Q(sreg[483]) );
  DFF \sreg_reg[482]  ( .D(c[498]), .CLK(clk), .RST(rst), .Q(sreg[482]) );
  DFF \sreg_reg[481]  ( .D(c[497]), .CLK(clk), .RST(rst), .Q(sreg[481]) );
  DFF \sreg_reg[480]  ( .D(c[496]), .CLK(clk), .RST(rst), .Q(sreg[480]) );
  DFF \sreg_reg[479]  ( .D(c[495]), .CLK(clk), .RST(rst), .Q(sreg[479]) );
  DFF \sreg_reg[478]  ( .D(c[494]), .CLK(clk), .RST(rst), .Q(sreg[478]) );
  DFF \sreg_reg[477]  ( .D(c[493]), .CLK(clk), .RST(rst), .Q(sreg[477]) );
  DFF \sreg_reg[476]  ( .D(c[492]), .CLK(clk), .RST(rst), .Q(sreg[476]) );
  DFF \sreg_reg[475]  ( .D(c[491]), .CLK(clk), .RST(rst), .Q(sreg[475]) );
  DFF \sreg_reg[474]  ( .D(c[490]), .CLK(clk), .RST(rst), .Q(sreg[474]) );
  DFF \sreg_reg[473]  ( .D(c[489]), .CLK(clk), .RST(rst), .Q(sreg[473]) );
  DFF \sreg_reg[472]  ( .D(c[488]), .CLK(clk), .RST(rst), .Q(sreg[472]) );
  DFF \sreg_reg[471]  ( .D(c[487]), .CLK(clk), .RST(rst), .Q(sreg[471]) );
  DFF \sreg_reg[470]  ( .D(c[486]), .CLK(clk), .RST(rst), .Q(sreg[470]) );
  DFF \sreg_reg[469]  ( .D(c[485]), .CLK(clk), .RST(rst), .Q(sreg[469]) );
  DFF \sreg_reg[468]  ( .D(c[484]), .CLK(clk), .RST(rst), .Q(sreg[468]) );
  DFF \sreg_reg[467]  ( .D(c[483]), .CLK(clk), .RST(rst), .Q(sreg[467]) );
  DFF \sreg_reg[466]  ( .D(c[482]), .CLK(clk), .RST(rst), .Q(sreg[466]) );
  DFF \sreg_reg[465]  ( .D(c[481]), .CLK(clk), .RST(rst), .Q(sreg[465]) );
  DFF \sreg_reg[464]  ( .D(c[480]), .CLK(clk), .RST(rst), .Q(sreg[464]) );
  DFF \sreg_reg[463]  ( .D(c[479]), .CLK(clk), .RST(rst), .Q(sreg[463]) );
  DFF \sreg_reg[462]  ( .D(c[478]), .CLK(clk), .RST(rst), .Q(sreg[462]) );
  DFF \sreg_reg[461]  ( .D(c[477]), .CLK(clk), .RST(rst), .Q(sreg[461]) );
  DFF \sreg_reg[460]  ( .D(c[476]), .CLK(clk), .RST(rst), .Q(sreg[460]) );
  DFF \sreg_reg[459]  ( .D(c[475]), .CLK(clk), .RST(rst), .Q(sreg[459]) );
  DFF \sreg_reg[458]  ( .D(c[474]), .CLK(clk), .RST(rst), .Q(sreg[458]) );
  DFF \sreg_reg[457]  ( .D(c[473]), .CLK(clk), .RST(rst), .Q(sreg[457]) );
  DFF \sreg_reg[456]  ( .D(c[472]), .CLK(clk), .RST(rst), .Q(sreg[456]) );
  DFF \sreg_reg[455]  ( .D(c[471]), .CLK(clk), .RST(rst), .Q(sreg[455]) );
  DFF \sreg_reg[454]  ( .D(c[470]), .CLK(clk), .RST(rst), .Q(sreg[454]) );
  DFF \sreg_reg[453]  ( .D(c[469]), .CLK(clk), .RST(rst), .Q(sreg[453]) );
  DFF \sreg_reg[452]  ( .D(c[468]), .CLK(clk), .RST(rst), .Q(sreg[452]) );
  DFF \sreg_reg[451]  ( .D(c[467]), .CLK(clk), .RST(rst), .Q(sreg[451]) );
  DFF \sreg_reg[450]  ( .D(c[466]), .CLK(clk), .RST(rst), .Q(sreg[450]) );
  DFF \sreg_reg[449]  ( .D(c[465]), .CLK(clk), .RST(rst), .Q(sreg[449]) );
  DFF \sreg_reg[448]  ( .D(c[464]), .CLK(clk), .RST(rst), .Q(sreg[448]) );
  DFF \sreg_reg[447]  ( .D(c[463]), .CLK(clk), .RST(rst), .Q(sreg[447]) );
  DFF \sreg_reg[446]  ( .D(c[462]), .CLK(clk), .RST(rst), .Q(sreg[446]) );
  DFF \sreg_reg[445]  ( .D(c[461]), .CLK(clk), .RST(rst), .Q(sreg[445]) );
  DFF \sreg_reg[444]  ( .D(c[460]), .CLK(clk), .RST(rst), .Q(sreg[444]) );
  DFF \sreg_reg[443]  ( .D(c[459]), .CLK(clk), .RST(rst), .Q(sreg[443]) );
  DFF \sreg_reg[442]  ( .D(c[458]), .CLK(clk), .RST(rst), .Q(sreg[442]) );
  DFF \sreg_reg[441]  ( .D(c[457]), .CLK(clk), .RST(rst), .Q(sreg[441]) );
  DFF \sreg_reg[440]  ( .D(c[456]), .CLK(clk), .RST(rst), .Q(sreg[440]) );
  DFF \sreg_reg[439]  ( .D(c[455]), .CLK(clk), .RST(rst), .Q(sreg[439]) );
  DFF \sreg_reg[438]  ( .D(c[454]), .CLK(clk), .RST(rst), .Q(sreg[438]) );
  DFF \sreg_reg[437]  ( .D(c[453]), .CLK(clk), .RST(rst), .Q(sreg[437]) );
  DFF \sreg_reg[436]  ( .D(c[452]), .CLK(clk), .RST(rst), .Q(sreg[436]) );
  DFF \sreg_reg[435]  ( .D(c[451]), .CLK(clk), .RST(rst), .Q(sreg[435]) );
  DFF \sreg_reg[434]  ( .D(c[450]), .CLK(clk), .RST(rst), .Q(sreg[434]) );
  DFF \sreg_reg[433]  ( .D(c[449]), .CLK(clk), .RST(rst), .Q(sreg[433]) );
  DFF \sreg_reg[432]  ( .D(c[448]), .CLK(clk), .RST(rst), .Q(sreg[432]) );
  DFF \sreg_reg[431]  ( .D(c[447]), .CLK(clk), .RST(rst), .Q(sreg[431]) );
  DFF \sreg_reg[430]  ( .D(c[446]), .CLK(clk), .RST(rst), .Q(sreg[430]) );
  DFF \sreg_reg[429]  ( .D(c[445]), .CLK(clk), .RST(rst), .Q(sreg[429]) );
  DFF \sreg_reg[428]  ( .D(c[444]), .CLK(clk), .RST(rst), .Q(sreg[428]) );
  DFF \sreg_reg[427]  ( .D(c[443]), .CLK(clk), .RST(rst), .Q(sreg[427]) );
  DFF \sreg_reg[426]  ( .D(c[442]), .CLK(clk), .RST(rst), .Q(sreg[426]) );
  DFF \sreg_reg[425]  ( .D(c[441]), .CLK(clk), .RST(rst), .Q(sreg[425]) );
  DFF \sreg_reg[424]  ( .D(c[440]), .CLK(clk), .RST(rst), .Q(sreg[424]) );
  DFF \sreg_reg[423]  ( .D(c[439]), .CLK(clk), .RST(rst), .Q(sreg[423]) );
  DFF \sreg_reg[422]  ( .D(c[438]), .CLK(clk), .RST(rst), .Q(sreg[422]) );
  DFF \sreg_reg[421]  ( .D(c[437]), .CLK(clk), .RST(rst), .Q(sreg[421]) );
  DFF \sreg_reg[420]  ( .D(c[436]), .CLK(clk), .RST(rst), .Q(sreg[420]) );
  DFF \sreg_reg[419]  ( .D(c[435]), .CLK(clk), .RST(rst), .Q(sreg[419]) );
  DFF \sreg_reg[418]  ( .D(c[434]), .CLK(clk), .RST(rst), .Q(sreg[418]) );
  DFF \sreg_reg[417]  ( .D(c[433]), .CLK(clk), .RST(rst), .Q(sreg[417]) );
  DFF \sreg_reg[416]  ( .D(c[432]), .CLK(clk), .RST(rst), .Q(sreg[416]) );
  DFF \sreg_reg[415]  ( .D(c[431]), .CLK(clk), .RST(rst), .Q(sreg[415]) );
  DFF \sreg_reg[414]  ( .D(c[430]), .CLK(clk), .RST(rst), .Q(sreg[414]) );
  DFF \sreg_reg[413]  ( .D(c[429]), .CLK(clk), .RST(rst), .Q(sreg[413]) );
  DFF \sreg_reg[412]  ( .D(c[428]), .CLK(clk), .RST(rst), .Q(sreg[412]) );
  DFF \sreg_reg[411]  ( .D(c[427]), .CLK(clk), .RST(rst), .Q(sreg[411]) );
  DFF \sreg_reg[410]  ( .D(c[426]), .CLK(clk), .RST(rst), .Q(sreg[410]) );
  DFF \sreg_reg[409]  ( .D(c[425]), .CLK(clk), .RST(rst), .Q(sreg[409]) );
  DFF \sreg_reg[408]  ( .D(c[424]), .CLK(clk), .RST(rst), .Q(sreg[408]) );
  DFF \sreg_reg[407]  ( .D(c[423]), .CLK(clk), .RST(rst), .Q(sreg[407]) );
  DFF \sreg_reg[406]  ( .D(c[422]), .CLK(clk), .RST(rst), .Q(sreg[406]) );
  DFF \sreg_reg[405]  ( .D(c[421]), .CLK(clk), .RST(rst), .Q(sreg[405]) );
  DFF \sreg_reg[404]  ( .D(c[420]), .CLK(clk), .RST(rst), .Q(sreg[404]) );
  DFF \sreg_reg[403]  ( .D(c[419]), .CLK(clk), .RST(rst), .Q(sreg[403]) );
  DFF \sreg_reg[402]  ( .D(c[418]), .CLK(clk), .RST(rst), .Q(sreg[402]) );
  DFF \sreg_reg[401]  ( .D(c[417]), .CLK(clk), .RST(rst), .Q(sreg[401]) );
  DFF \sreg_reg[400]  ( .D(c[416]), .CLK(clk), .RST(rst), .Q(sreg[400]) );
  DFF \sreg_reg[399]  ( .D(c[415]), .CLK(clk), .RST(rst), .Q(sreg[399]) );
  DFF \sreg_reg[398]  ( .D(c[414]), .CLK(clk), .RST(rst), .Q(sreg[398]) );
  DFF \sreg_reg[397]  ( .D(c[413]), .CLK(clk), .RST(rst), .Q(sreg[397]) );
  DFF \sreg_reg[396]  ( .D(c[412]), .CLK(clk), .RST(rst), .Q(sreg[396]) );
  DFF \sreg_reg[395]  ( .D(c[411]), .CLK(clk), .RST(rst), .Q(sreg[395]) );
  DFF \sreg_reg[394]  ( .D(c[410]), .CLK(clk), .RST(rst), .Q(sreg[394]) );
  DFF \sreg_reg[393]  ( .D(c[409]), .CLK(clk), .RST(rst), .Q(sreg[393]) );
  DFF \sreg_reg[392]  ( .D(c[408]), .CLK(clk), .RST(rst), .Q(sreg[392]) );
  DFF \sreg_reg[391]  ( .D(c[407]), .CLK(clk), .RST(rst), .Q(sreg[391]) );
  DFF \sreg_reg[390]  ( .D(c[406]), .CLK(clk), .RST(rst), .Q(sreg[390]) );
  DFF \sreg_reg[389]  ( .D(c[405]), .CLK(clk), .RST(rst), .Q(sreg[389]) );
  DFF \sreg_reg[388]  ( .D(c[404]), .CLK(clk), .RST(rst), .Q(sreg[388]) );
  DFF \sreg_reg[387]  ( .D(c[403]), .CLK(clk), .RST(rst), .Q(sreg[387]) );
  DFF \sreg_reg[386]  ( .D(c[402]), .CLK(clk), .RST(rst), .Q(sreg[386]) );
  DFF \sreg_reg[385]  ( .D(c[401]), .CLK(clk), .RST(rst), .Q(sreg[385]) );
  DFF \sreg_reg[384]  ( .D(c[400]), .CLK(clk), .RST(rst), .Q(sreg[384]) );
  DFF \sreg_reg[383]  ( .D(c[399]), .CLK(clk), .RST(rst), .Q(sreg[383]) );
  DFF \sreg_reg[382]  ( .D(c[398]), .CLK(clk), .RST(rst), .Q(sreg[382]) );
  DFF \sreg_reg[381]  ( .D(c[397]), .CLK(clk), .RST(rst), .Q(sreg[381]) );
  DFF \sreg_reg[380]  ( .D(c[396]), .CLK(clk), .RST(rst), .Q(sreg[380]) );
  DFF \sreg_reg[379]  ( .D(c[395]), .CLK(clk), .RST(rst), .Q(sreg[379]) );
  DFF \sreg_reg[378]  ( .D(c[394]), .CLK(clk), .RST(rst), .Q(sreg[378]) );
  DFF \sreg_reg[377]  ( .D(c[393]), .CLK(clk), .RST(rst), .Q(sreg[377]) );
  DFF \sreg_reg[376]  ( .D(c[392]), .CLK(clk), .RST(rst), .Q(sreg[376]) );
  DFF \sreg_reg[375]  ( .D(c[391]), .CLK(clk), .RST(rst), .Q(sreg[375]) );
  DFF \sreg_reg[374]  ( .D(c[390]), .CLK(clk), .RST(rst), .Q(sreg[374]) );
  DFF \sreg_reg[373]  ( .D(c[389]), .CLK(clk), .RST(rst), .Q(sreg[373]) );
  DFF \sreg_reg[372]  ( .D(c[388]), .CLK(clk), .RST(rst), .Q(sreg[372]) );
  DFF \sreg_reg[371]  ( .D(c[387]), .CLK(clk), .RST(rst), .Q(sreg[371]) );
  DFF \sreg_reg[370]  ( .D(c[386]), .CLK(clk), .RST(rst), .Q(sreg[370]) );
  DFF \sreg_reg[369]  ( .D(c[385]), .CLK(clk), .RST(rst), .Q(sreg[369]) );
  DFF \sreg_reg[368]  ( .D(c[384]), .CLK(clk), .RST(rst), .Q(sreg[368]) );
  DFF \sreg_reg[367]  ( .D(c[383]), .CLK(clk), .RST(rst), .Q(sreg[367]) );
  DFF \sreg_reg[366]  ( .D(c[382]), .CLK(clk), .RST(rst), .Q(sreg[366]) );
  DFF \sreg_reg[365]  ( .D(c[381]), .CLK(clk), .RST(rst), .Q(sreg[365]) );
  DFF \sreg_reg[364]  ( .D(c[380]), .CLK(clk), .RST(rst), .Q(sreg[364]) );
  DFF \sreg_reg[363]  ( .D(c[379]), .CLK(clk), .RST(rst), .Q(sreg[363]) );
  DFF \sreg_reg[362]  ( .D(c[378]), .CLK(clk), .RST(rst), .Q(sreg[362]) );
  DFF \sreg_reg[361]  ( .D(c[377]), .CLK(clk), .RST(rst), .Q(sreg[361]) );
  DFF \sreg_reg[360]  ( .D(c[376]), .CLK(clk), .RST(rst), .Q(sreg[360]) );
  DFF \sreg_reg[359]  ( .D(c[375]), .CLK(clk), .RST(rst), .Q(sreg[359]) );
  DFF \sreg_reg[358]  ( .D(c[374]), .CLK(clk), .RST(rst), .Q(sreg[358]) );
  DFF \sreg_reg[357]  ( .D(c[373]), .CLK(clk), .RST(rst), .Q(sreg[357]) );
  DFF \sreg_reg[356]  ( .D(c[372]), .CLK(clk), .RST(rst), .Q(sreg[356]) );
  DFF \sreg_reg[355]  ( .D(c[371]), .CLK(clk), .RST(rst), .Q(sreg[355]) );
  DFF \sreg_reg[354]  ( .D(c[370]), .CLK(clk), .RST(rst), .Q(sreg[354]) );
  DFF \sreg_reg[353]  ( .D(c[369]), .CLK(clk), .RST(rst), .Q(sreg[353]) );
  DFF \sreg_reg[352]  ( .D(c[368]), .CLK(clk), .RST(rst), .Q(sreg[352]) );
  DFF \sreg_reg[351]  ( .D(c[367]), .CLK(clk), .RST(rst), .Q(sreg[351]) );
  DFF \sreg_reg[350]  ( .D(c[366]), .CLK(clk), .RST(rst), .Q(sreg[350]) );
  DFF \sreg_reg[349]  ( .D(c[365]), .CLK(clk), .RST(rst), .Q(sreg[349]) );
  DFF \sreg_reg[348]  ( .D(c[364]), .CLK(clk), .RST(rst), .Q(sreg[348]) );
  DFF \sreg_reg[347]  ( .D(c[363]), .CLK(clk), .RST(rst), .Q(sreg[347]) );
  DFF \sreg_reg[346]  ( .D(c[362]), .CLK(clk), .RST(rst), .Q(sreg[346]) );
  DFF \sreg_reg[345]  ( .D(c[361]), .CLK(clk), .RST(rst), .Q(sreg[345]) );
  DFF \sreg_reg[344]  ( .D(c[360]), .CLK(clk), .RST(rst), .Q(sreg[344]) );
  DFF \sreg_reg[343]  ( .D(c[359]), .CLK(clk), .RST(rst), .Q(sreg[343]) );
  DFF \sreg_reg[342]  ( .D(c[358]), .CLK(clk), .RST(rst), .Q(sreg[342]) );
  DFF \sreg_reg[341]  ( .D(c[357]), .CLK(clk), .RST(rst), .Q(sreg[341]) );
  DFF \sreg_reg[340]  ( .D(c[356]), .CLK(clk), .RST(rst), .Q(sreg[340]) );
  DFF \sreg_reg[339]  ( .D(c[355]), .CLK(clk), .RST(rst), .Q(sreg[339]) );
  DFF \sreg_reg[338]  ( .D(c[354]), .CLK(clk), .RST(rst), .Q(sreg[338]) );
  DFF \sreg_reg[337]  ( .D(c[353]), .CLK(clk), .RST(rst), .Q(sreg[337]) );
  DFF \sreg_reg[336]  ( .D(c[352]), .CLK(clk), .RST(rst), .Q(sreg[336]) );
  DFF \sreg_reg[335]  ( .D(c[351]), .CLK(clk), .RST(rst), .Q(sreg[335]) );
  DFF \sreg_reg[334]  ( .D(c[350]), .CLK(clk), .RST(rst), .Q(sreg[334]) );
  DFF \sreg_reg[333]  ( .D(c[349]), .CLK(clk), .RST(rst), .Q(sreg[333]) );
  DFF \sreg_reg[332]  ( .D(c[348]), .CLK(clk), .RST(rst), .Q(sreg[332]) );
  DFF \sreg_reg[331]  ( .D(c[347]), .CLK(clk), .RST(rst), .Q(sreg[331]) );
  DFF \sreg_reg[330]  ( .D(c[346]), .CLK(clk), .RST(rst), .Q(sreg[330]) );
  DFF \sreg_reg[329]  ( .D(c[345]), .CLK(clk), .RST(rst), .Q(sreg[329]) );
  DFF \sreg_reg[328]  ( .D(c[344]), .CLK(clk), .RST(rst), .Q(sreg[328]) );
  DFF \sreg_reg[327]  ( .D(c[343]), .CLK(clk), .RST(rst), .Q(sreg[327]) );
  DFF \sreg_reg[326]  ( .D(c[342]), .CLK(clk), .RST(rst), .Q(sreg[326]) );
  DFF \sreg_reg[325]  ( .D(c[341]), .CLK(clk), .RST(rst), .Q(sreg[325]) );
  DFF \sreg_reg[324]  ( .D(c[340]), .CLK(clk), .RST(rst), .Q(sreg[324]) );
  DFF \sreg_reg[323]  ( .D(c[339]), .CLK(clk), .RST(rst), .Q(sreg[323]) );
  DFF \sreg_reg[322]  ( .D(c[338]), .CLK(clk), .RST(rst), .Q(sreg[322]) );
  DFF \sreg_reg[321]  ( .D(c[337]), .CLK(clk), .RST(rst), .Q(sreg[321]) );
  DFF \sreg_reg[320]  ( .D(c[336]), .CLK(clk), .RST(rst), .Q(sreg[320]) );
  DFF \sreg_reg[319]  ( .D(c[335]), .CLK(clk), .RST(rst), .Q(sreg[319]) );
  DFF \sreg_reg[318]  ( .D(c[334]), .CLK(clk), .RST(rst), .Q(sreg[318]) );
  DFF \sreg_reg[317]  ( .D(c[333]), .CLK(clk), .RST(rst), .Q(sreg[317]) );
  DFF \sreg_reg[316]  ( .D(c[332]), .CLK(clk), .RST(rst), .Q(sreg[316]) );
  DFF \sreg_reg[315]  ( .D(c[331]), .CLK(clk), .RST(rst), .Q(sreg[315]) );
  DFF \sreg_reg[314]  ( .D(c[330]), .CLK(clk), .RST(rst), .Q(sreg[314]) );
  DFF \sreg_reg[313]  ( .D(c[329]), .CLK(clk), .RST(rst), .Q(sreg[313]) );
  DFF \sreg_reg[312]  ( .D(c[328]), .CLK(clk), .RST(rst), .Q(sreg[312]) );
  DFF \sreg_reg[311]  ( .D(c[327]), .CLK(clk), .RST(rst), .Q(sreg[311]) );
  DFF \sreg_reg[310]  ( .D(c[326]), .CLK(clk), .RST(rst), .Q(sreg[310]) );
  DFF \sreg_reg[309]  ( .D(c[325]), .CLK(clk), .RST(rst), .Q(sreg[309]) );
  DFF \sreg_reg[308]  ( .D(c[324]), .CLK(clk), .RST(rst), .Q(sreg[308]) );
  DFF \sreg_reg[307]  ( .D(c[323]), .CLK(clk), .RST(rst), .Q(sreg[307]) );
  DFF \sreg_reg[306]  ( .D(c[322]), .CLK(clk), .RST(rst), .Q(sreg[306]) );
  DFF \sreg_reg[305]  ( .D(c[321]), .CLK(clk), .RST(rst), .Q(sreg[305]) );
  DFF \sreg_reg[304]  ( .D(c[320]), .CLK(clk), .RST(rst), .Q(sreg[304]) );
  DFF \sreg_reg[303]  ( .D(c[319]), .CLK(clk), .RST(rst), .Q(sreg[303]) );
  DFF \sreg_reg[302]  ( .D(c[318]), .CLK(clk), .RST(rst), .Q(sreg[302]) );
  DFF \sreg_reg[301]  ( .D(c[317]), .CLK(clk), .RST(rst), .Q(sreg[301]) );
  DFF \sreg_reg[300]  ( .D(c[316]), .CLK(clk), .RST(rst), .Q(sreg[300]) );
  DFF \sreg_reg[299]  ( .D(c[315]), .CLK(clk), .RST(rst), .Q(sreg[299]) );
  DFF \sreg_reg[298]  ( .D(c[314]), .CLK(clk), .RST(rst), .Q(sreg[298]) );
  DFF \sreg_reg[297]  ( .D(c[313]), .CLK(clk), .RST(rst), .Q(sreg[297]) );
  DFF \sreg_reg[296]  ( .D(c[312]), .CLK(clk), .RST(rst), .Q(sreg[296]) );
  DFF \sreg_reg[295]  ( .D(c[311]), .CLK(clk), .RST(rst), .Q(sreg[295]) );
  DFF \sreg_reg[294]  ( .D(c[310]), .CLK(clk), .RST(rst), .Q(sreg[294]) );
  DFF \sreg_reg[293]  ( .D(c[309]), .CLK(clk), .RST(rst), .Q(sreg[293]) );
  DFF \sreg_reg[292]  ( .D(c[308]), .CLK(clk), .RST(rst), .Q(sreg[292]) );
  DFF \sreg_reg[291]  ( .D(c[307]), .CLK(clk), .RST(rst), .Q(sreg[291]) );
  DFF \sreg_reg[290]  ( .D(c[306]), .CLK(clk), .RST(rst), .Q(sreg[290]) );
  DFF \sreg_reg[289]  ( .D(c[305]), .CLK(clk), .RST(rst), .Q(sreg[289]) );
  DFF \sreg_reg[288]  ( .D(c[304]), .CLK(clk), .RST(rst), .Q(sreg[288]) );
  DFF \sreg_reg[287]  ( .D(c[303]), .CLK(clk), .RST(rst), .Q(sreg[287]) );
  DFF \sreg_reg[286]  ( .D(c[302]), .CLK(clk), .RST(rst), .Q(sreg[286]) );
  DFF \sreg_reg[285]  ( .D(c[301]), .CLK(clk), .RST(rst), .Q(sreg[285]) );
  DFF \sreg_reg[284]  ( .D(c[300]), .CLK(clk), .RST(rst), .Q(sreg[284]) );
  DFF \sreg_reg[283]  ( .D(c[299]), .CLK(clk), .RST(rst), .Q(sreg[283]) );
  DFF \sreg_reg[282]  ( .D(c[298]), .CLK(clk), .RST(rst), .Q(sreg[282]) );
  DFF \sreg_reg[281]  ( .D(c[297]), .CLK(clk), .RST(rst), .Q(sreg[281]) );
  DFF \sreg_reg[280]  ( .D(c[296]), .CLK(clk), .RST(rst), .Q(sreg[280]) );
  DFF \sreg_reg[279]  ( .D(c[295]), .CLK(clk), .RST(rst), .Q(sreg[279]) );
  DFF \sreg_reg[278]  ( .D(c[294]), .CLK(clk), .RST(rst), .Q(sreg[278]) );
  DFF \sreg_reg[277]  ( .D(c[293]), .CLK(clk), .RST(rst), .Q(sreg[277]) );
  DFF \sreg_reg[276]  ( .D(c[292]), .CLK(clk), .RST(rst), .Q(sreg[276]) );
  DFF \sreg_reg[275]  ( .D(c[291]), .CLK(clk), .RST(rst), .Q(sreg[275]) );
  DFF \sreg_reg[274]  ( .D(c[290]), .CLK(clk), .RST(rst), .Q(sreg[274]) );
  DFF \sreg_reg[273]  ( .D(c[289]), .CLK(clk), .RST(rst), .Q(sreg[273]) );
  DFF \sreg_reg[272]  ( .D(c[288]), .CLK(clk), .RST(rst), .Q(sreg[272]) );
  DFF \sreg_reg[271]  ( .D(c[287]), .CLK(clk), .RST(rst), .Q(sreg[271]) );
  DFF \sreg_reg[270]  ( .D(c[286]), .CLK(clk), .RST(rst), .Q(sreg[270]) );
  DFF \sreg_reg[269]  ( .D(c[285]), .CLK(clk), .RST(rst), .Q(sreg[269]) );
  DFF \sreg_reg[268]  ( .D(c[284]), .CLK(clk), .RST(rst), .Q(sreg[268]) );
  DFF \sreg_reg[267]  ( .D(c[283]), .CLK(clk), .RST(rst), .Q(sreg[267]) );
  DFF \sreg_reg[266]  ( .D(c[282]), .CLK(clk), .RST(rst), .Q(sreg[266]) );
  DFF \sreg_reg[265]  ( .D(c[281]), .CLK(clk), .RST(rst), .Q(sreg[265]) );
  DFF \sreg_reg[264]  ( .D(c[280]), .CLK(clk), .RST(rst), .Q(sreg[264]) );
  DFF \sreg_reg[263]  ( .D(c[279]), .CLK(clk), .RST(rst), .Q(sreg[263]) );
  DFF \sreg_reg[262]  ( .D(c[278]), .CLK(clk), .RST(rst), .Q(sreg[262]) );
  DFF \sreg_reg[261]  ( .D(c[277]), .CLK(clk), .RST(rst), .Q(sreg[261]) );
  DFF \sreg_reg[260]  ( .D(c[276]), .CLK(clk), .RST(rst), .Q(sreg[260]) );
  DFF \sreg_reg[259]  ( .D(c[275]), .CLK(clk), .RST(rst), .Q(sreg[259]) );
  DFF \sreg_reg[258]  ( .D(c[274]), .CLK(clk), .RST(rst), .Q(sreg[258]) );
  DFF \sreg_reg[257]  ( .D(c[273]), .CLK(clk), .RST(rst), .Q(sreg[257]) );
  DFF \sreg_reg[256]  ( .D(c[272]), .CLK(clk), .RST(rst), .Q(sreg[256]) );
  DFF \sreg_reg[255]  ( .D(c[271]), .CLK(clk), .RST(rst), .Q(sreg[255]) );
  DFF \sreg_reg[254]  ( .D(c[270]), .CLK(clk), .RST(rst), .Q(sreg[254]) );
  DFF \sreg_reg[253]  ( .D(c[269]), .CLK(clk), .RST(rst), .Q(sreg[253]) );
  DFF \sreg_reg[252]  ( .D(c[268]), .CLK(clk), .RST(rst), .Q(sreg[252]) );
  DFF \sreg_reg[251]  ( .D(c[267]), .CLK(clk), .RST(rst), .Q(sreg[251]) );
  DFF \sreg_reg[250]  ( .D(c[266]), .CLK(clk), .RST(rst), .Q(sreg[250]) );
  DFF \sreg_reg[249]  ( .D(c[265]), .CLK(clk), .RST(rst), .Q(sreg[249]) );
  DFF \sreg_reg[248]  ( .D(c[264]), .CLK(clk), .RST(rst), .Q(sreg[248]) );
  DFF \sreg_reg[247]  ( .D(c[263]), .CLK(clk), .RST(rst), .Q(sreg[247]) );
  DFF \sreg_reg[246]  ( .D(c[262]), .CLK(clk), .RST(rst), .Q(sreg[246]) );
  DFF \sreg_reg[245]  ( .D(c[261]), .CLK(clk), .RST(rst), .Q(sreg[245]) );
  DFF \sreg_reg[244]  ( .D(c[260]), .CLK(clk), .RST(rst), .Q(sreg[244]) );
  DFF \sreg_reg[243]  ( .D(c[259]), .CLK(clk), .RST(rst), .Q(sreg[243]) );
  DFF \sreg_reg[242]  ( .D(c[258]), .CLK(clk), .RST(rst), .Q(sreg[242]) );
  DFF \sreg_reg[241]  ( .D(c[257]), .CLK(clk), .RST(rst), .Q(sreg[241]) );
  DFF \sreg_reg[240]  ( .D(c[256]), .CLK(clk), .RST(rst), .Q(sreg[240]) );
  DFF \sreg_reg[239]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(c[239]) );
  DFF \sreg_reg[238]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(c[238]) );
  DFF \sreg_reg[237]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(c[237]) );
  DFF \sreg_reg[236]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(c[236]) );
  DFF \sreg_reg[235]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(c[235]) );
  DFF \sreg_reg[234]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(c[234]) );
  DFF \sreg_reg[233]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(c[233]) );
  DFF \sreg_reg[232]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(c[232]) );
  DFF \sreg_reg[231]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(c[231]) );
  DFF \sreg_reg[230]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(c[230]) );
  DFF \sreg_reg[229]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(c[229]) );
  DFF \sreg_reg[228]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(c[228]) );
  DFF \sreg_reg[227]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(c[227]) );
  DFF \sreg_reg[226]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(c[226]) );
  DFF \sreg_reg[225]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(c[225]) );
  DFF \sreg_reg[224]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(c[224]) );
  DFF \sreg_reg[223]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(c[223]) );
  DFF \sreg_reg[222]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(c[222]) );
  DFF \sreg_reg[221]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(c[221]) );
  DFF \sreg_reg[220]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(c[220]) );
  DFF \sreg_reg[219]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(c[219]) );
  DFF \sreg_reg[218]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(c[218]) );
  DFF \sreg_reg[217]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(c[217]) );
  DFF \sreg_reg[216]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(c[216]) );
  DFF \sreg_reg[215]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(c[215]) );
  DFF \sreg_reg[214]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(c[214]) );
  DFF \sreg_reg[213]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(c[213]) );
  DFF \sreg_reg[212]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(c[212]) );
  DFF \sreg_reg[211]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(c[211]) );
  DFF \sreg_reg[210]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(c[210]) );
  DFF \sreg_reg[209]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(c[209]) );
  DFF \sreg_reg[208]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(c[208]) );
  DFF \sreg_reg[207]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(c[207]) );
  DFF \sreg_reg[206]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(c[206]) );
  DFF \sreg_reg[205]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(c[205]) );
  DFF \sreg_reg[204]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(c[204]) );
  DFF \sreg_reg[203]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(c[203]) );
  DFF \sreg_reg[202]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(c[202]) );
  DFF \sreg_reg[201]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(c[201]) );
  DFF \sreg_reg[200]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(c[200]) );
  DFF \sreg_reg[199]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(c[199]) );
  DFF \sreg_reg[198]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(c[198]) );
  DFF \sreg_reg[197]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(c[197]) );
  DFF \sreg_reg[196]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(c[196]) );
  DFF \sreg_reg[195]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(c[195]) );
  DFF \sreg_reg[194]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(c[194]) );
  DFF \sreg_reg[193]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(c[193]) );
  DFF \sreg_reg[192]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(c[192]) );
  DFF \sreg_reg[191]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(c[191]) );
  DFF \sreg_reg[190]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(c[190]) );
  DFF \sreg_reg[189]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(c[189]) );
  DFF \sreg_reg[188]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(c[188]) );
  DFF \sreg_reg[187]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(c[187]) );
  DFF \sreg_reg[186]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(c[186]) );
  DFF \sreg_reg[185]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(c[185]) );
  DFF \sreg_reg[184]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(c[184]) );
  DFF \sreg_reg[183]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(c[183]) );
  DFF \sreg_reg[182]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(c[182]) );
  DFF \sreg_reg[181]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(c[181]) );
  DFF \sreg_reg[180]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(c[180]) );
  DFF \sreg_reg[179]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(c[179]) );
  DFF \sreg_reg[178]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(c[178]) );
  DFF \sreg_reg[177]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(c[177]) );
  DFF \sreg_reg[176]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(c[176]) );
  DFF \sreg_reg[175]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(c[175]) );
  DFF \sreg_reg[174]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(c[174]) );
  DFF \sreg_reg[173]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(c[173]) );
  DFF \sreg_reg[172]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(c[172]) );
  DFF \sreg_reg[171]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(c[171]) );
  DFF \sreg_reg[170]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(c[170]) );
  DFF \sreg_reg[169]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(c[169]) );
  DFF \sreg_reg[168]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(c[168]) );
  DFF \sreg_reg[167]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(c[167]) );
  DFF \sreg_reg[166]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(c[166]) );
  DFF \sreg_reg[165]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(c[165]) );
  DFF \sreg_reg[164]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(c[164]) );
  DFF \sreg_reg[163]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(c[163]) );
  DFF \sreg_reg[162]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(c[162]) );
  DFF \sreg_reg[161]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(c[161]) );
  DFF \sreg_reg[160]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(c[160]) );
  DFF \sreg_reg[159]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(c[159]) );
  DFF \sreg_reg[158]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(c[158]) );
  DFF \sreg_reg[157]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(c[157]) );
  DFF \sreg_reg[156]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(c[156]) );
  DFF \sreg_reg[155]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(c[155]) );
  DFF \sreg_reg[154]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(c[154]) );
  DFF \sreg_reg[153]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(c[153]) );
  DFF \sreg_reg[152]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(c[152]) );
  DFF \sreg_reg[151]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(c[151]) );
  DFF \sreg_reg[150]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(c[150]) );
  DFF \sreg_reg[149]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(c[149]) );
  DFF \sreg_reg[148]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(c[148]) );
  DFF \sreg_reg[147]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(c[147]) );
  DFF \sreg_reg[146]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(c[146]) );
  DFF \sreg_reg[145]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(c[145]) );
  DFF \sreg_reg[144]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(c[144]) );
  DFF \sreg_reg[143]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(c[143]) );
  DFF \sreg_reg[142]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(c[142]) );
  DFF \sreg_reg[141]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(c[141]) );
  DFF \sreg_reg[140]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(c[140]) );
  DFF \sreg_reg[139]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(c[139]) );
  DFF \sreg_reg[138]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(c[138]) );
  DFF \sreg_reg[137]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(c[137]) );
  DFF \sreg_reg[136]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(c[136]) );
  DFF \sreg_reg[135]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(c[135]) );
  DFF \sreg_reg[134]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(c[134]) );
  DFF \sreg_reg[133]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(c[133]) );
  DFF \sreg_reg[132]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(c[132]) );
  DFF \sreg_reg[131]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(c[131]) );
  DFF \sreg_reg[130]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(c[130]) );
  DFF \sreg_reg[129]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(c[129]) );
  DFF \sreg_reg[128]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(c[128]) );
  DFF \sreg_reg[127]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(c[127]) );
  DFF \sreg_reg[126]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[125]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[124]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[123]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NANDN U19 ( .A(n19590), .B(n19589), .Z(n1) );
  NANDN U20 ( .A(n19644), .B(n19588), .Z(n2) );
  NAND U21 ( .A(n1), .B(n2), .Z(n19625) );
  NAND U22 ( .A(n19690), .B(n19689), .Z(n3) );
  NANDN U23 ( .A(n19732), .B(n19688), .Z(n4) );
  NAND U24 ( .A(n3), .B(n4), .Z(n19712) );
  XOR U25 ( .A(n18919), .B(n18918), .Z(n18920) );
  XOR U26 ( .A(n19146), .B(n19145), .Z(n19147) );
  XOR U27 ( .A(n19402), .B(n19401), .Z(n19435) );
  NAND U28 ( .A(n19433), .B(n19808), .Z(n5) );
  NANDN U29 ( .A(n19434), .B(n19496), .Z(n6) );
  AND U30 ( .A(n5), .B(n6), .Z(n19474) );
  XNOR U31 ( .A(n19054), .B(n19053), .Z(n19024) );
  XNOR U32 ( .A(n19133), .B(n19132), .Z(n19106) );
  XNOR U33 ( .A(n19225), .B(n19224), .Z(n19177) );
  XNOR U34 ( .A(n19294), .B(n19293), .Z(n19248) );
  NAND U35 ( .A(n19504), .B(n19503), .Z(n7) );
  NANDN U36 ( .A(n19554), .B(n19502), .Z(n8) );
  AND U37 ( .A(n7), .B(n8), .Z(n19520) );
  XOR U38 ( .A(n19659), .B(n19658), .Z(n19624) );
  XOR U39 ( .A(n19685), .B(n19684), .Z(n19678) );
  XOR U40 ( .A(n19710), .B(n19709), .Z(n19711) );
  XOR U41 ( .A(n19759), .B(n19758), .Z(n19760) );
  XNOR U42 ( .A(n19580), .B(n19581), .Z(n9) );
  XNOR U43 ( .A(n19579), .B(n9), .Z(n19573) );
  XOR U44 ( .A(n19827), .B(n19826), .Z(n19830) );
  NANDN U45 ( .A(b[0]), .B(a[255]), .Z(n10) );
  AND U46 ( .A(b[1]), .B(n10), .Z(n19205) );
  XOR U47 ( .A(n18990), .B(n18989), .Z(n18991) );
  XOR U48 ( .A(n18996), .B(n18995), .Z(n18997) );
  XOR U49 ( .A(n19067), .B(n19066), .Z(n19068) );
  XOR U50 ( .A(n19073), .B(n19072), .Z(n19074) );
  XOR U51 ( .A(n19324), .B(n19323), .Z(n19325) );
  XOR U52 ( .A(n19436), .B(n19435), .Z(n19438) );
  XOR U53 ( .A(n19480), .B(n19479), .Z(n19481) );
  XOR U54 ( .A(n19542), .B(n19541), .Z(n19543) );
  XOR U55 ( .A(n19548), .B(n19547), .Z(n19550) );
  NANDN U56 ( .A(n18902), .B(n18901), .Z(n11) );
  NANDN U57 ( .A(n18899), .B(n18900), .Z(n12) );
  AND U58 ( .A(n11), .B(n12), .Z(n18948) );
  XOR U59 ( .A(n19231), .B(n19230), .Z(n19179) );
  XOR U60 ( .A(n19300), .B(n19299), .Z(n19251) );
  XOR U61 ( .A(n19368), .B(n19367), .Z(n19369) );
  XOR U62 ( .A(n19444), .B(n19443), .Z(n19395) );
  XOR U63 ( .A(n19677), .B(n19676), .Z(n19679) );
  XOR U64 ( .A(n19775), .B(n19774), .Z(n19761) );
  XOR U65 ( .A(n19085), .B(n19084), .Z(n19086) );
  XOR U66 ( .A(n19164), .B(n19163), .Z(n19165) );
  XOR U67 ( .A(n19522), .B(n19521), .Z(n19513) );
  XOR U68 ( .A(n19574), .B(n19573), .Z(n19575) );
  XNOR U69 ( .A(n19627), .B(n19626), .Z(n19619) );
  XOR U70 ( .A(n19712), .B(n19711), .Z(n19738) );
  XOR U71 ( .A(n19793), .B(n19792), .Z(n19795) );
  XOR U72 ( .A(n19850), .B(n19849), .Z(n19851) );
  XOR U73 ( .A(n19205), .B(n19204), .Z(n19206) );
  XNOR U74 ( .A(n18921), .B(n18920), .Z(n18899) );
  XOR U75 ( .A(n19152), .B(n19151), .Z(n19153) );
  XOR U76 ( .A(n19193), .B(n19192), .Z(n19194) );
  XOR U77 ( .A(n19201), .B(n19200), .Z(n19222) );
  XOR U78 ( .A(n19276), .B(n19275), .Z(n19277) );
  XOR U79 ( .A(n19283), .B(n19282), .Z(n19291) );
  XOR U80 ( .A(n19356), .B(n19355), .Z(n19357) );
  XOR U81 ( .A(n19352), .B(n19351), .Z(n19323) );
  XOR U82 ( .A(n19412), .B(n19411), .Z(n19414) );
  XNOR U83 ( .A(n19482), .B(n19481), .Z(n19473) );
  XOR U84 ( .A(n19583), .B(n19582), .Z(n19584) );
  XOR U85 ( .A(n19631), .B(n19630), .Z(n19633) );
  XNOR U86 ( .A(n18992), .B(n18991), .Z(n19001) );
  XNOR U87 ( .A(n18977), .B(n18976), .Z(n18947) );
  XNOR U88 ( .A(n19069), .B(n19068), .Z(n19078) );
  XOR U89 ( .A(n19160), .B(n19159), .Z(n19108) );
  XOR U90 ( .A(n19544), .B(n19543), .Z(n19559) );
  XOR U91 ( .A(n19625), .B(n19624), .Z(n19626) );
  XOR U92 ( .A(n19235), .B(n19234), .Z(n19236) );
  XOR U93 ( .A(n19304), .B(n19303), .Z(n19305) );
  XNOR U94 ( .A(n19370), .B(n19369), .Z(n19373) );
  XOR U95 ( .A(n19388), .B(n19387), .Z(n19390) );
  XNOR U96 ( .A(n19464), .B(n19463), .Z(n19455) );
  XOR U97 ( .A(n19514), .B(n19513), .Z(n19515) );
  NAND U98 ( .A(n19580), .B(n19581), .Z(n13) );
  XOR U99 ( .A(n19580), .B(n19581), .Z(n14) );
  NANDN U100 ( .A(n19579), .B(n14), .Z(n15) );
  NAND U101 ( .A(n13), .B(n15), .Z(n19621) );
  XOR U102 ( .A(n19671), .B(n19670), .Z(n19672) );
  XOR U103 ( .A(n19739), .B(n19738), .Z(n19740) );
  XOR U104 ( .A(n19753), .B(n19752), .Z(n19754) );
  XOR U105 ( .A(n19787), .B(n19786), .Z(n19788) );
  XOR U106 ( .A(n19101), .B(n19100), .Z(n19102) );
  XOR U107 ( .A(n19576), .B(n19575), .Z(n19567) );
  XOR U108 ( .A(n19831), .B(n19830), .Z(n19832) );
  XOR U109 ( .A(n19856), .B(n19855), .Z(n19858) );
  NAND U110 ( .A(b[0]), .B(a[234]), .Z(n16) );
  XNOR U111 ( .A(b[1]), .B(n16), .Z(n17) );
  NANDN U112 ( .A(b[0]), .B(a[233]), .Z(n18) );
  AND U113 ( .A(n17), .B(n18), .Z(n17496) );
  XOR U114 ( .A(n18954), .B(n18953), .Z(n18955) );
  XOR U115 ( .A(n19031), .B(n19030), .Z(n19032) );
  XOR U116 ( .A(n19113), .B(n19112), .Z(n19114) );
  XOR U117 ( .A(n18998), .B(n18997), .Z(n18974) );
  XOR U118 ( .A(n19075), .B(n19074), .Z(n19051) );
  XOR U119 ( .A(n19154), .B(n19153), .Z(n19130) );
  XOR U120 ( .A(n19199), .B(n19198), .Z(n19200) );
  XOR U121 ( .A(n19207), .B(n19206), .Z(n19223) );
  XOR U122 ( .A(n19288), .B(n19287), .Z(n19292) );
  XOR U123 ( .A(n19350), .B(n19349), .Z(n19351) );
  XOR U124 ( .A(n19400), .B(n19399), .Z(n19401) );
  XNOR U125 ( .A(n19504), .B(n19503), .Z(n19475) );
  NANDN U126 ( .A(n612), .B(n613), .Z(n19) );
  NANDN U127 ( .A(n611), .B(n610), .Z(n20) );
  NAND U128 ( .A(n19), .B(n20), .Z(n636) );
  XOR U129 ( .A(n19004), .B(n19003), .Z(n18949) );
  NAND U130 ( .A(n18877), .B(n18876), .Z(n21) );
  NANDN U131 ( .A(n18874), .B(n18875), .Z(n22) );
  AND U132 ( .A(n21), .B(n22), .Z(n19010) );
  XOR U133 ( .A(n19081), .B(n19080), .Z(n19026) );
  XNOR U134 ( .A(n19148), .B(n19147), .Z(n19157) );
  XNOR U135 ( .A(n19195), .B(n19194), .Z(n19228) );
  XNOR U136 ( .A(n19278), .B(n19277), .Z(n19297) );
  XOR U137 ( .A(n19318), .B(n19317), .Z(n19319) );
  XOR U138 ( .A(n19442), .B(n19441), .Z(n19443) );
  XOR U139 ( .A(n19394), .B(n19393), .Z(n19396) );
  XOR U140 ( .A(n19468), .B(n19467), .Z(n19469) );
  XNOR U141 ( .A(n19562), .B(n19561), .Z(n19519) );
  XNOR U142 ( .A(n19585), .B(n19584), .Z(n19605) );
  XOR U143 ( .A(n19657), .B(n19656), .Z(n19658) );
  XOR U144 ( .A(n19683), .B(n19682), .Z(n19684) );
  XOR U145 ( .A(n19716), .B(n19715), .Z(n19718) );
  XNOR U146 ( .A(n19755), .B(n19754), .Z(n19746) );
  NAND U147 ( .A(n73), .B(n74), .Z(n23) );
  XOR U148 ( .A(n73), .B(n74), .Z(n24) );
  NANDN U149 ( .A(n72), .B(n24), .Z(n25) );
  NAND U150 ( .A(n23), .B(n25), .Z(n86) );
  XOR U151 ( .A(n19172), .B(n19171), .Z(n19173) );
  XOR U152 ( .A(n19103), .B(n19102), .Z(n19095) );
  XOR U153 ( .A(n19243), .B(n19242), .Z(n19244) );
  XOR U154 ( .A(n19312), .B(n19311), .Z(n19313) );
  XOR U155 ( .A(n19382), .B(n19381), .Z(n19383) );
  XOR U156 ( .A(n19508), .B(n19507), .Z(n19509) );
  XOR U157 ( .A(n19568), .B(n19567), .Z(n19569) );
  XOR U158 ( .A(n19613), .B(n19612), .Z(n19614) );
  XOR U159 ( .A(n19665), .B(n19664), .Z(n19666) );
  XOR U160 ( .A(n19704), .B(n19703), .Z(n19705) );
  XOR U161 ( .A(n19816), .B(n19815), .Z(n19817) );
  XOR U162 ( .A(n19863), .B(n19864), .Z(n19866) );
  NAND U163 ( .A(n202), .B(n415), .Z(n26) );
  NAND U164 ( .A(n123), .B(n463), .Z(n27) );
  NAND U165 ( .A(n296), .B(n678), .Z(n28) );
  NAND U166 ( .A(n75), .B(n30), .Z(n29) );
  XNOR U167 ( .A(b[1]), .B(b[2]), .Z(n30) );
  IV U168 ( .A(n29), .Z(n31) );
  IV U169 ( .A(n30), .Z(n32) );
  IV U170 ( .A(n27), .Z(n33) );
  IV U171 ( .A(n26), .Z(n34) );
  IV U172 ( .A(n28), .Z(n35) );
  AND U173 ( .A(b[0]), .B(a[0]), .Z(n37) );
  XOR U174 ( .A(n37), .B(sreg[240]), .Z(c[240]) );
  AND U175 ( .A(b[0]), .B(a[1]), .Z(n44) );
  NAND U176 ( .A(a[0]), .B(b[1]), .Z(n36) );
  XOR U177 ( .A(n44), .B(n36), .Z(n38) );
  XNOR U178 ( .A(sreg[241]), .B(n38), .Z(n40) );
  AND U179 ( .A(n37), .B(sreg[240]), .Z(n39) );
  XOR U180 ( .A(n40), .B(n39), .Z(c[241]) );
  NANDN U181 ( .A(n38), .B(sreg[241]), .Z(n42) );
  NAND U182 ( .A(n40), .B(n39), .Z(n41) );
  AND U183 ( .A(n42), .B(n41), .Z(n62) );
  XNOR U184 ( .A(n62), .B(sreg[242]), .Z(n64) );
  NAND U185 ( .A(a[0]), .B(b[2]), .Z(n43) );
  XNOR U186 ( .A(b[1]), .B(n43), .Z(n46) );
  NANDN U187 ( .A(a[0]), .B(n44), .Z(n45) );
  NAND U188 ( .A(n46), .B(n45), .Z(n51) );
  NAND U189 ( .A(b[0]), .B(a[2]), .Z(n47) );
  XNOR U190 ( .A(b[1]), .B(n47), .Z(n49) );
  NANDN U191 ( .A(b[0]), .B(a[1]), .Z(n48) );
  NAND U192 ( .A(n49), .B(n48), .Z(n50) );
  XOR U193 ( .A(n51), .B(n50), .Z(n63) );
  XOR U194 ( .A(n64), .B(n63), .Z(c[242]) );
  NOR U195 ( .A(n51), .B(n50), .Z(n74) );
  NAND U196 ( .A(n32), .B(a[0]), .Z(n53) );
  NAND U197 ( .A(b[1]), .B(b[2]), .Z(n52) );
  NAND U198 ( .A(b[3]), .B(n52), .Z(n19406) );
  IV U199 ( .A(n19406), .Z(n19348) );
  AND U200 ( .A(n53), .B(n19348), .Z(n73) );
  NAND U201 ( .A(b[0]), .B(a[3]), .Z(n54) );
  XNOR U202 ( .A(b[1]), .B(n54), .Z(n56) );
  NANDN U203 ( .A(b[0]), .B(a[2]), .Z(n55) );
  NAND U204 ( .A(n56), .B(n55), .Z(n83) );
  XOR U205 ( .A(b[3]), .B(b[2]), .Z(n75) );
  XOR U206 ( .A(b[3]), .B(a[0]), .Z(n57) );
  NAND U207 ( .A(n75), .B(n57), .Z(n58) );
  NANDN U208 ( .A(n58), .B(n30), .Z(n60) );
  XOR U209 ( .A(b[3]), .B(a[1]), .Z(n76) );
  NANDN U210 ( .A(n30), .B(n76), .Z(n59) );
  NAND U211 ( .A(n60), .B(n59), .Z(n82) );
  XOR U212 ( .A(n83), .B(n82), .Z(n72) );
  XOR U213 ( .A(n73), .B(n72), .Z(n61) );
  XOR U214 ( .A(n74), .B(n61), .Z(n67) );
  XNOR U215 ( .A(sreg[243]), .B(n67), .Z(n69) );
  NANDN U216 ( .A(n62), .B(sreg[242]), .Z(n66) );
  NAND U217 ( .A(n64), .B(n63), .Z(n65) );
  NAND U218 ( .A(n66), .B(n65), .Z(n68) );
  XOR U219 ( .A(n69), .B(n68), .Z(c[243]) );
  NANDN U220 ( .A(n67), .B(sreg[243]), .Z(n71) );
  NAND U221 ( .A(n69), .B(n68), .Z(n70) );
  AND U222 ( .A(n71), .B(n70), .Z(n107) );
  XNOR U223 ( .A(n107), .B(sreg[244]), .Z(n109) );
  NAND U224 ( .A(n31), .B(n76), .Z(n78) );
  XOR U225 ( .A(b[3]), .B(a[2]), .Z(n90) );
  NAND U226 ( .A(n32), .B(n90), .Z(n77) );
  AND U227 ( .A(n78), .B(n77), .Z(n104) );
  XNOR U228 ( .A(b[3]), .B(b[4]), .Z(n463) );
  IV U229 ( .A(n463), .Z(n19342) );
  AND U230 ( .A(a[0]), .B(n19342), .Z(n101) );
  NAND U231 ( .A(b[0]), .B(a[4]), .Z(n79) );
  XNOR U232 ( .A(b[1]), .B(n79), .Z(n81) );
  NANDN U233 ( .A(b[0]), .B(a[3]), .Z(n80) );
  NAND U234 ( .A(n81), .B(n80), .Z(n102) );
  XNOR U235 ( .A(n101), .B(n102), .Z(n103) );
  XNOR U236 ( .A(n104), .B(n103), .Z(n84) );
  NANDN U237 ( .A(n83), .B(n82), .Z(n85) );
  XOR U238 ( .A(n84), .B(n85), .Z(n87) );
  XNOR U239 ( .A(n86), .B(n87), .Z(n108) );
  XOR U240 ( .A(n109), .B(n108), .Z(c[244]) );
  NANDN U241 ( .A(n85), .B(n84), .Z(n89) );
  NANDN U242 ( .A(n87), .B(n86), .Z(n88) );
  AND U243 ( .A(n89), .B(n88), .Z(n120) );
  NAND U244 ( .A(n31), .B(n90), .Z(n92) );
  XOR U245 ( .A(b[3]), .B(a[3]), .Z(n129) );
  NAND U246 ( .A(n32), .B(n129), .Z(n91) );
  AND U247 ( .A(n92), .B(n91), .Z(n136) );
  NAND U248 ( .A(b[3]), .B(b[4]), .Z(n93) );
  AND U249 ( .A(b[5]), .B(n93), .Z(n19492) );
  IV U250 ( .A(n19492), .Z(n19553) );
  NOR U251 ( .A(n19553), .B(n101), .Z(n135) );
  XNOR U252 ( .A(n136), .B(n135), .Z(n138) );
  NAND U253 ( .A(b[0]), .B(a[5]), .Z(n94) );
  XNOR U254 ( .A(b[1]), .B(n94), .Z(n96) );
  NANDN U255 ( .A(b[0]), .B(a[4]), .Z(n95) );
  NAND U256 ( .A(n96), .B(n95), .Z(n127) );
  XOR U257 ( .A(b[5]), .B(b[4]), .Z(n123) );
  XOR U258 ( .A(b[5]), .B(a[0]), .Z(n97) );
  NAND U259 ( .A(n123), .B(n97), .Z(n98) );
  NANDN U260 ( .A(n98), .B(n463), .Z(n100) );
  XOR U261 ( .A(b[5]), .B(a[1]), .Z(n124) );
  NANDN U262 ( .A(n463), .B(n124), .Z(n99) );
  NAND U263 ( .A(n100), .B(n99), .Z(n128) );
  XNOR U264 ( .A(n127), .B(n128), .Z(n137) );
  XOR U265 ( .A(n138), .B(n137), .Z(n118) );
  NANDN U266 ( .A(n102), .B(n101), .Z(n106) );
  NANDN U267 ( .A(n104), .B(n103), .Z(n105) );
  AND U268 ( .A(n106), .B(n105), .Z(n117) );
  XNOR U269 ( .A(n118), .B(n117), .Z(n119) );
  XOR U270 ( .A(n120), .B(n119), .Z(n112) );
  XNOR U271 ( .A(n112), .B(sreg[245]), .Z(n114) );
  NANDN U272 ( .A(n107), .B(sreg[244]), .Z(n111) );
  NAND U273 ( .A(n109), .B(n108), .Z(n110) );
  NAND U274 ( .A(n111), .B(n110), .Z(n113) );
  XOR U275 ( .A(n114), .B(n113), .Z(c[245]) );
  NANDN U276 ( .A(n112), .B(sreg[245]), .Z(n116) );
  NAND U277 ( .A(n114), .B(n113), .Z(n115) );
  AND U278 ( .A(n116), .B(n115), .Z(n174) );
  XNOR U279 ( .A(n174), .B(sreg[246]), .Z(n176) );
  NANDN U280 ( .A(n118), .B(n117), .Z(n122) );
  NAND U281 ( .A(n120), .B(n119), .Z(n121) );
  AND U282 ( .A(n122), .B(n121), .Z(n143) );
  NAND U283 ( .A(n33), .B(n124), .Z(n126) );
  XOR U284 ( .A(b[5]), .B(a[2]), .Z(n152) );
  NAND U285 ( .A(n19342), .B(n152), .Z(n125) );
  AND U286 ( .A(n126), .B(n125), .Z(n169) );
  ANDN U287 ( .B(n128), .A(n127), .Z(n168) );
  XNOR U288 ( .A(n169), .B(n168), .Z(n171) );
  NAND U289 ( .A(n31), .B(n129), .Z(n131) );
  XOR U290 ( .A(b[3]), .B(a[4]), .Z(n159) );
  NAND U291 ( .A(n32), .B(n159), .Z(n130) );
  AND U292 ( .A(n131), .B(n130), .Z(n165) );
  XNOR U293 ( .A(b[5]), .B(b[6]), .Z(n415) );
  IV U294 ( .A(n415), .Z(n19486) );
  AND U295 ( .A(a[0]), .B(n19486), .Z(n162) );
  NAND U296 ( .A(b[0]), .B(a[6]), .Z(n132) );
  XNOR U297 ( .A(b[1]), .B(n132), .Z(n134) );
  NANDN U298 ( .A(b[0]), .B(a[5]), .Z(n133) );
  NAND U299 ( .A(n134), .B(n133), .Z(n163) );
  XNOR U300 ( .A(n162), .B(n163), .Z(n164) );
  XNOR U301 ( .A(n165), .B(n164), .Z(n170) );
  XOR U302 ( .A(n171), .B(n170), .Z(n142) );
  NANDN U303 ( .A(n136), .B(n135), .Z(n140) );
  NAND U304 ( .A(n138), .B(n137), .Z(n139) );
  AND U305 ( .A(n140), .B(n139), .Z(n141) );
  XOR U306 ( .A(n142), .B(n141), .Z(n144) );
  XNOR U307 ( .A(n143), .B(n144), .Z(n175) );
  XOR U308 ( .A(n176), .B(n175), .Z(c[246]) );
  NANDN U309 ( .A(n142), .B(n141), .Z(n146) );
  OR U310 ( .A(n144), .B(n143), .Z(n145) );
  AND U311 ( .A(n146), .B(n145), .Z(n186) );
  XOR U312 ( .A(b[7]), .B(a[0]), .Z(n149) );
  XOR U313 ( .A(b[7]), .B(b[5]), .Z(n147) );
  XOR U314 ( .A(b[7]), .B(b[6]), .Z(n202) );
  AND U315 ( .A(n147), .B(n202), .Z(n148) );
  NAND U316 ( .A(n149), .B(n148), .Z(n151) );
  XNOR U317 ( .A(b[7]), .B(a[1]), .Z(n203) );
  OR U318 ( .A(n203), .B(n415), .Z(n150) );
  AND U319 ( .A(n151), .B(n150), .Z(n209) );
  NAND U320 ( .A(n33), .B(n152), .Z(n154) );
  XOR U321 ( .A(b[5]), .B(a[3]), .Z(n214) );
  NAND U322 ( .A(n19342), .B(n214), .Z(n153) );
  AND U323 ( .A(n154), .B(n153), .Z(n210) );
  XOR U324 ( .A(n209), .B(n210), .Z(n199) );
  NAND U325 ( .A(b[5]), .B(b[6]), .Z(n155) );
  NAND U326 ( .A(b[7]), .B(n155), .Z(n19646) );
  NOR U327 ( .A(n19646), .B(n162), .Z(n197) );
  NAND U328 ( .A(b[0]), .B(a[7]), .Z(n156) );
  XNOR U329 ( .A(b[1]), .B(n156), .Z(n158) );
  NANDN U330 ( .A(b[0]), .B(a[6]), .Z(n157) );
  NAND U331 ( .A(n158), .B(n157), .Z(n196) );
  XNOR U332 ( .A(n197), .B(n196), .Z(n198) );
  XNOR U333 ( .A(n199), .B(n198), .Z(n190) );
  NANDN U334 ( .A(n29), .B(n159), .Z(n161) );
  XNOR U335 ( .A(b[3]), .B(a[5]), .Z(n206) );
  OR U336 ( .A(n206), .B(n30), .Z(n160) );
  NAND U337 ( .A(n161), .B(n160), .Z(n191) );
  XNOR U338 ( .A(n190), .B(n191), .Z(n192) );
  NANDN U339 ( .A(n163), .B(n162), .Z(n167) );
  NANDN U340 ( .A(n165), .B(n164), .Z(n166) );
  NAND U341 ( .A(n167), .B(n166), .Z(n193) );
  XNOR U342 ( .A(n192), .B(n193), .Z(n184) );
  NANDN U343 ( .A(n169), .B(n168), .Z(n173) );
  NAND U344 ( .A(n171), .B(n170), .Z(n172) );
  NAND U345 ( .A(n173), .B(n172), .Z(n185) );
  XOR U346 ( .A(n184), .B(n185), .Z(n187) );
  XOR U347 ( .A(n186), .B(n187), .Z(n179) );
  XNOR U348 ( .A(n179), .B(sreg[247]), .Z(n181) );
  NANDN U349 ( .A(n174), .B(sreg[246]), .Z(n178) );
  NAND U350 ( .A(n176), .B(n175), .Z(n177) );
  NAND U351 ( .A(n178), .B(n177), .Z(n180) );
  XOR U352 ( .A(n181), .B(n180), .Z(c[247]) );
  NANDN U353 ( .A(n179), .B(sreg[247]), .Z(n183) );
  NAND U354 ( .A(n181), .B(n180), .Z(n182) );
  AND U355 ( .A(n183), .B(n182), .Z(n259) );
  XNOR U356 ( .A(n259), .B(sreg[248]), .Z(n261) );
  NANDN U357 ( .A(n185), .B(n184), .Z(n189) );
  OR U358 ( .A(n187), .B(n186), .Z(n188) );
  AND U359 ( .A(n189), .B(n188), .Z(n255) );
  NANDN U360 ( .A(n191), .B(n190), .Z(n195) );
  NANDN U361 ( .A(n193), .B(n192), .Z(n194) );
  AND U362 ( .A(n195), .B(n194), .Z(n254) );
  NANDN U363 ( .A(n197), .B(n196), .Z(n201) );
  NANDN U364 ( .A(n199), .B(n198), .Z(n200) );
  AND U365 ( .A(n201), .B(n200), .Z(n220) );
  OR U366 ( .A(n203), .B(n26), .Z(n205) );
  XOR U367 ( .A(b[7]), .B(a[2]), .Z(n239) );
  NAND U368 ( .A(n19486), .B(n239), .Z(n204) );
  AND U369 ( .A(n205), .B(n204), .Z(n224) );
  OR U370 ( .A(n206), .B(n29), .Z(n208) );
  XOR U371 ( .A(b[3]), .B(a[6]), .Z(n250) );
  NAND U372 ( .A(n32), .B(n250), .Z(n207) );
  NAND U373 ( .A(n208), .B(n207), .Z(n223) );
  XNOR U374 ( .A(n224), .B(n223), .Z(n226) );
  NOR U375 ( .A(n210), .B(n209), .Z(n225) );
  XOR U376 ( .A(n226), .B(n225), .Z(n218) );
  NAND U377 ( .A(b[0]), .B(a[8]), .Z(n211) );
  XNOR U378 ( .A(b[1]), .B(n211), .Z(n213) );
  NANDN U379 ( .A(b[0]), .B(a[7]), .Z(n212) );
  NAND U380 ( .A(n213), .B(n212), .Z(n231) );
  XNOR U381 ( .A(b[7]), .B(b[8]), .Z(n678) );
  IV U382 ( .A(n678), .Z(n19598) );
  AND U383 ( .A(a[0]), .B(n19598), .Z(n243) );
  NAND U384 ( .A(n33), .B(n214), .Z(n216) );
  XOR U385 ( .A(b[5]), .B(a[4]), .Z(n244) );
  NAND U386 ( .A(n19342), .B(n244), .Z(n215) );
  AND U387 ( .A(n216), .B(n215), .Z(n229) );
  XOR U388 ( .A(n243), .B(n229), .Z(n230) );
  XNOR U389 ( .A(n231), .B(n230), .Z(n217) );
  XNOR U390 ( .A(n218), .B(n217), .Z(n219) );
  XNOR U391 ( .A(n220), .B(n219), .Z(n253) );
  XOR U392 ( .A(n254), .B(n253), .Z(n256) );
  XNOR U393 ( .A(n255), .B(n256), .Z(n260) );
  XOR U394 ( .A(n261), .B(n260), .Z(c[248]) );
  NANDN U395 ( .A(n218), .B(n217), .Z(n222) );
  NANDN U396 ( .A(n220), .B(n219), .Z(n221) );
  AND U397 ( .A(n222), .B(n221), .Z(n269) );
  NANDN U398 ( .A(n224), .B(n223), .Z(n228) );
  NAND U399 ( .A(n226), .B(n225), .Z(n227) );
  AND U400 ( .A(n228), .B(n227), .Z(n308) );
  NANDN U401 ( .A(n229), .B(n243), .Z(n233) );
  OR U402 ( .A(n231), .B(n230), .Z(n232) );
  AND U403 ( .A(n233), .B(n232), .Z(n306) );
  XOR U404 ( .A(b[9]), .B(a[0]), .Z(n236) );
  XOR U405 ( .A(b[9]), .B(b[7]), .Z(n234) );
  XOR U406 ( .A(b[9]), .B(b[8]), .Z(n296) );
  AND U407 ( .A(n234), .B(n296), .Z(n235) );
  NAND U408 ( .A(n236), .B(n235), .Z(n238) );
  XNOR U409 ( .A(b[9]), .B(a[1]), .Z(n297) );
  OR U410 ( .A(n297), .B(n678), .Z(n237) );
  AND U411 ( .A(n238), .B(n237), .Z(n300) );
  NAND U412 ( .A(n34), .B(n239), .Z(n241) );
  XOR U413 ( .A(b[7]), .B(a[3]), .Z(n290) );
  NAND U414 ( .A(n19486), .B(n290), .Z(n240) );
  NAND U415 ( .A(n241), .B(n240), .Z(n301) );
  XOR U416 ( .A(n300), .B(n301), .Z(n277) );
  NAND U417 ( .A(b[7]), .B(b[8]), .Z(n242) );
  NAND U418 ( .A(b[9]), .B(n242), .Z(n19734) );
  NOR U419 ( .A(n19734), .B(n243), .Z(n276) );
  NAND U420 ( .A(n33), .B(n244), .Z(n246) );
  XOR U421 ( .A(b[5]), .B(a[5]), .Z(n293) );
  NAND U422 ( .A(n19342), .B(n293), .Z(n245) );
  AND U423 ( .A(n246), .B(n245), .Z(n275) );
  XOR U424 ( .A(n276), .B(n275), .Z(n278) );
  XOR U425 ( .A(n277), .B(n278), .Z(n284) );
  NAND U426 ( .A(b[0]), .B(a[9]), .Z(n247) );
  XNOR U427 ( .A(b[1]), .B(n247), .Z(n249) );
  NANDN U428 ( .A(b[0]), .B(a[8]), .Z(n248) );
  NAND U429 ( .A(n249), .B(n248), .Z(n282) );
  NAND U430 ( .A(n31), .B(n250), .Z(n252) );
  XOR U431 ( .A(b[3]), .B(a[7]), .Z(n302) );
  NAND U432 ( .A(n32), .B(n302), .Z(n251) );
  NAND U433 ( .A(n252), .B(n251), .Z(n281) );
  XNOR U434 ( .A(n282), .B(n281), .Z(n283) );
  XOR U435 ( .A(n284), .B(n283), .Z(n305) );
  XNOR U436 ( .A(n306), .B(n305), .Z(n307) );
  XOR U437 ( .A(n308), .B(n307), .Z(n270) );
  XNOR U438 ( .A(n269), .B(n270), .Z(n271) );
  NANDN U439 ( .A(n254), .B(n253), .Z(n258) );
  OR U440 ( .A(n256), .B(n255), .Z(n257) );
  NAND U441 ( .A(n258), .B(n257), .Z(n272) );
  XOR U442 ( .A(n271), .B(n272), .Z(n264) );
  XNOR U443 ( .A(sreg[249]), .B(n264), .Z(n266) );
  NANDN U444 ( .A(n259), .B(sreg[248]), .Z(n263) );
  NAND U445 ( .A(n261), .B(n260), .Z(n262) );
  NAND U446 ( .A(n263), .B(n262), .Z(n265) );
  XOR U447 ( .A(n266), .B(n265), .Z(c[249]) );
  NANDN U448 ( .A(n264), .B(sreg[249]), .Z(n268) );
  NAND U449 ( .A(n266), .B(n265), .Z(n267) );
  AND U450 ( .A(n268), .B(n267), .Z(n311) );
  XNOR U451 ( .A(n311), .B(sreg[250]), .Z(n313) );
  NANDN U452 ( .A(n270), .B(n269), .Z(n274) );
  NANDN U453 ( .A(n272), .B(n271), .Z(n273) );
  AND U454 ( .A(n274), .B(n273), .Z(n319) );
  NANDN U455 ( .A(n276), .B(n275), .Z(n280) );
  NANDN U456 ( .A(n278), .B(n277), .Z(n279) );
  AND U457 ( .A(n280), .B(n279), .Z(n361) );
  NANDN U458 ( .A(n282), .B(n281), .Z(n286) );
  NAND U459 ( .A(n284), .B(n283), .Z(n285) );
  AND U460 ( .A(n286), .B(n285), .Z(n360) );
  XNOR U461 ( .A(n361), .B(n360), .Z(n362) );
  NAND U462 ( .A(b[0]), .B(a[10]), .Z(n287) );
  XNOR U463 ( .A(b[1]), .B(n287), .Z(n289) );
  NANDN U464 ( .A(b[0]), .B(a[9]), .Z(n288) );
  NAND U465 ( .A(n289), .B(n288), .Z(n330) );
  XNOR U466 ( .A(b[9]), .B(b[10]), .Z(n401) );
  IV U467 ( .A(n401), .Z(n19692) );
  AND U468 ( .A(a[0]), .B(n19692), .Z(n353) );
  NAND U469 ( .A(n34), .B(n290), .Z(n292) );
  XOR U470 ( .A(b[7]), .B(a[4]), .Z(n354) );
  NAND U471 ( .A(n19486), .B(n354), .Z(n291) );
  AND U472 ( .A(n292), .B(n291), .Z(n328) );
  XOR U473 ( .A(n353), .B(n328), .Z(n329) );
  XOR U474 ( .A(n330), .B(n329), .Z(n325) );
  NAND U475 ( .A(n33), .B(n293), .Z(n295) );
  XOR U476 ( .A(b[5]), .B(a[6]), .Z(n349) );
  NAND U477 ( .A(n19342), .B(n349), .Z(n294) );
  AND U478 ( .A(n295), .B(n294), .Z(n334) );
  OR U479 ( .A(n297), .B(n28), .Z(n299) );
  XOR U480 ( .A(b[9]), .B(a[2]), .Z(n339) );
  NAND U481 ( .A(n19598), .B(n339), .Z(n298) );
  NAND U482 ( .A(n299), .B(n298), .Z(n333) );
  XNOR U483 ( .A(n334), .B(n333), .Z(n336) );
  ANDN U484 ( .B(n301), .A(n300), .Z(n335) );
  XOR U485 ( .A(n336), .B(n335), .Z(n323) );
  NANDN U486 ( .A(n29), .B(n302), .Z(n304) );
  XNOR U487 ( .A(b[3]), .B(a[8]), .Z(n357) );
  OR U488 ( .A(n357), .B(n30), .Z(n303) );
  AND U489 ( .A(n304), .B(n303), .Z(n322) );
  XNOR U490 ( .A(n323), .B(n322), .Z(n324) );
  XOR U491 ( .A(n325), .B(n324), .Z(n363) );
  XNOR U492 ( .A(n362), .B(n363), .Z(n316) );
  NANDN U493 ( .A(n306), .B(n305), .Z(n310) );
  NANDN U494 ( .A(n308), .B(n307), .Z(n309) );
  NAND U495 ( .A(n310), .B(n309), .Z(n317) );
  XNOR U496 ( .A(n316), .B(n317), .Z(n318) );
  XNOR U497 ( .A(n319), .B(n318), .Z(n312) );
  XOR U498 ( .A(n313), .B(n312), .Z(c[250]) );
  NANDN U499 ( .A(n311), .B(sreg[250]), .Z(n315) );
  NAND U500 ( .A(n313), .B(n312), .Z(n314) );
  AND U501 ( .A(n315), .B(n314), .Z(n368) );
  NANDN U502 ( .A(n317), .B(n316), .Z(n321) );
  NAND U503 ( .A(n319), .B(n318), .Z(n320) );
  AND U504 ( .A(n321), .B(n320), .Z(n374) );
  NANDN U505 ( .A(n323), .B(n322), .Z(n327) );
  NANDN U506 ( .A(n325), .B(n324), .Z(n326) );
  AND U507 ( .A(n327), .B(n326), .Z(n421) );
  NANDN U508 ( .A(n328), .B(n353), .Z(n332) );
  OR U509 ( .A(n330), .B(n329), .Z(n331) );
  AND U510 ( .A(n332), .B(n331), .Z(n419) );
  NANDN U511 ( .A(n334), .B(n333), .Z(n338) );
  NAND U512 ( .A(n336), .B(n335), .Z(n337) );
  AND U513 ( .A(n338), .B(n337), .Z(n380) );
  NAND U514 ( .A(n35), .B(n339), .Z(n341) );
  XOR U515 ( .A(b[9]), .B(a[3]), .Z(n392) );
  NAND U516 ( .A(n19598), .B(n392), .Z(n340) );
  AND U517 ( .A(n341), .B(n340), .Z(n409) );
  XOR U518 ( .A(b[11]), .B(b[10]), .Z(n402) );
  XOR U519 ( .A(b[11]), .B(a[0]), .Z(n342) );
  NAND U520 ( .A(n402), .B(n342), .Z(n343) );
  NANDN U521 ( .A(n343), .B(n401), .Z(n345) );
  XOR U522 ( .A(b[11]), .B(a[1]), .Z(n403) );
  NANDN U523 ( .A(n401), .B(n403), .Z(n344) );
  AND U524 ( .A(n345), .B(n344), .Z(n410) );
  XOR U525 ( .A(n409), .B(n410), .Z(n397) );
  NAND U526 ( .A(b[0]), .B(a[11]), .Z(n346) );
  XNOR U527 ( .A(b[1]), .B(n346), .Z(n348) );
  NANDN U528 ( .A(b[0]), .B(a[10]), .Z(n347) );
  NAND U529 ( .A(n348), .B(n347), .Z(n395) );
  NANDN U530 ( .A(n27), .B(n349), .Z(n351) );
  XNOR U531 ( .A(b[5]), .B(a[7]), .Z(n406) );
  OR U532 ( .A(n406), .B(n463), .Z(n350) );
  NAND U533 ( .A(n351), .B(n350), .Z(n396) );
  XOR U534 ( .A(n395), .B(n396), .Z(n398) );
  XOR U535 ( .A(n397), .B(n398), .Z(n378) );
  NAND U536 ( .A(b[9]), .B(b[10]), .Z(n352) );
  AND U537 ( .A(b[11]), .B(n352), .Z(n19771) );
  IV U538 ( .A(n19771), .Z(n19801) );
  NOR U539 ( .A(n19801), .B(n353), .Z(n384) );
  NANDN U540 ( .A(n26), .B(n354), .Z(n356) );
  XNOR U541 ( .A(b[7]), .B(a[5]), .Z(n414) );
  OR U542 ( .A(n414), .B(n415), .Z(n355) );
  NAND U543 ( .A(n356), .B(n355), .Z(n383) );
  XOR U544 ( .A(n384), .B(n383), .Z(n386) );
  OR U545 ( .A(n357), .B(n29), .Z(n359) );
  XNOR U546 ( .A(b[3]), .B(a[9]), .Z(n411) );
  OR U547 ( .A(n411), .B(n30), .Z(n358) );
  NAND U548 ( .A(n359), .B(n358), .Z(n385) );
  XOR U549 ( .A(n386), .B(n385), .Z(n377) );
  XNOR U550 ( .A(n378), .B(n377), .Z(n379) );
  XNOR U551 ( .A(n380), .B(n379), .Z(n418) );
  XNOR U552 ( .A(n419), .B(n418), .Z(n420) );
  XOR U553 ( .A(n421), .B(n420), .Z(n372) );
  NANDN U554 ( .A(n361), .B(n360), .Z(n365) );
  NANDN U555 ( .A(n363), .B(n362), .Z(n364) );
  NAND U556 ( .A(n365), .B(n364), .Z(n371) );
  XNOR U557 ( .A(n372), .B(n371), .Z(n373) );
  XNOR U558 ( .A(n374), .B(n373), .Z(n366) );
  XNOR U559 ( .A(sreg[251]), .B(n366), .Z(n367) );
  XNOR U560 ( .A(n368), .B(n367), .Z(c[251]) );
  NANDN U561 ( .A(sreg[251]), .B(n366), .Z(n370) );
  NAND U562 ( .A(n368), .B(n367), .Z(n369) );
  NAND U563 ( .A(n370), .B(n369), .Z(n484) );
  XNOR U564 ( .A(sreg[252]), .B(n484), .Z(n486) );
  NANDN U565 ( .A(n372), .B(n371), .Z(n376) );
  NANDN U566 ( .A(n374), .B(n373), .Z(n375) );
  AND U567 ( .A(n376), .B(n375), .Z(n427) );
  NANDN U568 ( .A(n378), .B(n377), .Z(n382) );
  NANDN U569 ( .A(n380), .B(n379), .Z(n381) );
  AND U570 ( .A(n382), .B(n381), .Z(n479) );
  NAND U571 ( .A(n384), .B(n383), .Z(n388) );
  NAND U572 ( .A(n386), .B(n385), .Z(n387) );
  NAND U573 ( .A(n388), .B(n387), .Z(n478) );
  XNOR U574 ( .A(n479), .B(n478), .Z(n481) );
  NAND U575 ( .A(b[0]), .B(a[12]), .Z(n389) );
  XNOR U576 ( .A(b[1]), .B(n389), .Z(n391) );
  NANDN U577 ( .A(b[0]), .B(a[11]), .Z(n390) );
  NAND U578 ( .A(n391), .B(n390), .Z(n469) );
  XNOR U579 ( .A(b[11]), .B(b[12]), .Z(n19434) );
  IV U580 ( .A(n19434), .Z(n19768) );
  AND U581 ( .A(a[0]), .B(n19768), .Z(n466) );
  NAND U582 ( .A(n35), .B(n392), .Z(n394) );
  XOR U583 ( .A(b[9]), .B(a[4]), .Z(n458) );
  NAND U584 ( .A(n19598), .B(n458), .Z(n393) );
  AND U585 ( .A(n394), .B(n393), .Z(n467) );
  XNOR U586 ( .A(n466), .B(n467), .Z(n468) );
  XNOR U587 ( .A(n469), .B(n468), .Z(n430) );
  NANDN U588 ( .A(n396), .B(n395), .Z(n400) );
  OR U589 ( .A(n398), .B(n397), .Z(n399) );
  NAND U590 ( .A(n400), .B(n399), .Z(n431) );
  XNOR U591 ( .A(n430), .B(n431), .Z(n432) );
  AND U592 ( .A(n402), .B(n401), .Z(n19724) );
  NAND U593 ( .A(n403), .B(n19724), .Z(n405) );
  XOR U594 ( .A(b[11]), .B(a[2]), .Z(n448) );
  NAND U595 ( .A(n19692), .B(n448), .Z(n404) );
  AND U596 ( .A(n405), .B(n404), .Z(n439) );
  OR U597 ( .A(n406), .B(n27), .Z(n408) );
  XOR U598 ( .A(b[5]), .B(a[8]), .Z(n462) );
  NAND U599 ( .A(n19342), .B(n462), .Z(n407) );
  AND U600 ( .A(n408), .B(n407), .Z(n437) );
  NOR U601 ( .A(n410), .B(n409), .Z(n474) );
  OR U602 ( .A(n411), .B(n29), .Z(n413) );
  XNOR U603 ( .A(b[3]), .B(a[10]), .Z(n455) );
  OR U604 ( .A(n455), .B(n30), .Z(n412) );
  AND U605 ( .A(n413), .B(n412), .Z(n472) );
  OR U606 ( .A(n414), .B(n26), .Z(n417) );
  XNOR U607 ( .A(b[7]), .B(a[6]), .Z(n445) );
  OR U608 ( .A(n445), .B(n415), .Z(n416) );
  NAND U609 ( .A(n417), .B(n416), .Z(n473) );
  XOR U610 ( .A(n472), .B(n473), .Z(n475) );
  XNOR U611 ( .A(n474), .B(n475), .Z(n436) );
  XNOR U612 ( .A(n437), .B(n436), .Z(n438) );
  XOR U613 ( .A(n439), .B(n438), .Z(n433) );
  XNOR U614 ( .A(n432), .B(n433), .Z(n480) );
  XOR U615 ( .A(n481), .B(n480), .Z(n425) );
  NANDN U616 ( .A(n419), .B(n418), .Z(n423) );
  NAND U617 ( .A(n421), .B(n420), .Z(n422) );
  AND U618 ( .A(n423), .B(n422), .Z(n424) );
  XNOR U619 ( .A(n425), .B(n424), .Z(n426) );
  XNOR U620 ( .A(n427), .B(n426), .Z(n485) );
  XNOR U621 ( .A(n486), .B(n485), .Z(c[252]) );
  NANDN U622 ( .A(n425), .B(n424), .Z(n429) );
  NANDN U623 ( .A(n427), .B(n426), .Z(n428) );
  AND U624 ( .A(n429), .B(n428), .Z(n496) );
  NANDN U625 ( .A(n431), .B(n430), .Z(n435) );
  NANDN U626 ( .A(n433), .B(n432), .Z(n434) );
  AND U627 ( .A(n435), .B(n434), .Z(n550) );
  NANDN U628 ( .A(n437), .B(n436), .Z(n441) );
  NANDN U629 ( .A(n439), .B(n438), .Z(n440) );
  AND U630 ( .A(n441), .B(n440), .Z(n549) );
  NAND U631 ( .A(b[0]), .B(a[13]), .Z(n442) );
  XNOR U632 ( .A(b[1]), .B(n442), .Z(n444) );
  NANDN U633 ( .A(b[0]), .B(a[12]), .Z(n443) );
  NAND U634 ( .A(n444), .B(n443), .Z(n534) );
  OR U635 ( .A(n445), .B(n26), .Z(n447) );
  XOR U636 ( .A(b[7]), .B(a[7]), .Z(n527) );
  NAND U637 ( .A(n19486), .B(n527), .Z(n446) );
  NAND U638 ( .A(n447), .B(n446), .Z(n533) );
  XNOR U639 ( .A(n534), .B(n533), .Z(n536) );
  NAND U640 ( .A(n448), .B(n19724), .Z(n450) );
  XOR U641 ( .A(b[11]), .B(a[3]), .Z(n518) );
  NAND U642 ( .A(n19692), .B(n518), .Z(n449) );
  AND U643 ( .A(n450), .B(n449), .Z(n547) );
  XOR U644 ( .A(b[13]), .B(b[12]), .Z(n539) );
  XOR U645 ( .A(b[13]), .B(a[0]), .Z(n451) );
  NAND U646 ( .A(n539), .B(n451), .Z(n452) );
  NANDN U647 ( .A(n452), .B(n19434), .Z(n454) );
  XOR U648 ( .A(b[13]), .B(a[1]), .Z(n540) );
  NANDN U649 ( .A(n19434), .B(n540), .Z(n453) );
  NAND U650 ( .A(n454), .B(n453), .Z(n546) );
  XNOR U651 ( .A(n547), .B(n546), .Z(n535) );
  XOR U652 ( .A(n536), .B(n535), .Z(n508) );
  OR U653 ( .A(n455), .B(n29), .Z(n457) );
  XOR U654 ( .A(b[3]), .B(a[11]), .Z(n530) );
  NAND U655 ( .A(n32), .B(n530), .Z(n456) );
  AND U656 ( .A(n457), .B(n456), .Z(n513) );
  NAND U657 ( .A(n35), .B(n458), .Z(n460) );
  XOR U658 ( .A(b[9]), .B(a[5]), .Z(n543) );
  NAND U659 ( .A(n19598), .B(n543), .Z(n459) );
  NAND U660 ( .A(n460), .B(n459), .Z(n512) );
  XNOR U661 ( .A(n513), .B(n512), .Z(n515) );
  NAND U662 ( .A(b[11]), .B(b[12]), .Z(n461) );
  AND U663 ( .A(b[13]), .B(n461), .Z(n19821) );
  IV U664 ( .A(n19821), .Z(n19846) );
  NOR U665 ( .A(n19846), .B(n466), .Z(n514) );
  XOR U666 ( .A(n515), .B(n514), .Z(n507) );
  NANDN U667 ( .A(n27), .B(n462), .Z(n465) );
  XNOR U668 ( .A(b[5]), .B(a[9]), .Z(n524) );
  OR U669 ( .A(n524), .B(n463), .Z(n464) );
  AND U670 ( .A(n465), .B(n464), .Z(n506) );
  XOR U671 ( .A(n507), .B(n506), .Z(n509) );
  XOR U672 ( .A(n508), .B(n509), .Z(n503) );
  NANDN U673 ( .A(n467), .B(n466), .Z(n471) );
  NANDN U674 ( .A(n469), .B(n468), .Z(n470) );
  AND U675 ( .A(n471), .B(n470), .Z(n501) );
  NANDN U676 ( .A(n473), .B(n472), .Z(n477) );
  OR U677 ( .A(n475), .B(n474), .Z(n476) );
  AND U678 ( .A(n477), .B(n476), .Z(n500) );
  XNOR U679 ( .A(n501), .B(n500), .Z(n502) );
  XNOR U680 ( .A(n503), .B(n502), .Z(n548) );
  XOR U681 ( .A(n549), .B(n548), .Z(n551) );
  XOR U682 ( .A(n550), .B(n551), .Z(n495) );
  NANDN U683 ( .A(n479), .B(n478), .Z(n483) );
  NAND U684 ( .A(n481), .B(n480), .Z(n482) );
  AND U685 ( .A(n483), .B(n482), .Z(n494) );
  XOR U686 ( .A(n495), .B(n494), .Z(n497) );
  XOR U687 ( .A(n496), .B(n497), .Z(n489) );
  XNOR U688 ( .A(n489), .B(sreg[253]), .Z(n491) );
  NANDN U689 ( .A(sreg[252]), .B(n484), .Z(n488) );
  NAND U690 ( .A(n486), .B(n485), .Z(n487) );
  AND U691 ( .A(n488), .B(n487), .Z(n490) );
  XOR U692 ( .A(n491), .B(n490), .Z(c[253]) );
  NANDN U693 ( .A(n489), .B(sreg[253]), .Z(n493) );
  NAND U694 ( .A(n491), .B(n490), .Z(n492) );
  AND U695 ( .A(n493), .B(n492), .Z(n620) );
  XNOR U696 ( .A(sreg[254]), .B(n620), .Z(n622) );
  NANDN U697 ( .A(n495), .B(n494), .Z(n499) );
  OR U698 ( .A(n497), .B(n496), .Z(n498) );
  AND U699 ( .A(n499), .B(n498), .Z(n557) );
  NANDN U700 ( .A(n501), .B(n500), .Z(n505) );
  NANDN U701 ( .A(n503), .B(n502), .Z(n504) );
  AND U702 ( .A(n505), .B(n504), .Z(n616) );
  NANDN U703 ( .A(n507), .B(n506), .Z(n511) );
  OR U704 ( .A(n509), .B(n508), .Z(n510) );
  AND U705 ( .A(n511), .B(n510), .Z(n614) );
  NANDN U706 ( .A(n513), .B(n512), .Z(n517) );
  NAND U707 ( .A(n515), .B(n514), .Z(n516) );
  AND U708 ( .A(n517), .B(n516), .Z(n601) );
  XNOR U709 ( .A(b[13]), .B(b[14]), .Z(n19840) );
  IV U710 ( .A(n19840), .Z(n19805) );
  AND U711 ( .A(a[0]), .B(n19805), .Z(n604) );
  NAND U712 ( .A(n518), .B(n19724), .Z(n520) );
  XOR U713 ( .A(b[11]), .B(a[4]), .Z(n576) );
  NAND U714 ( .A(n19692), .B(n576), .Z(n519) );
  AND U715 ( .A(n520), .B(n519), .Z(n605) );
  XNOR U716 ( .A(n604), .B(n605), .Z(n606) );
  NAND U717 ( .A(b[0]), .B(a[14]), .Z(n521) );
  XNOR U718 ( .A(b[1]), .B(n521), .Z(n523) );
  NANDN U719 ( .A(b[0]), .B(a[13]), .Z(n522) );
  NAND U720 ( .A(n523), .B(n522), .Z(n607) );
  XNOR U721 ( .A(n606), .B(n607), .Z(n598) );
  OR U722 ( .A(n524), .B(n27), .Z(n526) );
  XOR U723 ( .A(b[5]), .B(a[10]), .Z(n570) );
  NAND U724 ( .A(n19342), .B(n570), .Z(n525) );
  AND U725 ( .A(n526), .B(n525), .Z(n582) );
  NAND U726 ( .A(n34), .B(n527), .Z(n529) );
  XOR U727 ( .A(b[7]), .B(a[8]), .Z(n566) );
  NAND U728 ( .A(n19486), .B(n566), .Z(n528) );
  AND U729 ( .A(n529), .B(n528), .Z(n580) );
  NAND U730 ( .A(n31), .B(n530), .Z(n532) );
  XOR U731 ( .A(b[3]), .B(a[12]), .Z(n573) );
  NAND U732 ( .A(n32), .B(n573), .Z(n531) );
  NAND U733 ( .A(n532), .B(n531), .Z(n579) );
  XNOR U734 ( .A(n580), .B(n579), .Z(n581) );
  XOR U735 ( .A(n582), .B(n581), .Z(n599) );
  XNOR U736 ( .A(n598), .B(n599), .Z(n600) );
  XNOR U737 ( .A(n601), .B(n600), .Z(n562) );
  NANDN U738 ( .A(n534), .B(n533), .Z(n538) );
  NAND U739 ( .A(n536), .B(n535), .Z(n537) );
  AND U740 ( .A(n538), .B(n537), .Z(n561) );
  AND U741 ( .A(n539), .B(n19434), .Z(n19808) );
  NAND U742 ( .A(n19808), .B(n540), .Z(n542) );
  XOR U743 ( .A(b[13]), .B(a[2]), .Z(n585) );
  NAND U744 ( .A(n19768), .B(n585), .Z(n541) );
  AND U745 ( .A(n542), .B(n541), .Z(n611) );
  NAND U746 ( .A(n35), .B(n543), .Z(n545) );
  XOR U747 ( .A(b[9]), .B(a[6]), .Z(n595) );
  NAND U748 ( .A(n19598), .B(n595), .Z(n544) );
  NAND U749 ( .A(n545), .B(n544), .Z(n610) );
  XNOR U750 ( .A(n611), .B(n610), .Z(n613) );
  NANDN U751 ( .A(n547), .B(n546), .Z(n612) );
  XNOR U752 ( .A(n613), .B(n612), .Z(n560) );
  XOR U753 ( .A(n561), .B(n560), .Z(n563) );
  XOR U754 ( .A(n562), .B(n563), .Z(n615) );
  XOR U755 ( .A(n614), .B(n615), .Z(n617) );
  XOR U756 ( .A(n616), .B(n617), .Z(n555) );
  NANDN U757 ( .A(n549), .B(n548), .Z(n553) );
  OR U758 ( .A(n551), .B(n550), .Z(n552) );
  AND U759 ( .A(n553), .B(n552), .Z(n554) );
  XNOR U760 ( .A(n555), .B(n554), .Z(n556) );
  XNOR U761 ( .A(n557), .B(n556), .Z(n621) );
  XNOR U762 ( .A(n622), .B(n621), .Z(c[254]) );
  NANDN U763 ( .A(n555), .B(n554), .Z(n559) );
  NANDN U764 ( .A(n557), .B(n556), .Z(n558) );
  AND U765 ( .A(n559), .B(n558), .Z(n633) );
  NANDN U766 ( .A(n561), .B(n560), .Z(n565) );
  NANDN U767 ( .A(n563), .B(n562), .Z(n564) );
  AND U768 ( .A(n565), .B(n564), .Z(n694) );
  NAND U769 ( .A(n34), .B(n566), .Z(n568) );
  XOR U770 ( .A(b[7]), .B(a[9]), .Z(n681) );
  NAND U771 ( .A(n19486), .B(n681), .Z(n567) );
  AND U772 ( .A(n568), .B(n567), .Z(n667) );
  NAND U773 ( .A(b[13]), .B(b[14]), .Z(n19878) );
  ANDN U774 ( .B(n19878), .A(n604), .Z(n569) );
  AND U775 ( .A(b[15]), .B(n569), .Z(n666) );
  XNOR U776 ( .A(n667), .B(n666), .Z(n669) );
  NAND U777 ( .A(n33), .B(n570), .Z(n572) );
  XOR U778 ( .A(b[5]), .B(a[11]), .Z(n690) );
  NAND U779 ( .A(n19342), .B(n690), .Z(n571) );
  AND U780 ( .A(n572), .B(n571), .Z(n663) );
  NAND U781 ( .A(n31), .B(n573), .Z(n575) );
  XOR U782 ( .A(b[3]), .B(a[13]), .Z(n674) );
  NAND U783 ( .A(n32), .B(n674), .Z(n574) );
  AND U784 ( .A(n575), .B(n574), .Z(n661) );
  NAND U785 ( .A(n576), .B(n19724), .Z(n578) );
  XOR U786 ( .A(b[11]), .B(a[5]), .Z(n684) );
  NAND U787 ( .A(n19692), .B(n684), .Z(n577) );
  NAND U788 ( .A(n578), .B(n577), .Z(n660) );
  XNOR U789 ( .A(n661), .B(n660), .Z(n662) );
  XNOR U790 ( .A(n663), .B(n662), .Z(n668) );
  XOR U791 ( .A(n669), .B(n668), .Z(n644) );
  NANDN U792 ( .A(n580), .B(n579), .Z(n584) );
  NANDN U793 ( .A(n582), .B(n581), .Z(n583) );
  AND U794 ( .A(n584), .B(n583), .Z(n642) );
  NAND U795 ( .A(n19808), .B(n585), .Z(n587) );
  XOR U796 ( .A(b[13]), .B(a[3]), .Z(n657) );
  NAND U797 ( .A(n19768), .B(n657), .Z(n586) );
  AND U798 ( .A(n587), .B(n586), .Z(n673) );
  XOR U799 ( .A(b[14]), .B(b[15]), .Z(n588) );
  AND U800 ( .A(n588), .B(n19840), .Z(n19838) );
  XOR U801 ( .A(a[0]), .B(b[15]), .Z(n589) );
  NAND U802 ( .A(n19838), .B(n589), .Z(n591) );
  XOR U803 ( .A(b[15]), .B(a[1]), .Z(n687) );
  AND U804 ( .A(n687), .B(n19805), .Z(n590) );
  ANDN U805 ( .B(n591), .A(n590), .Z(n672) );
  XOR U806 ( .A(n673), .B(n672), .Z(n651) );
  NAND U807 ( .A(b[0]), .B(a[15]), .Z(n592) );
  XNOR U808 ( .A(b[1]), .B(n592), .Z(n594) );
  NANDN U809 ( .A(b[0]), .B(a[14]), .Z(n593) );
  NAND U810 ( .A(n594), .B(n593), .Z(n648) );
  NANDN U811 ( .A(n28), .B(n595), .Z(n597) );
  XNOR U812 ( .A(b[9]), .B(a[7]), .Z(n677) );
  OR U813 ( .A(n677), .B(n678), .Z(n596) );
  NAND U814 ( .A(n597), .B(n596), .Z(n649) );
  XNOR U815 ( .A(n648), .B(n649), .Z(n650) );
  XOR U816 ( .A(n651), .B(n650), .Z(n643) );
  XOR U817 ( .A(n642), .B(n643), .Z(n645) );
  XNOR U818 ( .A(n644), .B(n645), .Z(n693) );
  XNOR U819 ( .A(n694), .B(n693), .Z(n696) );
  NANDN U820 ( .A(n599), .B(n598), .Z(n603) );
  NANDN U821 ( .A(n601), .B(n600), .Z(n602) );
  AND U822 ( .A(n603), .B(n602), .Z(n639) );
  NANDN U823 ( .A(n605), .B(n604), .Z(n609) );
  NANDN U824 ( .A(n607), .B(n606), .Z(n608) );
  AND U825 ( .A(n609), .B(n608), .Z(n637) );
  XNOR U826 ( .A(n637), .B(n636), .Z(n638) );
  XNOR U827 ( .A(n639), .B(n638), .Z(n695) );
  XOR U828 ( .A(n696), .B(n695), .Z(n631) );
  NANDN U829 ( .A(n615), .B(n614), .Z(n619) );
  OR U830 ( .A(n617), .B(n616), .Z(n618) );
  AND U831 ( .A(n619), .B(n618), .Z(n630) );
  XNOR U832 ( .A(n631), .B(n630), .Z(n632) );
  XNOR U833 ( .A(n633), .B(n632), .Z(n625) );
  XNOR U834 ( .A(sreg[255]), .B(n625), .Z(n627) );
  NANDN U835 ( .A(sreg[254]), .B(n620), .Z(n624) );
  NAND U836 ( .A(n622), .B(n621), .Z(n623) );
  NAND U837 ( .A(n624), .B(n623), .Z(n626) );
  XNOR U838 ( .A(n627), .B(n626), .Z(c[255]) );
  NANDN U839 ( .A(sreg[255]), .B(n625), .Z(n629) );
  NAND U840 ( .A(n627), .B(n626), .Z(n628) );
  NAND U841 ( .A(n629), .B(n628), .Z(n771) );
  XNOR U842 ( .A(sreg[256]), .B(n771), .Z(n773) );
  NANDN U843 ( .A(n631), .B(n630), .Z(n635) );
  NANDN U844 ( .A(n633), .B(n632), .Z(n634) );
  AND U845 ( .A(n635), .B(n634), .Z(n701) );
  NANDN U846 ( .A(n637), .B(n636), .Z(n641) );
  NANDN U847 ( .A(n639), .B(n638), .Z(n640) );
  AND U848 ( .A(n641), .B(n640), .Z(n767) );
  NANDN U849 ( .A(n643), .B(n642), .Z(n647) );
  OR U850 ( .A(n645), .B(n644), .Z(n646) );
  AND U851 ( .A(n647), .B(n646), .Z(n765) );
  NANDN U852 ( .A(n649), .B(n648), .Z(n653) );
  NANDN U853 ( .A(n651), .B(n650), .Z(n652) );
  AND U854 ( .A(n653), .B(n652), .Z(n760) );
  NAND U855 ( .A(b[0]), .B(a[16]), .Z(n654) );
  XNOR U856 ( .A(b[1]), .B(n654), .Z(n656) );
  NANDN U857 ( .A(b[0]), .B(a[15]), .Z(n655) );
  NAND U858 ( .A(n656), .B(n655), .Z(n729) );
  NAND U859 ( .A(n19808), .B(n657), .Z(n659) );
  XOR U860 ( .A(b[13]), .B(a[4]), .Z(n735) );
  NAND U861 ( .A(n19768), .B(n735), .Z(n658) );
  AND U862 ( .A(n659), .B(n658), .Z(n727) );
  AND U863 ( .A(b[15]), .B(a[0]), .Z(n726) );
  XOR U864 ( .A(n727), .B(n726), .Z(n728) );
  XNOR U865 ( .A(n729), .B(n728), .Z(n759) );
  XNOR U866 ( .A(n760), .B(n759), .Z(n762) );
  NANDN U867 ( .A(n661), .B(n660), .Z(n665) );
  NANDN U868 ( .A(n663), .B(n662), .Z(n664) );
  AND U869 ( .A(n665), .B(n664), .Z(n761) );
  XOR U870 ( .A(n762), .B(n761), .Z(n756) );
  NANDN U871 ( .A(n667), .B(n666), .Z(n671) );
  NAND U872 ( .A(n669), .B(n668), .Z(n670) );
  AND U873 ( .A(n671), .B(n670), .Z(n754) );
  NOR U874 ( .A(n673), .B(n672), .Z(n707) );
  NANDN U875 ( .A(n29), .B(n674), .Z(n676) );
  XNOR U876 ( .A(b[3]), .B(a[14]), .Z(n744) );
  OR U877 ( .A(n744), .B(n30), .Z(n675) );
  AND U878 ( .A(n676), .B(n675), .Z(n705) );
  OR U879 ( .A(n677), .B(n28), .Z(n680) );
  XNOR U880 ( .A(b[9]), .B(a[8]), .Z(n717) );
  OR U881 ( .A(n717), .B(n678), .Z(n679) );
  NAND U882 ( .A(n680), .B(n679), .Z(n706) );
  XOR U883 ( .A(n705), .B(n706), .Z(n708) );
  XOR U884 ( .A(n707), .B(n708), .Z(n750) );
  NAND U885 ( .A(n34), .B(n681), .Z(n683) );
  XOR U886 ( .A(b[7]), .B(a[10]), .Z(n741) );
  NAND U887 ( .A(n19486), .B(n741), .Z(n682) );
  AND U888 ( .A(n683), .B(n682), .Z(n748) );
  NAND U889 ( .A(n684), .B(n19724), .Z(n686) );
  XOR U890 ( .A(b[11]), .B(a[6]), .Z(n711) );
  NAND U891 ( .A(n19692), .B(n711), .Z(n685) );
  AND U892 ( .A(n686), .B(n685), .Z(n723) );
  NAND U893 ( .A(n19838), .B(n687), .Z(n689) );
  XOR U894 ( .A(b[15]), .B(a[2]), .Z(n714) );
  NAND U895 ( .A(n19805), .B(n714), .Z(n688) );
  AND U896 ( .A(n689), .B(n688), .Z(n721) );
  NAND U897 ( .A(n33), .B(n690), .Z(n692) );
  XOR U898 ( .A(b[5]), .B(a[12]), .Z(n738) );
  NAND U899 ( .A(n19342), .B(n738), .Z(n691) );
  NAND U900 ( .A(n692), .B(n691), .Z(n720) );
  XNOR U901 ( .A(n721), .B(n720), .Z(n722) );
  XNOR U902 ( .A(n723), .B(n722), .Z(n747) );
  XNOR U903 ( .A(n748), .B(n747), .Z(n749) );
  XNOR U904 ( .A(n750), .B(n749), .Z(n753) );
  XNOR U905 ( .A(n754), .B(n753), .Z(n755) );
  XOR U906 ( .A(n756), .B(n755), .Z(n766) );
  XOR U907 ( .A(n765), .B(n766), .Z(n768) );
  XOR U908 ( .A(n767), .B(n768), .Z(n700) );
  NANDN U909 ( .A(n694), .B(n693), .Z(n698) );
  NAND U910 ( .A(n696), .B(n695), .Z(n697) );
  AND U911 ( .A(n698), .B(n697), .Z(n699) );
  XOR U912 ( .A(n700), .B(n699), .Z(n702) );
  XNOR U913 ( .A(n701), .B(n702), .Z(n772) );
  XOR U914 ( .A(n773), .B(n772), .Z(c[256]) );
  NANDN U915 ( .A(n700), .B(n699), .Z(n704) );
  OR U916 ( .A(n702), .B(n701), .Z(n703) );
  AND U917 ( .A(n704), .B(n703), .Z(n779) );
  NANDN U918 ( .A(n706), .B(n705), .Z(n710) );
  OR U919 ( .A(n708), .B(n707), .Z(n709) );
  AND U920 ( .A(n710), .B(n709), .Z(n837) );
  NAND U921 ( .A(n711), .B(n19724), .Z(n713) );
  XOR U922 ( .A(b[11]), .B(a[7]), .Z(n788) );
  NAND U923 ( .A(n19692), .B(n788), .Z(n712) );
  AND U924 ( .A(n713), .B(n712), .Z(n799) );
  NAND U925 ( .A(n19838), .B(n714), .Z(n716) );
  XOR U926 ( .A(b[15]), .B(a[3]), .Z(n791) );
  NAND U927 ( .A(n19805), .B(n791), .Z(n715) );
  AND U928 ( .A(n716), .B(n715), .Z(n798) );
  OR U929 ( .A(n717), .B(n28), .Z(n719) );
  XOR U930 ( .A(b[9]), .B(a[9]), .Z(n794) );
  NAND U931 ( .A(n19598), .B(n794), .Z(n718) );
  NAND U932 ( .A(n719), .B(n718), .Z(n797) );
  XOR U933 ( .A(n798), .B(n797), .Z(n800) );
  XNOR U934 ( .A(n799), .B(n800), .Z(n836) );
  XNOR U935 ( .A(n837), .B(n836), .Z(n838) );
  NANDN U936 ( .A(n721), .B(n720), .Z(n725) );
  NANDN U937 ( .A(n723), .B(n722), .Z(n724) );
  NAND U938 ( .A(n725), .B(n724), .Z(n839) );
  XNOR U939 ( .A(n838), .B(n839), .Z(n785) );
  NANDN U940 ( .A(n727), .B(n726), .Z(n731) );
  OR U941 ( .A(n729), .B(n728), .Z(n730) );
  AND U942 ( .A(n731), .B(n730), .Z(n832) );
  NAND U943 ( .A(b[0]), .B(a[17]), .Z(n732) );
  XNOR U944 ( .A(b[1]), .B(n732), .Z(n734) );
  NANDN U945 ( .A(b[0]), .B(a[16]), .Z(n733) );
  NAND U946 ( .A(n734), .B(n733), .Z(n812) );
  NAND U947 ( .A(n19808), .B(n735), .Z(n737) );
  XOR U948 ( .A(b[13]), .B(a[5]), .Z(n815) );
  NAND U949 ( .A(n19768), .B(n815), .Z(n736) );
  AND U950 ( .A(n737), .B(n736), .Z(n810) );
  AND U951 ( .A(b[15]), .B(a[1]), .Z(n809) );
  XNOR U952 ( .A(n810), .B(n809), .Z(n811) );
  XNOR U953 ( .A(n812), .B(n811), .Z(n830) );
  NAND U954 ( .A(n33), .B(n738), .Z(n740) );
  XOR U955 ( .A(b[5]), .B(a[13]), .Z(n821) );
  NAND U956 ( .A(n19342), .B(n821), .Z(n739) );
  AND U957 ( .A(n740), .B(n739), .Z(n806) );
  NAND U958 ( .A(n34), .B(n741), .Z(n743) );
  XOR U959 ( .A(b[7]), .B(a[11]), .Z(n824) );
  NAND U960 ( .A(n19486), .B(n824), .Z(n742) );
  AND U961 ( .A(n743), .B(n742), .Z(n804) );
  OR U962 ( .A(n744), .B(n29), .Z(n746) );
  XOR U963 ( .A(b[3]), .B(a[15]), .Z(n827) );
  NAND U964 ( .A(n32), .B(n827), .Z(n745) );
  NAND U965 ( .A(n746), .B(n745), .Z(n803) );
  XNOR U966 ( .A(n804), .B(n803), .Z(n805) );
  XOR U967 ( .A(n806), .B(n805), .Z(n831) );
  XOR U968 ( .A(n830), .B(n831), .Z(n833) );
  XOR U969 ( .A(n832), .B(n833), .Z(n783) );
  NANDN U970 ( .A(n748), .B(n747), .Z(n752) );
  NANDN U971 ( .A(n750), .B(n749), .Z(n751) );
  AND U972 ( .A(n752), .B(n751), .Z(n782) );
  XNOR U973 ( .A(n783), .B(n782), .Z(n784) );
  XOR U974 ( .A(n785), .B(n784), .Z(n844) );
  NANDN U975 ( .A(n754), .B(n753), .Z(n758) );
  NANDN U976 ( .A(n756), .B(n755), .Z(n757) );
  AND U977 ( .A(n758), .B(n757), .Z(n843) );
  NANDN U978 ( .A(n760), .B(n759), .Z(n764) );
  NAND U979 ( .A(n762), .B(n761), .Z(n763) );
  AND U980 ( .A(n764), .B(n763), .Z(n842) );
  XOR U981 ( .A(n843), .B(n842), .Z(n845) );
  XOR U982 ( .A(n844), .B(n845), .Z(n777) );
  NANDN U983 ( .A(n766), .B(n765), .Z(n770) );
  OR U984 ( .A(n768), .B(n767), .Z(n769) );
  AND U985 ( .A(n770), .B(n769), .Z(n776) );
  XNOR U986 ( .A(n777), .B(n776), .Z(n778) );
  XNOR U987 ( .A(n779), .B(n778), .Z(n848) );
  XNOR U988 ( .A(sreg[257]), .B(n848), .Z(n850) );
  NANDN U989 ( .A(n771), .B(sreg[256]), .Z(n775) );
  NAND U990 ( .A(n773), .B(n772), .Z(n774) );
  AND U991 ( .A(n775), .B(n774), .Z(n849) );
  XNOR U992 ( .A(n850), .B(n849), .Z(c[257]) );
  NANDN U993 ( .A(n777), .B(n776), .Z(n781) );
  NANDN U994 ( .A(n779), .B(n778), .Z(n780) );
  AND U995 ( .A(n781), .B(n780), .Z(n856) );
  NANDN U996 ( .A(n783), .B(n782), .Z(n787) );
  NAND U997 ( .A(n785), .B(n784), .Z(n786) );
  AND U998 ( .A(n787), .B(n786), .Z(n922) );
  NAND U999 ( .A(n788), .B(n19724), .Z(n790) );
  XOR U1000 ( .A(b[11]), .B(a[8]), .Z(n892) );
  NAND U1001 ( .A(n19692), .B(n892), .Z(n789) );
  AND U1002 ( .A(n790), .B(n789), .Z(n903) );
  NAND U1003 ( .A(n19838), .B(n791), .Z(n793) );
  XOR U1004 ( .A(b[15]), .B(a[4]), .Z(n895) );
  NAND U1005 ( .A(n19805), .B(n895), .Z(n792) );
  AND U1006 ( .A(n793), .B(n792), .Z(n902) );
  NAND U1007 ( .A(n35), .B(n794), .Z(n796) );
  XOR U1008 ( .A(b[9]), .B(a[10]), .Z(n898) );
  NAND U1009 ( .A(n19598), .B(n898), .Z(n795) );
  NAND U1010 ( .A(n796), .B(n795), .Z(n901) );
  XOR U1011 ( .A(n902), .B(n901), .Z(n904) );
  XOR U1012 ( .A(n903), .B(n904), .Z(n914) );
  NANDN U1013 ( .A(n798), .B(n797), .Z(n802) );
  OR U1014 ( .A(n800), .B(n799), .Z(n801) );
  AND U1015 ( .A(n802), .B(n801), .Z(n913) );
  XNOR U1016 ( .A(n914), .B(n913), .Z(n915) );
  NANDN U1017 ( .A(n804), .B(n803), .Z(n808) );
  NANDN U1018 ( .A(n806), .B(n805), .Z(n807) );
  NAND U1019 ( .A(n808), .B(n807), .Z(n916) );
  XNOR U1020 ( .A(n915), .B(n916), .Z(n862) );
  NANDN U1021 ( .A(n810), .B(n809), .Z(n814) );
  NANDN U1022 ( .A(n812), .B(n811), .Z(n813) );
  AND U1023 ( .A(n814), .B(n813), .Z(n888) );
  NAND U1024 ( .A(n19808), .B(n815), .Z(n817) );
  XOR U1025 ( .A(b[13]), .B(a[6]), .Z(n871) );
  NAND U1026 ( .A(n19768), .B(n871), .Z(n816) );
  AND U1027 ( .A(n817), .B(n816), .Z(n866) );
  AND U1028 ( .A(b[15]), .B(a[2]), .Z(n865) );
  XNOR U1029 ( .A(n866), .B(n865), .Z(n867) );
  NAND U1030 ( .A(b[0]), .B(a[18]), .Z(n818) );
  XNOR U1031 ( .A(b[1]), .B(n818), .Z(n820) );
  NANDN U1032 ( .A(b[0]), .B(a[17]), .Z(n819) );
  NAND U1033 ( .A(n820), .B(n819), .Z(n868) );
  XNOR U1034 ( .A(n867), .B(n868), .Z(n886) );
  NAND U1035 ( .A(n33), .B(n821), .Z(n823) );
  XOR U1036 ( .A(b[5]), .B(a[14]), .Z(n877) );
  NAND U1037 ( .A(n19342), .B(n877), .Z(n822) );
  AND U1038 ( .A(n823), .B(n822), .Z(n910) );
  NAND U1039 ( .A(n34), .B(n824), .Z(n826) );
  XOR U1040 ( .A(b[7]), .B(a[12]), .Z(n880) );
  NAND U1041 ( .A(n19486), .B(n880), .Z(n825) );
  AND U1042 ( .A(n826), .B(n825), .Z(n908) );
  NAND U1043 ( .A(n31), .B(n827), .Z(n829) );
  XOR U1044 ( .A(b[3]), .B(a[16]), .Z(n883) );
  NAND U1045 ( .A(n32), .B(n883), .Z(n828) );
  NAND U1046 ( .A(n829), .B(n828), .Z(n907) );
  XNOR U1047 ( .A(n908), .B(n907), .Z(n909) );
  XOR U1048 ( .A(n910), .B(n909), .Z(n887) );
  XOR U1049 ( .A(n886), .B(n887), .Z(n889) );
  XOR U1050 ( .A(n888), .B(n889), .Z(n860) );
  NANDN U1051 ( .A(n831), .B(n830), .Z(n835) );
  OR U1052 ( .A(n833), .B(n832), .Z(n834) );
  AND U1053 ( .A(n835), .B(n834), .Z(n859) );
  XNOR U1054 ( .A(n860), .B(n859), .Z(n861) );
  XOR U1055 ( .A(n862), .B(n861), .Z(n920) );
  NANDN U1056 ( .A(n837), .B(n836), .Z(n841) );
  NANDN U1057 ( .A(n839), .B(n838), .Z(n840) );
  AND U1058 ( .A(n841), .B(n840), .Z(n919) );
  XNOR U1059 ( .A(n920), .B(n919), .Z(n921) );
  XOR U1060 ( .A(n922), .B(n921), .Z(n854) );
  NANDN U1061 ( .A(n843), .B(n842), .Z(n847) );
  OR U1062 ( .A(n845), .B(n844), .Z(n846) );
  AND U1063 ( .A(n847), .B(n846), .Z(n853) );
  XNOR U1064 ( .A(n854), .B(n853), .Z(n855) );
  XNOR U1065 ( .A(n856), .B(n855), .Z(n925) );
  XNOR U1066 ( .A(sreg[258]), .B(n925), .Z(n927) );
  NANDN U1067 ( .A(sreg[257]), .B(n848), .Z(n852) );
  NAND U1068 ( .A(n850), .B(n849), .Z(n851) );
  NAND U1069 ( .A(n852), .B(n851), .Z(n926) );
  XNOR U1070 ( .A(n927), .B(n926), .Z(c[258]) );
  NANDN U1071 ( .A(n854), .B(n853), .Z(n858) );
  NANDN U1072 ( .A(n856), .B(n855), .Z(n857) );
  AND U1073 ( .A(n858), .B(n857), .Z(n932) );
  NANDN U1074 ( .A(n860), .B(n859), .Z(n864) );
  NAND U1075 ( .A(n862), .B(n861), .Z(n863) );
  AND U1076 ( .A(n864), .B(n863), .Z(n999) );
  NANDN U1077 ( .A(n866), .B(n865), .Z(n870) );
  NANDN U1078 ( .A(n868), .B(n867), .Z(n869) );
  AND U1079 ( .A(n870), .B(n869), .Z(n965) );
  NAND U1080 ( .A(n19808), .B(n871), .Z(n873) );
  XOR U1081 ( .A(b[13]), .B(a[7]), .Z(n951) );
  NAND U1082 ( .A(n19768), .B(n951), .Z(n872) );
  AND U1083 ( .A(n873), .B(n872), .Z(n943) );
  AND U1084 ( .A(b[15]), .B(a[3]), .Z(n942) );
  XNOR U1085 ( .A(n943), .B(n942), .Z(n944) );
  NAND U1086 ( .A(b[0]), .B(a[19]), .Z(n874) );
  XNOR U1087 ( .A(b[1]), .B(n874), .Z(n876) );
  NANDN U1088 ( .A(b[0]), .B(a[18]), .Z(n875) );
  NAND U1089 ( .A(n876), .B(n875), .Z(n945) );
  XNOR U1090 ( .A(n944), .B(n945), .Z(n963) );
  NAND U1091 ( .A(n33), .B(n877), .Z(n879) );
  XOR U1092 ( .A(b[5]), .B(a[15]), .Z(n954) );
  NAND U1093 ( .A(n19342), .B(n954), .Z(n878) );
  AND U1094 ( .A(n879), .B(n878), .Z(n987) );
  NAND U1095 ( .A(n34), .B(n880), .Z(n882) );
  XOR U1096 ( .A(b[7]), .B(a[13]), .Z(n957) );
  NAND U1097 ( .A(n19486), .B(n957), .Z(n881) );
  AND U1098 ( .A(n882), .B(n881), .Z(n985) );
  NAND U1099 ( .A(n31), .B(n883), .Z(n885) );
  XOR U1100 ( .A(b[3]), .B(a[17]), .Z(n960) );
  NAND U1101 ( .A(n32), .B(n960), .Z(n884) );
  NAND U1102 ( .A(n885), .B(n884), .Z(n984) );
  XNOR U1103 ( .A(n985), .B(n984), .Z(n986) );
  XOR U1104 ( .A(n987), .B(n986), .Z(n964) );
  XOR U1105 ( .A(n963), .B(n964), .Z(n966) );
  XOR U1106 ( .A(n965), .B(n966), .Z(n937) );
  NANDN U1107 ( .A(n887), .B(n886), .Z(n891) );
  OR U1108 ( .A(n889), .B(n888), .Z(n890) );
  AND U1109 ( .A(n891), .B(n890), .Z(n936) );
  XNOR U1110 ( .A(n937), .B(n936), .Z(n939) );
  NAND U1111 ( .A(n892), .B(n19724), .Z(n894) );
  XOR U1112 ( .A(b[11]), .B(a[9]), .Z(n969) );
  NAND U1113 ( .A(n19692), .B(n969), .Z(n893) );
  AND U1114 ( .A(n894), .B(n893), .Z(n980) );
  NAND U1115 ( .A(n19838), .B(n895), .Z(n897) );
  XOR U1116 ( .A(b[15]), .B(a[5]), .Z(n972) );
  NAND U1117 ( .A(n19805), .B(n972), .Z(n896) );
  AND U1118 ( .A(n897), .B(n896), .Z(n979) );
  NAND U1119 ( .A(n35), .B(n898), .Z(n900) );
  XOR U1120 ( .A(b[9]), .B(a[11]), .Z(n975) );
  NAND U1121 ( .A(n19598), .B(n975), .Z(n899) );
  NAND U1122 ( .A(n900), .B(n899), .Z(n978) );
  XOR U1123 ( .A(n979), .B(n978), .Z(n981) );
  XOR U1124 ( .A(n980), .B(n981), .Z(n991) );
  NANDN U1125 ( .A(n902), .B(n901), .Z(n906) );
  OR U1126 ( .A(n904), .B(n903), .Z(n905) );
  AND U1127 ( .A(n906), .B(n905), .Z(n990) );
  XNOR U1128 ( .A(n991), .B(n990), .Z(n992) );
  NANDN U1129 ( .A(n908), .B(n907), .Z(n912) );
  NANDN U1130 ( .A(n910), .B(n909), .Z(n911) );
  NAND U1131 ( .A(n912), .B(n911), .Z(n993) );
  XNOR U1132 ( .A(n992), .B(n993), .Z(n938) );
  XOR U1133 ( .A(n939), .B(n938), .Z(n997) );
  NANDN U1134 ( .A(n914), .B(n913), .Z(n918) );
  NANDN U1135 ( .A(n916), .B(n915), .Z(n917) );
  AND U1136 ( .A(n918), .B(n917), .Z(n996) );
  XNOR U1137 ( .A(n997), .B(n996), .Z(n998) );
  XOR U1138 ( .A(n999), .B(n998), .Z(n931) );
  NANDN U1139 ( .A(n920), .B(n919), .Z(n924) );
  NAND U1140 ( .A(n922), .B(n921), .Z(n923) );
  AND U1141 ( .A(n924), .B(n923), .Z(n930) );
  XOR U1142 ( .A(n931), .B(n930), .Z(n933) );
  XOR U1143 ( .A(n932), .B(n933), .Z(n1002) );
  XNOR U1144 ( .A(n1002), .B(sreg[259]), .Z(n1004) );
  NANDN U1145 ( .A(sreg[258]), .B(n925), .Z(n929) );
  NAND U1146 ( .A(n927), .B(n926), .Z(n928) );
  AND U1147 ( .A(n929), .B(n928), .Z(n1003) );
  XOR U1148 ( .A(n1004), .B(n1003), .Z(c[259]) );
  NANDN U1149 ( .A(n931), .B(n930), .Z(n935) );
  OR U1150 ( .A(n933), .B(n932), .Z(n934) );
  AND U1151 ( .A(n935), .B(n934), .Z(n1010) );
  NANDN U1152 ( .A(n937), .B(n936), .Z(n941) );
  NAND U1153 ( .A(n939), .B(n938), .Z(n940) );
  AND U1154 ( .A(n941), .B(n940), .Z(n1076) );
  NANDN U1155 ( .A(n943), .B(n942), .Z(n947) );
  NANDN U1156 ( .A(n945), .B(n944), .Z(n946) );
  AND U1157 ( .A(n947), .B(n946), .Z(n1042) );
  NAND U1158 ( .A(b[0]), .B(a[20]), .Z(n948) );
  XNOR U1159 ( .A(b[1]), .B(n948), .Z(n950) );
  NANDN U1160 ( .A(b[0]), .B(a[19]), .Z(n949) );
  NAND U1161 ( .A(n950), .B(n949), .Z(n1022) );
  NAND U1162 ( .A(n19808), .B(n951), .Z(n953) );
  XOR U1163 ( .A(b[13]), .B(a[8]), .Z(n1025) );
  NAND U1164 ( .A(n19768), .B(n1025), .Z(n952) );
  AND U1165 ( .A(n953), .B(n952), .Z(n1020) );
  AND U1166 ( .A(b[15]), .B(a[4]), .Z(n1019) );
  XNOR U1167 ( .A(n1020), .B(n1019), .Z(n1021) );
  XNOR U1168 ( .A(n1022), .B(n1021), .Z(n1040) );
  NAND U1169 ( .A(n33), .B(n954), .Z(n956) );
  XOR U1170 ( .A(b[5]), .B(a[16]), .Z(n1031) );
  NAND U1171 ( .A(n19342), .B(n1031), .Z(n955) );
  AND U1172 ( .A(n956), .B(n955), .Z(n1064) );
  NAND U1173 ( .A(n34), .B(n957), .Z(n959) );
  XOR U1174 ( .A(b[7]), .B(a[14]), .Z(n1034) );
  NAND U1175 ( .A(n19486), .B(n1034), .Z(n958) );
  AND U1176 ( .A(n959), .B(n958), .Z(n1062) );
  NAND U1177 ( .A(n31), .B(n960), .Z(n962) );
  XOR U1178 ( .A(b[3]), .B(a[18]), .Z(n1037) );
  NAND U1179 ( .A(n32), .B(n1037), .Z(n961) );
  NAND U1180 ( .A(n962), .B(n961), .Z(n1061) );
  XNOR U1181 ( .A(n1062), .B(n1061), .Z(n1063) );
  XOR U1182 ( .A(n1064), .B(n1063), .Z(n1041) );
  XOR U1183 ( .A(n1040), .B(n1041), .Z(n1043) );
  XOR U1184 ( .A(n1042), .B(n1043), .Z(n1014) );
  NANDN U1185 ( .A(n964), .B(n963), .Z(n968) );
  OR U1186 ( .A(n966), .B(n965), .Z(n967) );
  AND U1187 ( .A(n968), .B(n967), .Z(n1013) );
  XNOR U1188 ( .A(n1014), .B(n1013), .Z(n1016) );
  NAND U1189 ( .A(n969), .B(n19724), .Z(n971) );
  XOR U1190 ( .A(b[11]), .B(a[10]), .Z(n1046) );
  NAND U1191 ( .A(n19692), .B(n1046), .Z(n970) );
  AND U1192 ( .A(n971), .B(n970), .Z(n1057) );
  NAND U1193 ( .A(n19838), .B(n972), .Z(n974) );
  XOR U1194 ( .A(b[15]), .B(a[6]), .Z(n1049) );
  NAND U1195 ( .A(n19805), .B(n1049), .Z(n973) );
  AND U1196 ( .A(n974), .B(n973), .Z(n1056) );
  NAND U1197 ( .A(n35), .B(n975), .Z(n977) );
  XOR U1198 ( .A(b[9]), .B(a[12]), .Z(n1052) );
  NAND U1199 ( .A(n19598), .B(n1052), .Z(n976) );
  NAND U1200 ( .A(n977), .B(n976), .Z(n1055) );
  XOR U1201 ( .A(n1056), .B(n1055), .Z(n1058) );
  XOR U1202 ( .A(n1057), .B(n1058), .Z(n1068) );
  NANDN U1203 ( .A(n979), .B(n978), .Z(n983) );
  OR U1204 ( .A(n981), .B(n980), .Z(n982) );
  AND U1205 ( .A(n983), .B(n982), .Z(n1067) );
  XNOR U1206 ( .A(n1068), .B(n1067), .Z(n1069) );
  NANDN U1207 ( .A(n985), .B(n984), .Z(n989) );
  NANDN U1208 ( .A(n987), .B(n986), .Z(n988) );
  NAND U1209 ( .A(n989), .B(n988), .Z(n1070) );
  XNOR U1210 ( .A(n1069), .B(n1070), .Z(n1015) );
  XOR U1211 ( .A(n1016), .B(n1015), .Z(n1074) );
  NANDN U1212 ( .A(n991), .B(n990), .Z(n995) );
  NANDN U1213 ( .A(n993), .B(n992), .Z(n994) );
  AND U1214 ( .A(n995), .B(n994), .Z(n1073) );
  XNOR U1215 ( .A(n1074), .B(n1073), .Z(n1075) );
  XOR U1216 ( .A(n1076), .B(n1075), .Z(n1008) );
  NANDN U1217 ( .A(n997), .B(n996), .Z(n1001) );
  NAND U1218 ( .A(n999), .B(n998), .Z(n1000) );
  AND U1219 ( .A(n1001), .B(n1000), .Z(n1007) );
  XNOR U1220 ( .A(n1008), .B(n1007), .Z(n1009) );
  XNOR U1221 ( .A(n1010), .B(n1009), .Z(n1079) );
  XNOR U1222 ( .A(sreg[260]), .B(n1079), .Z(n1081) );
  NANDN U1223 ( .A(n1002), .B(sreg[259]), .Z(n1006) );
  NAND U1224 ( .A(n1004), .B(n1003), .Z(n1005) );
  AND U1225 ( .A(n1006), .B(n1005), .Z(n1080) );
  XNOR U1226 ( .A(n1081), .B(n1080), .Z(c[260]) );
  NANDN U1227 ( .A(n1008), .B(n1007), .Z(n1012) );
  NANDN U1228 ( .A(n1010), .B(n1009), .Z(n1011) );
  AND U1229 ( .A(n1012), .B(n1011), .Z(n1087) );
  NANDN U1230 ( .A(n1014), .B(n1013), .Z(n1018) );
  NAND U1231 ( .A(n1016), .B(n1015), .Z(n1017) );
  AND U1232 ( .A(n1018), .B(n1017), .Z(n1153) );
  NANDN U1233 ( .A(n1020), .B(n1019), .Z(n1024) );
  NANDN U1234 ( .A(n1022), .B(n1021), .Z(n1023) );
  AND U1235 ( .A(n1024), .B(n1023), .Z(n1119) );
  NAND U1236 ( .A(n19808), .B(n1025), .Z(n1027) );
  XOR U1237 ( .A(b[13]), .B(a[9]), .Z(n1105) );
  NAND U1238 ( .A(n19768), .B(n1105), .Z(n1026) );
  AND U1239 ( .A(n1027), .B(n1026), .Z(n1097) );
  AND U1240 ( .A(b[15]), .B(a[5]), .Z(n1096) );
  XNOR U1241 ( .A(n1097), .B(n1096), .Z(n1098) );
  NAND U1242 ( .A(b[0]), .B(a[21]), .Z(n1028) );
  XNOR U1243 ( .A(b[1]), .B(n1028), .Z(n1030) );
  NANDN U1244 ( .A(b[0]), .B(a[20]), .Z(n1029) );
  NAND U1245 ( .A(n1030), .B(n1029), .Z(n1099) );
  XNOR U1246 ( .A(n1098), .B(n1099), .Z(n1117) );
  NAND U1247 ( .A(n33), .B(n1031), .Z(n1033) );
  XOR U1248 ( .A(b[5]), .B(a[17]), .Z(n1108) );
  NAND U1249 ( .A(n19342), .B(n1108), .Z(n1032) );
  AND U1250 ( .A(n1033), .B(n1032), .Z(n1141) );
  NAND U1251 ( .A(n34), .B(n1034), .Z(n1036) );
  XOR U1252 ( .A(b[7]), .B(a[15]), .Z(n1111) );
  NAND U1253 ( .A(n19486), .B(n1111), .Z(n1035) );
  AND U1254 ( .A(n1036), .B(n1035), .Z(n1139) );
  NAND U1255 ( .A(n31), .B(n1037), .Z(n1039) );
  XOR U1256 ( .A(b[3]), .B(a[19]), .Z(n1114) );
  NAND U1257 ( .A(n32), .B(n1114), .Z(n1038) );
  NAND U1258 ( .A(n1039), .B(n1038), .Z(n1138) );
  XNOR U1259 ( .A(n1139), .B(n1138), .Z(n1140) );
  XOR U1260 ( .A(n1141), .B(n1140), .Z(n1118) );
  XOR U1261 ( .A(n1117), .B(n1118), .Z(n1120) );
  XOR U1262 ( .A(n1119), .B(n1120), .Z(n1091) );
  NANDN U1263 ( .A(n1041), .B(n1040), .Z(n1045) );
  OR U1264 ( .A(n1043), .B(n1042), .Z(n1044) );
  AND U1265 ( .A(n1045), .B(n1044), .Z(n1090) );
  XNOR U1266 ( .A(n1091), .B(n1090), .Z(n1093) );
  NAND U1267 ( .A(n1046), .B(n19724), .Z(n1048) );
  XOR U1268 ( .A(b[11]), .B(a[11]), .Z(n1123) );
  NAND U1269 ( .A(n19692), .B(n1123), .Z(n1047) );
  AND U1270 ( .A(n1048), .B(n1047), .Z(n1134) );
  NAND U1271 ( .A(n19838), .B(n1049), .Z(n1051) );
  XOR U1272 ( .A(b[15]), .B(a[7]), .Z(n1126) );
  NAND U1273 ( .A(n19805), .B(n1126), .Z(n1050) );
  AND U1274 ( .A(n1051), .B(n1050), .Z(n1133) );
  NAND U1275 ( .A(n35), .B(n1052), .Z(n1054) );
  XOR U1276 ( .A(b[9]), .B(a[13]), .Z(n1129) );
  NAND U1277 ( .A(n19598), .B(n1129), .Z(n1053) );
  NAND U1278 ( .A(n1054), .B(n1053), .Z(n1132) );
  XOR U1279 ( .A(n1133), .B(n1132), .Z(n1135) );
  XOR U1280 ( .A(n1134), .B(n1135), .Z(n1145) );
  NANDN U1281 ( .A(n1056), .B(n1055), .Z(n1060) );
  OR U1282 ( .A(n1058), .B(n1057), .Z(n1059) );
  AND U1283 ( .A(n1060), .B(n1059), .Z(n1144) );
  XNOR U1284 ( .A(n1145), .B(n1144), .Z(n1146) );
  NANDN U1285 ( .A(n1062), .B(n1061), .Z(n1066) );
  NANDN U1286 ( .A(n1064), .B(n1063), .Z(n1065) );
  NAND U1287 ( .A(n1066), .B(n1065), .Z(n1147) );
  XNOR U1288 ( .A(n1146), .B(n1147), .Z(n1092) );
  XOR U1289 ( .A(n1093), .B(n1092), .Z(n1151) );
  NANDN U1290 ( .A(n1068), .B(n1067), .Z(n1072) );
  NANDN U1291 ( .A(n1070), .B(n1069), .Z(n1071) );
  AND U1292 ( .A(n1072), .B(n1071), .Z(n1150) );
  XNOR U1293 ( .A(n1151), .B(n1150), .Z(n1152) );
  XOR U1294 ( .A(n1153), .B(n1152), .Z(n1085) );
  NANDN U1295 ( .A(n1074), .B(n1073), .Z(n1078) );
  NAND U1296 ( .A(n1076), .B(n1075), .Z(n1077) );
  AND U1297 ( .A(n1078), .B(n1077), .Z(n1084) );
  XNOR U1298 ( .A(n1085), .B(n1084), .Z(n1086) );
  XNOR U1299 ( .A(n1087), .B(n1086), .Z(n1156) );
  XNOR U1300 ( .A(sreg[261]), .B(n1156), .Z(n1158) );
  NANDN U1301 ( .A(sreg[260]), .B(n1079), .Z(n1083) );
  NAND U1302 ( .A(n1081), .B(n1080), .Z(n1082) );
  NAND U1303 ( .A(n1083), .B(n1082), .Z(n1157) );
  XNOR U1304 ( .A(n1158), .B(n1157), .Z(c[261]) );
  NANDN U1305 ( .A(n1085), .B(n1084), .Z(n1089) );
  NANDN U1306 ( .A(n1087), .B(n1086), .Z(n1088) );
  AND U1307 ( .A(n1089), .B(n1088), .Z(n1164) );
  NANDN U1308 ( .A(n1091), .B(n1090), .Z(n1095) );
  NAND U1309 ( .A(n1093), .B(n1092), .Z(n1094) );
  AND U1310 ( .A(n1095), .B(n1094), .Z(n1230) );
  NANDN U1311 ( .A(n1097), .B(n1096), .Z(n1101) );
  NANDN U1312 ( .A(n1099), .B(n1098), .Z(n1100) );
  AND U1313 ( .A(n1101), .B(n1100), .Z(n1217) );
  NAND U1314 ( .A(b[0]), .B(a[22]), .Z(n1102) );
  XNOR U1315 ( .A(b[1]), .B(n1102), .Z(n1104) );
  NANDN U1316 ( .A(b[0]), .B(a[21]), .Z(n1103) );
  NAND U1317 ( .A(n1104), .B(n1103), .Z(n1197) );
  NAND U1318 ( .A(n19808), .B(n1105), .Z(n1107) );
  XOR U1319 ( .A(b[13]), .B(a[10]), .Z(n1203) );
  NAND U1320 ( .A(n19768), .B(n1203), .Z(n1106) );
  AND U1321 ( .A(n1107), .B(n1106), .Z(n1195) );
  AND U1322 ( .A(b[15]), .B(a[6]), .Z(n1194) );
  XNOR U1323 ( .A(n1195), .B(n1194), .Z(n1196) );
  XNOR U1324 ( .A(n1197), .B(n1196), .Z(n1215) );
  NAND U1325 ( .A(n33), .B(n1108), .Z(n1110) );
  XOR U1326 ( .A(b[5]), .B(a[18]), .Z(n1206) );
  NAND U1327 ( .A(n19342), .B(n1206), .Z(n1109) );
  AND U1328 ( .A(n1110), .B(n1109), .Z(n1191) );
  NAND U1329 ( .A(n34), .B(n1111), .Z(n1113) );
  XOR U1330 ( .A(b[7]), .B(a[16]), .Z(n1209) );
  NAND U1331 ( .A(n19486), .B(n1209), .Z(n1112) );
  AND U1332 ( .A(n1113), .B(n1112), .Z(n1189) );
  NAND U1333 ( .A(n31), .B(n1114), .Z(n1116) );
  XOR U1334 ( .A(b[3]), .B(a[20]), .Z(n1212) );
  NAND U1335 ( .A(n32), .B(n1212), .Z(n1115) );
  NAND U1336 ( .A(n1116), .B(n1115), .Z(n1188) );
  XNOR U1337 ( .A(n1189), .B(n1188), .Z(n1190) );
  XOR U1338 ( .A(n1191), .B(n1190), .Z(n1216) );
  XOR U1339 ( .A(n1215), .B(n1216), .Z(n1218) );
  XOR U1340 ( .A(n1217), .B(n1218), .Z(n1168) );
  NANDN U1341 ( .A(n1118), .B(n1117), .Z(n1122) );
  OR U1342 ( .A(n1120), .B(n1119), .Z(n1121) );
  AND U1343 ( .A(n1122), .B(n1121), .Z(n1167) );
  XNOR U1344 ( .A(n1168), .B(n1167), .Z(n1170) );
  NAND U1345 ( .A(n1123), .B(n19724), .Z(n1125) );
  XOR U1346 ( .A(b[11]), .B(a[12]), .Z(n1173) );
  NAND U1347 ( .A(n19692), .B(n1173), .Z(n1124) );
  AND U1348 ( .A(n1125), .B(n1124), .Z(n1184) );
  NAND U1349 ( .A(n19838), .B(n1126), .Z(n1128) );
  XOR U1350 ( .A(b[15]), .B(a[8]), .Z(n1176) );
  NAND U1351 ( .A(n19805), .B(n1176), .Z(n1127) );
  AND U1352 ( .A(n1128), .B(n1127), .Z(n1183) );
  NAND U1353 ( .A(n35), .B(n1129), .Z(n1131) );
  XOR U1354 ( .A(b[9]), .B(a[14]), .Z(n1179) );
  NAND U1355 ( .A(n19598), .B(n1179), .Z(n1130) );
  NAND U1356 ( .A(n1131), .B(n1130), .Z(n1182) );
  XOR U1357 ( .A(n1183), .B(n1182), .Z(n1185) );
  XOR U1358 ( .A(n1184), .B(n1185), .Z(n1222) );
  NANDN U1359 ( .A(n1133), .B(n1132), .Z(n1137) );
  OR U1360 ( .A(n1135), .B(n1134), .Z(n1136) );
  AND U1361 ( .A(n1137), .B(n1136), .Z(n1221) );
  XNOR U1362 ( .A(n1222), .B(n1221), .Z(n1223) );
  NANDN U1363 ( .A(n1139), .B(n1138), .Z(n1143) );
  NANDN U1364 ( .A(n1141), .B(n1140), .Z(n1142) );
  NAND U1365 ( .A(n1143), .B(n1142), .Z(n1224) );
  XNOR U1366 ( .A(n1223), .B(n1224), .Z(n1169) );
  XOR U1367 ( .A(n1170), .B(n1169), .Z(n1228) );
  NANDN U1368 ( .A(n1145), .B(n1144), .Z(n1149) );
  NANDN U1369 ( .A(n1147), .B(n1146), .Z(n1148) );
  AND U1370 ( .A(n1149), .B(n1148), .Z(n1227) );
  XNOR U1371 ( .A(n1228), .B(n1227), .Z(n1229) );
  XOR U1372 ( .A(n1230), .B(n1229), .Z(n1162) );
  NANDN U1373 ( .A(n1151), .B(n1150), .Z(n1155) );
  NAND U1374 ( .A(n1153), .B(n1152), .Z(n1154) );
  AND U1375 ( .A(n1155), .B(n1154), .Z(n1161) );
  XNOR U1376 ( .A(n1162), .B(n1161), .Z(n1163) );
  XNOR U1377 ( .A(n1164), .B(n1163), .Z(n1233) );
  XNOR U1378 ( .A(sreg[262]), .B(n1233), .Z(n1235) );
  NANDN U1379 ( .A(sreg[261]), .B(n1156), .Z(n1160) );
  NAND U1380 ( .A(n1158), .B(n1157), .Z(n1159) );
  NAND U1381 ( .A(n1160), .B(n1159), .Z(n1234) );
  XNOR U1382 ( .A(n1235), .B(n1234), .Z(c[262]) );
  NANDN U1383 ( .A(n1162), .B(n1161), .Z(n1166) );
  NANDN U1384 ( .A(n1164), .B(n1163), .Z(n1165) );
  AND U1385 ( .A(n1166), .B(n1165), .Z(n1241) );
  NANDN U1386 ( .A(n1168), .B(n1167), .Z(n1172) );
  NAND U1387 ( .A(n1170), .B(n1169), .Z(n1171) );
  AND U1388 ( .A(n1172), .B(n1171), .Z(n1307) );
  NAND U1389 ( .A(n1173), .B(n19724), .Z(n1175) );
  XOR U1390 ( .A(b[11]), .B(a[13]), .Z(n1250) );
  NAND U1391 ( .A(n19692), .B(n1250), .Z(n1174) );
  AND U1392 ( .A(n1175), .B(n1174), .Z(n1261) );
  NAND U1393 ( .A(n19838), .B(n1176), .Z(n1178) );
  XOR U1394 ( .A(b[15]), .B(a[9]), .Z(n1253) );
  NAND U1395 ( .A(n19805), .B(n1253), .Z(n1177) );
  AND U1396 ( .A(n1178), .B(n1177), .Z(n1260) );
  NAND U1397 ( .A(n35), .B(n1179), .Z(n1181) );
  XOR U1398 ( .A(b[9]), .B(a[15]), .Z(n1256) );
  NAND U1399 ( .A(n19598), .B(n1256), .Z(n1180) );
  NAND U1400 ( .A(n1181), .B(n1180), .Z(n1259) );
  XOR U1401 ( .A(n1260), .B(n1259), .Z(n1262) );
  XOR U1402 ( .A(n1261), .B(n1262), .Z(n1299) );
  NANDN U1403 ( .A(n1183), .B(n1182), .Z(n1187) );
  OR U1404 ( .A(n1185), .B(n1184), .Z(n1186) );
  AND U1405 ( .A(n1187), .B(n1186), .Z(n1298) );
  XNOR U1406 ( .A(n1299), .B(n1298), .Z(n1300) );
  NANDN U1407 ( .A(n1189), .B(n1188), .Z(n1193) );
  NANDN U1408 ( .A(n1191), .B(n1190), .Z(n1192) );
  NAND U1409 ( .A(n1193), .B(n1192), .Z(n1301) );
  XNOR U1410 ( .A(n1300), .B(n1301), .Z(n1247) );
  NANDN U1411 ( .A(n1195), .B(n1194), .Z(n1199) );
  NANDN U1412 ( .A(n1197), .B(n1196), .Z(n1198) );
  AND U1413 ( .A(n1199), .B(n1198), .Z(n1294) );
  NAND U1414 ( .A(b[0]), .B(a[23]), .Z(n1200) );
  XNOR U1415 ( .A(b[1]), .B(n1200), .Z(n1202) );
  NANDN U1416 ( .A(b[0]), .B(a[22]), .Z(n1201) );
  NAND U1417 ( .A(n1202), .B(n1201), .Z(n1274) );
  NAND U1418 ( .A(n19808), .B(n1203), .Z(n1205) );
  XOR U1419 ( .A(b[13]), .B(a[11]), .Z(n1277) );
  NAND U1420 ( .A(n19768), .B(n1277), .Z(n1204) );
  AND U1421 ( .A(n1205), .B(n1204), .Z(n1272) );
  AND U1422 ( .A(b[15]), .B(a[7]), .Z(n1271) );
  XNOR U1423 ( .A(n1272), .B(n1271), .Z(n1273) );
  XNOR U1424 ( .A(n1274), .B(n1273), .Z(n1292) );
  NAND U1425 ( .A(n33), .B(n1206), .Z(n1208) );
  XOR U1426 ( .A(b[5]), .B(a[19]), .Z(n1283) );
  NAND U1427 ( .A(n19342), .B(n1283), .Z(n1207) );
  AND U1428 ( .A(n1208), .B(n1207), .Z(n1268) );
  NAND U1429 ( .A(n34), .B(n1209), .Z(n1211) );
  XOR U1430 ( .A(b[7]), .B(a[17]), .Z(n1286) );
  NAND U1431 ( .A(n19486), .B(n1286), .Z(n1210) );
  AND U1432 ( .A(n1211), .B(n1210), .Z(n1266) );
  NAND U1433 ( .A(n31), .B(n1212), .Z(n1214) );
  XOR U1434 ( .A(b[3]), .B(a[21]), .Z(n1289) );
  NAND U1435 ( .A(n32), .B(n1289), .Z(n1213) );
  NAND U1436 ( .A(n1214), .B(n1213), .Z(n1265) );
  XNOR U1437 ( .A(n1266), .B(n1265), .Z(n1267) );
  XOR U1438 ( .A(n1268), .B(n1267), .Z(n1293) );
  XOR U1439 ( .A(n1292), .B(n1293), .Z(n1295) );
  XOR U1440 ( .A(n1294), .B(n1295), .Z(n1245) );
  NANDN U1441 ( .A(n1216), .B(n1215), .Z(n1220) );
  OR U1442 ( .A(n1218), .B(n1217), .Z(n1219) );
  AND U1443 ( .A(n1220), .B(n1219), .Z(n1244) );
  XNOR U1444 ( .A(n1245), .B(n1244), .Z(n1246) );
  XOR U1445 ( .A(n1247), .B(n1246), .Z(n1305) );
  NANDN U1446 ( .A(n1222), .B(n1221), .Z(n1226) );
  NANDN U1447 ( .A(n1224), .B(n1223), .Z(n1225) );
  AND U1448 ( .A(n1226), .B(n1225), .Z(n1304) );
  XNOR U1449 ( .A(n1305), .B(n1304), .Z(n1306) );
  XOR U1450 ( .A(n1307), .B(n1306), .Z(n1239) );
  NANDN U1451 ( .A(n1228), .B(n1227), .Z(n1232) );
  NAND U1452 ( .A(n1230), .B(n1229), .Z(n1231) );
  AND U1453 ( .A(n1232), .B(n1231), .Z(n1238) );
  XNOR U1454 ( .A(n1239), .B(n1238), .Z(n1240) );
  XNOR U1455 ( .A(n1241), .B(n1240), .Z(n1310) );
  XNOR U1456 ( .A(sreg[263]), .B(n1310), .Z(n1312) );
  NANDN U1457 ( .A(sreg[262]), .B(n1233), .Z(n1237) );
  NAND U1458 ( .A(n1235), .B(n1234), .Z(n1236) );
  NAND U1459 ( .A(n1237), .B(n1236), .Z(n1311) );
  XNOR U1460 ( .A(n1312), .B(n1311), .Z(c[263]) );
  NANDN U1461 ( .A(n1239), .B(n1238), .Z(n1243) );
  NANDN U1462 ( .A(n1241), .B(n1240), .Z(n1242) );
  AND U1463 ( .A(n1243), .B(n1242), .Z(n1318) );
  NANDN U1464 ( .A(n1245), .B(n1244), .Z(n1249) );
  NAND U1465 ( .A(n1247), .B(n1246), .Z(n1248) );
  AND U1466 ( .A(n1249), .B(n1248), .Z(n1384) );
  NAND U1467 ( .A(n1250), .B(n19724), .Z(n1252) );
  XOR U1468 ( .A(b[11]), .B(a[14]), .Z(n1354) );
  NAND U1469 ( .A(n19692), .B(n1354), .Z(n1251) );
  AND U1470 ( .A(n1252), .B(n1251), .Z(n1365) );
  NAND U1471 ( .A(n19838), .B(n1253), .Z(n1255) );
  XOR U1472 ( .A(b[15]), .B(a[10]), .Z(n1357) );
  NAND U1473 ( .A(n19805), .B(n1357), .Z(n1254) );
  AND U1474 ( .A(n1255), .B(n1254), .Z(n1364) );
  NAND U1475 ( .A(n35), .B(n1256), .Z(n1258) );
  XOR U1476 ( .A(b[9]), .B(a[16]), .Z(n1360) );
  NAND U1477 ( .A(n19598), .B(n1360), .Z(n1257) );
  NAND U1478 ( .A(n1258), .B(n1257), .Z(n1363) );
  XOR U1479 ( .A(n1364), .B(n1363), .Z(n1366) );
  XOR U1480 ( .A(n1365), .B(n1366), .Z(n1376) );
  NANDN U1481 ( .A(n1260), .B(n1259), .Z(n1264) );
  OR U1482 ( .A(n1262), .B(n1261), .Z(n1263) );
  AND U1483 ( .A(n1264), .B(n1263), .Z(n1375) );
  XNOR U1484 ( .A(n1376), .B(n1375), .Z(n1377) );
  NANDN U1485 ( .A(n1266), .B(n1265), .Z(n1270) );
  NANDN U1486 ( .A(n1268), .B(n1267), .Z(n1269) );
  NAND U1487 ( .A(n1270), .B(n1269), .Z(n1378) );
  XNOR U1488 ( .A(n1377), .B(n1378), .Z(n1324) );
  NANDN U1489 ( .A(n1272), .B(n1271), .Z(n1276) );
  NANDN U1490 ( .A(n1274), .B(n1273), .Z(n1275) );
  AND U1491 ( .A(n1276), .B(n1275), .Z(n1350) );
  NAND U1492 ( .A(n19808), .B(n1277), .Z(n1279) );
  XOR U1493 ( .A(b[13]), .B(a[12]), .Z(n1336) );
  NAND U1494 ( .A(n19768), .B(n1336), .Z(n1278) );
  AND U1495 ( .A(n1279), .B(n1278), .Z(n1328) );
  AND U1496 ( .A(b[15]), .B(a[8]), .Z(n1327) );
  XNOR U1497 ( .A(n1328), .B(n1327), .Z(n1329) );
  NAND U1498 ( .A(b[0]), .B(a[24]), .Z(n1280) );
  XNOR U1499 ( .A(b[1]), .B(n1280), .Z(n1282) );
  NANDN U1500 ( .A(b[0]), .B(a[23]), .Z(n1281) );
  NAND U1501 ( .A(n1282), .B(n1281), .Z(n1330) );
  XNOR U1502 ( .A(n1329), .B(n1330), .Z(n1348) );
  NAND U1503 ( .A(n33), .B(n1283), .Z(n1285) );
  XOR U1504 ( .A(b[5]), .B(a[20]), .Z(n1339) );
  NAND U1505 ( .A(n19342), .B(n1339), .Z(n1284) );
  AND U1506 ( .A(n1285), .B(n1284), .Z(n1372) );
  NAND U1507 ( .A(n34), .B(n1286), .Z(n1288) );
  XOR U1508 ( .A(b[7]), .B(a[18]), .Z(n1342) );
  NAND U1509 ( .A(n19486), .B(n1342), .Z(n1287) );
  AND U1510 ( .A(n1288), .B(n1287), .Z(n1370) );
  NAND U1511 ( .A(n31), .B(n1289), .Z(n1291) );
  XOR U1512 ( .A(b[3]), .B(a[22]), .Z(n1345) );
  NAND U1513 ( .A(n32), .B(n1345), .Z(n1290) );
  NAND U1514 ( .A(n1291), .B(n1290), .Z(n1369) );
  XNOR U1515 ( .A(n1370), .B(n1369), .Z(n1371) );
  XOR U1516 ( .A(n1372), .B(n1371), .Z(n1349) );
  XOR U1517 ( .A(n1348), .B(n1349), .Z(n1351) );
  XOR U1518 ( .A(n1350), .B(n1351), .Z(n1322) );
  NANDN U1519 ( .A(n1293), .B(n1292), .Z(n1297) );
  OR U1520 ( .A(n1295), .B(n1294), .Z(n1296) );
  AND U1521 ( .A(n1297), .B(n1296), .Z(n1321) );
  XNOR U1522 ( .A(n1322), .B(n1321), .Z(n1323) );
  XOR U1523 ( .A(n1324), .B(n1323), .Z(n1382) );
  NANDN U1524 ( .A(n1299), .B(n1298), .Z(n1303) );
  NANDN U1525 ( .A(n1301), .B(n1300), .Z(n1302) );
  AND U1526 ( .A(n1303), .B(n1302), .Z(n1381) );
  XNOR U1527 ( .A(n1382), .B(n1381), .Z(n1383) );
  XOR U1528 ( .A(n1384), .B(n1383), .Z(n1316) );
  NANDN U1529 ( .A(n1305), .B(n1304), .Z(n1309) );
  NAND U1530 ( .A(n1307), .B(n1306), .Z(n1308) );
  AND U1531 ( .A(n1309), .B(n1308), .Z(n1315) );
  XNOR U1532 ( .A(n1316), .B(n1315), .Z(n1317) );
  XNOR U1533 ( .A(n1318), .B(n1317), .Z(n1387) );
  XNOR U1534 ( .A(sreg[264]), .B(n1387), .Z(n1389) );
  NANDN U1535 ( .A(sreg[263]), .B(n1310), .Z(n1314) );
  NAND U1536 ( .A(n1312), .B(n1311), .Z(n1313) );
  NAND U1537 ( .A(n1314), .B(n1313), .Z(n1388) );
  XNOR U1538 ( .A(n1389), .B(n1388), .Z(c[264]) );
  NANDN U1539 ( .A(n1316), .B(n1315), .Z(n1320) );
  NANDN U1540 ( .A(n1318), .B(n1317), .Z(n1319) );
  AND U1541 ( .A(n1320), .B(n1319), .Z(n1395) );
  NANDN U1542 ( .A(n1322), .B(n1321), .Z(n1326) );
  NAND U1543 ( .A(n1324), .B(n1323), .Z(n1325) );
  AND U1544 ( .A(n1326), .B(n1325), .Z(n1461) );
  NANDN U1545 ( .A(n1328), .B(n1327), .Z(n1332) );
  NANDN U1546 ( .A(n1330), .B(n1329), .Z(n1331) );
  AND U1547 ( .A(n1332), .B(n1331), .Z(n1427) );
  NAND U1548 ( .A(b[0]), .B(a[25]), .Z(n1333) );
  XNOR U1549 ( .A(b[1]), .B(n1333), .Z(n1335) );
  NANDN U1550 ( .A(b[0]), .B(a[24]), .Z(n1334) );
  NAND U1551 ( .A(n1335), .B(n1334), .Z(n1407) );
  NAND U1552 ( .A(n19808), .B(n1336), .Z(n1338) );
  XOR U1553 ( .A(b[13]), .B(a[13]), .Z(n1410) );
  NAND U1554 ( .A(n19768), .B(n1410), .Z(n1337) );
  AND U1555 ( .A(n1338), .B(n1337), .Z(n1405) );
  AND U1556 ( .A(b[15]), .B(a[9]), .Z(n1404) );
  XNOR U1557 ( .A(n1405), .B(n1404), .Z(n1406) );
  XNOR U1558 ( .A(n1407), .B(n1406), .Z(n1425) );
  NAND U1559 ( .A(n33), .B(n1339), .Z(n1341) );
  XOR U1560 ( .A(b[5]), .B(a[21]), .Z(n1416) );
  NAND U1561 ( .A(n19342), .B(n1416), .Z(n1340) );
  AND U1562 ( .A(n1341), .B(n1340), .Z(n1449) );
  NAND U1563 ( .A(n34), .B(n1342), .Z(n1344) );
  XOR U1564 ( .A(b[7]), .B(a[19]), .Z(n1419) );
  NAND U1565 ( .A(n19486), .B(n1419), .Z(n1343) );
  AND U1566 ( .A(n1344), .B(n1343), .Z(n1447) );
  NAND U1567 ( .A(n31), .B(n1345), .Z(n1347) );
  XOR U1568 ( .A(b[3]), .B(a[23]), .Z(n1422) );
  NAND U1569 ( .A(n32), .B(n1422), .Z(n1346) );
  NAND U1570 ( .A(n1347), .B(n1346), .Z(n1446) );
  XNOR U1571 ( .A(n1447), .B(n1446), .Z(n1448) );
  XOR U1572 ( .A(n1449), .B(n1448), .Z(n1426) );
  XOR U1573 ( .A(n1425), .B(n1426), .Z(n1428) );
  XOR U1574 ( .A(n1427), .B(n1428), .Z(n1399) );
  NANDN U1575 ( .A(n1349), .B(n1348), .Z(n1353) );
  OR U1576 ( .A(n1351), .B(n1350), .Z(n1352) );
  AND U1577 ( .A(n1353), .B(n1352), .Z(n1398) );
  XNOR U1578 ( .A(n1399), .B(n1398), .Z(n1401) );
  NAND U1579 ( .A(n1354), .B(n19724), .Z(n1356) );
  XOR U1580 ( .A(b[11]), .B(a[15]), .Z(n1431) );
  NAND U1581 ( .A(n19692), .B(n1431), .Z(n1355) );
  AND U1582 ( .A(n1356), .B(n1355), .Z(n1442) );
  NAND U1583 ( .A(n19838), .B(n1357), .Z(n1359) );
  XOR U1584 ( .A(b[15]), .B(a[11]), .Z(n1434) );
  NAND U1585 ( .A(n19805), .B(n1434), .Z(n1358) );
  AND U1586 ( .A(n1359), .B(n1358), .Z(n1441) );
  NAND U1587 ( .A(n35), .B(n1360), .Z(n1362) );
  XOR U1588 ( .A(b[9]), .B(a[17]), .Z(n1437) );
  NAND U1589 ( .A(n19598), .B(n1437), .Z(n1361) );
  NAND U1590 ( .A(n1362), .B(n1361), .Z(n1440) );
  XOR U1591 ( .A(n1441), .B(n1440), .Z(n1443) );
  XOR U1592 ( .A(n1442), .B(n1443), .Z(n1453) );
  NANDN U1593 ( .A(n1364), .B(n1363), .Z(n1368) );
  OR U1594 ( .A(n1366), .B(n1365), .Z(n1367) );
  AND U1595 ( .A(n1368), .B(n1367), .Z(n1452) );
  XNOR U1596 ( .A(n1453), .B(n1452), .Z(n1454) );
  NANDN U1597 ( .A(n1370), .B(n1369), .Z(n1374) );
  NANDN U1598 ( .A(n1372), .B(n1371), .Z(n1373) );
  NAND U1599 ( .A(n1374), .B(n1373), .Z(n1455) );
  XNOR U1600 ( .A(n1454), .B(n1455), .Z(n1400) );
  XOR U1601 ( .A(n1401), .B(n1400), .Z(n1459) );
  NANDN U1602 ( .A(n1376), .B(n1375), .Z(n1380) );
  NANDN U1603 ( .A(n1378), .B(n1377), .Z(n1379) );
  AND U1604 ( .A(n1380), .B(n1379), .Z(n1458) );
  XNOR U1605 ( .A(n1459), .B(n1458), .Z(n1460) );
  XOR U1606 ( .A(n1461), .B(n1460), .Z(n1393) );
  NANDN U1607 ( .A(n1382), .B(n1381), .Z(n1386) );
  NAND U1608 ( .A(n1384), .B(n1383), .Z(n1385) );
  AND U1609 ( .A(n1386), .B(n1385), .Z(n1392) );
  XNOR U1610 ( .A(n1393), .B(n1392), .Z(n1394) );
  XNOR U1611 ( .A(n1395), .B(n1394), .Z(n1464) );
  XNOR U1612 ( .A(sreg[265]), .B(n1464), .Z(n1466) );
  NANDN U1613 ( .A(sreg[264]), .B(n1387), .Z(n1391) );
  NAND U1614 ( .A(n1389), .B(n1388), .Z(n1390) );
  NAND U1615 ( .A(n1391), .B(n1390), .Z(n1465) );
  XNOR U1616 ( .A(n1466), .B(n1465), .Z(c[265]) );
  NANDN U1617 ( .A(n1393), .B(n1392), .Z(n1397) );
  NANDN U1618 ( .A(n1395), .B(n1394), .Z(n1396) );
  AND U1619 ( .A(n1397), .B(n1396), .Z(n1472) );
  NANDN U1620 ( .A(n1399), .B(n1398), .Z(n1403) );
  NAND U1621 ( .A(n1401), .B(n1400), .Z(n1402) );
  AND U1622 ( .A(n1403), .B(n1402), .Z(n1538) );
  NANDN U1623 ( .A(n1405), .B(n1404), .Z(n1409) );
  NANDN U1624 ( .A(n1407), .B(n1406), .Z(n1408) );
  AND U1625 ( .A(n1409), .B(n1408), .Z(n1504) );
  NAND U1626 ( .A(n19808), .B(n1410), .Z(n1412) );
  XOR U1627 ( .A(b[13]), .B(a[14]), .Z(n1490) );
  NAND U1628 ( .A(n19768), .B(n1490), .Z(n1411) );
  AND U1629 ( .A(n1412), .B(n1411), .Z(n1482) );
  AND U1630 ( .A(b[15]), .B(a[10]), .Z(n1481) );
  XNOR U1631 ( .A(n1482), .B(n1481), .Z(n1483) );
  NAND U1632 ( .A(b[0]), .B(a[26]), .Z(n1413) );
  XNOR U1633 ( .A(b[1]), .B(n1413), .Z(n1415) );
  NANDN U1634 ( .A(b[0]), .B(a[25]), .Z(n1414) );
  NAND U1635 ( .A(n1415), .B(n1414), .Z(n1484) );
  XNOR U1636 ( .A(n1483), .B(n1484), .Z(n1502) );
  NAND U1637 ( .A(n33), .B(n1416), .Z(n1418) );
  XOR U1638 ( .A(b[5]), .B(a[22]), .Z(n1493) );
  NAND U1639 ( .A(n19342), .B(n1493), .Z(n1417) );
  AND U1640 ( .A(n1418), .B(n1417), .Z(n1526) );
  NAND U1641 ( .A(n34), .B(n1419), .Z(n1421) );
  XOR U1642 ( .A(b[7]), .B(a[20]), .Z(n1496) );
  NAND U1643 ( .A(n19486), .B(n1496), .Z(n1420) );
  AND U1644 ( .A(n1421), .B(n1420), .Z(n1524) );
  NAND U1645 ( .A(n31), .B(n1422), .Z(n1424) );
  XOR U1646 ( .A(b[3]), .B(a[24]), .Z(n1499) );
  NAND U1647 ( .A(n32), .B(n1499), .Z(n1423) );
  NAND U1648 ( .A(n1424), .B(n1423), .Z(n1523) );
  XNOR U1649 ( .A(n1524), .B(n1523), .Z(n1525) );
  XOR U1650 ( .A(n1526), .B(n1525), .Z(n1503) );
  XOR U1651 ( .A(n1502), .B(n1503), .Z(n1505) );
  XOR U1652 ( .A(n1504), .B(n1505), .Z(n1476) );
  NANDN U1653 ( .A(n1426), .B(n1425), .Z(n1430) );
  OR U1654 ( .A(n1428), .B(n1427), .Z(n1429) );
  AND U1655 ( .A(n1430), .B(n1429), .Z(n1475) );
  XNOR U1656 ( .A(n1476), .B(n1475), .Z(n1478) );
  NAND U1657 ( .A(n1431), .B(n19724), .Z(n1433) );
  XOR U1658 ( .A(b[11]), .B(a[16]), .Z(n1508) );
  NAND U1659 ( .A(n19692), .B(n1508), .Z(n1432) );
  AND U1660 ( .A(n1433), .B(n1432), .Z(n1519) );
  NAND U1661 ( .A(n19838), .B(n1434), .Z(n1436) );
  XOR U1662 ( .A(b[15]), .B(a[12]), .Z(n1511) );
  NAND U1663 ( .A(n19805), .B(n1511), .Z(n1435) );
  AND U1664 ( .A(n1436), .B(n1435), .Z(n1518) );
  NAND U1665 ( .A(n35), .B(n1437), .Z(n1439) );
  XOR U1666 ( .A(b[9]), .B(a[18]), .Z(n1514) );
  NAND U1667 ( .A(n19598), .B(n1514), .Z(n1438) );
  NAND U1668 ( .A(n1439), .B(n1438), .Z(n1517) );
  XOR U1669 ( .A(n1518), .B(n1517), .Z(n1520) );
  XOR U1670 ( .A(n1519), .B(n1520), .Z(n1530) );
  NANDN U1671 ( .A(n1441), .B(n1440), .Z(n1445) );
  OR U1672 ( .A(n1443), .B(n1442), .Z(n1444) );
  AND U1673 ( .A(n1445), .B(n1444), .Z(n1529) );
  XNOR U1674 ( .A(n1530), .B(n1529), .Z(n1531) );
  NANDN U1675 ( .A(n1447), .B(n1446), .Z(n1451) );
  NANDN U1676 ( .A(n1449), .B(n1448), .Z(n1450) );
  NAND U1677 ( .A(n1451), .B(n1450), .Z(n1532) );
  XNOR U1678 ( .A(n1531), .B(n1532), .Z(n1477) );
  XOR U1679 ( .A(n1478), .B(n1477), .Z(n1536) );
  NANDN U1680 ( .A(n1453), .B(n1452), .Z(n1457) );
  NANDN U1681 ( .A(n1455), .B(n1454), .Z(n1456) );
  AND U1682 ( .A(n1457), .B(n1456), .Z(n1535) );
  XNOR U1683 ( .A(n1536), .B(n1535), .Z(n1537) );
  XOR U1684 ( .A(n1538), .B(n1537), .Z(n1470) );
  NANDN U1685 ( .A(n1459), .B(n1458), .Z(n1463) );
  NAND U1686 ( .A(n1461), .B(n1460), .Z(n1462) );
  AND U1687 ( .A(n1463), .B(n1462), .Z(n1469) );
  XNOR U1688 ( .A(n1470), .B(n1469), .Z(n1471) );
  XNOR U1689 ( .A(n1472), .B(n1471), .Z(n1541) );
  XNOR U1690 ( .A(sreg[266]), .B(n1541), .Z(n1543) );
  NANDN U1691 ( .A(sreg[265]), .B(n1464), .Z(n1468) );
  NAND U1692 ( .A(n1466), .B(n1465), .Z(n1467) );
  NAND U1693 ( .A(n1468), .B(n1467), .Z(n1542) );
  XNOR U1694 ( .A(n1543), .B(n1542), .Z(c[266]) );
  NANDN U1695 ( .A(n1470), .B(n1469), .Z(n1474) );
  NANDN U1696 ( .A(n1472), .B(n1471), .Z(n1473) );
  AND U1697 ( .A(n1474), .B(n1473), .Z(n1549) );
  NANDN U1698 ( .A(n1476), .B(n1475), .Z(n1480) );
  NAND U1699 ( .A(n1478), .B(n1477), .Z(n1479) );
  AND U1700 ( .A(n1480), .B(n1479), .Z(n1615) );
  NANDN U1701 ( .A(n1482), .B(n1481), .Z(n1486) );
  NANDN U1702 ( .A(n1484), .B(n1483), .Z(n1485) );
  AND U1703 ( .A(n1486), .B(n1485), .Z(n1581) );
  NAND U1704 ( .A(b[0]), .B(a[27]), .Z(n1487) );
  XNOR U1705 ( .A(b[1]), .B(n1487), .Z(n1489) );
  NANDN U1706 ( .A(b[0]), .B(a[26]), .Z(n1488) );
  NAND U1707 ( .A(n1489), .B(n1488), .Z(n1561) );
  NAND U1708 ( .A(n19808), .B(n1490), .Z(n1492) );
  XOR U1709 ( .A(b[13]), .B(a[15]), .Z(n1567) );
  NAND U1710 ( .A(n19768), .B(n1567), .Z(n1491) );
  AND U1711 ( .A(n1492), .B(n1491), .Z(n1559) );
  AND U1712 ( .A(b[15]), .B(a[11]), .Z(n1558) );
  XNOR U1713 ( .A(n1559), .B(n1558), .Z(n1560) );
  XNOR U1714 ( .A(n1561), .B(n1560), .Z(n1579) );
  NAND U1715 ( .A(n33), .B(n1493), .Z(n1495) );
  XOR U1716 ( .A(b[5]), .B(a[23]), .Z(n1570) );
  NAND U1717 ( .A(n19342), .B(n1570), .Z(n1494) );
  AND U1718 ( .A(n1495), .B(n1494), .Z(n1603) );
  NAND U1719 ( .A(n34), .B(n1496), .Z(n1498) );
  XOR U1720 ( .A(b[7]), .B(a[21]), .Z(n1573) );
  NAND U1721 ( .A(n19486), .B(n1573), .Z(n1497) );
  AND U1722 ( .A(n1498), .B(n1497), .Z(n1601) );
  NAND U1723 ( .A(n31), .B(n1499), .Z(n1501) );
  XOR U1724 ( .A(b[3]), .B(a[25]), .Z(n1576) );
  NAND U1725 ( .A(n32), .B(n1576), .Z(n1500) );
  NAND U1726 ( .A(n1501), .B(n1500), .Z(n1600) );
  XNOR U1727 ( .A(n1601), .B(n1600), .Z(n1602) );
  XOR U1728 ( .A(n1603), .B(n1602), .Z(n1580) );
  XOR U1729 ( .A(n1579), .B(n1580), .Z(n1582) );
  XOR U1730 ( .A(n1581), .B(n1582), .Z(n1553) );
  NANDN U1731 ( .A(n1503), .B(n1502), .Z(n1507) );
  OR U1732 ( .A(n1505), .B(n1504), .Z(n1506) );
  AND U1733 ( .A(n1507), .B(n1506), .Z(n1552) );
  XNOR U1734 ( .A(n1553), .B(n1552), .Z(n1555) );
  NAND U1735 ( .A(n1508), .B(n19724), .Z(n1510) );
  XOR U1736 ( .A(b[11]), .B(a[17]), .Z(n1585) );
  NAND U1737 ( .A(n19692), .B(n1585), .Z(n1509) );
  AND U1738 ( .A(n1510), .B(n1509), .Z(n1596) );
  NAND U1739 ( .A(n19838), .B(n1511), .Z(n1513) );
  XOR U1740 ( .A(b[15]), .B(a[13]), .Z(n1588) );
  NAND U1741 ( .A(n19805), .B(n1588), .Z(n1512) );
  AND U1742 ( .A(n1513), .B(n1512), .Z(n1595) );
  NAND U1743 ( .A(n35), .B(n1514), .Z(n1516) );
  XOR U1744 ( .A(b[9]), .B(a[19]), .Z(n1591) );
  NAND U1745 ( .A(n19598), .B(n1591), .Z(n1515) );
  NAND U1746 ( .A(n1516), .B(n1515), .Z(n1594) );
  XOR U1747 ( .A(n1595), .B(n1594), .Z(n1597) );
  XOR U1748 ( .A(n1596), .B(n1597), .Z(n1607) );
  NANDN U1749 ( .A(n1518), .B(n1517), .Z(n1522) );
  OR U1750 ( .A(n1520), .B(n1519), .Z(n1521) );
  AND U1751 ( .A(n1522), .B(n1521), .Z(n1606) );
  XNOR U1752 ( .A(n1607), .B(n1606), .Z(n1608) );
  NANDN U1753 ( .A(n1524), .B(n1523), .Z(n1528) );
  NANDN U1754 ( .A(n1526), .B(n1525), .Z(n1527) );
  NAND U1755 ( .A(n1528), .B(n1527), .Z(n1609) );
  XNOR U1756 ( .A(n1608), .B(n1609), .Z(n1554) );
  XOR U1757 ( .A(n1555), .B(n1554), .Z(n1613) );
  NANDN U1758 ( .A(n1530), .B(n1529), .Z(n1534) );
  NANDN U1759 ( .A(n1532), .B(n1531), .Z(n1533) );
  AND U1760 ( .A(n1534), .B(n1533), .Z(n1612) );
  XNOR U1761 ( .A(n1613), .B(n1612), .Z(n1614) );
  XOR U1762 ( .A(n1615), .B(n1614), .Z(n1547) );
  NANDN U1763 ( .A(n1536), .B(n1535), .Z(n1540) );
  NAND U1764 ( .A(n1538), .B(n1537), .Z(n1539) );
  AND U1765 ( .A(n1540), .B(n1539), .Z(n1546) );
  XNOR U1766 ( .A(n1547), .B(n1546), .Z(n1548) );
  XNOR U1767 ( .A(n1549), .B(n1548), .Z(n1618) );
  XNOR U1768 ( .A(sreg[267]), .B(n1618), .Z(n1620) );
  NANDN U1769 ( .A(sreg[266]), .B(n1541), .Z(n1545) );
  NAND U1770 ( .A(n1543), .B(n1542), .Z(n1544) );
  NAND U1771 ( .A(n1545), .B(n1544), .Z(n1619) );
  XNOR U1772 ( .A(n1620), .B(n1619), .Z(c[267]) );
  NANDN U1773 ( .A(n1547), .B(n1546), .Z(n1551) );
  NANDN U1774 ( .A(n1549), .B(n1548), .Z(n1550) );
  AND U1775 ( .A(n1551), .B(n1550), .Z(n1626) );
  NANDN U1776 ( .A(n1553), .B(n1552), .Z(n1557) );
  NAND U1777 ( .A(n1555), .B(n1554), .Z(n1556) );
  AND U1778 ( .A(n1557), .B(n1556), .Z(n1692) );
  NANDN U1779 ( .A(n1559), .B(n1558), .Z(n1563) );
  NANDN U1780 ( .A(n1561), .B(n1560), .Z(n1562) );
  AND U1781 ( .A(n1563), .B(n1562), .Z(n1658) );
  NAND U1782 ( .A(b[0]), .B(a[28]), .Z(n1564) );
  XNOR U1783 ( .A(b[1]), .B(n1564), .Z(n1566) );
  NANDN U1784 ( .A(b[0]), .B(a[27]), .Z(n1565) );
  NAND U1785 ( .A(n1566), .B(n1565), .Z(n1638) );
  NAND U1786 ( .A(n19808), .B(n1567), .Z(n1569) );
  XOR U1787 ( .A(b[13]), .B(a[16]), .Z(n1644) );
  NAND U1788 ( .A(n19768), .B(n1644), .Z(n1568) );
  AND U1789 ( .A(n1569), .B(n1568), .Z(n1636) );
  AND U1790 ( .A(b[15]), .B(a[12]), .Z(n1635) );
  XNOR U1791 ( .A(n1636), .B(n1635), .Z(n1637) );
  XNOR U1792 ( .A(n1638), .B(n1637), .Z(n1656) );
  NAND U1793 ( .A(n33), .B(n1570), .Z(n1572) );
  XOR U1794 ( .A(b[5]), .B(a[24]), .Z(n1647) );
  NAND U1795 ( .A(n19342), .B(n1647), .Z(n1571) );
  AND U1796 ( .A(n1572), .B(n1571), .Z(n1680) );
  NAND U1797 ( .A(n34), .B(n1573), .Z(n1575) );
  XOR U1798 ( .A(b[7]), .B(a[22]), .Z(n1650) );
  NAND U1799 ( .A(n19486), .B(n1650), .Z(n1574) );
  AND U1800 ( .A(n1575), .B(n1574), .Z(n1678) );
  NAND U1801 ( .A(n31), .B(n1576), .Z(n1578) );
  XOR U1802 ( .A(b[3]), .B(a[26]), .Z(n1653) );
  NAND U1803 ( .A(n32), .B(n1653), .Z(n1577) );
  NAND U1804 ( .A(n1578), .B(n1577), .Z(n1677) );
  XNOR U1805 ( .A(n1678), .B(n1677), .Z(n1679) );
  XOR U1806 ( .A(n1680), .B(n1679), .Z(n1657) );
  XOR U1807 ( .A(n1656), .B(n1657), .Z(n1659) );
  XOR U1808 ( .A(n1658), .B(n1659), .Z(n1630) );
  NANDN U1809 ( .A(n1580), .B(n1579), .Z(n1584) );
  OR U1810 ( .A(n1582), .B(n1581), .Z(n1583) );
  AND U1811 ( .A(n1584), .B(n1583), .Z(n1629) );
  XNOR U1812 ( .A(n1630), .B(n1629), .Z(n1632) );
  NAND U1813 ( .A(n1585), .B(n19724), .Z(n1587) );
  XOR U1814 ( .A(b[11]), .B(a[18]), .Z(n1662) );
  NAND U1815 ( .A(n19692), .B(n1662), .Z(n1586) );
  AND U1816 ( .A(n1587), .B(n1586), .Z(n1673) );
  NAND U1817 ( .A(n19838), .B(n1588), .Z(n1590) );
  XOR U1818 ( .A(b[15]), .B(a[14]), .Z(n1665) );
  NAND U1819 ( .A(n19805), .B(n1665), .Z(n1589) );
  AND U1820 ( .A(n1590), .B(n1589), .Z(n1672) );
  NAND U1821 ( .A(n35), .B(n1591), .Z(n1593) );
  XOR U1822 ( .A(b[9]), .B(a[20]), .Z(n1668) );
  NAND U1823 ( .A(n19598), .B(n1668), .Z(n1592) );
  NAND U1824 ( .A(n1593), .B(n1592), .Z(n1671) );
  XOR U1825 ( .A(n1672), .B(n1671), .Z(n1674) );
  XOR U1826 ( .A(n1673), .B(n1674), .Z(n1684) );
  NANDN U1827 ( .A(n1595), .B(n1594), .Z(n1599) );
  OR U1828 ( .A(n1597), .B(n1596), .Z(n1598) );
  AND U1829 ( .A(n1599), .B(n1598), .Z(n1683) );
  XNOR U1830 ( .A(n1684), .B(n1683), .Z(n1685) );
  NANDN U1831 ( .A(n1601), .B(n1600), .Z(n1605) );
  NANDN U1832 ( .A(n1603), .B(n1602), .Z(n1604) );
  NAND U1833 ( .A(n1605), .B(n1604), .Z(n1686) );
  XNOR U1834 ( .A(n1685), .B(n1686), .Z(n1631) );
  XOR U1835 ( .A(n1632), .B(n1631), .Z(n1690) );
  NANDN U1836 ( .A(n1607), .B(n1606), .Z(n1611) );
  NANDN U1837 ( .A(n1609), .B(n1608), .Z(n1610) );
  AND U1838 ( .A(n1611), .B(n1610), .Z(n1689) );
  XNOR U1839 ( .A(n1690), .B(n1689), .Z(n1691) );
  XOR U1840 ( .A(n1692), .B(n1691), .Z(n1624) );
  NANDN U1841 ( .A(n1613), .B(n1612), .Z(n1617) );
  NAND U1842 ( .A(n1615), .B(n1614), .Z(n1616) );
  AND U1843 ( .A(n1617), .B(n1616), .Z(n1623) );
  XNOR U1844 ( .A(n1624), .B(n1623), .Z(n1625) );
  XNOR U1845 ( .A(n1626), .B(n1625), .Z(n1695) );
  XNOR U1846 ( .A(sreg[268]), .B(n1695), .Z(n1697) );
  NANDN U1847 ( .A(sreg[267]), .B(n1618), .Z(n1622) );
  NAND U1848 ( .A(n1620), .B(n1619), .Z(n1621) );
  NAND U1849 ( .A(n1622), .B(n1621), .Z(n1696) );
  XNOR U1850 ( .A(n1697), .B(n1696), .Z(c[268]) );
  NANDN U1851 ( .A(n1624), .B(n1623), .Z(n1628) );
  NANDN U1852 ( .A(n1626), .B(n1625), .Z(n1627) );
  AND U1853 ( .A(n1628), .B(n1627), .Z(n1703) );
  NANDN U1854 ( .A(n1630), .B(n1629), .Z(n1634) );
  NAND U1855 ( .A(n1632), .B(n1631), .Z(n1633) );
  AND U1856 ( .A(n1634), .B(n1633), .Z(n1769) );
  NANDN U1857 ( .A(n1636), .B(n1635), .Z(n1640) );
  NANDN U1858 ( .A(n1638), .B(n1637), .Z(n1639) );
  AND U1859 ( .A(n1640), .B(n1639), .Z(n1735) );
  NAND U1860 ( .A(b[0]), .B(a[29]), .Z(n1641) );
  XNOR U1861 ( .A(b[1]), .B(n1641), .Z(n1643) );
  NANDN U1862 ( .A(b[0]), .B(a[28]), .Z(n1642) );
  NAND U1863 ( .A(n1643), .B(n1642), .Z(n1715) );
  NAND U1864 ( .A(n19808), .B(n1644), .Z(n1646) );
  XOR U1865 ( .A(b[13]), .B(a[17]), .Z(n1721) );
  NAND U1866 ( .A(n19768), .B(n1721), .Z(n1645) );
  AND U1867 ( .A(n1646), .B(n1645), .Z(n1713) );
  AND U1868 ( .A(b[15]), .B(a[13]), .Z(n1712) );
  XNOR U1869 ( .A(n1713), .B(n1712), .Z(n1714) );
  XNOR U1870 ( .A(n1715), .B(n1714), .Z(n1733) );
  NAND U1871 ( .A(n33), .B(n1647), .Z(n1649) );
  XOR U1872 ( .A(b[5]), .B(a[25]), .Z(n1724) );
  NAND U1873 ( .A(n19342), .B(n1724), .Z(n1648) );
  AND U1874 ( .A(n1649), .B(n1648), .Z(n1757) );
  NAND U1875 ( .A(n34), .B(n1650), .Z(n1652) );
  XOR U1876 ( .A(b[7]), .B(a[23]), .Z(n1727) );
  NAND U1877 ( .A(n19486), .B(n1727), .Z(n1651) );
  AND U1878 ( .A(n1652), .B(n1651), .Z(n1755) );
  NAND U1879 ( .A(n31), .B(n1653), .Z(n1655) );
  XOR U1880 ( .A(b[3]), .B(a[27]), .Z(n1730) );
  NAND U1881 ( .A(n32), .B(n1730), .Z(n1654) );
  NAND U1882 ( .A(n1655), .B(n1654), .Z(n1754) );
  XNOR U1883 ( .A(n1755), .B(n1754), .Z(n1756) );
  XOR U1884 ( .A(n1757), .B(n1756), .Z(n1734) );
  XOR U1885 ( .A(n1733), .B(n1734), .Z(n1736) );
  XOR U1886 ( .A(n1735), .B(n1736), .Z(n1707) );
  NANDN U1887 ( .A(n1657), .B(n1656), .Z(n1661) );
  OR U1888 ( .A(n1659), .B(n1658), .Z(n1660) );
  AND U1889 ( .A(n1661), .B(n1660), .Z(n1706) );
  XNOR U1890 ( .A(n1707), .B(n1706), .Z(n1709) );
  NAND U1891 ( .A(n1662), .B(n19724), .Z(n1664) );
  XOR U1892 ( .A(b[11]), .B(a[19]), .Z(n1739) );
  NAND U1893 ( .A(n19692), .B(n1739), .Z(n1663) );
  AND U1894 ( .A(n1664), .B(n1663), .Z(n1750) );
  NAND U1895 ( .A(n19838), .B(n1665), .Z(n1667) );
  XOR U1896 ( .A(b[15]), .B(a[15]), .Z(n1742) );
  NAND U1897 ( .A(n19805), .B(n1742), .Z(n1666) );
  AND U1898 ( .A(n1667), .B(n1666), .Z(n1749) );
  NAND U1899 ( .A(n35), .B(n1668), .Z(n1670) );
  XOR U1900 ( .A(b[9]), .B(a[21]), .Z(n1745) );
  NAND U1901 ( .A(n19598), .B(n1745), .Z(n1669) );
  NAND U1902 ( .A(n1670), .B(n1669), .Z(n1748) );
  XOR U1903 ( .A(n1749), .B(n1748), .Z(n1751) );
  XOR U1904 ( .A(n1750), .B(n1751), .Z(n1761) );
  NANDN U1905 ( .A(n1672), .B(n1671), .Z(n1676) );
  OR U1906 ( .A(n1674), .B(n1673), .Z(n1675) );
  AND U1907 ( .A(n1676), .B(n1675), .Z(n1760) );
  XNOR U1908 ( .A(n1761), .B(n1760), .Z(n1762) );
  NANDN U1909 ( .A(n1678), .B(n1677), .Z(n1682) );
  NANDN U1910 ( .A(n1680), .B(n1679), .Z(n1681) );
  NAND U1911 ( .A(n1682), .B(n1681), .Z(n1763) );
  XNOR U1912 ( .A(n1762), .B(n1763), .Z(n1708) );
  XOR U1913 ( .A(n1709), .B(n1708), .Z(n1767) );
  NANDN U1914 ( .A(n1684), .B(n1683), .Z(n1688) );
  NANDN U1915 ( .A(n1686), .B(n1685), .Z(n1687) );
  AND U1916 ( .A(n1688), .B(n1687), .Z(n1766) );
  XNOR U1917 ( .A(n1767), .B(n1766), .Z(n1768) );
  XOR U1918 ( .A(n1769), .B(n1768), .Z(n1701) );
  NANDN U1919 ( .A(n1690), .B(n1689), .Z(n1694) );
  NAND U1920 ( .A(n1692), .B(n1691), .Z(n1693) );
  AND U1921 ( .A(n1694), .B(n1693), .Z(n1700) );
  XNOR U1922 ( .A(n1701), .B(n1700), .Z(n1702) );
  XNOR U1923 ( .A(n1703), .B(n1702), .Z(n1772) );
  XNOR U1924 ( .A(sreg[269]), .B(n1772), .Z(n1774) );
  NANDN U1925 ( .A(sreg[268]), .B(n1695), .Z(n1699) );
  NAND U1926 ( .A(n1697), .B(n1696), .Z(n1698) );
  NAND U1927 ( .A(n1699), .B(n1698), .Z(n1773) );
  XNOR U1928 ( .A(n1774), .B(n1773), .Z(c[269]) );
  NANDN U1929 ( .A(n1701), .B(n1700), .Z(n1705) );
  NANDN U1930 ( .A(n1703), .B(n1702), .Z(n1704) );
  AND U1931 ( .A(n1705), .B(n1704), .Z(n1780) );
  NANDN U1932 ( .A(n1707), .B(n1706), .Z(n1711) );
  NAND U1933 ( .A(n1709), .B(n1708), .Z(n1710) );
  AND U1934 ( .A(n1711), .B(n1710), .Z(n1846) );
  NANDN U1935 ( .A(n1713), .B(n1712), .Z(n1717) );
  NANDN U1936 ( .A(n1715), .B(n1714), .Z(n1716) );
  AND U1937 ( .A(n1717), .B(n1716), .Z(n1812) );
  NAND U1938 ( .A(b[0]), .B(a[30]), .Z(n1718) );
  XNOR U1939 ( .A(b[1]), .B(n1718), .Z(n1720) );
  NANDN U1940 ( .A(b[0]), .B(a[29]), .Z(n1719) );
  NAND U1941 ( .A(n1720), .B(n1719), .Z(n1792) );
  NAND U1942 ( .A(n19808), .B(n1721), .Z(n1723) );
  XOR U1943 ( .A(b[13]), .B(a[18]), .Z(n1798) );
  NAND U1944 ( .A(n19768), .B(n1798), .Z(n1722) );
  AND U1945 ( .A(n1723), .B(n1722), .Z(n1790) );
  AND U1946 ( .A(b[15]), .B(a[14]), .Z(n1789) );
  XNOR U1947 ( .A(n1790), .B(n1789), .Z(n1791) );
  XNOR U1948 ( .A(n1792), .B(n1791), .Z(n1810) );
  NAND U1949 ( .A(n33), .B(n1724), .Z(n1726) );
  XOR U1950 ( .A(b[5]), .B(a[26]), .Z(n1801) );
  NAND U1951 ( .A(n19342), .B(n1801), .Z(n1725) );
  AND U1952 ( .A(n1726), .B(n1725), .Z(n1834) );
  NAND U1953 ( .A(n34), .B(n1727), .Z(n1729) );
  XOR U1954 ( .A(b[7]), .B(a[24]), .Z(n1804) );
  NAND U1955 ( .A(n19486), .B(n1804), .Z(n1728) );
  AND U1956 ( .A(n1729), .B(n1728), .Z(n1832) );
  NAND U1957 ( .A(n31), .B(n1730), .Z(n1732) );
  XOR U1958 ( .A(b[3]), .B(a[28]), .Z(n1807) );
  NAND U1959 ( .A(n32), .B(n1807), .Z(n1731) );
  NAND U1960 ( .A(n1732), .B(n1731), .Z(n1831) );
  XNOR U1961 ( .A(n1832), .B(n1831), .Z(n1833) );
  XOR U1962 ( .A(n1834), .B(n1833), .Z(n1811) );
  XOR U1963 ( .A(n1810), .B(n1811), .Z(n1813) );
  XOR U1964 ( .A(n1812), .B(n1813), .Z(n1784) );
  NANDN U1965 ( .A(n1734), .B(n1733), .Z(n1738) );
  OR U1966 ( .A(n1736), .B(n1735), .Z(n1737) );
  AND U1967 ( .A(n1738), .B(n1737), .Z(n1783) );
  XNOR U1968 ( .A(n1784), .B(n1783), .Z(n1786) );
  NAND U1969 ( .A(n1739), .B(n19724), .Z(n1741) );
  XOR U1970 ( .A(b[11]), .B(a[20]), .Z(n1816) );
  NAND U1971 ( .A(n19692), .B(n1816), .Z(n1740) );
  AND U1972 ( .A(n1741), .B(n1740), .Z(n1827) );
  NAND U1973 ( .A(n19838), .B(n1742), .Z(n1744) );
  XOR U1974 ( .A(b[15]), .B(a[16]), .Z(n1819) );
  NAND U1975 ( .A(n19805), .B(n1819), .Z(n1743) );
  AND U1976 ( .A(n1744), .B(n1743), .Z(n1826) );
  NAND U1977 ( .A(n35), .B(n1745), .Z(n1747) );
  XOR U1978 ( .A(b[9]), .B(a[22]), .Z(n1822) );
  NAND U1979 ( .A(n19598), .B(n1822), .Z(n1746) );
  NAND U1980 ( .A(n1747), .B(n1746), .Z(n1825) );
  XOR U1981 ( .A(n1826), .B(n1825), .Z(n1828) );
  XOR U1982 ( .A(n1827), .B(n1828), .Z(n1838) );
  NANDN U1983 ( .A(n1749), .B(n1748), .Z(n1753) );
  OR U1984 ( .A(n1751), .B(n1750), .Z(n1752) );
  AND U1985 ( .A(n1753), .B(n1752), .Z(n1837) );
  XNOR U1986 ( .A(n1838), .B(n1837), .Z(n1839) );
  NANDN U1987 ( .A(n1755), .B(n1754), .Z(n1759) );
  NANDN U1988 ( .A(n1757), .B(n1756), .Z(n1758) );
  NAND U1989 ( .A(n1759), .B(n1758), .Z(n1840) );
  XNOR U1990 ( .A(n1839), .B(n1840), .Z(n1785) );
  XOR U1991 ( .A(n1786), .B(n1785), .Z(n1844) );
  NANDN U1992 ( .A(n1761), .B(n1760), .Z(n1765) );
  NANDN U1993 ( .A(n1763), .B(n1762), .Z(n1764) );
  AND U1994 ( .A(n1765), .B(n1764), .Z(n1843) );
  XNOR U1995 ( .A(n1844), .B(n1843), .Z(n1845) );
  XOR U1996 ( .A(n1846), .B(n1845), .Z(n1778) );
  NANDN U1997 ( .A(n1767), .B(n1766), .Z(n1771) );
  NAND U1998 ( .A(n1769), .B(n1768), .Z(n1770) );
  AND U1999 ( .A(n1771), .B(n1770), .Z(n1777) );
  XNOR U2000 ( .A(n1778), .B(n1777), .Z(n1779) );
  XNOR U2001 ( .A(n1780), .B(n1779), .Z(n1849) );
  XNOR U2002 ( .A(sreg[270]), .B(n1849), .Z(n1851) );
  NANDN U2003 ( .A(sreg[269]), .B(n1772), .Z(n1776) );
  NAND U2004 ( .A(n1774), .B(n1773), .Z(n1775) );
  NAND U2005 ( .A(n1776), .B(n1775), .Z(n1850) );
  XNOR U2006 ( .A(n1851), .B(n1850), .Z(c[270]) );
  NANDN U2007 ( .A(n1778), .B(n1777), .Z(n1782) );
  NANDN U2008 ( .A(n1780), .B(n1779), .Z(n1781) );
  AND U2009 ( .A(n1782), .B(n1781), .Z(n1857) );
  NANDN U2010 ( .A(n1784), .B(n1783), .Z(n1788) );
  NAND U2011 ( .A(n1786), .B(n1785), .Z(n1787) );
  AND U2012 ( .A(n1788), .B(n1787), .Z(n1923) );
  NANDN U2013 ( .A(n1790), .B(n1789), .Z(n1794) );
  NANDN U2014 ( .A(n1792), .B(n1791), .Z(n1793) );
  AND U2015 ( .A(n1794), .B(n1793), .Z(n1889) );
  NAND U2016 ( .A(b[0]), .B(a[31]), .Z(n1795) );
  XNOR U2017 ( .A(b[1]), .B(n1795), .Z(n1797) );
  NANDN U2018 ( .A(b[0]), .B(a[30]), .Z(n1796) );
  NAND U2019 ( .A(n1797), .B(n1796), .Z(n1869) );
  NAND U2020 ( .A(n19808), .B(n1798), .Z(n1800) );
  XOR U2021 ( .A(b[13]), .B(a[19]), .Z(n1875) );
  NAND U2022 ( .A(n19768), .B(n1875), .Z(n1799) );
  AND U2023 ( .A(n1800), .B(n1799), .Z(n1867) );
  AND U2024 ( .A(b[15]), .B(a[15]), .Z(n1866) );
  XNOR U2025 ( .A(n1867), .B(n1866), .Z(n1868) );
  XNOR U2026 ( .A(n1869), .B(n1868), .Z(n1887) );
  NAND U2027 ( .A(n33), .B(n1801), .Z(n1803) );
  XOR U2028 ( .A(b[5]), .B(a[27]), .Z(n1878) );
  NAND U2029 ( .A(n19342), .B(n1878), .Z(n1802) );
  AND U2030 ( .A(n1803), .B(n1802), .Z(n1911) );
  NAND U2031 ( .A(n34), .B(n1804), .Z(n1806) );
  XOR U2032 ( .A(b[7]), .B(a[25]), .Z(n1881) );
  NAND U2033 ( .A(n19486), .B(n1881), .Z(n1805) );
  AND U2034 ( .A(n1806), .B(n1805), .Z(n1909) );
  NAND U2035 ( .A(n31), .B(n1807), .Z(n1809) );
  XOR U2036 ( .A(b[3]), .B(a[29]), .Z(n1884) );
  NAND U2037 ( .A(n32), .B(n1884), .Z(n1808) );
  NAND U2038 ( .A(n1809), .B(n1808), .Z(n1908) );
  XNOR U2039 ( .A(n1909), .B(n1908), .Z(n1910) );
  XOR U2040 ( .A(n1911), .B(n1910), .Z(n1888) );
  XOR U2041 ( .A(n1887), .B(n1888), .Z(n1890) );
  XOR U2042 ( .A(n1889), .B(n1890), .Z(n1861) );
  NANDN U2043 ( .A(n1811), .B(n1810), .Z(n1815) );
  OR U2044 ( .A(n1813), .B(n1812), .Z(n1814) );
  AND U2045 ( .A(n1815), .B(n1814), .Z(n1860) );
  XNOR U2046 ( .A(n1861), .B(n1860), .Z(n1863) );
  NAND U2047 ( .A(n1816), .B(n19724), .Z(n1818) );
  XOR U2048 ( .A(b[11]), .B(a[21]), .Z(n1893) );
  NAND U2049 ( .A(n19692), .B(n1893), .Z(n1817) );
  AND U2050 ( .A(n1818), .B(n1817), .Z(n1904) );
  NAND U2051 ( .A(n19838), .B(n1819), .Z(n1821) );
  XOR U2052 ( .A(b[15]), .B(a[17]), .Z(n1896) );
  NAND U2053 ( .A(n19805), .B(n1896), .Z(n1820) );
  AND U2054 ( .A(n1821), .B(n1820), .Z(n1903) );
  NAND U2055 ( .A(n35), .B(n1822), .Z(n1824) );
  XOR U2056 ( .A(b[9]), .B(a[23]), .Z(n1899) );
  NAND U2057 ( .A(n19598), .B(n1899), .Z(n1823) );
  NAND U2058 ( .A(n1824), .B(n1823), .Z(n1902) );
  XOR U2059 ( .A(n1903), .B(n1902), .Z(n1905) );
  XOR U2060 ( .A(n1904), .B(n1905), .Z(n1915) );
  NANDN U2061 ( .A(n1826), .B(n1825), .Z(n1830) );
  OR U2062 ( .A(n1828), .B(n1827), .Z(n1829) );
  AND U2063 ( .A(n1830), .B(n1829), .Z(n1914) );
  XNOR U2064 ( .A(n1915), .B(n1914), .Z(n1916) );
  NANDN U2065 ( .A(n1832), .B(n1831), .Z(n1836) );
  NANDN U2066 ( .A(n1834), .B(n1833), .Z(n1835) );
  NAND U2067 ( .A(n1836), .B(n1835), .Z(n1917) );
  XNOR U2068 ( .A(n1916), .B(n1917), .Z(n1862) );
  XOR U2069 ( .A(n1863), .B(n1862), .Z(n1921) );
  NANDN U2070 ( .A(n1838), .B(n1837), .Z(n1842) );
  NANDN U2071 ( .A(n1840), .B(n1839), .Z(n1841) );
  AND U2072 ( .A(n1842), .B(n1841), .Z(n1920) );
  XNOR U2073 ( .A(n1921), .B(n1920), .Z(n1922) );
  XOR U2074 ( .A(n1923), .B(n1922), .Z(n1855) );
  NANDN U2075 ( .A(n1844), .B(n1843), .Z(n1848) );
  NAND U2076 ( .A(n1846), .B(n1845), .Z(n1847) );
  AND U2077 ( .A(n1848), .B(n1847), .Z(n1854) );
  XNOR U2078 ( .A(n1855), .B(n1854), .Z(n1856) );
  XNOR U2079 ( .A(n1857), .B(n1856), .Z(n1926) );
  XNOR U2080 ( .A(sreg[271]), .B(n1926), .Z(n1928) );
  NANDN U2081 ( .A(sreg[270]), .B(n1849), .Z(n1853) );
  NAND U2082 ( .A(n1851), .B(n1850), .Z(n1852) );
  NAND U2083 ( .A(n1853), .B(n1852), .Z(n1927) );
  XNOR U2084 ( .A(n1928), .B(n1927), .Z(c[271]) );
  NANDN U2085 ( .A(n1855), .B(n1854), .Z(n1859) );
  NANDN U2086 ( .A(n1857), .B(n1856), .Z(n1858) );
  AND U2087 ( .A(n1859), .B(n1858), .Z(n1934) );
  NANDN U2088 ( .A(n1861), .B(n1860), .Z(n1865) );
  NAND U2089 ( .A(n1863), .B(n1862), .Z(n1864) );
  AND U2090 ( .A(n1865), .B(n1864), .Z(n2000) );
  NANDN U2091 ( .A(n1867), .B(n1866), .Z(n1871) );
  NANDN U2092 ( .A(n1869), .B(n1868), .Z(n1870) );
  AND U2093 ( .A(n1871), .B(n1870), .Z(n1966) );
  NAND U2094 ( .A(b[0]), .B(a[32]), .Z(n1872) );
  XNOR U2095 ( .A(b[1]), .B(n1872), .Z(n1874) );
  NANDN U2096 ( .A(b[0]), .B(a[31]), .Z(n1873) );
  NAND U2097 ( .A(n1874), .B(n1873), .Z(n1946) );
  NAND U2098 ( .A(n19808), .B(n1875), .Z(n1877) );
  XOR U2099 ( .A(b[13]), .B(a[20]), .Z(n1952) );
  NAND U2100 ( .A(n19768), .B(n1952), .Z(n1876) );
  AND U2101 ( .A(n1877), .B(n1876), .Z(n1944) );
  AND U2102 ( .A(b[15]), .B(a[16]), .Z(n1943) );
  XNOR U2103 ( .A(n1944), .B(n1943), .Z(n1945) );
  XNOR U2104 ( .A(n1946), .B(n1945), .Z(n1964) );
  NAND U2105 ( .A(n33), .B(n1878), .Z(n1880) );
  XOR U2106 ( .A(b[5]), .B(a[28]), .Z(n1955) );
  NAND U2107 ( .A(n19342), .B(n1955), .Z(n1879) );
  AND U2108 ( .A(n1880), .B(n1879), .Z(n1988) );
  NAND U2109 ( .A(n34), .B(n1881), .Z(n1883) );
  XOR U2110 ( .A(b[7]), .B(a[26]), .Z(n1958) );
  NAND U2111 ( .A(n19486), .B(n1958), .Z(n1882) );
  AND U2112 ( .A(n1883), .B(n1882), .Z(n1986) );
  NAND U2113 ( .A(n31), .B(n1884), .Z(n1886) );
  XOR U2114 ( .A(b[3]), .B(a[30]), .Z(n1961) );
  NAND U2115 ( .A(n32), .B(n1961), .Z(n1885) );
  NAND U2116 ( .A(n1886), .B(n1885), .Z(n1985) );
  XNOR U2117 ( .A(n1986), .B(n1985), .Z(n1987) );
  XOR U2118 ( .A(n1988), .B(n1987), .Z(n1965) );
  XOR U2119 ( .A(n1964), .B(n1965), .Z(n1967) );
  XOR U2120 ( .A(n1966), .B(n1967), .Z(n1938) );
  NANDN U2121 ( .A(n1888), .B(n1887), .Z(n1892) );
  OR U2122 ( .A(n1890), .B(n1889), .Z(n1891) );
  AND U2123 ( .A(n1892), .B(n1891), .Z(n1937) );
  XNOR U2124 ( .A(n1938), .B(n1937), .Z(n1940) );
  NAND U2125 ( .A(n1893), .B(n19724), .Z(n1895) );
  XOR U2126 ( .A(b[11]), .B(a[22]), .Z(n1970) );
  NAND U2127 ( .A(n19692), .B(n1970), .Z(n1894) );
  AND U2128 ( .A(n1895), .B(n1894), .Z(n1981) );
  NAND U2129 ( .A(n19838), .B(n1896), .Z(n1898) );
  XOR U2130 ( .A(b[15]), .B(a[18]), .Z(n1973) );
  NAND U2131 ( .A(n19805), .B(n1973), .Z(n1897) );
  AND U2132 ( .A(n1898), .B(n1897), .Z(n1980) );
  NAND U2133 ( .A(n35), .B(n1899), .Z(n1901) );
  XOR U2134 ( .A(b[9]), .B(a[24]), .Z(n1976) );
  NAND U2135 ( .A(n19598), .B(n1976), .Z(n1900) );
  NAND U2136 ( .A(n1901), .B(n1900), .Z(n1979) );
  XOR U2137 ( .A(n1980), .B(n1979), .Z(n1982) );
  XOR U2138 ( .A(n1981), .B(n1982), .Z(n1992) );
  NANDN U2139 ( .A(n1903), .B(n1902), .Z(n1907) );
  OR U2140 ( .A(n1905), .B(n1904), .Z(n1906) );
  AND U2141 ( .A(n1907), .B(n1906), .Z(n1991) );
  XNOR U2142 ( .A(n1992), .B(n1991), .Z(n1993) );
  NANDN U2143 ( .A(n1909), .B(n1908), .Z(n1913) );
  NANDN U2144 ( .A(n1911), .B(n1910), .Z(n1912) );
  NAND U2145 ( .A(n1913), .B(n1912), .Z(n1994) );
  XNOR U2146 ( .A(n1993), .B(n1994), .Z(n1939) );
  XOR U2147 ( .A(n1940), .B(n1939), .Z(n1998) );
  NANDN U2148 ( .A(n1915), .B(n1914), .Z(n1919) );
  NANDN U2149 ( .A(n1917), .B(n1916), .Z(n1918) );
  AND U2150 ( .A(n1919), .B(n1918), .Z(n1997) );
  XNOR U2151 ( .A(n1998), .B(n1997), .Z(n1999) );
  XOR U2152 ( .A(n2000), .B(n1999), .Z(n1932) );
  NANDN U2153 ( .A(n1921), .B(n1920), .Z(n1925) );
  NAND U2154 ( .A(n1923), .B(n1922), .Z(n1924) );
  AND U2155 ( .A(n1925), .B(n1924), .Z(n1931) );
  XNOR U2156 ( .A(n1932), .B(n1931), .Z(n1933) );
  XNOR U2157 ( .A(n1934), .B(n1933), .Z(n2003) );
  XNOR U2158 ( .A(sreg[272]), .B(n2003), .Z(n2005) );
  NANDN U2159 ( .A(sreg[271]), .B(n1926), .Z(n1930) );
  NAND U2160 ( .A(n1928), .B(n1927), .Z(n1929) );
  NAND U2161 ( .A(n1930), .B(n1929), .Z(n2004) );
  XNOR U2162 ( .A(n2005), .B(n2004), .Z(c[272]) );
  NANDN U2163 ( .A(n1932), .B(n1931), .Z(n1936) );
  NANDN U2164 ( .A(n1934), .B(n1933), .Z(n1935) );
  AND U2165 ( .A(n1936), .B(n1935), .Z(n2011) );
  NANDN U2166 ( .A(n1938), .B(n1937), .Z(n1942) );
  NAND U2167 ( .A(n1940), .B(n1939), .Z(n1941) );
  AND U2168 ( .A(n1942), .B(n1941), .Z(n2077) );
  NANDN U2169 ( .A(n1944), .B(n1943), .Z(n1948) );
  NANDN U2170 ( .A(n1946), .B(n1945), .Z(n1947) );
  AND U2171 ( .A(n1948), .B(n1947), .Z(n2043) );
  NAND U2172 ( .A(b[0]), .B(a[33]), .Z(n1949) );
  XNOR U2173 ( .A(b[1]), .B(n1949), .Z(n1951) );
  NANDN U2174 ( .A(b[0]), .B(a[32]), .Z(n1950) );
  NAND U2175 ( .A(n1951), .B(n1950), .Z(n2023) );
  NAND U2176 ( .A(n19808), .B(n1952), .Z(n1954) );
  XOR U2177 ( .A(b[13]), .B(a[21]), .Z(n2026) );
  NAND U2178 ( .A(n19768), .B(n2026), .Z(n1953) );
  AND U2179 ( .A(n1954), .B(n1953), .Z(n2021) );
  AND U2180 ( .A(b[15]), .B(a[17]), .Z(n2020) );
  XNOR U2181 ( .A(n2021), .B(n2020), .Z(n2022) );
  XNOR U2182 ( .A(n2023), .B(n2022), .Z(n2041) );
  NAND U2183 ( .A(n33), .B(n1955), .Z(n1957) );
  XOR U2184 ( .A(b[5]), .B(a[29]), .Z(n2032) );
  NAND U2185 ( .A(n19342), .B(n2032), .Z(n1956) );
  AND U2186 ( .A(n1957), .B(n1956), .Z(n2065) );
  NAND U2187 ( .A(n34), .B(n1958), .Z(n1960) );
  XOR U2188 ( .A(b[7]), .B(a[27]), .Z(n2035) );
  NAND U2189 ( .A(n19486), .B(n2035), .Z(n1959) );
  AND U2190 ( .A(n1960), .B(n1959), .Z(n2063) );
  NAND U2191 ( .A(n31), .B(n1961), .Z(n1963) );
  XOR U2192 ( .A(b[3]), .B(a[31]), .Z(n2038) );
  NAND U2193 ( .A(n32), .B(n2038), .Z(n1962) );
  NAND U2194 ( .A(n1963), .B(n1962), .Z(n2062) );
  XNOR U2195 ( .A(n2063), .B(n2062), .Z(n2064) );
  XOR U2196 ( .A(n2065), .B(n2064), .Z(n2042) );
  XOR U2197 ( .A(n2041), .B(n2042), .Z(n2044) );
  XOR U2198 ( .A(n2043), .B(n2044), .Z(n2015) );
  NANDN U2199 ( .A(n1965), .B(n1964), .Z(n1969) );
  OR U2200 ( .A(n1967), .B(n1966), .Z(n1968) );
  AND U2201 ( .A(n1969), .B(n1968), .Z(n2014) );
  XNOR U2202 ( .A(n2015), .B(n2014), .Z(n2017) );
  NAND U2203 ( .A(n1970), .B(n19724), .Z(n1972) );
  XOR U2204 ( .A(b[11]), .B(a[23]), .Z(n2047) );
  NAND U2205 ( .A(n19692), .B(n2047), .Z(n1971) );
  AND U2206 ( .A(n1972), .B(n1971), .Z(n2058) );
  NAND U2207 ( .A(n19838), .B(n1973), .Z(n1975) );
  XOR U2208 ( .A(b[15]), .B(a[19]), .Z(n2050) );
  NAND U2209 ( .A(n19805), .B(n2050), .Z(n1974) );
  AND U2210 ( .A(n1975), .B(n1974), .Z(n2057) );
  NAND U2211 ( .A(n35), .B(n1976), .Z(n1978) );
  XOR U2212 ( .A(b[9]), .B(a[25]), .Z(n2053) );
  NAND U2213 ( .A(n19598), .B(n2053), .Z(n1977) );
  NAND U2214 ( .A(n1978), .B(n1977), .Z(n2056) );
  XOR U2215 ( .A(n2057), .B(n2056), .Z(n2059) );
  XOR U2216 ( .A(n2058), .B(n2059), .Z(n2069) );
  NANDN U2217 ( .A(n1980), .B(n1979), .Z(n1984) );
  OR U2218 ( .A(n1982), .B(n1981), .Z(n1983) );
  AND U2219 ( .A(n1984), .B(n1983), .Z(n2068) );
  XNOR U2220 ( .A(n2069), .B(n2068), .Z(n2070) );
  NANDN U2221 ( .A(n1986), .B(n1985), .Z(n1990) );
  NANDN U2222 ( .A(n1988), .B(n1987), .Z(n1989) );
  NAND U2223 ( .A(n1990), .B(n1989), .Z(n2071) );
  XNOR U2224 ( .A(n2070), .B(n2071), .Z(n2016) );
  XOR U2225 ( .A(n2017), .B(n2016), .Z(n2075) );
  NANDN U2226 ( .A(n1992), .B(n1991), .Z(n1996) );
  NANDN U2227 ( .A(n1994), .B(n1993), .Z(n1995) );
  AND U2228 ( .A(n1996), .B(n1995), .Z(n2074) );
  XNOR U2229 ( .A(n2075), .B(n2074), .Z(n2076) );
  XOR U2230 ( .A(n2077), .B(n2076), .Z(n2009) );
  NANDN U2231 ( .A(n1998), .B(n1997), .Z(n2002) );
  NAND U2232 ( .A(n2000), .B(n1999), .Z(n2001) );
  AND U2233 ( .A(n2002), .B(n2001), .Z(n2008) );
  XNOR U2234 ( .A(n2009), .B(n2008), .Z(n2010) );
  XNOR U2235 ( .A(n2011), .B(n2010), .Z(n2080) );
  XNOR U2236 ( .A(sreg[273]), .B(n2080), .Z(n2082) );
  NANDN U2237 ( .A(sreg[272]), .B(n2003), .Z(n2007) );
  NAND U2238 ( .A(n2005), .B(n2004), .Z(n2006) );
  NAND U2239 ( .A(n2007), .B(n2006), .Z(n2081) );
  XNOR U2240 ( .A(n2082), .B(n2081), .Z(c[273]) );
  NANDN U2241 ( .A(n2009), .B(n2008), .Z(n2013) );
  NANDN U2242 ( .A(n2011), .B(n2010), .Z(n2012) );
  AND U2243 ( .A(n2013), .B(n2012), .Z(n2088) );
  NANDN U2244 ( .A(n2015), .B(n2014), .Z(n2019) );
  NAND U2245 ( .A(n2017), .B(n2016), .Z(n2018) );
  AND U2246 ( .A(n2019), .B(n2018), .Z(n2154) );
  NANDN U2247 ( .A(n2021), .B(n2020), .Z(n2025) );
  NANDN U2248 ( .A(n2023), .B(n2022), .Z(n2024) );
  AND U2249 ( .A(n2025), .B(n2024), .Z(n2120) );
  NAND U2250 ( .A(n19808), .B(n2026), .Z(n2028) );
  XOR U2251 ( .A(b[13]), .B(a[22]), .Z(n2106) );
  NAND U2252 ( .A(n19768), .B(n2106), .Z(n2027) );
  AND U2253 ( .A(n2028), .B(n2027), .Z(n2098) );
  AND U2254 ( .A(b[15]), .B(a[18]), .Z(n2097) );
  XNOR U2255 ( .A(n2098), .B(n2097), .Z(n2099) );
  NAND U2256 ( .A(b[0]), .B(a[34]), .Z(n2029) );
  XNOR U2257 ( .A(b[1]), .B(n2029), .Z(n2031) );
  NANDN U2258 ( .A(b[0]), .B(a[33]), .Z(n2030) );
  NAND U2259 ( .A(n2031), .B(n2030), .Z(n2100) );
  XNOR U2260 ( .A(n2099), .B(n2100), .Z(n2118) );
  NAND U2261 ( .A(n33), .B(n2032), .Z(n2034) );
  XOR U2262 ( .A(b[5]), .B(a[30]), .Z(n2109) );
  NAND U2263 ( .A(n19342), .B(n2109), .Z(n2033) );
  AND U2264 ( .A(n2034), .B(n2033), .Z(n2142) );
  NAND U2265 ( .A(n34), .B(n2035), .Z(n2037) );
  XOR U2266 ( .A(b[7]), .B(a[28]), .Z(n2112) );
  NAND U2267 ( .A(n19486), .B(n2112), .Z(n2036) );
  AND U2268 ( .A(n2037), .B(n2036), .Z(n2140) );
  NAND U2269 ( .A(n31), .B(n2038), .Z(n2040) );
  XOR U2270 ( .A(b[3]), .B(a[32]), .Z(n2115) );
  NAND U2271 ( .A(n32), .B(n2115), .Z(n2039) );
  NAND U2272 ( .A(n2040), .B(n2039), .Z(n2139) );
  XNOR U2273 ( .A(n2140), .B(n2139), .Z(n2141) );
  XOR U2274 ( .A(n2142), .B(n2141), .Z(n2119) );
  XOR U2275 ( .A(n2118), .B(n2119), .Z(n2121) );
  XOR U2276 ( .A(n2120), .B(n2121), .Z(n2092) );
  NANDN U2277 ( .A(n2042), .B(n2041), .Z(n2046) );
  OR U2278 ( .A(n2044), .B(n2043), .Z(n2045) );
  AND U2279 ( .A(n2046), .B(n2045), .Z(n2091) );
  XNOR U2280 ( .A(n2092), .B(n2091), .Z(n2094) );
  NAND U2281 ( .A(n2047), .B(n19724), .Z(n2049) );
  XOR U2282 ( .A(b[11]), .B(a[24]), .Z(n2124) );
  NAND U2283 ( .A(n19692), .B(n2124), .Z(n2048) );
  AND U2284 ( .A(n2049), .B(n2048), .Z(n2135) );
  NAND U2285 ( .A(n19838), .B(n2050), .Z(n2052) );
  XOR U2286 ( .A(b[15]), .B(a[20]), .Z(n2127) );
  NAND U2287 ( .A(n19805), .B(n2127), .Z(n2051) );
  AND U2288 ( .A(n2052), .B(n2051), .Z(n2134) );
  NAND U2289 ( .A(n35), .B(n2053), .Z(n2055) );
  XOR U2290 ( .A(b[9]), .B(a[26]), .Z(n2130) );
  NAND U2291 ( .A(n19598), .B(n2130), .Z(n2054) );
  NAND U2292 ( .A(n2055), .B(n2054), .Z(n2133) );
  XOR U2293 ( .A(n2134), .B(n2133), .Z(n2136) );
  XOR U2294 ( .A(n2135), .B(n2136), .Z(n2146) );
  NANDN U2295 ( .A(n2057), .B(n2056), .Z(n2061) );
  OR U2296 ( .A(n2059), .B(n2058), .Z(n2060) );
  AND U2297 ( .A(n2061), .B(n2060), .Z(n2145) );
  XNOR U2298 ( .A(n2146), .B(n2145), .Z(n2147) );
  NANDN U2299 ( .A(n2063), .B(n2062), .Z(n2067) );
  NANDN U2300 ( .A(n2065), .B(n2064), .Z(n2066) );
  NAND U2301 ( .A(n2067), .B(n2066), .Z(n2148) );
  XNOR U2302 ( .A(n2147), .B(n2148), .Z(n2093) );
  XOR U2303 ( .A(n2094), .B(n2093), .Z(n2152) );
  NANDN U2304 ( .A(n2069), .B(n2068), .Z(n2073) );
  NANDN U2305 ( .A(n2071), .B(n2070), .Z(n2072) );
  AND U2306 ( .A(n2073), .B(n2072), .Z(n2151) );
  XNOR U2307 ( .A(n2152), .B(n2151), .Z(n2153) );
  XOR U2308 ( .A(n2154), .B(n2153), .Z(n2086) );
  NANDN U2309 ( .A(n2075), .B(n2074), .Z(n2079) );
  NAND U2310 ( .A(n2077), .B(n2076), .Z(n2078) );
  AND U2311 ( .A(n2079), .B(n2078), .Z(n2085) );
  XNOR U2312 ( .A(n2086), .B(n2085), .Z(n2087) );
  XNOR U2313 ( .A(n2088), .B(n2087), .Z(n2157) );
  XNOR U2314 ( .A(sreg[274]), .B(n2157), .Z(n2159) );
  NANDN U2315 ( .A(sreg[273]), .B(n2080), .Z(n2084) );
  NAND U2316 ( .A(n2082), .B(n2081), .Z(n2083) );
  NAND U2317 ( .A(n2084), .B(n2083), .Z(n2158) );
  XNOR U2318 ( .A(n2159), .B(n2158), .Z(c[274]) );
  NANDN U2319 ( .A(n2086), .B(n2085), .Z(n2090) );
  NANDN U2320 ( .A(n2088), .B(n2087), .Z(n2089) );
  AND U2321 ( .A(n2090), .B(n2089), .Z(n2165) );
  NANDN U2322 ( .A(n2092), .B(n2091), .Z(n2096) );
  NAND U2323 ( .A(n2094), .B(n2093), .Z(n2095) );
  AND U2324 ( .A(n2096), .B(n2095), .Z(n2231) );
  NANDN U2325 ( .A(n2098), .B(n2097), .Z(n2102) );
  NANDN U2326 ( .A(n2100), .B(n2099), .Z(n2101) );
  AND U2327 ( .A(n2102), .B(n2101), .Z(n2197) );
  NAND U2328 ( .A(b[0]), .B(a[35]), .Z(n2103) );
  XNOR U2329 ( .A(b[1]), .B(n2103), .Z(n2105) );
  NANDN U2330 ( .A(b[0]), .B(a[34]), .Z(n2104) );
  NAND U2331 ( .A(n2105), .B(n2104), .Z(n2177) );
  NAND U2332 ( .A(n19808), .B(n2106), .Z(n2108) );
  XOR U2333 ( .A(b[13]), .B(a[23]), .Z(n2183) );
  NAND U2334 ( .A(n19768), .B(n2183), .Z(n2107) );
  AND U2335 ( .A(n2108), .B(n2107), .Z(n2175) );
  AND U2336 ( .A(b[15]), .B(a[19]), .Z(n2174) );
  XNOR U2337 ( .A(n2175), .B(n2174), .Z(n2176) );
  XNOR U2338 ( .A(n2177), .B(n2176), .Z(n2195) );
  NAND U2339 ( .A(n33), .B(n2109), .Z(n2111) );
  XOR U2340 ( .A(b[5]), .B(a[31]), .Z(n2186) );
  NAND U2341 ( .A(n19342), .B(n2186), .Z(n2110) );
  AND U2342 ( .A(n2111), .B(n2110), .Z(n2219) );
  NAND U2343 ( .A(n34), .B(n2112), .Z(n2114) );
  XOR U2344 ( .A(b[7]), .B(a[29]), .Z(n2189) );
  NAND U2345 ( .A(n19486), .B(n2189), .Z(n2113) );
  AND U2346 ( .A(n2114), .B(n2113), .Z(n2217) );
  NAND U2347 ( .A(n31), .B(n2115), .Z(n2117) );
  XOR U2348 ( .A(b[3]), .B(a[33]), .Z(n2192) );
  NAND U2349 ( .A(n32), .B(n2192), .Z(n2116) );
  NAND U2350 ( .A(n2117), .B(n2116), .Z(n2216) );
  XNOR U2351 ( .A(n2217), .B(n2216), .Z(n2218) );
  XOR U2352 ( .A(n2219), .B(n2218), .Z(n2196) );
  XOR U2353 ( .A(n2195), .B(n2196), .Z(n2198) );
  XOR U2354 ( .A(n2197), .B(n2198), .Z(n2169) );
  NANDN U2355 ( .A(n2119), .B(n2118), .Z(n2123) );
  OR U2356 ( .A(n2121), .B(n2120), .Z(n2122) );
  AND U2357 ( .A(n2123), .B(n2122), .Z(n2168) );
  XNOR U2358 ( .A(n2169), .B(n2168), .Z(n2171) );
  NAND U2359 ( .A(n2124), .B(n19724), .Z(n2126) );
  XOR U2360 ( .A(b[11]), .B(a[25]), .Z(n2201) );
  NAND U2361 ( .A(n19692), .B(n2201), .Z(n2125) );
  AND U2362 ( .A(n2126), .B(n2125), .Z(n2212) );
  NAND U2363 ( .A(n19838), .B(n2127), .Z(n2129) );
  XOR U2364 ( .A(b[15]), .B(a[21]), .Z(n2204) );
  NAND U2365 ( .A(n19805), .B(n2204), .Z(n2128) );
  AND U2366 ( .A(n2129), .B(n2128), .Z(n2211) );
  NAND U2367 ( .A(n35), .B(n2130), .Z(n2132) );
  XOR U2368 ( .A(b[9]), .B(a[27]), .Z(n2207) );
  NAND U2369 ( .A(n19598), .B(n2207), .Z(n2131) );
  NAND U2370 ( .A(n2132), .B(n2131), .Z(n2210) );
  XOR U2371 ( .A(n2211), .B(n2210), .Z(n2213) );
  XOR U2372 ( .A(n2212), .B(n2213), .Z(n2223) );
  NANDN U2373 ( .A(n2134), .B(n2133), .Z(n2138) );
  OR U2374 ( .A(n2136), .B(n2135), .Z(n2137) );
  AND U2375 ( .A(n2138), .B(n2137), .Z(n2222) );
  XNOR U2376 ( .A(n2223), .B(n2222), .Z(n2224) );
  NANDN U2377 ( .A(n2140), .B(n2139), .Z(n2144) );
  NANDN U2378 ( .A(n2142), .B(n2141), .Z(n2143) );
  NAND U2379 ( .A(n2144), .B(n2143), .Z(n2225) );
  XNOR U2380 ( .A(n2224), .B(n2225), .Z(n2170) );
  XOR U2381 ( .A(n2171), .B(n2170), .Z(n2229) );
  NANDN U2382 ( .A(n2146), .B(n2145), .Z(n2150) );
  NANDN U2383 ( .A(n2148), .B(n2147), .Z(n2149) );
  AND U2384 ( .A(n2150), .B(n2149), .Z(n2228) );
  XNOR U2385 ( .A(n2229), .B(n2228), .Z(n2230) );
  XOR U2386 ( .A(n2231), .B(n2230), .Z(n2163) );
  NANDN U2387 ( .A(n2152), .B(n2151), .Z(n2156) );
  NAND U2388 ( .A(n2154), .B(n2153), .Z(n2155) );
  AND U2389 ( .A(n2156), .B(n2155), .Z(n2162) );
  XNOR U2390 ( .A(n2163), .B(n2162), .Z(n2164) );
  XNOR U2391 ( .A(n2165), .B(n2164), .Z(n2234) );
  XNOR U2392 ( .A(sreg[275]), .B(n2234), .Z(n2236) );
  NANDN U2393 ( .A(sreg[274]), .B(n2157), .Z(n2161) );
  NAND U2394 ( .A(n2159), .B(n2158), .Z(n2160) );
  NAND U2395 ( .A(n2161), .B(n2160), .Z(n2235) );
  XNOR U2396 ( .A(n2236), .B(n2235), .Z(c[275]) );
  NANDN U2397 ( .A(n2163), .B(n2162), .Z(n2167) );
  NANDN U2398 ( .A(n2165), .B(n2164), .Z(n2166) );
  AND U2399 ( .A(n2167), .B(n2166), .Z(n2242) );
  NANDN U2400 ( .A(n2169), .B(n2168), .Z(n2173) );
  NAND U2401 ( .A(n2171), .B(n2170), .Z(n2172) );
  AND U2402 ( .A(n2173), .B(n2172), .Z(n2308) );
  NANDN U2403 ( .A(n2175), .B(n2174), .Z(n2179) );
  NANDN U2404 ( .A(n2177), .B(n2176), .Z(n2178) );
  AND U2405 ( .A(n2179), .B(n2178), .Z(n2274) );
  NAND U2406 ( .A(b[0]), .B(a[36]), .Z(n2180) );
  XNOR U2407 ( .A(b[1]), .B(n2180), .Z(n2182) );
  NANDN U2408 ( .A(b[0]), .B(a[35]), .Z(n2181) );
  NAND U2409 ( .A(n2182), .B(n2181), .Z(n2254) );
  NAND U2410 ( .A(n19808), .B(n2183), .Z(n2185) );
  XOR U2411 ( .A(b[13]), .B(a[24]), .Z(n2260) );
  NAND U2412 ( .A(n19768), .B(n2260), .Z(n2184) );
  AND U2413 ( .A(n2185), .B(n2184), .Z(n2252) );
  AND U2414 ( .A(b[15]), .B(a[20]), .Z(n2251) );
  XNOR U2415 ( .A(n2252), .B(n2251), .Z(n2253) );
  XNOR U2416 ( .A(n2254), .B(n2253), .Z(n2272) );
  NAND U2417 ( .A(n33), .B(n2186), .Z(n2188) );
  XOR U2418 ( .A(b[5]), .B(a[32]), .Z(n2263) );
  NAND U2419 ( .A(n19342), .B(n2263), .Z(n2187) );
  AND U2420 ( .A(n2188), .B(n2187), .Z(n2296) );
  NAND U2421 ( .A(n34), .B(n2189), .Z(n2191) );
  XOR U2422 ( .A(b[7]), .B(a[30]), .Z(n2266) );
  NAND U2423 ( .A(n19486), .B(n2266), .Z(n2190) );
  AND U2424 ( .A(n2191), .B(n2190), .Z(n2294) );
  NAND U2425 ( .A(n31), .B(n2192), .Z(n2194) );
  XOR U2426 ( .A(b[3]), .B(a[34]), .Z(n2269) );
  NAND U2427 ( .A(n32), .B(n2269), .Z(n2193) );
  NAND U2428 ( .A(n2194), .B(n2193), .Z(n2293) );
  XNOR U2429 ( .A(n2294), .B(n2293), .Z(n2295) );
  XOR U2430 ( .A(n2296), .B(n2295), .Z(n2273) );
  XOR U2431 ( .A(n2272), .B(n2273), .Z(n2275) );
  XOR U2432 ( .A(n2274), .B(n2275), .Z(n2246) );
  NANDN U2433 ( .A(n2196), .B(n2195), .Z(n2200) );
  OR U2434 ( .A(n2198), .B(n2197), .Z(n2199) );
  AND U2435 ( .A(n2200), .B(n2199), .Z(n2245) );
  XNOR U2436 ( .A(n2246), .B(n2245), .Z(n2248) );
  NAND U2437 ( .A(n2201), .B(n19724), .Z(n2203) );
  XOR U2438 ( .A(b[11]), .B(a[26]), .Z(n2278) );
  NAND U2439 ( .A(n19692), .B(n2278), .Z(n2202) );
  AND U2440 ( .A(n2203), .B(n2202), .Z(n2289) );
  NAND U2441 ( .A(n19838), .B(n2204), .Z(n2206) );
  XOR U2442 ( .A(b[15]), .B(a[22]), .Z(n2281) );
  NAND U2443 ( .A(n19805), .B(n2281), .Z(n2205) );
  AND U2444 ( .A(n2206), .B(n2205), .Z(n2288) );
  NAND U2445 ( .A(n35), .B(n2207), .Z(n2209) );
  XOR U2446 ( .A(b[9]), .B(a[28]), .Z(n2284) );
  NAND U2447 ( .A(n19598), .B(n2284), .Z(n2208) );
  NAND U2448 ( .A(n2209), .B(n2208), .Z(n2287) );
  XOR U2449 ( .A(n2288), .B(n2287), .Z(n2290) );
  XOR U2450 ( .A(n2289), .B(n2290), .Z(n2300) );
  NANDN U2451 ( .A(n2211), .B(n2210), .Z(n2215) );
  OR U2452 ( .A(n2213), .B(n2212), .Z(n2214) );
  AND U2453 ( .A(n2215), .B(n2214), .Z(n2299) );
  XNOR U2454 ( .A(n2300), .B(n2299), .Z(n2301) );
  NANDN U2455 ( .A(n2217), .B(n2216), .Z(n2221) );
  NANDN U2456 ( .A(n2219), .B(n2218), .Z(n2220) );
  NAND U2457 ( .A(n2221), .B(n2220), .Z(n2302) );
  XNOR U2458 ( .A(n2301), .B(n2302), .Z(n2247) );
  XOR U2459 ( .A(n2248), .B(n2247), .Z(n2306) );
  NANDN U2460 ( .A(n2223), .B(n2222), .Z(n2227) );
  NANDN U2461 ( .A(n2225), .B(n2224), .Z(n2226) );
  AND U2462 ( .A(n2227), .B(n2226), .Z(n2305) );
  XNOR U2463 ( .A(n2306), .B(n2305), .Z(n2307) );
  XOR U2464 ( .A(n2308), .B(n2307), .Z(n2240) );
  NANDN U2465 ( .A(n2229), .B(n2228), .Z(n2233) );
  NAND U2466 ( .A(n2231), .B(n2230), .Z(n2232) );
  AND U2467 ( .A(n2233), .B(n2232), .Z(n2239) );
  XNOR U2468 ( .A(n2240), .B(n2239), .Z(n2241) );
  XNOR U2469 ( .A(n2242), .B(n2241), .Z(n2311) );
  XNOR U2470 ( .A(sreg[276]), .B(n2311), .Z(n2313) );
  NANDN U2471 ( .A(sreg[275]), .B(n2234), .Z(n2238) );
  NAND U2472 ( .A(n2236), .B(n2235), .Z(n2237) );
  NAND U2473 ( .A(n2238), .B(n2237), .Z(n2312) );
  XNOR U2474 ( .A(n2313), .B(n2312), .Z(c[276]) );
  NANDN U2475 ( .A(n2240), .B(n2239), .Z(n2244) );
  NANDN U2476 ( .A(n2242), .B(n2241), .Z(n2243) );
  AND U2477 ( .A(n2244), .B(n2243), .Z(n2324) );
  NANDN U2478 ( .A(n2246), .B(n2245), .Z(n2250) );
  NAND U2479 ( .A(n2248), .B(n2247), .Z(n2249) );
  AND U2480 ( .A(n2250), .B(n2249), .Z(n2390) );
  NANDN U2481 ( .A(n2252), .B(n2251), .Z(n2256) );
  NANDN U2482 ( .A(n2254), .B(n2253), .Z(n2255) );
  AND U2483 ( .A(n2256), .B(n2255), .Z(n2356) );
  NAND U2484 ( .A(b[0]), .B(a[37]), .Z(n2257) );
  XNOR U2485 ( .A(b[1]), .B(n2257), .Z(n2259) );
  NANDN U2486 ( .A(b[0]), .B(a[36]), .Z(n2258) );
  NAND U2487 ( .A(n2259), .B(n2258), .Z(n2336) );
  NAND U2488 ( .A(n19808), .B(n2260), .Z(n2262) );
  XOR U2489 ( .A(b[13]), .B(a[25]), .Z(n2339) );
  NAND U2490 ( .A(n19768), .B(n2339), .Z(n2261) );
  AND U2491 ( .A(n2262), .B(n2261), .Z(n2334) );
  AND U2492 ( .A(b[15]), .B(a[21]), .Z(n2333) );
  XNOR U2493 ( .A(n2334), .B(n2333), .Z(n2335) );
  XNOR U2494 ( .A(n2336), .B(n2335), .Z(n2354) );
  NAND U2495 ( .A(n33), .B(n2263), .Z(n2265) );
  XOR U2496 ( .A(b[5]), .B(a[33]), .Z(n2345) );
  NAND U2497 ( .A(n19342), .B(n2345), .Z(n2264) );
  AND U2498 ( .A(n2265), .B(n2264), .Z(n2378) );
  NAND U2499 ( .A(n34), .B(n2266), .Z(n2268) );
  XOR U2500 ( .A(b[7]), .B(a[31]), .Z(n2348) );
  NAND U2501 ( .A(n19486), .B(n2348), .Z(n2267) );
  AND U2502 ( .A(n2268), .B(n2267), .Z(n2376) );
  NAND U2503 ( .A(n31), .B(n2269), .Z(n2271) );
  XOR U2504 ( .A(b[3]), .B(a[35]), .Z(n2351) );
  NAND U2505 ( .A(n32), .B(n2351), .Z(n2270) );
  NAND U2506 ( .A(n2271), .B(n2270), .Z(n2375) );
  XNOR U2507 ( .A(n2376), .B(n2375), .Z(n2377) );
  XOR U2508 ( .A(n2378), .B(n2377), .Z(n2355) );
  XOR U2509 ( .A(n2354), .B(n2355), .Z(n2357) );
  XOR U2510 ( .A(n2356), .B(n2357), .Z(n2328) );
  NANDN U2511 ( .A(n2273), .B(n2272), .Z(n2277) );
  OR U2512 ( .A(n2275), .B(n2274), .Z(n2276) );
  AND U2513 ( .A(n2277), .B(n2276), .Z(n2327) );
  XNOR U2514 ( .A(n2328), .B(n2327), .Z(n2330) );
  NAND U2515 ( .A(n2278), .B(n19724), .Z(n2280) );
  XOR U2516 ( .A(b[11]), .B(a[27]), .Z(n2360) );
  NAND U2517 ( .A(n19692), .B(n2360), .Z(n2279) );
  AND U2518 ( .A(n2280), .B(n2279), .Z(n2371) );
  NAND U2519 ( .A(n19838), .B(n2281), .Z(n2283) );
  XOR U2520 ( .A(b[15]), .B(a[23]), .Z(n2363) );
  NAND U2521 ( .A(n19805), .B(n2363), .Z(n2282) );
  AND U2522 ( .A(n2283), .B(n2282), .Z(n2370) );
  NAND U2523 ( .A(n35), .B(n2284), .Z(n2286) );
  XOR U2524 ( .A(b[9]), .B(a[29]), .Z(n2366) );
  NAND U2525 ( .A(n19598), .B(n2366), .Z(n2285) );
  NAND U2526 ( .A(n2286), .B(n2285), .Z(n2369) );
  XOR U2527 ( .A(n2370), .B(n2369), .Z(n2372) );
  XOR U2528 ( .A(n2371), .B(n2372), .Z(n2382) );
  NANDN U2529 ( .A(n2288), .B(n2287), .Z(n2292) );
  OR U2530 ( .A(n2290), .B(n2289), .Z(n2291) );
  AND U2531 ( .A(n2292), .B(n2291), .Z(n2381) );
  XNOR U2532 ( .A(n2382), .B(n2381), .Z(n2383) );
  NANDN U2533 ( .A(n2294), .B(n2293), .Z(n2298) );
  NANDN U2534 ( .A(n2296), .B(n2295), .Z(n2297) );
  NAND U2535 ( .A(n2298), .B(n2297), .Z(n2384) );
  XNOR U2536 ( .A(n2383), .B(n2384), .Z(n2329) );
  XOR U2537 ( .A(n2330), .B(n2329), .Z(n2388) );
  NANDN U2538 ( .A(n2300), .B(n2299), .Z(n2304) );
  NANDN U2539 ( .A(n2302), .B(n2301), .Z(n2303) );
  AND U2540 ( .A(n2304), .B(n2303), .Z(n2387) );
  XNOR U2541 ( .A(n2388), .B(n2387), .Z(n2389) );
  XOR U2542 ( .A(n2390), .B(n2389), .Z(n2322) );
  NANDN U2543 ( .A(n2306), .B(n2305), .Z(n2310) );
  NAND U2544 ( .A(n2308), .B(n2307), .Z(n2309) );
  AND U2545 ( .A(n2310), .B(n2309), .Z(n2321) );
  XNOR U2546 ( .A(n2322), .B(n2321), .Z(n2323) );
  XNOR U2547 ( .A(n2324), .B(n2323), .Z(n2316) );
  XNOR U2548 ( .A(sreg[277]), .B(n2316), .Z(n2318) );
  NANDN U2549 ( .A(sreg[276]), .B(n2311), .Z(n2315) );
  NAND U2550 ( .A(n2313), .B(n2312), .Z(n2314) );
  NAND U2551 ( .A(n2315), .B(n2314), .Z(n2317) );
  XNOR U2552 ( .A(n2318), .B(n2317), .Z(c[277]) );
  NANDN U2553 ( .A(sreg[277]), .B(n2316), .Z(n2320) );
  NAND U2554 ( .A(n2318), .B(n2317), .Z(n2319) );
  AND U2555 ( .A(n2320), .B(n2319), .Z(n2395) );
  NANDN U2556 ( .A(n2322), .B(n2321), .Z(n2326) );
  NANDN U2557 ( .A(n2324), .B(n2323), .Z(n2325) );
  AND U2558 ( .A(n2326), .B(n2325), .Z(n2400) );
  NANDN U2559 ( .A(n2328), .B(n2327), .Z(n2332) );
  NAND U2560 ( .A(n2330), .B(n2329), .Z(n2331) );
  AND U2561 ( .A(n2332), .B(n2331), .Z(n2467) );
  NANDN U2562 ( .A(n2334), .B(n2333), .Z(n2338) );
  NANDN U2563 ( .A(n2336), .B(n2335), .Z(n2337) );
  AND U2564 ( .A(n2338), .B(n2337), .Z(n2433) );
  NAND U2565 ( .A(n19808), .B(n2339), .Z(n2341) );
  XOR U2566 ( .A(b[13]), .B(a[26]), .Z(n2419) );
  NAND U2567 ( .A(n19768), .B(n2419), .Z(n2340) );
  AND U2568 ( .A(n2341), .B(n2340), .Z(n2411) );
  AND U2569 ( .A(b[15]), .B(a[22]), .Z(n2410) );
  XNOR U2570 ( .A(n2411), .B(n2410), .Z(n2412) );
  NAND U2571 ( .A(b[0]), .B(a[38]), .Z(n2342) );
  XNOR U2572 ( .A(b[1]), .B(n2342), .Z(n2344) );
  NANDN U2573 ( .A(b[0]), .B(a[37]), .Z(n2343) );
  NAND U2574 ( .A(n2344), .B(n2343), .Z(n2413) );
  XNOR U2575 ( .A(n2412), .B(n2413), .Z(n2431) );
  NAND U2576 ( .A(n33), .B(n2345), .Z(n2347) );
  XOR U2577 ( .A(b[5]), .B(a[34]), .Z(n2422) );
  NAND U2578 ( .A(n19342), .B(n2422), .Z(n2346) );
  AND U2579 ( .A(n2347), .B(n2346), .Z(n2455) );
  NAND U2580 ( .A(n34), .B(n2348), .Z(n2350) );
  XOR U2581 ( .A(b[7]), .B(a[32]), .Z(n2425) );
  NAND U2582 ( .A(n19486), .B(n2425), .Z(n2349) );
  AND U2583 ( .A(n2350), .B(n2349), .Z(n2453) );
  NAND U2584 ( .A(n31), .B(n2351), .Z(n2353) );
  XOR U2585 ( .A(b[3]), .B(a[36]), .Z(n2428) );
  NAND U2586 ( .A(n32), .B(n2428), .Z(n2352) );
  NAND U2587 ( .A(n2353), .B(n2352), .Z(n2452) );
  XNOR U2588 ( .A(n2453), .B(n2452), .Z(n2454) );
  XOR U2589 ( .A(n2455), .B(n2454), .Z(n2432) );
  XOR U2590 ( .A(n2431), .B(n2432), .Z(n2434) );
  XOR U2591 ( .A(n2433), .B(n2434), .Z(n2405) );
  NANDN U2592 ( .A(n2355), .B(n2354), .Z(n2359) );
  OR U2593 ( .A(n2357), .B(n2356), .Z(n2358) );
  AND U2594 ( .A(n2359), .B(n2358), .Z(n2404) );
  XNOR U2595 ( .A(n2405), .B(n2404), .Z(n2407) );
  NAND U2596 ( .A(n2360), .B(n19724), .Z(n2362) );
  XOR U2597 ( .A(b[11]), .B(a[28]), .Z(n2437) );
  NAND U2598 ( .A(n19692), .B(n2437), .Z(n2361) );
  AND U2599 ( .A(n2362), .B(n2361), .Z(n2448) );
  NAND U2600 ( .A(n19838), .B(n2363), .Z(n2365) );
  XOR U2601 ( .A(b[15]), .B(a[24]), .Z(n2440) );
  NAND U2602 ( .A(n19805), .B(n2440), .Z(n2364) );
  AND U2603 ( .A(n2365), .B(n2364), .Z(n2447) );
  NAND U2604 ( .A(n35), .B(n2366), .Z(n2368) );
  XOR U2605 ( .A(b[9]), .B(a[30]), .Z(n2443) );
  NAND U2606 ( .A(n19598), .B(n2443), .Z(n2367) );
  NAND U2607 ( .A(n2368), .B(n2367), .Z(n2446) );
  XOR U2608 ( .A(n2447), .B(n2446), .Z(n2449) );
  XOR U2609 ( .A(n2448), .B(n2449), .Z(n2459) );
  NANDN U2610 ( .A(n2370), .B(n2369), .Z(n2374) );
  OR U2611 ( .A(n2372), .B(n2371), .Z(n2373) );
  AND U2612 ( .A(n2374), .B(n2373), .Z(n2458) );
  XNOR U2613 ( .A(n2459), .B(n2458), .Z(n2460) );
  NANDN U2614 ( .A(n2376), .B(n2375), .Z(n2380) );
  NANDN U2615 ( .A(n2378), .B(n2377), .Z(n2379) );
  NAND U2616 ( .A(n2380), .B(n2379), .Z(n2461) );
  XNOR U2617 ( .A(n2460), .B(n2461), .Z(n2406) );
  XOR U2618 ( .A(n2407), .B(n2406), .Z(n2465) );
  NANDN U2619 ( .A(n2382), .B(n2381), .Z(n2386) );
  NANDN U2620 ( .A(n2384), .B(n2383), .Z(n2385) );
  AND U2621 ( .A(n2386), .B(n2385), .Z(n2464) );
  XNOR U2622 ( .A(n2465), .B(n2464), .Z(n2466) );
  XOR U2623 ( .A(n2467), .B(n2466), .Z(n2399) );
  NANDN U2624 ( .A(n2388), .B(n2387), .Z(n2392) );
  NAND U2625 ( .A(n2390), .B(n2389), .Z(n2391) );
  AND U2626 ( .A(n2392), .B(n2391), .Z(n2398) );
  XOR U2627 ( .A(n2399), .B(n2398), .Z(n2401) );
  XOR U2628 ( .A(n2400), .B(n2401), .Z(n2393) );
  XNOR U2629 ( .A(n2393), .B(sreg[278]), .Z(n2394) );
  XOR U2630 ( .A(n2395), .B(n2394), .Z(c[278]) );
  NANDN U2631 ( .A(n2393), .B(sreg[278]), .Z(n2397) );
  NAND U2632 ( .A(n2395), .B(n2394), .Z(n2396) );
  AND U2633 ( .A(n2397), .B(n2396), .Z(n2544) );
  NANDN U2634 ( .A(n2399), .B(n2398), .Z(n2403) );
  OR U2635 ( .A(n2401), .B(n2400), .Z(n2402) );
  AND U2636 ( .A(n2403), .B(n2402), .Z(n2473) );
  NANDN U2637 ( .A(n2405), .B(n2404), .Z(n2409) );
  NAND U2638 ( .A(n2407), .B(n2406), .Z(n2408) );
  AND U2639 ( .A(n2409), .B(n2408), .Z(n2539) );
  NANDN U2640 ( .A(n2411), .B(n2410), .Z(n2415) );
  NANDN U2641 ( .A(n2413), .B(n2412), .Z(n2414) );
  AND U2642 ( .A(n2415), .B(n2414), .Z(n2505) );
  NAND U2643 ( .A(b[0]), .B(a[39]), .Z(n2416) );
  XNOR U2644 ( .A(b[1]), .B(n2416), .Z(n2418) );
  NANDN U2645 ( .A(b[0]), .B(a[38]), .Z(n2417) );
  NAND U2646 ( .A(n2418), .B(n2417), .Z(n2485) );
  NAND U2647 ( .A(n19808), .B(n2419), .Z(n2421) );
  XOR U2648 ( .A(b[13]), .B(a[27]), .Z(n2491) );
  NAND U2649 ( .A(n19768), .B(n2491), .Z(n2420) );
  AND U2650 ( .A(n2421), .B(n2420), .Z(n2483) );
  AND U2651 ( .A(b[15]), .B(a[23]), .Z(n2482) );
  XNOR U2652 ( .A(n2483), .B(n2482), .Z(n2484) );
  XNOR U2653 ( .A(n2485), .B(n2484), .Z(n2503) );
  NAND U2654 ( .A(n33), .B(n2422), .Z(n2424) );
  XOR U2655 ( .A(b[5]), .B(a[35]), .Z(n2494) );
  NAND U2656 ( .A(n19342), .B(n2494), .Z(n2423) );
  AND U2657 ( .A(n2424), .B(n2423), .Z(n2527) );
  NAND U2658 ( .A(n34), .B(n2425), .Z(n2427) );
  XOR U2659 ( .A(b[7]), .B(a[33]), .Z(n2497) );
  NAND U2660 ( .A(n19486), .B(n2497), .Z(n2426) );
  AND U2661 ( .A(n2427), .B(n2426), .Z(n2525) );
  NAND U2662 ( .A(n31), .B(n2428), .Z(n2430) );
  XOR U2663 ( .A(b[3]), .B(a[37]), .Z(n2500) );
  NAND U2664 ( .A(n32), .B(n2500), .Z(n2429) );
  NAND U2665 ( .A(n2430), .B(n2429), .Z(n2524) );
  XNOR U2666 ( .A(n2525), .B(n2524), .Z(n2526) );
  XOR U2667 ( .A(n2527), .B(n2526), .Z(n2504) );
  XOR U2668 ( .A(n2503), .B(n2504), .Z(n2506) );
  XOR U2669 ( .A(n2505), .B(n2506), .Z(n2477) );
  NANDN U2670 ( .A(n2432), .B(n2431), .Z(n2436) );
  OR U2671 ( .A(n2434), .B(n2433), .Z(n2435) );
  AND U2672 ( .A(n2436), .B(n2435), .Z(n2476) );
  XNOR U2673 ( .A(n2477), .B(n2476), .Z(n2479) );
  NAND U2674 ( .A(n2437), .B(n19724), .Z(n2439) );
  XOR U2675 ( .A(b[11]), .B(a[29]), .Z(n2509) );
  NAND U2676 ( .A(n19692), .B(n2509), .Z(n2438) );
  AND U2677 ( .A(n2439), .B(n2438), .Z(n2520) );
  NAND U2678 ( .A(n19838), .B(n2440), .Z(n2442) );
  XOR U2679 ( .A(b[15]), .B(a[25]), .Z(n2512) );
  NAND U2680 ( .A(n19805), .B(n2512), .Z(n2441) );
  AND U2681 ( .A(n2442), .B(n2441), .Z(n2519) );
  NAND U2682 ( .A(n35), .B(n2443), .Z(n2445) );
  XOR U2683 ( .A(b[9]), .B(a[31]), .Z(n2515) );
  NAND U2684 ( .A(n19598), .B(n2515), .Z(n2444) );
  NAND U2685 ( .A(n2445), .B(n2444), .Z(n2518) );
  XOR U2686 ( .A(n2519), .B(n2518), .Z(n2521) );
  XOR U2687 ( .A(n2520), .B(n2521), .Z(n2531) );
  NANDN U2688 ( .A(n2447), .B(n2446), .Z(n2451) );
  OR U2689 ( .A(n2449), .B(n2448), .Z(n2450) );
  AND U2690 ( .A(n2451), .B(n2450), .Z(n2530) );
  XNOR U2691 ( .A(n2531), .B(n2530), .Z(n2532) );
  NANDN U2692 ( .A(n2453), .B(n2452), .Z(n2457) );
  NANDN U2693 ( .A(n2455), .B(n2454), .Z(n2456) );
  NAND U2694 ( .A(n2457), .B(n2456), .Z(n2533) );
  XNOR U2695 ( .A(n2532), .B(n2533), .Z(n2478) );
  XOR U2696 ( .A(n2479), .B(n2478), .Z(n2537) );
  NANDN U2697 ( .A(n2459), .B(n2458), .Z(n2463) );
  NANDN U2698 ( .A(n2461), .B(n2460), .Z(n2462) );
  AND U2699 ( .A(n2463), .B(n2462), .Z(n2536) );
  XNOR U2700 ( .A(n2537), .B(n2536), .Z(n2538) );
  XOR U2701 ( .A(n2539), .B(n2538), .Z(n2471) );
  NANDN U2702 ( .A(n2465), .B(n2464), .Z(n2469) );
  NAND U2703 ( .A(n2467), .B(n2466), .Z(n2468) );
  AND U2704 ( .A(n2469), .B(n2468), .Z(n2470) );
  XNOR U2705 ( .A(n2471), .B(n2470), .Z(n2472) );
  XNOR U2706 ( .A(n2473), .B(n2472), .Z(n2542) );
  XNOR U2707 ( .A(sreg[279]), .B(n2542), .Z(n2543) );
  XNOR U2708 ( .A(n2544), .B(n2543), .Z(c[279]) );
  NANDN U2709 ( .A(n2471), .B(n2470), .Z(n2475) );
  NANDN U2710 ( .A(n2473), .B(n2472), .Z(n2474) );
  AND U2711 ( .A(n2475), .B(n2474), .Z(n2550) );
  NANDN U2712 ( .A(n2477), .B(n2476), .Z(n2481) );
  NAND U2713 ( .A(n2479), .B(n2478), .Z(n2480) );
  AND U2714 ( .A(n2481), .B(n2480), .Z(n2616) );
  NANDN U2715 ( .A(n2483), .B(n2482), .Z(n2487) );
  NANDN U2716 ( .A(n2485), .B(n2484), .Z(n2486) );
  AND U2717 ( .A(n2487), .B(n2486), .Z(n2582) );
  NAND U2718 ( .A(b[0]), .B(a[40]), .Z(n2488) );
  XNOR U2719 ( .A(b[1]), .B(n2488), .Z(n2490) );
  NANDN U2720 ( .A(b[0]), .B(a[39]), .Z(n2489) );
  NAND U2721 ( .A(n2490), .B(n2489), .Z(n2562) );
  NAND U2722 ( .A(n19808), .B(n2491), .Z(n2493) );
  XOR U2723 ( .A(b[13]), .B(a[28]), .Z(n2568) );
  NAND U2724 ( .A(n19768), .B(n2568), .Z(n2492) );
  AND U2725 ( .A(n2493), .B(n2492), .Z(n2560) );
  AND U2726 ( .A(b[15]), .B(a[24]), .Z(n2559) );
  XNOR U2727 ( .A(n2560), .B(n2559), .Z(n2561) );
  XNOR U2728 ( .A(n2562), .B(n2561), .Z(n2580) );
  NAND U2729 ( .A(n33), .B(n2494), .Z(n2496) );
  XOR U2730 ( .A(b[5]), .B(a[36]), .Z(n2571) );
  NAND U2731 ( .A(n19342), .B(n2571), .Z(n2495) );
  AND U2732 ( .A(n2496), .B(n2495), .Z(n2604) );
  NAND U2733 ( .A(n34), .B(n2497), .Z(n2499) );
  XOR U2734 ( .A(b[7]), .B(a[34]), .Z(n2574) );
  NAND U2735 ( .A(n19486), .B(n2574), .Z(n2498) );
  AND U2736 ( .A(n2499), .B(n2498), .Z(n2602) );
  NAND U2737 ( .A(n31), .B(n2500), .Z(n2502) );
  XOR U2738 ( .A(b[3]), .B(a[38]), .Z(n2577) );
  NAND U2739 ( .A(n32), .B(n2577), .Z(n2501) );
  NAND U2740 ( .A(n2502), .B(n2501), .Z(n2601) );
  XNOR U2741 ( .A(n2602), .B(n2601), .Z(n2603) );
  XOR U2742 ( .A(n2604), .B(n2603), .Z(n2581) );
  XOR U2743 ( .A(n2580), .B(n2581), .Z(n2583) );
  XOR U2744 ( .A(n2582), .B(n2583), .Z(n2554) );
  NANDN U2745 ( .A(n2504), .B(n2503), .Z(n2508) );
  OR U2746 ( .A(n2506), .B(n2505), .Z(n2507) );
  AND U2747 ( .A(n2508), .B(n2507), .Z(n2553) );
  XNOR U2748 ( .A(n2554), .B(n2553), .Z(n2556) );
  NAND U2749 ( .A(n2509), .B(n19724), .Z(n2511) );
  XOR U2750 ( .A(b[11]), .B(a[30]), .Z(n2586) );
  NAND U2751 ( .A(n19692), .B(n2586), .Z(n2510) );
  AND U2752 ( .A(n2511), .B(n2510), .Z(n2597) );
  NAND U2753 ( .A(n19838), .B(n2512), .Z(n2514) );
  XOR U2754 ( .A(b[15]), .B(a[26]), .Z(n2589) );
  NAND U2755 ( .A(n19805), .B(n2589), .Z(n2513) );
  AND U2756 ( .A(n2514), .B(n2513), .Z(n2596) );
  NAND U2757 ( .A(n35), .B(n2515), .Z(n2517) );
  XOR U2758 ( .A(b[9]), .B(a[32]), .Z(n2592) );
  NAND U2759 ( .A(n19598), .B(n2592), .Z(n2516) );
  NAND U2760 ( .A(n2517), .B(n2516), .Z(n2595) );
  XOR U2761 ( .A(n2596), .B(n2595), .Z(n2598) );
  XOR U2762 ( .A(n2597), .B(n2598), .Z(n2608) );
  NANDN U2763 ( .A(n2519), .B(n2518), .Z(n2523) );
  OR U2764 ( .A(n2521), .B(n2520), .Z(n2522) );
  AND U2765 ( .A(n2523), .B(n2522), .Z(n2607) );
  XNOR U2766 ( .A(n2608), .B(n2607), .Z(n2609) );
  NANDN U2767 ( .A(n2525), .B(n2524), .Z(n2529) );
  NANDN U2768 ( .A(n2527), .B(n2526), .Z(n2528) );
  NAND U2769 ( .A(n2529), .B(n2528), .Z(n2610) );
  XNOR U2770 ( .A(n2609), .B(n2610), .Z(n2555) );
  XOR U2771 ( .A(n2556), .B(n2555), .Z(n2614) );
  NANDN U2772 ( .A(n2531), .B(n2530), .Z(n2535) );
  NANDN U2773 ( .A(n2533), .B(n2532), .Z(n2534) );
  AND U2774 ( .A(n2535), .B(n2534), .Z(n2613) );
  XNOR U2775 ( .A(n2614), .B(n2613), .Z(n2615) );
  XOR U2776 ( .A(n2616), .B(n2615), .Z(n2548) );
  NANDN U2777 ( .A(n2537), .B(n2536), .Z(n2541) );
  NAND U2778 ( .A(n2539), .B(n2538), .Z(n2540) );
  AND U2779 ( .A(n2541), .B(n2540), .Z(n2547) );
  XNOR U2780 ( .A(n2548), .B(n2547), .Z(n2549) );
  XNOR U2781 ( .A(n2550), .B(n2549), .Z(n2619) );
  XNOR U2782 ( .A(sreg[280]), .B(n2619), .Z(n2621) );
  NANDN U2783 ( .A(sreg[279]), .B(n2542), .Z(n2546) );
  NAND U2784 ( .A(n2544), .B(n2543), .Z(n2545) );
  NAND U2785 ( .A(n2546), .B(n2545), .Z(n2620) );
  XNOR U2786 ( .A(n2621), .B(n2620), .Z(c[280]) );
  NANDN U2787 ( .A(n2548), .B(n2547), .Z(n2552) );
  NANDN U2788 ( .A(n2550), .B(n2549), .Z(n2551) );
  AND U2789 ( .A(n2552), .B(n2551), .Z(n2627) );
  NANDN U2790 ( .A(n2554), .B(n2553), .Z(n2558) );
  NAND U2791 ( .A(n2556), .B(n2555), .Z(n2557) );
  AND U2792 ( .A(n2558), .B(n2557), .Z(n2693) );
  NANDN U2793 ( .A(n2560), .B(n2559), .Z(n2564) );
  NANDN U2794 ( .A(n2562), .B(n2561), .Z(n2563) );
  AND U2795 ( .A(n2564), .B(n2563), .Z(n2659) );
  NAND U2796 ( .A(b[0]), .B(a[41]), .Z(n2565) );
  XNOR U2797 ( .A(b[1]), .B(n2565), .Z(n2567) );
  NANDN U2798 ( .A(b[0]), .B(a[40]), .Z(n2566) );
  NAND U2799 ( .A(n2567), .B(n2566), .Z(n2639) );
  NAND U2800 ( .A(n19808), .B(n2568), .Z(n2570) );
  XOR U2801 ( .A(b[13]), .B(a[29]), .Z(n2645) );
  NAND U2802 ( .A(n19768), .B(n2645), .Z(n2569) );
  AND U2803 ( .A(n2570), .B(n2569), .Z(n2637) );
  AND U2804 ( .A(b[15]), .B(a[25]), .Z(n2636) );
  XNOR U2805 ( .A(n2637), .B(n2636), .Z(n2638) );
  XNOR U2806 ( .A(n2639), .B(n2638), .Z(n2657) );
  NAND U2807 ( .A(n33), .B(n2571), .Z(n2573) );
  XOR U2808 ( .A(b[5]), .B(a[37]), .Z(n2648) );
  NAND U2809 ( .A(n19342), .B(n2648), .Z(n2572) );
  AND U2810 ( .A(n2573), .B(n2572), .Z(n2681) );
  NAND U2811 ( .A(n34), .B(n2574), .Z(n2576) );
  XOR U2812 ( .A(b[7]), .B(a[35]), .Z(n2651) );
  NAND U2813 ( .A(n19486), .B(n2651), .Z(n2575) );
  AND U2814 ( .A(n2576), .B(n2575), .Z(n2679) );
  NAND U2815 ( .A(n31), .B(n2577), .Z(n2579) );
  XOR U2816 ( .A(b[3]), .B(a[39]), .Z(n2654) );
  NAND U2817 ( .A(n32), .B(n2654), .Z(n2578) );
  NAND U2818 ( .A(n2579), .B(n2578), .Z(n2678) );
  XNOR U2819 ( .A(n2679), .B(n2678), .Z(n2680) );
  XOR U2820 ( .A(n2681), .B(n2680), .Z(n2658) );
  XOR U2821 ( .A(n2657), .B(n2658), .Z(n2660) );
  XOR U2822 ( .A(n2659), .B(n2660), .Z(n2631) );
  NANDN U2823 ( .A(n2581), .B(n2580), .Z(n2585) );
  OR U2824 ( .A(n2583), .B(n2582), .Z(n2584) );
  AND U2825 ( .A(n2585), .B(n2584), .Z(n2630) );
  XNOR U2826 ( .A(n2631), .B(n2630), .Z(n2633) );
  NAND U2827 ( .A(n2586), .B(n19724), .Z(n2588) );
  XOR U2828 ( .A(b[11]), .B(a[31]), .Z(n2663) );
  NAND U2829 ( .A(n19692), .B(n2663), .Z(n2587) );
  AND U2830 ( .A(n2588), .B(n2587), .Z(n2674) );
  NAND U2831 ( .A(n19838), .B(n2589), .Z(n2591) );
  XOR U2832 ( .A(b[15]), .B(a[27]), .Z(n2666) );
  NAND U2833 ( .A(n19805), .B(n2666), .Z(n2590) );
  AND U2834 ( .A(n2591), .B(n2590), .Z(n2673) );
  NAND U2835 ( .A(n35), .B(n2592), .Z(n2594) );
  XOR U2836 ( .A(b[9]), .B(a[33]), .Z(n2669) );
  NAND U2837 ( .A(n19598), .B(n2669), .Z(n2593) );
  NAND U2838 ( .A(n2594), .B(n2593), .Z(n2672) );
  XOR U2839 ( .A(n2673), .B(n2672), .Z(n2675) );
  XOR U2840 ( .A(n2674), .B(n2675), .Z(n2685) );
  NANDN U2841 ( .A(n2596), .B(n2595), .Z(n2600) );
  OR U2842 ( .A(n2598), .B(n2597), .Z(n2599) );
  AND U2843 ( .A(n2600), .B(n2599), .Z(n2684) );
  XNOR U2844 ( .A(n2685), .B(n2684), .Z(n2686) );
  NANDN U2845 ( .A(n2602), .B(n2601), .Z(n2606) );
  NANDN U2846 ( .A(n2604), .B(n2603), .Z(n2605) );
  NAND U2847 ( .A(n2606), .B(n2605), .Z(n2687) );
  XNOR U2848 ( .A(n2686), .B(n2687), .Z(n2632) );
  XOR U2849 ( .A(n2633), .B(n2632), .Z(n2691) );
  NANDN U2850 ( .A(n2608), .B(n2607), .Z(n2612) );
  NANDN U2851 ( .A(n2610), .B(n2609), .Z(n2611) );
  AND U2852 ( .A(n2612), .B(n2611), .Z(n2690) );
  XNOR U2853 ( .A(n2691), .B(n2690), .Z(n2692) );
  XOR U2854 ( .A(n2693), .B(n2692), .Z(n2625) );
  NANDN U2855 ( .A(n2614), .B(n2613), .Z(n2618) );
  NAND U2856 ( .A(n2616), .B(n2615), .Z(n2617) );
  AND U2857 ( .A(n2618), .B(n2617), .Z(n2624) );
  XNOR U2858 ( .A(n2625), .B(n2624), .Z(n2626) );
  XNOR U2859 ( .A(n2627), .B(n2626), .Z(n2696) );
  XNOR U2860 ( .A(sreg[281]), .B(n2696), .Z(n2698) );
  NANDN U2861 ( .A(sreg[280]), .B(n2619), .Z(n2623) );
  NAND U2862 ( .A(n2621), .B(n2620), .Z(n2622) );
  NAND U2863 ( .A(n2623), .B(n2622), .Z(n2697) );
  XNOR U2864 ( .A(n2698), .B(n2697), .Z(c[281]) );
  NANDN U2865 ( .A(n2625), .B(n2624), .Z(n2629) );
  NANDN U2866 ( .A(n2627), .B(n2626), .Z(n2628) );
  AND U2867 ( .A(n2629), .B(n2628), .Z(n2704) );
  NANDN U2868 ( .A(n2631), .B(n2630), .Z(n2635) );
  NAND U2869 ( .A(n2633), .B(n2632), .Z(n2634) );
  AND U2870 ( .A(n2635), .B(n2634), .Z(n2770) );
  NANDN U2871 ( .A(n2637), .B(n2636), .Z(n2641) );
  NANDN U2872 ( .A(n2639), .B(n2638), .Z(n2640) );
  AND U2873 ( .A(n2641), .B(n2640), .Z(n2736) );
  NAND U2874 ( .A(b[0]), .B(a[42]), .Z(n2642) );
  XNOR U2875 ( .A(b[1]), .B(n2642), .Z(n2644) );
  NANDN U2876 ( .A(b[0]), .B(a[41]), .Z(n2643) );
  NAND U2877 ( .A(n2644), .B(n2643), .Z(n2716) );
  NAND U2878 ( .A(n19808), .B(n2645), .Z(n2647) );
  XOR U2879 ( .A(b[13]), .B(a[30]), .Z(n2722) );
  NAND U2880 ( .A(n19768), .B(n2722), .Z(n2646) );
  AND U2881 ( .A(n2647), .B(n2646), .Z(n2714) );
  AND U2882 ( .A(b[15]), .B(a[26]), .Z(n2713) );
  XNOR U2883 ( .A(n2714), .B(n2713), .Z(n2715) );
  XNOR U2884 ( .A(n2716), .B(n2715), .Z(n2734) );
  NAND U2885 ( .A(n33), .B(n2648), .Z(n2650) );
  XOR U2886 ( .A(b[5]), .B(a[38]), .Z(n2725) );
  NAND U2887 ( .A(n19342), .B(n2725), .Z(n2649) );
  AND U2888 ( .A(n2650), .B(n2649), .Z(n2758) );
  NAND U2889 ( .A(n34), .B(n2651), .Z(n2653) );
  XOR U2890 ( .A(b[7]), .B(a[36]), .Z(n2728) );
  NAND U2891 ( .A(n19486), .B(n2728), .Z(n2652) );
  AND U2892 ( .A(n2653), .B(n2652), .Z(n2756) );
  NAND U2893 ( .A(n31), .B(n2654), .Z(n2656) );
  XOR U2894 ( .A(b[3]), .B(a[40]), .Z(n2731) );
  NAND U2895 ( .A(n32), .B(n2731), .Z(n2655) );
  NAND U2896 ( .A(n2656), .B(n2655), .Z(n2755) );
  XNOR U2897 ( .A(n2756), .B(n2755), .Z(n2757) );
  XOR U2898 ( .A(n2758), .B(n2757), .Z(n2735) );
  XOR U2899 ( .A(n2734), .B(n2735), .Z(n2737) );
  XOR U2900 ( .A(n2736), .B(n2737), .Z(n2708) );
  NANDN U2901 ( .A(n2658), .B(n2657), .Z(n2662) );
  OR U2902 ( .A(n2660), .B(n2659), .Z(n2661) );
  AND U2903 ( .A(n2662), .B(n2661), .Z(n2707) );
  XNOR U2904 ( .A(n2708), .B(n2707), .Z(n2710) );
  NAND U2905 ( .A(n2663), .B(n19724), .Z(n2665) );
  XOR U2906 ( .A(b[11]), .B(a[32]), .Z(n2740) );
  NAND U2907 ( .A(n19692), .B(n2740), .Z(n2664) );
  AND U2908 ( .A(n2665), .B(n2664), .Z(n2751) );
  NAND U2909 ( .A(n19838), .B(n2666), .Z(n2668) );
  XOR U2910 ( .A(b[15]), .B(a[28]), .Z(n2743) );
  NAND U2911 ( .A(n19805), .B(n2743), .Z(n2667) );
  AND U2912 ( .A(n2668), .B(n2667), .Z(n2750) );
  NAND U2913 ( .A(n35), .B(n2669), .Z(n2671) );
  XOR U2914 ( .A(b[9]), .B(a[34]), .Z(n2746) );
  NAND U2915 ( .A(n19598), .B(n2746), .Z(n2670) );
  NAND U2916 ( .A(n2671), .B(n2670), .Z(n2749) );
  XOR U2917 ( .A(n2750), .B(n2749), .Z(n2752) );
  XOR U2918 ( .A(n2751), .B(n2752), .Z(n2762) );
  NANDN U2919 ( .A(n2673), .B(n2672), .Z(n2677) );
  OR U2920 ( .A(n2675), .B(n2674), .Z(n2676) );
  AND U2921 ( .A(n2677), .B(n2676), .Z(n2761) );
  XNOR U2922 ( .A(n2762), .B(n2761), .Z(n2763) );
  NANDN U2923 ( .A(n2679), .B(n2678), .Z(n2683) );
  NANDN U2924 ( .A(n2681), .B(n2680), .Z(n2682) );
  NAND U2925 ( .A(n2683), .B(n2682), .Z(n2764) );
  XNOR U2926 ( .A(n2763), .B(n2764), .Z(n2709) );
  XOR U2927 ( .A(n2710), .B(n2709), .Z(n2768) );
  NANDN U2928 ( .A(n2685), .B(n2684), .Z(n2689) );
  NANDN U2929 ( .A(n2687), .B(n2686), .Z(n2688) );
  AND U2930 ( .A(n2689), .B(n2688), .Z(n2767) );
  XNOR U2931 ( .A(n2768), .B(n2767), .Z(n2769) );
  XOR U2932 ( .A(n2770), .B(n2769), .Z(n2702) );
  NANDN U2933 ( .A(n2691), .B(n2690), .Z(n2695) );
  NAND U2934 ( .A(n2693), .B(n2692), .Z(n2694) );
  AND U2935 ( .A(n2695), .B(n2694), .Z(n2701) );
  XNOR U2936 ( .A(n2702), .B(n2701), .Z(n2703) );
  XNOR U2937 ( .A(n2704), .B(n2703), .Z(n2773) );
  XNOR U2938 ( .A(sreg[282]), .B(n2773), .Z(n2775) );
  NANDN U2939 ( .A(sreg[281]), .B(n2696), .Z(n2700) );
  NAND U2940 ( .A(n2698), .B(n2697), .Z(n2699) );
  NAND U2941 ( .A(n2700), .B(n2699), .Z(n2774) );
  XNOR U2942 ( .A(n2775), .B(n2774), .Z(c[282]) );
  NANDN U2943 ( .A(n2702), .B(n2701), .Z(n2706) );
  NANDN U2944 ( .A(n2704), .B(n2703), .Z(n2705) );
  AND U2945 ( .A(n2706), .B(n2705), .Z(n2781) );
  NANDN U2946 ( .A(n2708), .B(n2707), .Z(n2712) );
  NAND U2947 ( .A(n2710), .B(n2709), .Z(n2711) );
  AND U2948 ( .A(n2712), .B(n2711), .Z(n2847) );
  NANDN U2949 ( .A(n2714), .B(n2713), .Z(n2718) );
  NANDN U2950 ( .A(n2716), .B(n2715), .Z(n2717) );
  AND U2951 ( .A(n2718), .B(n2717), .Z(n2813) );
  NAND U2952 ( .A(b[0]), .B(a[43]), .Z(n2719) );
  XNOR U2953 ( .A(b[1]), .B(n2719), .Z(n2721) );
  NANDN U2954 ( .A(b[0]), .B(a[42]), .Z(n2720) );
  NAND U2955 ( .A(n2721), .B(n2720), .Z(n2793) );
  NAND U2956 ( .A(n19808), .B(n2722), .Z(n2724) );
  XOR U2957 ( .A(b[13]), .B(a[31]), .Z(n2796) );
  NAND U2958 ( .A(n19768), .B(n2796), .Z(n2723) );
  AND U2959 ( .A(n2724), .B(n2723), .Z(n2791) );
  AND U2960 ( .A(b[15]), .B(a[27]), .Z(n2790) );
  XNOR U2961 ( .A(n2791), .B(n2790), .Z(n2792) );
  XNOR U2962 ( .A(n2793), .B(n2792), .Z(n2811) );
  NAND U2963 ( .A(n33), .B(n2725), .Z(n2727) );
  XOR U2964 ( .A(b[5]), .B(a[39]), .Z(n2802) );
  NAND U2965 ( .A(n19342), .B(n2802), .Z(n2726) );
  AND U2966 ( .A(n2727), .B(n2726), .Z(n2835) );
  NAND U2967 ( .A(n34), .B(n2728), .Z(n2730) );
  XOR U2968 ( .A(b[7]), .B(a[37]), .Z(n2805) );
  NAND U2969 ( .A(n19486), .B(n2805), .Z(n2729) );
  AND U2970 ( .A(n2730), .B(n2729), .Z(n2833) );
  NAND U2971 ( .A(n31), .B(n2731), .Z(n2733) );
  XOR U2972 ( .A(b[3]), .B(a[41]), .Z(n2808) );
  NAND U2973 ( .A(n32), .B(n2808), .Z(n2732) );
  NAND U2974 ( .A(n2733), .B(n2732), .Z(n2832) );
  XNOR U2975 ( .A(n2833), .B(n2832), .Z(n2834) );
  XOR U2976 ( .A(n2835), .B(n2834), .Z(n2812) );
  XOR U2977 ( .A(n2811), .B(n2812), .Z(n2814) );
  XOR U2978 ( .A(n2813), .B(n2814), .Z(n2785) );
  NANDN U2979 ( .A(n2735), .B(n2734), .Z(n2739) );
  OR U2980 ( .A(n2737), .B(n2736), .Z(n2738) );
  AND U2981 ( .A(n2739), .B(n2738), .Z(n2784) );
  XNOR U2982 ( .A(n2785), .B(n2784), .Z(n2787) );
  NAND U2983 ( .A(n2740), .B(n19724), .Z(n2742) );
  XOR U2984 ( .A(b[11]), .B(a[33]), .Z(n2817) );
  NAND U2985 ( .A(n19692), .B(n2817), .Z(n2741) );
  AND U2986 ( .A(n2742), .B(n2741), .Z(n2828) );
  NAND U2987 ( .A(n19838), .B(n2743), .Z(n2745) );
  XOR U2988 ( .A(b[15]), .B(a[29]), .Z(n2820) );
  NAND U2989 ( .A(n19805), .B(n2820), .Z(n2744) );
  AND U2990 ( .A(n2745), .B(n2744), .Z(n2827) );
  NAND U2991 ( .A(n35), .B(n2746), .Z(n2748) );
  XOR U2992 ( .A(b[9]), .B(a[35]), .Z(n2823) );
  NAND U2993 ( .A(n19598), .B(n2823), .Z(n2747) );
  NAND U2994 ( .A(n2748), .B(n2747), .Z(n2826) );
  XOR U2995 ( .A(n2827), .B(n2826), .Z(n2829) );
  XOR U2996 ( .A(n2828), .B(n2829), .Z(n2839) );
  NANDN U2997 ( .A(n2750), .B(n2749), .Z(n2754) );
  OR U2998 ( .A(n2752), .B(n2751), .Z(n2753) );
  AND U2999 ( .A(n2754), .B(n2753), .Z(n2838) );
  XNOR U3000 ( .A(n2839), .B(n2838), .Z(n2840) );
  NANDN U3001 ( .A(n2756), .B(n2755), .Z(n2760) );
  NANDN U3002 ( .A(n2758), .B(n2757), .Z(n2759) );
  NAND U3003 ( .A(n2760), .B(n2759), .Z(n2841) );
  XNOR U3004 ( .A(n2840), .B(n2841), .Z(n2786) );
  XOR U3005 ( .A(n2787), .B(n2786), .Z(n2845) );
  NANDN U3006 ( .A(n2762), .B(n2761), .Z(n2766) );
  NANDN U3007 ( .A(n2764), .B(n2763), .Z(n2765) );
  AND U3008 ( .A(n2766), .B(n2765), .Z(n2844) );
  XNOR U3009 ( .A(n2845), .B(n2844), .Z(n2846) );
  XOR U3010 ( .A(n2847), .B(n2846), .Z(n2779) );
  NANDN U3011 ( .A(n2768), .B(n2767), .Z(n2772) );
  NAND U3012 ( .A(n2770), .B(n2769), .Z(n2771) );
  AND U3013 ( .A(n2772), .B(n2771), .Z(n2778) );
  XNOR U3014 ( .A(n2779), .B(n2778), .Z(n2780) );
  XNOR U3015 ( .A(n2781), .B(n2780), .Z(n2850) );
  XNOR U3016 ( .A(sreg[283]), .B(n2850), .Z(n2852) );
  NANDN U3017 ( .A(sreg[282]), .B(n2773), .Z(n2777) );
  NAND U3018 ( .A(n2775), .B(n2774), .Z(n2776) );
  NAND U3019 ( .A(n2777), .B(n2776), .Z(n2851) );
  XNOR U3020 ( .A(n2852), .B(n2851), .Z(c[283]) );
  NANDN U3021 ( .A(n2779), .B(n2778), .Z(n2783) );
  NANDN U3022 ( .A(n2781), .B(n2780), .Z(n2782) );
  AND U3023 ( .A(n2783), .B(n2782), .Z(n2858) );
  NANDN U3024 ( .A(n2785), .B(n2784), .Z(n2789) );
  NAND U3025 ( .A(n2787), .B(n2786), .Z(n2788) );
  AND U3026 ( .A(n2789), .B(n2788), .Z(n2924) );
  NANDN U3027 ( .A(n2791), .B(n2790), .Z(n2795) );
  NANDN U3028 ( .A(n2793), .B(n2792), .Z(n2794) );
  AND U3029 ( .A(n2795), .B(n2794), .Z(n2890) );
  NAND U3030 ( .A(n19808), .B(n2796), .Z(n2798) );
  XOR U3031 ( .A(b[13]), .B(a[32]), .Z(n2876) );
  NAND U3032 ( .A(n19768), .B(n2876), .Z(n2797) );
  AND U3033 ( .A(n2798), .B(n2797), .Z(n2868) );
  AND U3034 ( .A(b[15]), .B(a[28]), .Z(n2867) );
  XNOR U3035 ( .A(n2868), .B(n2867), .Z(n2869) );
  NAND U3036 ( .A(b[0]), .B(a[44]), .Z(n2799) );
  XNOR U3037 ( .A(b[1]), .B(n2799), .Z(n2801) );
  NANDN U3038 ( .A(b[0]), .B(a[43]), .Z(n2800) );
  NAND U3039 ( .A(n2801), .B(n2800), .Z(n2870) );
  XNOR U3040 ( .A(n2869), .B(n2870), .Z(n2888) );
  NAND U3041 ( .A(n33), .B(n2802), .Z(n2804) );
  XOR U3042 ( .A(b[5]), .B(a[40]), .Z(n2879) );
  NAND U3043 ( .A(n19342), .B(n2879), .Z(n2803) );
  AND U3044 ( .A(n2804), .B(n2803), .Z(n2912) );
  NAND U3045 ( .A(n34), .B(n2805), .Z(n2807) );
  XOR U3046 ( .A(b[7]), .B(a[38]), .Z(n2882) );
  NAND U3047 ( .A(n19486), .B(n2882), .Z(n2806) );
  AND U3048 ( .A(n2807), .B(n2806), .Z(n2910) );
  NAND U3049 ( .A(n31), .B(n2808), .Z(n2810) );
  XOR U3050 ( .A(b[3]), .B(a[42]), .Z(n2885) );
  NAND U3051 ( .A(n32), .B(n2885), .Z(n2809) );
  NAND U3052 ( .A(n2810), .B(n2809), .Z(n2909) );
  XNOR U3053 ( .A(n2910), .B(n2909), .Z(n2911) );
  XOR U3054 ( .A(n2912), .B(n2911), .Z(n2889) );
  XOR U3055 ( .A(n2888), .B(n2889), .Z(n2891) );
  XOR U3056 ( .A(n2890), .B(n2891), .Z(n2862) );
  NANDN U3057 ( .A(n2812), .B(n2811), .Z(n2816) );
  OR U3058 ( .A(n2814), .B(n2813), .Z(n2815) );
  AND U3059 ( .A(n2816), .B(n2815), .Z(n2861) );
  XNOR U3060 ( .A(n2862), .B(n2861), .Z(n2864) );
  NAND U3061 ( .A(n2817), .B(n19724), .Z(n2819) );
  XOR U3062 ( .A(b[11]), .B(a[34]), .Z(n2894) );
  NAND U3063 ( .A(n19692), .B(n2894), .Z(n2818) );
  AND U3064 ( .A(n2819), .B(n2818), .Z(n2905) );
  NAND U3065 ( .A(n19838), .B(n2820), .Z(n2822) );
  XOR U3066 ( .A(b[15]), .B(a[30]), .Z(n2897) );
  NAND U3067 ( .A(n19805), .B(n2897), .Z(n2821) );
  AND U3068 ( .A(n2822), .B(n2821), .Z(n2904) );
  NAND U3069 ( .A(n35), .B(n2823), .Z(n2825) );
  XOR U3070 ( .A(b[9]), .B(a[36]), .Z(n2900) );
  NAND U3071 ( .A(n19598), .B(n2900), .Z(n2824) );
  NAND U3072 ( .A(n2825), .B(n2824), .Z(n2903) );
  XOR U3073 ( .A(n2904), .B(n2903), .Z(n2906) );
  XOR U3074 ( .A(n2905), .B(n2906), .Z(n2916) );
  NANDN U3075 ( .A(n2827), .B(n2826), .Z(n2831) );
  OR U3076 ( .A(n2829), .B(n2828), .Z(n2830) );
  AND U3077 ( .A(n2831), .B(n2830), .Z(n2915) );
  XNOR U3078 ( .A(n2916), .B(n2915), .Z(n2917) );
  NANDN U3079 ( .A(n2833), .B(n2832), .Z(n2837) );
  NANDN U3080 ( .A(n2835), .B(n2834), .Z(n2836) );
  NAND U3081 ( .A(n2837), .B(n2836), .Z(n2918) );
  XNOR U3082 ( .A(n2917), .B(n2918), .Z(n2863) );
  XOR U3083 ( .A(n2864), .B(n2863), .Z(n2922) );
  NANDN U3084 ( .A(n2839), .B(n2838), .Z(n2843) );
  NANDN U3085 ( .A(n2841), .B(n2840), .Z(n2842) );
  AND U3086 ( .A(n2843), .B(n2842), .Z(n2921) );
  XNOR U3087 ( .A(n2922), .B(n2921), .Z(n2923) );
  XOR U3088 ( .A(n2924), .B(n2923), .Z(n2856) );
  NANDN U3089 ( .A(n2845), .B(n2844), .Z(n2849) );
  NAND U3090 ( .A(n2847), .B(n2846), .Z(n2848) );
  AND U3091 ( .A(n2849), .B(n2848), .Z(n2855) );
  XNOR U3092 ( .A(n2856), .B(n2855), .Z(n2857) );
  XNOR U3093 ( .A(n2858), .B(n2857), .Z(n2927) );
  XNOR U3094 ( .A(sreg[284]), .B(n2927), .Z(n2929) );
  NANDN U3095 ( .A(sreg[283]), .B(n2850), .Z(n2854) );
  NAND U3096 ( .A(n2852), .B(n2851), .Z(n2853) );
  NAND U3097 ( .A(n2854), .B(n2853), .Z(n2928) );
  XNOR U3098 ( .A(n2929), .B(n2928), .Z(c[284]) );
  NANDN U3099 ( .A(n2856), .B(n2855), .Z(n2860) );
  NANDN U3100 ( .A(n2858), .B(n2857), .Z(n2859) );
  AND U3101 ( .A(n2860), .B(n2859), .Z(n2935) );
  NANDN U3102 ( .A(n2862), .B(n2861), .Z(n2866) );
  NAND U3103 ( .A(n2864), .B(n2863), .Z(n2865) );
  AND U3104 ( .A(n2866), .B(n2865), .Z(n3001) );
  NANDN U3105 ( .A(n2868), .B(n2867), .Z(n2872) );
  NANDN U3106 ( .A(n2870), .B(n2869), .Z(n2871) );
  AND U3107 ( .A(n2872), .B(n2871), .Z(n2967) );
  NAND U3108 ( .A(b[0]), .B(a[45]), .Z(n2873) );
  XNOR U3109 ( .A(b[1]), .B(n2873), .Z(n2875) );
  NANDN U3110 ( .A(b[0]), .B(a[44]), .Z(n2874) );
  NAND U3111 ( .A(n2875), .B(n2874), .Z(n2947) );
  NAND U3112 ( .A(n19808), .B(n2876), .Z(n2878) );
  XOR U3113 ( .A(b[13]), .B(a[33]), .Z(n2950) );
  NAND U3114 ( .A(n19768), .B(n2950), .Z(n2877) );
  AND U3115 ( .A(n2878), .B(n2877), .Z(n2945) );
  AND U3116 ( .A(b[15]), .B(a[29]), .Z(n2944) );
  XNOR U3117 ( .A(n2945), .B(n2944), .Z(n2946) );
  XNOR U3118 ( .A(n2947), .B(n2946), .Z(n2965) );
  NAND U3119 ( .A(n33), .B(n2879), .Z(n2881) );
  XOR U3120 ( .A(b[5]), .B(a[41]), .Z(n2956) );
  NAND U3121 ( .A(n19342), .B(n2956), .Z(n2880) );
  AND U3122 ( .A(n2881), .B(n2880), .Z(n2989) );
  NAND U3123 ( .A(n34), .B(n2882), .Z(n2884) );
  XOR U3124 ( .A(b[7]), .B(a[39]), .Z(n2959) );
  NAND U3125 ( .A(n19486), .B(n2959), .Z(n2883) );
  AND U3126 ( .A(n2884), .B(n2883), .Z(n2987) );
  NAND U3127 ( .A(n31), .B(n2885), .Z(n2887) );
  XOR U3128 ( .A(b[3]), .B(a[43]), .Z(n2962) );
  NAND U3129 ( .A(n32), .B(n2962), .Z(n2886) );
  NAND U3130 ( .A(n2887), .B(n2886), .Z(n2986) );
  XNOR U3131 ( .A(n2987), .B(n2986), .Z(n2988) );
  XOR U3132 ( .A(n2989), .B(n2988), .Z(n2966) );
  XOR U3133 ( .A(n2965), .B(n2966), .Z(n2968) );
  XOR U3134 ( .A(n2967), .B(n2968), .Z(n2939) );
  NANDN U3135 ( .A(n2889), .B(n2888), .Z(n2893) );
  OR U3136 ( .A(n2891), .B(n2890), .Z(n2892) );
  AND U3137 ( .A(n2893), .B(n2892), .Z(n2938) );
  XNOR U3138 ( .A(n2939), .B(n2938), .Z(n2941) );
  NAND U3139 ( .A(n2894), .B(n19724), .Z(n2896) );
  XOR U3140 ( .A(b[11]), .B(a[35]), .Z(n2971) );
  NAND U3141 ( .A(n19692), .B(n2971), .Z(n2895) );
  AND U3142 ( .A(n2896), .B(n2895), .Z(n2982) );
  NAND U3143 ( .A(n19838), .B(n2897), .Z(n2899) );
  XOR U3144 ( .A(b[15]), .B(a[31]), .Z(n2974) );
  NAND U3145 ( .A(n19805), .B(n2974), .Z(n2898) );
  AND U3146 ( .A(n2899), .B(n2898), .Z(n2981) );
  NAND U3147 ( .A(n35), .B(n2900), .Z(n2902) );
  XOR U3148 ( .A(b[9]), .B(a[37]), .Z(n2977) );
  NAND U3149 ( .A(n19598), .B(n2977), .Z(n2901) );
  NAND U3150 ( .A(n2902), .B(n2901), .Z(n2980) );
  XOR U3151 ( .A(n2981), .B(n2980), .Z(n2983) );
  XOR U3152 ( .A(n2982), .B(n2983), .Z(n2993) );
  NANDN U3153 ( .A(n2904), .B(n2903), .Z(n2908) );
  OR U3154 ( .A(n2906), .B(n2905), .Z(n2907) );
  AND U3155 ( .A(n2908), .B(n2907), .Z(n2992) );
  XNOR U3156 ( .A(n2993), .B(n2992), .Z(n2994) );
  NANDN U3157 ( .A(n2910), .B(n2909), .Z(n2914) );
  NANDN U3158 ( .A(n2912), .B(n2911), .Z(n2913) );
  NAND U3159 ( .A(n2914), .B(n2913), .Z(n2995) );
  XNOR U3160 ( .A(n2994), .B(n2995), .Z(n2940) );
  XOR U3161 ( .A(n2941), .B(n2940), .Z(n2999) );
  NANDN U3162 ( .A(n2916), .B(n2915), .Z(n2920) );
  NANDN U3163 ( .A(n2918), .B(n2917), .Z(n2919) );
  AND U3164 ( .A(n2920), .B(n2919), .Z(n2998) );
  XNOR U3165 ( .A(n2999), .B(n2998), .Z(n3000) );
  XOR U3166 ( .A(n3001), .B(n3000), .Z(n2933) );
  NANDN U3167 ( .A(n2922), .B(n2921), .Z(n2926) );
  NAND U3168 ( .A(n2924), .B(n2923), .Z(n2925) );
  AND U3169 ( .A(n2926), .B(n2925), .Z(n2932) );
  XNOR U3170 ( .A(n2933), .B(n2932), .Z(n2934) );
  XNOR U3171 ( .A(n2935), .B(n2934), .Z(n3004) );
  XNOR U3172 ( .A(sreg[285]), .B(n3004), .Z(n3006) );
  NANDN U3173 ( .A(sreg[284]), .B(n2927), .Z(n2931) );
  NAND U3174 ( .A(n2929), .B(n2928), .Z(n2930) );
  NAND U3175 ( .A(n2931), .B(n2930), .Z(n3005) );
  XNOR U3176 ( .A(n3006), .B(n3005), .Z(c[285]) );
  NANDN U3177 ( .A(n2933), .B(n2932), .Z(n2937) );
  NANDN U3178 ( .A(n2935), .B(n2934), .Z(n2936) );
  AND U3179 ( .A(n2937), .B(n2936), .Z(n3012) );
  NANDN U3180 ( .A(n2939), .B(n2938), .Z(n2943) );
  NAND U3181 ( .A(n2941), .B(n2940), .Z(n2942) );
  AND U3182 ( .A(n2943), .B(n2942), .Z(n3078) );
  NANDN U3183 ( .A(n2945), .B(n2944), .Z(n2949) );
  NANDN U3184 ( .A(n2947), .B(n2946), .Z(n2948) );
  AND U3185 ( .A(n2949), .B(n2948), .Z(n3065) );
  NAND U3186 ( .A(n19808), .B(n2950), .Z(n2952) );
  XOR U3187 ( .A(b[13]), .B(a[34]), .Z(n3051) );
  NAND U3188 ( .A(n19768), .B(n3051), .Z(n2951) );
  AND U3189 ( .A(n2952), .B(n2951), .Z(n3043) );
  AND U3190 ( .A(b[15]), .B(a[30]), .Z(n3042) );
  XNOR U3191 ( .A(n3043), .B(n3042), .Z(n3044) );
  NAND U3192 ( .A(b[0]), .B(a[46]), .Z(n2953) );
  XNOR U3193 ( .A(b[1]), .B(n2953), .Z(n2955) );
  NANDN U3194 ( .A(b[0]), .B(a[45]), .Z(n2954) );
  NAND U3195 ( .A(n2955), .B(n2954), .Z(n3045) );
  XNOR U3196 ( .A(n3044), .B(n3045), .Z(n3063) );
  NAND U3197 ( .A(n33), .B(n2956), .Z(n2958) );
  XOR U3198 ( .A(b[5]), .B(a[42]), .Z(n3054) );
  NAND U3199 ( .A(n19342), .B(n3054), .Z(n2957) );
  AND U3200 ( .A(n2958), .B(n2957), .Z(n3039) );
  NAND U3201 ( .A(n34), .B(n2959), .Z(n2961) );
  XOR U3202 ( .A(b[7]), .B(a[40]), .Z(n3057) );
  NAND U3203 ( .A(n19486), .B(n3057), .Z(n2960) );
  AND U3204 ( .A(n2961), .B(n2960), .Z(n3037) );
  NAND U3205 ( .A(n31), .B(n2962), .Z(n2964) );
  XOR U3206 ( .A(b[3]), .B(a[44]), .Z(n3060) );
  NAND U3207 ( .A(n32), .B(n3060), .Z(n2963) );
  NAND U3208 ( .A(n2964), .B(n2963), .Z(n3036) );
  XNOR U3209 ( .A(n3037), .B(n3036), .Z(n3038) );
  XOR U3210 ( .A(n3039), .B(n3038), .Z(n3064) );
  XOR U3211 ( .A(n3063), .B(n3064), .Z(n3066) );
  XOR U3212 ( .A(n3065), .B(n3066), .Z(n3016) );
  NANDN U3213 ( .A(n2966), .B(n2965), .Z(n2970) );
  OR U3214 ( .A(n2968), .B(n2967), .Z(n2969) );
  AND U3215 ( .A(n2970), .B(n2969), .Z(n3015) );
  XNOR U3216 ( .A(n3016), .B(n3015), .Z(n3018) );
  NAND U3217 ( .A(n2971), .B(n19724), .Z(n2973) );
  XOR U3218 ( .A(b[11]), .B(a[36]), .Z(n3021) );
  NAND U3219 ( .A(n19692), .B(n3021), .Z(n2972) );
  AND U3220 ( .A(n2973), .B(n2972), .Z(n3032) );
  NAND U3221 ( .A(n19838), .B(n2974), .Z(n2976) );
  XOR U3222 ( .A(b[15]), .B(a[32]), .Z(n3024) );
  NAND U3223 ( .A(n19805), .B(n3024), .Z(n2975) );
  AND U3224 ( .A(n2976), .B(n2975), .Z(n3031) );
  NAND U3225 ( .A(n35), .B(n2977), .Z(n2979) );
  XOR U3226 ( .A(b[9]), .B(a[38]), .Z(n3027) );
  NAND U3227 ( .A(n19598), .B(n3027), .Z(n2978) );
  NAND U3228 ( .A(n2979), .B(n2978), .Z(n3030) );
  XOR U3229 ( .A(n3031), .B(n3030), .Z(n3033) );
  XOR U3230 ( .A(n3032), .B(n3033), .Z(n3070) );
  NANDN U3231 ( .A(n2981), .B(n2980), .Z(n2985) );
  OR U3232 ( .A(n2983), .B(n2982), .Z(n2984) );
  AND U3233 ( .A(n2985), .B(n2984), .Z(n3069) );
  XNOR U3234 ( .A(n3070), .B(n3069), .Z(n3071) );
  NANDN U3235 ( .A(n2987), .B(n2986), .Z(n2991) );
  NANDN U3236 ( .A(n2989), .B(n2988), .Z(n2990) );
  NAND U3237 ( .A(n2991), .B(n2990), .Z(n3072) );
  XNOR U3238 ( .A(n3071), .B(n3072), .Z(n3017) );
  XOR U3239 ( .A(n3018), .B(n3017), .Z(n3076) );
  NANDN U3240 ( .A(n2993), .B(n2992), .Z(n2997) );
  NANDN U3241 ( .A(n2995), .B(n2994), .Z(n2996) );
  AND U3242 ( .A(n2997), .B(n2996), .Z(n3075) );
  XNOR U3243 ( .A(n3076), .B(n3075), .Z(n3077) );
  XOR U3244 ( .A(n3078), .B(n3077), .Z(n3010) );
  NANDN U3245 ( .A(n2999), .B(n2998), .Z(n3003) );
  NAND U3246 ( .A(n3001), .B(n3000), .Z(n3002) );
  AND U3247 ( .A(n3003), .B(n3002), .Z(n3009) );
  XNOR U3248 ( .A(n3010), .B(n3009), .Z(n3011) );
  XNOR U3249 ( .A(n3012), .B(n3011), .Z(n3081) );
  XNOR U3250 ( .A(sreg[286]), .B(n3081), .Z(n3083) );
  NANDN U3251 ( .A(sreg[285]), .B(n3004), .Z(n3008) );
  NAND U3252 ( .A(n3006), .B(n3005), .Z(n3007) );
  NAND U3253 ( .A(n3008), .B(n3007), .Z(n3082) );
  XNOR U3254 ( .A(n3083), .B(n3082), .Z(c[286]) );
  NANDN U3255 ( .A(n3010), .B(n3009), .Z(n3014) );
  NANDN U3256 ( .A(n3012), .B(n3011), .Z(n3013) );
  AND U3257 ( .A(n3014), .B(n3013), .Z(n3089) );
  NANDN U3258 ( .A(n3016), .B(n3015), .Z(n3020) );
  NAND U3259 ( .A(n3018), .B(n3017), .Z(n3019) );
  AND U3260 ( .A(n3020), .B(n3019), .Z(n3155) );
  NAND U3261 ( .A(n3021), .B(n19724), .Z(n3023) );
  XOR U3262 ( .A(b[11]), .B(a[37]), .Z(n3125) );
  NAND U3263 ( .A(n19692), .B(n3125), .Z(n3022) );
  AND U3264 ( .A(n3023), .B(n3022), .Z(n3136) );
  NAND U3265 ( .A(n19838), .B(n3024), .Z(n3026) );
  XOR U3266 ( .A(b[15]), .B(a[33]), .Z(n3128) );
  NAND U3267 ( .A(n19805), .B(n3128), .Z(n3025) );
  AND U3268 ( .A(n3026), .B(n3025), .Z(n3135) );
  NAND U3269 ( .A(n35), .B(n3027), .Z(n3029) );
  XOR U3270 ( .A(b[9]), .B(a[39]), .Z(n3131) );
  NAND U3271 ( .A(n19598), .B(n3131), .Z(n3028) );
  NAND U3272 ( .A(n3029), .B(n3028), .Z(n3134) );
  XOR U3273 ( .A(n3135), .B(n3134), .Z(n3137) );
  XOR U3274 ( .A(n3136), .B(n3137), .Z(n3147) );
  NANDN U3275 ( .A(n3031), .B(n3030), .Z(n3035) );
  OR U3276 ( .A(n3033), .B(n3032), .Z(n3034) );
  AND U3277 ( .A(n3035), .B(n3034), .Z(n3146) );
  XNOR U3278 ( .A(n3147), .B(n3146), .Z(n3148) );
  NANDN U3279 ( .A(n3037), .B(n3036), .Z(n3041) );
  NANDN U3280 ( .A(n3039), .B(n3038), .Z(n3040) );
  NAND U3281 ( .A(n3041), .B(n3040), .Z(n3149) );
  XNOR U3282 ( .A(n3148), .B(n3149), .Z(n3095) );
  NANDN U3283 ( .A(n3043), .B(n3042), .Z(n3047) );
  NANDN U3284 ( .A(n3045), .B(n3044), .Z(n3046) );
  AND U3285 ( .A(n3047), .B(n3046), .Z(n3121) );
  AND U3286 ( .A(b[0]), .B(a[47]), .Z(n3048) );
  XOR U3287 ( .A(b[1]), .B(n3048), .Z(n3050) );
  NANDN U3288 ( .A(b[0]), .B(a[46]), .Z(n3049) );
  AND U3289 ( .A(n3050), .B(n3049), .Z(n3100) );
  NAND U3290 ( .A(n19808), .B(n3051), .Z(n3053) );
  XOR U3291 ( .A(b[13]), .B(a[35]), .Z(n3104) );
  NAND U3292 ( .A(n19768), .B(n3104), .Z(n3052) );
  AND U3293 ( .A(n3053), .B(n3052), .Z(n3099) );
  AND U3294 ( .A(b[15]), .B(a[31]), .Z(n3098) );
  XOR U3295 ( .A(n3099), .B(n3098), .Z(n3101) );
  XNOR U3296 ( .A(n3100), .B(n3101), .Z(n3119) );
  NAND U3297 ( .A(n33), .B(n3054), .Z(n3056) );
  XOR U3298 ( .A(b[5]), .B(a[43]), .Z(n3110) );
  NAND U3299 ( .A(n19342), .B(n3110), .Z(n3055) );
  AND U3300 ( .A(n3056), .B(n3055), .Z(n3143) );
  NAND U3301 ( .A(n34), .B(n3057), .Z(n3059) );
  XOR U3302 ( .A(b[7]), .B(a[41]), .Z(n3113) );
  NAND U3303 ( .A(n19486), .B(n3113), .Z(n3058) );
  AND U3304 ( .A(n3059), .B(n3058), .Z(n3141) );
  NAND U3305 ( .A(n31), .B(n3060), .Z(n3062) );
  XOR U3306 ( .A(b[3]), .B(a[45]), .Z(n3116) );
  NAND U3307 ( .A(n32), .B(n3116), .Z(n3061) );
  NAND U3308 ( .A(n3062), .B(n3061), .Z(n3140) );
  XNOR U3309 ( .A(n3141), .B(n3140), .Z(n3142) );
  XOR U3310 ( .A(n3143), .B(n3142), .Z(n3120) );
  XOR U3311 ( .A(n3119), .B(n3120), .Z(n3122) );
  XOR U3312 ( .A(n3121), .B(n3122), .Z(n3093) );
  NANDN U3313 ( .A(n3064), .B(n3063), .Z(n3068) );
  OR U3314 ( .A(n3066), .B(n3065), .Z(n3067) );
  AND U3315 ( .A(n3068), .B(n3067), .Z(n3092) );
  XNOR U3316 ( .A(n3093), .B(n3092), .Z(n3094) );
  XOR U3317 ( .A(n3095), .B(n3094), .Z(n3153) );
  NANDN U3318 ( .A(n3070), .B(n3069), .Z(n3074) );
  NANDN U3319 ( .A(n3072), .B(n3071), .Z(n3073) );
  AND U3320 ( .A(n3074), .B(n3073), .Z(n3152) );
  XNOR U3321 ( .A(n3153), .B(n3152), .Z(n3154) );
  XOR U3322 ( .A(n3155), .B(n3154), .Z(n3087) );
  NANDN U3323 ( .A(n3076), .B(n3075), .Z(n3080) );
  NAND U3324 ( .A(n3078), .B(n3077), .Z(n3079) );
  AND U3325 ( .A(n3080), .B(n3079), .Z(n3086) );
  XNOR U3326 ( .A(n3087), .B(n3086), .Z(n3088) );
  XNOR U3327 ( .A(n3089), .B(n3088), .Z(n3158) );
  XNOR U3328 ( .A(sreg[287]), .B(n3158), .Z(n3160) );
  NANDN U3329 ( .A(sreg[286]), .B(n3081), .Z(n3085) );
  NAND U3330 ( .A(n3083), .B(n3082), .Z(n3084) );
  NAND U3331 ( .A(n3085), .B(n3084), .Z(n3159) );
  XNOR U3332 ( .A(n3160), .B(n3159), .Z(c[287]) );
  NANDN U3333 ( .A(n3087), .B(n3086), .Z(n3091) );
  NANDN U3334 ( .A(n3089), .B(n3088), .Z(n3090) );
  AND U3335 ( .A(n3091), .B(n3090), .Z(n3166) );
  NANDN U3336 ( .A(n3093), .B(n3092), .Z(n3097) );
  NAND U3337 ( .A(n3095), .B(n3094), .Z(n3096) );
  AND U3338 ( .A(n3097), .B(n3096), .Z(n3232) );
  NANDN U3339 ( .A(n3099), .B(n3098), .Z(n3103) );
  NANDN U3340 ( .A(n3101), .B(n3100), .Z(n3102) );
  AND U3341 ( .A(n3103), .B(n3102), .Z(n3198) );
  NAND U3342 ( .A(n19808), .B(n3104), .Z(n3106) );
  XOR U3343 ( .A(b[13]), .B(a[36]), .Z(n3184) );
  NAND U3344 ( .A(n19768), .B(n3184), .Z(n3105) );
  AND U3345 ( .A(n3106), .B(n3105), .Z(n3176) );
  AND U3346 ( .A(b[15]), .B(a[32]), .Z(n3175) );
  XNOR U3347 ( .A(n3176), .B(n3175), .Z(n3177) );
  NAND U3348 ( .A(b[0]), .B(a[48]), .Z(n3107) );
  XNOR U3349 ( .A(b[1]), .B(n3107), .Z(n3109) );
  NANDN U3350 ( .A(b[0]), .B(a[47]), .Z(n3108) );
  NAND U3351 ( .A(n3109), .B(n3108), .Z(n3178) );
  XNOR U3352 ( .A(n3177), .B(n3178), .Z(n3196) );
  NAND U3353 ( .A(n33), .B(n3110), .Z(n3112) );
  XOR U3354 ( .A(b[5]), .B(a[44]), .Z(n3187) );
  NAND U3355 ( .A(n19342), .B(n3187), .Z(n3111) );
  AND U3356 ( .A(n3112), .B(n3111), .Z(n3220) );
  NAND U3357 ( .A(n34), .B(n3113), .Z(n3115) );
  XOR U3358 ( .A(b[7]), .B(a[42]), .Z(n3190) );
  NAND U3359 ( .A(n19486), .B(n3190), .Z(n3114) );
  AND U3360 ( .A(n3115), .B(n3114), .Z(n3218) );
  NAND U3361 ( .A(n31), .B(n3116), .Z(n3118) );
  XOR U3362 ( .A(b[3]), .B(a[46]), .Z(n3193) );
  NAND U3363 ( .A(n32), .B(n3193), .Z(n3117) );
  NAND U3364 ( .A(n3118), .B(n3117), .Z(n3217) );
  XNOR U3365 ( .A(n3218), .B(n3217), .Z(n3219) );
  XOR U3366 ( .A(n3220), .B(n3219), .Z(n3197) );
  XOR U3367 ( .A(n3196), .B(n3197), .Z(n3199) );
  XOR U3368 ( .A(n3198), .B(n3199), .Z(n3170) );
  NANDN U3369 ( .A(n3120), .B(n3119), .Z(n3124) );
  OR U3370 ( .A(n3122), .B(n3121), .Z(n3123) );
  AND U3371 ( .A(n3124), .B(n3123), .Z(n3169) );
  XNOR U3372 ( .A(n3170), .B(n3169), .Z(n3172) );
  NAND U3373 ( .A(n3125), .B(n19724), .Z(n3127) );
  XOR U3374 ( .A(b[11]), .B(a[38]), .Z(n3202) );
  NAND U3375 ( .A(n19692), .B(n3202), .Z(n3126) );
  AND U3376 ( .A(n3127), .B(n3126), .Z(n3213) );
  NAND U3377 ( .A(n19838), .B(n3128), .Z(n3130) );
  XOR U3378 ( .A(b[15]), .B(a[34]), .Z(n3205) );
  NAND U3379 ( .A(n19805), .B(n3205), .Z(n3129) );
  AND U3380 ( .A(n3130), .B(n3129), .Z(n3212) );
  NAND U3381 ( .A(n35), .B(n3131), .Z(n3133) );
  XOR U3382 ( .A(b[9]), .B(a[40]), .Z(n3208) );
  NAND U3383 ( .A(n19598), .B(n3208), .Z(n3132) );
  NAND U3384 ( .A(n3133), .B(n3132), .Z(n3211) );
  XOR U3385 ( .A(n3212), .B(n3211), .Z(n3214) );
  XOR U3386 ( .A(n3213), .B(n3214), .Z(n3224) );
  NANDN U3387 ( .A(n3135), .B(n3134), .Z(n3139) );
  OR U3388 ( .A(n3137), .B(n3136), .Z(n3138) );
  AND U3389 ( .A(n3139), .B(n3138), .Z(n3223) );
  XNOR U3390 ( .A(n3224), .B(n3223), .Z(n3225) );
  NANDN U3391 ( .A(n3141), .B(n3140), .Z(n3145) );
  NANDN U3392 ( .A(n3143), .B(n3142), .Z(n3144) );
  NAND U3393 ( .A(n3145), .B(n3144), .Z(n3226) );
  XNOR U3394 ( .A(n3225), .B(n3226), .Z(n3171) );
  XOR U3395 ( .A(n3172), .B(n3171), .Z(n3230) );
  NANDN U3396 ( .A(n3147), .B(n3146), .Z(n3151) );
  NANDN U3397 ( .A(n3149), .B(n3148), .Z(n3150) );
  AND U3398 ( .A(n3151), .B(n3150), .Z(n3229) );
  XNOR U3399 ( .A(n3230), .B(n3229), .Z(n3231) );
  XOR U3400 ( .A(n3232), .B(n3231), .Z(n3164) );
  NANDN U3401 ( .A(n3153), .B(n3152), .Z(n3157) );
  NAND U3402 ( .A(n3155), .B(n3154), .Z(n3156) );
  AND U3403 ( .A(n3157), .B(n3156), .Z(n3163) );
  XNOR U3404 ( .A(n3164), .B(n3163), .Z(n3165) );
  XNOR U3405 ( .A(n3166), .B(n3165), .Z(n3235) );
  XNOR U3406 ( .A(sreg[288]), .B(n3235), .Z(n3237) );
  NANDN U3407 ( .A(sreg[287]), .B(n3158), .Z(n3162) );
  NAND U3408 ( .A(n3160), .B(n3159), .Z(n3161) );
  NAND U3409 ( .A(n3162), .B(n3161), .Z(n3236) );
  XNOR U3410 ( .A(n3237), .B(n3236), .Z(c[288]) );
  NANDN U3411 ( .A(n3164), .B(n3163), .Z(n3168) );
  NANDN U3412 ( .A(n3166), .B(n3165), .Z(n3167) );
  AND U3413 ( .A(n3168), .B(n3167), .Z(n3243) );
  NANDN U3414 ( .A(n3170), .B(n3169), .Z(n3174) );
  NAND U3415 ( .A(n3172), .B(n3171), .Z(n3173) );
  AND U3416 ( .A(n3174), .B(n3173), .Z(n3309) );
  NANDN U3417 ( .A(n3176), .B(n3175), .Z(n3180) );
  NANDN U3418 ( .A(n3178), .B(n3177), .Z(n3179) );
  AND U3419 ( .A(n3180), .B(n3179), .Z(n3275) );
  NAND U3420 ( .A(b[0]), .B(a[49]), .Z(n3181) );
  XNOR U3421 ( .A(b[1]), .B(n3181), .Z(n3183) );
  NANDN U3422 ( .A(b[0]), .B(a[48]), .Z(n3182) );
  NAND U3423 ( .A(n3183), .B(n3182), .Z(n3255) );
  NAND U3424 ( .A(n19808), .B(n3184), .Z(n3186) );
  XOR U3425 ( .A(b[13]), .B(a[37]), .Z(n3258) );
  NAND U3426 ( .A(n19768), .B(n3258), .Z(n3185) );
  AND U3427 ( .A(n3186), .B(n3185), .Z(n3253) );
  AND U3428 ( .A(b[15]), .B(a[33]), .Z(n3252) );
  XNOR U3429 ( .A(n3253), .B(n3252), .Z(n3254) );
  XNOR U3430 ( .A(n3255), .B(n3254), .Z(n3273) );
  NAND U3431 ( .A(n33), .B(n3187), .Z(n3189) );
  XOR U3432 ( .A(b[5]), .B(a[45]), .Z(n3264) );
  NAND U3433 ( .A(n19342), .B(n3264), .Z(n3188) );
  AND U3434 ( .A(n3189), .B(n3188), .Z(n3297) );
  NAND U3435 ( .A(n34), .B(n3190), .Z(n3192) );
  XOR U3436 ( .A(b[7]), .B(a[43]), .Z(n3267) );
  NAND U3437 ( .A(n19486), .B(n3267), .Z(n3191) );
  AND U3438 ( .A(n3192), .B(n3191), .Z(n3295) );
  NAND U3439 ( .A(n31), .B(n3193), .Z(n3195) );
  XOR U3440 ( .A(b[3]), .B(a[47]), .Z(n3270) );
  NAND U3441 ( .A(n32), .B(n3270), .Z(n3194) );
  NAND U3442 ( .A(n3195), .B(n3194), .Z(n3294) );
  XNOR U3443 ( .A(n3295), .B(n3294), .Z(n3296) );
  XOR U3444 ( .A(n3297), .B(n3296), .Z(n3274) );
  XOR U3445 ( .A(n3273), .B(n3274), .Z(n3276) );
  XOR U3446 ( .A(n3275), .B(n3276), .Z(n3247) );
  NANDN U3447 ( .A(n3197), .B(n3196), .Z(n3201) );
  OR U3448 ( .A(n3199), .B(n3198), .Z(n3200) );
  AND U3449 ( .A(n3201), .B(n3200), .Z(n3246) );
  XNOR U3450 ( .A(n3247), .B(n3246), .Z(n3249) );
  NAND U3451 ( .A(n3202), .B(n19724), .Z(n3204) );
  XOR U3452 ( .A(b[11]), .B(a[39]), .Z(n3279) );
  NAND U3453 ( .A(n19692), .B(n3279), .Z(n3203) );
  AND U3454 ( .A(n3204), .B(n3203), .Z(n3290) );
  NAND U3455 ( .A(n19838), .B(n3205), .Z(n3207) );
  XOR U3456 ( .A(b[15]), .B(a[35]), .Z(n3282) );
  NAND U3457 ( .A(n19805), .B(n3282), .Z(n3206) );
  AND U3458 ( .A(n3207), .B(n3206), .Z(n3289) );
  NAND U3459 ( .A(n35), .B(n3208), .Z(n3210) );
  XOR U3460 ( .A(b[9]), .B(a[41]), .Z(n3285) );
  NAND U3461 ( .A(n19598), .B(n3285), .Z(n3209) );
  NAND U3462 ( .A(n3210), .B(n3209), .Z(n3288) );
  XOR U3463 ( .A(n3289), .B(n3288), .Z(n3291) );
  XOR U3464 ( .A(n3290), .B(n3291), .Z(n3301) );
  NANDN U3465 ( .A(n3212), .B(n3211), .Z(n3216) );
  OR U3466 ( .A(n3214), .B(n3213), .Z(n3215) );
  AND U3467 ( .A(n3216), .B(n3215), .Z(n3300) );
  XNOR U3468 ( .A(n3301), .B(n3300), .Z(n3302) );
  NANDN U3469 ( .A(n3218), .B(n3217), .Z(n3222) );
  NANDN U3470 ( .A(n3220), .B(n3219), .Z(n3221) );
  NAND U3471 ( .A(n3222), .B(n3221), .Z(n3303) );
  XNOR U3472 ( .A(n3302), .B(n3303), .Z(n3248) );
  XOR U3473 ( .A(n3249), .B(n3248), .Z(n3307) );
  NANDN U3474 ( .A(n3224), .B(n3223), .Z(n3228) );
  NANDN U3475 ( .A(n3226), .B(n3225), .Z(n3227) );
  AND U3476 ( .A(n3228), .B(n3227), .Z(n3306) );
  XNOR U3477 ( .A(n3307), .B(n3306), .Z(n3308) );
  XOR U3478 ( .A(n3309), .B(n3308), .Z(n3241) );
  NANDN U3479 ( .A(n3230), .B(n3229), .Z(n3234) );
  NAND U3480 ( .A(n3232), .B(n3231), .Z(n3233) );
  AND U3481 ( .A(n3234), .B(n3233), .Z(n3240) );
  XNOR U3482 ( .A(n3241), .B(n3240), .Z(n3242) );
  XNOR U3483 ( .A(n3243), .B(n3242), .Z(n3312) );
  XNOR U3484 ( .A(sreg[289]), .B(n3312), .Z(n3314) );
  NANDN U3485 ( .A(sreg[288]), .B(n3235), .Z(n3239) );
  NAND U3486 ( .A(n3237), .B(n3236), .Z(n3238) );
  NAND U3487 ( .A(n3239), .B(n3238), .Z(n3313) );
  XNOR U3488 ( .A(n3314), .B(n3313), .Z(c[289]) );
  NANDN U3489 ( .A(n3241), .B(n3240), .Z(n3245) );
  NANDN U3490 ( .A(n3243), .B(n3242), .Z(n3244) );
  AND U3491 ( .A(n3245), .B(n3244), .Z(n3320) );
  NANDN U3492 ( .A(n3247), .B(n3246), .Z(n3251) );
  NAND U3493 ( .A(n3249), .B(n3248), .Z(n3250) );
  AND U3494 ( .A(n3251), .B(n3250), .Z(n3386) );
  NANDN U3495 ( .A(n3253), .B(n3252), .Z(n3257) );
  NANDN U3496 ( .A(n3255), .B(n3254), .Z(n3256) );
  AND U3497 ( .A(n3257), .B(n3256), .Z(n3352) );
  NAND U3498 ( .A(n19808), .B(n3258), .Z(n3260) );
  XOR U3499 ( .A(b[13]), .B(a[38]), .Z(n3338) );
  NAND U3500 ( .A(n19768), .B(n3338), .Z(n3259) );
  AND U3501 ( .A(n3260), .B(n3259), .Z(n3330) );
  AND U3502 ( .A(b[15]), .B(a[34]), .Z(n3329) );
  XNOR U3503 ( .A(n3330), .B(n3329), .Z(n3331) );
  NAND U3504 ( .A(b[0]), .B(a[50]), .Z(n3261) );
  XNOR U3505 ( .A(b[1]), .B(n3261), .Z(n3263) );
  NANDN U3506 ( .A(b[0]), .B(a[49]), .Z(n3262) );
  NAND U3507 ( .A(n3263), .B(n3262), .Z(n3332) );
  XNOR U3508 ( .A(n3331), .B(n3332), .Z(n3350) );
  NAND U3509 ( .A(n33), .B(n3264), .Z(n3266) );
  XOR U3510 ( .A(b[5]), .B(a[46]), .Z(n3341) );
  NAND U3511 ( .A(n19342), .B(n3341), .Z(n3265) );
  AND U3512 ( .A(n3266), .B(n3265), .Z(n3374) );
  NAND U3513 ( .A(n34), .B(n3267), .Z(n3269) );
  XOR U3514 ( .A(b[7]), .B(a[44]), .Z(n3344) );
  NAND U3515 ( .A(n19486), .B(n3344), .Z(n3268) );
  AND U3516 ( .A(n3269), .B(n3268), .Z(n3372) );
  NAND U3517 ( .A(n31), .B(n3270), .Z(n3272) );
  XOR U3518 ( .A(b[3]), .B(a[48]), .Z(n3347) );
  NAND U3519 ( .A(n32), .B(n3347), .Z(n3271) );
  NAND U3520 ( .A(n3272), .B(n3271), .Z(n3371) );
  XNOR U3521 ( .A(n3372), .B(n3371), .Z(n3373) );
  XOR U3522 ( .A(n3374), .B(n3373), .Z(n3351) );
  XOR U3523 ( .A(n3350), .B(n3351), .Z(n3353) );
  XOR U3524 ( .A(n3352), .B(n3353), .Z(n3324) );
  NANDN U3525 ( .A(n3274), .B(n3273), .Z(n3278) );
  OR U3526 ( .A(n3276), .B(n3275), .Z(n3277) );
  AND U3527 ( .A(n3278), .B(n3277), .Z(n3323) );
  XNOR U3528 ( .A(n3324), .B(n3323), .Z(n3326) );
  NAND U3529 ( .A(n3279), .B(n19724), .Z(n3281) );
  XOR U3530 ( .A(b[11]), .B(a[40]), .Z(n3356) );
  NAND U3531 ( .A(n19692), .B(n3356), .Z(n3280) );
  AND U3532 ( .A(n3281), .B(n3280), .Z(n3367) );
  NAND U3533 ( .A(n19838), .B(n3282), .Z(n3284) );
  XOR U3534 ( .A(b[15]), .B(a[36]), .Z(n3359) );
  NAND U3535 ( .A(n19805), .B(n3359), .Z(n3283) );
  AND U3536 ( .A(n3284), .B(n3283), .Z(n3366) );
  NAND U3537 ( .A(n35), .B(n3285), .Z(n3287) );
  XOR U3538 ( .A(b[9]), .B(a[42]), .Z(n3362) );
  NAND U3539 ( .A(n19598), .B(n3362), .Z(n3286) );
  NAND U3540 ( .A(n3287), .B(n3286), .Z(n3365) );
  XOR U3541 ( .A(n3366), .B(n3365), .Z(n3368) );
  XOR U3542 ( .A(n3367), .B(n3368), .Z(n3378) );
  NANDN U3543 ( .A(n3289), .B(n3288), .Z(n3293) );
  OR U3544 ( .A(n3291), .B(n3290), .Z(n3292) );
  AND U3545 ( .A(n3293), .B(n3292), .Z(n3377) );
  XNOR U3546 ( .A(n3378), .B(n3377), .Z(n3379) );
  NANDN U3547 ( .A(n3295), .B(n3294), .Z(n3299) );
  NANDN U3548 ( .A(n3297), .B(n3296), .Z(n3298) );
  NAND U3549 ( .A(n3299), .B(n3298), .Z(n3380) );
  XNOR U3550 ( .A(n3379), .B(n3380), .Z(n3325) );
  XOR U3551 ( .A(n3326), .B(n3325), .Z(n3384) );
  NANDN U3552 ( .A(n3301), .B(n3300), .Z(n3305) );
  NANDN U3553 ( .A(n3303), .B(n3302), .Z(n3304) );
  AND U3554 ( .A(n3305), .B(n3304), .Z(n3383) );
  XNOR U3555 ( .A(n3384), .B(n3383), .Z(n3385) );
  XOR U3556 ( .A(n3386), .B(n3385), .Z(n3318) );
  NANDN U3557 ( .A(n3307), .B(n3306), .Z(n3311) );
  NAND U3558 ( .A(n3309), .B(n3308), .Z(n3310) );
  AND U3559 ( .A(n3311), .B(n3310), .Z(n3317) );
  XNOR U3560 ( .A(n3318), .B(n3317), .Z(n3319) );
  XNOR U3561 ( .A(n3320), .B(n3319), .Z(n3389) );
  XNOR U3562 ( .A(sreg[290]), .B(n3389), .Z(n3391) );
  NANDN U3563 ( .A(sreg[289]), .B(n3312), .Z(n3316) );
  NAND U3564 ( .A(n3314), .B(n3313), .Z(n3315) );
  NAND U3565 ( .A(n3316), .B(n3315), .Z(n3390) );
  XNOR U3566 ( .A(n3391), .B(n3390), .Z(c[290]) );
  NANDN U3567 ( .A(n3318), .B(n3317), .Z(n3322) );
  NANDN U3568 ( .A(n3320), .B(n3319), .Z(n3321) );
  AND U3569 ( .A(n3322), .B(n3321), .Z(n3397) );
  NANDN U3570 ( .A(n3324), .B(n3323), .Z(n3328) );
  NAND U3571 ( .A(n3326), .B(n3325), .Z(n3327) );
  AND U3572 ( .A(n3328), .B(n3327), .Z(n3463) );
  NANDN U3573 ( .A(n3330), .B(n3329), .Z(n3334) );
  NANDN U3574 ( .A(n3332), .B(n3331), .Z(n3333) );
  AND U3575 ( .A(n3334), .B(n3333), .Z(n3429) );
  NAND U3576 ( .A(b[0]), .B(a[51]), .Z(n3335) );
  XNOR U3577 ( .A(b[1]), .B(n3335), .Z(n3337) );
  NANDN U3578 ( .A(b[0]), .B(a[50]), .Z(n3336) );
  NAND U3579 ( .A(n3337), .B(n3336), .Z(n3409) );
  NAND U3580 ( .A(n19808), .B(n3338), .Z(n3340) );
  XOR U3581 ( .A(b[13]), .B(a[39]), .Z(n3412) );
  NAND U3582 ( .A(n19768), .B(n3412), .Z(n3339) );
  AND U3583 ( .A(n3340), .B(n3339), .Z(n3407) );
  AND U3584 ( .A(b[15]), .B(a[35]), .Z(n3406) );
  XNOR U3585 ( .A(n3407), .B(n3406), .Z(n3408) );
  XNOR U3586 ( .A(n3409), .B(n3408), .Z(n3427) );
  NAND U3587 ( .A(n33), .B(n3341), .Z(n3343) );
  XOR U3588 ( .A(b[5]), .B(a[47]), .Z(n3418) );
  NAND U3589 ( .A(n19342), .B(n3418), .Z(n3342) );
  AND U3590 ( .A(n3343), .B(n3342), .Z(n3451) );
  NAND U3591 ( .A(n34), .B(n3344), .Z(n3346) );
  XOR U3592 ( .A(b[7]), .B(a[45]), .Z(n3421) );
  NAND U3593 ( .A(n19486), .B(n3421), .Z(n3345) );
  AND U3594 ( .A(n3346), .B(n3345), .Z(n3449) );
  NAND U3595 ( .A(n31), .B(n3347), .Z(n3349) );
  XOR U3596 ( .A(b[3]), .B(a[49]), .Z(n3424) );
  NAND U3597 ( .A(n32), .B(n3424), .Z(n3348) );
  NAND U3598 ( .A(n3349), .B(n3348), .Z(n3448) );
  XNOR U3599 ( .A(n3449), .B(n3448), .Z(n3450) );
  XOR U3600 ( .A(n3451), .B(n3450), .Z(n3428) );
  XOR U3601 ( .A(n3427), .B(n3428), .Z(n3430) );
  XOR U3602 ( .A(n3429), .B(n3430), .Z(n3401) );
  NANDN U3603 ( .A(n3351), .B(n3350), .Z(n3355) );
  OR U3604 ( .A(n3353), .B(n3352), .Z(n3354) );
  AND U3605 ( .A(n3355), .B(n3354), .Z(n3400) );
  XNOR U3606 ( .A(n3401), .B(n3400), .Z(n3403) );
  NAND U3607 ( .A(n3356), .B(n19724), .Z(n3358) );
  XOR U3608 ( .A(b[11]), .B(a[41]), .Z(n3433) );
  NAND U3609 ( .A(n19692), .B(n3433), .Z(n3357) );
  AND U3610 ( .A(n3358), .B(n3357), .Z(n3444) );
  NAND U3611 ( .A(n19838), .B(n3359), .Z(n3361) );
  XOR U3612 ( .A(b[15]), .B(a[37]), .Z(n3436) );
  NAND U3613 ( .A(n19805), .B(n3436), .Z(n3360) );
  AND U3614 ( .A(n3361), .B(n3360), .Z(n3443) );
  NAND U3615 ( .A(n35), .B(n3362), .Z(n3364) );
  XOR U3616 ( .A(b[9]), .B(a[43]), .Z(n3439) );
  NAND U3617 ( .A(n19598), .B(n3439), .Z(n3363) );
  NAND U3618 ( .A(n3364), .B(n3363), .Z(n3442) );
  XOR U3619 ( .A(n3443), .B(n3442), .Z(n3445) );
  XOR U3620 ( .A(n3444), .B(n3445), .Z(n3455) );
  NANDN U3621 ( .A(n3366), .B(n3365), .Z(n3370) );
  OR U3622 ( .A(n3368), .B(n3367), .Z(n3369) );
  AND U3623 ( .A(n3370), .B(n3369), .Z(n3454) );
  XNOR U3624 ( .A(n3455), .B(n3454), .Z(n3456) );
  NANDN U3625 ( .A(n3372), .B(n3371), .Z(n3376) );
  NANDN U3626 ( .A(n3374), .B(n3373), .Z(n3375) );
  NAND U3627 ( .A(n3376), .B(n3375), .Z(n3457) );
  XNOR U3628 ( .A(n3456), .B(n3457), .Z(n3402) );
  XOR U3629 ( .A(n3403), .B(n3402), .Z(n3461) );
  NANDN U3630 ( .A(n3378), .B(n3377), .Z(n3382) );
  NANDN U3631 ( .A(n3380), .B(n3379), .Z(n3381) );
  AND U3632 ( .A(n3382), .B(n3381), .Z(n3460) );
  XNOR U3633 ( .A(n3461), .B(n3460), .Z(n3462) );
  XOR U3634 ( .A(n3463), .B(n3462), .Z(n3395) );
  NANDN U3635 ( .A(n3384), .B(n3383), .Z(n3388) );
  NAND U3636 ( .A(n3386), .B(n3385), .Z(n3387) );
  AND U3637 ( .A(n3388), .B(n3387), .Z(n3394) );
  XNOR U3638 ( .A(n3395), .B(n3394), .Z(n3396) );
  XNOR U3639 ( .A(n3397), .B(n3396), .Z(n3466) );
  XNOR U3640 ( .A(sreg[291]), .B(n3466), .Z(n3468) );
  NANDN U3641 ( .A(sreg[290]), .B(n3389), .Z(n3393) );
  NAND U3642 ( .A(n3391), .B(n3390), .Z(n3392) );
  NAND U3643 ( .A(n3393), .B(n3392), .Z(n3467) );
  XNOR U3644 ( .A(n3468), .B(n3467), .Z(c[291]) );
  NANDN U3645 ( .A(n3395), .B(n3394), .Z(n3399) );
  NANDN U3646 ( .A(n3397), .B(n3396), .Z(n3398) );
  AND U3647 ( .A(n3399), .B(n3398), .Z(n3474) );
  NANDN U3648 ( .A(n3401), .B(n3400), .Z(n3405) );
  NAND U3649 ( .A(n3403), .B(n3402), .Z(n3404) );
  AND U3650 ( .A(n3405), .B(n3404), .Z(n3540) );
  NANDN U3651 ( .A(n3407), .B(n3406), .Z(n3411) );
  NANDN U3652 ( .A(n3409), .B(n3408), .Z(n3410) );
  AND U3653 ( .A(n3411), .B(n3410), .Z(n3506) );
  NAND U3654 ( .A(n19808), .B(n3412), .Z(n3414) );
  XOR U3655 ( .A(b[13]), .B(a[40]), .Z(n3489) );
  NAND U3656 ( .A(n19768), .B(n3489), .Z(n3413) );
  AND U3657 ( .A(n3414), .B(n3413), .Z(n3484) );
  AND U3658 ( .A(b[15]), .B(a[36]), .Z(n3483) );
  XNOR U3659 ( .A(n3484), .B(n3483), .Z(n3485) );
  NAND U3660 ( .A(b[0]), .B(a[52]), .Z(n3415) );
  XNOR U3661 ( .A(b[1]), .B(n3415), .Z(n3417) );
  NANDN U3662 ( .A(b[0]), .B(a[51]), .Z(n3416) );
  NAND U3663 ( .A(n3417), .B(n3416), .Z(n3486) );
  XNOR U3664 ( .A(n3485), .B(n3486), .Z(n3504) );
  NAND U3665 ( .A(n33), .B(n3418), .Z(n3420) );
  XOR U3666 ( .A(b[5]), .B(a[48]), .Z(n3495) );
  NAND U3667 ( .A(n19342), .B(n3495), .Z(n3419) );
  AND U3668 ( .A(n3420), .B(n3419), .Z(n3528) );
  NAND U3669 ( .A(n34), .B(n3421), .Z(n3423) );
  XOR U3670 ( .A(b[7]), .B(a[46]), .Z(n3498) );
  NAND U3671 ( .A(n19486), .B(n3498), .Z(n3422) );
  AND U3672 ( .A(n3423), .B(n3422), .Z(n3526) );
  NAND U3673 ( .A(n31), .B(n3424), .Z(n3426) );
  XOR U3674 ( .A(b[3]), .B(a[50]), .Z(n3501) );
  NAND U3675 ( .A(n32), .B(n3501), .Z(n3425) );
  NAND U3676 ( .A(n3426), .B(n3425), .Z(n3525) );
  XNOR U3677 ( .A(n3526), .B(n3525), .Z(n3527) );
  XOR U3678 ( .A(n3528), .B(n3527), .Z(n3505) );
  XOR U3679 ( .A(n3504), .B(n3505), .Z(n3507) );
  XOR U3680 ( .A(n3506), .B(n3507), .Z(n3478) );
  NANDN U3681 ( .A(n3428), .B(n3427), .Z(n3432) );
  OR U3682 ( .A(n3430), .B(n3429), .Z(n3431) );
  AND U3683 ( .A(n3432), .B(n3431), .Z(n3477) );
  XNOR U3684 ( .A(n3478), .B(n3477), .Z(n3480) );
  NAND U3685 ( .A(n3433), .B(n19724), .Z(n3435) );
  XOR U3686 ( .A(b[11]), .B(a[42]), .Z(n3510) );
  NAND U3687 ( .A(n19692), .B(n3510), .Z(n3434) );
  AND U3688 ( .A(n3435), .B(n3434), .Z(n3521) );
  NAND U3689 ( .A(n19838), .B(n3436), .Z(n3438) );
  XOR U3690 ( .A(b[15]), .B(a[38]), .Z(n3513) );
  NAND U3691 ( .A(n19805), .B(n3513), .Z(n3437) );
  AND U3692 ( .A(n3438), .B(n3437), .Z(n3520) );
  NAND U3693 ( .A(n35), .B(n3439), .Z(n3441) );
  XOR U3694 ( .A(b[9]), .B(a[44]), .Z(n3516) );
  NAND U3695 ( .A(n19598), .B(n3516), .Z(n3440) );
  NAND U3696 ( .A(n3441), .B(n3440), .Z(n3519) );
  XOR U3697 ( .A(n3520), .B(n3519), .Z(n3522) );
  XOR U3698 ( .A(n3521), .B(n3522), .Z(n3532) );
  NANDN U3699 ( .A(n3443), .B(n3442), .Z(n3447) );
  OR U3700 ( .A(n3445), .B(n3444), .Z(n3446) );
  AND U3701 ( .A(n3447), .B(n3446), .Z(n3531) );
  XNOR U3702 ( .A(n3532), .B(n3531), .Z(n3533) );
  NANDN U3703 ( .A(n3449), .B(n3448), .Z(n3453) );
  NANDN U3704 ( .A(n3451), .B(n3450), .Z(n3452) );
  NAND U3705 ( .A(n3453), .B(n3452), .Z(n3534) );
  XNOR U3706 ( .A(n3533), .B(n3534), .Z(n3479) );
  XOR U3707 ( .A(n3480), .B(n3479), .Z(n3538) );
  NANDN U3708 ( .A(n3455), .B(n3454), .Z(n3459) );
  NANDN U3709 ( .A(n3457), .B(n3456), .Z(n3458) );
  AND U3710 ( .A(n3459), .B(n3458), .Z(n3537) );
  XNOR U3711 ( .A(n3538), .B(n3537), .Z(n3539) );
  XOR U3712 ( .A(n3540), .B(n3539), .Z(n3472) );
  NANDN U3713 ( .A(n3461), .B(n3460), .Z(n3465) );
  NAND U3714 ( .A(n3463), .B(n3462), .Z(n3464) );
  AND U3715 ( .A(n3465), .B(n3464), .Z(n3471) );
  XNOR U3716 ( .A(n3472), .B(n3471), .Z(n3473) );
  XNOR U3717 ( .A(n3474), .B(n3473), .Z(n3543) );
  XNOR U3718 ( .A(sreg[292]), .B(n3543), .Z(n3545) );
  NANDN U3719 ( .A(sreg[291]), .B(n3466), .Z(n3470) );
  NAND U3720 ( .A(n3468), .B(n3467), .Z(n3469) );
  NAND U3721 ( .A(n3470), .B(n3469), .Z(n3544) );
  XNOR U3722 ( .A(n3545), .B(n3544), .Z(c[292]) );
  NANDN U3723 ( .A(n3472), .B(n3471), .Z(n3476) );
  NANDN U3724 ( .A(n3474), .B(n3473), .Z(n3475) );
  AND U3725 ( .A(n3476), .B(n3475), .Z(n3551) );
  NANDN U3726 ( .A(n3478), .B(n3477), .Z(n3482) );
  NAND U3727 ( .A(n3480), .B(n3479), .Z(n3481) );
  AND U3728 ( .A(n3482), .B(n3481), .Z(n3617) );
  NANDN U3729 ( .A(n3484), .B(n3483), .Z(n3488) );
  NANDN U3730 ( .A(n3486), .B(n3485), .Z(n3487) );
  AND U3731 ( .A(n3488), .B(n3487), .Z(n3604) );
  NAND U3732 ( .A(n19808), .B(n3489), .Z(n3491) );
  XOR U3733 ( .A(b[13]), .B(a[41]), .Z(n3590) );
  NAND U3734 ( .A(n19768), .B(n3590), .Z(n3490) );
  AND U3735 ( .A(n3491), .B(n3490), .Z(n3582) );
  AND U3736 ( .A(b[15]), .B(a[37]), .Z(n3581) );
  XNOR U3737 ( .A(n3582), .B(n3581), .Z(n3583) );
  NAND U3738 ( .A(b[0]), .B(a[53]), .Z(n3492) );
  XNOR U3739 ( .A(b[1]), .B(n3492), .Z(n3494) );
  NANDN U3740 ( .A(b[0]), .B(a[52]), .Z(n3493) );
  NAND U3741 ( .A(n3494), .B(n3493), .Z(n3584) );
  XNOR U3742 ( .A(n3583), .B(n3584), .Z(n3602) );
  NAND U3743 ( .A(n33), .B(n3495), .Z(n3497) );
  XOR U3744 ( .A(b[5]), .B(a[49]), .Z(n3593) );
  NAND U3745 ( .A(n19342), .B(n3593), .Z(n3496) );
  AND U3746 ( .A(n3497), .B(n3496), .Z(n3578) );
  NAND U3747 ( .A(n34), .B(n3498), .Z(n3500) );
  XOR U3748 ( .A(b[7]), .B(a[47]), .Z(n3596) );
  NAND U3749 ( .A(n19486), .B(n3596), .Z(n3499) );
  AND U3750 ( .A(n3500), .B(n3499), .Z(n3576) );
  NAND U3751 ( .A(n31), .B(n3501), .Z(n3503) );
  XOR U3752 ( .A(b[3]), .B(a[51]), .Z(n3599) );
  NAND U3753 ( .A(n32), .B(n3599), .Z(n3502) );
  NAND U3754 ( .A(n3503), .B(n3502), .Z(n3575) );
  XNOR U3755 ( .A(n3576), .B(n3575), .Z(n3577) );
  XOR U3756 ( .A(n3578), .B(n3577), .Z(n3603) );
  XOR U3757 ( .A(n3602), .B(n3603), .Z(n3605) );
  XOR U3758 ( .A(n3604), .B(n3605), .Z(n3555) );
  NANDN U3759 ( .A(n3505), .B(n3504), .Z(n3509) );
  OR U3760 ( .A(n3507), .B(n3506), .Z(n3508) );
  AND U3761 ( .A(n3509), .B(n3508), .Z(n3554) );
  XNOR U3762 ( .A(n3555), .B(n3554), .Z(n3557) );
  NAND U3763 ( .A(n3510), .B(n19724), .Z(n3512) );
  XOR U3764 ( .A(b[11]), .B(a[43]), .Z(n3560) );
  NAND U3765 ( .A(n19692), .B(n3560), .Z(n3511) );
  AND U3766 ( .A(n3512), .B(n3511), .Z(n3571) );
  NAND U3767 ( .A(n19838), .B(n3513), .Z(n3515) );
  XOR U3768 ( .A(b[15]), .B(a[39]), .Z(n3563) );
  NAND U3769 ( .A(n19805), .B(n3563), .Z(n3514) );
  AND U3770 ( .A(n3515), .B(n3514), .Z(n3570) );
  NAND U3771 ( .A(n35), .B(n3516), .Z(n3518) );
  XOR U3772 ( .A(b[9]), .B(a[45]), .Z(n3566) );
  NAND U3773 ( .A(n19598), .B(n3566), .Z(n3517) );
  NAND U3774 ( .A(n3518), .B(n3517), .Z(n3569) );
  XOR U3775 ( .A(n3570), .B(n3569), .Z(n3572) );
  XOR U3776 ( .A(n3571), .B(n3572), .Z(n3609) );
  NANDN U3777 ( .A(n3520), .B(n3519), .Z(n3524) );
  OR U3778 ( .A(n3522), .B(n3521), .Z(n3523) );
  AND U3779 ( .A(n3524), .B(n3523), .Z(n3608) );
  XNOR U3780 ( .A(n3609), .B(n3608), .Z(n3610) );
  NANDN U3781 ( .A(n3526), .B(n3525), .Z(n3530) );
  NANDN U3782 ( .A(n3528), .B(n3527), .Z(n3529) );
  NAND U3783 ( .A(n3530), .B(n3529), .Z(n3611) );
  XNOR U3784 ( .A(n3610), .B(n3611), .Z(n3556) );
  XOR U3785 ( .A(n3557), .B(n3556), .Z(n3615) );
  NANDN U3786 ( .A(n3532), .B(n3531), .Z(n3536) );
  NANDN U3787 ( .A(n3534), .B(n3533), .Z(n3535) );
  AND U3788 ( .A(n3536), .B(n3535), .Z(n3614) );
  XNOR U3789 ( .A(n3615), .B(n3614), .Z(n3616) );
  XOR U3790 ( .A(n3617), .B(n3616), .Z(n3549) );
  NANDN U3791 ( .A(n3538), .B(n3537), .Z(n3542) );
  NAND U3792 ( .A(n3540), .B(n3539), .Z(n3541) );
  AND U3793 ( .A(n3542), .B(n3541), .Z(n3548) );
  XNOR U3794 ( .A(n3549), .B(n3548), .Z(n3550) );
  XNOR U3795 ( .A(n3551), .B(n3550), .Z(n3620) );
  XNOR U3796 ( .A(sreg[293]), .B(n3620), .Z(n3622) );
  NANDN U3797 ( .A(sreg[292]), .B(n3543), .Z(n3547) );
  NAND U3798 ( .A(n3545), .B(n3544), .Z(n3546) );
  NAND U3799 ( .A(n3547), .B(n3546), .Z(n3621) );
  XNOR U3800 ( .A(n3622), .B(n3621), .Z(c[293]) );
  NANDN U3801 ( .A(n3549), .B(n3548), .Z(n3553) );
  NANDN U3802 ( .A(n3551), .B(n3550), .Z(n3552) );
  AND U3803 ( .A(n3553), .B(n3552), .Z(n3628) );
  NANDN U3804 ( .A(n3555), .B(n3554), .Z(n3559) );
  NAND U3805 ( .A(n3557), .B(n3556), .Z(n3558) );
  AND U3806 ( .A(n3559), .B(n3558), .Z(n3694) );
  NAND U3807 ( .A(n3560), .B(n19724), .Z(n3562) );
  XOR U3808 ( .A(b[11]), .B(a[44]), .Z(n3664) );
  NAND U3809 ( .A(n19692), .B(n3664), .Z(n3561) );
  AND U3810 ( .A(n3562), .B(n3561), .Z(n3675) );
  NAND U3811 ( .A(n19838), .B(n3563), .Z(n3565) );
  XOR U3812 ( .A(b[15]), .B(a[40]), .Z(n3667) );
  NAND U3813 ( .A(n19805), .B(n3667), .Z(n3564) );
  AND U3814 ( .A(n3565), .B(n3564), .Z(n3674) );
  NAND U3815 ( .A(n35), .B(n3566), .Z(n3568) );
  XOR U3816 ( .A(b[9]), .B(a[46]), .Z(n3670) );
  NAND U3817 ( .A(n19598), .B(n3670), .Z(n3567) );
  NAND U3818 ( .A(n3568), .B(n3567), .Z(n3673) );
  XOR U3819 ( .A(n3674), .B(n3673), .Z(n3676) );
  XOR U3820 ( .A(n3675), .B(n3676), .Z(n3686) );
  NANDN U3821 ( .A(n3570), .B(n3569), .Z(n3574) );
  OR U3822 ( .A(n3572), .B(n3571), .Z(n3573) );
  AND U3823 ( .A(n3574), .B(n3573), .Z(n3685) );
  XNOR U3824 ( .A(n3686), .B(n3685), .Z(n3687) );
  NANDN U3825 ( .A(n3576), .B(n3575), .Z(n3580) );
  NANDN U3826 ( .A(n3578), .B(n3577), .Z(n3579) );
  NAND U3827 ( .A(n3580), .B(n3579), .Z(n3688) );
  XNOR U3828 ( .A(n3687), .B(n3688), .Z(n3634) );
  NANDN U3829 ( .A(n3582), .B(n3581), .Z(n3586) );
  NANDN U3830 ( .A(n3584), .B(n3583), .Z(n3585) );
  AND U3831 ( .A(n3586), .B(n3585), .Z(n3660) );
  NAND U3832 ( .A(b[0]), .B(a[54]), .Z(n3587) );
  XNOR U3833 ( .A(b[1]), .B(n3587), .Z(n3589) );
  NANDN U3834 ( .A(b[0]), .B(a[53]), .Z(n3588) );
  NAND U3835 ( .A(n3589), .B(n3588), .Z(n3640) );
  NAND U3836 ( .A(n19808), .B(n3590), .Z(n3592) );
  XOR U3837 ( .A(b[13]), .B(a[42]), .Z(n3646) );
  NAND U3838 ( .A(n19768), .B(n3646), .Z(n3591) );
  AND U3839 ( .A(n3592), .B(n3591), .Z(n3638) );
  AND U3840 ( .A(b[15]), .B(a[38]), .Z(n3637) );
  XNOR U3841 ( .A(n3638), .B(n3637), .Z(n3639) );
  XNOR U3842 ( .A(n3640), .B(n3639), .Z(n3658) );
  NAND U3843 ( .A(n33), .B(n3593), .Z(n3595) );
  XOR U3844 ( .A(b[5]), .B(a[50]), .Z(n3649) );
  NAND U3845 ( .A(n19342), .B(n3649), .Z(n3594) );
  AND U3846 ( .A(n3595), .B(n3594), .Z(n3682) );
  NAND U3847 ( .A(n34), .B(n3596), .Z(n3598) );
  XOR U3848 ( .A(b[7]), .B(a[48]), .Z(n3652) );
  NAND U3849 ( .A(n19486), .B(n3652), .Z(n3597) );
  AND U3850 ( .A(n3598), .B(n3597), .Z(n3680) );
  NAND U3851 ( .A(n31), .B(n3599), .Z(n3601) );
  XOR U3852 ( .A(b[3]), .B(a[52]), .Z(n3655) );
  NAND U3853 ( .A(n32), .B(n3655), .Z(n3600) );
  NAND U3854 ( .A(n3601), .B(n3600), .Z(n3679) );
  XNOR U3855 ( .A(n3680), .B(n3679), .Z(n3681) );
  XOR U3856 ( .A(n3682), .B(n3681), .Z(n3659) );
  XOR U3857 ( .A(n3658), .B(n3659), .Z(n3661) );
  XOR U3858 ( .A(n3660), .B(n3661), .Z(n3632) );
  NANDN U3859 ( .A(n3603), .B(n3602), .Z(n3607) );
  OR U3860 ( .A(n3605), .B(n3604), .Z(n3606) );
  AND U3861 ( .A(n3607), .B(n3606), .Z(n3631) );
  XNOR U3862 ( .A(n3632), .B(n3631), .Z(n3633) );
  XOR U3863 ( .A(n3634), .B(n3633), .Z(n3692) );
  NANDN U3864 ( .A(n3609), .B(n3608), .Z(n3613) );
  NANDN U3865 ( .A(n3611), .B(n3610), .Z(n3612) );
  AND U3866 ( .A(n3613), .B(n3612), .Z(n3691) );
  XNOR U3867 ( .A(n3692), .B(n3691), .Z(n3693) );
  XOR U3868 ( .A(n3694), .B(n3693), .Z(n3626) );
  NANDN U3869 ( .A(n3615), .B(n3614), .Z(n3619) );
  NAND U3870 ( .A(n3617), .B(n3616), .Z(n3618) );
  AND U3871 ( .A(n3619), .B(n3618), .Z(n3625) );
  XNOR U3872 ( .A(n3626), .B(n3625), .Z(n3627) );
  XNOR U3873 ( .A(n3628), .B(n3627), .Z(n3697) );
  XNOR U3874 ( .A(sreg[294]), .B(n3697), .Z(n3699) );
  NANDN U3875 ( .A(sreg[293]), .B(n3620), .Z(n3624) );
  NAND U3876 ( .A(n3622), .B(n3621), .Z(n3623) );
  NAND U3877 ( .A(n3624), .B(n3623), .Z(n3698) );
  XNOR U3878 ( .A(n3699), .B(n3698), .Z(c[294]) );
  NANDN U3879 ( .A(n3626), .B(n3625), .Z(n3630) );
  NANDN U3880 ( .A(n3628), .B(n3627), .Z(n3629) );
  AND U3881 ( .A(n3630), .B(n3629), .Z(n3705) );
  NANDN U3882 ( .A(n3632), .B(n3631), .Z(n3636) );
  NAND U3883 ( .A(n3634), .B(n3633), .Z(n3635) );
  AND U3884 ( .A(n3636), .B(n3635), .Z(n3771) );
  NANDN U3885 ( .A(n3638), .B(n3637), .Z(n3642) );
  NANDN U3886 ( .A(n3640), .B(n3639), .Z(n3641) );
  AND U3887 ( .A(n3642), .B(n3641), .Z(n3758) );
  NAND U3888 ( .A(b[0]), .B(a[55]), .Z(n3643) );
  XNOR U3889 ( .A(b[1]), .B(n3643), .Z(n3645) );
  NANDN U3890 ( .A(b[0]), .B(a[54]), .Z(n3644) );
  NAND U3891 ( .A(n3645), .B(n3644), .Z(n3738) );
  NAND U3892 ( .A(n19808), .B(n3646), .Z(n3648) );
  XOR U3893 ( .A(b[13]), .B(a[43]), .Z(n3744) );
  NAND U3894 ( .A(n19768), .B(n3744), .Z(n3647) );
  AND U3895 ( .A(n3648), .B(n3647), .Z(n3736) );
  AND U3896 ( .A(b[15]), .B(a[39]), .Z(n3735) );
  XNOR U3897 ( .A(n3736), .B(n3735), .Z(n3737) );
  XNOR U3898 ( .A(n3738), .B(n3737), .Z(n3756) );
  NAND U3899 ( .A(n33), .B(n3649), .Z(n3651) );
  XOR U3900 ( .A(b[5]), .B(a[51]), .Z(n3747) );
  NAND U3901 ( .A(n19342), .B(n3747), .Z(n3650) );
  AND U3902 ( .A(n3651), .B(n3650), .Z(n3732) );
  NAND U3903 ( .A(n34), .B(n3652), .Z(n3654) );
  XOR U3904 ( .A(b[7]), .B(a[49]), .Z(n3750) );
  NAND U3905 ( .A(n19486), .B(n3750), .Z(n3653) );
  AND U3906 ( .A(n3654), .B(n3653), .Z(n3730) );
  NAND U3907 ( .A(n31), .B(n3655), .Z(n3657) );
  XOR U3908 ( .A(b[3]), .B(a[53]), .Z(n3753) );
  NAND U3909 ( .A(n32), .B(n3753), .Z(n3656) );
  NAND U3910 ( .A(n3657), .B(n3656), .Z(n3729) );
  XNOR U3911 ( .A(n3730), .B(n3729), .Z(n3731) );
  XOR U3912 ( .A(n3732), .B(n3731), .Z(n3757) );
  XOR U3913 ( .A(n3756), .B(n3757), .Z(n3759) );
  XOR U3914 ( .A(n3758), .B(n3759), .Z(n3709) );
  NANDN U3915 ( .A(n3659), .B(n3658), .Z(n3663) );
  OR U3916 ( .A(n3661), .B(n3660), .Z(n3662) );
  AND U3917 ( .A(n3663), .B(n3662), .Z(n3708) );
  XNOR U3918 ( .A(n3709), .B(n3708), .Z(n3711) );
  NAND U3919 ( .A(n3664), .B(n19724), .Z(n3666) );
  XOR U3920 ( .A(b[11]), .B(a[45]), .Z(n3714) );
  NAND U3921 ( .A(n19692), .B(n3714), .Z(n3665) );
  AND U3922 ( .A(n3666), .B(n3665), .Z(n3725) );
  NAND U3923 ( .A(n19838), .B(n3667), .Z(n3669) );
  XOR U3924 ( .A(b[15]), .B(a[41]), .Z(n3717) );
  NAND U3925 ( .A(n19805), .B(n3717), .Z(n3668) );
  AND U3926 ( .A(n3669), .B(n3668), .Z(n3724) );
  NAND U3927 ( .A(n35), .B(n3670), .Z(n3672) );
  XOR U3928 ( .A(b[9]), .B(a[47]), .Z(n3720) );
  NAND U3929 ( .A(n19598), .B(n3720), .Z(n3671) );
  NAND U3930 ( .A(n3672), .B(n3671), .Z(n3723) );
  XOR U3931 ( .A(n3724), .B(n3723), .Z(n3726) );
  XOR U3932 ( .A(n3725), .B(n3726), .Z(n3763) );
  NANDN U3933 ( .A(n3674), .B(n3673), .Z(n3678) );
  OR U3934 ( .A(n3676), .B(n3675), .Z(n3677) );
  AND U3935 ( .A(n3678), .B(n3677), .Z(n3762) );
  XNOR U3936 ( .A(n3763), .B(n3762), .Z(n3764) );
  NANDN U3937 ( .A(n3680), .B(n3679), .Z(n3684) );
  NANDN U3938 ( .A(n3682), .B(n3681), .Z(n3683) );
  NAND U3939 ( .A(n3684), .B(n3683), .Z(n3765) );
  XNOR U3940 ( .A(n3764), .B(n3765), .Z(n3710) );
  XOR U3941 ( .A(n3711), .B(n3710), .Z(n3769) );
  NANDN U3942 ( .A(n3686), .B(n3685), .Z(n3690) );
  NANDN U3943 ( .A(n3688), .B(n3687), .Z(n3689) );
  AND U3944 ( .A(n3690), .B(n3689), .Z(n3768) );
  XNOR U3945 ( .A(n3769), .B(n3768), .Z(n3770) );
  XOR U3946 ( .A(n3771), .B(n3770), .Z(n3703) );
  NANDN U3947 ( .A(n3692), .B(n3691), .Z(n3696) );
  NAND U3948 ( .A(n3694), .B(n3693), .Z(n3695) );
  AND U3949 ( .A(n3696), .B(n3695), .Z(n3702) );
  XNOR U3950 ( .A(n3703), .B(n3702), .Z(n3704) );
  XNOR U3951 ( .A(n3705), .B(n3704), .Z(n3774) );
  XNOR U3952 ( .A(sreg[295]), .B(n3774), .Z(n3776) );
  NANDN U3953 ( .A(sreg[294]), .B(n3697), .Z(n3701) );
  NAND U3954 ( .A(n3699), .B(n3698), .Z(n3700) );
  NAND U3955 ( .A(n3701), .B(n3700), .Z(n3775) );
  XNOR U3956 ( .A(n3776), .B(n3775), .Z(c[295]) );
  NANDN U3957 ( .A(n3703), .B(n3702), .Z(n3707) );
  NANDN U3958 ( .A(n3705), .B(n3704), .Z(n3706) );
  AND U3959 ( .A(n3707), .B(n3706), .Z(n3782) );
  NANDN U3960 ( .A(n3709), .B(n3708), .Z(n3713) );
  NAND U3961 ( .A(n3711), .B(n3710), .Z(n3712) );
  AND U3962 ( .A(n3713), .B(n3712), .Z(n3848) );
  NAND U3963 ( .A(n3714), .B(n19724), .Z(n3716) );
  XOR U3964 ( .A(b[11]), .B(a[46]), .Z(n3818) );
  NAND U3965 ( .A(n19692), .B(n3818), .Z(n3715) );
  AND U3966 ( .A(n3716), .B(n3715), .Z(n3829) );
  NAND U3967 ( .A(n19838), .B(n3717), .Z(n3719) );
  XOR U3968 ( .A(b[15]), .B(a[42]), .Z(n3821) );
  NAND U3969 ( .A(n19805), .B(n3821), .Z(n3718) );
  AND U3970 ( .A(n3719), .B(n3718), .Z(n3828) );
  NAND U3971 ( .A(n35), .B(n3720), .Z(n3722) );
  XOR U3972 ( .A(b[9]), .B(a[48]), .Z(n3824) );
  NAND U3973 ( .A(n19598), .B(n3824), .Z(n3721) );
  NAND U3974 ( .A(n3722), .B(n3721), .Z(n3827) );
  XOR U3975 ( .A(n3828), .B(n3827), .Z(n3830) );
  XOR U3976 ( .A(n3829), .B(n3830), .Z(n3840) );
  NANDN U3977 ( .A(n3724), .B(n3723), .Z(n3728) );
  OR U3978 ( .A(n3726), .B(n3725), .Z(n3727) );
  AND U3979 ( .A(n3728), .B(n3727), .Z(n3839) );
  XNOR U3980 ( .A(n3840), .B(n3839), .Z(n3841) );
  NANDN U3981 ( .A(n3730), .B(n3729), .Z(n3734) );
  NANDN U3982 ( .A(n3732), .B(n3731), .Z(n3733) );
  NAND U3983 ( .A(n3734), .B(n3733), .Z(n3842) );
  XNOR U3984 ( .A(n3841), .B(n3842), .Z(n3788) );
  NANDN U3985 ( .A(n3736), .B(n3735), .Z(n3740) );
  NANDN U3986 ( .A(n3738), .B(n3737), .Z(n3739) );
  AND U3987 ( .A(n3740), .B(n3739), .Z(n3814) );
  NAND U3988 ( .A(b[0]), .B(a[56]), .Z(n3741) );
  XNOR U3989 ( .A(b[1]), .B(n3741), .Z(n3743) );
  NANDN U3990 ( .A(b[0]), .B(a[55]), .Z(n3742) );
  NAND U3991 ( .A(n3743), .B(n3742), .Z(n3794) );
  NAND U3992 ( .A(n19808), .B(n3744), .Z(n3746) );
  XOR U3993 ( .A(b[13]), .B(a[44]), .Z(n3800) );
  NAND U3994 ( .A(n19768), .B(n3800), .Z(n3745) );
  AND U3995 ( .A(n3746), .B(n3745), .Z(n3792) );
  AND U3996 ( .A(b[15]), .B(a[40]), .Z(n3791) );
  XNOR U3997 ( .A(n3792), .B(n3791), .Z(n3793) );
  XNOR U3998 ( .A(n3794), .B(n3793), .Z(n3812) );
  NAND U3999 ( .A(n33), .B(n3747), .Z(n3749) );
  XOR U4000 ( .A(b[5]), .B(a[52]), .Z(n3803) );
  NAND U4001 ( .A(n19342), .B(n3803), .Z(n3748) );
  AND U4002 ( .A(n3749), .B(n3748), .Z(n3836) );
  NAND U4003 ( .A(n34), .B(n3750), .Z(n3752) );
  XOR U4004 ( .A(b[7]), .B(a[50]), .Z(n3806) );
  NAND U4005 ( .A(n19486), .B(n3806), .Z(n3751) );
  AND U4006 ( .A(n3752), .B(n3751), .Z(n3834) );
  NAND U4007 ( .A(n31), .B(n3753), .Z(n3755) );
  XOR U4008 ( .A(b[3]), .B(a[54]), .Z(n3809) );
  NAND U4009 ( .A(n32), .B(n3809), .Z(n3754) );
  NAND U4010 ( .A(n3755), .B(n3754), .Z(n3833) );
  XNOR U4011 ( .A(n3834), .B(n3833), .Z(n3835) );
  XOR U4012 ( .A(n3836), .B(n3835), .Z(n3813) );
  XOR U4013 ( .A(n3812), .B(n3813), .Z(n3815) );
  XOR U4014 ( .A(n3814), .B(n3815), .Z(n3786) );
  NANDN U4015 ( .A(n3757), .B(n3756), .Z(n3761) );
  OR U4016 ( .A(n3759), .B(n3758), .Z(n3760) );
  AND U4017 ( .A(n3761), .B(n3760), .Z(n3785) );
  XNOR U4018 ( .A(n3786), .B(n3785), .Z(n3787) );
  XOR U4019 ( .A(n3788), .B(n3787), .Z(n3846) );
  NANDN U4020 ( .A(n3763), .B(n3762), .Z(n3767) );
  NANDN U4021 ( .A(n3765), .B(n3764), .Z(n3766) );
  AND U4022 ( .A(n3767), .B(n3766), .Z(n3845) );
  XNOR U4023 ( .A(n3846), .B(n3845), .Z(n3847) );
  XOR U4024 ( .A(n3848), .B(n3847), .Z(n3780) );
  NANDN U4025 ( .A(n3769), .B(n3768), .Z(n3773) );
  NAND U4026 ( .A(n3771), .B(n3770), .Z(n3772) );
  AND U4027 ( .A(n3773), .B(n3772), .Z(n3779) );
  XNOR U4028 ( .A(n3780), .B(n3779), .Z(n3781) );
  XNOR U4029 ( .A(n3782), .B(n3781), .Z(n3851) );
  XNOR U4030 ( .A(sreg[296]), .B(n3851), .Z(n3853) );
  NANDN U4031 ( .A(sreg[295]), .B(n3774), .Z(n3778) );
  NAND U4032 ( .A(n3776), .B(n3775), .Z(n3777) );
  NAND U4033 ( .A(n3778), .B(n3777), .Z(n3852) );
  XNOR U4034 ( .A(n3853), .B(n3852), .Z(c[296]) );
  NANDN U4035 ( .A(n3780), .B(n3779), .Z(n3784) );
  NANDN U4036 ( .A(n3782), .B(n3781), .Z(n3783) );
  AND U4037 ( .A(n3784), .B(n3783), .Z(n3859) );
  NANDN U4038 ( .A(n3786), .B(n3785), .Z(n3790) );
  NAND U4039 ( .A(n3788), .B(n3787), .Z(n3789) );
  AND U4040 ( .A(n3790), .B(n3789), .Z(n3925) );
  NANDN U4041 ( .A(n3792), .B(n3791), .Z(n3796) );
  NANDN U4042 ( .A(n3794), .B(n3793), .Z(n3795) );
  AND U4043 ( .A(n3796), .B(n3795), .Z(n3891) );
  NAND U4044 ( .A(b[0]), .B(a[57]), .Z(n3797) );
  XNOR U4045 ( .A(b[1]), .B(n3797), .Z(n3799) );
  NANDN U4046 ( .A(b[0]), .B(a[56]), .Z(n3798) );
  NAND U4047 ( .A(n3799), .B(n3798), .Z(n3871) );
  NAND U4048 ( .A(n19808), .B(n3800), .Z(n3802) );
  XOR U4049 ( .A(b[13]), .B(a[45]), .Z(n3877) );
  NAND U4050 ( .A(n19768), .B(n3877), .Z(n3801) );
  AND U4051 ( .A(n3802), .B(n3801), .Z(n3869) );
  AND U4052 ( .A(b[15]), .B(a[41]), .Z(n3868) );
  XNOR U4053 ( .A(n3869), .B(n3868), .Z(n3870) );
  XNOR U4054 ( .A(n3871), .B(n3870), .Z(n3889) );
  NAND U4055 ( .A(n33), .B(n3803), .Z(n3805) );
  XOR U4056 ( .A(b[5]), .B(a[53]), .Z(n3880) );
  NAND U4057 ( .A(n19342), .B(n3880), .Z(n3804) );
  AND U4058 ( .A(n3805), .B(n3804), .Z(n3913) );
  NAND U4059 ( .A(n34), .B(n3806), .Z(n3808) );
  XOR U4060 ( .A(b[7]), .B(a[51]), .Z(n3883) );
  NAND U4061 ( .A(n19486), .B(n3883), .Z(n3807) );
  AND U4062 ( .A(n3808), .B(n3807), .Z(n3911) );
  NAND U4063 ( .A(n31), .B(n3809), .Z(n3811) );
  XOR U4064 ( .A(b[3]), .B(a[55]), .Z(n3886) );
  NAND U4065 ( .A(n32), .B(n3886), .Z(n3810) );
  NAND U4066 ( .A(n3811), .B(n3810), .Z(n3910) );
  XNOR U4067 ( .A(n3911), .B(n3910), .Z(n3912) );
  XOR U4068 ( .A(n3913), .B(n3912), .Z(n3890) );
  XOR U4069 ( .A(n3889), .B(n3890), .Z(n3892) );
  XOR U4070 ( .A(n3891), .B(n3892), .Z(n3863) );
  NANDN U4071 ( .A(n3813), .B(n3812), .Z(n3817) );
  OR U4072 ( .A(n3815), .B(n3814), .Z(n3816) );
  AND U4073 ( .A(n3817), .B(n3816), .Z(n3862) );
  XNOR U4074 ( .A(n3863), .B(n3862), .Z(n3865) );
  NAND U4075 ( .A(n3818), .B(n19724), .Z(n3820) );
  XOR U4076 ( .A(b[11]), .B(a[47]), .Z(n3895) );
  NAND U4077 ( .A(n19692), .B(n3895), .Z(n3819) );
  AND U4078 ( .A(n3820), .B(n3819), .Z(n3906) );
  NAND U4079 ( .A(n19838), .B(n3821), .Z(n3823) );
  XOR U4080 ( .A(b[15]), .B(a[43]), .Z(n3898) );
  NAND U4081 ( .A(n19805), .B(n3898), .Z(n3822) );
  AND U4082 ( .A(n3823), .B(n3822), .Z(n3905) );
  NAND U4083 ( .A(n35), .B(n3824), .Z(n3826) );
  XOR U4084 ( .A(b[9]), .B(a[49]), .Z(n3901) );
  NAND U4085 ( .A(n19598), .B(n3901), .Z(n3825) );
  NAND U4086 ( .A(n3826), .B(n3825), .Z(n3904) );
  XOR U4087 ( .A(n3905), .B(n3904), .Z(n3907) );
  XOR U4088 ( .A(n3906), .B(n3907), .Z(n3917) );
  NANDN U4089 ( .A(n3828), .B(n3827), .Z(n3832) );
  OR U4090 ( .A(n3830), .B(n3829), .Z(n3831) );
  AND U4091 ( .A(n3832), .B(n3831), .Z(n3916) );
  XNOR U4092 ( .A(n3917), .B(n3916), .Z(n3918) );
  NANDN U4093 ( .A(n3834), .B(n3833), .Z(n3838) );
  NANDN U4094 ( .A(n3836), .B(n3835), .Z(n3837) );
  NAND U4095 ( .A(n3838), .B(n3837), .Z(n3919) );
  XNOR U4096 ( .A(n3918), .B(n3919), .Z(n3864) );
  XOR U4097 ( .A(n3865), .B(n3864), .Z(n3923) );
  NANDN U4098 ( .A(n3840), .B(n3839), .Z(n3844) );
  NANDN U4099 ( .A(n3842), .B(n3841), .Z(n3843) );
  AND U4100 ( .A(n3844), .B(n3843), .Z(n3922) );
  XNOR U4101 ( .A(n3923), .B(n3922), .Z(n3924) );
  XOR U4102 ( .A(n3925), .B(n3924), .Z(n3857) );
  NANDN U4103 ( .A(n3846), .B(n3845), .Z(n3850) );
  NAND U4104 ( .A(n3848), .B(n3847), .Z(n3849) );
  AND U4105 ( .A(n3850), .B(n3849), .Z(n3856) );
  XNOR U4106 ( .A(n3857), .B(n3856), .Z(n3858) );
  XNOR U4107 ( .A(n3859), .B(n3858), .Z(n3928) );
  XNOR U4108 ( .A(sreg[297]), .B(n3928), .Z(n3930) );
  NANDN U4109 ( .A(sreg[296]), .B(n3851), .Z(n3855) );
  NAND U4110 ( .A(n3853), .B(n3852), .Z(n3854) );
  NAND U4111 ( .A(n3855), .B(n3854), .Z(n3929) );
  XNOR U4112 ( .A(n3930), .B(n3929), .Z(c[297]) );
  NANDN U4113 ( .A(n3857), .B(n3856), .Z(n3861) );
  NANDN U4114 ( .A(n3859), .B(n3858), .Z(n3860) );
  AND U4115 ( .A(n3861), .B(n3860), .Z(n3936) );
  NANDN U4116 ( .A(n3863), .B(n3862), .Z(n3867) );
  NAND U4117 ( .A(n3865), .B(n3864), .Z(n3866) );
  AND U4118 ( .A(n3867), .B(n3866), .Z(n4002) );
  NANDN U4119 ( .A(n3869), .B(n3868), .Z(n3873) );
  NANDN U4120 ( .A(n3871), .B(n3870), .Z(n3872) );
  AND U4121 ( .A(n3873), .B(n3872), .Z(n3968) );
  NAND U4122 ( .A(b[0]), .B(a[58]), .Z(n3874) );
  XNOR U4123 ( .A(b[1]), .B(n3874), .Z(n3876) );
  NANDN U4124 ( .A(b[0]), .B(a[57]), .Z(n3875) );
  NAND U4125 ( .A(n3876), .B(n3875), .Z(n3948) );
  NAND U4126 ( .A(n19808), .B(n3877), .Z(n3879) );
  XOR U4127 ( .A(b[13]), .B(a[46]), .Z(n3951) );
  NAND U4128 ( .A(n19768), .B(n3951), .Z(n3878) );
  AND U4129 ( .A(n3879), .B(n3878), .Z(n3946) );
  AND U4130 ( .A(b[15]), .B(a[42]), .Z(n3945) );
  XNOR U4131 ( .A(n3946), .B(n3945), .Z(n3947) );
  XNOR U4132 ( .A(n3948), .B(n3947), .Z(n3966) );
  NAND U4133 ( .A(n33), .B(n3880), .Z(n3882) );
  XOR U4134 ( .A(b[5]), .B(a[54]), .Z(n3957) );
  NAND U4135 ( .A(n19342), .B(n3957), .Z(n3881) );
  AND U4136 ( .A(n3882), .B(n3881), .Z(n3990) );
  NAND U4137 ( .A(n34), .B(n3883), .Z(n3885) );
  XOR U4138 ( .A(b[7]), .B(a[52]), .Z(n3960) );
  NAND U4139 ( .A(n19486), .B(n3960), .Z(n3884) );
  AND U4140 ( .A(n3885), .B(n3884), .Z(n3988) );
  NAND U4141 ( .A(n31), .B(n3886), .Z(n3888) );
  XOR U4142 ( .A(b[3]), .B(a[56]), .Z(n3963) );
  NAND U4143 ( .A(n32), .B(n3963), .Z(n3887) );
  NAND U4144 ( .A(n3888), .B(n3887), .Z(n3987) );
  XNOR U4145 ( .A(n3988), .B(n3987), .Z(n3989) );
  XOR U4146 ( .A(n3990), .B(n3989), .Z(n3967) );
  XOR U4147 ( .A(n3966), .B(n3967), .Z(n3969) );
  XOR U4148 ( .A(n3968), .B(n3969), .Z(n3940) );
  NANDN U4149 ( .A(n3890), .B(n3889), .Z(n3894) );
  OR U4150 ( .A(n3892), .B(n3891), .Z(n3893) );
  AND U4151 ( .A(n3894), .B(n3893), .Z(n3939) );
  XNOR U4152 ( .A(n3940), .B(n3939), .Z(n3942) );
  NAND U4153 ( .A(n3895), .B(n19724), .Z(n3897) );
  XOR U4154 ( .A(b[11]), .B(a[48]), .Z(n3972) );
  NAND U4155 ( .A(n19692), .B(n3972), .Z(n3896) );
  AND U4156 ( .A(n3897), .B(n3896), .Z(n3983) );
  NAND U4157 ( .A(n19838), .B(n3898), .Z(n3900) );
  XOR U4158 ( .A(b[15]), .B(a[44]), .Z(n3975) );
  NAND U4159 ( .A(n19805), .B(n3975), .Z(n3899) );
  AND U4160 ( .A(n3900), .B(n3899), .Z(n3982) );
  NAND U4161 ( .A(n35), .B(n3901), .Z(n3903) );
  XOR U4162 ( .A(b[9]), .B(a[50]), .Z(n3978) );
  NAND U4163 ( .A(n19598), .B(n3978), .Z(n3902) );
  NAND U4164 ( .A(n3903), .B(n3902), .Z(n3981) );
  XOR U4165 ( .A(n3982), .B(n3981), .Z(n3984) );
  XOR U4166 ( .A(n3983), .B(n3984), .Z(n3994) );
  NANDN U4167 ( .A(n3905), .B(n3904), .Z(n3909) );
  OR U4168 ( .A(n3907), .B(n3906), .Z(n3908) );
  AND U4169 ( .A(n3909), .B(n3908), .Z(n3993) );
  XNOR U4170 ( .A(n3994), .B(n3993), .Z(n3995) );
  NANDN U4171 ( .A(n3911), .B(n3910), .Z(n3915) );
  NANDN U4172 ( .A(n3913), .B(n3912), .Z(n3914) );
  NAND U4173 ( .A(n3915), .B(n3914), .Z(n3996) );
  XNOR U4174 ( .A(n3995), .B(n3996), .Z(n3941) );
  XOR U4175 ( .A(n3942), .B(n3941), .Z(n4000) );
  NANDN U4176 ( .A(n3917), .B(n3916), .Z(n3921) );
  NANDN U4177 ( .A(n3919), .B(n3918), .Z(n3920) );
  AND U4178 ( .A(n3921), .B(n3920), .Z(n3999) );
  XNOR U4179 ( .A(n4000), .B(n3999), .Z(n4001) );
  XOR U4180 ( .A(n4002), .B(n4001), .Z(n3934) );
  NANDN U4181 ( .A(n3923), .B(n3922), .Z(n3927) );
  NAND U4182 ( .A(n3925), .B(n3924), .Z(n3926) );
  AND U4183 ( .A(n3927), .B(n3926), .Z(n3933) );
  XNOR U4184 ( .A(n3934), .B(n3933), .Z(n3935) );
  XNOR U4185 ( .A(n3936), .B(n3935), .Z(n4005) );
  XNOR U4186 ( .A(sreg[298]), .B(n4005), .Z(n4007) );
  NANDN U4187 ( .A(sreg[297]), .B(n3928), .Z(n3932) );
  NAND U4188 ( .A(n3930), .B(n3929), .Z(n3931) );
  NAND U4189 ( .A(n3932), .B(n3931), .Z(n4006) );
  XNOR U4190 ( .A(n4007), .B(n4006), .Z(c[298]) );
  NANDN U4191 ( .A(n3934), .B(n3933), .Z(n3938) );
  NANDN U4192 ( .A(n3936), .B(n3935), .Z(n3937) );
  AND U4193 ( .A(n3938), .B(n3937), .Z(n4013) );
  NANDN U4194 ( .A(n3940), .B(n3939), .Z(n3944) );
  NAND U4195 ( .A(n3942), .B(n3941), .Z(n3943) );
  AND U4196 ( .A(n3944), .B(n3943), .Z(n4079) );
  NANDN U4197 ( .A(n3946), .B(n3945), .Z(n3950) );
  NANDN U4198 ( .A(n3948), .B(n3947), .Z(n3949) );
  AND U4199 ( .A(n3950), .B(n3949), .Z(n4045) );
  NAND U4200 ( .A(n19808), .B(n3951), .Z(n3953) );
  XOR U4201 ( .A(b[13]), .B(a[47]), .Z(n4031) );
  NAND U4202 ( .A(n19768), .B(n4031), .Z(n3952) );
  AND U4203 ( .A(n3953), .B(n3952), .Z(n4023) );
  AND U4204 ( .A(b[15]), .B(a[43]), .Z(n4022) );
  XNOR U4205 ( .A(n4023), .B(n4022), .Z(n4024) );
  NAND U4206 ( .A(b[0]), .B(a[59]), .Z(n3954) );
  XNOR U4207 ( .A(b[1]), .B(n3954), .Z(n3956) );
  NANDN U4208 ( .A(b[0]), .B(a[58]), .Z(n3955) );
  NAND U4209 ( .A(n3956), .B(n3955), .Z(n4025) );
  XNOR U4210 ( .A(n4024), .B(n4025), .Z(n4043) );
  NAND U4211 ( .A(n33), .B(n3957), .Z(n3959) );
  XOR U4212 ( .A(b[5]), .B(a[55]), .Z(n4034) );
  NAND U4213 ( .A(n19342), .B(n4034), .Z(n3958) );
  AND U4214 ( .A(n3959), .B(n3958), .Z(n4067) );
  NAND U4215 ( .A(n34), .B(n3960), .Z(n3962) );
  XOR U4216 ( .A(b[7]), .B(a[53]), .Z(n4037) );
  NAND U4217 ( .A(n19486), .B(n4037), .Z(n3961) );
  AND U4218 ( .A(n3962), .B(n3961), .Z(n4065) );
  NAND U4219 ( .A(n31), .B(n3963), .Z(n3965) );
  XOR U4220 ( .A(b[3]), .B(a[57]), .Z(n4040) );
  NAND U4221 ( .A(n32), .B(n4040), .Z(n3964) );
  NAND U4222 ( .A(n3965), .B(n3964), .Z(n4064) );
  XNOR U4223 ( .A(n4065), .B(n4064), .Z(n4066) );
  XOR U4224 ( .A(n4067), .B(n4066), .Z(n4044) );
  XOR U4225 ( .A(n4043), .B(n4044), .Z(n4046) );
  XOR U4226 ( .A(n4045), .B(n4046), .Z(n4017) );
  NANDN U4227 ( .A(n3967), .B(n3966), .Z(n3971) );
  OR U4228 ( .A(n3969), .B(n3968), .Z(n3970) );
  AND U4229 ( .A(n3971), .B(n3970), .Z(n4016) );
  XNOR U4230 ( .A(n4017), .B(n4016), .Z(n4019) );
  NAND U4231 ( .A(n3972), .B(n19724), .Z(n3974) );
  XOR U4232 ( .A(b[11]), .B(a[49]), .Z(n4049) );
  NAND U4233 ( .A(n19692), .B(n4049), .Z(n3973) );
  AND U4234 ( .A(n3974), .B(n3973), .Z(n4060) );
  NAND U4235 ( .A(n19838), .B(n3975), .Z(n3977) );
  XOR U4236 ( .A(b[15]), .B(a[45]), .Z(n4052) );
  NAND U4237 ( .A(n19805), .B(n4052), .Z(n3976) );
  AND U4238 ( .A(n3977), .B(n3976), .Z(n4059) );
  NAND U4239 ( .A(n35), .B(n3978), .Z(n3980) );
  XOR U4240 ( .A(b[9]), .B(a[51]), .Z(n4055) );
  NAND U4241 ( .A(n19598), .B(n4055), .Z(n3979) );
  NAND U4242 ( .A(n3980), .B(n3979), .Z(n4058) );
  XOR U4243 ( .A(n4059), .B(n4058), .Z(n4061) );
  XOR U4244 ( .A(n4060), .B(n4061), .Z(n4071) );
  NANDN U4245 ( .A(n3982), .B(n3981), .Z(n3986) );
  OR U4246 ( .A(n3984), .B(n3983), .Z(n3985) );
  AND U4247 ( .A(n3986), .B(n3985), .Z(n4070) );
  XNOR U4248 ( .A(n4071), .B(n4070), .Z(n4072) );
  NANDN U4249 ( .A(n3988), .B(n3987), .Z(n3992) );
  NANDN U4250 ( .A(n3990), .B(n3989), .Z(n3991) );
  NAND U4251 ( .A(n3992), .B(n3991), .Z(n4073) );
  XNOR U4252 ( .A(n4072), .B(n4073), .Z(n4018) );
  XOR U4253 ( .A(n4019), .B(n4018), .Z(n4077) );
  NANDN U4254 ( .A(n3994), .B(n3993), .Z(n3998) );
  NANDN U4255 ( .A(n3996), .B(n3995), .Z(n3997) );
  AND U4256 ( .A(n3998), .B(n3997), .Z(n4076) );
  XNOR U4257 ( .A(n4077), .B(n4076), .Z(n4078) );
  XOR U4258 ( .A(n4079), .B(n4078), .Z(n4011) );
  NANDN U4259 ( .A(n4000), .B(n3999), .Z(n4004) );
  NAND U4260 ( .A(n4002), .B(n4001), .Z(n4003) );
  AND U4261 ( .A(n4004), .B(n4003), .Z(n4010) );
  XNOR U4262 ( .A(n4011), .B(n4010), .Z(n4012) );
  XNOR U4263 ( .A(n4013), .B(n4012), .Z(n4082) );
  XNOR U4264 ( .A(sreg[299]), .B(n4082), .Z(n4084) );
  NANDN U4265 ( .A(sreg[298]), .B(n4005), .Z(n4009) );
  NAND U4266 ( .A(n4007), .B(n4006), .Z(n4008) );
  NAND U4267 ( .A(n4009), .B(n4008), .Z(n4083) );
  XNOR U4268 ( .A(n4084), .B(n4083), .Z(c[299]) );
  NANDN U4269 ( .A(n4011), .B(n4010), .Z(n4015) );
  NANDN U4270 ( .A(n4013), .B(n4012), .Z(n4014) );
  AND U4271 ( .A(n4015), .B(n4014), .Z(n4090) );
  NANDN U4272 ( .A(n4017), .B(n4016), .Z(n4021) );
  NAND U4273 ( .A(n4019), .B(n4018), .Z(n4020) );
  AND U4274 ( .A(n4021), .B(n4020), .Z(n4156) );
  NANDN U4275 ( .A(n4023), .B(n4022), .Z(n4027) );
  NANDN U4276 ( .A(n4025), .B(n4024), .Z(n4026) );
  AND U4277 ( .A(n4027), .B(n4026), .Z(n4122) );
  NAND U4278 ( .A(b[0]), .B(a[60]), .Z(n4028) );
  XNOR U4279 ( .A(b[1]), .B(n4028), .Z(n4030) );
  NANDN U4280 ( .A(b[0]), .B(a[59]), .Z(n4029) );
  NAND U4281 ( .A(n4030), .B(n4029), .Z(n4102) );
  NAND U4282 ( .A(n19808), .B(n4031), .Z(n4033) );
  XOR U4283 ( .A(b[13]), .B(a[48]), .Z(n4105) );
  NAND U4284 ( .A(n19768), .B(n4105), .Z(n4032) );
  AND U4285 ( .A(n4033), .B(n4032), .Z(n4100) );
  AND U4286 ( .A(b[15]), .B(a[44]), .Z(n4099) );
  XNOR U4287 ( .A(n4100), .B(n4099), .Z(n4101) );
  XNOR U4288 ( .A(n4102), .B(n4101), .Z(n4120) );
  NAND U4289 ( .A(n33), .B(n4034), .Z(n4036) );
  XOR U4290 ( .A(b[5]), .B(a[56]), .Z(n4111) );
  NAND U4291 ( .A(n19342), .B(n4111), .Z(n4035) );
  AND U4292 ( .A(n4036), .B(n4035), .Z(n4144) );
  NAND U4293 ( .A(n34), .B(n4037), .Z(n4039) );
  XOR U4294 ( .A(b[7]), .B(a[54]), .Z(n4114) );
  NAND U4295 ( .A(n19486), .B(n4114), .Z(n4038) );
  AND U4296 ( .A(n4039), .B(n4038), .Z(n4142) );
  NAND U4297 ( .A(n31), .B(n4040), .Z(n4042) );
  XOR U4298 ( .A(b[3]), .B(a[58]), .Z(n4117) );
  NAND U4299 ( .A(n32), .B(n4117), .Z(n4041) );
  NAND U4300 ( .A(n4042), .B(n4041), .Z(n4141) );
  XNOR U4301 ( .A(n4142), .B(n4141), .Z(n4143) );
  XOR U4302 ( .A(n4144), .B(n4143), .Z(n4121) );
  XOR U4303 ( .A(n4120), .B(n4121), .Z(n4123) );
  XOR U4304 ( .A(n4122), .B(n4123), .Z(n4094) );
  NANDN U4305 ( .A(n4044), .B(n4043), .Z(n4048) );
  OR U4306 ( .A(n4046), .B(n4045), .Z(n4047) );
  AND U4307 ( .A(n4048), .B(n4047), .Z(n4093) );
  XNOR U4308 ( .A(n4094), .B(n4093), .Z(n4096) );
  NAND U4309 ( .A(n4049), .B(n19724), .Z(n4051) );
  XOR U4310 ( .A(b[11]), .B(a[50]), .Z(n4126) );
  NAND U4311 ( .A(n19692), .B(n4126), .Z(n4050) );
  AND U4312 ( .A(n4051), .B(n4050), .Z(n4137) );
  NAND U4313 ( .A(n19838), .B(n4052), .Z(n4054) );
  XOR U4314 ( .A(b[15]), .B(a[46]), .Z(n4129) );
  NAND U4315 ( .A(n19805), .B(n4129), .Z(n4053) );
  AND U4316 ( .A(n4054), .B(n4053), .Z(n4136) );
  NAND U4317 ( .A(n35), .B(n4055), .Z(n4057) );
  XOR U4318 ( .A(b[9]), .B(a[52]), .Z(n4132) );
  NAND U4319 ( .A(n19598), .B(n4132), .Z(n4056) );
  NAND U4320 ( .A(n4057), .B(n4056), .Z(n4135) );
  XOR U4321 ( .A(n4136), .B(n4135), .Z(n4138) );
  XOR U4322 ( .A(n4137), .B(n4138), .Z(n4148) );
  NANDN U4323 ( .A(n4059), .B(n4058), .Z(n4063) );
  OR U4324 ( .A(n4061), .B(n4060), .Z(n4062) );
  AND U4325 ( .A(n4063), .B(n4062), .Z(n4147) );
  XNOR U4326 ( .A(n4148), .B(n4147), .Z(n4149) );
  NANDN U4327 ( .A(n4065), .B(n4064), .Z(n4069) );
  NANDN U4328 ( .A(n4067), .B(n4066), .Z(n4068) );
  NAND U4329 ( .A(n4069), .B(n4068), .Z(n4150) );
  XNOR U4330 ( .A(n4149), .B(n4150), .Z(n4095) );
  XOR U4331 ( .A(n4096), .B(n4095), .Z(n4154) );
  NANDN U4332 ( .A(n4071), .B(n4070), .Z(n4075) );
  NANDN U4333 ( .A(n4073), .B(n4072), .Z(n4074) );
  AND U4334 ( .A(n4075), .B(n4074), .Z(n4153) );
  XNOR U4335 ( .A(n4154), .B(n4153), .Z(n4155) );
  XOR U4336 ( .A(n4156), .B(n4155), .Z(n4088) );
  NANDN U4337 ( .A(n4077), .B(n4076), .Z(n4081) );
  NAND U4338 ( .A(n4079), .B(n4078), .Z(n4080) );
  AND U4339 ( .A(n4081), .B(n4080), .Z(n4087) );
  XNOR U4340 ( .A(n4088), .B(n4087), .Z(n4089) );
  XNOR U4341 ( .A(n4090), .B(n4089), .Z(n4159) );
  XNOR U4342 ( .A(sreg[300]), .B(n4159), .Z(n4161) );
  NANDN U4343 ( .A(sreg[299]), .B(n4082), .Z(n4086) );
  NAND U4344 ( .A(n4084), .B(n4083), .Z(n4085) );
  NAND U4345 ( .A(n4086), .B(n4085), .Z(n4160) );
  XNOR U4346 ( .A(n4161), .B(n4160), .Z(c[300]) );
  NANDN U4347 ( .A(n4088), .B(n4087), .Z(n4092) );
  NANDN U4348 ( .A(n4090), .B(n4089), .Z(n4091) );
  AND U4349 ( .A(n4092), .B(n4091), .Z(n4167) );
  NANDN U4350 ( .A(n4094), .B(n4093), .Z(n4098) );
  NAND U4351 ( .A(n4096), .B(n4095), .Z(n4097) );
  AND U4352 ( .A(n4098), .B(n4097), .Z(n4233) );
  NANDN U4353 ( .A(n4100), .B(n4099), .Z(n4104) );
  NANDN U4354 ( .A(n4102), .B(n4101), .Z(n4103) );
  AND U4355 ( .A(n4104), .B(n4103), .Z(n4199) );
  NAND U4356 ( .A(n19808), .B(n4105), .Z(n4107) );
  XOR U4357 ( .A(b[13]), .B(a[49]), .Z(n4185) );
  NAND U4358 ( .A(n19768), .B(n4185), .Z(n4106) );
  AND U4359 ( .A(n4107), .B(n4106), .Z(n4177) );
  AND U4360 ( .A(b[15]), .B(a[45]), .Z(n4176) );
  XNOR U4361 ( .A(n4177), .B(n4176), .Z(n4178) );
  NAND U4362 ( .A(b[0]), .B(a[61]), .Z(n4108) );
  XNOR U4363 ( .A(b[1]), .B(n4108), .Z(n4110) );
  NANDN U4364 ( .A(b[0]), .B(a[60]), .Z(n4109) );
  NAND U4365 ( .A(n4110), .B(n4109), .Z(n4179) );
  XNOR U4366 ( .A(n4178), .B(n4179), .Z(n4197) );
  NAND U4367 ( .A(n33), .B(n4111), .Z(n4113) );
  XOR U4368 ( .A(b[5]), .B(a[57]), .Z(n4188) );
  NAND U4369 ( .A(n19342), .B(n4188), .Z(n4112) );
  AND U4370 ( .A(n4113), .B(n4112), .Z(n4221) );
  NAND U4371 ( .A(n34), .B(n4114), .Z(n4116) );
  XOR U4372 ( .A(b[7]), .B(a[55]), .Z(n4191) );
  NAND U4373 ( .A(n19486), .B(n4191), .Z(n4115) );
  AND U4374 ( .A(n4116), .B(n4115), .Z(n4219) );
  NAND U4375 ( .A(n31), .B(n4117), .Z(n4119) );
  XOR U4376 ( .A(b[3]), .B(a[59]), .Z(n4194) );
  NAND U4377 ( .A(n32), .B(n4194), .Z(n4118) );
  NAND U4378 ( .A(n4119), .B(n4118), .Z(n4218) );
  XNOR U4379 ( .A(n4219), .B(n4218), .Z(n4220) );
  XOR U4380 ( .A(n4221), .B(n4220), .Z(n4198) );
  XOR U4381 ( .A(n4197), .B(n4198), .Z(n4200) );
  XOR U4382 ( .A(n4199), .B(n4200), .Z(n4171) );
  NANDN U4383 ( .A(n4121), .B(n4120), .Z(n4125) );
  OR U4384 ( .A(n4123), .B(n4122), .Z(n4124) );
  AND U4385 ( .A(n4125), .B(n4124), .Z(n4170) );
  XNOR U4386 ( .A(n4171), .B(n4170), .Z(n4173) );
  NAND U4387 ( .A(n4126), .B(n19724), .Z(n4128) );
  XOR U4388 ( .A(b[11]), .B(a[51]), .Z(n4203) );
  NAND U4389 ( .A(n19692), .B(n4203), .Z(n4127) );
  AND U4390 ( .A(n4128), .B(n4127), .Z(n4214) );
  NAND U4391 ( .A(n19838), .B(n4129), .Z(n4131) );
  XOR U4392 ( .A(b[15]), .B(a[47]), .Z(n4206) );
  NAND U4393 ( .A(n19805), .B(n4206), .Z(n4130) );
  AND U4394 ( .A(n4131), .B(n4130), .Z(n4213) );
  NAND U4395 ( .A(n35), .B(n4132), .Z(n4134) );
  XOR U4396 ( .A(b[9]), .B(a[53]), .Z(n4209) );
  NAND U4397 ( .A(n19598), .B(n4209), .Z(n4133) );
  NAND U4398 ( .A(n4134), .B(n4133), .Z(n4212) );
  XOR U4399 ( .A(n4213), .B(n4212), .Z(n4215) );
  XOR U4400 ( .A(n4214), .B(n4215), .Z(n4225) );
  NANDN U4401 ( .A(n4136), .B(n4135), .Z(n4140) );
  OR U4402 ( .A(n4138), .B(n4137), .Z(n4139) );
  AND U4403 ( .A(n4140), .B(n4139), .Z(n4224) );
  XNOR U4404 ( .A(n4225), .B(n4224), .Z(n4226) );
  NANDN U4405 ( .A(n4142), .B(n4141), .Z(n4146) );
  NANDN U4406 ( .A(n4144), .B(n4143), .Z(n4145) );
  NAND U4407 ( .A(n4146), .B(n4145), .Z(n4227) );
  XNOR U4408 ( .A(n4226), .B(n4227), .Z(n4172) );
  XOR U4409 ( .A(n4173), .B(n4172), .Z(n4231) );
  NANDN U4410 ( .A(n4148), .B(n4147), .Z(n4152) );
  NANDN U4411 ( .A(n4150), .B(n4149), .Z(n4151) );
  AND U4412 ( .A(n4152), .B(n4151), .Z(n4230) );
  XNOR U4413 ( .A(n4231), .B(n4230), .Z(n4232) );
  XOR U4414 ( .A(n4233), .B(n4232), .Z(n4165) );
  NANDN U4415 ( .A(n4154), .B(n4153), .Z(n4158) );
  NAND U4416 ( .A(n4156), .B(n4155), .Z(n4157) );
  AND U4417 ( .A(n4158), .B(n4157), .Z(n4164) );
  XNOR U4418 ( .A(n4165), .B(n4164), .Z(n4166) );
  XNOR U4419 ( .A(n4167), .B(n4166), .Z(n4236) );
  XNOR U4420 ( .A(sreg[301]), .B(n4236), .Z(n4238) );
  NANDN U4421 ( .A(sreg[300]), .B(n4159), .Z(n4163) );
  NAND U4422 ( .A(n4161), .B(n4160), .Z(n4162) );
  NAND U4423 ( .A(n4163), .B(n4162), .Z(n4237) );
  XNOR U4424 ( .A(n4238), .B(n4237), .Z(c[301]) );
  NANDN U4425 ( .A(n4165), .B(n4164), .Z(n4169) );
  NANDN U4426 ( .A(n4167), .B(n4166), .Z(n4168) );
  AND U4427 ( .A(n4169), .B(n4168), .Z(n4244) );
  NANDN U4428 ( .A(n4171), .B(n4170), .Z(n4175) );
  NAND U4429 ( .A(n4173), .B(n4172), .Z(n4174) );
  AND U4430 ( .A(n4175), .B(n4174), .Z(n4310) );
  NANDN U4431 ( .A(n4177), .B(n4176), .Z(n4181) );
  NANDN U4432 ( .A(n4179), .B(n4178), .Z(n4180) );
  AND U4433 ( .A(n4181), .B(n4180), .Z(n4276) );
  NAND U4434 ( .A(b[0]), .B(a[62]), .Z(n4182) );
  XNOR U4435 ( .A(b[1]), .B(n4182), .Z(n4184) );
  NANDN U4436 ( .A(b[0]), .B(a[61]), .Z(n4183) );
  NAND U4437 ( .A(n4184), .B(n4183), .Z(n4256) );
  NAND U4438 ( .A(n19808), .B(n4185), .Z(n4187) );
  XOR U4439 ( .A(b[13]), .B(a[50]), .Z(n4262) );
  NAND U4440 ( .A(n19768), .B(n4262), .Z(n4186) );
  AND U4441 ( .A(n4187), .B(n4186), .Z(n4254) );
  AND U4442 ( .A(b[15]), .B(a[46]), .Z(n4253) );
  XNOR U4443 ( .A(n4254), .B(n4253), .Z(n4255) );
  XNOR U4444 ( .A(n4256), .B(n4255), .Z(n4274) );
  NAND U4445 ( .A(n33), .B(n4188), .Z(n4190) );
  XOR U4446 ( .A(b[5]), .B(a[58]), .Z(n4265) );
  NAND U4447 ( .A(n19342), .B(n4265), .Z(n4189) );
  AND U4448 ( .A(n4190), .B(n4189), .Z(n4298) );
  NAND U4449 ( .A(n34), .B(n4191), .Z(n4193) );
  XOR U4450 ( .A(b[7]), .B(a[56]), .Z(n4268) );
  NAND U4451 ( .A(n19486), .B(n4268), .Z(n4192) );
  AND U4452 ( .A(n4193), .B(n4192), .Z(n4296) );
  NAND U4453 ( .A(n31), .B(n4194), .Z(n4196) );
  XOR U4454 ( .A(b[3]), .B(a[60]), .Z(n4271) );
  NAND U4455 ( .A(n32), .B(n4271), .Z(n4195) );
  NAND U4456 ( .A(n4196), .B(n4195), .Z(n4295) );
  XNOR U4457 ( .A(n4296), .B(n4295), .Z(n4297) );
  XOR U4458 ( .A(n4298), .B(n4297), .Z(n4275) );
  XOR U4459 ( .A(n4274), .B(n4275), .Z(n4277) );
  XOR U4460 ( .A(n4276), .B(n4277), .Z(n4248) );
  NANDN U4461 ( .A(n4198), .B(n4197), .Z(n4202) );
  OR U4462 ( .A(n4200), .B(n4199), .Z(n4201) );
  AND U4463 ( .A(n4202), .B(n4201), .Z(n4247) );
  XNOR U4464 ( .A(n4248), .B(n4247), .Z(n4250) );
  NAND U4465 ( .A(n4203), .B(n19724), .Z(n4205) );
  XOR U4466 ( .A(b[11]), .B(a[52]), .Z(n4280) );
  NAND U4467 ( .A(n19692), .B(n4280), .Z(n4204) );
  AND U4468 ( .A(n4205), .B(n4204), .Z(n4291) );
  NAND U4469 ( .A(n19838), .B(n4206), .Z(n4208) );
  XOR U4470 ( .A(b[15]), .B(a[48]), .Z(n4283) );
  NAND U4471 ( .A(n19805), .B(n4283), .Z(n4207) );
  AND U4472 ( .A(n4208), .B(n4207), .Z(n4290) );
  NAND U4473 ( .A(n35), .B(n4209), .Z(n4211) );
  XOR U4474 ( .A(b[9]), .B(a[54]), .Z(n4286) );
  NAND U4475 ( .A(n19598), .B(n4286), .Z(n4210) );
  NAND U4476 ( .A(n4211), .B(n4210), .Z(n4289) );
  XOR U4477 ( .A(n4290), .B(n4289), .Z(n4292) );
  XOR U4478 ( .A(n4291), .B(n4292), .Z(n4302) );
  NANDN U4479 ( .A(n4213), .B(n4212), .Z(n4217) );
  OR U4480 ( .A(n4215), .B(n4214), .Z(n4216) );
  AND U4481 ( .A(n4217), .B(n4216), .Z(n4301) );
  XNOR U4482 ( .A(n4302), .B(n4301), .Z(n4303) );
  NANDN U4483 ( .A(n4219), .B(n4218), .Z(n4223) );
  NANDN U4484 ( .A(n4221), .B(n4220), .Z(n4222) );
  NAND U4485 ( .A(n4223), .B(n4222), .Z(n4304) );
  XNOR U4486 ( .A(n4303), .B(n4304), .Z(n4249) );
  XOR U4487 ( .A(n4250), .B(n4249), .Z(n4308) );
  NANDN U4488 ( .A(n4225), .B(n4224), .Z(n4229) );
  NANDN U4489 ( .A(n4227), .B(n4226), .Z(n4228) );
  AND U4490 ( .A(n4229), .B(n4228), .Z(n4307) );
  XNOR U4491 ( .A(n4308), .B(n4307), .Z(n4309) );
  XOR U4492 ( .A(n4310), .B(n4309), .Z(n4242) );
  NANDN U4493 ( .A(n4231), .B(n4230), .Z(n4235) );
  NAND U4494 ( .A(n4233), .B(n4232), .Z(n4234) );
  AND U4495 ( .A(n4235), .B(n4234), .Z(n4241) );
  XNOR U4496 ( .A(n4242), .B(n4241), .Z(n4243) );
  XNOR U4497 ( .A(n4244), .B(n4243), .Z(n4313) );
  XNOR U4498 ( .A(sreg[302]), .B(n4313), .Z(n4315) );
  NANDN U4499 ( .A(sreg[301]), .B(n4236), .Z(n4240) );
  NAND U4500 ( .A(n4238), .B(n4237), .Z(n4239) );
  NAND U4501 ( .A(n4240), .B(n4239), .Z(n4314) );
  XNOR U4502 ( .A(n4315), .B(n4314), .Z(c[302]) );
  NANDN U4503 ( .A(n4242), .B(n4241), .Z(n4246) );
  NANDN U4504 ( .A(n4244), .B(n4243), .Z(n4245) );
  AND U4505 ( .A(n4246), .B(n4245), .Z(n4321) );
  NANDN U4506 ( .A(n4248), .B(n4247), .Z(n4252) );
  NAND U4507 ( .A(n4250), .B(n4249), .Z(n4251) );
  AND U4508 ( .A(n4252), .B(n4251), .Z(n4387) );
  NANDN U4509 ( .A(n4254), .B(n4253), .Z(n4258) );
  NANDN U4510 ( .A(n4256), .B(n4255), .Z(n4257) );
  AND U4511 ( .A(n4258), .B(n4257), .Z(n4353) );
  NAND U4512 ( .A(b[0]), .B(a[63]), .Z(n4259) );
  XNOR U4513 ( .A(b[1]), .B(n4259), .Z(n4261) );
  NANDN U4514 ( .A(b[0]), .B(a[62]), .Z(n4260) );
  NAND U4515 ( .A(n4261), .B(n4260), .Z(n4333) );
  NAND U4516 ( .A(n19808), .B(n4262), .Z(n4264) );
  XOR U4517 ( .A(b[13]), .B(a[51]), .Z(n4339) );
  NAND U4518 ( .A(n19768), .B(n4339), .Z(n4263) );
  AND U4519 ( .A(n4264), .B(n4263), .Z(n4331) );
  AND U4520 ( .A(b[15]), .B(a[47]), .Z(n4330) );
  XNOR U4521 ( .A(n4331), .B(n4330), .Z(n4332) );
  XNOR U4522 ( .A(n4333), .B(n4332), .Z(n4351) );
  NAND U4523 ( .A(n33), .B(n4265), .Z(n4267) );
  XOR U4524 ( .A(b[5]), .B(a[59]), .Z(n4342) );
  NAND U4525 ( .A(n19342), .B(n4342), .Z(n4266) );
  AND U4526 ( .A(n4267), .B(n4266), .Z(n4375) );
  NAND U4527 ( .A(n34), .B(n4268), .Z(n4270) );
  XOR U4528 ( .A(b[7]), .B(a[57]), .Z(n4345) );
  NAND U4529 ( .A(n19486), .B(n4345), .Z(n4269) );
  AND U4530 ( .A(n4270), .B(n4269), .Z(n4373) );
  NAND U4531 ( .A(n31), .B(n4271), .Z(n4273) );
  XOR U4532 ( .A(b[3]), .B(a[61]), .Z(n4348) );
  NAND U4533 ( .A(n32), .B(n4348), .Z(n4272) );
  NAND U4534 ( .A(n4273), .B(n4272), .Z(n4372) );
  XNOR U4535 ( .A(n4373), .B(n4372), .Z(n4374) );
  XOR U4536 ( .A(n4375), .B(n4374), .Z(n4352) );
  XOR U4537 ( .A(n4351), .B(n4352), .Z(n4354) );
  XOR U4538 ( .A(n4353), .B(n4354), .Z(n4325) );
  NANDN U4539 ( .A(n4275), .B(n4274), .Z(n4279) );
  OR U4540 ( .A(n4277), .B(n4276), .Z(n4278) );
  AND U4541 ( .A(n4279), .B(n4278), .Z(n4324) );
  XNOR U4542 ( .A(n4325), .B(n4324), .Z(n4327) );
  NAND U4543 ( .A(n4280), .B(n19724), .Z(n4282) );
  XOR U4544 ( .A(b[11]), .B(a[53]), .Z(n4357) );
  NAND U4545 ( .A(n19692), .B(n4357), .Z(n4281) );
  AND U4546 ( .A(n4282), .B(n4281), .Z(n4368) );
  NAND U4547 ( .A(n19838), .B(n4283), .Z(n4285) );
  XOR U4548 ( .A(b[15]), .B(a[49]), .Z(n4360) );
  NAND U4549 ( .A(n19805), .B(n4360), .Z(n4284) );
  AND U4550 ( .A(n4285), .B(n4284), .Z(n4367) );
  NAND U4551 ( .A(n35), .B(n4286), .Z(n4288) );
  XOR U4552 ( .A(b[9]), .B(a[55]), .Z(n4363) );
  NAND U4553 ( .A(n19598), .B(n4363), .Z(n4287) );
  NAND U4554 ( .A(n4288), .B(n4287), .Z(n4366) );
  XOR U4555 ( .A(n4367), .B(n4366), .Z(n4369) );
  XOR U4556 ( .A(n4368), .B(n4369), .Z(n4379) );
  NANDN U4557 ( .A(n4290), .B(n4289), .Z(n4294) );
  OR U4558 ( .A(n4292), .B(n4291), .Z(n4293) );
  AND U4559 ( .A(n4294), .B(n4293), .Z(n4378) );
  XNOR U4560 ( .A(n4379), .B(n4378), .Z(n4380) );
  NANDN U4561 ( .A(n4296), .B(n4295), .Z(n4300) );
  NANDN U4562 ( .A(n4298), .B(n4297), .Z(n4299) );
  NAND U4563 ( .A(n4300), .B(n4299), .Z(n4381) );
  XNOR U4564 ( .A(n4380), .B(n4381), .Z(n4326) );
  XOR U4565 ( .A(n4327), .B(n4326), .Z(n4385) );
  NANDN U4566 ( .A(n4302), .B(n4301), .Z(n4306) );
  NANDN U4567 ( .A(n4304), .B(n4303), .Z(n4305) );
  AND U4568 ( .A(n4306), .B(n4305), .Z(n4384) );
  XNOR U4569 ( .A(n4385), .B(n4384), .Z(n4386) );
  XOR U4570 ( .A(n4387), .B(n4386), .Z(n4319) );
  NANDN U4571 ( .A(n4308), .B(n4307), .Z(n4312) );
  NAND U4572 ( .A(n4310), .B(n4309), .Z(n4311) );
  AND U4573 ( .A(n4312), .B(n4311), .Z(n4318) );
  XNOR U4574 ( .A(n4319), .B(n4318), .Z(n4320) );
  XNOR U4575 ( .A(n4321), .B(n4320), .Z(n4390) );
  XNOR U4576 ( .A(sreg[303]), .B(n4390), .Z(n4392) );
  NANDN U4577 ( .A(sreg[302]), .B(n4313), .Z(n4317) );
  NAND U4578 ( .A(n4315), .B(n4314), .Z(n4316) );
  NAND U4579 ( .A(n4317), .B(n4316), .Z(n4391) );
  XNOR U4580 ( .A(n4392), .B(n4391), .Z(c[303]) );
  NANDN U4581 ( .A(n4319), .B(n4318), .Z(n4323) );
  NANDN U4582 ( .A(n4321), .B(n4320), .Z(n4322) );
  AND U4583 ( .A(n4323), .B(n4322), .Z(n4398) );
  NANDN U4584 ( .A(n4325), .B(n4324), .Z(n4329) );
  NAND U4585 ( .A(n4327), .B(n4326), .Z(n4328) );
  AND U4586 ( .A(n4329), .B(n4328), .Z(n4464) );
  NANDN U4587 ( .A(n4331), .B(n4330), .Z(n4335) );
  NANDN U4588 ( .A(n4333), .B(n4332), .Z(n4334) );
  AND U4589 ( .A(n4335), .B(n4334), .Z(n4451) );
  NAND U4590 ( .A(b[0]), .B(a[64]), .Z(n4336) );
  XNOR U4591 ( .A(b[1]), .B(n4336), .Z(n4338) );
  NANDN U4592 ( .A(b[0]), .B(a[63]), .Z(n4337) );
  NAND U4593 ( .A(n4338), .B(n4337), .Z(n4431) );
  NAND U4594 ( .A(n19808), .B(n4339), .Z(n4341) );
  XOR U4595 ( .A(b[13]), .B(a[52]), .Z(n4437) );
  NAND U4596 ( .A(n19768), .B(n4437), .Z(n4340) );
  AND U4597 ( .A(n4341), .B(n4340), .Z(n4429) );
  AND U4598 ( .A(b[15]), .B(a[48]), .Z(n4428) );
  XNOR U4599 ( .A(n4429), .B(n4428), .Z(n4430) );
  XNOR U4600 ( .A(n4431), .B(n4430), .Z(n4449) );
  NAND U4601 ( .A(n33), .B(n4342), .Z(n4344) );
  XOR U4602 ( .A(b[5]), .B(a[60]), .Z(n4440) );
  NAND U4603 ( .A(n19342), .B(n4440), .Z(n4343) );
  AND U4604 ( .A(n4344), .B(n4343), .Z(n4425) );
  NAND U4605 ( .A(n34), .B(n4345), .Z(n4347) );
  XOR U4606 ( .A(b[7]), .B(a[58]), .Z(n4443) );
  NAND U4607 ( .A(n19486), .B(n4443), .Z(n4346) );
  AND U4608 ( .A(n4347), .B(n4346), .Z(n4423) );
  NAND U4609 ( .A(n31), .B(n4348), .Z(n4350) );
  XOR U4610 ( .A(b[3]), .B(a[62]), .Z(n4446) );
  NAND U4611 ( .A(n32), .B(n4446), .Z(n4349) );
  NAND U4612 ( .A(n4350), .B(n4349), .Z(n4422) );
  XNOR U4613 ( .A(n4423), .B(n4422), .Z(n4424) );
  XOR U4614 ( .A(n4425), .B(n4424), .Z(n4450) );
  XOR U4615 ( .A(n4449), .B(n4450), .Z(n4452) );
  XOR U4616 ( .A(n4451), .B(n4452), .Z(n4402) );
  NANDN U4617 ( .A(n4352), .B(n4351), .Z(n4356) );
  OR U4618 ( .A(n4354), .B(n4353), .Z(n4355) );
  AND U4619 ( .A(n4356), .B(n4355), .Z(n4401) );
  XNOR U4620 ( .A(n4402), .B(n4401), .Z(n4404) );
  NAND U4621 ( .A(n4357), .B(n19724), .Z(n4359) );
  XOR U4622 ( .A(b[11]), .B(a[54]), .Z(n4407) );
  NAND U4623 ( .A(n19692), .B(n4407), .Z(n4358) );
  AND U4624 ( .A(n4359), .B(n4358), .Z(n4418) );
  NAND U4625 ( .A(n19838), .B(n4360), .Z(n4362) );
  XOR U4626 ( .A(b[15]), .B(a[50]), .Z(n4410) );
  NAND U4627 ( .A(n19805), .B(n4410), .Z(n4361) );
  AND U4628 ( .A(n4362), .B(n4361), .Z(n4417) );
  NAND U4629 ( .A(n35), .B(n4363), .Z(n4365) );
  XOR U4630 ( .A(b[9]), .B(a[56]), .Z(n4413) );
  NAND U4631 ( .A(n19598), .B(n4413), .Z(n4364) );
  NAND U4632 ( .A(n4365), .B(n4364), .Z(n4416) );
  XOR U4633 ( .A(n4417), .B(n4416), .Z(n4419) );
  XOR U4634 ( .A(n4418), .B(n4419), .Z(n4456) );
  NANDN U4635 ( .A(n4367), .B(n4366), .Z(n4371) );
  OR U4636 ( .A(n4369), .B(n4368), .Z(n4370) );
  AND U4637 ( .A(n4371), .B(n4370), .Z(n4455) );
  XNOR U4638 ( .A(n4456), .B(n4455), .Z(n4457) );
  NANDN U4639 ( .A(n4373), .B(n4372), .Z(n4377) );
  NANDN U4640 ( .A(n4375), .B(n4374), .Z(n4376) );
  NAND U4641 ( .A(n4377), .B(n4376), .Z(n4458) );
  XNOR U4642 ( .A(n4457), .B(n4458), .Z(n4403) );
  XOR U4643 ( .A(n4404), .B(n4403), .Z(n4462) );
  NANDN U4644 ( .A(n4379), .B(n4378), .Z(n4383) );
  NANDN U4645 ( .A(n4381), .B(n4380), .Z(n4382) );
  AND U4646 ( .A(n4383), .B(n4382), .Z(n4461) );
  XNOR U4647 ( .A(n4462), .B(n4461), .Z(n4463) );
  XOR U4648 ( .A(n4464), .B(n4463), .Z(n4396) );
  NANDN U4649 ( .A(n4385), .B(n4384), .Z(n4389) );
  NAND U4650 ( .A(n4387), .B(n4386), .Z(n4388) );
  AND U4651 ( .A(n4389), .B(n4388), .Z(n4395) );
  XNOR U4652 ( .A(n4396), .B(n4395), .Z(n4397) );
  XNOR U4653 ( .A(n4398), .B(n4397), .Z(n4467) );
  XNOR U4654 ( .A(sreg[304]), .B(n4467), .Z(n4469) );
  NANDN U4655 ( .A(sreg[303]), .B(n4390), .Z(n4394) );
  NAND U4656 ( .A(n4392), .B(n4391), .Z(n4393) );
  NAND U4657 ( .A(n4394), .B(n4393), .Z(n4468) );
  XNOR U4658 ( .A(n4469), .B(n4468), .Z(c[304]) );
  NANDN U4659 ( .A(n4396), .B(n4395), .Z(n4400) );
  NANDN U4660 ( .A(n4398), .B(n4397), .Z(n4399) );
  AND U4661 ( .A(n4400), .B(n4399), .Z(n4475) );
  NANDN U4662 ( .A(n4402), .B(n4401), .Z(n4406) );
  NAND U4663 ( .A(n4404), .B(n4403), .Z(n4405) );
  AND U4664 ( .A(n4406), .B(n4405), .Z(n4541) );
  NAND U4665 ( .A(n4407), .B(n19724), .Z(n4409) );
  XOR U4666 ( .A(b[11]), .B(a[55]), .Z(n4511) );
  NAND U4667 ( .A(n19692), .B(n4511), .Z(n4408) );
  AND U4668 ( .A(n4409), .B(n4408), .Z(n4522) );
  NAND U4669 ( .A(n19838), .B(n4410), .Z(n4412) );
  XOR U4670 ( .A(b[15]), .B(a[51]), .Z(n4514) );
  NAND U4671 ( .A(n19805), .B(n4514), .Z(n4411) );
  AND U4672 ( .A(n4412), .B(n4411), .Z(n4521) );
  NAND U4673 ( .A(n35), .B(n4413), .Z(n4415) );
  XOR U4674 ( .A(b[9]), .B(a[57]), .Z(n4517) );
  NAND U4675 ( .A(n19598), .B(n4517), .Z(n4414) );
  NAND U4676 ( .A(n4415), .B(n4414), .Z(n4520) );
  XOR U4677 ( .A(n4521), .B(n4520), .Z(n4523) );
  XOR U4678 ( .A(n4522), .B(n4523), .Z(n4533) );
  NANDN U4679 ( .A(n4417), .B(n4416), .Z(n4421) );
  OR U4680 ( .A(n4419), .B(n4418), .Z(n4420) );
  AND U4681 ( .A(n4421), .B(n4420), .Z(n4532) );
  XNOR U4682 ( .A(n4533), .B(n4532), .Z(n4534) );
  NANDN U4683 ( .A(n4423), .B(n4422), .Z(n4427) );
  NANDN U4684 ( .A(n4425), .B(n4424), .Z(n4426) );
  NAND U4685 ( .A(n4427), .B(n4426), .Z(n4535) );
  XNOR U4686 ( .A(n4534), .B(n4535), .Z(n4481) );
  NANDN U4687 ( .A(n4429), .B(n4428), .Z(n4433) );
  NANDN U4688 ( .A(n4431), .B(n4430), .Z(n4432) );
  AND U4689 ( .A(n4433), .B(n4432), .Z(n4507) );
  NAND U4690 ( .A(b[0]), .B(a[65]), .Z(n4434) );
  XNOR U4691 ( .A(b[1]), .B(n4434), .Z(n4436) );
  NANDN U4692 ( .A(b[0]), .B(a[64]), .Z(n4435) );
  NAND U4693 ( .A(n4436), .B(n4435), .Z(n4487) );
  NAND U4694 ( .A(n19808), .B(n4437), .Z(n4439) );
  XOR U4695 ( .A(b[13]), .B(a[53]), .Z(n4493) );
  NAND U4696 ( .A(n19768), .B(n4493), .Z(n4438) );
  AND U4697 ( .A(n4439), .B(n4438), .Z(n4485) );
  AND U4698 ( .A(b[15]), .B(a[49]), .Z(n4484) );
  XNOR U4699 ( .A(n4485), .B(n4484), .Z(n4486) );
  XNOR U4700 ( .A(n4487), .B(n4486), .Z(n4505) );
  NAND U4701 ( .A(n33), .B(n4440), .Z(n4442) );
  XOR U4702 ( .A(b[5]), .B(a[61]), .Z(n4496) );
  NAND U4703 ( .A(n19342), .B(n4496), .Z(n4441) );
  AND U4704 ( .A(n4442), .B(n4441), .Z(n4529) );
  NAND U4705 ( .A(n34), .B(n4443), .Z(n4445) );
  XOR U4706 ( .A(b[7]), .B(a[59]), .Z(n4499) );
  NAND U4707 ( .A(n19486), .B(n4499), .Z(n4444) );
  AND U4708 ( .A(n4445), .B(n4444), .Z(n4527) );
  NAND U4709 ( .A(n31), .B(n4446), .Z(n4448) );
  XOR U4710 ( .A(b[3]), .B(a[63]), .Z(n4502) );
  NAND U4711 ( .A(n32), .B(n4502), .Z(n4447) );
  NAND U4712 ( .A(n4448), .B(n4447), .Z(n4526) );
  XNOR U4713 ( .A(n4527), .B(n4526), .Z(n4528) );
  XOR U4714 ( .A(n4529), .B(n4528), .Z(n4506) );
  XOR U4715 ( .A(n4505), .B(n4506), .Z(n4508) );
  XOR U4716 ( .A(n4507), .B(n4508), .Z(n4479) );
  NANDN U4717 ( .A(n4450), .B(n4449), .Z(n4454) );
  OR U4718 ( .A(n4452), .B(n4451), .Z(n4453) );
  AND U4719 ( .A(n4454), .B(n4453), .Z(n4478) );
  XNOR U4720 ( .A(n4479), .B(n4478), .Z(n4480) );
  XOR U4721 ( .A(n4481), .B(n4480), .Z(n4539) );
  NANDN U4722 ( .A(n4456), .B(n4455), .Z(n4460) );
  NANDN U4723 ( .A(n4458), .B(n4457), .Z(n4459) );
  AND U4724 ( .A(n4460), .B(n4459), .Z(n4538) );
  XNOR U4725 ( .A(n4539), .B(n4538), .Z(n4540) );
  XOR U4726 ( .A(n4541), .B(n4540), .Z(n4473) );
  NANDN U4727 ( .A(n4462), .B(n4461), .Z(n4466) );
  NAND U4728 ( .A(n4464), .B(n4463), .Z(n4465) );
  AND U4729 ( .A(n4466), .B(n4465), .Z(n4472) );
  XNOR U4730 ( .A(n4473), .B(n4472), .Z(n4474) );
  XNOR U4731 ( .A(n4475), .B(n4474), .Z(n4544) );
  XNOR U4732 ( .A(sreg[305]), .B(n4544), .Z(n4546) );
  NANDN U4733 ( .A(sreg[304]), .B(n4467), .Z(n4471) );
  NAND U4734 ( .A(n4469), .B(n4468), .Z(n4470) );
  NAND U4735 ( .A(n4471), .B(n4470), .Z(n4545) );
  XNOR U4736 ( .A(n4546), .B(n4545), .Z(c[305]) );
  NANDN U4737 ( .A(n4473), .B(n4472), .Z(n4477) );
  NANDN U4738 ( .A(n4475), .B(n4474), .Z(n4476) );
  AND U4739 ( .A(n4477), .B(n4476), .Z(n4552) );
  NANDN U4740 ( .A(n4479), .B(n4478), .Z(n4483) );
  NAND U4741 ( .A(n4481), .B(n4480), .Z(n4482) );
  AND U4742 ( .A(n4483), .B(n4482), .Z(n4618) );
  NANDN U4743 ( .A(n4485), .B(n4484), .Z(n4489) );
  NANDN U4744 ( .A(n4487), .B(n4486), .Z(n4488) );
  AND U4745 ( .A(n4489), .B(n4488), .Z(n4584) );
  NAND U4746 ( .A(b[0]), .B(a[66]), .Z(n4490) );
  XNOR U4747 ( .A(b[1]), .B(n4490), .Z(n4492) );
  NANDN U4748 ( .A(b[0]), .B(a[65]), .Z(n4491) );
  NAND U4749 ( .A(n4492), .B(n4491), .Z(n4564) );
  NAND U4750 ( .A(n19808), .B(n4493), .Z(n4495) );
  XOR U4751 ( .A(b[13]), .B(a[54]), .Z(n4567) );
  NAND U4752 ( .A(n19768), .B(n4567), .Z(n4494) );
  AND U4753 ( .A(n4495), .B(n4494), .Z(n4562) );
  AND U4754 ( .A(b[15]), .B(a[50]), .Z(n4561) );
  XNOR U4755 ( .A(n4562), .B(n4561), .Z(n4563) );
  XNOR U4756 ( .A(n4564), .B(n4563), .Z(n4582) );
  NAND U4757 ( .A(n33), .B(n4496), .Z(n4498) );
  XOR U4758 ( .A(b[5]), .B(a[62]), .Z(n4573) );
  NAND U4759 ( .A(n19342), .B(n4573), .Z(n4497) );
  AND U4760 ( .A(n4498), .B(n4497), .Z(n4606) );
  NAND U4761 ( .A(n34), .B(n4499), .Z(n4501) );
  XOR U4762 ( .A(b[7]), .B(a[60]), .Z(n4576) );
  NAND U4763 ( .A(n19486), .B(n4576), .Z(n4500) );
  AND U4764 ( .A(n4501), .B(n4500), .Z(n4604) );
  NAND U4765 ( .A(n31), .B(n4502), .Z(n4504) );
  XOR U4766 ( .A(b[3]), .B(a[64]), .Z(n4579) );
  NAND U4767 ( .A(n32), .B(n4579), .Z(n4503) );
  NAND U4768 ( .A(n4504), .B(n4503), .Z(n4603) );
  XNOR U4769 ( .A(n4604), .B(n4603), .Z(n4605) );
  XOR U4770 ( .A(n4606), .B(n4605), .Z(n4583) );
  XOR U4771 ( .A(n4582), .B(n4583), .Z(n4585) );
  XOR U4772 ( .A(n4584), .B(n4585), .Z(n4556) );
  NANDN U4773 ( .A(n4506), .B(n4505), .Z(n4510) );
  OR U4774 ( .A(n4508), .B(n4507), .Z(n4509) );
  AND U4775 ( .A(n4510), .B(n4509), .Z(n4555) );
  XNOR U4776 ( .A(n4556), .B(n4555), .Z(n4558) );
  NAND U4777 ( .A(n4511), .B(n19724), .Z(n4513) );
  XOR U4778 ( .A(b[11]), .B(a[56]), .Z(n4588) );
  NAND U4779 ( .A(n19692), .B(n4588), .Z(n4512) );
  AND U4780 ( .A(n4513), .B(n4512), .Z(n4599) );
  NAND U4781 ( .A(n19838), .B(n4514), .Z(n4516) );
  XOR U4782 ( .A(b[15]), .B(a[52]), .Z(n4591) );
  NAND U4783 ( .A(n19805), .B(n4591), .Z(n4515) );
  AND U4784 ( .A(n4516), .B(n4515), .Z(n4598) );
  NAND U4785 ( .A(n35), .B(n4517), .Z(n4519) );
  XOR U4786 ( .A(b[9]), .B(a[58]), .Z(n4594) );
  NAND U4787 ( .A(n19598), .B(n4594), .Z(n4518) );
  NAND U4788 ( .A(n4519), .B(n4518), .Z(n4597) );
  XOR U4789 ( .A(n4598), .B(n4597), .Z(n4600) );
  XOR U4790 ( .A(n4599), .B(n4600), .Z(n4610) );
  NANDN U4791 ( .A(n4521), .B(n4520), .Z(n4525) );
  OR U4792 ( .A(n4523), .B(n4522), .Z(n4524) );
  AND U4793 ( .A(n4525), .B(n4524), .Z(n4609) );
  XNOR U4794 ( .A(n4610), .B(n4609), .Z(n4611) );
  NANDN U4795 ( .A(n4527), .B(n4526), .Z(n4531) );
  NANDN U4796 ( .A(n4529), .B(n4528), .Z(n4530) );
  NAND U4797 ( .A(n4531), .B(n4530), .Z(n4612) );
  XNOR U4798 ( .A(n4611), .B(n4612), .Z(n4557) );
  XOR U4799 ( .A(n4558), .B(n4557), .Z(n4616) );
  NANDN U4800 ( .A(n4533), .B(n4532), .Z(n4537) );
  NANDN U4801 ( .A(n4535), .B(n4534), .Z(n4536) );
  AND U4802 ( .A(n4537), .B(n4536), .Z(n4615) );
  XNOR U4803 ( .A(n4616), .B(n4615), .Z(n4617) );
  XOR U4804 ( .A(n4618), .B(n4617), .Z(n4550) );
  NANDN U4805 ( .A(n4539), .B(n4538), .Z(n4543) );
  NAND U4806 ( .A(n4541), .B(n4540), .Z(n4542) );
  AND U4807 ( .A(n4543), .B(n4542), .Z(n4549) );
  XNOR U4808 ( .A(n4550), .B(n4549), .Z(n4551) );
  XNOR U4809 ( .A(n4552), .B(n4551), .Z(n4621) );
  XNOR U4810 ( .A(sreg[306]), .B(n4621), .Z(n4623) );
  NANDN U4811 ( .A(sreg[305]), .B(n4544), .Z(n4548) );
  NAND U4812 ( .A(n4546), .B(n4545), .Z(n4547) );
  NAND U4813 ( .A(n4548), .B(n4547), .Z(n4622) );
  XNOR U4814 ( .A(n4623), .B(n4622), .Z(c[306]) );
  NANDN U4815 ( .A(n4550), .B(n4549), .Z(n4554) );
  NANDN U4816 ( .A(n4552), .B(n4551), .Z(n4553) );
  AND U4817 ( .A(n4554), .B(n4553), .Z(n4629) );
  NANDN U4818 ( .A(n4556), .B(n4555), .Z(n4560) );
  NAND U4819 ( .A(n4558), .B(n4557), .Z(n4559) );
  AND U4820 ( .A(n4560), .B(n4559), .Z(n4695) );
  NANDN U4821 ( .A(n4562), .B(n4561), .Z(n4566) );
  NANDN U4822 ( .A(n4564), .B(n4563), .Z(n4565) );
  AND U4823 ( .A(n4566), .B(n4565), .Z(n4661) );
  NAND U4824 ( .A(n19808), .B(n4567), .Z(n4569) );
  XOR U4825 ( .A(b[13]), .B(a[55]), .Z(n4647) );
  NAND U4826 ( .A(n19768), .B(n4647), .Z(n4568) );
  AND U4827 ( .A(n4569), .B(n4568), .Z(n4639) );
  AND U4828 ( .A(b[15]), .B(a[51]), .Z(n4638) );
  XNOR U4829 ( .A(n4639), .B(n4638), .Z(n4640) );
  NAND U4830 ( .A(b[0]), .B(a[67]), .Z(n4570) );
  XNOR U4831 ( .A(b[1]), .B(n4570), .Z(n4572) );
  NANDN U4832 ( .A(b[0]), .B(a[66]), .Z(n4571) );
  NAND U4833 ( .A(n4572), .B(n4571), .Z(n4641) );
  XNOR U4834 ( .A(n4640), .B(n4641), .Z(n4659) );
  NAND U4835 ( .A(n33), .B(n4573), .Z(n4575) );
  XOR U4836 ( .A(b[5]), .B(a[63]), .Z(n4650) );
  NAND U4837 ( .A(n19342), .B(n4650), .Z(n4574) );
  AND U4838 ( .A(n4575), .B(n4574), .Z(n4683) );
  NAND U4839 ( .A(n34), .B(n4576), .Z(n4578) );
  XOR U4840 ( .A(b[7]), .B(a[61]), .Z(n4653) );
  NAND U4841 ( .A(n19486), .B(n4653), .Z(n4577) );
  AND U4842 ( .A(n4578), .B(n4577), .Z(n4681) );
  NAND U4843 ( .A(n31), .B(n4579), .Z(n4581) );
  XOR U4844 ( .A(b[3]), .B(a[65]), .Z(n4656) );
  NAND U4845 ( .A(n32), .B(n4656), .Z(n4580) );
  NAND U4846 ( .A(n4581), .B(n4580), .Z(n4680) );
  XNOR U4847 ( .A(n4681), .B(n4680), .Z(n4682) );
  XOR U4848 ( .A(n4683), .B(n4682), .Z(n4660) );
  XOR U4849 ( .A(n4659), .B(n4660), .Z(n4662) );
  XOR U4850 ( .A(n4661), .B(n4662), .Z(n4633) );
  NANDN U4851 ( .A(n4583), .B(n4582), .Z(n4587) );
  OR U4852 ( .A(n4585), .B(n4584), .Z(n4586) );
  AND U4853 ( .A(n4587), .B(n4586), .Z(n4632) );
  XNOR U4854 ( .A(n4633), .B(n4632), .Z(n4635) );
  NAND U4855 ( .A(n4588), .B(n19724), .Z(n4590) );
  XOR U4856 ( .A(b[11]), .B(a[57]), .Z(n4665) );
  NAND U4857 ( .A(n19692), .B(n4665), .Z(n4589) );
  AND U4858 ( .A(n4590), .B(n4589), .Z(n4676) );
  NAND U4859 ( .A(n19838), .B(n4591), .Z(n4593) );
  XOR U4860 ( .A(b[15]), .B(a[53]), .Z(n4668) );
  NAND U4861 ( .A(n19805), .B(n4668), .Z(n4592) );
  AND U4862 ( .A(n4593), .B(n4592), .Z(n4675) );
  NAND U4863 ( .A(n35), .B(n4594), .Z(n4596) );
  XOR U4864 ( .A(b[9]), .B(a[59]), .Z(n4671) );
  NAND U4865 ( .A(n19598), .B(n4671), .Z(n4595) );
  NAND U4866 ( .A(n4596), .B(n4595), .Z(n4674) );
  XOR U4867 ( .A(n4675), .B(n4674), .Z(n4677) );
  XOR U4868 ( .A(n4676), .B(n4677), .Z(n4687) );
  NANDN U4869 ( .A(n4598), .B(n4597), .Z(n4602) );
  OR U4870 ( .A(n4600), .B(n4599), .Z(n4601) );
  AND U4871 ( .A(n4602), .B(n4601), .Z(n4686) );
  XNOR U4872 ( .A(n4687), .B(n4686), .Z(n4688) );
  NANDN U4873 ( .A(n4604), .B(n4603), .Z(n4608) );
  NANDN U4874 ( .A(n4606), .B(n4605), .Z(n4607) );
  NAND U4875 ( .A(n4608), .B(n4607), .Z(n4689) );
  XNOR U4876 ( .A(n4688), .B(n4689), .Z(n4634) );
  XOR U4877 ( .A(n4635), .B(n4634), .Z(n4693) );
  NANDN U4878 ( .A(n4610), .B(n4609), .Z(n4614) );
  NANDN U4879 ( .A(n4612), .B(n4611), .Z(n4613) );
  AND U4880 ( .A(n4614), .B(n4613), .Z(n4692) );
  XNOR U4881 ( .A(n4693), .B(n4692), .Z(n4694) );
  XOR U4882 ( .A(n4695), .B(n4694), .Z(n4627) );
  NANDN U4883 ( .A(n4616), .B(n4615), .Z(n4620) );
  NAND U4884 ( .A(n4618), .B(n4617), .Z(n4619) );
  AND U4885 ( .A(n4620), .B(n4619), .Z(n4626) );
  XNOR U4886 ( .A(n4627), .B(n4626), .Z(n4628) );
  XNOR U4887 ( .A(n4629), .B(n4628), .Z(n4698) );
  XNOR U4888 ( .A(sreg[307]), .B(n4698), .Z(n4700) );
  NANDN U4889 ( .A(sreg[306]), .B(n4621), .Z(n4625) );
  NAND U4890 ( .A(n4623), .B(n4622), .Z(n4624) );
  NAND U4891 ( .A(n4625), .B(n4624), .Z(n4699) );
  XNOR U4892 ( .A(n4700), .B(n4699), .Z(c[307]) );
  NANDN U4893 ( .A(n4627), .B(n4626), .Z(n4631) );
  NANDN U4894 ( .A(n4629), .B(n4628), .Z(n4630) );
  AND U4895 ( .A(n4631), .B(n4630), .Z(n4706) );
  NANDN U4896 ( .A(n4633), .B(n4632), .Z(n4637) );
  NAND U4897 ( .A(n4635), .B(n4634), .Z(n4636) );
  AND U4898 ( .A(n4637), .B(n4636), .Z(n4772) );
  NANDN U4899 ( .A(n4639), .B(n4638), .Z(n4643) );
  NANDN U4900 ( .A(n4641), .B(n4640), .Z(n4642) );
  AND U4901 ( .A(n4643), .B(n4642), .Z(n4738) );
  NAND U4902 ( .A(b[0]), .B(a[68]), .Z(n4644) );
  XNOR U4903 ( .A(b[1]), .B(n4644), .Z(n4646) );
  NANDN U4904 ( .A(b[0]), .B(a[67]), .Z(n4645) );
  NAND U4905 ( .A(n4646), .B(n4645), .Z(n4718) );
  NAND U4906 ( .A(n19808), .B(n4647), .Z(n4649) );
  XOR U4907 ( .A(b[13]), .B(a[56]), .Z(n4724) );
  NAND U4908 ( .A(n19768), .B(n4724), .Z(n4648) );
  AND U4909 ( .A(n4649), .B(n4648), .Z(n4716) );
  AND U4910 ( .A(b[15]), .B(a[52]), .Z(n4715) );
  XNOR U4911 ( .A(n4716), .B(n4715), .Z(n4717) );
  XNOR U4912 ( .A(n4718), .B(n4717), .Z(n4736) );
  NAND U4913 ( .A(n33), .B(n4650), .Z(n4652) );
  XOR U4914 ( .A(b[5]), .B(a[64]), .Z(n4727) );
  NAND U4915 ( .A(n19342), .B(n4727), .Z(n4651) );
  AND U4916 ( .A(n4652), .B(n4651), .Z(n4760) );
  NAND U4917 ( .A(n34), .B(n4653), .Z(n4655) );
  XOR U4918 ( .A(b[7]), .B(a[62]), .Z(n4730) );
  NAND U4919 ( .A(n19486), .B(n4730), .Z(n4654) );
  AND U4920 ( .A(n4655), .B(n4654), .Z(n4758) );
  NAND U4921 ( .A(n31), .B(n4656), .Z(n4658) );
  XOR U4922 ( .A(b[3]), .B(a[66]), .Z(n4733) );
  NAND U4923 ( .A(n32), .B(n4733), .Z(n4657) );
  NAND U4924 ( .A(n4658), .B(n4657), .Z(n4757) );
  XNOR U4925 ( .A(n4758), .B(n4757), .Z(n4759) );
  XOR U4926 ( .A(n4760), .B(n4759), .Z(n4737) );
  XOR U4927 ( .A(n4736), .B(n4737), .Z(n4739) );
  XOR U4928 ( .A(n4738), .B(n4739), .Z(n4710) );
  NANDN U4929 ( .A(n4660), .B(n4659), .Z(n4664) );
  OR U4930 ( .A(n4662), .B(n4661), .Z(n4663) );
  AND U4931 ( .A(n4664), .B(n4663), .Z(n4709) );
  XNOR U4932 ( .A(n4710), .B(n4709), .Z(n4712) );
  NAND U4933 ( .A(n4665), .B(n19724), .Z(n4667) );
  XOR U4934 ( .A(b[11]), .B(a[58]), .Z(n4742) );
  NAND U4935 ( .A(n19692), .B(n4742), .Z(n4666) );
  AND U4936 ( .A(n4667), .B(n4666), .Z(n4753) );
  NAND U4937 ( .A(n19838), .B(n4668), .Z(n4670) );
  XOR U4938 ( .A(b[15]), .B(a[54]), .Z(n4745) );
  NAND U4939 ( .A(n19805), .B(n4745), .Z(n4669) );
  AND U4940 ( .A(n4670), .B(n4669), .Z(n4752) );
  NAND U4941 ( .A(n35), .B(n4671), .Z(n4673) );
  XOR U4942 ( .A(b[9]), .B(a[60]), .Z(n4748) );
  NAND U4943 ( .A(n19598), .B(n4748), .Z(n4672) );
  NAND U4944 ( .A(n4673), .B(n4672), .Z(n4751) );
  XOR U4945 ( .A(n4752), .B(n4751), .Z(n4754) );
  XOR U4946 ( .A(n4753), .B(n4754), .Z(n4764) );
  NANDN U4947 ( .A(n4675), .B(n4674), .Z(n4679) );
  OR U4948 ( .A(n4677), .B(n4676), .Z(n4678) );
  AND U4949 ( .A(n4679), .B(n4678), .Z(n4763) );
  XNOR U4950 ( .A(n4764), .B(n4763), .Z(n4765) );
  NANDN U4951 ( .A(n4681), .B(n4680), .Z(n4685) );
  NANDN U4952 ( .A(n4683), .B(n4682), .Z(n4684) );
  NAND U4953 ( .A(n4685), .B(n4684), .Z(n4766) );
  XNOR U4954 ( .A(n4765), .B(n4766), .Z(n4711) );
  XOR U4955 ( .A(n4712), .B(n4711), .Z(n4770) );
  NANDN U4956 ( .A(n4687), .B(n4686), .Z(n4691) );
  NANDN U4957 ( .A(n4689), .B(n4688), .Z(n4690) );
  AND U4958 ( .A(n4691), .B(n4690), .Z(n4769) );
  XNOR U4959 ( .A(n4770), .B(n4769), .Z(n4771) );
  XOR U4960 ( .A(n4772), .B(n4771), .Z(n4704) );
  NANDN U4961 ( .A(n4693), .B(n4692), .Z(n4697) );
  NAND U4962 ( .A(n4695), .B(n4694), .Z(n4696) );
  AND U4963 ( .A(n4697), .B(n4696), .Z(n4703) );
  XNOR U4964 ( .A(n4704), .B(n4703), .Z(n4705) );
  XNOR U4965 ( .A(n4706), .B(n4705), .Z(n4775) );
  XNOR U4966 ( .A(sreg[308]), .B(n4775), .Z(n4777) );
  NANDN U4967 ( .A(sreg[307]), .B(n4698), .Z(n4702) );
  NAND U4968 ( .A(n4700), .B(n4699), .Z(n4701) );
  NAND U4969 ( .A(n4702), .B(n4701), .Z(n4776) );
  XNOR U4970 ( .A(n4777), .B(n4776), .Z(c[308]) );
  NANDN U4971 ( .A(n4704), .B(n4703), .Z(n4708) );
  NANDN U4972 ( .A(n4706), .B(n4705), .Z(n4707) );
  AND U4973 ( .A(n4708), .B(n4707), .Z(n4783) );
  NANDN U4974 ( .A(n4710), .B(n4709), .Z(n4714) );
  NAND U4975 ( .A(n4712), .B(n4711), .Z(n4713) );
  AND U4976 ( .A(n4714), .B(n4713), .Z(n4849) );
  NANDN U4977 ( .A(n4716), .B(n4715), .Z(n4720) );
  NANDN U4978 ( .A(n4718), .B(n4717), .Z(n4719) );
  AND U4979 ( .A(n4720), .B(n4719), .Z(n4815) );
  NAND U4980 ( .A(b[0]), .B(a[69]), .Z(n4721) );
  XNOR U4981 ( .A(b[1]), .B(n4721), .Z(n4723) );
  NANDN U4982 ( .A(b[0]), .B(a[68]), .Z(n4722) );
  NAND U4983 ( .A(n4723), .B(n4722), .Z(n4795) );
  NAND U4984 ( .A(n19808), .B(n4724), .Z(n4726) );
  XOR U4985 ( .A(b[13]), .B(a[57]), .Z(n4801) );
  NAND U4986 ( .A(n19768), .B(n4801), .Z(n4725) );
  AND U4987 ( .A(n4726), .B(n4725), .Z(n4793) );
  AND U4988 ( .A(b[15]), .B(a[53]), .Z(n4792) );
  XNOR U4989 ( .A(n4793), .B(n4792), .Z(n4794) );
  XNOR U4990 ( .A(n4795), .B(n4794), .Z(n4813) );
  NAND U4991 ( .A(n33), .B(n4727), .Z(n4729) );
  XOR U4992 ( .A(b[5]), .B(a[65]), .Z(n4804) );
  NAND U4993 ( .A(n19342), .B(n4804), .Z(n4728) );
  AND U4994 ( .A(n4729), .B(n4728), .Z(n4837) );
  NAND U4995 ( .A(n34), .B(n4730), .Z(n4732) );
  XOR U4996 ( .A(b[7]), .B(a[63]), .Z(n4807) );
  NAND U4997 ( .A(n19486), .B(n4807), .Z(n4731) );
  AND U4998 ( .A(n4732), .B(n4731), .Z(n4835) );
  NAND U4999 ( .A(n31), .B(n4733), .Z(n4735) );
  XOR U5000 ( .A(b[3]), .B(a[67]), .Z(n4810) );
  NAND U5001 ( .A(n32), .B(n4810), .Z(n4734) );
  NAND U5002 ( .A(n4735), .B(n4734), .Z(n4834) );
  XNOR U5003 ( .A(n4835), .B(n4834), .Z(n4836) );
  XOR U5004 ( .A(n4837), .B(n4836), .Z(n4814) );
  XOR U5005 ( .A(n4813), .B(n4814), .Z(n4816) );
  XOR U5006 ( .A(n4815), .B(n4816), .Z(n4787) );
  NANDN U5007 ( .A(n4737), .B(n4736), .Z(n4741) );
  OR U5008 ( .A(n4739), .B(n4738), .Z(n4740) );
  AND U5009 ( .A(n4741), .B(n4740), .Z(n4786) );
  XNOR U5010 ( .A(n4787), .B(n4786), .Z(n4789) );
  NAND U5011 ( .A(n4742), .B(n19724), .Z(n4744) );
  XOR U5012 ( .A(b[11]), .B(a[59]), .Z(n4819) );
  NAND U5013 ( .A(n19692), .B(n4819), .Z(n4743) );
  AND U5014 ( .A(n4744), .B(n4743), .Z(n4830) );
  NAND U5015 ( .A(n19838), .B(n4745), .Z(n4747) );
  XOR U5016 ( .A(b[15]), .B(a[55]), .Z(n4822) );
  NAND U5017 ( .A(n19805), .B(n4822), .Z(n4746) );
  AND U5018 ( .A(n4747), .B(n4746), .Z(n4829) );
  NAND U5019 ( .A(n35), .B(n4748), .Z(n4750) );
  XOR U5020 ( .A(b[9]), .B(a[61]), .Z(n4825) );
  NAND U5021 ( .A(n19598), .B(n4825), .Z(n4749) );
  NAND U5022 ( .A(n4750), .B(n4749), .Z(n4828) );
  XOR U5023 ( .A(n4829), .B(n4828), .Z(n4831) );
  XOR U5024 ( .A(n4830), .B(n4831), .Z(n4841) );
  NANDN U5025 ( .A(n4752), .B(n4751), .Z(n4756) );
  OR U5026 ( .A(n4754), .B(n4753), .Z(n4755) );
  AND U5027 ( .A(n4756), .B(n4755), .Z(n4840) );
  XNOR U5028 ( .A(n4841), .B(n4840), .Z(n4842) );
  NANDN U5029 ( .A(n4758), .B(n4757), .Z(n4762) );
  NANDN U5030 ( .A(n4760), .B(n4759), .Z(n4761) );
  NAND U5031 ( .A(n4762), .B(n4761), .Z(n4843) );
  XNOR U5032 ( .A(n4842), .B(n4843), .Z(n4788) );
  XOR U5033 ( .A(n4789), .B(n4788), .Z(n4847) );
  NANDN U5034 ( .A(n4764), .B(n4763), .Z(n4768) );
  NANDN U5035 ( .A(n4766), .B(n4765), .Z(n4767) );
  AND U5036 ( .A(n4768), .B(n4767), .Z(n4846) );
  XNOR U5037 ( .A(n4847), .B(n4846), .Z(n4848) );
  XOR U5038 ( .A(n4849), .B(n4848), .Z(n4781) );
  NANDN U5039 ( .A(n4770), .B(n4769), .Z(n4774) );
  NAND U5040 ( .A(n4772), .B(n4771), .Z(n4773) );
  AND U5041 ( .A(n4774), .B(n4773), .Z(n4780) );
  XNOR U5042 ( .A(n4781), .B(n4780), .Z(n4782) );
  XNOR U5043 ( .A(n4783), .B(n4782), .Z(n4852) );
  XNOR U5044 ( .A(sreg[309]), .B(n4852), .Z(n4854) );
  NANDN U5045 ( .A(sreg[308]), .B(n4775), .Z(n4779) );
  NAND U5046 ( .A(n4777), .B(n4776), .Z(n4778) );
  NAND U5047 ( .A(n4779), .B(n4778), .Z(n4853) );
  XNOR U5048 ( .A(n4854), .B(n4853), .Z(c[309]) );
  NANDN U5049 ( .A(n4781), .B(n4780), .Z(n4785) );
  NANDN U5050 ( .A(n4783), .B(n4782), .Z(n4784) );
  AND U5051 ( .A(n4785), .B(n4784), .Z(n4860) );
  NANDN U5052 ( .A(n4787), .B(n4786), .Z(n4791) );
  NAND U5053 ( .A(n4789), .B(n4788), .Z(n4790) );
  AND U5054 ( .A(n4791), .B(n4790), .Z(n4926) );
  NANDN U5055 ( .A(n4793), .B(n4792), .Z(n4797) );
  NANDN U5056 ( .A(n4795), .B(n4794), .Z(n4796) );
  AND U5057 ( .A(n4797), .B(n4796), .Z(n4892) );
  NAND U5058 ( .A(b[0]), .B(a[70]), .Z(n4798) );
  XNOR U5059 ( .A(b[1]), .B(n4798), .Z(n4800) );
  NANDN U5060 ( .A(b[0]), .B(a[69]), .Z(n4799) );
  NAND U5061 ( .A(n4800), .B(n4799), .Z(n4872) );
  NAND U5062 ( .A(n19808), .B(n4801), .Z(n4803) );
  XOR U5063 ( .A(b[13]), .B(a[58]), .Z(n4878) );
  NAND U5064 ( .A(n19768), .B(n4878), .Z(n4802) );
  AND U5065 ( .A(n4803), .B(n4802), .Z(n4870) );
  AND U5066 ( .A(b[15]), .B(a[54]), .Z(n4869) );
  XNOR U5067 ( .A(n4870), .B(n4869), .Z(n4871) );
  XNOR U5068 ( .A(n4872), .B(n4871), .Z(n4890) );
  NAND U5069 ( .A(n33), .B(n4804), .Z(n4806) );
  XOR U5070 ( .A(b[5]), .B(a[66]), .Z(n4881) );
  NAND U5071 ( .A(n19342), .B(n4881), .Z(n4805) );
  AND U5072 ( .A(n4806), .B(n4805), .Z(n4914) );
  NAND U5073 ( .A(n34), .B(n4807), .Z(n4809) );
  XOR U5074 ( .A(b[7]), .B(a[64]), .Z(n4884) );
  NAND U5075 ( .A(n19486), .B(n4884), .Z(n4808) );
  AND U5076 ( .A(n4809), .B(n4808), .Z(n4912) );
  NAND U5077 ( .A(n31), .B(n4810), .Z(n4812) );
  XOR U5078 ( .A(b[3]), .B(a[68]), .Z(n4887) );
  NAND U5079 ( .A(n32), .B(n4887), .Z(n4811) );
  NAND U5080 ( .A(n4812), .B(n4811), .Z(n4911) );
  XNOR U5081 ( .A(n4912), .B(n4911), .Z(n4913) );
  XOR U5082 ( .A(n4914), .B(n4913), .Z(n4891) );
  XOR U5083 ( .A(n4890), .B(n4891), .Z(n4893) );
  XOR U5084 ( .A(n4892), .B(n4893), .Z(n4864) );
  NANDN U5085 ( .A(n4814), .B(n4813), .Z(n4818) );
  OR U5086 ( .A(n4816), .B(n4815), .Z(n4817) );
  AND U5087 ( .A(n4818), .B(n4817), .Z(n4863) );
  XNOR U5088 ( .A(n4864), .B(n4863), .Z(n4866) );
  NAND U5089 ( .A(n4819), .B(n19724), .Z(n4821) );
  XOR U5090 ( .A(b[11]), .B(a[60]), .Z(n4896) );
  NAND U5091 ( .A(n19692), .B(n4896), .Z(n4820) );
  AND U5092 ( .A(n4821), .B(n4820), .Z(n4907) );
  NAND U5093 ( .A(n19838), .B(n4822), .Z(n4824) );
  XOR U5094 ( .A(b[15]), .B(a[56]), .Z(n4899) );
  NAND U5095 ( .A(n19805), .B(n4899), .Z(n4823) );
  AND U5096 ( .A(n4824), .B(n4823), .Z(n4906) );
  NAND U5097 ( .A(n35), .B(n4825), .Z(n4827) );
  XOR U5098 ( .A(b[9]), .B(a[62]), .Z(n4902) );
  NAND U5099 ( .A(n19598), .B(n4902), .Z(n4826) );
  NAND U5100 ( .A(n4827), .B(n4826), .Z(n4905) );
  XOR U5101 ( .A(n4906), .B(n4905), .Z(n4908) );
  XOR U5102 ( .A(n4907), .B(n4908), .Z(n4918) );
  NANDN U5103 ( .A(n4829), .B(n4828), .Z(n4833) );
  OR U5104 ( .A(n4831), .B(n4830), .Z(n4832) );
  AND U5105 ( .A(n4833), .B(n4832), .Z(n4917) );
  XNOR U5106 ( .A(n4918), .B(n4917), .Z(n4919) );
  NANDN U5107 ( .A(n4835), .B(n4834), .Z(n4839) );
  NANDN U5108 ( .A(n4837), .B(n4836), .Z(n4838) );
  NAND U5109 ( .A(n4839), .B(n4838), .Z(n4920) );
  XNOR U5110 ( .A(n4919), .B(n4920), .Z(n4865) );
  XOR U5111 ( .A(n4866), .B(n4865), .Z(n4924) );
  NANDN U5112 ( .A(n4841), .B(n4840), .Z(n4845) );
  NANDN U5113 ( .A(n4843), .B(n4842), .Z(n4844) );
  AND U5114 ( .A(n4845), .B(n4844), .Z(n4923) );
  XNOR U5115 ( .A(n4924), .B(n4923), .Z(n4925) );
  XOR U5116 ( .A(n4926), .B(n4925), .Z(n4858) );
  NANDN U5117 ( .A(n4847), .B(n4846), .Z(n4851) );
  NAND U5118 ( .A(n4849), .B(n4848), .Z(n4850) );
  AND U5119 ( .A(n4851), .B(n4850), .Z(n4857) );
  XNOR U5120 ( .A(n4858), .B(n4857), .Z(n4859) );
  XNOR U5121 ( .A(n4860), .B(n4859), .Z(n4929) );
  XNOR U5122 ( .A(sreg[310]), .B(n4929), .Z(n4931) );
  NANDN U5123 ( .A(sreg[309]), .B(n4852), .Z(n4856) );
  NAND U5124 ( .A(n4854), .B(n4853), .Z(n4855) );
  NAND U5125 ( .A(n4856), .B(n4855), .Z(n4930) );
  XNOR U5126 ( .A(n4931), .B(n4930), .Z(c[310]) );
  NANDN U5127 ( .A(n4858), .B(n4857), .Z(n4862) );
  NANDN U5128 ( .A(n4860), .B(n4859), .Z(n4861) );
  AND U5129 ( .A(n4862), .B(n4861), .Z(n4937) );
  NANDN U5130 ( .A(n4864), .B(n4863), .Z(n4868) );
  NAND U5131 ( .A(n4866), .B(n4865), .Z(n4867) );
  AND U5132 ( .A(n4868), .B(n4867), .Z(n5003) );
  NANDN U5133 ( .A(n4870), .B(n4869), .Z(n4874) );
  NANDN U5134 ( .A(n4872), .B(n4871), .Z(n4873) );
  AND U5135 ( .A(n4874), .B(n4873), .Z(n4969) );
  NAND U5136 ( .A(b[0]), .B(a[71]), .Z(n4875) );
  XNOR U5137 ( .A(b[1]), .B(n4875), .Z(n4877) );
  NANDN U5138 ( .A(b[0]), .B(a[70]), .Z(n4876) );
  NAND U5139 ( .A(n4877), .B(n4876), .Z(n4949) );
  NAND U5140 ( .A(n19808), .B(n4878), .Z(n4880) );
  XOR U5141 ( .A(b[13]), .B(a[59]), .Z(n4955) );
  NAND U5142 ( .A(n19768), .B(n4955), .Z(n4879) );
  AND U5143 ( .A(n4880), .B(n4879), .Z(n4947) );
  AND U5144 ( .A(b[15]), .B(a[55]), .Z(n4946) );
  XNOR U5145 ( .A(n4947), .B(n4946), .Z(n4948) );
  XNOR U5146 ( .A(n4949), .B(n4948), .Z(n4967) );
  NAND U5147 ( .A(n33), .B(n4881), .Z(n4883) );
  XOR U5148 ( .A(b[5]), .B(a[67]), .Z(n4958) );
  NAND U5149 ( .A(n19342), .B(n4958), .Z(n4882) );
  AND U5150 ( .A(n4883), .B(n4882), .Z(n4991) );
  NAND U5151 ( .A(n34), .B(n4884), .Z(n4886) );
  XOR U5152 ( .A(b[7]), .B(a[65]), .Z(n4961) );
  NAND U5153 ( .A(n19486), .B(n4961), .Z(n4885) );
  AND U5154 ( .A(n4886), .B(n4885), .Z(n4989) );
  NAND U5155 ( .A(n31), .B(n4887), .Z(n4889) );
  XOR U5156 ( .A(b[3]), .B(a[69]), .Z(n4964) );
  NAND U5157 ( .A(n32), .B(n4964), .Z(n4888) );
  NAND U5158 ( .A(n4889), .B(n4888), .Z(n4988) );
  XNOR U5159 ( .A(n4989), .B(n4988), .Z(n4990) );
  XOR U5160 ( .A(n4991), .B(n4990), .Z(n4968) );
  XOR U5161 ( .A(n4967), .B(n4968), .Z(n4970) );
  XOR U5162 ( .A(n4969), .B(n4970), .Z(n4941) );
  NANDN U5163 ( .A(n4891), .B(n4890), .Z(n4895) );
  OR U5164 ( .A(n4893), .B(n4892), .Z(n4894) );
  AND U5165 ( .A(n4895), .B(n4894), .Z(n4940) );
  XNOR U5166 ( .A(n4941), .B(n4940), .Z(n4943) );
  NAND U5167 ( .A(n4896), .B(n19724), .Z(n4898) );
  XOR U5168 ( .A(b[11]), .B(a[61]), .Z(n4973) );
  NAND U5169 ( .A(n19692), .B(n4973), .Z(n4897) );
  AND U5170 ( .A(n4898), .B(n4897), .Z(n4984) );
  NAND U5171 ( .A(n19838), .B(n4899), .Z(n4901) );
  XOR U5172 ( .A(b[15]), .B(a[57]), .Z(n4976) );
  NAND U5173 ( .A(n19805), .B(n4976), .Z(n4900) );
  AND U5174 ( .A(n4901), .B(n4900), .Z(n4983) );
  NAND U5175 ( .A(n35), .B(n4902), .Z(n4904) );
  XOR U5176 ( .A(b[9]), .B(a[63]), .Z(n4979) );
  NAND U5177 ( .A(n19598), .B(n4979), .Z(n4903) );
  NAND U5178 ( .A(n4904), .B(n4903), .Z(n4982) );
  XOR U5179 ( .A(n4983), .B(n4982), .Z(n4985) );
  XOR U5180 ( .A(n4984), .B(n4985), .Z(n4995) );
  NANDN U5181 ( .A(n4906), .B(n4905), .Z(n4910) );
  OR U5182 ( .A(n4908), .B(n4907), .Z(n4909) );
  AND U5183 ( .A(n4910), .B(n4909), .Z(n4994) );
  XNOR U5184 ( .A(n4995), .B(n4994), .Z(n4996) );
  NANDN U5185 ( .A(n4912), .B(n4911), .Z(n4916) );
  NANDN U5186 ( .A(n4914), .B(n4913), .Z(n4915) );
  NAND U5187 ( .A(n4916), .B(n4915), .Z(n4997) );
  XNOR U5188 ( .A(n4996), .B(n4997), .Z(n4942) );
  XOR U5189 ( .A(n4943), .B(n4942), .Z(n5001) );
  NANDN U5190 ( .A(n4918), .B(n4917), .Z(n4922) );
  NANDN U5191 ( .A(n4920), .B(n4919), .Z(n4921) );
  AND U5192 ( .A(n4922), .B(n4921), .Z(n5000) );
  XNOR U5193 ( .A(n5001), .B(n5000), .Z(n5002) );
  XOR U5194 ( .A(n5003), .B(n5002), .Z(n4935) );
  NANDN U5195 ( .A(n4924), .B(n4923), .Z(n4928) );
  NAND U5196 ( .A(n4926), .B(n4925), .Z(n4927) );
  AND U5197 ( .A(n4928), .B(n4927), .Z(n4934) );
  XNOR U5198 ( .A(n4935), .B(n4934), .Z(n4936) );
  XNOR U5199 ( .A(n4937), .B(n4936), .Z(n5006) );
  XNOR U5200 ( .A(sreg[311]), .B(n5006), .Z(n5008) );
  NANDN U5201 ( .A(sreg[310]), .B(n4929), .Z(n4933) );
  NAND U5202 ( .A(n4931), .B(n4930), .Z(n4932) );
  NAND U5203 ( .A(n4933), .B(n4932), .Z(n5007) );
  XNOR U5204 ( .A(n5008), .B(n5007), .Z(c[311]) );
  NANDN U5205 ( .A(n4935), .B(n4934), .Z(n4939) );
  NANDN U5206 ( .A(n4937), .B(n4936), .Z(n4938) );
  AND U5207 ( .A(n4939), .B(n4938), .Z(n5014) );
  NANDN U5208 ( .A(n4941), .B(n4940), .Z(n4945) );
  NAND U5209 ( .A(n4943), .B(n4942), .Z(n4944) );
  AND U5210 ( .A(n4945), .B(n4944), .Z(n5080) );
  NANDN U5211 ( .A(n4947), .B(n4946), .Z(n4951) );
  NANDN U5212 ( .A(n4949), .B(n4948), .Z(n4950) );
  AND U5213 ( .A(n4951), .B(n4950), .Z(n5067) );
  NAND U5214 ( .A(b[0]), .B(a[72]), .Z(n4952) );
  XNOR U5215 ( .A(b[1]), .B(n4952), .Z(n4954) );
  NANDN U5216 ( .A(b[0]), .B(a[71]), .Z(n4953) );
  NAND U5217 ( .A(n4954), .B(n4953), .Z(n5047) );
  NAND U5218 ( .A(n19808), .B(n4955), .Z(n4957) );
  XOR U5219 ( .A(b[13]), .B(a[60]), .Z(n5053) );
  NAND U5220 ( .A(n19768), .B(n5053), .Z(n4956) );
  AND U5221 ( .A(n4957), .B(n4956), .Z(n5045) );
  AND U5222 ( .A(b[15]), .B(a[56]), .Z(n5044) );
  XNOR U5223 ( .A(n5045), .B(n5044), .Z(n5046) );
  XNOR U5224 ( .A(n5047), .B(n5046), .Z(n5065) );
  NAND U5225 ( .A(n33), .B(n4958), .Z(n4960) );
  XOR U5226 ( .A(b[5]), .B(a[68]), .Z(n5056) );
  NAND U5227 ( .A(n19342), .B(n5056), .Z(n4959) );
  AND U5228 ( .A(n4960), .B(n4959), .Z(n5041) );
  NAND U5229 ( .A(n34), .B(n4961), .Z(n4963) );
  XOR U5230 ( .A(b[7]), .B(a[66]), .Z(n5059) );
  NAND U5231 ( .A(n19486), .B(n5059), .Z(n4962) );
  AND U5232 ( .A(n4963), .B(n4962), .Z(n5039) );
  NAND U5233 ( .A(n31), .B(n4964), .Z(n4966) );
  XOR U5234 ( .A(b[3]), .B(a[70]), .Z(n5062) );
  NAND U5235 ( .A(n32), .B(n5062), .Z(n4965) );
  NAND U5236 ( .A(n4966), .B(n4965), .Z(n5038) );
  XNOR U5237 ( .A(n5039), .B(n5038), .Z(n5040) );
  XOR U5238 ( .A(n5041), .B(n5040), .Z(n5066) );
  XOR U5239 ( .A(n5065), .B(n5066), .Z(n5068) );
  XOR U5240 ( .A(n5067), .B(n5068), .Z(n5018) );
  NANDN U5241 ( .A(n4968), .B(n4967), .Z(n4972) );
  OR U5242 ( .A(n4970), .B(n4969), .Z(n4971) );
  AND U5243 ( .A(n4972), .B(n4971), .Z(n5017) );
  XNOR U5244 ( .A(n5018), .B(n5017), .Z(n5020) );
  NAND U5245 ( .A(n4973), .B(n19724), .Z(n4975) );
  XOR U5246 ( .A(b[11]), .B(a[62]), .Z(n5023) );
  NAND U5247 ( .A(n19692), .B(n5023), .Z(n4974) );
  AND U5248 ( .A(n4975), .B(n4974), .Z(n5034) );
  NAND U5249 ( .A(n19838), .B(n4976), .Z(n4978) );
  XOR U5250 ( .A(b[15]), .B(a[58]), .Z(n5026) );
  NAND U5251 ( .A(n19805), .B(n5026), .Z(n4977) );
  AND U5252 ( .A(n4978), .B(n4977), .Z(n5033) );
  NAND U5253 ( .A(n35), .B(n4979), .Z(n4981) );
  XOR U5254 ( .A(b[9]), .B(a[64]), .Z(n5029) );
  NAND U5255 ( .A(n19598), .B(n5029), .Z(n4980) );
  NAND U5256 ( .A(n4981), .B(n4980), .Z(n5032) );
  XOR U5257 ( .A(n5033), .B(n5032), .Z(n5035) );
  XOR U5258 ( .A(n5034), .B(n5035), .Z(n5072) );
  NANDN U5259 ( .A(n4983), .B(n4982), .Z(n4987) );
  OR U5260 ( .A(n4985), .B(n4984), .Z(n4986) );
  AND U5261 ( .A(n4987), .B(n4986), .Z(n5071) );
  XNOR U5262 ( .A(n5072), .B(n5071), .Z(n5073) );
  NANDN U5263 ( .A(n4989), .B(n4988), .Z(n4993) );
  NANDN U5264 ( .A(n4991), .B(n4990), .Z(n4992) );
  NAND U5265 ( .A(n4993), .B(n4992), .Z(n5074) );
  XNOR U5266 ( .A(n5073), .B(n5074), .Z(n5019) );
  XOR U5267 ( .A(n5020), .B(n5019), .Z(n5078) );
  NANDN U5268 ( .A(n4995), .B(n4994), .Z(n4999) );
  NANDN U5269 ( .A(n4997), .B(n4996), .Z(n4998) );
  AND U5270 ( .A(n4999), .B(n4998), .Z(n5077) );
  XNOR U5271 ( .A(n5078), .B(n5077), .Z(n5079) );
  XOR U5272 ( .A(n5080), .B(n5079), .Z(n5012) );
  NANDN U5273 ( .A(n5001), .B(n5000), .Z(n5005) );
  NAND U5274 ( .A(n5003), .B(n5002), .Z(n5004) );
  AND U5275 ( .A(n5005), .B(n5004), .Z(n5011) );
  XNOR U5276 ( .A(n5012), .B(n5011), .Z(n5013) );
  XNOR U5277 ( .A(n5014), .B(n5013), .Z(n5083) );
  XNOR U5278 ( .A(sreg[312]), .B(n5083), .Z(n5085) );
  NANDN U5279 ( .A(sreg[311]), .B(n5006), .Z(n5010) );
  NAND U5280 ( .A(n5008), .B(n5007), .Z(n5009) );
  NAND U5281 ( .A(n5010), .B(n5009), .Z(n5084) );
  XNOR U5282 ( .A(n5085), .B(n5084), .Z(c[312]) );
  NANDN U5283 ( .A(n5012), .B(n5011), .Z(n5016) );
  NANDN U5284 ( .A(n5014), .B(n5013), .Z(n5015) );
  AND U5285 ( .A(n5016), .B(n5015), .Z(n5091) );
  NANDN U5286 ( .A(n5018), .B(n5017), .Z(n5022) );
  NAND U5287 ( .A(n5020), .B(n5019), .Z(n5021) );
  AND U5288 ( .A(n5022), .B(n5021), .Z(n5157) );
  NAND U5289 ( .A(n5023), .B(n19724), .Z(n5025) );
  XOR U5290 ( .A(b[11]), .B(a[63]), .Z(n5127) );
  NAND U5291 ( .A(n19692), .B(n5127), .Z(n5024) );
  AND U5292 ( .A(n5025), .B(n5024), .Z(n5138) );
  NAND U5293 ( .A(n19838), .B(n5026), .Z(n5028) );
  XOR U5294 ( .A(b[15]), .B(a[59]), .Z(n5130) );
  NAND U5295 ( .A(n19805), .B(n5130), .Z(n5027) );
  AND U5296 ( .A(n5028), .B(n5027), .Z(n5137) );
  NAND U5297 ( .A(n35), .B(n5029), .Z(n5031) );
  XOR U5298 ( .A(b[9]), .B(a[65]), .Z(n5133) );
  NAND U5299 ( .A(n19598), .B(n5133), .Z(n5030) );
  NAND U5300 ( .A(n5031), .B(n5030), .Z(n5136) );
  XOR U5301 ( .A(n5137), .B(n5136), .Z(n5139) );
  XOR U5302 ( .A(n5138), .B(n5139), .Z(n5149) );
  NANDN U5303 ( .A(n5033), .B(n5032), .Z(n5037) );
  OR U5304 ( .A(n5035), .B(n5034), .Z(n5036) );
  AND U5305 ( .A(n5037), .B(n5036), .Z(n5148) );
  XNOR U5306 ( .A(n5149), .B(n5148), .Z(n5150) );
  NANDN U5307 ( .A(n5039), .B(n5038), .Z(n5043) );
  NANDN U5308 ( .A(n5041), .B(n5040), .Z(n5042) );
  NAND U5309 ( .A(n5043), .B(n5042), .Z(n5151) );
  XNOR U5310 ( .A(n5150), .B(n5151), .Z(n5097) );
  NANDN U5311 ( .A(n5045), .B(n5044), .Z(n5049) );
  NANDN U5312 ( .A(n5047), .B(n5046), .Z(n5048) );
  AND U5313 ( .A(n5049), .B(n5048), .Z(n5123) );
  AND U5314 ( .A(b[0]), .B(a[73]), .Z(n5050) );
  XOR U5315 ( .A(b[1]), .B(n5050), .Z(n5052) );
  NANDN U5316 ( .A(b[0]), .B(a[72]), .Z(n5051) );
  AND U5317 ( .A(n5052), .B(n5051), .Z(n5102) );
  NAND U5318 ( .A(n19808), .B(n5053), .Z(n5055) );
  XOR U5319 ( .A(b[13]), .B(a[61]), .Z(n5109) );
  NAND U5320 ( .A(n19768), .B(n5109), .Z(n5054) );
  AND U5321 ( .A(n5055), .B(n5054), .Z(n5101) );
  AND U5322 ( .A(b[15]), .B(a[57]), .Z(n5100) );
  XOR U5323 ( .A(n5101), .B(n5100), .Z(n5103) );
  XNOR U5324 ( .A(n5102), .B(n5103), .Z(n5121) );
  NAND U5325 ( .A(n33), .B(n5056), .Z(n5058) );
  XOR U5326 ( .A(b[5]), .B(a[69]), .Z(n5112) );
  NAND U5327 ( .A(n19342), .B(n5112), .Z(n5057) );
  AND U5328 ( .A(n5058), .B(n5057), .Z(n5145) );
  NAND U5329 ( .A(n34), .B(n5059), .Z(n5061) );
  XOR U5330 ( .A(b[7]), .B(a[67]), .Z(n5115) );
  NAND U5331 ( .A(n19486), .B(n5115), .Z(n5060) );
  AND U5332 ( .A(n5061), .B(n5060), .Z(n5143) );
  NAND U5333 ( .A(n31), .B(n5062), .Z(n5064) );
  XOR U5334 ( .A(b[3]), .B(a[71]), .Z(n5118) );
  NAND U5335 ( .A(n32), .B(n5118), .Z(n5063) );
  NAND U5336 ( .A(n5064), .B(n5063), .Z(n5142) );
  XNOR U5337 ( .A(n5143), .B(n5142), .Z(n5144) );
  XOR U5338 ( .A(n5145), .B(n5144), .Z(n5122) );
  XOR U5339 ( .A(n5121), .B(n5122), .Z(n5124) );
  XOR U5340 ( .A(n5123), .B(n5124), .Z(n5095) );
  NANDN U5341 ( .A(n5066), .B(n5065), .Z(n5070) );
  OR U5342 ( .A(n5068), .B(n5067), .Z(n5069) );
  AND U5343 ( .A(n5070), .B(n5069), .Z(n5094) );
  XNOR U5344 ( .A(n5095), .B(n5094), .Z(n5096) );
  XOR U5345 ( .A(n5097), .B(n5096), .Z(n5155) );
  NANDN U5346 ( .A(n5072), .B(n5071), .Z(n5076) );
  NANDN U5347 ( .A(n5074), .B(n5073), .Z(n5075) );
  AND U5348 ( .A(n5076), .B(n5075), .Z(n5154) );
  XNOR U5349 ( .A(n5155), .B(n5154), .Z(n5156) );
  XOR U5350 ( .A(n5157), .B(n5156), .Z(n5089) );
  NANDN U5351 ( .A(n5078), .B(n5077), .Z(n5082) );
  NAND U5352 ( .A(n5080), .B(n5079), .Z(n5081) );
  AND U5353 ( .A(n5082), .B(n5081), .Z(n5088) );
  XNOR U5354 ( .A(n5089), .B(n5088), .Z(n5090) );
  XNOR U5355 ( .A(n5091), .B(n5090), .Z(n5160) );
  XNOR U5356 ( .A(sreg[313]), .B(n5160), .Z(n5162) );
  NANDN U5357 ( .A(sreg[312]), .B(n5083), .Z(n5087) );
  NAND U5358 ( .A(n5085), .B(n5084), .Z(n5086) );
  NAND U5359 ( .A(n5087), .B(n5086), .Z(n5161) );
  XNOR U5360 ( .A(n5162), .B(n5161), .Z(c[313]) );
  NANDN U5361 ( .A(n5089), .B(n5088), .Z(n5093) );
  NANDN U5362 ( .A(n5091), .B(n5090), .Z(n5092) );
  AND U5363 ( .A(n5093), .B(n5092), .Z(n5168) );
  NANDN U5364 ( .A(n5095), .B(n5094), .Z(n5099) );
  NAND U5365 ( .A(n5097), .B(n5096), .Z(n5098) );
  AND U5366 ( .A(n5099), .B(n5098), .Z(n5234) );
  NANDN U5367 ( .A(n5101), .B(n5100), .Z(n5105) );
  NANDN U5368 ( .A(n5103), .B(n5102), .Z(n5104) );
  AND U5369 ( .A(n5105), .B(n5104), .Z(n5200) );
  NAND U5370 ( .A(b[0]), .B(a[74]), .Z(n5106) );
  XNOR U5371 ( .A(b[1]), .B(n5106), .Z(n5108) );
  NANDN U5372 ( .A(b[0]), .B(a[73]), .Z(n5107) );
  NAND U5373 ( .A(n5108), .B(n5107), .Z(n5180) );
  NAND U5374 ( .A(n19808), .B(n5109), .Z(n5111) );
  XOR U5375 ( .A(b[13]), .B(a[62]), .Z(n5186) );
  NAND U5376 ( .A(n19768), .B(n5186), .Z(n5110) );
  AND U5377 ( .A(n5111), .B(n5110), .Z(n5178) );
  AND U5378 ( .A(b[15]), .B(a[58]), .Z(n5177) );
  XNOR U5379 ( .A(n5178), .B(n5177), .Z(n5179) );
  XNOR U5380 ( .A(n5180), .B(n5179), .Z(n5198) );
  NAND U5381 ( .A(n33), .B(n5112), .Z(n5114) );
  XOR U5382 ( .A(b[5]), .B(a[70]), .Z(n5189) );
  NAND U5383 ( .A(n19342), .B(n5189), .Z(n5113) );
  AND U5384 ( .A(n5114), .B(n5113), .Z(n5222) );
  NAND U5385 ( .A(n34), .B(n5115), .Z(n5117) );
  XOR U5386 ( .A(b[7]), .B(a[68]), .Z(n5192) );
  NAND U5387 ( .A(n19486), .B(n5192), .Z(n5116) );
  AND U5388 ( .A(n5117), .B(n5116), .Z(n5220) );
  NAND U5389 ( .A(n31), .B(n5118), .Z(n5120) );
  XOR U5390 ( .A(b[3]), .B(a[72]), .Z(n5195) );
  NAND U5391 ( .A(n32), .B(n5195), .Z(n5119) );
  NAND U5392 ( .A(n5120), .B(n5119), .Z(n5219) );
  XNOR U5393 ( .A(n5220), .B(n5219), .Z(n5221) );
  XOR U5394 ( .A(n5222), .B(n5221), .Z(n5199) );
  XOR U5395 ( .A(n5198), .B(n5199), .Z(n5201) );
  XOR U5396 ( .A(n5200), .B(n5201), .Z(n5172) );
  NANDN U5397 ( .A(n5122), .B(n5121), .Z(n5126) );
  OR U5398 ( .A(n5124), .B(n5123), .Z(n5125) );
  AND U5399 ( .A(n5126), .B(n5125), .Z(n5171) );
  XNOR U5400 ( .A(n5172), .B(n5171), .Z(n5174) );
  NAND U5401 ( .A(n5127), .B(n19724), .Z(n5129) );
  XOR U5402 ( .A(b[11]), .B(a[64]), .Z(n5204) );
  NAND U5403 ( .A(n19692), .B(n5204), .Z(n5128) );
  AND U5404 ( .A(n5129), .B(n5128), .Z(n5215) );
  NAND U5405 ( .A(n19838), .B(n5130), .Z(n5132) );
  XOR U5406 ( .A(b[15]), .B(a[60]), .Z(n5207) );
  NAND U5407 ( .A(n19805), .B(n5207), .Z(n5131) );
  AND U5408 ( .A(n5132), .B(n5131), .Z(n5214) );
  NAND U5409 ( .A(n35), .B(n5133), .Z(n5135) );
  XOR U5410 ( .A(b[9]), .B(a[66]), .Z(n5210) );
  NAND U5411 ( .A(n19598), .B(n5210), .Z(n5134) );
  NAND U5412 ( .A(n5135), .B(n5134), .Z(n5213) );
  XOR U5413 ( .A(n5214), .B(n5213), .Z(n5216) );
  XOR U5414 ( .A(n5215), .B(n5216), .Z(n5226) );
  NANDN U5415 ( .A(n5137), .B(n5136), .Z(n5141) );
  OR U5416 ( .A(n5139), .B(n5138), .Z(n5140) );
  AND U5417 ( .A(n5141), .B(n5140), .Z(n5225) );
  XNOR U5418 ( .A(n5226), .B(n5225), .Z(n5227) );
  NANDN U5419 ( .A(n5143), .B(n5142), .Z(n5147) );
  NANDN U5420 ( .A(n5145), .B(n5144), .Z(n5146) );
  NAND U5421 ( .A(n5147), .B(n5146), .Z(n5228) );
  XNOR U5422 ( .A(n5227), .B(n5228), .Z(n5173) );
  XOR U5423 ( .A(n5174), .B(n5173), .Z(n5232) );
  NANDN U5424 ( .A(n5149), .B(n5148), .Z(n5153) );
  NANDN U5425 ( .A(n5151), .B(n5150), .Z(n5152) );
  AND U5426 ( .A(n5153), .B(n5152), .Z(n5231) );
  XNOR U5427 ( .A(n5232), .B(n5231), .Z(n5233) );
  XOR U5428 ( .A(n5234), .B(n5233), .Z(n5166) );
  NANDN U5429 ( .A(n5155), .B(n5154), .Z(n5159) );
  NAND U5430 ( .A(n5157), .B(n5156), .Z(n5158) );
  AND U5431 ( .A(n5159), .B(n5158), .Z(n5165) );
  XNOR U5432 ( .A(n5166), .B(n5165), .Z(n5167) );
  XNOR U5433 ( .A(n5168), .B(n5167), .Z(n5237) );
  XNOR U5434 ( .A(sreg[314]), .B(n5237), .Z(n5239) );
  NANDN U5435 ( .A(sreg[313]), .B(n5160), .Z(n5164) );
  NAND U5436 ( .A(n5162), .B(n5161), .Z(n5163) );
  NAND U5437 ( .A(n5164), .B(n5163), .Z(n5238) );
  XNOR U5438 ( .A(n5239), .B(n5238), .Z(c[314]) );
  NANDN U5439 ( .A(n5166), .B(n5165), .Z(n5170) );
  NANDN U5440 ( .A(n5168), .B(n5167), .Z(n5169) );
  AND U5441 ( .A(n5170), .B(n5169), .Z(n5245) );
  NANDN U5442 ( .A(n5172), .B(n5171), .Z(n5176) );
  NAND U5443 ( .A(n5174), .B(n5173), .Z(n5175) );
  AND U5444 ( .A(n5176), .B(n5175), .Z(n5311) );
  NANDN U5445 ( .A(n5178), .B(n5177), .Z(n5182) );
  NANDN U5446 ( .A(n5180), .B(n5179), .Z(n5181) );
  AND U5447 ( .A(n5182), .B(n5181), .Z(n5277) );
  NAND U5448 ( .A(b[0]), .B(a[75]), .Z(n5183) );
  XNOR U5449 ( .A(b[1]), .B(n5183), .Z(n5185) );
  NANDN U5450 ( .A(b[0]), .B(a[74]), .Z(n5184) );
  NAND U5451 ( .A(n5185), .B(n5184), .Z(n5257) );
  NAND U5452 ( .A(n19808), .B(n5186), .Z(n5188) );
  XOR U5453 ( .A(b[13]), .B(a[63]), .Z(n5263) );
  NAND U5454 ( .A(n19768), .B(n5263), .Z(n5187) );
  AND U5455 ( .A(n5188), .B(n5187), .Z(n5255) );
  AND U5456 ( .A(b[15]), .B(a[59]), .Z(n5254) );
  XNOR U5457 ( .A(n5255), .B(n5254), .Z(n5256) );
  XNOR U5458 ( .A(n5257), .B(n5256), .Z(n5275) );
  NAND U5459 ( .A(n33), .B(n5189), .Z(n5191) );
  XOR U5460 ( .A(b[5]), .B(a[71]), .Z(n5266) );
  NAND U5461 ( .A(n19342), .B(n5266), .Z(n5190) );
  AND U5462 ( .A(n5191), .B(n5190), .Z(n5299) );
  NAND U5463 ( .A(n34), .B(n5192), .Z(n5194) );
  XOR U5464 ( .A(b[7]), .B(a[69]), .Z(n5269) );
  NAND U5465 ( .A(n19486), .B(n5269), .Z(n5193) );
  AND U5466 ( .A(n5194), .B(n5193), .Z(n5297) );
  NAND U5467 ( .A(n31), .B(n5195), .Z(n5197) );
  XOR U5468 ( .A(b[3]), .B(a[73]), .Z(n5272) );
  NAND U5469 ( .A(n32), .B(n5272), .Z(n5196) );
  NAND U5470 ( .A(n5197), .B(n5196), .Z(n5296) );
  XNOR U5471 ( .A(n5297), .B(n5296), .Z(n5298) );
  XOR U5472 ( .A(n5299), .B(n5298), .Z(n5276) );
  XOR U5473 ( .A(n5275), .B(n5276), .Z(n5278) );
  XOR U5474 ( .A(n5277), .B(n5278), .Z(n5249) );
  NANDN U5475 ( .A(n5199), .B(n5198), .Z(n5203) );
  OR U5476 ( .A(n5201), .B(n5200), .Z(n5202) );
  AND U5477 ( .A(n5203), .B(n5202), .Z(n5248) );
  XNOR U5478 ( .A(n5249), .B(n5248), .Z(n5251) );
  NAND U5479 ( .A(n5204), .B(n19724), .Z(n5206) );
  XOR U5480 ( .A(b[11]), .B(a[65]), .Z(n5281) );
  NAND U5481 ( .A(n19692), .B(n5281), .Z(n5205) );
  AND U5482 ( .A(n5206), .B(n5205), .Z(n5292) );
  NAND U5483 ( .A(n19838), .B(n5207), .Z(n5209) );
  XOR U5484 ( .A(b[15]), .B(a[61]), .Z(n5284) );
  NAND U5485 ( .A(n19805), .B(n5284), .Z(n5208) );
  AND U5486 ( .A(n5209), .B(n5208), .Z(n5291) );
  NAND U5487 ( .A(n35), .B(n5210), .Z(n5212) );
  XOR U5488 ( .A(b[9]), .B(a[67]), .Z(n5287) );
  NAND U5489 ( .A(n19598), .B(n5287), .Z(n5211) );
  NAND U5490 ( .A(n5212), .B(n5211), .Z(n5290) );
  XOR U5491 ( .A(n5291), .B(n5290), .Z(n5293) );
  XOR U5492 ( .A(n5292), .B(n5293), .Z(n5303) );
  NANDN U5493 ( .A(n5214), .B(n5213), .Z(n5218) );
  OR U5494 ( .A(n5216), .B(n5215), .Z(n5217) );
  AND U5495 ( .A(n5218), .B(n5217), .Z(n5302) );
  XNOR U5496 ( .A(n5303), .B(n5302), .Z(n5304) );
  NANDN U5497 ( .A(n5220), .B(n5219), .Z(n5224) );
  NANDN U5498 ( .A(n5222), .B(n5221), .Z(n5223) );
  NAND U5499 ( .A(n5224), .B(n5223), .Z(n5305) );
  XNOR U5500 ( .A(n5304), .B(n5305), .Z(n5250) );
  XOR U5501 ( .A(n5251), .B(n5250), .Z(n5309) );
  NANDN U5502 ( .A(n5226), .B(n5225), .Z(n5230) );
  NANDN U5503 ( .A(n5228), .B(n5227), .Z(n5229) );
  AND U5504 ( .A(n5230), .B(n5229), .Z(n5308) );
  XNOR U5505 ( .A(n5309), .B(n5308), .Z(n5310) );
  XOR U5506 ( .A(n5311), .B(n5310), .Z(n5243) );
  NANDN U5507 ( .A(n5232), .B(n5231), .Z(n5236) );
  NAND U5508 ( .A(n5234), .B(n5233), .Z(n5235) );
  AND U5509 ( .A(n5236), .B(n5235), .Z(n5242) );
  XNOR U5510 ( .A(n5243), .B(n5242), .Z(n5244) );
  XNOR U5511 ( .A(n5245), .B(n5244), .Z(n5314) );
  XNOR U5512 ( .A(sreg[315]), .B(n5314), .Z(n5316) );
  NANDN U5513 ( .A(sreg[314]), .B(n5237), .Z(n5241) );
  NAND U5514 ( .A(n5239), .B(n5238), .Z(n5240) );
  NAND U5515 ( .A(n5241), .B(n5240), .Z(n5315) );
  XNOR U5516 ( .A(n5316), .B(n5315), .Z(c[315]) );
  NANDN U5517 ( .A(n5243), .B(n5242), .Z(n5247) );
  NANDN U5518 ( .A(n5245), .B(n5244), .Z(n5246) );
  AND U5519 ( .A(n5247), .B(n5246), .Z(n5322) );
  NANDN U5520 ( .A(n5249), .B(n5248), .Z(n5253) );
  NAND U5521 ( .A(n5251), .B(n5250), .Z(n5252) );
  AND U5522 ( .A(n5253), .B(n5252), .Z(n5388) );
  NANDN U5523 ( .A(n5255), .B(n5254), .Z(n5259) );
  NANDN U5524 ( .A(n5257), .B(n5256), .Z(n5258) );
  AND U5525 ( .A(n5259), .B(n5258), .Z(n5354) );
  NAND U5526 ( .A(b[0]), .B(a[76]), .Z(n5260) );
  XNOR U5527 ( .A(b[1]), .B(n5260), .Z(n5262) );
  NANDN U5528 ( .A(b[0]), .B(a[75]), .Z(n5261) );
  NAND U5529 ( .A(n5262), .B(n5261), .Z(n5334) );
  NAND U5530 ( .A(n19808), .B(n5263), .Z(n5265) );
  XOR U5531 ( .A(b[13]), .B(a[64]), .Z(n5337) );
  NAND U5532 ( .A(n19768), .B(n5337), .Z(n5264) );
  AND U5533 ( .A(n5265), .B(n5264), .Z(n5332) );
  AND U5534 ( .A(b[15]), .B(a[60]), .Z(n5331) );
  XNOR U5535 ( .A(n5332), .B(n5331), .Z(n5333) );
  XNOR U5536 ( .A(n5334), .B(n5333), .Z(n5352) );
  NAND U5537 ( .A(n33), .B(n5266), .Z(n5268) );
  XOR U5538 ( .A(b[5]), .B(a[72]), .Z(n5343) );
  NAND U5539 ( .A(n19342), .B(n5343), .Z(n5267) );
  AND U5540 ( .A(n5268), .B(n5267), .Z(n5376) );
  NAND U5541 ( .A(n34), .B(n5269), .Z(n5271) );
  XOR U5542 ( .A(b[7]), .B(a[70]), .Z(n5346) );
  NAND U5543 ( .A(n19486), .B(n5346), .Z(n5270) );
  AND U5544 ( .A(n5271), .B(n5270), .Z(n5374) );
  NAND U5545 ( .A(n31), .B(n5272), .Z(n5274) );
  XOR U5546 ( .A(b[3]), .B(a[74]), .Z(n5349) );
  NAND U5547 ( .A(n32), .B(n5349), .Z(n5273) );
  NAND U5548 ( .A(n5274), .B(n5273), .Z(n5373) );
  XNOR U5549 ( .A(n5374), .B(n5373), .Z(n5375) );
  XOR U5550 ( .A(n5376), .B(n5375), .Z(n5353) );
  XOR U5551 ( .A(n5352), .B(n5353), .Z(n5355) );
  XOR U5552 ( .A(n5354), .B(n5355), .Z(n5326) );
  NANDN U5553 ( .A(n5276), .B(n5275), .Z(n5280) );
  OR U5554 ( .A(n5278), .B(n5277), .Z(n5279) );
  AND U5555 ( .A(n5280), .B(n5279), .Z(n5325) );
  XNOR U5556 ( .A(n5326), .B(n5325), .Z(n5328) );
  NAND U5557 ( .A(n5281), .B(n19724), .Z(n5283) );
  XOR U5558 ( .A(b[11]), .B(a[66]), .Z(n5358) );
  NAND U5559 ( .A(n19692), .B(n5358), .Z(n5282) );
  AND U5560 ( .A(n5283), .B(n5282), .Z(n5369) );
  NAND U5561 ( .A(n19838), .B(n5284), .Z(n5286) );
  XOR U5562 ( .A(b[15]), .B(a[62]), .Z(n5361) );
  NAND U5563 ( .A(n19805), .B(n5361), .Z(n5285) );
  AND U5564 ( .A(n5286), .B(n5285), .Z(n5368) );
  NAND U5565 ( .A(n35), .B(n5287), .Z(n5289) );
  XOR U5566 ( .A(b[9]), .B(a[68]), .Z(n5364) );
  NAND U5567 ( .A(n19598), .B(n5364), .Z(n5288) );
  NAND U5568 ( .A(n5289), .B(n5288), .Z(n5367) );
  XOR U5569 ( .A(n5368), .B(n5367), .Z(n5370) );
  XOR U5570 ( .A(n5369), .B(n5370), .Z(n5380) );
  NANDN U5571 ( .A(n5291), .B(n5290), .Z(n5295) );
  OR U5572 ( .A(n5293), .B(n5292), .Z(n5294) );
  AND U5573 ( .A(n5295), .B(n5294), .Z(n5379) );
  XNOR U5574 ( .A(n5380), .B(n5379), .Z(n5381) );
  NANDN U5575 ( .A(n5297), .B(n5296), .Z(n5301) );
  NANDN U5576 ( .A(n5299), .B(n5298), .Z(n5300) );
  NAND U5577 ( .A(n5301), .B(n5300), .Z(n5382) );
  XNOR U5578 ( .A(n5381), .B(n5382), .Z(n5327) );
  XOR U5579 ( .A(n5328), .B(n5327), .Z(n5386) );
  NANDN U5580 ( .A(n5303), .B(n5302), .Z(n5307) );
  NANDN U5581 ( .A(n5305), .B(n5304), .Z(n5306) );
  AND U5582 ( .A(n5307), .B(n5306), .Z(n5385) );
  XNOR U5583 ( .A(n5386), .B(n5385), .Z(n5387) );
  XOR U5584 ( .A(n5388), .B(n5387), .Z(n5320) );
  NANDN U5585 ( .A(n5309), .B(n5308), .Z(n5313) );
  NAND U5586 ( .A(n5311), .B(n5310), .Z(n5312) );
  AND U5587 ( .A(n5313), .B(n5312), .Z(n5319) );
  XNOR U5588 ( .A(n5320), .B(n5319), .Z(n5321) );
  XNOR U5589 ( .A(n5322), .B(n5321), .Z(n5391) );
  XNOR U5590 ( .A(sreg[316]), .B(n5391), .Z(n5393) );
  NANDN U5591 ( .A(sreg[315]), .B(n5314), .Z(n5318) );
  NAND U5592 ( .A(n5316), .B(n5315), .Z(n5317) );
  NAND U5593 ( .A(n5318), .B(n5317), .Z(n5392) );
  XNOR U5594 ( .A(n5393), .B(n5392), .Z(c[316]) );
  NANDN U5595 ( .A(n5320), .B(n5319), .Z(n5324) );
  NANDN U5596 ( .A(n5322), .B(n5321), .Z(n5323) );
  AND U5597 ( .A(n5324), .B(n5323), .Z(n5399) );
  NANDN U5598 ( .A(n5326), .B(n5325), .Z(n5330) );
  NAND U5599 ( .A(n5328), .B(n5327), .Z(n5329) );
  AND U5600 ( .A(n5330), .B(n5329), .Z(n5465) );
  NANDN U5601 ( .A(n5332), .B(n5331), .Z(n5336) );
  NANDN U5602 ( .A(n5334), .B(n5333), .Z(n5335) );
  AND U5603 ( .A(n5336), .B(n5335), .Z(n5431) );
  NAND U5604 ( .A(n19808), .B(n5337), .Z(n5339) );
  XOR U5605 ( .A(b[13]), .B(a[65]), .Z(n5417) );
  NAND U5606 ( .A(n19768), .B(n5417), .Z(n5338) );
  AND U5607 ( .A(n5339), .B(n5338), .Z(n5409) );
  AND U5608 ( .A(b[15]), .B(a[61]), .Z(n5408) );
  XNOR U5609 ( .A(n5409), .B(n5408), .Z(n5410) );
  NAND U5610 ( .A(b[0]), .B(a[77]), .Z(n5340) );
  XNOR U5611 ( .A(b[1]), .B(n5340), .Z(n5342) );
  NANDN U5612 ( .A(b[0]), .B(a[76]), .Z(n5341) );
  NAND U5613 ( .A(n5342), .B(n5341), .Z(n5411) );
  XNOR U5614 ( .A(n5410), .B(n5411), .Z(n5429) );
  NAND U5615 ( .A(n33), .B(n5343), .Z(n5345) );
  XOR U5616 ( .A(b[5]), .B(a[73]), .Z(n5420) );
  NAND U5617 ( .A(n19342), .B(n5420), .Z(n5344) );
  AND U5618 ( .A(n5345), .B(n5344), .Z(n5453) );
  NAND U5619 ( .A(n34), .B(n5346), .Z(n5348) );
  XOR U5620 ( .A(b[7]), .B(a[71]), .Z(n5423) );
  NAND U5621 ( .A(n19486), .B(n5423), .Z(n5347) );
  AND U5622 ( .A(n5348), .B(n5347), .Z(n5451) );
  NAND U5623 ( .A(n31), .B(n5349), .Z(n5351) );
  XOR U5624 ( .A(b[3]), .B(a[75]), .Z(n5426) );
  NAND U5625 ( .A(n32), .B(n5426), .Z(n5350) );
  NAND U5626 ( .A(n5351), .B(n5350), .Z(n5450) );
  XNOR U5627 ( .A(n5451), .B(n5450), .Z(n5452) );
  XOR U5628 ( .A(n5453), .B(n5452), .Z(n5430) );
  XOR U5629 ( .A(n5429), .B(n5430), .Z(n5432) );
  XOR U5630 ( .A(n5431), .B(n5432), .Z(n5403) );
  NANDN U5631 ( .A(n5353), .B(n5352), .Z(n5357) );
  OR U5632 ( .A(n5355), .B(n5354), .Z(n5356) );
  AND U5633 ( .A(n5357), .B(n5356), .Z(n5402) );
  XNOR U5634 ( .A(n5403), .B(n5402), .Z(n5405) );
  NAND U5635 ( .A(n5358), .B(n19724), .Z(n5360) );
  XOR U5636 ( .A(b[11]), .B(a[67]), .Z(n5435) );
  NAND U5637 ( .A(n19692), .B(n5435), .Z(n5359) );
  AND U5638 ( .A(n5360), .B(n5359), .Z(n5446) );
  NAND U5639 ( .A(n19838), .B(n5361), .Z(n5363) );
  XOR U5640 ( .A(b[15]), .B(a[63]), .Z(n5438) );
  NAND U5641 ( .A(n19805), .B(n5438), .Z(n5362) );
  AND U5642 ( .A(n5363), .B(n5362), .Z(n5445) );
  NAND U5643 ( .A(n35), .B(n5364), .Z(n5366) );
  XOR U5644 ( .A(b[9]), .B(a[69]), .Z(n5441) );
  NAND U5645 ( .A(n19598), .B(n5441), .Z(n5365) );
  NAND U5646 ( .A(n5366), .B(n5365), .Z(n5444) );
  XOR U5647 ( .A(n5445), .B(n5444), .Z(n5447) );
  XOR U5648 ( .A(n5446), .B(n5447), .Z(n5457) );
  NANDN U5649 ( .A(n5368), .B(n5367), .Z(n5372) );
  OR U5650 ( .A(n5370), .B(n5369), .Z(n5371) );
  AND U5651 ( .A(n5372), .B(n5371), .Z(n5456) );
  XNOR U5652 ( .A(n5457), .B(n5456), .Z(n5458) );
  NANDN U5653 ( .A(n5374), .B(n5373), .Z(n5378) );
  NANDN U5654 ( .A(n5376), .B(n5375), .Z(n5377) );
  NAND U5655 ( .A(n5378), .B(n5377), .Z(n5459) );
  XNOR U5656 ( .A(n5458), .B(n5459), .Z(n5404) );
  XOR U5657 ( .A(n5405), .B(n5404), .Z(n5463) );
  NANDN U5658 ( .A(n5380), .B(n5379), .Z(n5384) );
  NANDN U5659 ( .A(n5382), .B(n5381), .Z(n5383) );
  AND U5660 ( .A(n5384), .B(n5383), .Z(n5462) );
  XNOR U5661 ( .A(n5463), .B(n5462), .Z(n5464) );
  XOR U5662 ( .A(n5465), .B(n5464), .Z(n5397) );
  NANDN U5663 ( .A(n5386), .B(n5385), .Z(n5390) );
  NAND U5664 ( .A(n5388), .B(n5387), .Z(n5389) );
  AND U5665 ( .A(n5390), .B(n5389), .Z(n5396) );
  XNOR U5666 ( .A(n5397), .B(n5396), .Z(n5398) );
  XNOR U5667 ( .A(n5399), .B(n5398), .Z(n5468) );
  XNOR U5668 ( .A(sreg[317]), .B(n5468), .Z(n5470) );
  NANDN U5669 ( .A(sreg[316]), .B(n5391), .Z(n5395) );
  NAND U5670 ( .A(n5393), .B(n5392), .Z(n5394) );
  NAND U5671 ( .A(n5395), .B(n5394), .Z(n5469) );
  XNOR U5672 ( .A(n5470), .B(n5469), .Z(c[317]) );
  NANDN U5673 ( .A(n5397), .B(n5396), .Z(n5401) );
  NANDN U5674 ( .A(n5399), .B(n5398), .Z(n5400) );
  AND U5675 ( .A(n5401), .B(n5400), .Z(n5476) );
  NANDN U5676 ( .A(n5403), .B(n5402), .Z(n5407) );
  NAND U5677 ( .A(n5405), .B(n5404), .Z(n5406) );
  AND U5678 ( .A(n5407), .B(n5406), .Z(n5542) );
  NANDN U5679 ( .A(n5409), .B(n5408), .Z(n5413) );
  NANDN U5680 ( .A(n5411), .B(n5410), .Z(n5412) );
  AND U5681 ( .A(n5413), .B(n5412), .Z(n5508) );
  NAND U5682 ( .A(b[0]), .B(a[78]), .Z(n5414) );
  XNOR U5683 ( .A(b[1]), .B(n5414), .Z(n5416) );
  NANDN U5684 ( .A(b[0]), .B(a[77]), .Z(n5415) );
  NAND U5685 ( .A(n5416), .B(n5415), .Z(n5488) );
  NAND U5686 ( .A(n19808), .B(n5417), .Z(n5419) );
  XOR U5687 ( .A(b[13]), .B(a[66]), .Z(n5494) );
  NAND U5688 ( .A(n19768), .B(n5494), .Z(n5418) );
  AND U5689 ( .A(n5419), .B(n5418), .Z(n5486) );
  AND U5690 ( .A(b[15]), .B(a[62]), .Z(n5485) );
  XNOR U5691 ( .A(n5486), .B(n5485), .Z(n5487) );
  XNOR U5692 ( .A(n5488), .B(n5487), .Z(n5506) );
  NAND U5693 ( .A(n33), .B(n5420), .Z(n5422) );
  XOR U5694 ( .A(b[5]), .B(a[74]), .Z(n5497) );
  NAND U5695 ( .A(n19342), .B(n5497), .Z(n5421) );
  AND U5696 ( .A(n5422), .B(n5421), .Z(n5530) );
  NAND U5697 ( .A(n34), .B(n5423), .Z(n5425) );
  XOR U5698 ( .A(b[7]), .B(a[72]), .Z(n5500) );
  NAND U5699 ( .A(n19486), .B(n5500), .Z(n5424) );
  AND U5700 ( .A(n5425), .B(n5424), .Z(n5528) );
  NAND U5701 ( .A(n31), .B(n5426), .Z(n5428) );
  XOR U5702 ( .A(b[3]), .B(a[76]), .Z(n5503) );
  NAND U5703 ( .A(n32), .B(n5503), .Z(n5427) );
  NAND U5704 ( .A(n5428), .B(n5427), .Z(n5527) );
  XNOR U5705 ( .A(n5528), .B(n5527), .Z(n5529) );
  XOR U5706 ( .A(n5530), .B(n5529), .Z(n5507) );
  XOR U5707 ( .A(n5506), .B(n5507), .Z(n5509) );
  XOR U5708 ( .A(n5508), .B(n5509), .Z(n5480) );
  NANDN U5709 ( .A(n5430), .B(n5429), .Z(n5434) );
  OR U5710 ( .A(n5432), .B(n5431), .Z(n5433) );
  AND U5711 ( .A(n5434), .B(n5433), .Z(n5479) );
  XNOR U5712 ( .A(n5480), .B(n5479), .Z(n5482) );
  NAND U5713 ( .A(n5435), .B(n19724), .Z(n5437) );
  XOR U5714 ( .A(b[11]), .B(a[68]), .Z(n5512) );
  NAND U5715 ( .A(n19692), .B(n5512), .Z(n5436) );
  AND U5716 ( .A(n5437), .B(n5436), .Z(n5523) );
  NAND U5717 ( .A(n19838), .B(n5438), .Z(n5440) );
  XOR U5718 ( .A(b[15]), .B(a[64]), .Z(n5515) );
  NAND U5719 ( .A(n19805), .B(n5515), .Z(n5439) );
  AND U5720 ( .A(n5440), .B(n5439), .Z(n5522) );
  NAND U5721 ( .A(n35), .B(n5441), .Z(n5443) );
  XOR U5722 ( .A(b[9]), .B(a[70]), .Z(n5518) );
  NAND U5723 ( .A(n19598), .B(n5518), .Z(n5442) );
  NAND U5724 ( .A(n5443), .B(n5442), .Z(n5521) );
  XOR U5725 ( .A(n5522), .B(n5521), .Z(n5524) );
  XOR U5726 ( .A(n5523), .B(n5524), .Z(n5534) );
  NANDN U5727 ( .A(n5445), .B(n5444), .Z(n5449) );
  OR U5728 ( .A(n5447), .B(n5446), .Z(n5448) );
  AND U5729 ( .A(n5449), .B(n5448), .Z(n5533) );
  XNOR U5730 ( .A(n5534), .B(n5533), .Z(n5535) );
  NANDN U5731 ( .A(n5451), .B(n5450), .Z(n5455) );
  NANDN U5732 ( .A(n5453), .B(n5452), .Z(n5454) );
  NAND U5733 ( .A(n5455), .B(n5454), .Z(n5536) );
  XNOR U5734 ( .A(n5535), .B(n5536), .Z(n5481) );
  XOR U5735 ( .A(n5482), .B(n5481), .Z(n5540) );
  NANDN U5736 ( .A(n5457), .B(n5456), .Z(n5461) );
  NANDN U5737 ( .A(n5459), .B(n5458), .Z(n5460) );
  AND U5738 ( .A(n5461), .B(n5460), .Z(n5539) );
  XNOR U5739 ( .A(n5540), .B(n5539), .Z(n5541) );
  XOR U5740 ( .A(n5542), .B(n5541), .Z(n5474) );
  NANDN U5741 ( .A(n5463), .B(n5462), .Z(n5467) );
  NAND U5742 ( .A(n5465), .B(n5464), .Z(n5466) );
  AND U5743 ( .A(n5467), .B(n5466), .Z(n5473) );
  XNOR U5744 ( .A(n5474), .B(n5473), .Z(n5475) );
  XNOR U5745 ( .A(n5476), .B(n5475), .Z(n5545) );
  XNOR U5746 ( .A(sreg[318]), .B(n5545), .Z(n5547) );
  NANDN U5747 ( .A(sreg[317]), .B(n5468), .Z(n5472) );
  NAND U5748 ( .A(n5470), .B(n5469), .Z(n5471) );
  NAND U5749 ( .A(n5472), .B(n5471), .Z(n5546) );
  XNOR U5750 ( .A(n5547), .B(n5546), .Z(c[318]) );
  NANDN U5751 ( .A(n5474), .B(n5473), .Z(n5478) );
  NANDN U5752 ( .A(n5476), .B(n5475), .Z(n5477) );
  AND U5753 ( .A(n5478), .B(n5477), .Z(n5553) );
  NANDN U5754 ( .A(n5480), .B(n5479), .Z(n5484) );
  NAND U5755 ( .A(n5482), .B(n5481), .Z(n5483) );
  AND U5756 ( .A(n5484), .B(n5483), .Z(n5619) );
  NANDN U5757 ( .A(n5486), .B(n5485), .Z(n5490) );
  NANDN U5758 ( .A(n5488), .B(n5487), .Z(n5489) );
  AND U5759 ( .A(n5490), .B(n5489), .Z(n5585) );
  NAND U5760 ( .A(b[0]), .B(a[79]), .Z(n5491) );
  XNOR U5761 ( .A(b[1]), .B(n5491), .Z(n5493) );
  NANDN U5762 ( .A(b[0]), .B(a[78]), .Z(n5492) );
  NAND U5763 ( .A(n5493), .B(n5492), .Z(n5565) );
  NAND U5764 ( .A(n19808), .B(n5494), .Z(n5496) );
  XOR U5765 ( .A(b[13]), .B(a[67]), .Z(n5571) );
  NAND U5766 ( .A(n19768), .B(n5571), .Z(n5495) );
  AND U5767 ( .A(n5496), .B(n5495), .Z(n5563) );
  AND U5768 ( .A(b[15]), .B(a[63]), .Z(n5562) );
  XNOR U5769 ( .A(n5563), .B(n5562), .Z(n5564) );
  XNOR U5770 ( .A(n5565), .B(n5564), .Z(n5583) );
  NAND U5771 ( .A(n33), .B(n5497), .Z(n5499) );
  XOR U5772 ( .A(b[5]), .B(a[75]), .Z(n5574) );
  NAND U5773 ( .A(n19342), .B(n5574), .Z(n5498) );
  AND U5774 ( .A(n5499), .B(n5498), .Z(n5607) );
  NAND U5775 ( .A(n34), .B(n5500), .Z(n5502) );
  XOR U5776 ( .A(b[7]), .B(a[73]), .Z(n5577) );
  NAND U5777 ( .A(n19486), .B(n5577), .Z(n5501) );
  AND U5778 ( .A(n5502), .B(n5501), .Z(n5605) );
  NAND U5779 ( .A(n31), .B(n5503), .Z(n5505) );
  XOR U5780 ( .A(b[3]), .B(a[77]), .Z(n5580) );
  NAND U5781 ( .A(n32), .B(n5580), .Z(n5504) );
  NAND U5782 ( .A(n5505), .B(n5504), .Z(n5604) );
  XNOR U5783 ( .A(n5605), .B(n5604), .Z(n5606) );
  XOR U5784 ( .A(n5607), .B(n5606), .Z(n5584) );
  XOR U5785 ( .A(n5583), .B(n5584), .Z(n5586) );
  XOR U5786 ( .A(n5585), .B(n5586), .Z(n5557) );
  NANDN U5787 ( .A(n5507), .B(n5506), .Z(n5511) );
  OR U5788 ( .A(n5509), .B(n5508), .Z(n5510) );
  AND U5789 ( .A(n5511), .B(n5510), .Z(n5556) );
  XNOR U5790 ( .A(n5557), .B(n5556), .Z(n5559) );
  NAND U5791 ( .A(n5512), .B(n19724), .Z(n5514) );
  XOR U5792 ( .A(b[11]), .B(a[69]), .Z(n5589) );
  NAND U5793 ( .A(n19692), .B(n5589), .Z(n5513) );
  AND U5794 ( .A(n5514), .B(n5513), .Z(n5600) );
  NAND U5795 ( .A(n19838), .B(n5515), .Z(n5517) );
  XOR U5796 ( .A(b[15]), .B(a[65]), .Z(n5592) );
  NAND U5797 ( .A(n19805), .B(n5592), .Z(n5516) );
  AND U5798 ( .A(n5517), .B(n5516), .Z(n5599) );
  NAND U5799 ( .A(n35), .B(n5518), .Z(n5520) );
  XOR U5800 ( .A(b[9]), .B(a[71]), .Z(n5595) );
  NAND U5801 ( .A(n19598), .B(n5595), .Z(n5519) );
  NAND U5802 ( .A(n5520), .B(n5519), .Z(n5598) );
  XOR U5803 ( .A(n5599), .B(n5598), .Z(n5601) );
  XOR U5804 ( .A(n5600), .B(n5601), .Z(n5611) );
  NANDN U5805 ( .A(n5522), .B(n5521), .Z(n5526) );
  OR U5806 ( .A(n5524), .B(n5523), .Z(n5525) );
  AND U5807 ( .A(n5526), .B(n5525), .Z(n5610) );
  XNOR U5808 ( .A(n5611), .B(n5610), .Z(n5612) );
  NANDN U5809 ( .A(n5528), .B(n5527), .Z(n5532) );
  NANDN U5810 ( .A(n5530), .B(n5529), .Z(n5531) );
  NAND U5811 ( .A(n5532), .B(n5531), .Z(n5613) );
  XNOR U5812 ( .A(n5612), .B(n5613), .Z(n5558) );
  XOR U5813 ( .A(n5559), .B(n5558), .Z(n5617) );
  NANDN U5814 ( .A(n5534), .B(n5533), .Z(n5538) );
  NANDN U5815 ( .A(n5536), .B(n5535), .Z(n5537) );
  AND U5816 ( .A(n5538), .B(n5537), .Z(n5616) );
  XNOR U5817 ( .A(n5617), .B(n5616), .Z(n5618) );
  XOR U5818 ( .A(n5619), .B(n5618), .Z(n5551) );
  NANDN U5819 ( .A(n5540), .B(n5539), .Z(n5544) );
  NAND U5820 ( .A(n5542), .B(n5541), .Z(n5543) );
  AND U5821 ( .A(n5544), .B(n5543), .Z(n5550) );
  XNOR U5822 ( .A(n5551), .B(n5550), .Z(n5552) );
  XNOR U5823 ( .A(n5553), .B(n5552), .Z(n5622) );
  XNOR U5824 ( .A(sreg[319]), .B(n5622), .Z(n5624) );
  NANDN U5825 ( .A(sreg[318]), .B(n5545), .Z(n5549) );
  NAND U5826 ( .A(n5547), .B(n5546), .Z(n5548) );
  NAND U5827 ( .A(n5549), .B(n5548), .Z(n5623) );
  XNOR U5828 ( .A(n5624), .B(n5623), .Z(c[319]) );
  NANDN U5829 ( .A(n5551), .B(n5550), .Z(n5555) );
  NANDN U5830 ( .A(n5553), .B(n5552), .Z(n5554) );
  AND U5831 ( .A(n5555), .B(n5554), .Z(n5630) );
  NANDN U5832 ( .A(n5557), .B(n5556), .Z(n5561) );
  NAND U5833 ( .A(n5559), .B(n5558), .Z(n5560) );
  AND U5834 ( .A(n5561), .B(n5560), .Z(n5696) );
  NANDN U5835 ( .A(n5563), .B(n5562), .Z(n5567) );
  NANDN U5836 ( .A(n5565), .B(n5564), .Z(n5566) );
  AND U5837 ( .A(n5567), .B(n5566), .Z(n5662) );
  NAND U5838 ( .A(b[0]), .B(a[80]), .Z(n5568) );
  XNOR U5839 ( .A(b[1]), .B(n5568), .Z(n5570) );
  NANDN U5840 ( .A(b[0]), .B(a[79]), .Z(n5569) );
  NAND U5841 ( .A(n5570), .B(n5569), .Z(n5642) );
  NAND U5842 ( .A(n19808), .B(n5571), .Z(n5573) );
  XOR U5843 ( .A(b[13]), .B(a[68]), .Z(n5648) );
  NAND U5844 ( .A(n19768), .B(n5648), .Z(n5572) );
  AND U5845 ( .A(n5573), .B(n5572), .Z(n5640) );
  AND U5846 ( .A(b[15]), .B(a[64]), .Z(n5639) );
  XNOR U5847 ( .A(n5640), .B(n5639), .Z(n5641) );
  XNOR U5848 ( .A(n5642), .B(n5641), .Z(n5660) );
  NAND U5849 ( .A(n33), .B(n5574), .Z(n5576) );
  XOR U5850 ( .A(b[5]), .B(a[76]), .Z(n5651) );
  NAND U5851 ( .A(n19342), .B(n5651), .Z(n5575) );
  AND U5852 ( .A(n5576), .B(n5575), .Z(n5684) );
  NAND U5853 ( .A(n34), .B(n5577), .Z(n5579) );
  XOR U5854 ( .A(b[7]), .B(a[74]), .Z(n5654) );
  NAND U5855 ( .A(n19486), .B(n5654), .Z(n5578) );
  AND U5856 ( .A(n5579), .B(n5578), .Z(n5682) );
  NAND U5857 ( .A(n31), .B(n5580), .Z(n5582) );
  XOR U5858 ( .A(b[3]), .B(a[78]), .Z(n5657) );
  NAND U5859 ( .A(n32), .B(n5657), .Z(n5581) );
  NAND U5860 ( .A(n5582), .B(n5581), .Z(n5681) );
  XNOR U5861 ( .A(n5682), .B(n5681), .Z(n5683) );
  XOR U5862 ( .A(n5684), .B(n5683), .Z(n5661) );
  XOR U5863 ( .A(n5660), .B(n5661), .Z(n5663) );
  XOR U5864 ( .A(n5662), .B(n5663), .Z(n5634) );
  NANDN U5865 ( .A(n5584), .B(n5583), .Z(n5588) );
  OR U5866 ( .A(n5586), .B(n5585), .Z(n5587) );
  AND U5867 ( .A(n5588), .B(n5587), .Z(n5633) );
  XNOR U5868 ( .A(n5634), .B(n5633), .Z(n5636) );
  NAND U5869 ( .A(n5589), .B(n19724), .Z(n5591) );
  XOR U5870 ( .A(b[11]), .B(a[70]), .Z(n5666) );
  NAND U5871 ( .A(n19692), .B(n5666), .Z(n5590) );
  AND U5872 ( .A(n5591), .B(n5590), .Z(n5677) );
  NAND U5873 ( .A(n19838), .B(n5592), .Z(n5594) );
  XOR U5874 ( .A(b[15]), .B(a[66]), .Z(n5669) );
  NAND U5875 ( .A(n19805), .B(n5669), .Z(n5593) );
  AND U5876 ( .A(n5594), .B(n5593), .Z(n5676) );
  NAND U5877 ( .A(n35), .B(n5595), .Z(n5597) );
  XOR U5878 ( .A(b[9]), .B(a[72]), .Z(n5672) );
  NAND U5879 ( .A(n19598), .B(n5672), .Z(n5596) );
  NAND U5880 ( .A(n5597), .B(n5596), .Z(n5675) );
  XOR U5881 ( .A(n5676), .B(n5675), .Z(n5678) );
  XOR U5882 ( .A(n5677), .B(n5678), .Z(n5688) );
  NANDN U5883 ( .A(n5599), .B(n5598), .Z(n5603) );
  OR U5884 ( .A(n5601), .B(n5600), .Z(n5602) );
  AND U5885 ( .A(n5603), .B(n5602), .Z(n5687) );
  XNOR U5886 ( .A(n5688), .B(n5687), .Z(n5689) );
  NANDN U5887 ( .A(n5605), .B(n5604), .Z(n5609) );
  NANDN U5888 ( .A(n5607), .B(n5606), .Z(n5608) );
  NAND U5889 ( .A(n5609), .B(n5608), .Z(n5690) );
  XNOR U5890 ( .A(n5689), .B(n5690), .Z(n5635) );
  XOR U5891 ( .A(n5636), .B(n5635), .Z(n5694) );
  NANDN U5892 ( .A(n5611), .B(n5610), .Z(n5615) );
  NANDN U5893 ( .A(n5613), .B(n5612), .Z(n5614) );
  AND U5894 ( .A(n5615), .B(n5614), .Z(n5693) );
  XNOR U5895 ( .A(n5694), .B(n5693), .Z(n5695) );
  XOR U5896 ( .A(n5696), .B(n5695), .Z(n5628) );
  NANDN U5897 ( .A(n5617), .B(n5616), .Z(n5621) );
  NAND U5898 ( .A(n5619), .B(n5618), .Z(n5620) );
  AND U5899 ( .A(n5621), .B(n5620), .Z(n5627) );
  XNOR U5900 ( .A(n5628), .B(n5627), .Z(n5629) );
  XNOR U5901 ( .A(n5630), .B(n5629), .Z(n5699) );
  XNOR U5902 ( .A(sreg[320]), .B(n5699), .Z(n5701) );
  NANDN U5903 ( .A(sreg[319]), .B(n5622), .Z(n5626) );
  NAND U5904 ( .A(n5624), .B(n5623), .Z(n5625) );
  NAND U5905 ( .A(n5626), .B(n5625), .Z(n5700) );
  XNOR U5906 ( .A(n5701), .B(n5700), .Z(c[320]) );
  NANDN U5907 ( .A(n5628), .B(n5627), .Z(n5632) );
  NANDN U5908 ( .A(n5630), .B(n5629), .Z(n5631) );
  AND U5909 ( .A(n5632), .B(n5631), .Z(n5707) );
  NANDN U5910 ( .A(n5634), .B(n5633), .Z(n5638) );
  NAND U5911 ( .A(n5636), .B(n5635), .Z(n5637) );
  AND U5912 ( .A(n5638), .B(n5637), .Z(n5773) );
  NANDN U5913 ( .A(n5640), .B(n5639), .Z(n5644) );
  NANDN U5914 ( .A(n5642), .B(n5641), .Z(n5643) );
  AND U5915 ( .A(n5644), .B(n5643), .Z(n5760) );
  NAND U5916 ( .A(b[0]), .B(a[81]), .Z(n5645) );
  XNOR U5917 ( .A(b[1]), .B(n5645), .Z(n5647) );
  NANDN U5918 ( .A(b[0]), .B(a[80]), .Z(n5646) );
  NAND U5919 ( .A(n5647), .B(n5646), .Z(n5740) );
  NAND U5920 ( .A(n19808), .B(n5648), .Z(n5650) );
  XOR U5921 ( .A(b[13]), .B(a[69]), .Z(n5746) );
  NAND U5922 ( .A(n19768), .B(n5746), .Z(n5649) );
  AND U5923 ( .A(n5650), .B(n5649), .Z(n5738) );
  AND U5924 ( .A(b[15]), .B(a[65]), .Z(n5737) );
  XNOR U5925 ( .A(n5738), .B(n5737), .Z(n5739) );
  XNOR U5926 ( .A(n5740), .B(n5739), .Z(n5758) );
  NAND U5927 ( .A(n33), .B(n5651), .Z(n5653) );
  XOR U5928 ( .A(b[5]), .B(a[77]), .Z(n5749) );
  NAND U5929 ( .A(n19342), .B(n5749), .Z(n5652) );
  AND U5930 ( .A(n5653), .B(n5652), .Z(n5734) );
  NAND U5931 ( .A(n34), .B(n5654), .Z(n5656) );
  XOR U5932 ( .A(b[7]), .B(a[75]), .Z(n5752) );
  NAND U5933 ( .A(n19486), .B(n5752), .Z(n5655) );
  AND U5934 ( .A(n5656), .B(n5655), .Z(n5732) );
  NAND U5935 ( .A(n31), .B(n5657), .Z(n5659) );
  XOR U5936 ( .A(b[3]), .B(a[79]), .Z(n5755) );
  NAND U5937 ( .A(n32), .B(n5755), .Z(n5658) );
  NAND U5938 ( .A(n5659), .B(n5658), .Z(n5731) );
  XNOR U5939 ( .A(n5732), .B(n5731), .Z(n5733) );
  XOR U5940 ( .A(n5734), .B(n5733), .Z(n5759) );
  XOR U5941 ( .A(n5758), .B(n5759), .Z(n5761) );
  XOR U5942 ( .A(n5760), .B(n5761), .Z(n5711) );
  NANDN U5943 ( .A(n5661), .B(n5660), .Z(n5665) );
  OR U5944 ( .A(n5663), .B(n5662), .Z(n5664) );
  AND U5945 ( .A(n5665), .B(n5664), .Z(n5710) );
  XNOR U5946 ( .A(n5711), .B(n5710), .Z(n5713) );
  NAND U5947 ( .A(n5666), .B(n19724), .Z(n5668) );
  XOR U5948 ( .A(b[11]), .B(a[71]), .Z(n5716) );
  NAND U5949 ( .A(n19692), .B(n5716), .Z(n5667) );
  AND U5950 ( .A(n5668), .B(n5667), .Z(n5727) );
  NAND U5951 ( .A(n19838), .B(n5669), .Z(n5671) );
  XOR U5952 ( .A(b[15]), .B(a[67]), .Z(n5719) );
  NAND U5953 ( .A(n19805), .B(n5719), .Z(n5670) );
  AND U5954 ( .A(n5671), .B(n5670), .Z(n5726) );
  NAND U5955 ( .A(n35), .B(n5672), .Z(n5674) );
  XOR U5956 ( .A(b[9]), .B(a[73]), .Z(n5722) );
  NAND U5957 ( .A(n19598), .B(n5722), .Z(n5673) );
  NAND U5958 ( .A(n5674), .B(n5673), .Z(n5725) );
  XOR U5959 ( .A(n5726), .B(n5725), .Z(n5728) );
  XOR U5960 ( .A(n5727), .B(n5728), .Z(n5765) );
  NANDN U5961 ( .A(n5676), .B(n5675), .Z(n5680) );
  OR U5962 ( .A(n5678), .B(n5677), .Z(n5679) );
  AND U5963 ( .A(n5680), .B(n5679), .Z(n5764) );
  XNOR U5964 ( .A(n5765), .B(n5764), .Z(n5766) );
  NANDN U5965 ( .A(n5682), .B(n5681), .Z(n5686) );
  NANDN U5966 ( .A(n5684), .B(n5683), .Z(n5685) );
  NAND U5967 ( .A(n5686), .B(n5685), .Z(n5767) );
  XNOR U5968 ( .A(n5766), .B(n5767), .Z(n5712) );
  XOR U5969 ( .A(n5713), .B(n5712), .Z(n5771) );
  NANDN U5970 ( .A(n5688), .B(n5687), .Z(n5692) );
  NANDN U5971 ( .A(n5690), .B(n5689), .Z(n5691) );
  AND U5972 ( .A(n5692), .B(n5691), .Z(n5770) );
  XNOR U5973 ( .A(n5771), .B(n5770), .Z(n5772) );
  XOR U5974 ( .A(n5773), .B(n5772), .Z(n5705) );
  NANDN U5975 ( .A(n5694), .B(n5693), .Z(n5698) );
  NAND U5976 ( .A(n5696), .B(n5695), .Z(n5697) );
  AND U5977 ( .A(n5698), .B(n5697), .Z(n5704) );
  XNOR U5978 ( .A(n5705), .B(n5704), .Z(n5706) );
  XNOR U5979 ( .A(n5707), .B(n5706), .Z(n5776) );
  XNOR U5980 ( .A(sreg[321]), .B(n5776), .Z(n5778) );
  NANDN U5981 ( .A(sreg[320]), .B(n5699), .Z(n5703) );
  NAND U5982 ( .A(n5701), .B(n5700), .Z(n5702) );
  NAND U5983 ( .A(n5703), .B(n5702), .Z(n5777) );
  XNOR U5984 ( .A(n5778), .B(n5777), .Z(c[321]) );
  NANDN U5985 ( .A(n5705), .B(n5704), .Z(n5709) );
  NANDN U5986 ( .A(n5707), .B(n5706), .Z(n5708) );
  AND U5987 ( .A(n5709), .B(n5708), .Z(n5784) );
  NANDN U5988 ( .A(n5711), .B(n5710), .Z(n5715) );
  NAND U5989 ( .A(n5713), .B(n5712), .Z(n5714) );
  AND U5990 ( .A(n5715), .B(n5714), .Z(n5850) );
  NAND U5991 ( .A(n5716), .B(n19724), .Z(n5718) );
  XOR U5992 ( .A(b[11]), .B(a[72]), .Z(n5793) );
  NAND U5993 ( .A(n19692), .B(n5793), .Z(n5717) );
  AND U5994 ( .A(n5718), .B(n5717), .Z(n5804) );
  NAND U5995 ( .A(n19838), .B(n5719), .Z(n5721) );
  XOR U5996 ( .A(b[15]), .B(a[68]), .Z(n5796) );
  NAND U5997 ( .A(n19805), .B(n5796), .Z(n5720) );
  AND U5998 ( .A(n5721), .B(n5720), .Z(n5803) );
  NAND U5999 ( .A(n35), .B(n5722), .Z(n5724) );
  XOR U6000 ( .A(b[9]), .B(a[74]), .Z(n5799) );
  NAND U6001 ( .A(n19598), .B(n5799), .Z(n5723) );
  NAND U6002 ( .A(n5724), .B(n5723), .Z(n5802) );
  XOR U6003 ( .A(n5803), .B(n5802), .Z(n5805) );
  XOR U6004 ( .A(n5804), .B(n5805), .Z(n5842) );
  NANDN U6005 ( .A(n5726), .B(n5725), .Z(n5730) );
  OR U6006 ( .A(n5728), .B(n5727), .Z(n5729) );
  AND U6007 ( .A(n5730), .B(n5729), .Z(n5841) );
  XNOR U6008 ( .A(n5842), .B(n5841), .Z(n5843) );
  NANDN U6009 ( .A(n5732), .B(n5731), .Z(n5736) );
  NANDN U6010 ( .A(n5734), .B(n5733), .Z(n5735) );
  NAND U6011 ( .A(n5736), .B(n5735), .Z(n5844) );
  XNOR U6012 ( .A(n5843), .B(n5844), .Z(n5790) );
  NANDN U6013 ( .A(n5738), .B(n5737), .Z(n5742) );
  NANDN U6014 ( .A(n5740), .B(n5739), .Z(n5741) );
  AND U6015 ( .A(n5742), .B(n5741), .Z(n5837) );
  NAND U6016 ( .A(b[0]), .B(a[82]), .Z(n5743) );
  XNOR U6017 ( .A(b[1]), .B(n5743), .Z(n5745) );
  NANDN U6018 ( .A(b[0]), .B(a[81]), .Z(n5744) );
  NAND U6019 ( .A(n5745), .B(n5744), .Z(n5817) );
  NAND U6020 ( .A(n19808), .B(n5746), .Z(n5748) );
  XOR U6021 ( .A(b[13]), .B(a[70]), .Z(n5823) );
  NAND U6022 ( .A(n19768), .B(n5823), .Z(n5747) );
  AND U6023 ( .A(n5748), .B(n5747), .Z(n5815) );
  AND U6024 ( .A(b[15]), .B(a[66]), .Z(n5814) );
  XNOR U6025 ( .A(n5815), .B(n5814), .Z(n5816) );
  XNOR U6026 ( .A(n5817), .B(n5816), .Z(n5835) );
  NAND U6027 ( .A(n33), .B(n5749), .Z(n5751) );
  XOR U6028 ( .A(b[5]), .B(a[78]), .Z(n5826) );
  NAND U6029 ( .A(n19342), .B(n5826), .Z(n5750) );
  AND U6030 ( .A(n5751), .B(n5750), .Z(n5811) );
  NAND U6031 ( .A(n34), .B(n5752), .Z(n5754) );
  XOR U6032 ( .A(b[7]), .B(a[76]), .Z(n5829) );
  NAND U6033 ( .A(n19486), .B(n5829), .Z(n5753) );
  AND U6034 ( .A(n5754), .B(n5753), .Z(n5809) );
  NAND U6035 ( .A(n31), .B(n5755), .Z(n5757) );
  XOR U6036 ( .A(b[3]), .B(a[80]), .Z(n5832) );
  NAND U6037 ( .A(n32), .B(n5832), .Z(n5756) );
  NAND U6038 ( .A(n5757), .B(n5756), .Z(n5808) );
  XNOR U6039 ( .A(n5809), .B(n5808), .Z(n5810) );
  XOR U6040 ( .A(n5811), .B(n5810), .Z(n5836) );
  XOR U6041 ( .A(n5835), .B(n5836), .Z(n5838) );
  XOR U6042 ( .A(n5837), .B(n5838), .Z(n5788) );
  NANDN U6043 ( .A(n5759), .B(n5758), .Z(n5763) );
  OR U6044 ( .A(n5761), .B(n5760), .Z(n5762) );
  AND U6045 ( .A(n5763), .B(n5762), .Z(n5787) );
  XNOR U6046 ( .A(n5788), .B(n5787), .Z(n5789) );
  XOR U6047 ( .A(n5790), .B(n5789), .Z(n5848) );
  NANDN U6048 ( .A(n5765), .B(n5764), .Z(n5769) );
  NANDN U6049 ( .A(n5767), .B(n5766), .Z(n5768) );
  AND U6050 ( .A(n5769), .B(n5768), .Z(n5847) );
  XNOR U6051 ( .A(n5848), .B(n5847), .Z(n5849) );
  XOR U6052 ( .A(n5850), .B(n5849), .Z(n5782) );
  NANDN U6053 ( .A(n5771), .B(n5770), .Z(n5775) );
  NAND U6054 ( .A(n5773), .B(n5772), .Z(n5774) );
  AND U6055 ( .A(n5775), .B(n5774), .Z(n5781) );
  XNOR U6056 ( .A(n5782), .B(n5781), .Z(n5783) );
  XNOR U6057 ( .A(n5784), .B(n5783), .Z(n5853) );
  XNOR U6058 ( .A(sreg[322]), .B(n5853), .Z(n5855) );
  NANDN U6059 ( .A(sreg[321]), .B(n5776), .Z(n5780) );
  NAND U6060 ( .A(n5778), .B(n5777), .Z(n5779) );
  NAND U6061 ( .A(n5780), .B(n5779), .Z(n5854) );
  XNOR U6062 ( .A(n5855), .B(n5854), .Z(c[322]) );
  NANDN U6063 ( .A(n5782), .B(n5781), .Z(n5786) );
  NANDN U6064 ( .A(n5784), .B(n5783), .Z(n5785) );
  AND U6065 ( .A(n5786), .B(n5785), .Z(n5861) );
  NANDN U6066 ( .A(n5788), .B(n5787), .Z(n5792) );
  NAND U6067 ( .A(n5790), .B(n5789), .Z(n5791) );
  AND U6068 ( .A(n5792), .B(n5791), .Z(n5927) );
  NAND U6069 ( .A(n5793), .B(n19724), .Z(n5795) );
  XOR U6070 ( .A(b[11]), .B(a[73]), .Z(n5897) );
  NAND U6071 ( .A(n19692), .B(n5897), .Z(n5794) );
  AND U6072 ( .A(n5795), .B(n5794), .Z(n5908) );
  NAND U6073 ( .A(n19838), .B(n5796), .Z(n5798) );
  XOR U6074 ( .A(b[15]), .B(a[69]), .Z(n5900) );
  NAND U6075 ( .A(n19805), .B(n5900), .Z(n5797) );
  AND U6076 ( .A(n5798), .B(n5797), .Z(n5907) );
  NAND U6077 ( .A(n35), .B(n5799), .Z(n5801) );
  XOR U6078 ( .A(b[9]), .B(a[75]), .Z(n5903) );
  NAND U6079 ( .A(n19598), .B(n5903), .Z(n5800) );
  NAND U6080 ( .A(n5801), .B(n5800), .Z(n5906) );
  XOR U6081 ( .A(n5907), .B(n5906), .Z(n5909) );
  XOR U6082 ( .A(n5908), .B(n5909), .Z(n5919) );
  NANDN U6083 ( .A(n5803), .B(n5802), .Z(n5807) );
  OR U6084 ( .A(n5805), .B(n5804), .Z(n5806) );
  AND U6085 ( .A(n5807), .B(n5806), .Z(n5918) );
  XNOR U6086 ( .A(n5919), .B(n5918), .Z(n5920) );
  NANDN U6087 ( .A(n5809), .B(n5808), .Z(n5813) );
  NANDN U6088 ( .A(n5811), .B(n5810), .Z(n5812) );
  NAND U6089 ( .A(n5813), .B(n5812), .Z(n5921) );
  XNOR U6090 ( .A(n5920), .B(n5921), .Z(n5867) );
  NANDN U6091 ( .A(n5815), .B(n5814), .Z(n5819) );
  NANDN U6092 ( .A(n5817), .B(n5816), .Z(n5818) );
  AND U6093 ( .A(n5819), .B(n5818), .Z(n5893) );
  NAND U6094 ( .A(b[0]), .B(a[83]), .Z(n5820) );
  XNOR U6095 ( .A(b[1]), .B(n5820), .Z(n5822) );
  NANDN U6096 ( .A(b[0]), .B(a[82]), .Z(n5821) );
  NAND U6097 ( .A(n5822), .B(n5821), .Z(n5873) );
  NAND U6098 ( .A(n19808), .B(n5823), .Z(n5825) );
  XOR U6099 ( .A(b[13]), .B(a[71]), .Z(n5876) );
  NAND U6100 ( .A(n19768), .B(n5876), .Z(n5824) );
  AND U6101 ( .A(n5825), .B(n5824), .Z(n5871) );
  AND U6102 ( .A(b[15]), .B(a[67]), .Z(n5870) );
  XNOR U6103 ( .A(n5871), .B(n5870), .Z(n5872) );
  XNOR U6104 ( .A(n5873), .B(n5872), .Z(n5891) );
  NAND U6105 ( .A(n33), .B(n5826), .Z(n5828) );
  XOR U6106 ( .A(b[5]), .B(a[79]), .Z(n5882) );
  NAND U6107 ( .A(n19342), .B(n5882), .Z(n5827) );
  AND U6108 ( .A(n5828), .B(n5827), .Z(n5915) );
  NAND U6109 ( .A(n34), .B(n5829), .Z(n5831) );
  XOR U6110 ( .A(b[7]), .B(a[77]), .Z(n5885) );
  NAND U6111 ( .A(n19486), .B(n5885), .Z(n5830) );
  AND U6112 ( .A(n5831), .B(n5830), .Z(n5913) );
  NAND U6113 ( .A(n31), .B(n5832), .Z(n5834) );
  XOR U6114 ( .A(b[3]), .B(a[81]), .Z(n5888) );
  NAND U6115 ( .A(n32), .B(n5888), .Z(n5833) );
  NAND U6116 ( .A(n5834), .B(n5833), .Z(n5912) );
  XNOR U6117 ( .A(n5913), .B(n5912), .Z(n5914) );
  XOR U6118 ( .A(n5915), .B(n5914), .Z(n5892) );
  XOR U6119 ( .A(n5891), .B(n5892), .Z(n5894) );
  XOR U6120 ( .A(n5893), .B(n5894), .Z(n5865) );
  NANDN U6121 ( .A(n5836), .B(n5835), .Z(n5840) );
  OR U6122 ( .A(n5838), .B(n5837), .Z(n5839) );
  AND U6123 ( .A(n5840), .B(n5839), .Z(n5864) );
  XNOR U6124 ( .A(n5865), .B(n5864), .Z(n5866) );
  XOR U6125 ( .A(n5867), .B(n5866), .Z(n5925) );
  NANDN U6126 ( .A(n5842), .B(n5841), .Z(n5846) );
  NANDN U6127 ( .A(n5844), .B(n5843), .Z(n5845) );
  AND U6128 ( .A(n5846), .B(n5845), .Z(n5924) );
  XNOR U6129 ( .A(n5925), .B(n5924), .Z(n5926) );
  XOR U6130 ( .A(n5927), .B(n5926), .Z(n5859) );
  NANDN U6131 ( .A(n5848), .B(n5847), .Z(n5852) );
  NAND U6132 ( .A(n5850), .B(n5849), .Z(n5851) );
  AND U6133 ( .A(n5852), .B(n5851), .Z(n5858) );
  XNOR U6134 ( .A(n5859), .B(n5858), .Z(n5860) );
  XNOR U6135 ( .A(n5861), .B(n5860), .Z(n5930) );
  XNOR U6136 ( .A(sreg[323]), .B(n5930), .Z(n5932) );
  NANDN U6137 ( .A(sreg[322]), .B(n5853), .Z(n5857) );
  NAND U6138 ( .A(n5855), .B(n5854), .Z(n5856) );
  NAND U6139 ( .A(n5857), .B(n5856), .Z(n5931) );
  XNOR U6140 ( .A(n5932), .B(n5931), .Z(c[323]) );
  NANDN U6141 ( .A(n5859), .B(n5858), .Z(n5863) );
  NANDN U6142 ( .A(n5861), .B(n5860), .Z(n5862) );
  AND U6143 ( .A(n5863), .B(n5862), .Z(n5938) );
  NANDN U6144 ( .A(n5865), .B(n5864), .Z(n5869) );
  NAND U6145 ( .A(n5867), .B(n5866), .Z(n5868) );
  AND U6146 ( .A(n5869), .B(n5868), .Z(n6004) );
  NANDN U6147 ( .A(n5871), .B(n5870), .Z(n5875) );
  NANDN U6148 ( .A(n5873), .B(n5872), .Z(n5874) );
  AND U6149 ( .A(n5875), .B(n5874), .Z(n5970) );
  NAND U6150 ( .A(n19808), .B(n5876), .Z(n5878) );
  XOR U6151 ( .A(b[13]), .B(a[72]), .Z(n5956) );
  NAND U6152 ( .A(n19768), .B(n5956), .Z(n5877) );
  AND U6153 ( .A(n5878), .B(n5877), .Z(n5948) );
  AND U6154 ( .A(b[15]), .B(a[68]), .Z(n5947) );
  XNOR U6155 ( .A(n5948), .B(n5947), .Z(n5949) );
  NAND U6156 ( .A(b[0]), .B(a[84]), .Z(n5879) );
  XNOR U6157 ( .A(b[1]), .B(n5879), .Z(n5881) );
  NANDN U6158 ( .A(b[0]), .B(a[83]), .Z(n5880) );
  NAND U6159 ( .A(n5881), .B(n5880), .Z(n5950) );
  XNOR U6160 ( .A(n5949), .B(n5950), .Z(n5968) );
  NAND U6161 ( .A(n33), .B(n5882), .Z(n5884) );
  XOR U6162 ( .A(b[5]), .B(a[80]), .Z(n5959) );
  NAND U6163 ( .A(n19342), .B(n5959), .Z(n5883) );
  AND U6164 ( .A(n5884), .B(n5883), .Z(n5992) );
  NAND U6165 ( .A(n34), .B(n5885), .Z(n5887) );
  XOR U6166 ( .A(b[7]), .B(a[78]), .Z(n5962) );
  NAND U6167 ( .A(n19486), .B(n5962), .Z(n5886) );
  AND U6168 ( .A(n5887), .B(n5886), .Z(n5990) );
  NAND U6169 ( .A(n31), .B(n5888), .Z(n5890) );
  XOR U6170 ( .A(b[3]), .B(a[82]), .Z(n5965) );
  NAND U6171 ( .A(n32), .B(n5965), .Z(n5889) );
  NAND U6172 ( .A(n5890), .B(n5889), .Z(n5989) );
  XNOR U6173 ( .A(n5990), .B(n5989), .Z(n5991) );
  XOR U6174 ( .A(n5992), .B(n5991), .Z(n5969) );
  XOR U6175 ( .A(n5968), .B(n5969), .Z(n5971) );
  XOR U6176 ( .A(n5970), .B(n5971), .Z(n5942) );
  NANDN U6177 ( .A(n5892), .B(n5891), .Z(n5896) );
  OR U6178 ( .A(n5894), .B(n5893), .Z(n5895) );
  AND U6179 ( .A(n5896), .B(n5895), .Z(n5941) );
  XNOR U6180 ( .A(n5942), .B(n5941), .Z(n5944) );
  NAND U6181 ( .A(n5897), .B(n19724), .Z(n5899) );
  XOR U6182 ( .A(b[11]), .B(a[74]), .Z(n5974) );
  NAND U6183 ( .A(n19692), .B(n5974), .Z(n5898) );
  AND U6184 ( .A(n5899), .B(n5898), .Z(n5985) );
  NAND U6185 ( .A(n19838), .B(n5900), .Z(n5902) );
  XOR U6186 ( .A(b[15]), .B(a[70]), .Z(n5977) );
  NAND U6187 ( .A(n19805), .B(n5977), .Z(n5901) );
  AND U6188 ( .A(n5902), .B(n5901), .Z(n5984) );
  NAND U6189 ( .A(n35), .B(n5903), .Z(n5905) );
  XOR U6190 ( .A(b[9]), .B(a[76]), .Z(n5980) );
  NAND U6191 ( .A(n19598), .B(n5980), .Z(n5904) );
  NAND U6192 ( .A(n5905), .B(n5904), .Z(n5983) );
  XOR U6193 ( .A(n5984), .B(n5983), .Z(n5986) );
  XOR U6194 ( .A(n5985), .B(n5986), .Z(n5996) );
  NANDN U6195 ( .A(n5907), .B(n5906), .Z(n5911) );
  OR U6196 ( .A(n5909), .B(n5908), .Z(n5910) );
  AND U6197 ( .A(n5911), .B(n5910), .Z(n5995) );
  XNOR U6198 ( .A(n5996), .B(n5995), .Z(n5997) );
  NANDN U6199 ( .A(n5913), .B(n5912), .Z(n5917) );
  NANDN U6200 ( .A(n5915), .B(n5914), .Z(n5916) );
  NAND U6201 ( .A(n5917), .B(n5916), .Z(n5998) );
  XNOR U6202 ( .A(n5997), .B(n5998), .Z(n5943) );
  XOR U6203 ( .A(n5944), .B(n5943), .Z(n6002) );
  NANDN U6204 ( .A(n5919), .B(n5918), .Z(n5923) );
  NANDN U6205 ( .A(n5921), .B(n5920), .Z(n5922) );
  AND U6206 ( .A(n5923), .B(n5922), .Z(n6001) );
  XNOR U6207 ( .A(n6002), .B(n6001), .Z(n6003) );
  XOR U6208 ( .A(n6004), .B(n6003), .Z(n5936) );
  NANDN U6209 ( .A(n5925), .B(n5924), .Z(n5929) );
  NAND U6210 ( .A(n5927), .B(n5926), .Z(n5928) );
  AND U6211 ( .A(n5929), .B(n5928), .Z(n5935) );
  XNOR U6212 ( .A(n5936), .B(n5935), .Z(n5937) );
  XNOR U6213 ( .A(n5938), .B(n5937), .Z(n6007) );
  XNOR U6214 ( .A(sreg[324]), .B(n6007), .Z(n6009) );
  NANDN U6215 ( .A(sreg[323]), .B(n5930), .Z(n5934) );
  NAND U6216 ( .A(n5932), .B(n5931), .Z(n5933) );
  NAND U6217 ( .A(n5934), .B(n5933), .Z(n6008) );
  XNOR U6218 ( .A(n6009), .B(n6008), .Z(c[324]) );
  NANDN U6219 ( .A(n5936), .B(n5935), .Z(n5940) );
  NANDN U6220 ( .A(n5938), .B(n5937), .Z(n5939) );
  AND U6221 ( .A(n5940), .B(n5939), .Z(n6015) );
  NANDN U6222 ( .A(n5942), .B(n5941), .Z(n5946) );
  NAND U6223 ( .A(n5944), .B(n5943), .Z(n5945) );
  AND U6224 ( .A(n5946), .B(n5945), .Z(n6081) );
  NANDN U6225 ( .A(n5948), .B(n5947), .Z(n5952) );
  NANDN U6226 ( .A(n5950), .B(n5949), .Z(n5951) );
  AND U6227 ( .A(n5952), .B(n5951), .Z(n6047) );
  NAND U6228 ( .A(b[0]), .B(a[85]), .Z(n5953) );
  XNOR U6229 ( .A(b[1]), .B(n5953), .Z(n5955) );
  NANDN U6230 ( .A(b[0]), .B(a[84]), .Z(n5954) );
  NAND U6231 ( .A(n5955), .B(n5954), .Z(n6027) );
  NAND U6232 ( .A(n19808), .B(n5956), .Z(n5958) );
  XOR U6233 ( .A(b[13]), .B(a[73]), .Z(n6033) );
  NAND U6234 ( .A(n19768), .B(n6033), .Z(n5957) );
  AND U6235 ( .A(n5958), .B(n5957), .Z(n6025) );
  AND U6236 ( .A(b[15]), .B(a[69]), .Z(n6024) );
  XNOR U6237 ( .A(n6025), .B(n6024), .Z(n6026) );
  XNOR U6238 ( .A(n6027), .B(n6026), .Z(n6045) );
  NAND U6239 ( .A(n33), .B(n5959), .Z(n5961) );
  XOR U6240 ( .A(b[5]), .B(a[81]), .Z(n6036) );
  NAND U6241 ( .A(n19342), .B(n6036), .Z(n5960) );
  AND U6242 ( .A(n5961), .B(n5960), .Z(n6069) );
  NAND U6243 ( .A(n34), .B(n5962), .Z(n5964) );
  XOR U6244 ( .A(b[7]), .B(a[79]), .Z(n6039) );
  NAND U6245 ( .A(n19486), .B(n6039), .Z(n5963) );
  AND U6246 ( .A(n5964), .B(n5963), .Z(n6067) );
  NAND U6247 ( .A(n31), .B(n5965), .Z(n5967) );
  XOR U6248 ( .A(b[3]), .B(a[83]), .Z(n6042) );
  NAND U6249 ( .A(n32), .B(n6042), .Z(n5966) );
  NAND U6250 ( .A(n5967), .B(n5966), .Z(n6066) );
  XNOR U6251 ( .A(n6067), .B(n6066), .Z(n6068) );
  XOR U6252 ( .A(n6069), .B(n6068), .Z(n6046) );
  XOR U6253 ( .A(n6045), .B(n6046), .Z(n6048) );
  XOR U6254 ( .A(n6047), .B(n6048), .Z(n6019) );
  NANDN U6255 ( .A(n5969), .B(n5968), .Z(n5973) );
  OR U6256 ( .A(n5971), .B(n5970), .Z(n5972) );
  AND U6257 ( .A(n5973), .B(n5972), .Z(n6018) );
  XNOR U6258 ( .A(n6019), .B(n6018), .Z(n6021) );
  NAND U6259 ( .A(n5974), .B(n19724), .Z(n5976) );
  XOR U6260 ( .A(b[11]), .B(a[75]), .Z(n6051) );
  NAND U6261 ( .A(n19692), .B(n6051), .Z(n5975) );
  AND U6262 ( .A(n5976), .B(n5975), .Z(n6062) );
  NAND U6263 ( .A(n19838), .B(n5977), .Z(n5979) );
  XOR U6264 ( .A(b[15]), .B(a[71]), .Z(n6054) );
  NAND U6265 ( .A(n19805), .B(n6054), .Z(n5978) );
  AND U6266 ( .A(n5979), .B(n5978), .Z(n6061) );
  NAND U6267 ( .A(n35), .B(n5980), .Z(n5982) );
  XOR U6268 ( .A(b[9]), .B(a[77]), .Z(n6057) );
  NAND U6269 ( .A(n19598), .B(n6057), .Z(n5981) );
  NAND U6270 ( .A(n5982), .B(n5981), .Z(n6060) );
  XOR U6271 ( .A(n6061), .B(n6060), .Z(n6063) );
  XOR U6272 ( .A(n6062), .B(n6063), .Z(n6073) );
  NANDN U6273 ( .A(n5984), .B(n5983), .Z(n5988) );
  OR U6274 ( .A(n5986), .B(n5985), .Z(n5987) );
  AND U6275 ( .A(n5988), .B(n5987), .Z(n6072) );
  XNOR U6276 ( .A(n6073), .B(n6072), .Z(n6074) );
  NANDN U6277 ( .A(n5990), .B(n5989), .Z(n5994) );
  NANDN U6278 ( .A(n5992), .B(n5991), .Z(n5993) );
  NAND U6279 ( .A(n5994), .B(n5993), .Z(n6075) );
  XNOR U6280 ( .A(n6074), .B(n6075), .Z(n6020) );
  XOR U6281 ( .A(n6021), .B(n6020), .Z(n6079) );
  NANDN U6282 ( .A(n5996), .B(n5995), .Z(n6000) );
  NANDN U6283 ( .A(n5998), .B(n5997), .Z(n5999) );
  AND U6284 ( .A(n6000), .B(n5999), .Z(n6078) );
  XNOR U6285 ( .A(n6079), .B(n6078), .Z(n6080) );
  XOR U6286 ( .A(n6081), .B(n6080), .Z(n6013) );
  NANDN U6287 ( .A(n6002), .B(n6001), .Z(n6006) );
  NAND U6288 ( .A(n6004), .B(n6003), .Z(n6005) );
  AND U6289 ( .A(n6006), .B(n6005), .Z(n6012) );
  XNOR U6290 ( .A(n6013), .B(n6012), .Z(n6014) );
  XNOR U6291 ( .A(n6015), .B(n6014), .Z(n6084) );
  XNOR U6292 ( .A(sreg[325]), .B(n6084), .Z(n6086) );
  NANDN U6293 ( .A(sreg[324]), .B(n6007), .Z(n6011) );
  NAND U6294 ( .A(n6009), .B(n6008), .Z(n6010) );
  NAND U6295 ( .A(n6011), .B(n6010), .Z(n6085) );
  XNOR U6296 ( .A(n6086), .B(n6085), .Z(c[325]) );
  NANDN U6297 ( .A(n6013), .B(n6012), .Z(n6017) );
  NANDN U6298 ( .A(n6015), .B(n6014), .Z(n6016) );
  AND U6299 ( .A(n6017), .B(n6016), .Z(n6092) );
  NANDN U6300 ( .A(n6019), .B(n6018), .Z(n6023) );
  NAND U6301 ( .A(n6021), .B(n6020), .Z(n6022) );
  AND U6302 ( .A(n6023), .B(n6022), .Z(n6158) );
  NANDN U6303 ( .A(n6025), .B(n6024), .Z(n6029) );
  NANDN U6304 ( .A(n6027), .B(n6026), .Z(n6028) );
  AND U6305 ( .A(n6029), .B(n6028), .Z(n6124) );
  NAND U6306 ( .A(b[0]), .B(a[86]), .Z(n6030) );
  XNOR U6307 ( .A(b[1]), .B(n6030), .Z(n6032) );
  NANDN U6308 ( .A(b[0]), .B(a[85]), .Z(n6031) );
  NAND U6309 ( .A(n6032), .B(n6031), .Z(n6104) );
  NAND U6310 ( .A(n19808), .B(n6033), .Z(n6035) );
  XOR U6311 ( .A(b[13]), .B(a[74]), .Z(n6107) );
  NAND U6312 ( .A(n19768), .B(n6107), .Z(n6034) );
  AND U6313 ( .A(n6035), .B(n6034), .Z(n6102) );
  AND U6314 ( .A(b[15]), .B(a[70]), .Z(n6101) );
  XNOR U6315 ( .A(n6102), .B(n6101), .Z(n6103) );
  XNOR U6316 ( .A(n6104), .B(n6103), .Z(n6122) );
  NAND U6317 ( .A(n33), .B(n6036), .Z(n6038) );
  XOR U6318 ( .A(b[5]), .B(a[82]), .Z(n6113) );
  NAND U6319 ( .A(n19342), .B(n6113), .Z(n6037) );
  AND U6320 ( .A(n6038), .B(n6037), .Z(n6146) );
  NAND U6321 ( .A(n34), .B(n6039), .Z(n6041) );
  XOR U6322 ( .A(b[7]), .B(a[80]), .Z(n6116) );
  NAND U6323 ( .A(n19486), .B(n6116), .Z(n6040) );
  AND U6324 ( .A(n6041), .B(n6040), .Z(n6144) );
  NAND U6325 ( .A(n31), .B(n6042), .Z(n6044) );
  XOR U6326 ( .A(b[3]), .B(a[84]), .Z(n6119) );
  NAND U6327 ( .A(n32), .B(n6119), .Z(n6043) );
  NAND U6328 ( .A(n6044), .B(n6043), .Z(n6143) );
  XNOR U6329 ( .A(n6144), .B(n6143), .Z(n6145) );
  XOR U6330 ( .A(n6146), .B(n6145), .Z(n6123) );
  XOR U6331 ( .A(n6122), .B(n6123), .Z(n6125) );
  XOR U6332 ( .A(n6124), .B(n6125), .Z(n6096) );
  NANDN U6333 ( .A(n6046), .B(n6045), .Z(n6050) );
  OR U6334 ( .A(n6048), .B(n6047), .Z(n6049) );
  AND U6335 ( .A(n6050), .B(n6049), .Z(n6095) );
  XNOR U6336 ( .A(n6096), .B(n6095), .Z(n6098) );
  NAND U6337 ( .A(n6051), .B(n19724), .Z(n6053) );
  XOR U6338 ( .A(b[11]), .B(a[76]), .Z(n6128) );
  NAND U6339 ( .A(n19692), .B(n6128), .Z(n6052) );
  AND U6340 ( .A(n6053), .B(n6052), .Z(n6139) );
  NAND U6341 ( .A(n19838), .B(n6054), .Z(n6056) );
  XOR U6342 ( .A(b[15]), .B(a[72]), .Z(n6131) );
  NAND U6343 ( .A(n19805), .B(n6131), .Z(n6055) );
  AND U6344 ( .A(n6056), .B(n6055), .Z(n6138) );
  NAND U6345 ( .A(n35), .B(n6057), .Z(n6059) );
  XOR U6346 ( .A(b[9]), .B(a[78]), .Z(n6134) );
  NAND U6347 ( .A(n19598), .B(n6134), .Z(n6058) );
  NAND U6348 ( .A(n6059), .B(n6058), .Z(n6137) );
  XOR U6349 ( .A(n6138), .B(n6137), .Z(n6140) );
  XOR U6350 ( .A(n6139), .B(n6140), .Z(n6150) );
  NANDN U6351 ( .A(n6061), .B(n6060), .Z(n6065) );
  OR U6352 ( .A(n6063), .B(n6062), .Z(n6064) );
  AND U6353 ( .A(n6065), .B(n6064), .Z(n6149) );
  XNOR U6354 ( .A(n6150), .B(n6149), .Z(n6151) );
  NANDN U6355 ( .A(n6067), .B(n6066), .Z(n6071) );
  NANDN U6356 ( .A(n6069), .B(n6068), .Z(n6070) );
  NAND U6357 ( .A(n6071), .B(n6070), .Z(n6152) );
  XNOR U6358 ( .A(n6151), .B(n6152), .Z(n6097) );
  XOR U6359 ( .A(n6098), .B(n6097), .Z(n6156) );
  NANDN U6360 ( .A(n6073), .B(n6072), .Z(n6077) );
  NANDN U6361 ( .A(n6075), .B(n6074), .Z(n6076) );
  AND U6362 ( .A(n6077), .B(n6076), .Z(n6155) );
  XNOR U6363 ( .A(n6156), .B(n6155), .Z(n6157) );
  XOR U6364 ( .A(n6158), .B(n6157), .Z(n6090) );
  NANDN U6365 ( .A(n6079), .B(n6078), .Z(n6083) );
  NAND U6366 ( .A(n6081), .B(n6080), .Z(n6082) );
  AND U6367 ( .A(n6083), .B(n6082), .Z(n6089) );
  XNOR U6368 ( .A(n6090), .B(n6089), .Z(n6091) );
  XNOR U6369 ( .A(n6092), .B(n6091), .Z(n6161) );
  XNOR U6370 ( .A(sreg[326]), .B(n6161), .Z(n6163) );
  NANDN U6371 ( .A(sreg[325]), .B(n6084), .Z(n6088) );
  NAND U6372 ( .A(n6086), .B(n6085), .Z(n6087) );
  NAND U6373 ( .A(n6088), .B(n6087), .Z(n6162) );
  XNOR U6374 ( .A(n6163), .B(n6162), .Z(c[326]) );
  NANDN U6375 ( .A(n6090), .B(n6089), .Z(n6094) );
  NANDN U6376 ( .A(n6092), .B(n6091), .Z(n6093) );
  AND U6377 ( .A(n6094), .B(n6093), .Z(n6169) );
  NANDN U6378 ( .A(n6096), .B(n6095), .Z(n6100) );
  NAND U6379 ( .A(n6098), .B(n6097), .Z(n6099) );
  AND U6380 ( .A(n6100), .B(n6099), .Z(n6235) );
  NANDN U6381 ( .A(n6102), .B(n6101), .Z(n6106) );
  NANDN U6382 ( .A(n6104), .B(n6103), .Z(n6105) );
  AND U6383 ( .A(n6106), .B(n6105), .Z(n6201) );
  NAND U6384 ( .A(n19808), .B(n6107), .Z(n6109) );
  XOR U6385 ( .A(b[13]), .B(a[75]), .Z(n6187) );
  NAND U6386 ( .A(n19768), .B(n6187), .Z(n6108) );
  AND U6387 ( .A(n6109), .B(n6108), .Z(n6179) );
  AND U6388 ( .A(b[15]), .B(a[71]), .Z(n6178) );
  XNOR U6389 ( .A(n6179), .B(n6178), .Z(n6180) );
  NAND U6390 ( .A(b[0]), .B(a[87]), .Z(n6110) );
  XNOR U6391 ( .A(b[1]), .B(n6110), .Z(n6112) );
  NANDN U6392 ( .A(b[0]), .B(a[86]), .Z(n6111) );
  NAND U6393 ( .A(n6112), .B(n6111), .Z(n6181) );
  XNOR U6394 ( .A(n6180), .B(n6181), .Z(n6199) );
  NAND U6395 ( .A(n33), .B(n6113), .Z(n6115) );
  XOR U6396 ( .A(b[5]), .B(a[83]), .Z(n6190) );
  NAND U6397 ( .A(n19342), .B(n6190), .Z(n6114) );
  AND U6398 ( .A(n6115), .B(n6114), .Z(n6223) );
  NAND U6399 ( .A(n34), .B(n6116), .Z(n6118) );
  XOR U6400 ( .A(b[7]), .B(a[81]), .Z(n6193) );
  NAND U6401 ( .A(n19486), .B(n6193), .Z(n6117) );
  AND U6402 ( .A(n6118), .B(n6117), .Z(n6221) );
  NAND U6403 ( .A(n31), .B(n6119), .Z(n6121) );
  XOR U6404 ( .A(b[3]), .B(a[85]), .Z(n6196) );
  NAND U6405 ( .A(n32), .B(n6196), .Z(n6120) );
  NAND U6406 ( .A(n6121), .B(n6120), .Z(n6220) );
  XNOR U6407 ( .A(n6221), .B(n6220), .Z(n6222) );
  XOR U6408 ( .A(n6223), .B(n6222), .Z(n6200) );
  XOR U6409 ( .A(n6199), .B(n6200), .Z(n6202) );
  XOR U6410 ( .A(n6201), .B(n6202), .Z(n6173) );
  NANDN U6411 ( .A(n6123), .B(n6122), .Z(n6127) );
  OR U6412 ( .A(n6125), .B(n6124), .Z(n6126) );
  AND U6413 ( .A(n6127), .B(n6126), .Z(n6172) );
  XNOR U6414 ( .A(n6173), .B(n6172), .Z(n6175) );
  NAND U6415 ( .A(n6128), .B(n19724), .Z(n6130) );
  XOR U6416 ( .A(b[11]), .B(a[77]), .Z(n6205) );
  NAND U6417 ( .A(n19692), .B(n6205), .Z(n6129) );
  AND U6418 ( .A(n6130), .B(n6129), .Z(n6216) );
  NAND U6419 ( .A(n19838), .B(n6131), .Z(n6133) );
  XOR U6420 ( .A(b[15]), .B(a[73]), .Z(n6208) );
  NAND U6421 ( .A(n19805), .B(n6208), .Z(n6132) );
  AND U6422 ( .A(n6133), .B(n6132), .Z(n6215) );
  NAND U6423 ( .A(n35), .B(n6134), .Z(n6136) );
  XOR U6424 ( .A(b[9]), .B(a[79]), .Z(n6211) );
  NAND U6425 ( .A(n19598), .B(n6211), .Z(n6135) );
  NAND U6426 ( .A(n6136), .B(n6135), .Z(n6214) );
  XOR U6427 ( .A(n6215), .B(n6214), .Z(n6217) );
  XOR U6428 ( .A(n6216), .B(n6217), .Z(n6227) );
  NANDN U6429 ( .A(n6138), .B(n6137), .Z(n6142) );
  OR U6430 ( .A(n6140), .B(n6139), .Z(n6141) );
  AND U6431 ( .A(n6142), .B(n6141), .Z(n6226) );
  XNOR U6432 ( .A(n6227), .B(n6226), .Z(n6228) );
  NANDN U6433 ( .A(n6144), .B(n6143), .Z(n6148) );
  NANDN U6434 ( .A(n6146), .B(n6145), .Z(n6147) );
  NAND U6435 ( .A(n6148), .B(n6147), .Z(n6229) );
  XNOR U6436 ( .A(n6228), .B(n6229), .Z(n6174) );
  XOR U6437 ( .A(n6175), .B(n6174), .Z(n6233) );
  NANDN U6438 ( .A(n6150), .B(n6149), .Z(n6154) );
  NANDN U6439 ( .A(n6152), .B(n6151), .Z(n6153) );
  AND U6440 ( .A(n6154), .B(n6153), .Z(n6232) );
  XNOR U6441 ( .A(n6233), .B(n6232), .Z(n6234) );
  XOR U6442 ( .A(n6235), .B(n6234), .Z(n6167) );
  NANDN U6443 ( .A(n6156), .B(n6155), .Z(n6160) );
  NAND U6444 ( .A(n6158), .B(n6157), .Z(n6159) );
  AND U6445 ( .A(n6160), .B(n6159), .Z(n6166) );
  XNOR U6446 ( .A(n6167), .B(n6166), .Z(n6168) );
  XNOR U6447 ( .A(n6169), .B(n6168), .Z(n6238) );
  XNOR U6448 ( .A(sreg[327]), .B(n6238), .Z(n6240) );
  NANDN U6449 ( .A(sreg[326]), .B(n6161), .Z(n6165) );
  NAND U6450 ( .A(n6163), .B(n6162), .Z(n6164) );
  NAND U6451 ( .A(n6165), .B(n6164), .Z(n6239) );
  XNOR U6452 ( .A(n6240), .B(n6239), .Z(c[327]) );
  NANDN U6453 ( .A(n6167), .B(n6166), .Z(n6171) );
  NANDN U6454 ( .A(n6169), .B(n6168), .Z(n6170) );
  AND U6455 ( .A(n6171), .B(n6170), .Z(n6246) );
  NANDN U6456 ( .A(n6173), .B(n6172), .Z(n6177) );
  NAND U6457 ( .A(n6175), .B(n6174), .Z(n6176) );
  AND U6458 ( .A(n6177), .B(n6176), .Z(n6312) );
  NANDN U6459 ( .A(n6179), .B(n6178), .Z(n6183) );
  NANDN U6460 ( .A(n6181), .B(n6180), .Z(n6182) );
  AND U6461 ( .A(n6183), .B(n6182), .Z(n6278) );
  NAND U6462 ( .A(b[0]), .B(a[88]), .Z(n6184) );
  XNOR U6463 ( .A(b[1]), .B(n6184), .Z(n6186) );
  NANDN U6464 ( .A(b[0]), .B(a[87]), .Z(n6185) );
  NAND U6465 ( .A(n6186), .B(n6185), .Z(n6258) );
  NAND U6466 ( .A(n19808), .B(n6187), .Z(n6189) );
  XOR U6467 ( .A(b[13]), .B(a[76]), .Z(n6261) );
  NAND U6468 ( .A(n19768), .B(n6261), .Z(n6188) );
  AND U6469 ( .A(n6189), .B(n6188), .Z(n6256) );
  AND U6470 ( .A(b[15]), .B(a[72]), .Z(n6255) );
  XNOR U6471 ( .A(n6256), .B(n6255), .Z(n6257) );
  XNOR U6472 ( .A(n6258), .B(n6257), .Z(n6276) );
  NAND U6473 ( .A(n33), .B(n6190), .Z(n6192) );
  XOR U6474 ( .A(b[5]), .B(a[84]), .Z(n6267) );
  NAND U6475 ( .A(n19342), .B(n6267), .Z(n6191) );
  AND U6476 ( .A(n6192), .B(n6191), .Z(n6300) );
  NAND U6477 ( .A(n34), .B(n6193), .Z(n6195) );
  XOR U6478 ( .A(b[7]), .B(a[82]), .Z(n6270) );
  NAND U6479 ( .A(n19486), .B(n6270), .Z(n6194) );
  AND U6480 ( .A(n6195), .B(n6194), .Z(n6298) );
  NAND U6481 ( .A(n31), .B(n6196), .Z(n6198) );
  XOR U6482 ( .A(b[3]), .B(a[86]), .Z(n6273) );
  NAND U6483 ( .A(n32), .B(n6273), .Z(n6197) );
  NAND U6484 ( .A(n6198), .B(n6197), .Z(n6297) );
  XNOR U6485 ( .A(n6298), .B(n6297), .Z(n6299) );
  XOR U6486 ( .A(n6300), .B(n6299), .Z(n6277) );
  XOR U6487 ( .A(n6276), .B(n6277), .Z(n6279) );
  XOR U6488 ( .A(n6278), .B(n6279), .Z(n6250) );
  NANDN U6489 ( .A(n6200), .B(n6199), .Z(n6204) );
  OR U6490 ( .A(n6202), .B(n6201), .Z(n6203) );
  AND U6491 ( .A(n6204), .B(n6203), .Z(n6249) );
  XNOR U6492 ( .A(n6250), .B(n6249), .Z(n6252) );
  NAND U6493 ( .A(n6205), .B(n19724), .Z(n6207) );
  XOR U6494 ( .A(b[11]), .B(a[78]), .Z(n6282) );
  NAND U6495 ( .A(n19692), .B(n6282), .Z(n6206) );
  AND U6496 ( .A(n6207), .B(n6206), .Z(n6293) );
  NAND U6497 ( .A(n19838), .B(n6208), .Z(n6210) );
  XOR U6498 ( .A(b[15]), .B(a[74]), .Z(n6285) );
  NAND U6499 ( .A(n19805), .B(n6285), .Z(n6209) );
  AND U6500 ( .A(n6210), .B(n6209), .Z(n6292) );
  NAND U6501 ( .A(n35), .B(n6211), .Z(n6213) );
  XOR U6502 ( .A(b[9]), .B(a[80]), .Z(n6288) );
  NAND U6503 ( .A(n19598), .B(n6288), .Z(n6212) );
  NAND U6504 ( .A(n6213), .B(n6212), .Z(n6291) );
  XOR U6505 ( .A(n6292), .B(n6291), .Z(n6294) );
  XOR U6506 ( .A(n6293), .B(n6294), .Z(n6304) );
  NANDN U6507 ( .A(n6215), .B(n6214), .Z(n6219) );
  OR U6508 ( .A(n6217), .B(n6216), .Z(n6218) );
  AND U6509 ( .A(n6219), .B(n6218), .Z(n6303) );
  XNOR U6510 ( .A(n6304), .B(n6303), .Z(n6305) );
  NANDN U6511 ( .A(n6221), .B(n6220), .Z(n6225) );
  NANDN U6512 ( .A(n6223), .B(n6222), .Z(n6224) );
  NAND U6513 ( .A(n6225), .B(n6224), .Z(n6306) );
  XNOR U6514 ( .A(n6305), .B(n6306), .Z(n6251) );
  XOR U6515 ( .A(n6252), .B(n6251), .Z(n6310) );
  NANDN U6516 ( .A(n6227), .B(n6226), .Z(n6231) );
  NANDN U6517 ( .A(n6229), .B(n6228), .Z(n6230) );
  AND U6518 ( .A(n6231), .B(n6230), .Z(n6309) );
  XNOR U6519 ( .A(n6310), .B(n6309), .Z(n6311) );
  XOR U6520 ( .A(n6312), .B(n6311), .Z(n6244) );
  NANDN U6521 ( .A(n6233), .B(n6232), .Z(n6237) );
  NAND U6522 ( .A(n6235), .B(n6234), .Z(n6236) );
  AND U6523 ( .A(n6237), .B(n6236), .Z(n6243) );
  XNOR U6524 ( .A(n6244), .B(n6243), .Z(n6245) );
  XNOR U6525 ( .A(n6246), .B(n6245), .Z(n6315) );
  XNOR U6526 ( .A(sreg[328]), .B(n6315), .Z(n6317) );
  NANDN U6527 ( .A(sreg[327]), .B(n6238), .Z(n6242) );
  NAND U6528 ( .A(n6240), .B(n6239), .Z(n6241) );
  NAND U6529 ( .A(n6242), .B(n6241), .Z(n6316) );
  XNOR U6530 ( .A(n6317), .B(n6316), .Z(c[328]) );
  NANDN U6531 ( .A(n6244), .B(n6243), .Z(n6248) );
  NANDN U6532 ( .A(n6246), .B(n6245), .Z(n6247) );
  AND U6533 ( .A(n6248), .B(n6247), .Z(n6323) );
  NANDN U6534 ( .A(n6250), .B(n6249), .Z(n6254) );
  NAND U6535 ( .A(n6252), .B(n6251), .Z(n6253) );
  AND U6536 ( .A(n6254), .B(n6253), .Z(n6389) );
  NANDN U6537 ( .A(n6256), .B(n6255), .Z(n6260) );
  NANDN U6538 ( .A(n6258), .B(n6257), .Z(n6259) );
  AND U6539 ( .A(n6260), .B(n6259), .Z(n6355) );
  NAND U6540 ( .A(n19808), .B(n6261), .Z(n6263) );
  XOR U6541 ( .A(b[13]), .B(a[77]), .Z(n6341) );
  NAND U6542 ( .A(n19768), .B(n6341), .Z(n6262) );
  AND U6543 ( .A(n6263), .B(n6262), .Z(n6333) );
  AND U6544 ( .A(b[15]), .B(a[73]), .Z(n6332) );
  XNOR U6545 ( .A(n6333), .B(n6332), .Z(n6334) );
  NAND U6546 ( .A(b[0]), .B(a[89]), .Z(n6264) );
  XNOR U6547 ( .A(b[1]), .B(n6264), .Z(n6266) );
  NANDN U6548 ( .A(b[0]), .B(a[88]), .Z(n6265) );
  NAND U6549 ( .A(n6266), .B(n6265), .Z(n6335) );
  XNOR U6550 ( .A(n6334), .B(n6335), .Z(n6353) );
  NAND U6551 ( .A(n33), .B(n6267), .Z(n6269) );
  XOR U6552 ( .A(b[5]), .B(a[85]), .Z(n6344) );
  NAND U6553 ( .A(n19342), .B(n6344), .Z(n6268) );
  AND U6554 ( .A(n6269), .B(n6268), .Z(n6377) );
  NAND U6555 ( .A(n34), .B(n6270), .Z(n6272) );
  XOR U6556 ( .A(b[7]), .B(a[83]), .Z(n6347) );
  NAND U6557 ( .A(n19486), .B(n6347), .Z(n6271) );
  AND U6558 ( .A(n6272), .B(n6271), .Z(n6375) );
  NAND U6559 ( .A(n31), .B(n6273), .Z(n6275) );
  XOR U6560 ( .A(b[3]), .B(a[87]), .Z(n6350) );
  NAND U6561 ( .A(n32), .B(n6350), .Z(n6274) );
  NAND U6562 ( .A(n6275), .B(n6274), .Z(n6374) );
  XNOR U6563 ( .A(n6375), .B(n6374), .Z(n6376) );
  XOR U6564 ( .A(n6377), .B(n6376), .Z(n6354) );
  XOR U6565 ( .A(n6353), .B(n6354), .Z(n6356) );
  XOR U6566 ( .A(n6355), .B(n6356), .Z(n6327) );
  NANDN U6567 ( .A(n6277), .B(n6276), .Z(n6281) );
  OR U6568 ( .A(n6279), .B(n6278), .Z(n6280) );
  AND U6569 ( .A(n6281), .B(n6280), .Z(n6326) );
  XNOR U6570 ( .A(n6327), .B(n6326), .Z(n6329) );
  NAND U6571 ( .A(n6282), .B(n19724), .Z(n6284) );
  XOR U6572 ( .A(b[11]), .B(a[79]), .Z(n6359) );
  NAND U6573 ( .A(n19692), .B(n6359), .Z(n6283) );
  AND U6574 ( .A(n6284), .B(n6283), .Z(n6370) );
  NAND U6575 ( .A(n19838), .B(n6285), .Z(n6287) );
  XOR U6576 ( .A(b[15]), .B(a[75]), .Z(n6362) );
  NAND U6577 ( .A(n19805), .B(n6362), .Z(n6286) );
  AND U6578 ( .A(n6287), .B(n6286), .Z(n6369) );
  NAND U6579 ( .A(n35), .B(n6288), .Z(n6290) );
  XOR U6580 ( .A(b[9]), .B(a[81]), .Z(n6365) );
  NAND U6581 ( .A(n19598), .B(n6365), .Z(n6289) );
  NAND U6582 ( .A(n6290), .B(n6289), .Z(n6368) );
  XOR U6583 ( .A(n6369), .B(n6368), .Z(n6371) );
  XOR U6584 ( .A(n6370), .B(n6371), .Z(n6381) );
  NANDN U6585 ( .A(n6292), .B(n6291), .Z(n6296) );
  OR U6586 ( .A(n6294), .B(n6293), .Z(n6295) );
  AND U6587 ( .A(n6296), .B(n6295), .Z(n6380) );
  XNOR U6588 ( .A(n6381), .B(n6380), .Z(n6382) );
  NANDN U6589 ( .A(n6298), .B(n6297), .Z(n6302) );
  NANDN U6590 ( .A(n6300), .B(n6299), .Z(n6301) );
  NAND U6591 ( .A(n6302), .B(n6301), .Z(n6383) );
  XNOR U6592 ( .A(n6382), .B(n6383), .Z(n6328) );
  XOR U6593 ( .A(n6329), .B(n6328), .Z(n6387) );
  NANDN U6594 ( .A(n6304), .B(n6303), .Z(n6308) );
  NANDN U6595 ( .A(n6306), .B(n6305), .Z(n6307) );
  AND U6596 ( .A(n6308), .B(n6307), .Z(n6386) );
  XNOR U6597 ( .A(n6387), .B(n6386), .Z(n6388) );
  XOR U6598 ( .A(n6389), .B(n6388), .Z(n6321) );
  NANDN U6599 ( .A(n6310), .B(n6309), .Z(n6314) );
  NAND U6600 ( .A(n6312), .B(n6311), .Z(n6313) );
  AND U6601 ( .A(n6314), .B(n6313), .Z(n6320) );
  XNOR U6602 ( .A(n6321), .B(n6320), .Z(n6322) );
  XNOR U6603 ( .A(n6323), .B(n6322), .Z(n6392) );
  XNOR U6604 ( .A(sreg[329]), .B(n6392), .Z(n6394) );
  NANDN U6605 ( .A(sreg[328]), .B(n6315), .Z(n6319) );
  NAND U6606 ( .A(n6317), .B(n6316), .Z(n6318) );
  NAND U6607 ( .A(n6319), .B(n6318), .Z(n6393) );
  XNOR U6608 ( .A(n6394), .B(n6393), .Z(c[329]) );
  NANDN U6609 ( .A(n6321), .B(n6320), .Z(n6325) );
  NANDN U6610 ( .A(n6323), .B(n6322), .Z(n6324) );
  AND U6611 ( .A(n6325), .B(n6324), .Z(n6400) );
  NANDN U6612 ( .A(n6327), .B(n6326), .Z(n6331) );
  NAND U6613 ( .A(n6329), .B(n6328), .Z(n6330) );
  AND U6614 ( .A(n6331), .B(n6330), .Z(n6466) );
  NANDN U6615 ( .A(n6333), .B(n6332), .Z(n6337) );
  NANDN U6616 ( .A(n6335), .B(n6334), .Z(n6336) );
  AND U6617 ( .A(n6337), .B(n6336), .Z(n6432) );
  NAND U6618 ( .A(b[0]), .B(a[90]), .Z(n6338) );
  XNOR U6619 ( .A(b[1]), .B(n6338), .Z(n6340) );
  NANDN U6620 ( .A(b[0]), .B(a[89]), .Z(n6339) );
  NAND U6621 ( .A(n6340), .B(n6339), .Z(n6412) );
  NAND U6622 ( .A(n19808), .B(n6341), .Z(n6343) );
  XOR U6623 ( .A(b[13]), .B(a[78]), .Z(n6418) );
  NAND U6624 ( .A(n19768), .B(n6418), .Z(n6342) );
  AND U6625 ( .A(n6343), .B(n6342), .Z(n6410) );
  AND U6626 ( .A(b[15]), .B(a[74]), .Z(n6409) );
  XNOR U6627 ( .A(n6410), .B(n6409), .Z(n6411) );
  XNOR U6628 ( .A(n6412), .B(n6411), .Z(n6430) );
  NAND U6629 ( .A(n33), .B(n6344), .Z(n6346) );
  XOR U6630 ( .A(b[5]), .B(a[86]), .Z(n6421) );
  NAND U6631 ( .A(n19342), .B(n6421), .Z(n6345) );
  AND U6632 ( .A(n6346), .B(n6345), .Z(n6454) );
  NAND U6633 ( .A(n34), .B(n6347), .Z(n6349) );
  XOR U6634 ( .A(b[7]), .B(a[84]), .Z(n6424) );
  NAND U6635 ( .A(n19486), .B(n6424), .Z(n6348) );
  AND U6636 ( .A(n6349), .B(n6348), .Z(n6452) );
  NAND U6637 ( .A(n31), .B(n6350), .Z(n6352) );
  XOR U6638 ( .A(b[3]), .B(a[88]), .Z(n6427) );
  NAND U6639 ( .A(n32), .B(n6427), .Z(n6351) );
  NAND U6640 ( .A(n6352), .B(n6351), .Z(n6451) );
  XNOR U6641 ( .A(n6452), .B(n6451), .Z(n6453) );
  XOR U6642 ( .A(n6454), .B(n6453), .Z(n6431) );
  XOR U6643 ( .A(n6430), .B(n6431), .Z(n6433) );
  XOR U6644 ( .A(n6432), .B(n6433), .Z(n6404) );
  NANDN U6645 ( .A(n6354), .B(n6353), .Z(n6358) );
  OR U6646 ( .A(n6356), .B(n6355), .Z(n6357) );
  AND U6647 ( .A(n6358), .B(n6357), .Z(n6403) );
  XNOR U6648 ( .A(n6404), .B(n6403), .Z(n6406) );
  NAND U6649 ( .A(n6359), .B(n19724), .Z(n6361) );
  XOR U6650 ( .A(b[11]), .B(a[80]), .Z(n6436) );
  NAND U6651 ( .A(n19692), .B(n6436), .Z(n6360) );
  AND U6652 ( .A(n6361), .B(n6360), .Z(n6447) );
  NAND U6653 ( .A(n19838), .B(n6362), .Z(n6364) );
  XOR U6654 ( .A(b[15]), .B(a[76]), .Z(n6439) );
  NAND U6655 ( .A(n19805), .B(n6439), .Z(n6363) );
  AND U6656 ( .A(n6364), .B(n6363), .Z(n6446) );
  NAND U6657 ( .A(n35), .B(n6365), .Z(n6367) );
  XOR U6658 ( .A(b[9]), .B(a[82]), .Z(n6442) );
  NAND U6659 ( .A(n19598), .B(n6442), .Z(n6366) );
  NAND U6660 ( .A(n6367), .B(n6366), .Z(n6445) );
  XOR U6661 ( .A(n6446), .B(n6445), .Z(n6448) );
  XOR U6662 ( .A(n6447), .B(n6448), .Z(n6458) );
  NANDN U6663 ( .A(n6369), .B(n6368), .Z(n6373) );
  OR U6664 ( .A(n6371), .B(n6370), .Z(n6372) );
  AND U6665 ( .A(n6373), .B(n6372), .Z(n6457) );
  XNOR U6666 ( .A(n6458), .B(n6457), .Z(n6459) );
  NANDN U6667 ( .A(n6375), .B(n6374), .Z(n6379) );
  NANDN U6668 ( .A(n6377), .B(n6376), .Z(n6378) );
  NAND U6669 ( .A(n6379), .B(n6378), .Z(n6460) );
  XNOR U6670 ( .A(n6459), .B(n6460), .Z(n6405) );
  XOR U6671 ( .A(n6406), .B(n6405), .Z(n6464) );
  NANDN U6672 ( .A(n6381), .B(n6380), .Z(n6385) );
  NANDN U6673 ( .A(n6383), .B(n6382), .Z(n6384) );
  AND U6674 ( .A(n6385), .B(n6384), .Z(n6463) );
  XNOR U6675 ( .A(n6464), .B(n6463), .Z(n6465) );
  XOR U6676 ( .A(n6466), .B(n6465), .Z(n6398) );
  NANDN U6677 ( .A(n6387), .B(n6386), .Z(n6391) );
  NAND U6678 ( .A(n6389), .B(n6388), .Z(n6390) );
  AND U6679 ( .A(n6391), .B(n6390), .Z(n6397) );
  XNOR U6680 ( .A(n6398), .B(n6397), .Z(n6399) );
  XNOR U6681 ( .A(n6400), .B(n6399), .Z(n6469) );
  XNOR U6682 ( .A(sreg[330]), .B(n6469), .Z(n6471) );
  NANDN U6683 ( .A(sreg[329]), .B(n6392), .Z(n6396) );
  NAND U6684 ( .A(n6394), .B(n6393), .Z(n6395) );
  NAND U6685 ( .A(n6396), .B(n6395), .Z(n6470) );
  XNOR U6686 ( .A(n6471), .B(n6470), .Z(c[330]) );
  NANDN U6687 ( .A(n6398), .B(n6397), .Z(n6402) );
  NANDN U6688 ( .A(n6400), .B(n6399), .Z(n6401) );
  AND U6689 ( .A(n6402), .B(n6401), .Z(n6477) );
  NANDN U6690 ( .A(n6404), .B(n6403), .Z(n6408) );
  NAND U6691 ( .A(n6406), .B(n6405), .Z(n6407) );
  AND U6692 ( .A(n6408), .B(n6407), .Z(n6543) );
  NANDN U6693 ( .A(n6410), .B(n6409), .Z(n6414) );
  NANDN U6694 ( .A(n6412), .B(n6411), .Z(n6413) );
  AND U6695 ( .A(n6414), .B(n6413), .Z(n6509) );
  NAND U6696 ( .A(b[0]), .B(a[91]), .Z(n6415) );
  XNOR U6697 ( .A(b[1]), .B(n6415), .Z(n6417) );
  NANDN U6698 ( .A(b[0]), .B(a[90]), .Z(n6416) );
  NAND U6699 ( .A(n6417), .B(n6416), .Z(n6489) );
  NAND U6700 ( .A(n19808), .B(n6418), .Z(n6420) );
  XOR U6701 ( .A(b[13]), .B(a[79]), .Z(n6495) );
  NAND U6702 ( .A(n19768), .B(n6495), .Z(n6419) );
  AND U6703 ( .A(n6420), .B(n6419), .Z(n6487) );
  AND U6704 ( .A(b[15]), .B(a[75]), .Z(n6486) );
  XNOR U6705 ( .A(n6487), .B(n6486), .Z(n6488) );
  XNOR U6706 ( .A(n6489), .B(n6488), .Z(n6507) );
  NAND U6707 ( .A(n33), .B(n6421), .Z(n6423) );
  XOR U6708 ( .A(b[5]), .B(a[87]), .Z(n6498) );
  NAND U6709 ( .A(n19342), .B(n6498), .Z(n6422) );
  AND U6710 ( .A(n6423), .B(n6422), .Z(n6531) );
  NAND U6711 ( .A(n34), .B(n6424), .Z(n6426) );
  XOR U6712 ( .A(b[7]), .B(a[85]), .Z(n6501) );
  NAND U6713 ( .A(n19486), .B(n6501), .Z(n6425) );
  AND U6714 ( .A(n6426), .B(n6425), .Z(n6529) );
  NAND U6715 ( .A(n31), .B(n6427), .Z(n6429) );
  XOR U6716 ( .A(b[3]), .B(a[89]), .Z(n6504) );
  NAND U6717 ( .A(n32), .B(n6504), .Z(n6428) );
  NAND U6718 ( .A(n6429), .B(n6428), .Z(n6528) );
  XNOR U6719 ( .A(n6529), .B(n6528), .Z(n6530) );
  XOR U6720 ( .A(n6531), .B(n6530), .Z(n6508) );
  XOR U6721 ( .A(n6507), .B(n6508), .Z(n6510) );
  XOR U6722 ( .A(n6509), .B(n6510), .Z(n6481) );
  NANDN U6723 ( .A(n6431), .B(n6430), .Z(n6435) );
  OR U6724 ( .A(n6433), .B(n6432), .Z(n6434) );
  AND U6725 ( .A(n6435), .B(n6434), .Z(n6480) );
  XNOR U6726 ( .A(n6481), .B(n6480), .Z(n6483) );
  NAND U6727 ( .A(n6436), .B(n19724), .Z(n6438) );
  XOR U6728 ( .A(b[11]), .B(a[81]), .Z(n6513) );
  NAND U6729 ( .A(n19692), .B(n6513), .Z(n6437) );
  AND U6730 ( .A(n6438), .B(n6437), .Z(n6524) );
  NAND U6731 ( .A(n19838), .B(n6439), .Z(n6441) );
  XOR U6732 ( .A(b[15]), .B(a[77]), .Z(n6516) );
  NAND U6733 ( .A(n19805), .B(n6516), .Z(n6440) );
  AND U6734 ( .A(n6441), .B(n6440), .Z(n6523) );
  NAND U6735 ( .A(n35), .B(n6442), .Z(n6444) );
  XOR U6736 ( .A(b[9]), .B(a[83]), .Z(n6519) );
  NAND U6737 ( .A(n19598), .B(n6519), .Z(n6443) );
  NAND U6738 ( .A(n6444), .B(n6443), .Z(n6522) );
  XOR U6739 ( .A(n6523), .B(n6522), .Z(n6525) );
  XOR U6740 ( .A(n6524), .B(n6525), .Z(n6535) );
  NANDN U6741 ( .A(n6446), .B(n6445), .Z(n6450) );
  OR U6742 ( .A(n6448), .B(n6447), .Z(n6449) );
  AND U6743 ( .A(n6450), .B(n6449), .Z(n6534) );
  XNOR U6744 ( .A(n6535), .B(n6534), .Z(n6536) );
  NANDN U6745 ( .A(n6452), .B(n6451), .Z(n6456) );
  NANDN U6746 ( .A(n6454), .B(n6453), .Z(n6455) );
  NAND U6747 ( .A(n6456), .B(n6455), .Z(n6537) );
  XNOR U6748 ( .A(n6536), .B(n6537), .Z(n6482) );
  XOR U6749 ( .A(n6483), .B(n6482), .Z(n6541) );
  NANDN U6750 ( .A(n6458), .B(n6457), .Z(n6462) );
  NANDN U6751 ( .A(n6460), .B(n6459), .Z(n6461) );
  AND U6752 ( .A(n6462), .B(n6461), .Z(n6540) );
  XNOR U6753 ( .A(n6541), .B(n6540), .Z(n6542) );
  XOR U6754 ( .A(n6543), .B(n6542), .Z(n6475) );
  NANDN U6755 ( .A(n6464), .B(n6463), .Z(n6468) );
  NAND U6756 ( .A(n6466), .B(n6465), .Z(n6467) );
  AND U6757 ( .A(n6468), .B(n6467), .Z(n6474) );
  XNOR U6758 ( .A(n6475), .B(n6474), .Z(n6476) );
  XNOR U6759 ( .A(n6477), .B(n6476), .Z(n6546) );
  XNOR U6760 ( .A(sreg[331]), .B(n6546), .Z(n6548) );
  NANDN U6761 ( .A(sreg[330]), .B(n6469), .Z(n6473) );
  NAND U6762 ( .A(n6471), .B(n6470), .Z(n6472) );
  NAND U6763 ( .A(n6473), .B(n6472), .Z(n6547) );
  XNOR U6764 ( .A(n6548), .B(n6547), .Z(c[331]) );
  NANDN U6765 ( .A(n6475), .B(n6474), .Z(n6479) );
  NANDN U6766 ( .A(n6477), .B(n6476), .Z(n6478) );
  AND U6767 ( .A(n6479), .B(n6478), .Z(n6554) );
  NANDN U6768 ( .A(n6481), .B(n6480), .Z(n6485) );
  NAND U6769 ( .A(n6483), .B(n6482), .Z(n6484) );
  AND U6770 ( .A(n6485), .B(n6484), .Z(n6620) );
  NANDN U6771 ( .A(n6487), .B(n6486), .Z(n6491) );
  NANDN U6772 ( .A(n6489), .B(n6488), .Z(n6490) );
  AND U6773 ( .A(n6491), .B(n6490), .Z(n6607) );
  NAND U6774 ( .A(b[0]), .B(a[92]), .Z(n6492) );
  XNOR U6775 ( .A(b[1]), .B(n6492), .Z(n6494) );
  NANDN U6776 ( .A(b[0]), .B(a[91]), .Z(n6493) );
  NAND U6777 ( .A(n6494), .B(n6493), .Z(n6587) );
  NAND U6778 ( .A(n19808), .B(n6495), .Z(n6497) );
  XOR U6779 ( .A(b[13]), .B(a[80]), .Z(n6590) );
  NAND U6780 ( .A(n19768), .B(n6590), .Z(n6496) );
  AND U6781 ( .A(n6497), .B(n6496), .Z(n6585) );
  AND U6782 ( .A(b[15]), .B(a[76]), .Z(n6584) );
  XNOR U6783 ( .A(n6585), .B(n6584), .Z(n6586) );
  XNOR U6784 ( .A(n6587), .B(n6586), .Z(n6605) );
  NAND U6785 ( .A(n33), .B(n6498), .Z(n6500) );
  XOR U6786 ( .A(b[5]), .B(a[88]), .Z(n6596) );
  NAND U6787 ( .A(n19342), .B(n6596), .Z(n6499) );
  AND U6788 ( .A(n6500), .B(n6499), .Z(n6581) );
  NAND U6789 ( .A(n34), .B(n6501), .Z(n6503) );
  XOR U6790 ( .A(b[7]), .B(a[86]), .Z(n6599) );
  NAND U6791 ( .A(n19486), .B(n6599), .Z(n6502) );
  AND U6792 ( .A(n6503), .B(n6502), .Z(n6579) );
  NAND U6793 ( .A(n31), .B(n6504), .Z(n6506) );
  XOR U6794 ( .A(b[3]), .B(a[90]), .Z(n6602) );
  NAND U6795 ( .A(n32), .B(n6602), .Z(n6505) );
  NAND U6796 ( .A(n6506), .B(n6505), .Z(n6578) );
  XNOR U6797 ( .A(n6579), .B(n6578), .Z(n6580) );
  XOR U6798 ( .A(n6581), .B(n6580), .Z(n6606) );
  XOR U6799 ( .A(n6605), .B(n6606), .Z(n6608) );
  XOR U6800 ( .A(n6607), .B(n6608), .Z(n6558) );
  NANDN U6801 ( .A(n6508), .B(n6507), .Z(n6512) );
  OR U6802 ( .A(n6510), .B(n6509), .Z(n6511) );
  AND U6803 ( .A(n6512), .B(n6511), .Z(n6557) );
  XNOR U6804 ( .A(n6558), .B(n6557), .Z(n6560) );
  NAND U6805 ( .A(n6513), .B(n19724), .Z(n6515) );
  XOR U6806 ( .A(b[11]), .B(a[82]), .Z(n6563) );
  NAND U6807 ( .A(n19692), .B(n6563), .Z(n6514) );
  AND U6808 ( .A(n6515), .B(n6514), .Z(n6574) );
  NAND U6809 ( .A(n19838), .B(n6516), .Z(n6518) );
  XOR U6810 ( .A(b[15]), .B(a[78]), .Z(n6566) );
  NAND U6811 ( .A(n19805), .B(n6566), .Z(n6517) );
  AND U6812 ( .A(n6518), .B(n6517), .Z(n6573) );
  NAND U6813 ( .A(n35), .B(n6519), .Z(n6521) );
  XOR U6814 ( .A(b[9]), .B(a[84]), .Z(n6569) );
  NAND U6815 ( .A(n19598), .B(n6569), .Z(n6520) );
  NAND U6816 ( .A(n6521), .B(n6520), .Z(n6572) );
  XOR U6817 ( .A(n6573), .B(n6572), .Z(n6575) );
  XOR U6818 ( .A(n6574), .B(n6575), .Z(n6612) );
  NANDN U6819 ( .A(n6523), .B(n6522), .Z(n6527) );
  OR U6820 ( .A(n6525), .B(n6524), .Z(n6526) );
  AND U6821 ( .A(n6527), .B(n6526), .Z(n6611) );
  XNOR U6822 ( .A(n6612), .B(n6611), .Z(n6613) );
  NANDN U6823 ( .A(n6529), .B(n6528), .Z(n6533) );
  NANDN U6824 ( .A(n6531), .B(n6530), .Z(n6532) );
  NAND U6825 ( .A(n6533), .B(n6532), .Z(n6614) );
  XNOR U6826 ( .A(n6613), .B(n6614), .Z(n6559) );
  XOR U6827 ( .A(n6560), .B(n6559), .Z(n6618) );
  NANDN U6828 ( .A(n6535), .B(n6534), .Z(n6539) );
  NANDN U6829 ( .A(n6537), .B(n6536), .Z(n6538) );
  AND U6830 ( .A(n6539), .B(n6538), .Z(n6617) );
  XNOR U6831 ( .A(n6618), .B(n6617), .Z(n6619) );
  XOR U6832 ( .A(n6620), .B(n6619), .Z(n6552) );
  NANDN U6833 ( .A(n6541), .B(n6540), .Z(n6545) );
  NAND U6834 ( .A(n6543), .B(n6542), .Z(n6544) );
  AND U6835 ( .A(n6545), .B(n6544), .Z(n6551) );
  XNOR U6836 ( .A(n6552), .B(n6551), .Z(n6553) );
  XNOR U6837 ( .A(n6554), .B(n6553), .Z(n6623) );
  XNOR U6838 ( .A(sreg[332]), .B(n6623), .Z(n6625) );
  NANDN U6839 ( .A(sreg[331]), .B(n6546), .Z(n6550) );
  NAND U6840 ( .A(n6548), .B(n6547), .Z(n6549) );
  NAND U6841 ( .A(n6550), .B(n6549), .Z(n6624) );
  XNOR U6842 ( .A(n6625), .B(n6624), .Z(c[332]) );
  NANDN U6843 ( .A(n6552), .B(n6551), .Z(n6556) );
  NANDN U6844 ( .A(n6554), .B(n6553), .Z(n6555) );
  AND U6845 ( .A(n6556), .B(n6555), .Z(n6631) );
  NANDN U6846 ( .A(n6558), .B(n6557), .Z(n6562) );
  NAND U6847 ( .A(n6560), .B(n6559), .Z(n6561) );
  AND U6848 ( .A(n6562), .B(n6561), .Z(n6697) );
  NAND U6849 ( .A(n6563), .B(n19724), .Z(n6565) );
  XOR U6850 ( .A(b[11]), .B(a[83]), .Z(n6667) );
  NAND U6851 ( .A(n19692), .B(n6667), .Z(n6564) );
  AND U6852 ( .A(n6565), .B(n6564), .Z(n6678) );
  NAND U6853 ( .A(n19838), .B(n6566), .Z(n6568) );
  XOR U6854 ( .A(b[15]), .B(a[79]), .Z(n6670) );
  NAND U6855 ( .A(n19805), .B(n6670), .Z(n6567) );
  AND U6856 ( .A(n6568), .B(n6567), .Z(n6677) );
  NAND U6857 ( .A(n35), .B(n6569), .Z(n6571) );
  XOR U6858 ( .A(b[9]), .B(a[85]), .Z(n6673) );
  NAND U6859 ( .A(n19598), .B(n6673), .Z(n6570) );
  NAND U6860 ( .A(n6571), .B(n6570), .Z(n6676) );
  XOR U6861 ( .A(n6677), .B(n6676), .Z(n6679) );
  XOR U6862 ( .A(n6678), .B(n6679), .Z(n6689) );
  NANDN U6863 ( .A(n6573), .B(n6572), .Z(n6577) );
  OR U6864 ( .A(n6575), .B(n6574), .Z(n6576) );
  AND U6865 ( .A(n6577), .B(n6576), .Z(n6688) );
  XNOR U6866 ( .A(n6689), .B(n6688), .Z(n6690) );
  NANDN U6867 ( .A(n6579), .B(n6578), .Z(n6583) );
  NANDN U6868 ( .A(n6581), .B(n6580), .Z(n6582) );
  NAND U6869 ( .A(n6583), .B(n6582), .Z(n6691) );
  XNOR U6870 ( .A(n6690), .B(n6691), .Z(n6637) );
  NANDN U6871 ( .A(n6585), .B(n6584), .Z(n6589) );
  NANDN U6872 ( .A(n6587), .B(n6586), .Z(n6588) );
  AND U6873 ( .A(n6589), .B(n6588), .Z(n6663) );
  NAND U6874 ( .A(n19808), .B(n6590), .Z(n6592) );
  XOR U6875 ( .A(b[13]), .B(a[81]), .Z(n6649) );
  NAND U6876 ( .A(n19768), .B(n6649), .Z(n6591) );
  AND U6877 ( .A(n6592), .B(n6591), .Z(n6641) );
  AND U6878 ( .A(b[15]), .B(a[77]), .Z(n6640) );
  XNOR U6879 ( .A(n6641), .B(n6640), .Z(n6642) );
  NAND U6880 ( .A(b[0]), .B(a[93]), .Z(n6593) );
  XNOR U6881 ( .A(b[1]), .B(n6593), .Z(n6595) );
  NANDN U6882 ( .A(b[0]), .B(a[92]), .Z(n6594) );
  NAND U6883 ( .A(n6595), .B(n6594), .Z(n6643) );
  XNOR U6884 ( .A(n6642), .B(n6643), .Z(n6661) );
  NAND U6885 ( .A(n33), .B(n6596), .Z(n6598) );
  XOR U6886 ( .A(b[5]), .B(a[89]), .Z(n6652) );
  NAND U6887 ( .A(n19342), .B(n6652), .Z(n6597) );
  AND U6888 ( .A(n6598), .B(n6597), .Z(n6685) );
  NAND U6889 ( .A(n34), .B(n6599), .Z(n6601) );
  XOR U6890 ( .A(b[7]), .B(a[87]), .Z(n6655) );
  NAND U6891 ( .A(n19486), .B(n6655), .Z(n6600) );
  AND U6892 ( .A(n6601), .B(n6600), .Z(n6683) );
  NAND U6893 ( .A(n31), .B(n6602), .Z(n6604) );
  XOR U6894 ( .A(b[3]), .B(a[91]), .Z(n6658) );
  NAND U6895 ( .A(n32), .B(n6658), .Z(n6603) );
  NAND U6896 ( .A(n6604), .B(n6603), .Z(n6682) );
  XNOR U6897 ( .A(n6683), .B(n6682), .Z(n6684) );
  XOR U6898 ( .A(n6685), .B(n6684), .Z(n6662) );
  XOR U6899 ( .A(n6661), .B(n6662), .Z(n6664) );
  XOR U6900 ( .A(n6663), .B(n6664), .Z(n6635) );
  NANDN U6901 ( .A(n6606), .B(n6605), .Z(n6610) );
  OR U6902 ( .A(n6608), .B(n6607), .Z(n6609) );
  AND U6903 ( .A(n6610), .B(n6609), .Z(n6634) );
  XNOR U6904 ( .A(n6635), .B(n6634), .Z(n6636) );
  XOR U6905 ( .A(n6637), .B(n6636), .Z(n6695) );
  NANDN U6906 ( .A(n6612), .B(n6611), .Z(n6616) );
  NANDN U6907 ( .A(n6614), .B(n6613), .Z(n6615) );
  AND U6908 ( .A(n6616), .B(n6615), .Z(n6694) );
  XNOR U6909 ( .A(n6695), .B(n6694), .Z(n6696) );
  XOR U6910 ( .A(n6697), .B(n6696), .Z(n6629) );
  NANDN U6911 ( .A(n6618), .B(n6617), .Z(n6622) );
  NAND U6912 ( .A(n6620), .B(n6619), .Z(n6621) );
  AND U6913 ( .A(n6622), .B(n6621), .Z(n6628) );
  XNOR U6914 ( .A(n6629), .B(n6628), .Z(n6630) );
  XNOR U6915 ( .A(n6631), .B(n6630), .Z(n6700) );
  XNOR U6916 ( .A(sreg[333]), .B(n6700), .Z(n6702) );
  NANDN U6917 ( .A(sreg[332]), .B(n6623), .Z(n6627) );
  NAND U6918 ( .A(n6625), .B(n6624), .Z(n6626) );
  NAND U6919 ( .A(n6627), .B(n6626), .Z(n6701) );
  XNOR U6920 ( .A(n6702), .B(n6701), .Z(c[333]) );
  NANDN U6921 ( .A(n6629), .B(n6628), .Z(n6633) );
  NANDN U6922 ( .A(n6631), .B(n6630), .Z(n6632) );
  AND U6923 ( .A(n6633), .B(n6632), .Z(n6708) );
  NANDN U6924 ( .A(n6635), .B(n6634), .Z(n6639) );
  NAND U6925 ( .A(n6637), .B(n6636), .Z(n6638) );
  AND U6926 ( .A(n6639), .B(n6638), .Z(n6774) );
  NANDN U6927 ( .A(n6641), .B(n6640), .Z(n6645) );
  NANDN U6928 ( .A(n6643), .B(n6642), .Z(n6644) );
  AND U6929 ( .A(n6645), .B(n6644), .Z(n6740) );
  NAND U6930 ( .A(b[0]), .B(a[94]), .Z(n6646) );
  XNOR U6931 ( .A(b[1]), .B(n6646), .Z(n6648) );
  NANDN U6932 ( .A(b[0]), .B(a[93]), .Z(n6647) );
  NAND U6933 ( .A(n6648), .B(n6647), .Z(n6720) );
  NAND U6934 ( .A(n19808), .B(n6649), .Z(n6651) );
  XOR U6935 ( .A(b[13]), .B(a[82]), .Z(n6726) );
  NAND U6936 ( .A(n19768), .B(n6726), .Z(n6650) );
  AND U6937 ( .A(n6651), .B(n6650), .Z(n6718) );
  AND U6938 ( .A(b[15]), .B(a[78]), .Z(n6717) );
  XNOR U6939 ( .A(n6718), .B(n6717), .Z(n6719) );
  XNOR U6940 ( .A(n6720), .B(n6719), .Z(n6738) );
  NAND U6941 ( .A(n33), .B(n6652), .Z(n6654) );
  XOR U6942 ( .A(b[5]), .B(a[90]), .Z(n6729) );
  NAND U6943 ( .A(n19342), .B(n6729), .Z(n6653) );
  AND U6944 ( .A(n6654), .B(n6653), .Z(n6762) );
  NAND U6945 ( .A(n34), .B(n6655), .Z(n6657) );
  XOR U6946 ( .A(b[7]), .B(a[88]), .Z(n6732) );
  NAND U6947 ( .A(n19486), .B(n6732), .Z(n6656) );
  AND U6948 ( .A(n6657), .B(n6656), .Z(n6760) );
  NAND U6949 ( .A(n31), .B(n6658), .Z(n6660) );
  XOR U6950 ( .A(b[3]), .B(a[92]), .Z(n6735) );
  NAND U6951 ( .A(n32), .B(n6735), .Z(n6659) );
  NAND U6952 ( .A(n6660), .B(n6659), .Z(n6759) );
  XNOR U6953 ( .A(n6760), .B(n6759), .Z(n6761) );
  XOR U6954 ( .A(n6762), .B(n6761), .Z(n6739) );
  XOR U6955 ( .A(n6738), .B(n6739), .Z(n6741) );
  XOR U6956 ( .A(n6740), .B(n6741), .Z(n6712) );
  NANDN U6957 ( .A(n6662), .B(n6661), .Z(n6666) );
  OR U6958 ( .A(n6664), .B(n6663), .Z(n6665) );
  AND U6959 ( .A(n6666), .B(n6665), .Z(n6711) );
  XNOR U6960 ( .A(n6712), .B(n6711), .Z(n6714) );
  NAND U6961 ( .A(n6667), .B(n19724), .Z(n6669) );
  XOR U6962 ( .A(b[11]), .B(a[84]), .Z(n6744) );
  NAND U6963 ( .A(n19692), .B(n6744), .Z(n6668) );
  AND U6964 ( .A(n6669), .B(n6668), .Z(n6755) );
  NAND U6965 ( .A(n19838), .B(n6670), .Z(n6672) );
  XOR U6966 ( .A(b[15]), .B(a[80]), .Z(n6747) );
  NAND U6967 ( .A(n19805), .B(n6747), .Z(n6671) );
  AND U6968 ( .A(n6672), .B(n6671), .Z(n6754) );
  NAND U6969 ( .A(n35), .B(n6673), .Z(n6675) );
  XOR U6970 ( .A(b[9]), .B(a[86]), .Z(n6750) );
  NAND U6971 ( .A(n19598), .B(n6750), .Z(n6674) );
  NAND U6972 ( .A(n6675), .B(n6674), .Z(n6753) );
  XOR U6973 ( .A(n6754), .B(n6753), .Z(n6756) );
  XOR U6974 ( .A(n6755), .B(n6756), .Z(n6766) );
  NANDN U6975 ( .A(n6677), .B(n6676), .Z(n6681) );
  OR U6976 ( .A(n6679), .B(n6678), .Z(n6680) );
  AND U6977 ( .A(n6681), .B(n6680), .Z(n6765) );
  XNOR U6978 ( .A(n6766), .B(n6765), .Z(n6767) );
  NANDN U6979 ( .A(n6683), .B(n6682), .Z(n6687) );
  NANDN U6980 ( .A(n6685), .B(n6684), .Z(n6686) );
  NAND U6981 ( .A(n6687), .B(n6686), .Z(n6768) );
  XNOR U6982 ( .A(n6767), .B(n6768), .Z(n6713) );
  XOR U6983 ( .A(n6714), .B(n6713), .Z(n6772) );
  NANDN U6984 ( .A(n6689), .B(n6688), .Z(n6693) );
  NANDN U6985 ( .A(n6691), .B(n6690), .Z(n6692) );
  AND U6986 ( .A(n6693), .B(n6692), .Z(n6771) );
  XNOR U6987 ( .A(n6772), .B(n6771), .Z(n6773) );
  XOR U6988 ( .A(n6774), .B(n6773), .Z(n6706) );
  NANDN U6989 ( .A(n6695), .B(n6694), .Z(n6699) );
  NAND U6990 ( .A(n6697), .B(n6696), .Z(n6698) );
  AND U6991 ( .A(n6699), .B(n6698), .Z(n6705) );
  XNOR U6992 ( .A(n6706), .B(n6705), .Z(n6707) );
  XNOR U6993 ( .A(n6708), .B(n6707), .Z(n6777) );
  XNOR U6994 ( .A(sreg[334]), .B(n6777), .Z(n6779) );
  NANDN U6995 ( .A(sreg[333]), .B(n6700), .Z(n6704) );
  NAND U6996 ( .A(n6702), .B(n6701), .Z(n6703) );
  NAND U6997 ( .A(n6704), .B(n6703), .Z(n6778) );
  XNOR U6998 ( .A(n6779), .B(n6778), .Z(c[334]) );
  NANDN U6999 ( .A(n6706), .B(n6705), .Z(n6710) );
  NANDN U7000 ( .A(n6708), .B(n6707), .Z(n6709) );
  AND U7001 ( .A(n6710), .B(n6709), .Z(n6785) );
  NANDN U7002 ( .A(n6712), .B(n6711), .Z(n6716) );
  NAND U7003 ( .A(n6714), .B(n6713), .Z(n6715) );
  AND U7004 ( .A(n6716), .B(n6715), .Z(n6851) );
  NANDN U7005 ( .A(n6718), .B(n6717), .Z(n6722) );
  NANDN U7006 ( .A(n6720), .B(n6719), .Z(n6721) );
  AND U7007 ( .A(n6722), .B(n6721), .Z(n6817) );
  NAND U7008 ( .A(b[0]), .B(a[95]), .Z(n6723) );
  XNOR U7009 ( .A(b[1]), .B(n6723), .Z(n6725) );
  NANDN U7010 ( .A(b[0]), .B(a[94]), .Z(n6724) );
  NAND U7011 ( .A(n6725), .B(n6724), .Z(n6797) );
  NAND U7012 ( .A(n19808), .B(n6726), .Z(n6728) );
  XOR U7013 ( .A(b[13]), .B(a[83]), .Z(n6803) );
  NAND U7014 ( .A(n19768), .B(n6803), .Z(n6727) );
  AND U7015 ( .A(n6728), .B(n6727), .Z(n6795) );
  AND U7016 ( .A(b[15]), .B(a[79]), .Z(n6794) );
  XNOR U7017 ( .A(n6795), .B(n6794), .Z(n6796) );
  XNOR U7018 ( .A(n6797), .B(n6796), .Z(n6815) );
  NAND U7019 ( .A(n33), .B(n6729), .Z(n6731) );
  XOR U7020 ( .A(b[5]), .B(a[91]), .Z(n6806) );
  NAND U7021 ( .A(n19342), .B(n6806), .Z(n6730) );
  AND U7022 ( .A(n6731), .B(n6730), .Z(n6839) );
  NAND U7023 ( .A(n34), .B(n6732), .Z(n6734) );
  XOR U7024 ( .A(b[7]), .B(a[89]), .Z(n6809) );
  NAND U7025 ( .A(n19486), .B(n6809), .Z(n6733) );
  AND U7026 ( .A(n6734), .B(n6733), .Z(n6837) );
  NAND U7027 ( .A(n31), .B(n6735), .Z(n6737) );
  XOR U7028 ( .A(b[3]), .B(a[93]), .Z(n6812) );
  NAND U7029 ( .A(n32), .B(n6812), .Z(n6736) );
  NAND U7030 ( .A(n6737), .B(n6736), .Z(n6836) );
  XNOR U7031 ( .A(n6837), .B(n6836), .Z(n6838) );
  XOR U7032 ( .A(n6839), .B(n6838), .Z(n6816) );
  XOR U7033 ( .A(n6815), .B(n6816), .Z(n6818) );
  XOR U7034 ( .A(n6817), .B(n6818), .Z(n6789) );
  NANDN U7035 ( .A(n6739), .B(n6738), .Z(n6743) );
  OR U7036 ( .A(n6741), .B(n6740), .Z(n6742) );
  AND U7037 ( .A(n6743), .B(n6742), .Z(n6788) );
  XNOR U7038 ( .A(n6789), .B(n6788), .Z(n6791) );
  NAND U7039 ( .A(n6744), .B(n19724), .Z(n6746) );
  XOR U7040 ( .A(b[11]), .B(a[85]), .Z(n6821) );
  NAND U7041 ( .A(n19692), .B(n6821), .Z(n6745) );
  AND U7042 ( .A(n6746), .B(n6745), .Z(n6832) );
  NAND U7043 ( .A(n19838), .B(n6747), .Z(n6749) );
  XOR U7044 ( .A(b[15]), .B(a[81]), .Z(n6824) );
  NAND U7045 ( .A(n19805), .B(n6824), .Z(n6748) );
  AND U7046 ( .A(n6749), .B(n6748), .Z(n6831) );
  NAND U7047 ( .A(n35), .B(n6750), .Z(n6752) );
  XOR U7048 ( .A(b[9]), .B(a[87]), .Z(n6827) );
  NAND U7049 ( .A(n19598), .B(n6827), .Z(n6751) );
  NAND U7050 ( .A(n6752), .B(n6751), .Z(n6830) );
  XOR U7051 ( .A(n6831), .B(n6830), .Z(n6833) );
  XOR U7052 ( .A(n6832), .B(n6833), .Z(n6843) );
  NANDN U7053 ( .A(n6754), .B(n6753), .Z(n6758) );
  OR U7054 ( .A(n6756), .B(n6755), .Z(n6757) );
  AND U7055 ( .A(n6758), .B(n6757), .Z(n6842) );
  XNOR U7056 ( .A(n6843), .B(n6842), .Z(n6844) );
  NANDN U7057 ( .A(n6760), .B(n6759), .Z(n6764) );
  NANDN U7058 ( .A(n6762), .B(n6761), .Z(n6763) );
  NAND U7059 ( .A(n6764), .B(n6763), .Z(n6845) );
  XNOR U7060 ( .A(n6844), .B(n6845), .Z(n6790) );
  XOR U7061 ( .A(n6791), .B(n6790), .Z(n6849) );
  NANDN U7062 ( .A(n6766), .B(n6765), .Z(n6770) );
  NANDN U7063 ( .A(n6768), .B(n6767), .Z(n6769) );
  AND U7064 ( .A(n6770), .B(n6769), .Z(n6848) );
  XNOR U7065 ( .A(n6849), .B(n6848), .Z(n6850) );
  XOR U7066 ( .A(n6851), .B(n6850), .Z(n6783) );
  NANDN U7067 ( .A(n6772), .B(n6771), .Z(n6776) );
  NAND U7068 ( .A(n6774), .B(n6773), .Z(n6775) );
  AND U7069 ( .A(n6776), .B(n6775), .Z(n6782) );
  XNOR U7070 ( .A(n6783), .B(n6782), .Z(n6784) );
  XNOR U7071 ( .A(n6785), .B(n6784), .Z(n6854) );
  XNOR U7072 ( .A(sreg[335]), .B(n6854), .Z(n6856) );
  NANDN U7073 ( .A(sreg[334]), .B(n6777), .Z(n6781) );
  NAND U7074 ( .A(n6779), .B(n6778), .Z(n6780) );
  NAND U7075 ( .A(n6781), .B(n6780), .Z(n6855) );
  XNOR U7076 ( .A(n6856), .B(n6855), .Z(c[335]) );
  NANDN U7077 ( .A(n6783), .B(n6782), .Z(n6787) );
  NANDN U7078 ( .A(n6785), .B(n6784), .Z(n6786) );
  AND U7079 ( .A(n6787), .B(n6786), .Z(n6862) );
  NANDN U7080 ( .A(n6789), .B(n6788), .Z(n6793) );
  NAND U7081 ( .A(n6791), .B(n6790), .Z(n6792) );
  AND U7082 ( .A(n6793), .B(n6792), .Z(n6928) );
  NANDN U7083 ( .A(n6795), .B(n6794), .Z(n6799) );
  NANDN U7084 ( .A(n6797), .B(n6796), .Z(n6798) );
  AND U7085 ( .A(n6799), .B(n6798), .Z(n6894) );
  NAND U7086 ( .A(b[0]), .B(a[96]), .Z(n6800) );
  XNOR U7087 ( .A(b[1]), .B(n6800), .Z(n6802) );
  NANDN U7088 ( .A(b[0]), .B(a[95]), .Z(n6801) );
  NAND U7089 ( .A(n6802), .B(n6801), .Z(n6874) );
  NAND U7090 ( .A(n19808), .B(n6803), .Z(n6805) );
  XOR U7091 ( .A(b[13]), .B(a[84]), .Z(n6880) );
  NAND U7092 ( .A(n19768), .B(n6880), .Z(n6804) );
  AND U7093 ( .A(n6805), .B(n6804), .Z(n6872) );
  AND U7094 ( .A(b[15]), .B(a[80]), .Z(n6871) );
  XNOR U7095 ( .A(n6872), .B(n6871), .Z(n6873) );
  XNOR U7096 ( .A(n6874), .B(n6873), .Z(n6892) );
  NAND U7097 ( .A(n33), .B(n6806), .Z(n6808) );
  XOR U7098 ( .A(b[5]), .B(a[92]), .Z(n6883) );
  NAND U7099 ( .A(n19342), .B(n6883), .Z(n6807) );
  AND U7100 ( .A(n6808), .B(n6807), .Z(n6916) );
  NAND U7101 ( .A(n34), .B(n6809), .Z(n6811) );
  XOR U7102 ( .A(b[7]), .B(a[90]), .Z(n6886) );
  NAND U7103 ( .A(n19486), .B(n6886), .Z(n6810) );
  AND U7104 ( .A(n6811), .B(n6810), .Z(n6914) );
  NAND U7105 ( .A(n31), .B(n6812), .Z(n6814) );
  XOR U7106 ( .A(b[3]), .B(a[94]), .Z(n6889) );
  NAND U7107 ( .A(n32), .B(n6889), .Z(n6813) );
  NAND U7108 ( .A(n6814), .B(n6813), .Z(n6913) );
  XNOR U7109 ( .A(n6914), .B(n6913), .Z(n6915) );
  XOR U7110 ( .A(n6916), .B(n6915), .Z(n6893) );
  XOR U7111 ( .A(n6892), .B(n6893), .Z(n6895) );
  XOR U7112 ( .A(n6894), .B(n6895), .Z(n6866) );
  NANDN U7113 ( .A(n6816), .B(n6815), .Z(n6820) );
  OR U7114 ( .A(n6818), .B(n6817), .Z(n6819) );
  AND U7115 ( .A(n6820), .B(n6819), .Z(n6865) );
  XNOR U7116 ( .A(n6866), .B(n6865), .Z(n6868) );
  NAND U7117 ( .A(n6821), .B(n19724), .Z(n6823) );
  XOR U7118 ( .A(b[11]), .B(a[86]), .Z(n6898) );
  NAND U7119 ( .A(n19692), .B(n6898), .Z(n6822) );
  AND U7120 ( .A(n6823), .B(n6822), .Z(n6909) );
  NAND U7121 ( .A(n19838), .B(n6824), .Z(n6826) );
  XOR U7122 ( .A(b[15]), .B(a[82]), .Z(n6901) );
  NAND U7123 ( .A(n19805), .B(n6901), .Z(n6825) );
  AND U7124 ( .A(n6826), .B(n6825), .Z(n6908) );
  NAND U7125 ( .A(n35), .B(n6827), .Z(n6829) );
  XOR U7126 ( .A(b[9]), .B(a[88]), .Z(n6904) );
  NAND U7127 ( .A(n19598), .B(n6904), .Z(n6828) );
  NAND U7128 ( .A(n6829), .B(n6828), .Z(n6907) );
  XOR U7129 ( .A(n6908), .B(n6907), .Z(n6910) );
  XOR U7130 ( .A(n6909), .B(n6910), .Z(n6920) );
  NANDN U7131 ( .A(n6831), .B(n6830), .Z(n6835) );
  OR U7132 ( .A(n6833), .B(n6832), .Z(n6834) );
  AND U7133 ( .A(n6835), .B(n6834), .Z(n6919) );
  XNOR U7134 ( .A(n6920), .B(n6919), .Z(n6921) );
  NANDN U7135 ( .A(n6837), .B(n6836), .Z(n6841) );
  NANDN U7136 ( .A(n6839), .B(n6838), .Z(n6840) );
  NAND U7137 ( .A(n6841), .B(n6840), .Z(n6922) );
  XNOR U7138 ( .A(n6921), .B(n6922), .Z(n6867) );
  XOR U7139 ( .A(n6868), .B(n6867), .Z(n6926) );
  NANDN U7140 ( .A(n6843), .B(n6842), .Z(n6847) );
  NANDN U7141 ( .A(n6845), .B(n6844), .Z(n6846) );
  AND U7142 ( .A(n6847), .B(n6846), .Z(n6925) );
  XNOR U7143 ( .A(n6926), .B(n6925), .Z(n6927) );
  XOR U7144 ( .A(n6928), .B(n6927), .Z(n6860) );
  NANDN U7145 ( .A(n6849), .B(n6848), .Z(n6853) );
  NAND U7146 ( .A(n6851), .B(n6850), .Z(n6852) );
  AND U7147 ( .A(n6853), .B(n6852), .Z(n6859) );
  XNOR U7148 ( .A(n6860), .B(n6859), .Z(n6861) );
  XNOR U7149 ( .A(n6862), .B(n6861), .Z(n6931) );
  XNOR U7150 ( .A(sreg[336]), .B(n6931), .Z(n6933) );
  NANDN U7151 ( .A(sreg[335]), .B(n6854), .Z(n6858) );
  NAND U7152 ( .A(n6856), .B(n6855), .Z(n6857) );
  NAND U7153 ( .A(n6858), .B(n6857), .Z(n6932) );
  XNOR U7154 ( .A(n6933), .B(n6932), .Z(c[336]) );
  NANDN U7155 ( .A(n6860), .B(n6859), .Z(n6864) );
  NANDN U7156 ( .A(n6862), .B(n6861), .Z(n6863) );
  AND U7157 ( .A(n6864), .B(n6863), .Z(n6939) );
  NANDN U7158 ( .A(n6866), .B(n6865), .Z(n6870) );
  NAND U7159 ( .A(n6868), .B(n6867), .Z(n6869) );
  AND U7160 ( .A(n6870), .B(n6869), .Z(n7005) );
  NANDN U7161 ( .A(n6872), .B(n6871), .Z(n6876) );
  NANDN U7162 ( .A(n6874), .B(n6873), .Z(n6875) );
  AND U7163 ( .A(n6876), .B(n6875), .Z(n6971) );
  NAND U7164 ( .A(b[0]), .B(a[97]), .Z(n6877) );
  XNOR U7165 ( .A(b[1]), .B(n6877), .Z(n6879) );
  NANDN U7166 ( .A(b[0]), .B(a[96]), .Z(n6878) );
  NAND U7167 ( .A(n6879), .B(n6878), .Z(n6951) );
  NAND U7168 ( .A(n19808), .B(n6880), .Z(n6882) );
  XOR U7169 ( .A(b[13]), .B(a[85]), .Z(n6957) );
  NAND U7170 ( .A(n19768), .B(n6957), .Z(n6881) );
  AND U7171 ( .A(n6882), .B(n6881), .Z(n6949) );
  AND U7172 ( .A(b[15]), .B(a[81]), .Z(n6948) );
  XNOR U7173 ( .A(n6949), .B(n6948), .Z(n6950) );
  XNOR U7174 ( .A(n6951), .B(n6950), .Z(n6969) );
  NAND U7175 ( .A(n33), .B(n6883), .Z(n6885) );
  XOR U7176 ( .A(b[5]), .B(a[93]), .Z(n6960) );
  NAND U7177 ( .A(n19342), .B(n6960), .Z(n6884) );
  AND U7178 ( .A(n6885), .B(n6884), .Z(n6993) );
  NAND U7179 ( .A(n34), .B(n6886), .Z(n6888) );
  XOR U7180 ( .A(b[7]), .B(a[91]), .Z(n6963) );
  NAND U7181 ( .A(n19486), .B(n6963), .Z(n6887) );
  AND U7182 ( .A(n6888), .B(n6887), .Z(n6991) );
  NAND U7183 ( .A(n31), .B(n6889), .Z(n6891) );
  XOR U7184 ( .A(b[3]), .B(a[95]), .Z(n6966) );
  NAND U7185 ( .A(n32), .B(n6966), .Z(n6890) );
  NAND U7186 ( .A(n6891), .B(n6890), .Z(n6990) );
  XNOR U7187 ( .A(n6991), .B(n6990), .Z(n6992) );
  XOR U7188 ( .A(n6993), .B(n6992), .Z(n6970) );
  XOR U7189 ( .A(n6969), .B(n6970), .Z(n6972) );
  XOR U7190 ( .A(n6971), .B(n6972), .Z(n6943) );
  NANDN U7191 ( .A(n6893), .B(n6892), .Z(n6897) );
  OR U7192 ( .A(n6895), .B(n6894), .Z(n6896) );
  AND U7193 ( .A(n6897), .B(n6896), .Z(n6942) );
  XNOR U7194 ( .A(n6943), .B(n6942), .Z(n6945) );
  NAND U7195 ( .A(n6898), .B(n19724), .Z(n6900) );
  XOR U7196 ( .A(b[11]), .B(a[87]), .Z(n6975) );
  NAND U7197 ( .A(n19692), .B(n6975), .Z(n6899) );
  AND U7198 ( .A(n6900), .B(n6899), .Z(n6986) );
  NAND U7199 ( .A(n19838), .B(n6901), .Z(n6903) );
  XOR U7200 ( .A(b[15]), .B(a[83]), .Z(n6978) );
  NAND U7201 ( .A(n19805), .B(n6978), .Z(n6902) );
  AND U7202 ( .A(n6903), .B(n6902), .Z(n6985) );
  NAND U7203 ( .A(n35), .B(n6904), .Z(n6906) );
  XOR U7204 ( .A(b[9]), .B(a[89]), .Z(n6981) );
  NAND U7205 ( .A(n19598), .B(n6981), .Z(n6905) );
  NAND U7206 ( .A(n6906), .B(n6905), .Z(n6984) );
  XOR U7207 ( .A(n6985), .B(n6984), .Z(n6987) );
  XOR U7208 ( .A(n6986), .B(n6987), .Z(n6997) );
  NANDN U7209 ( .A(n6908), .B(n6907), .Z(n6912) );
  OR U7210 ( .A(n6910), .B(n6909), .Z(n6911) );
  AND U7211 ( .A(n6912), .B(n6911), .Z(n6996) );
  XNOR U7212 ( .A(n6997), .B(n6996), .Z(n6998) );
  NANDN U7213 ( .A(n6914), .B(n6913), .Z(n6918) );
  NANDN U7214 ( .A(n6916), .B(n6915), .Z(n6917) );
  NAND U7215 ( .A(n6918), .B(n6917), .Z(n6999) );
  XNOR U7216 ( .A(n6998), .B(n6999), .Z(n6944) );
  XOR U7217 ( .A(n6945), .B(n6944), .Z(n7003) );
  NANDN U7218 ( .A(n6920), .B(n6919), .Z(n6924) );
  NANDN U7219 ( .A(n6922), .B(n6921), .Z(n6923) );
  AND U7220 ( .A(n6924), .B(n6923), .Z(n7002) );
  XNOR U7221 ( .A(n7003), .B(n7002), .Z(n7004) );
  XOR U7222 ( .A(n7005), .B(n7004), .Z(n6937) );
  NANDN U7223 ( .A(n6926), .B(n6925), .Z(n6930) );
  NAND U7224 ( .A(n6928), .B(n6927), .Z(n6929) );
  AND U7225 ( .A(n6930), .B(n6929), .Z(n6936) );
  XNOR U7226 ( .A(n6937), .B(n6936), .Z(n6938) );
  XNOR U7227 ( .A(n6939), .B(n6938), .Z(n7008) );
  XNOR U7228 ( .A(sreg[337]), .B(n7008), .Z(n7010) );
  NANDN U7229 ( .A(sreg[336]), .B(n6931), .Z(n6935) );
  NAND U7230 ( .A(n6933), .B(n6932), .Z(n6934) );
  NAND U7231 ( .A(n6935), .B(n6934), .Z(n7009) );
  XNOR U7232 ( .A(n7010), .B(n7009), .Z(c[337]) );
  NANDN U7233 ( .A(n6937), .B(n6936), .Z(n6941) );
  NANDN U7234 ( .A(n6939), .B(n6938), .Z(n6940) );
  AND U7235 ( .A(n6941), .B(n6940), .Z(n7016) );
  NANDN U7236 ( .A(n6943), .B(n6942), .Z(n6947) );
  NAND U7237 ( .A(n6945), .B(n6944), .Z(n6946) );
  AND U7238 ( .A(n6947), .B(n6946), .Z(n7082) );
  NANDN U7239 ( .A(n6949), .B(n6948), .Z(n6953) );
  NANDN U7240 ( .A(n6951), .B(n6950), .Z(n6952) );
  AND U7241 ( .A(n6953), .B(n6952), .Z(n7069) );
  NAND U7242 ( .A(b[0]), .B(a[98]), .Z(n6954) );
  XNOR U7243 ( .A(b[1]), .B(n6954), .Z(n6956) );
  NANDN U7244 ( .A(b[0]), .B(a[97]), .Z(n6955) );
  NAND U7245 ( .A(n6956), .B(n6955), .Z(n7049) );
  NAND U7246 ( .A(n19808), .B(n6957), .Z(n6959) );
  XOR U7247 ( .A(b[13]), .B(a[86]), .Z(n7055) );
  NAND U7248 ( .A(n19768), .B(n7055), .Z(n6958) );
  AND U7249 ( .A(n6959), .B(n6958), .Z(n7047) );
  AND U7250 ( .A(b[15]), .B(a[82]), .Z(n7046) );
  XNOR U7251 ( .A(n7047), .B(n7046), .Z(n7048) );
  XNOR U7252 ( .A(n7049), .B(n7048), .Z(n7067) );
  NAND U7253 ( .A(n33), .B(n6960), .Z(n6962) );
  XOR U7254 ( .A(b[5]), .B(a[94]), .Z(n7058) );
  NAND U7255 ( .A(n19342), .B(n7058), .Z(n6961) );
  AND U7256 ( .A(n6962), .B(n6961), .Z(n7043) );
  NAND U7257 ( .A(n34), .B(n6963), .Z(n6965) );
  XOR U7258 ( .A(b[7]), .B(a[92]), .Z(n7061) );
  NAND U7259 ( .A(n19486), .B(n7061), .Z(n6964) );
  AND U7260 ( .A(n6965), .B(n6964), .Z(n7041) );
  NAND U7261 ( .A(n31), .B(n6966), .Z(n6968) );
  XOR U7262 ( .A(b[3]), .B(a[96]), .Z(n7064) );
  NAND U7263 ( .A(n32), .B(n7064), .Z(n6967) );
  NAND U7264 ( .A(n6968), .B(n6967), .Z(n7040) );
  XNOR U7265 ( .A(n7041), .B(n7040), .Z(n7042) );
  XOR U7266 ( .A(n7043), .B(n7042), .Z(n7068) );
  XOR U7267 ( .A(n7067), .B(n7068), .Z(n7070) );
  XOR U7268 ( .A(n7069), .B(n7070), .Z(n7020) );
  NANDN U7269 ( .A(n6970), .B(n6969), .Z(n6974) );
  OR U7270 ( .A(n6972), .B(n6971), .Z(n6973) );
  AND U7271 ( .A(n6974), .B(n6973), .Z(n7019) );
  XNOR U7272 ( .A(n7020), .B(n7019), .Z(n7022) );
  NAND U7273 ( .A(n6975), .B(n19724), .Z(n6977) );
  XOR U7274 ( .A(b[11]), .B(a[88]), .Z(n7025) );
  NAND U7275 ( .A(n19692), .B(n7025), .Z(n6976) );
  AND U7276 ( .A(n6977), .B(n6976), .Z(n7036) );
  NAND U7277 ( .A(n19838), .B(n6978), .Z(n6980) );
  XOR U7278 ( .A(b[15]), .B(a[84]), .Z(n7028) );
  NAND U7279 ( .A(n19805), .B(n7028), .Z(n6979) );
  AND U7280 ( .A(n6980), .B(n6979), .Z(n7035) );
  NAND U7281 ( .A(n35), .B(n6981), .Z(n6983) );
  XOR U7282 ( .A(b[9]), .B(a[90]), .Z(n7031) );
  NAND U7283 ( .A(n19598), .B(n7031), .Z(n6982) );
  NAND U7284 ( .A(n6983), .B(n6982), .Z(n7034) );
  XOR U7285 ( .A(n7035), .B(n7034), .Z(n7037) );
  XOR U7286 ( .A(n7036), .B(n7037), .Z(n7074) );
  NANDN U7287 ( .A(n6985), .B(n6984), .Z(n6989) );
  OR U7288 ( .A(n6987), .B(n6986), .Z(n6988) );
  AND U7289 ( .A(n6989), .B(n6988), .Z(n7073) );
  XNOR U7290 ( .A(n7074), .B(n7073), .Z(n7075) );
  NANDN U7291 ( .A(n6991), .B(n6990), .Z(n6995) );
  NANDN U7292 ( .A(n6993), .B(n6992), .Z(n6994) );
  NAND U7293 ( .A(n6995), .B(n6994), .Z(n7076) );
  XNOR U7294 ( .A(n7075), .B(n7076), .Z(n7021) );
  XOR U7295 ( .A(n7022), .B(n7021), .Z(n7080) );
  NANDN U7296 ( .A(n6997), .B(n6996), .Z(n7001) );
  NANDN U7297 ( .A(n6999), .B(n6998), .Z(n7000) );
  AND U7298 ( .A(n7001), .B(n7000), .Z(n7079) );
  XNOR U7299 ( .A(n7080), .B(n7079), .Z(n7081) );
  XOR U7300 ( .A(n7082), .B(n7081), .Z(n7014) );
  NANDN U7301 ( .A(n7003), .B(n7002), .Z(n7007) );
  NAND U7302 ( .A(n7005), .B(n7004), .Z(n7006) );
  AND U7303 ( .A(n7007), .B(n7006), .Z(n7013) );
  XNOR U7304 ( .A(n7014), .B(n7013), .Z(n7015) );
  XNOR U7305 ( .A(n7016), .B(n7015), .Z(n7085) );
  XNOR U7306 ( .A(sreg[338]), .B(n7085), .Z(n7087) );
  NANDN U7307 ( .A(sreg[337]), .B(n7008), .Z(n7012) );
  NAND U7308 ( .A(n7010), .B(n7009), .Z(n7011) );
  NAND U7309 ( .A(n7012), .B(n7011), .Z(n7086) );
  XNOR U7310 ( .A(n7087), .B(n7086), .Z(c[338]) );
  NANDN U7311 ( .A(n7014), .B(n7013), .Z(n7018) );
  NANDN U7312 ( .A(n7016), .B(n7015), .Z(n7017) );
  AND U7313 ( .A(n7018), .B(n7017), .Z(n7093) );
  NANDN U7314 ( .A(n7020), .B(n7019), .Z(n7024) );
  NAND U7315 ( .A(n7022), .B(n7021), .Z(n7023) );
  AND U7316 ( .A(n7024), .B(n7023), .Z(n7159) );
  NAND U7317 ( .A(n7025), .B(n19724), .Z(n7027) );
  XOR U7318 ( .A(b[11]), .B(a[89]), .Z(n7102) );
  NAND U7319 ( .A(n19692), .B(n7102), .Z(n7026) );
  AND U7320 ( .A(n7027), .B(n7026), .Z(n7113) );
  NAND U7321 ( .A(n19838), .B(n7028), .Z(n7030) );
  XOR U7322 ( .A(b[15]), .B(a[85]), .Z(n7105) );
  NAND U7323 ( .A(n19805), .B(n7105), .Z(n7029) );
  AND U7324 ( .A(n7030), .B(n7029), .Z(n7112) );
  NAND U7325 ( .A(n35), .B(n7031), .Z(n7033) );
  XOR U7326 ( .A(b[9]), .B(a[91]), .Z(n7108) );
  NAND U7327 ( .A(n19598), .B(n7108), .Z(n7032) );
  NAND U7328 ( .A(n7033), .B(n7032), .Z(n7111) );
  XOR U7329 ( .A(n7112), .B(n7111), .Z(n7114) );
  XOR U7330 ( .A(n7113), .B(n7114), .Z(n7151) );
  NANDN U7331 ( .A(n7035), .B(n7034), .Z(n7039) );
  OR U7332 ( .A(n7037), .B(n7036), .Z(n7038) );
  AND U7333 ( .A(n7039), .B(n7038), .Z(n7150) );
  XNOR U7334 ( .A(n7151), .B(n7150), .Z(n7152) );
  NANDN U7335 ( .A(n7041), .B(n7040), .Z(n7045) );
  NANDN U7336 ( .A(n7043), .B(n7042), .Z(n7044) );
  NAND U7337 ( .A(n7045), .B(n7044), .Z(n7153) );
  XNOR U7338 ( .A(n7152), .B(n7153), .Z(n7099) );
  NANDN U7339 ( .A(n7047), .B(n7046), .Z(n7051) );
  NANDN U7340 ( .A(n7049), .B(n7048), .Z(n7050) );
  AND U7341 ( .A(n7051), .B(n7050), .Z(n7146) );
  NAND U7342 ( .A(b[0]), .B(a[99]), .Z(n7052) );
  XNOR U7343 ( .A(b[1]), .B(n7052), .Z(n7054) );
  NANDN U7344 ( .A(b[0]), .B(a[98]), .Z(n7053) );
  NAND U7345 ( .A(n7054), .B(n7053), .Z(n7126) );
  NAND U7346 ( .A(n19808), .B(n7055), .Z(n7057) );
  XOR U7347 ( .A(b[13]), .B(a[87]), .Z(n7132) );
  NAND U7348 ( .A(n19768), .B(n7132), .Z(n7056) );
  AND U7349 ( .A(n7057), .B(n7056), .Z(n7124) );
  AND U7350 ( .A(b[15]), .B(a[83]), .Z(n7123) );
  XNOR U7351 ( .A(n7124), .B(n7123), .Z(n7125) );
  XNOR U7352 ( .A(n7126), .B(n7125), .Z(n7144) );
  NAND U7353 ( .A(n33), .B(n7058), .Z(n7060) );
  XOR U7354 ( .A(b[5]), .B(a[95]), .Z(n7135) );
  NAND U7355 ( .A(n19342), .B(n7135), .Z(n7059) );
  AND U7356 ( .A(n7060), .B(n7059), .Z(n7120) );
  NAND U7357 ( .A(n34), .B(n7061), .Z(n7063) );
  XOR U7358 ( .A(b[7]), .B(a[93]), .Z(n7138) );
  NAND U7359 ( .A(n19486), .B(n7138), .Z(n7062) );
  AND U7360 ( .A(n7063), .B(n7062), .Z(n7118) );
  NAND U7361 ( .A(n31), .B(n7064), .Z(n7066) );
  XOR U7362 ( .A(b[3]), .B(a[97]), .Z(n7141) );
  NAND U7363 ( .A(n32), .B(n7141), .Z(n7065) );
  NAND U7364 ( .A(n7066), .B(n7065), .Z(n7117) );
  XNOR U7365 ( .A(n7118), .B(n7117), .Z(n7119) );
  XOR U7366 ( .A(n7120), .B(n7119), .Z(n7145) );
  XOR U7367 ( .A(n7144), .B(n7145), .Z(n7147) );
  XOR U7368 ( .A(n7146), .B(n7147), .Z(n7097) );
  NANDN U7369 ( .A(n7068), .B(n7067), .Z(n7072) );
  OR U7370 ( .A(n7070), .B(n7069), .Z(n7071) );
  AND U7371 ( .A(n7072), .B(n7071), .Z(n7096) );
  XNOR U7372 ( .A(n7097), .B(n7096), .Z(n7098) );
  XOR U7373 ( .A(n7099), .B(n7098), .Z(n7157) );
  NANDN U7374 ( .A(n7074), .B(n7073), .Z(n7078) );
  NANDN U7375 ( .A(n7076), .B(n7075), .Z(n7077) );
  AND U7376 ( .A(n7078), .B(n7077), .Z(n7156) );
  XNOR U7377 ( .A(n7157), .B(n7156), .Z(n7158) );
  XOR U7378 ( .A(n7159), .B(n7158), .Z(n7091) );
  NANDN U7379 ( .A(n7080), .B(n7079), .Z(n7084) );
  NAND U7380 ( .A(n7082), .B(n7081), .Z(n7083) );
  AND U7381 ( .A(n7084), .B(n7083), .Z(n7090) );
  XNOR U7382 ( .A(n7091), .B(n7090), .Z(n7092) );
  XNOR U7383 ( .A(n7093), .B(n7092), .Z(n7162) );
  XNOR U7384 ( .A(sreg[339]), .B(n7162), .Z(n7164) );
  NANDN U7385 ( .A(sreg[338]), .B(n7085), .Z(n7089) );
  NAND U7386 ( .A(n7087), .B(n7086), .Z(n7088) );
  NAND U7387 ( .A(n7089), .B(n7088), .Z(n7163) );
  XNOR U7388 ( .A(n7164), .B(n7163), .Z(c[339]) );
  NANDN U7389 ( .A(n7091), .B(n7090), .Z(n7095) );
  NANDN U7390 ( .A(n7093), .B(n7092), .Z(n7094) );
  AND U7391 ( .A(n7095), .B(n7094), .Z(n7170) );
  NANDN U7392 ( .A(n7097), .B(n7096), .Z(n7101) );
  NAND U7393 ( .A(n7099), .B(n7098), .Z(n7100) );
  AND U7394 ( .A(n7101), .B(n7100), .Z(n7236) );
  NAND U7395 ( .A(n7102), .B(n19724), .Z(n7104) );
  XOR U7396 ( .A(b[11]), .B(a[90]), .Z(n7206) );
  NAND U7397 ( .A(n19692), .B(n7206), .Z(n7103) );
  AND U7398 ( .A(n7104), .B(n7103), .Z(n7217) );
  NAND U7399 ( .A(n19838), .B(n7105), .Z(n7107) );
  XOR U7400 ( .A(b[15]), .B(a[86]), .Z(n7209) );
  NAND U7401 ( .A(n19805), .B(n7209), .Z(n7106) );
  AND U7402 ( .A(n7107), .B(n7106), .Z(n7216) );
  NAND U7403 ( .A(n35), .B(n7108), .Z(n7110) );
  XOR U7404 ( .A(b[9]), .B(a[92]), .Z(n7212) );
  NAND U7405 ( .A(n19598), .B(n7212), .Z(n7109) );
  NAND U7406 ( .A(n7110), .B(n7109), .Z(n7215) );
  XOR U7407 ( .A(n7216), .B(n7215), .Z(n7218) );
  XOR U7408 ( .A(n7217), .B(n7218), .Z(n7228) );
  NANDN U7409 ( .A(n7112), .B(n7111), .Z(n7116) );
  OR U7410 ( .A(n7114), .B(n7113), .Z(n7115) );
  AND U7411 ( .A(n7116), .B(n7115), .Z(n7227) );
  XNOR U7412 ( .A(n7228), .B(n7227), .Z(n7229) );
  NANDN U7413 ( .A(n7118), .B(n7117), .Z(n7122) );
  NANDN U7414 ( .A(n7120), .B(n7119), .Z(n7121) );
  NAND U7415 ( .A(n7122), .B(n7121), .Z(n7230) );
  XNOR U7416 ( .A(n7229), .B(n7230), .Z(n7176) );
  NANDN U7417 ( .A(n7124), .B(n7123), .Z(n7128) );
  NANDN U7418 ( .A(n7126), .B(n7125), .Z(n7127) );
  AND U7419 ( .A(n7128), .B(n7127), .Z(n7202) );
  NAND U7420 ( .A(b[0]), .B(a[100]), .Z(n7129) );
  XNOR U7421 ( .A(b[1]), .B(n7129), .Z(n7131) );
  NANDN U7422 ( .A(b[0]), .B(a[99]), .Z(n7130) );
  NAND U7423 ( .A(n7131), .B(n7130), .Z(n7182) );
  NAND U7424 ( .A(n19808), .B(n7132), .Z(n7134) );
  XOR U7425 ( .A(b[13]), .B(a[88]), .Z(n7188) );
  NAND U7426 ( .A(n19768), .B(n7188), .Z(n7133) );
  AND U7427 ( .A(n7134), .B(n7133), .Z(n7180) );
  AND U7428 ( .A(b[15]), .B(a[84]), .Z(n7179) );
  XNOR U7429 ( .A(n7180), .B(n7179), .Z(n7181) );
  XNOR U7430 ( .A(n7182), .B(n7181), .Z(n7200) );
  NAND U7431 ( .A(n33), .B(n7135), .Z(n7137) );
  XOR U7432 ( .A(b[5]), .B(a[96]), .Z(n7191) );
  NAND U7433 ( .A(n19342), .B(n7191), .Z(n7136) );
  AND U7434 ( .A(n7137), .B(n7136), .Z(n7224) );
  NAND U7435 ( .A(n34), .B(n7138), .Z(n7140) );
  XOR U7436 ( .A(b[7]), .B(a[94]), .Z(n7194) );
  NAND U7437 ( .A(n19486), .B(n7194), .Z(n7139) );
  AND U7438 ( .A(n7140), .B(n7139), .Z(n7222) );
  NAND U7439 ( .A(n31), .B(n7141), .Z(n7143) );
  XOR U7440 ( .A(b[3]), .B(a[98]), .Z(n7197) );
  NAND U7441 ( .A(n32), .B(n7197), .Z(n7142) );
  NAND U7442 ( .A(n7143), .B(n7142), .Z(n7221) );
  XNOR U7443 ( .A(n7222), .B(n7221), .Z(n7223) );
  XOR U7444 ( .A(n7224), .B(n7223), .Z(n7201) );
  XOR U7445 ( .A(n7200), .B(n7201), .Z(n7203) );
  XOR U7446 ( .A(n7202), .B(n7203), .Z(n7174) );
  NANDN U7447 ( .A(n7145), .B(n7144), .Z(n7149) );
  OR U7448 ( .A(n7147), .B(n7146), .Z(n7148) );
  AND U7449 ( .A(n7149), .B(n7148), .Z(n7173) );
  XNOR U7450 ( .A(n7174), .B(n7173), .Z(n7175) );
  XOR U7451 ( .A(n7176), .B(n7175), .Z(n7234) );
  NANDN U7452 ( .A(n7151), .B(n7150), .Z(n7155) );
  NANDN U7453 ( .A(n7153), .B(n7152), .Z(n7154) );
  AND U7454 ( .A(n7155), .B(n7154), .Z(n7233) );
  XNOR U7455 ( .A(n7234), .B(n7233), .Z(n7235) );
  XOR U7456 ( .A(n7236), .B(n7235), .Z(n7168) );
  NANDN U7457 ( .A(n7157), .B(n7156), .Z(n7161) );
  NAND U7458 ( .A(n7159), .B(n7158), .Z(n7160) );
  AND U7459 ( .A(n7161), .B(n7160), .Z(n7167) );
  XNOR U7460 ( .A(n7168), .B(n7167), .Z(n7169) );
  XNOR U7461 ( .A(n7170), .B(n7169), .Z(n7239) );
  XNOR U7462 ( .A(sreg[340]), .B(n7239), .Z(n7241) );
  NANDN U7463 ( .A(sreg[339]), .B(n7162), .Z(n7166) );
  NAND U7464 ( .A(n7164), .B(n7163), .Z(n7165) );
  NAND U7465 ( .A(n7166), .B(n7165), .Z(n7240) );
  XNOR U7466 ( .A(n7241), .B(n7240), .Z(c[340]) );
  NANDN U7467 ( .A(n7168), .B(n7167), .Z(n7172) );
  NANDN U7468 ( .A(n7170), .B(n7169), .Z(n7171) );
  AND U7469 ( .A(n7172), .B(n7171), .Z(n7247) );
  NANDN U7470 ( .A(n7174), .B(n7173), .Z(n7178) );
  NAND U7471 ( .A(n7176), .B(n7175), .Z(n7177) );
  AND U7472 ( .A(n7178), .B(n7177), .Z(n7313) );
  NANDN U7473 ( .A(n7180), .B(n7179), .Z(n7184) );
  NANDN U7474 ( .A(n7182), .B(n7181), .Z(n7183) );
  AND U7475 ( .A(n7184), .B(n7183), .Z(n7279) );
  NAND U7476 ( .A(b[0]), .B(a[101]), .Z(n7185) );
  XNOR U7477 ( .A(b[1]), .B(n7185), .Z(n7187) );
  NANDN U7478 ( .A(b[0]), .B(a[100]), .Z(n7186) );
  NAND U7479 ( .A(n7187), .B(n7186), .Z(n7259) );
  NAND U7480 ( .A(n19808), .B(n7188), .Z(n7190) );
  XOR U7481 ( .A(b[13]), .B(a[89]), .Z(n7262) );
  NAND U7482 ( .A(n19768), .B(n7262), .Z(n7189) );
  AND U7483 ( .A(n7190), .B(n7189), .Z(n7257) );
  AND U7484 ( .A(b[15]), .B(a[85]), .Z(n7256) );
  XNOR U7485 ( .A(n7257), .B(n7256), .Z(n7258) );
  XNOR U7486 ( .A(n7259), .B(n7258), .Z(n7277) );
  NAND U7487 ( .A(n33), .B(n7191), .Z(n7193) );
  XOR U7488 ( .A(b[5]), .B(a[97]), .Z(n7268) );
  NAND U7489 ( .A(n19342), .B(n7268), .Z(n7192) );
  AND U7490 ( .A(n7193), .B(n7192), .Z(n7301) );
  NAND U7491 ( .A(n34), .B(n7194), .Z(n7196) );
  XOR U7492 ( .A(b[7]), .B(a[95]), .Z(n7271) );
  NAND U7493 ( .A(n19486), .B(n7271), .Z(n7195) );
  AND U7494 ( .A(n7196), .B(n7195), .Z(n7299) );
  NAND U7495 ( .A(n31), .B(n7197), .Z(n7199) );
  XOR U7496 ( .A(b[3]), .B(a[99]), .Z(n7274) );
  NAND U7497 ( .A(n32), .B(n7274), .Z(n7198) );
  NAND U7498 ( .A(n7199), .B(n7198), .Z(n7298) );
  XNOR U7499 ( .A(n7299), .B(n7298), .Z(n7300) );
  XOR U7500 ( .A(n7301), .B(n7300), .Z(n7278) );
  XOR U7501 ( .A(n7277), .B(n7278), .Z(n7280) );
  XOR U7502 ( .A(n7279), .B(n7280), .Z(n7251) );
  NANDN U7503 ( .A(n7201), .B(n7200), .Z(n7205) );
  OR U7504 ( .A(n7203), .B(n7202), .Z(n7204) );
  AND U7505 ( .A(n7205), .B(n7204), .Z(n7250) );
  XNOR U7506 ( .A(n7251), .B(n7250), .Z(n7253) );
  NAND U7507 ( .A(n7206), .B(n19724), .Z(n7208) );
  XOR U7508 ( .A(b[11]), .B(a[91]), .Z(n7283) );
  NAND U7509 ( .A(n19692), .B(n7283), .Z(n7207) );
  AND U7510 ( .A(n7208), .B(n7207), .Z(n7294) );
  NAND U7511 ( .A(n19838), .B(n7209), .Z(n7211) );
  XOR U7512 ( .A(b[15]), .B(a[87]), .Z(n7286) );
  NAND U7513 ( .A(n19805), .B(n7286), .Z(n7210) );
  AND U7514 ( .A(n7211), .B(n7210), .Z(n7293) );
  NAND U7515 ( .A(n35), .B(n7212), .Z(n7214) );
  XOR U7516 ( .A(b[9]), .B(a[93]), .Z(n7289) );
  NAND U7517 ( .A(n19598), .B(n7289), .Z(n7213) );
  NAND U7518 ( .A(n7214), .B(n7213), .Z(n7292) );
  XOR U7519 ( .A(n7293), .B(n7292), .Z(n7295) );
  XOR U7520 ( .A(n7294), .B(n7295), .Z(n7305) );
  NANDN U7521 ( .A(n7216), .B(n7215), .Z(n7220) );
  OR U7522 ( .A(n7218), .B(n7217), .Z(n7219) );
  AND U7523 ( .A(n7220), .B(n7219), .Z(n7304) );
  XNOR U7524 ( .A(n7305), .B(n7304), .Z(n7306) );
  NANDN U7525 ( .A(n7222), .B(n7221), .Z(n7226) );
  NANDN U7526 ( .A(n7224), .B(n7223), .Z(n7225) );
  NAND U7527 ( .A(n7226), .B(n7225), .Z(n7307) );
  XNOR U7528 ( .A(n7306), .B(n7307), .Z(n7252) );
  XOR U7529 ( .A(n7253), .B(n7252), .Z(n7311) );
  NANDN U7530 ( .A(n7228), .B(n7227), .Z(n7232) );
  NANDN U7531 ( .A(n7230), .B(n7229), .Z(n7231) );
  AND U7532 ( .A(n7232), .B(n7231), .Z(n7310) );
  XNOR U7533 ( .A(n7311), .B(n7310), .Z(n7312) );
  XOR U7534 ( .A(n7313), .B(n7312), .Z(n7245) );
  NANDN U7535 ( .A(n7234), .B(n7233), .Z(n7238) );
  NAND U7536 ( .A(n7236), .B(n7235), .Z(n7237) );
  AND U7537 ( .A(n7238), .B(n7237), .Z(n7244) );
  XNOR U7538 ( .A(n7245), .B(n7244), .Z(n7246) );
  XNOR U7539 ( .A(n7247), .B(n7246), .Z(n7316) );
  XNOR U7540 ( .A(sreg[341]), .B(n7316), .Z(n7318) );
  NANDN U7541 ( .A(sreg[340]), .B(n7239), .Z(n7243) );
  NAND U7542 ( .A(n7241), .B(n7240), .Z(n7242) );
  NAND U7543 ( .A(n7243), .B(n7242), .Z(n7317) );
  XNOR U7544 ( .A(n7318), .B(n7317), .Z(c[341]) );
  NANDN U7545 ( .A(n7245), .B(n7244), .Z(n7249) );
  NANDN U7546 ( .A(n7247), .B(n7246), .Z(n7248) );
  AND U7547 ( .A(n7249), .B(n7248), .Z(n7324) );
  NANDN U7548 ( .A(n7251), .B(n7250), .Z(n7255) );
  NAND U7549 ( .A(n7253), .B(n7252), .Z(n7254) );
  AND U7550 ( .A(n7255), .B(n7254), .Z(n7390) );
  NANDN U7551 ( .A(n7257), .B(n7256), .Z(n7261) );
  NANDN U7552 ( .A(n7259), .B(n7258), .Z(n7260) );
  AND U7553 ( .A(n7261), .B(n7260), .Z(n7356) );
  NAND U7554 ( .A(n19808), .B(n7262), .Z(n7264) );
  XOR U7555 ( .A(b[13]), .B(a[90]), .Z(n7339) );
  NAND U7556 ( .A(n19768), .B(n7339), .Z(n7263) );
  AND U7557 ( .A(n7264), .B(n7263), .Z(n7334) );
  AND U7558 ( .A(b[15]), .B(a[86]), .Z(n7333) );
  XNOR U7559 ( .A(n7334), .B(n7333), .Z(n7335) );
  NAND U7560 ( .A(b[0]), .B(a[102]), .Z(n7265) );
  XNOR U7561 ( .A(b[1]), .B(n7265), .Z(n7267) );
  NANDN U7562 ( .A(b[0]), .B(a[101]), .Z(n7266) );
  NAND U7563 ( .A(n7267), .B(n7266), .Z(n7336) );
  XNOR U7564 ( .A(n7335), .B(n7336), .Z(n7354) );
  NAND U7565 ( .A(n33), .B(n7268), .Z(n7270) );
  XOR U7566 ( .A(b[5]), .B(a[98]), .Z(n7345) );
  NAND U7567 ( .A(n19342), .B(n7345), .Z(n7269) );
  AND U7568 ( .A(n7270), .B(n7269), .Z(n7378) );
  NAND U7569 ( .A(n34), .B(n7271), .Z(n7273) );
  XOR U7570 ( .A(b[7]), .B(a[96]), .Z(n7348) );
  NAND U7571 ( .A(n19486), .B(n7348), .Z(n7272) );
  AND U7572 ( .A(n7273), .B(n7272), .Z(n7376) );
  NAND U7573 ( .A(n31), .B(n7274), .Z(n7276) );
  XOR U7574 ( .A(b[3]), .B(a[100]), .Z(n7351) );
  NAND U7575 ( .A(n32), .B(n7351), .Z(n7275) );
  NAND U7576 ( .A(n7276), .B(n7275), .Z(n7375) );
  XNOR U7577 ( .A(n7376), .B(n7375), .Z(n7377) );
  XOR U7578 ( .A(n7378), .B(n7377), .Z(n7355) );
  XOR U7579 ( .A(n7354), .B(n7355), .Z(n7357) );
  XOR U7580 ( .A(n7356), .B(n7357), .Z(n7328) );
  NANDN U7581 ( .A(n7278), .B(n7277), .Z(n7282) );
  OR U7582 ( .A(n7280), .B(n7279), .Z(n7281) );
  AND U7583 ( .A(n7282), .B(n7281), .Z(n7327) );
  XNOR U7584 ( .A(n7328), .B(n7327), .Z(n7330) );
  NAND U7585 ( .A(n7283), .B(n19724), .Z(n7285) );
  XOR U7586 ( .A(b[11]), .B(a[92]), .Z(n7360) );
  NAND U7587 ( .A(n19692), .B(n7360), .Z(n7284) );
  AND U7588 ( .A(n7285), .B(n7284), .Z(n7371) );
  NAND U7589 ( .A(n19838), .B(n7286), .Z(n7288) );
  XOR U7590 ( .A(b[15]), .B(a[88]), .Z(n7363) );
  NAND U7591 ( .A(n19805), .B(n7363), .Z(n7287) );
  AND U7592 ( .A(n7288), .B(n7287), .Z(n7370) );
  NAND U7593 ( .A(n35), .B(n7289), .Z(n7291) );
  XOR U7594 ( .A(b[9]), .B(a[94]), .Z(n7366) );
  NAND U7595 ( .A(n19598), .B(n7366), .Z(n7290) );
  NAND U7596 ( .A(n7291), .B(n7290), .Z(n7369) );
  XOR U7597 ( .A(n7370), .B(n7369), .Z(n7372) );
  XOR U7598 ( .A(n7371), .B(n7372), .Z(n7382) );
  NANDN U7599 ( .A(n7293), .B(n7292), .Z(n7297) );
  OR U7600 ( .A(n7295), .B(n7294), .Z(n7296) );
  AND U7601 ( .A(n7297), .B(n7296), .Z(n7381) );
  XNOR U7602 ( .A(n7382), .B(n7381), .Z(n7383) );
  NANDN U7603 ( .A(n7299), .B(n7298), .Z(n7303) );
  NANDN U7604 ( .A(n7301), .B(n7300), .Z(n7302) );
  NAND U7605 ( .A(n7303), .B(n7302), .Z(n7384) );
  XNOR U7606 ( .A(n7383), .B(n7384), .Z(n7329) );
  XOR U7607 ( .A(n7330), .B(n7329), .Z(n7388) );
  NANDN U7608 ( .A(n7305), .B(n7304), .Z(n7309) );
  NANDN U7609 ( .A(n7307), .B(n7306), .Z(n7308) );
  AND U7610 ( .A(n7309), .B(n7308), .Z(n7387) );
  XNOR U7611 ( .A(n7388), .B(n7387), .Z(n7389) );
  XOR U7612 ( .A(n7390), .B(n7389), .Z(n7322) );
  NANDN U7613 ( .A(n7311), .B(n7310), .Z(n7315) );
  NAND U7614 ( .A(n7313), .B(n7312), .Z(n7314) );
  AND U7615 ( .A(n7315), .B(n7314), .Z(n7321) );
  XNOR U7616 ( .A(n7322), .B(n7321), .Z(n7323) );
  XNOR U7617 ( .A(n7324), .B(n7323), .Z(n7393) );
  XNOR U7618 ( .A(sreg[342]), .B(n7393), .Z(n7395) );
  NANDN U7619 ( .A(sreg[341]), .B(n7316), .Z(n7320) );
  NAND U7620 ( .A(n7318), .B(n7317), .Z(n7319) );
  NAND U7621 ( .A(n7320), .B(n7319), .Z(n7394) );
  XNOR U7622 ( .A(n7395), .B(n7394), .Z(c[342]) );
  NANDN U7623 ( .A(n7322), .B(n7321), .Z(n7326) );
  NANDN U7624 ( .A(n7324), .B(n7323), .Z(n7325) );
  AND U7625 ( .A(n7326), .B(n7325), .Z(n7401) );
  NANDN U7626 ( .A(n7328), .B(n7327), .Z(n7332) );
  NAND U7627 ( .A(n7330), .B(n7329), .Z(n7331) );
  AND U7628 ( .A(n7332), .B(n7331), .Z(n7467) );
  NANDN U7629 ( .A(n7334), .B(n7333), .Z(n7338) );
  NANDN U7630 ( .A(n7336), .B(n7335), .Z(n7337) );
  AND U7631 ( .A(n7338), .B(n7337), .Z(n7433) );
  NAND U7632 ( .A(n19808), .B(n7339), .Z(n7341) );
  XOR U7633 ( .A(b[13]), .B(a[91]), .Z(n7416) );
  NAND U7634 ( .A(n19768), .B(n7416), .Z(n7340) );
  AND U7635 ( .A(n7341), .B(n7340), .Z(n7411) );
  AND U7636 ( .A(b[15]), .B(a[87]), .Z(n7410) );
  XNOR U7637 ( .A(n7411), .B(n7410), .Z(n7412) );
  NAND U7638 ( .A(b[0]), .B(a[103]), .Z(n7342) );
  XNOR U7639 ( .A(b[1]), .B(n7342), .Z(n7344) );
  NANDN U7640 ( .A(b[0]), .B(a[102]), .Z(n7343) );
  NAND U7641 ( .A(n7344), .B(n7343), .Z(n7413) );
  XNOR U7642 ( .A(n7412), .B(n7413), .Z(n7431) );
  NAND U7643 ( .A(n33), .B(n7345), .Z(n7347) );
  XOR U7644 ( .A(b[5]), .B(a[99]), .Z(n7422) );
  NAND U7645 ( .A(n19342), .B(n7422), .Z(n7346) );
  AND U7646 ( .A(n7347), .B(n7346), .Z(n7455) );
  NAND U7647 ( .A(n34), .B(n7348), .Z(n7350) );
  XOR U7648 ( .A(b[7]), .B(a[97]), .Z(n7425) );
  NAND U7649 ( .A(n19486), .B(n7425), .Z(n7349) );
  AND U7650 ( .A(n7350), .B(n7349), .Z(n7453) );
  NAND U7651 ( .A(n31), .B(n7351), .Z(n7353) );
  XOR U7652 ( .A(b[3]), .B(a[101]), .Z(n7428) );
  NAND U7653 ( .A(n32), .B(n7428), .Z(n7352) );
  NAND U7654 ( .A(n7353), .B(n7352), .Z(n7452) );
  XNOR U7655 ( .A(n7453), .B(n7452), .Z(n7454) );
  XOR U7656 ( .A(n7455), .B(n7454), .Z(n7432) );
  XOR U7657 ( .A(n7431), .B(n7432), .Z(n7434) );
  XOR U7658 ( .A(n7433), .B(n7434), .Z(n7405) );
  NANDN U7659 ( .A(n7355), .B(n7354), .Z(n7359) );
  OR U7660 ( .A(n7357), .B(n7356), .Z(n7358) );
  AND U7661 ( .A(n7359), .B(n7358), .Z(n7404) );
  XNOR U7662 ( .A(n7405), .B(n7404), .Z(n7407) );
  NAND U7663 ( .A(n7360), .B(n19724), .Z(n7362) );
  XOR U7664 ( .A(b[11]), .B(a[93]), .Z(n7437) );
  NAND U7665 ( .A(n19692), .B(n7437), .Z(n7361) );
  AND U7666 ( .A(n7362), .B(n7361), .Z(n7448) );
  NAND U7667 ( .A(n19838), .B(n7363), .Z(n7365) );
  XOR U7668 ( .A(b[15]), .B(a[89]), .Z(n7440) );
  NAND U7669 ( .A(n19805), .B(n7440), .Z(n7364) );
  AND U7670 ( .A(n7365), .B(n7364), .Z(n7447) );
  NAND U7671 ( .A(n35), .B(n7366), .Z(n7368) );
  XOR U7672 ( .A(b[9]), .B(a[95]), .Z(n7443) );
  NAND U7673 ( .A(n19598), .B(n7443), .Z(n7367) );
  NAND U7674 ( .A(n7368), .B(n7367), .Z(n7446) );
  XOR U7675 ( .A(n7447), .B(n7446), .Z(n7449) );
  XOR U7676 ( .A(n7448), .B(n7449), .Z(n7459) );
  NANDN U7677 ( .A(n7370), .B(n7369), .Z(n7374) );
  OR U7678 ( .A(n7372), .B(n7371), .Z(n7373) );
  AND U7679 ( .A(n7374), .B(n7373), .Z(n7458) );
  XNOR U7680 ( .A(n7459), .B(n7458), .Z(n7460) );
  NANDN U7681 ( .A(n7376), .B(n7375), .Z(n7380) );
  NANDN U7682 ( .A(n7378), .B(n7377), .Z(n7379) );
  NAND U7683 ( .A(n7380), .B(n7379), .Z(n7461) );
  XNOR U7684 ( .A(n7460), .B(n7461), .Z(n7406) );
  XOR U7685 ( .A(n7407), .B(n7406), .Z(n7465) );
  NANDN U7686 ( .A(n7382), .B(n7381), .Z(n7386) );
  NANDN U7687 ( .A(n7384), .B(n7383), .Z(n7385) );
  AND U7688 ( .A(n7386), .B(n7385), .Z(n7464) );
  XNOR U7689 ( .A(n7465), .B(n7464), .Z(n7466) );
  XOR U7690 ( .A(n7467), .B(n7466), .Z(n7399) );
  NANDN U7691 ( .A(n7388), .B(n7387), .Z(n7392) );
  NAND U7692 ( .A(n7390), .B(n7389), .Z(n7391) );
  AND U7693 ( .A(n7392), .B(n7391), .Z(n7398) );
  XNOR U7694 ( .A(n7399), .B(n7398), .Z(n7400) );
  XNOR U7695 ( .A(n7401), .B(n7400), .Z(n7470) );
  XNOR U7696 ( .A(sreg[343]), .B(n7470), .Z(n7472) );
  NANDN U7697 ( .A(sreg[342]), .B(n7393), .Z(n7397) );
  NAND U7698 ( .A(n7395), .B(n7394), .Z(n7396) );
  NAND U7699 ( .A(n7397), .B(n7396), .Z(n7471) );
  XNOR U7700 ( .A(n7472), .B(n7471), .Z(c[343]) );
  NANDN U7701 ( .A(n7399), .B(n7398), .Z(n7403) );
  NANDN U7702 ( .A(n7401), .B(n7400), .Z(n7402) );
  AND U7703 ( .A(n7403), .B(n7402), .Z(n7478) );
  NANDN U7704 ( .A(n7405), .B(n7404), .Z(n7409) );
  NAND U7705 ( .A(n7407), .B(n7406), .Z(n7408) );
  AND U7706 ( .A(n7409), .B(n7408), .Z(n7544) );
  NANDN U7707 ( .A(n7411), .B(n7410), .Z(n7415) );
  NANDN U7708 ( .A(n7413), .B(n7412), .Z(n7414) );
  AND U7709 ( .A(n7415), .B(n7414), .Z(n7510) );
  NAND U7710 ( .A(n19808), .B(n7416), .Z(n7418) );
  XOR U7711 ( .A(b[13]), .B(a[92]), .Z(n7496) );
  NAND U7712 ( .A(n19768), .B(n7496), .Z(n7417) );
  AND U7713 ( .A(n7418), .B(n7417), .Z(n7488) );
  AND U7714 ( .A(b[15]), .B(a[88]), .Z(n7487) );
  XNOR U7715 ( .A(n7488), .B(n7487), .Z(n7489) );
  NAND U7716 ( .A(b[0]), .B(a[104]), .Z(n7419) );
  XNOR U7717 ( .A(b[1]), .B(n7419), .Z(n7421) );
  NANDN U7718 ( .A(b[0]), .B(a[103]), .Z(n7420) );
  NAND U7719 ( .A(n7421), .B(n7420), .Z(n7490) );
  XNOR U7720 ( .A(n7489), .B(n7490), .Z(n7508) );
  NAND U7721 ( .A(n33), .B(n7422), .Z(n7424) );
  XOR U7722 ( .A(b[5]), .B(a[100]), .Z(n7499) );
  NAND U7723 ( .A(n19342), .B(n7499), .Z(n7423) );
  AND U7724 ( .A(n7424), .B(n7423), .Z(n7532) );
  NAND U7725 ( .A(n34), .B(n7425), .Z(n7427) );
  XOR U7726 ( .A(b[7]), .B(a[98]), .Z(n7502) );
  NAND U7727 ( .A(n19486), .B(n7502), .Z(n7426) );
  AND U7728 ( .A(n7427), .B(n7426), .Z(n7530) );
  NAND U7729 ( .A(n31), .B(n7428), .Z(n7430) );
  XOR U7730 ( .A(b[3]), .B(a[102]), .Z(n7505) );
  NAND U7731 ( .A(n32), .B(n7505), .Z(n7429) );
  NAND U7732 ( .A(n7430), .B(n7429), .Z(n7529) );
  XNOR U7733 ( .A(n7530), .B(n7529), .Z(n7531) );
  XOR U7734 ( .A(n7532), .B(n7531), .Z(n7509) );
  XOR U7735 ( .A(n7508), .B(n7509), .Z(n7511) );
  XOR U7736 ( .A(n7510), .B(n7511), .Z(n7482) );
  NANDN U7737 ( .A(n7432), .B(n7431), .Z(n7436) );
  OR U7738 ( .A(n7434), .B(n7433), .Z(n7435) );
  AND U7739 ( .A(n7436), .B(n7435), .Z(n7481) );
  XNOR U7740 ( .A(n7482), .B(n7481), .Z(n7484) );
  NAND U7741 ( .A(n7437), .B(n19724), .Z(n7439) );
  XOR U7742 ( .A(b[11]), .B(a[94]), .Z(n7514) );
  NAND U7743 ( .A(n19692), .B(n7514), .Z(n7438) );
  AND U7744 ( .A(n7439), .B(n7438), .Z(n7525) );
  NAND U7745 ( .A(n19838), .B(n7440), .Z(n7442) );
  XOR U7746 ( .A(b[15]), .B(a[90]), .Z(n7517) );
  NAND U7747 ( .A(n19805), .B(n7517), .Z(n7441) );
  AND U7748 ( .A(n7442), .B(n7441), .Z(n7524) );
  NAND U7749 ( .A(n35), .B(n7443), .Z(n7445) );
  XOR U7750 ( .A(b[9]), .B(a[96]), .Z(n7520) );
  NAND U7751 ( .A(n19598), .B(n7520), .Z(n7444) );
  NAND U7752 ( .A(n7445), .B(n7444), .Z(n7523) );
  XOR U7753 ( .A(n7524), .B(n7523), .Z(n7526) );
  XOR U7754 ( .A(n7525), .B(n7526), .Z(n7536) );
  NANDN U7755 ( .A(n7447), .B(n7446), .Z(n7451) );
  OR U7756 ( .A(n7449), .B(n7448), .Z(n7450) );
  AND U7757 ( .A(n7451), .B(n7450), .Z(n7535) );
  XNOR U7758 ( .A(n7536), .B(n7535), .Z(n7537) );
  NANDN U7759 ( .A(n7453), .B(n7452), .Z(n7457) );
  NANDN U7760 ( .A(n7455), .B(n7454), .Z(n7456) );
  NAND U7761 ( .A(n7457), .B(n7456), .Z(n7538) );
  XNOR U7762 ( .A(n7537), .B(n7538), .Z(n7483) );
  XOR U7763 ( .A(n7484), .B(n7483), .Z(n7542) );
  NANDN U7764 ( .A(n7459), .B(n7458), .Z(n7463) );
  NANDN U7765 ( .A(n7461), .B(n7460), .Z(n7462) );
  AND U7766 ( .A(n7463), .B(n7462), .Z(n7541) );
  XNOR U7767 ( .A(n7542), .B(n7541), .Z(n7543) );
  XOR U7768 ( .A(n7544), .B(n7543), .Z(n7476) );
  NANDN U7769 ( .A(n7465), .B(n7464), .Z(n7469) );
  NAND U7770 ( .A(n7467), .B(n7466), .Z(n7468) );
  AND U7771 ( .A(n7469), .B(n7468), .Z(n7475) );
  XNOR U7772 ( .A(n7476), .B(n7475), .Z(n7477) );
  XNOR U7773 ( .A(n7478), .B(n7477), .Z(n7547) );
  XNOR U7774 ( .A(sreg[344]), .B(n7547), .Z(n7549) );
  NANDN U7775 ( .A(sreg[343]), .B(n7470), .Z(n7474) );
  NAND U7776 ( .A(n7472), .B(n7471), .Z(n7473) );
  NAND U7777 ( .A(n7474), .B(n7473), .Z(n7548) );
  XNOR U7778 ( .A(n7549), .B(n7548), .Z(c[344]) );
  NANDN U7779 ( .A(n7476), .B(n7475), .Z(n7480) );
  NANDN U7780 ( .A(n7478), .B(n7477), .Z(n7479) );
  AND U7781 ( .A(n7480), .B(n7479), .Z(n7555) );
  NANDN U7782 ( .A(n7482), .B(n7481), .Z(n7486) );
  NAND U7783 ( .A(n7484), .B(n7483), .Z(n7485) );
  AND U7784 ( .A(n7486), .B(n7485), .Z(n7621) );
  NANDN U7785 ( .A(n7488), .B(n7487), .Z(n7492) );
  NANDN U7786 ( .A(n7490), .B(n7489), .Z(n7491) );
  AND U7787 ( .A(n7492), .B(n7491), .Z(n7608) );
  NAND U7788 ( .A(b[0]), .B(a[105]), .Z(n7493) );
  XNOR U7789 ( .A(b[1]), .B(n7493), .Z(n7495) );
  NANDN U7790 ( .A(b[0]), .B(a[104]), .Z(n7494) );
  NAND U7791 ( .A(n7495), .B(n7494), .Z(n7588) );
  NAND U7792 ( .A(n19808), .B(n7496), .Z(n7498) );
  XOR U7793 ( .A(b[13]), .B(a[93]), .Z(n7594) );
  NAND U7794 ( .A(n19768), .B(n7594), .Z(n7497) );
  AND U7795 ( .A(n7498), .B(n7497), .Z(n7586) );
  AND U7796 ( .A(b[15]), .B(a[89]), .Z(n7585) );
  XNOR U7797 ( .A(n7586), .B(n7585), .Z(n7587) );
  XNOR U7798 ( .A(n7588), .B(n7587), .Z(n7606) );
  NAND U7799 ( .A(n33), .B(n7499), .Z(n7501) );
  XOR U7800 ( .A(b[5]), .B(a[101]), .Z(n7597) );
  NAND U7801 ( .A(n19342), .B(n7597), .Z(n7500) );
  AND U7802 ( .A(n7501), .B(n7500), .Z(n7582) );
  NAND U7803 ( .A(n34), .B(n7502), .Z(n7504) );
  XOR U7804 ( .A(b[7]), .B(a[99]), .Z(n7600) );
  NAND U7805 ( .A(n19486), .B(n7600), .Z(n7503) );
  AND U7806 ( .A(n7504), .B(n7503), .Z(n7580) );
  NAND U7807 ( .A(n31), .B(n7505), .Z(n7507) );
  XOR U7808 ( .A(b[3]), .B(a[103]), .Z(n7603) );
  NAND U7809 ( .A(n32), .B(n7603), .Z(n7506) );
  NAND U7810 ( .A(n7507), .B(n7506), .Z(n7579) );
  XNOR U7811 ( .A(n7580), .B(n7579), .Z(n7581) );
  XOR U7812 ( .A(n7582), .B(n7581), .Z(n7607) );
  XOR U7813 ( .A(n7606), .B(n7607), .Z(n7609) );
  XOR U7814 ( .A(n7608), .B(n7609), .Z(n7559) );
  NANDN U7815 ( .A(n7509), .B(n7508), .Z(n7513) );
  OR U7816 ( .A(n7511), .B(n7510), .Z(n7512) );
  AND U7817 ( .A(n7513), .B(n7512), .Z(n7558) );
  XNOR U7818 ( .A(n7559), .B(n7558), .Z(n7561) );
  NAND U7819 ( .A(n7514), .B(n19724), .Z(n7516) );
  XOR U7820 ( .A(b[11]), .B(a[95]), .Z(n7564) );
  NAND U7821 ( .A(n19692), .B(n7564), .Z(n7515) );
  AND U7822 ( .A(n7516), .B(n7515), .Z(n7575) );
  NAND U7823 ( .A(n19838), .B(n7517), .Z(n7519) );
  XOR U7824 ( .A(b[15]), .B(a[91]), .Z(n7567) );
  NAND U7825 ( .A(n19805), .B(n7567), .Z(n7518) );
  AND U7826 ( .A(n7519), .B(n7518), .Z(n7574) );
  NAND U7827 ( .A(n35), .B(n7520), .Z(n7522) );
  XOR U7828 ( .A(b[9]), .B(a[97]), .Z(n7570) );
  NAND U7829 ( .A(n19598), .B(n7570), .Z(n7521) );
  NAND U7830 ( .A(n7522), .B(n7521), .Z(n7573) );
  XOR U7831 ( .A(n7574), .B(n7573), .Z(n7576) );
  XOR U7832 ( .A(n7575), .B(n7576), .Z(n7613) );
  NANDN U7833 ( .A(n7524), .B(n7523), .Z(n7528) );
  OR U7834 ( .A(n7526), .B(n7525), .Z(n7527) );
  AND U7835 ( .A(n7528), .B(n7527), .Z(n7612) );
  XNOR U7836 ( .A(n7613), .B(n7612), .Z(n7614) );
  NANDN U7837 ( .A(n7530), .B(n7529), .Z(n7534) );
  NANDN U7838 ( .A(n7532), .B(n7531), .Z(n7533) );
  NAND U7839 ( .A(n7534), .B(n7533), .Z(n7615) );
  XNOR U7840 ( .A(n7614), .B(n7615), .Z(n7560) );
  XOR U7841 ( .A(n7561), .B(n7560), .Z(n7619) );
  NANDN U7842 ( .A(n7536), .B(n7535), .Z(n7540) );
  NANDN U7843 ( .A(n7538), .B(n7537), .Z(n7539) );
  AND U7844 ( .A(n7540), .B(n7539), .Z(n7618) );
  XNOR U7845 ( .A(n7619), .B(n7618), .Z(n7620) );
  XOR U7846 ( .A(n7621), .B(n7620), .Z(n7553) );
  NANDN U7847 ( .A(n7542), .B(n7541), .Z(n7546) );
  NAND U7848 ( .A(n7544), .B(n7543), .Z(n7545) );
  AND U7849 ( .A(n7546), .B(n7545), .Z(n7552) );
  XNOR U7850 ( .A(n7553), .B(n7552), .Z(n7554) );
  XNOR U7851 ( .A(n7555), .B(n7554), .Z(n7624) );
  XNOR U7852 ( .A(sreg[345]), .B(n7624), .Z(n7626) );
  NANDN U7853 ( .A(sreg[344]), .B(n7547), .Z(n7551) );
  NAND U7854 ( .A(n7549), .B(n7548), .Z(n7550) );
  NAND U7855 ( .A(n7551), .B(n7550), .Z(n7625) );
  XNOR U7856 ( .A(n7626), .B(n7625), .Z(c[345]) );
  NANDN U7857 ( .A(n7553), .B(n7552), .Z(n7557) );
  NANDN U7858 ( .A(n7555), .B(n7554), .Z(n7556) );
  AND U7859 ( .A(n7557), .B(n7556), .Z(n7632) );
  NANDN U7860 ( .A(n7559), .B(n7558), .Z(n7563) );
  NAND U7861 ( .A(n7561), .B(n7560), .Z(n7562) );
  AND U7862 ( .A(n7563), .B(n7562), .Z(n7698) );
  NAND U7863 ( .A(n7564), .B(n19724), .Z(n7566) );
  XOR U7864 ( .A(b[11]), .B(a[96]), .Z(n7668) );
  NAND U7865 ( .A(n19692), .B(n7668), .Z(n7565) );
  AND U7866 ( .A(n7566), .B(n7565), .Z(n7679) );
  NAND U7867 ( .A(n19838), .B(n7567), .Z(n7569) );
  XOR U7868 ( .A(b[15]), .B(a[92]), .Z(n7671) );
  NAND U7869 ( .A(n19805), .B(n7671), .Z(n7568) );
  AND U7870 ( .A(n7569), .B(n7568), .Z(n7678) );
  NAND U7871 ( .A(n35), .B(n7570), .Z(n7572) );
  XOR U7872 ( .A(b[9]), .B(a[98]), .Z(n7674) );
  NAND U7873 ( .A(n19598), .B(n7674), .Z(n7571) );
  NAND U7874 ( .A(n7572), .B(n7571), .Z(n7677) );
  XOR U7875 ( .A(n7678), .B(n7677), .Z(n7680) );
  XOR U7876 ( .A(n7679), .B(n7680), .Z(n7690) );
  NANDN U7877 ( .A(n7574), .B(n7573), .Z(n7578) );
  OR U7878 ( .A(n7576), .B(n7575), .Z(n7577) );
  AND U7879 ( .A(n7578), .B(n7577), .Z(n7689) );
  XNOR U7880 ( .A(n7690), .B(n7689), .Z(n7691) );
  NANDN U7881 ( .A(n7580), .B(n7579), .Z(n7584) );
  NANDN U7882 ( .A(n7582), .B(n7581), .Z(n7583) );
  NAND U7883 ( .A(n7584), .B(n7583), .Z(n7692) );
  XNOR U7884 ( .A(n7691), .B(n7692), .Z(n7638) );
  NANDN U7885 ( .A(n7586), .B(n7585), .Z(n7590) );
  NANDN U7886 ( .A(n7588), .B(n7587), .Z(n7589) );
  AND U7887 ( .A(n7590), .B(n7589), .Z(n7664) );
  NAND U7888 ( .A(b[0]), .B(a[106]), .Z(n7591) );
  XNOR U7889 ( .A(b[1]), .B(n7591), .Z(n7593) );
  NANDN U7890 ( .A(b[0]), .B(a[105]), .Z(n7592) );
  NAND U7891 ( .A(n7593), .B(n7592), .Z(n7644) );
  NAND U7892 ( .A(n19808), .B(n7594), .Z(n7596) );
  XOR U7893 ( .A(b[13]), .B(a[94]), .Z(n7647) );
  NAND U7894 ( .A(n19768), .B(n7647), .Z(n7595) );
  AND U7895 ( .A(n7596), .B(n7595), .Z(n7642) );
  AND U7896 ( .A(b[15]), .B(a[90]), .Z(n7641) );
  XNOR U7897 ( .A(n7642), .B(n7641), .Z(n7643) );
  XNOR U7898 ( .A(n7644), .B(n7643), .Z(n7662) );
  NAND U7899 ( .A(n33), .B(n7597), .Z(n7599) );
  XOR U7900 ( .A(b[5]), .B(a[102]), .Z(n7653) );
  NAND U7901 ( .A(n19342), .B(n7653), .Z(n7598) );
  AND U7902 ( .A(n7599), .B(n7598), .Z(n7686) );
  NAND U7903 ( .A(n34), .B(n7600), .Z(n7602) );
  XOR U7904 ( .A(b[7]), .B(a[100]), .Z(n7656) );
  NAND U7905 ( .A(n19486), .B(n7656), .Z(n7601) );
  AND U7906 ( .A(n7602), .B(n7601), .Z(n7684) );
  NAND U7907 ( .A(n31), .B(n7603), .Z(n7605) );
  XOR U7908 ( .A(b[3]), .B(a[104]), .Z(n7659) );
  NAND U7909 ( .A(n32), .B(n7659), .Z(n7604) );
  NAND U7910 ( .A(n7605), .B(n7604), .Z(n7683) );
  XNOR U7911 ( .A(n7684), .B(n7683), .Z(n7685) );
  XOR U7912 ( .A(n7686), .B(n7685), .Z(n7663) );
  XOR U7913 ( .A(n7662), .B(n7663), .Z(n7665) );
  XOR U7914 ( .A(n7664), .B(n7665), .Z(n7636) );
  NANDN U7915 ( .A(n7607), .B(n7606), .Z(n7611) );
  OR U7916 ( .A(n7609), .B(n7608), .Z(n7610) );
  AND U7917 ( .A(n7611), .B(n7610), .Z(n7635) );
  XNOR U7918 ( .A(n7636), .B(n7635), .Z(n7637) );
  XOR U7919 ( .A(n7638), .B(n7637), .Z(n7696) );
  NANDN U7920 ( .A(n7613), .B(n7612), .Z(n7617) );
  NANDN U7921 ( .A(n7615), .B(n7614), .Z(n7616) );
  AND U7922 ( .A(n7617), .B(n7616), .Z(n7695) );
  XNOR U7923 ( .A(n7696), .B(n7695), .Z(n7697) );
  XOR U7924 ( .A(n7698), .B(n7697), .Z(n7630) );
  NANDN U7925 ( .A(n7619), .B(n7618), .Z(n7623) );
  NAND U7926 ( .A(n7621), .B(n7620), .Z(n7622) );
  AND U7927 ( .A(n7623), .B(n7622), .Z(n7629) );
  XNOR U7928 ( .A(n7630), .B(n7629), .Z(n7631) );
  XNOR U7929 ( .A(n7632), .B(n7631), .Z(n7701) );
  XNOR U7930 ( .A(sreg[346]), .B(n7701), .Z(n7703) );
  NANDN U7931 ( .A(sreg[345]), .B(n7624), .Z(n7628) );
  NAND U7932 ( .A(n7626), .B(n7625), .Z(n7627) );
  NAND U7933 ( .A(n7628), .B(n7627), .Z(n7702) );
  XNOR U7934 ( .A(n7703), .B(n7702), .Z(c[346]) );
  NANDN U7935 ( .A(n7630), .B(n7629), .Z(n7634) );
  NANDN U7936 ( .A(n7632), .B(n7631), .Z(n7633) );
  AND U7937 ( .A(n7634), .B(n7633), .Z(n7709) );
  NANDN U7938 ( .A(n7636), .B(n7635), .Z(n7640) );
  NAND U7939 ( .A(n7638), .B(n7637), .Z(n7639) );
  AND U7940 ( .A(n7640), .B(n7639), .Z(n7775) );
  NANDN U7941 ( .A(n7642), .B(n7641), .Z(n7646) );
  NANDN U7942 ( .A(n7644), .B(n7643), .Z(n7645) );
  AND U7943 ( .A(n7646), .B(n7645), .Z(n7741) );
  NAND U7944 ( .A(n19808), .B(n7647), .Z(n7649) );
  XOR U7945 ( .A(b[13]), .B(a[95]), .Z(n7727) );
  NAND U7946 ( .A(n19768), .B(n7727), .Z(n7648) );
  AND U7947 ( .A(n7649), .B(n7648), .Z(n7719) );
  AND U7948 ( .A(b[15]), .B(a[91]), .Z(n7718) );
  XNOR U7949 ( .A(n7719), .B(n7718), .Z(n7720) );
  NAND U7950 ( .A(b[0]), .B(a[107]), .Z(n7650) );
  XNOR U7951 ( .A(b[1]), .B(n7650), .Z(n7652) );
  NANDN U7952 ( .A(b[0]), .B(a[106]), .Z(n7651) );
  NAND U7953 ( .A(n7652), .B(n7651), .Z(n7721) );
  XNOR U7954 ( .A(n7720), .B(n7721), .Z(n7739) );
  NAND U7955 ( .A(n33), .B(n7653), .Z(n7655) );
  XOR U7956 ( .A(b[5]), .B(a[103]), .Z(n7730) );
  NAND U7957 ( .A(n19342), .B(n7730), .Z(n7654) );
  AND U7958 ( .A(n7655), .B(n7654), .Z(n7763) );
  NAND U7959 ( .A(n34), .B(n7656), .Z(n7658) );
  XOR U7960 ( .A(b[7]), .B(a[101]), .Z(n7733) );
  NAND U7961 ( .A(n19486), .B(n7733), .Z(n7657) );
  AND U7962 ( .A(n7658), .B(n7657), .Z(n7761) );
  NAND U7963 ( .A(n31), .B(n7659), .Z(n7661) );
  XOR U7964 ( .A(b[3]), .B(a[105]), .Z(n7736) );
  NAND U7965 ( .A(n32), .B(n7736), .Z(n7660) );
  NAND U7966 ( .A(n7661), .B(n7660), .Z(n7760) );
  XNOR U7967 ( .A(n7761), .B(n7760), .Z(n7762) );
  XOR U7968 ( .A(n7763), .B(n7762), .Z(n7740) );
  XOR U7969 ( .A(n7739), .B(n7740), .Z(n7742) );
  XOR U7970 ( .A(n7741), .B(n7742), .Z(n7713) );
  NANDN U7971 ( .A(n7663), .B(n7662), .Z(n7667) );
  OR U7972 ( .A(n7665), .B(n7664), .Z(n7666) );
  AND U7973 ( .A(n7667), .B(n7666), .Z(n7712) );
  XNOR U7974 ( .A(n7713), .B(n7712), .Z(n7715) );
  NAND U7975 ( .A(n7668), .B(n19724), .Z(n7670) );
  XOR U7976 ( .A(b[11]), .B(a[97]), .Z(n7745) );
  NAND U7977 ( .A(n19692), .B(n7745), .Z(n7669) );
  AND U7978 ( .A(n7670), .B(n7669), .Z(n7756) );
  NAND U7979 ( .A(n19838), .B(n7671), .Z(n7673) );
  XOR U7980 ( .A(b[15]), .B(a[93]), .Z(n7748) );
  NAND U7981 ( .A(n19805), .B(n7748), .Z(n7672) );
  AND U7982 ( .A(n7673), .B(n7672), .Z(n7755) );
  NAND U7983 ( .A(n35), .B(n7674), .Z(n7676) );
  XOR U7984 ( .A(b[9]), .B(a[99]), .Z(n7751) );
  NAND U7985 ( .A(n19598), .B(n7751), .Z(n7675) );
  NAND U7986 ( .A(n7676), .B(n7675), .Z(n7754) );
  XOR U7987 ( .A(n7755), .B(n7754), .Z(n7757) );
  XOR U7988 ( .A(n7756), .B(n7757), .Z(n7767) );
  NANDN U7989 ( .A(n7678), .B(n7677), .Z(n7682) );
  OR U7990 ( .A(n7680), .B(n7679), .Z(n7681) );
  AND U7991 ( .A(n7682), .B(n7681), .Z(n7766) );
  XNOR U7992 ( .A(n7767), .B(n7766), .Z(n7768) );
  NANDN U7993 ( .A(n7684), .B(n7683), .Z(n7688) );
  NANDN U7994 ( .A(n7686), .B(n7685), .Z(n7687) );
  NAND U7995 ( .A(n7688), .B(n7687), .Z(n7769) );
  XNOR U7996 ( .A(n7768), .B(n7769), .Z(n7714) );
  XOR U7997 ( .A(n7715), .B(n7714), .Z(n7773) );
  NANDN U7998 ( .A(n7690), .B(n7689), .Z(n7694) );
  NANDN U7999 ( .A(n7692), .B(n7691), .Z(n7693) );
  AND U8000 ( .A(n7694), .B(n7693), .Z(n7772) );
  XNOR U8001 ( .A(n7773), .B(n7772), .Z(n7774) );
  XOR U8002 ( .A(n7775), .B(n7774), .Z(n7707) );
  NANDN U8003 ( .A(n7696), .B(n7695), .Z(n7700) );
  NAND U8004 ( .A(n7698), .B(n7697), .Z(n7699) );
  AND U8005 ( .A(n7700), .B(n7699), .Z(n7706) );
  XNOR U8006 ( .A(n7707), .B(n7706), .Z(n7708) );
  XNOR U8007 ( .A(n7709), .B(n7708), .Z(n7778) );
  XNOR U8008 ( .A(sreg[347]), .B(n7778), .Z(n7780) );
  NANDN U8009 ( .A(sreg[346]), .B(n7701), .Z(n7705) );
  NAND U8010 ( .A(n7703), .B(n7702), .Z(n7704) );
  NAND U8011 ( .A(n7705), .B(n7704), .Z(n7779) );
  XNOR U8012 ( .A(n7780), .B(n7779), .Z(c[347]) );
  NANDN U8013 ( .A(n7707), .B(n7706), .Z(n7711) );
  NANDN U8014 ( .A(n7709), .B(n7708), .Z(n7710) );
  AND U8015 ( .A(n7711), .B(n7710), .Z(n7786) );
  NANDN U8016 ( .A(n7713), .B(n7712), .Z(n7717) );
  NAND U8017 ( .A(n7715), .B(n7714), .Z(n7716) );
  AND U8018 ( .A(n7717), .B(n7716), .Z(n7852) );
  NANDN U8019 ( .A(n7719), .B(n7718), .Z(n7723) );
  NANDN U8020 ( .A(n7721), .B(n7720), .Z(n7722) );
  AND U8021 ( .A(n7723), .B(n7722), .Z(n7818) );
  NAND U8022 ( .A(b[0]), .B(a[108]), .Z(n7724) );
  XNOR U8023 ( .A(b[1]), .B(n7724), .Z(n7726) );
  NANDN U8024 ( .A(b[0]), .B(a[107]), .Z(n7725) );
  NAND U8025 ( .A(n7726), .B(n7725), .Z(n7798) );
  NAND U8026 ( .A(n19808), .B(n7727), .Z(n7729) );
  XOR U8027 ( .A(b[13]), .B(a[96]), .Z(n7804) );
  NAND U8028 ( .A(n19768), .B(n7804), .Z(n7728) );
  AND U8029 ( .A(n7729), .B(n7728), .Z(n7796) );
  AND U8030 ( .A(b[15]), .B(a[92]), .Z(n7795) );
  XNOR U8031 ( .A(n7796), .B(n7795), .Z(n7797) );
  XNOR U8032 ( .A(n7798), .B(n7797), .Z(n7816) );
  NAND U8033 ( .A(n33), .B(n7730), .Z(n7732) );
  XOR U8034 ( .A(b[5]), .B(a[104]), .Z(n7807) );
  NAND U8035 ( .A(n19342), .B(n7807), .Z(n7731) );
  AND U8036 ( .A(n7732), .B(n7731), .Z(n7840) );
  NAND U8037 ( .A(n34), .B(n7733), .Z(n7735) );
  XOR U8038 ( .A(b[7]), .B(a[102]), .Z(n7810) );
  NAND U8039 ( .A(n19486), .B(n7810), .Z(n7734) );
  AND U8040 ( .A(n7735), .B(n7734), .Z(n7838) );
  NAND U8041 ( .A(n31), .B(n7736), .Z(n7738) );
  XOR U8042 ( .A(b[3]), .B(a[106]), .Z(n7813) );
  NAND U8043 ( .A(n32), .B(n7813), .Z(n7737) );
  NAND U8044 ( .A(n7738), .B(n7737), .Z(n7837) );
  XNOR U8045 ( .A(n7838), .B(n7837), .Z(n7839) );
  XOR U8046 ( .A(n7840), .B(n7839), .Z(n7817) );
  XOR U8047 ( .A(n7816), .B(n7817), .Z(n7819) );
  XOR U8048 ( .A(n7818), .B(n7819), .Z(n7790) );
  NANDN U8049 ( .A(n7740), .B(n7739), .Z(n7744) );
  OR U8050 ( .A(n7742), .B(n7741), .Z(n7743) );
  AND U8051 ( .A(n7744), .B(n7743), .Z(n7789) );
  XNOR U8052 ( .A(n7790), .B(n7789), .Z(n7792) );
  NAND U8053 ( .A(n7745), .B(n19724), .Z(n7747) );
  XOR U8054 ( .A(b[11]), .B(a[98]), .Z(n7822) );
  NAND U8055 ( .A(n19692), .B(n7822), .Z(n7746) );
  AND U8056 ( .A(n7747), .B(n7746), .Z(n7833) );
  NAND U8057 ( .A(n19838), .B(n7748), .Z(n7750) );
  XOR U8058 ( .A(b[15]), .B(a[94]), .Z(n7825) );
  NAND U8059 ( .A(n19805), .B(n7825), .Z(n7749) );
  AND U8060 ( .A(n7750), .B(n7749), .Z(n7832) );
  NAND U8061 ( .A(n35), .B(n7751), .Z(n7753) );
  XOR U8062 ( .A(b[9]), .B(a[100]), .Z(n7828) );
  NAND U8063 ( .A(n19598), .B(n7828), .Z(n7752) );
  NAND U8064 ( .A(n7753), .B(n7752), .Z(n7831) );
  XOR U8065 ( .A(n7832), .B(n7831), .Z(n7834) );
  XOR U8066 ( .A(n7833), .B(n7834), .Z(n7844) );
  NANDN U8067 ( .A(n7755), .B(n7754), .Z(n7759) );
  OR U8068 ( .A(n7757), .B(n7756), .Z(n7758) );
  AND U8069 ( .A(n7759), .B(n7758), .Z(n7843) );
  XNOR U8070 ( .A(n7844), .B(n7843), .Z(n7845) );
  NANDN U8071 ( .A(n7761), .B(n7760), .Z(n7765) );
  NANDN U8072 ( .A(n7763), .B(n7762), .Z(n7764) );
  NAND U8073 ( .A(n7765), .B(n7764), .Z(n7846) );
  XNOR U8074 ( .A(n7845), .B(n7846), .Z(n7791) );
  XOR U8075 ( .A(n7792), .B(n7791), .Z(n7850) );
  NANDN U8076 ( .A(n7767), .B(n7766), .Z(n7771) );
  NANDN U8077 ( .A(n7769), .B(n7768), .Z(n7770) );
  AND U8078 ( .A(n7771), .B(n7770), .Z(n7849) );
  XNOR U8079 ( .A(n7850), .B(n7849), .Z(n7851) );
  XOR U8080 ( .A(n7852), .B(n7851), .Z(n7784) );
  NANDN U8081 ( .A(n7773), .B(n7772), .Z(n7777) );
  NAND U8082 ( .A(n7775), .B(n7774), .Z(n7776) );
  AND U8083 ( .A(n7777), .B(n7776), .Z(n7783) );
  XNOR U8084 ( .A(n7784), .B(n7783), .Z(n7785) );
  XNOR U8085 ( .A(n7786), .B(n7785), .Z(n7855) );
  XNOR U8086 ( .A(sreg[348]), .B(n7855), .Z(n7857) );
  NANDN U8087 ( .A(sreg[347]), .B(n7778), .Z(n7782) );
  NAND U8088 ( .A(n7780), .B(n7779), .Z(n7781) );
  NAND U8089 ( .A(n7782), .B(n7781), .Z(n7856) );
  XNOR U8090 ( .A(n7857), .B(n7856), .Z(c[348]) );
  NANDN U8091 ( .A(n7784), .B(n7783), .Z(n7788) );
  NANDN U8092 ( .A(n7786), .B(n7785), .Z(n7787) );
  AND U8093 ( .A(n7788), .B(n7787), .Z(n7863) );
  NANDN U8094 ( .A(n7790), .B(n7789), .Z(n7794) );
  NAND U8095 ( .A(n7792), .B(n7791), .Z(n7793) );
  AND U8096 ( .A(n7794), .B(n7793), .Z(n7929) );
  NANDN U8097 ( .A(n7796), .B(n7795), .Z(n7800) );
  NANDN U8098 ( .A(n7798), .B(n7797), .Z(n7799) );
  AND U8099 ( .A(n7800), .B(n7799), .Z(n7895) );
  NAND U8100 ( .A(b[0]), .B(a[109]), .Z(n7801) );
  XNOR U8101 ( .A(b[1]), .B(n7801), .Z(n7803) );
  NANDN U8102 ( .A(b[0]), .B(a[108]), .Z(n7802) );
  NAND U8103 ( .A(n7803), .B(n7802), .Z(n7875) );
  NAND U8104 ( .A(n19808), .B(n7804), .Z(n7806) );
  XOR U8105 ( .A(b[13]), .B(a[97]), .Z(n7881) );
  NAND U8106 ( .A(n19768), .B(n7881), .Z(n7805) );
  AND U8107 ( .A(n7806), .B(n7805), .Z(n7873) );
  AND U8108 ( .A(b[15]), .B(a[93]), .Z(n7872) );
  XNOR U8109 ( .A(n7873), .B(n7872), .Z(n7874) );
  XNOR U8110 ( .A(n7875), .B(n7874), .Z(n7893) );
  NAND U8111 ( .A(n33), .B(n7807), .Z(n7809) );
  XOR U8112 ( .A(b[5]), .B(a[105]), .Z(n7884) );
  NAND U8113 ( .A(n19342), .B(n7884), .Z(n7808) );
  AND U8114 ( .A(n7809), .B(n7808), .Z(n7917) );
  NAND U8115 ( .A(n34), .B(n7810), .Z(n7812) );
  XOR U8116 ( .A(b[7]), .B(a[103]), .Z(n7887) );
  NAND U8117 ( .A(n19486), .B(n7887), .Z(n7811) );
  AND U8118 ( .A(n7812), .B(n7811), .Z(n7915) );
  NAND U8119 ( .A(n31), .B(n7813), .Z(n7815) );
  XOR U8120 ( .A(b[3]), .B(a[107]), .Z(n7890) );
  NAND U8121 ( .A(n32), .B(n7890), .Z(n7814) );
  NAND U8122 ( .A(n7815), .B(n7814), .Z(n7914) );
  XNOR U8123 ( .A(n7915), .B(n7914), .Z(n7916) );
  XOR U8124 ( .A(n7917), .B(n7916), .Z(n7894) );
  XOR U8125 ( .A(n7893), .B(n7894), .Z(n7896) );
  XOR U8126 ( .A(n7895), .B(n7896), .Z(n7867) );
  NANDN U8127 ( .A(n7817), .B(n7816), .Z(n7821) );
  OR U8128 ( .A(n7819), .B(n7818), .Z(n7820) );
  AND U8129 ( .A(n7821), .B(n7820), .Z(n7866) );
  XNOR U8130 ( .A(n7867), .B(n7866), .Z(n7869) );
  NAND U8131 ( .A(n7822), .B(n19724), .Z(n7824) );
  XOR U8132 ( .A(b[11]), .B(a[99]), .Z(n7899) );
  NAND U8133 ( .A(n19692), .B(n7899), .Z(n7823) );
  AND U8134 ( .A(n7824), .B(n7823), .Z(n7910) );
  NAND U8135 ( .A(n19838), .B(n7825), .Z(n7827) );
  XOR U8136 ( .A(b[15]), .B(a[95]), .Z(n7902) );
  NAND U8137 ( .A(n19805), .B(n7902), .Z(n7826) );
  AND U8138 ( .A(n7827), .B(n7826), .Z(n7909) );
  NAND U8139 ( .A(n35), .B(n7828), .Z(n7830) );
  XOR U8140 ( .A(b[9]), .B(a[101]), .Z(n7905) );
  NAND U8141 ( .A(n19598), .B(n7905), .Z(n7829) );
  NAND U8142 ( .A(n7830), .B(n7829), .Z(n7908) );
  XOR U8143 ( .A(n7909), .B(n7908), .Z(n7911) );
  XOR U8144 ( .A(n7910), .B(n7911), .Z(n7921) );
  NANDN U8145 ( .A(n7832), .B(n7831), .Z(n7836) );
  OR U8146 ( .A(n7834), .B(n7833), .Z(n7835) );
  AND U8147 ( .A(n7836), .B(n7835), .Z(n7920) );
  XNOR U8148 ( .A(n7921), .B(n7920), .Z(n7922) );
  NANDN U8149 ( .A(n7838), .B(n7837), .Z(n7842) );
  NANDN U8150 ( .A(n7840), .B(n7839), .Z(n7841) );
  NAND U8151 ( .A(n7842), .B(n7841), .Z(n7923) );
  XNOR U8152 ( .A(n7922), .B(n7923), .Z(n7868) );
  XOR U8153 ( .A(n7869), .B(n7868), .Z(n7927) );
  NANDN U8154 ( .A(n7844), .B(n7843), .Z(n7848) );
  NANDN U8155 ( .A(n7846), .B(n7845), .Z(n7847) );
  AND U8156 ( .A(n7848), .B(n7847), .Z(n7926) );
  XNOR U8157 ( .A(n7927), .B(n7926), .Z(n7928) );
  XOR U8158 ( .A(n7929), .B(n7928), .Z(n7861) );
  NANDN U8159 ( .A(n7850), .B(n7849), .Z(n7854) );
  NAND U8160 ( .A(n7852), .B(n7851), .Z(n7853) );
  AND U8161 ( .A(n7854), .B(n7853), .Z(n7860) );
  XNOR U8162 ( .A(n7861), .B(n7860), .Z(n7862) );
  XNOR U8163 ( .A(n7863), .B(n7862), .Z(n7932) );
  XNOR U8164 ( .A(sreg[349]), .B(n7932), .Z(n7934) );
  NANDN U8165 ( .A(sreg[348]), .B(n7855), .Z(n7859) );
  NAND U8166 ( .A(n7857), .B(n7856), .Z(n7858) );
  NAND U8167 ( .A(n7859), .B(n7858), .Z(n7933) );
  XNOR U8168 ( .A(n7934), .B(n7933), .Z(c[349]) );
  NANDN U8169 ( .A(n7861), .B(n7860), .Z(n7865) );
  NANDN U8170 ( .A(n7863), .B(n7862), .Z(n7864) );
  AND U8171 ( .A(n7865), .B(n7864), .Z(n7940) );
  NANDN U8172 ( .A(n7867), .B(n7866), .Z(n7871) );
  NAND U8173 ( .A(n7869), .B(n7868), .Z(n7870) );
  AND U8174 ( .A(n7871), .B(n7870), .Z(n8006) );
  NANDN U8175 ( .A(n7873), .B(n7872), .Z(n7877) );
  NANDN U8176 ( .A(n7875), .B(n7874), .Z(n7876) );
  AND U8177 ( .A(n7877), .B(n7876), .Z(n7972) );
  NAND U8178 ( .A(b[0]), .B(a[110]), .Z(n7878) );
  XNOR U8179 ( .A(b[1]), .B(n7878), .Z(n7880) );
  NANDN U8180 ( .A(b[0]), .B(a[109]), .Z(n7879) );
  NAND U8181 ( .A(n7880), .B(n7879), .Z(n7952) );
  NAND U8182 ( .A(n19808), .B(n7881), .Z(n7883) );
  XOR U8183 ( .A(b[13]), .B(a[98]), .Z(n7955) );
  NAND U8184 ( .A(n19768), .B(n7955), .Z(n7882) );
  AND U8185 ( .A(n7883), .B(n7882), .Z(n7950) );
  AND U8186 ( .A(b[15]), .B(a[94]), .Z(n7949) );
  XNOR U8187 ( .A(n7950), .B(n7949), .Z(n7951) );
  XNOR U8188 ( .A(n7952), .B(n7951), .Z(n7970) );
  NAND U8189 ( .A(n33), .B(n7884), .Z(n7886) );
  XOR U8190 ( .A(b[5]), .B(a[106]), .Z(n7961) );
  NAND U8191 ( .A(n19342), .B(n7961), .Z(n7885) );
  AND U8192 ( .A(n7886), .B(n7885), .Z(n7994) );
  NAND U8193 ( .A(n34), .B(n7887), .Z(n7889) );
  XOR U8194 ( .A(b[7]), .B(a[104]), .Z(n7964) );
  NAND U8195 ( .A(n19486), .B(n7964), .Z(n7888) );
  AND U8196 ( .A(n7889), .B(n7888), .Z(n7992) );
  NAND U8197 ( .A(n31), .B(n7890), .Z(n7892) );
  XOR U8198 ( .A(b[3]), .B(a[108]), .Z(n7967) );
  NAND U8199 ( .A(n32), .B(n7967), .Z(n7891) );
  NAND U8200 ( .A(n7892), .B(n7891), .Z(n7991) );
  XNOR U8201 ( .A(n7992), .B(n7991), .Z(n7993) );
  XOR U8202 ( .A(n7994), .B(n7993), .Z(n7971) );
  XOR U8203 ( .A(n7970), .B(n7971), .Z(n7973) );
  XOR U8204 ( .A(n7972), .B(n7973), .Z(n7944) );
  NANDN U8205 ( .A(n7894), .B(n7893), .Z(n7898) );
  OR U8206 ( .A(n7896), .B(n7895), .Z(n7897) );
  AND U8207 ( .A(n7898), .B(n7897), .Z(n7943) );
  XNOR U8208 ( .A(n7944), .B(n7943), .Z(n7946) );
  NAND U8209 ( .A(n7899), .B(n19724), .Z(n7901) );
  XOR U8210 ( .A(b[11]), .B(a[100]), .Z(n7976) );
  NAND U8211 ( .A(n19692), .B(n7976), .Z(n7900) );
  AND U8212 ( .A(n7901), .B(n7900), .Z(n7987) );
  NAND U8213 ( .A(n19838), .B(n7902), .Z(n7904) );
  XOR U8214 ( .A(b[15]), .B(a[96]), .Z(n7979) );
  NAND U8215 ( .A(n19805), .B(n7979), .Z(n7903) );
  AND U8216 ( .A(n7904), .B(n7903), .Z(n7986) );
  NAND U8217 ( .A(n35), .B(n7905), .Z(n7907) );
  XOR U8218 ( .A(b[9]), .B(a[102]), .Z(n7982) );
  NAND U8219 ( .A(n19598), .B(n7982), .Z(n7906) );
  NAND U8220 ( .A(n7907), .B(n7906), .Z(n7985) );
  XOR U8221 ( .A(n7986), .B(n7985), .Z(n7988) );
  XOR U8222 ( .A(n7987), .B(n7988), .Z(n7998) );
  NANDN U8223 ( .A(n7909), .B(n7908), .Z(n7913) );
  OR U8224 ( .A(n7911), .B(n7910), .Z(n7912) );
  AND U8225 ( .A(n7913), .B(n7912), .Z(n7997) );
  XNOR U8226 ( .A(n7998), .B(n7997), .Z(n7999) );
  NANDN U8227 ( .A(n7915), .B(n7914), .Z(n7919) );
  NANDN U8228 ( .A(n7917), .B(n7916), .Z(n7918) );
  NAND U8229 ( .A(n7919), .B(n7918), .Z(n8000) );
  XNOR U8230 ( .A(n7999), .B(n8000), .Z(n7945) );
  XOR U8231 ( .A(n7946), .B(n7945), .Z(n8004) );
  NANDN U8232 ( .A(n7921), .B(n7920), .Z(n7925) );
  NANDN U8233 ( .A(n7923), .B(n7922), .Z(n7924) );
  AND U8234 ( .A(n7925), .B(n7924), .Z(n8003) );
  XNOR U8235 ( .A(n8004), .B(n8003), .Z(n8005) );
  XOR U8236 ( .A(n8006), .B(n8005), .Z(n7938) );
  NANDN U8237 ( .A(n7927), .B(n7926), .Z(n7931) );
  NAND U8238 ( .A(n7929), .B(n7928), .Z(n7930) );
  AND U8239 ( .A(n7931), .B(n7930), .Z(n7937) );
  XNOR U8240 ( .A(n7938), .B(n7937), .Z(n7939) );
  XNOR U8241 ( .A(n7940), .B(n7939), .Z(n8009) );
  XNOR U8242 ( .A(sreg[350]), .B(n8009), .Z(n8011) );
  NANDN U8243 ( .A(sreg[349]), .B(n7932), .Z(n7936) );
  NAND U8244 ( .A(n7934), .B(n7933), .Z(n7935) );
  NAND U8245 ( .A(n7936), .B(n7935), .Z(n8010) );
  XNOR U8246 ( .A(n8011), .B(n8010), .Z(c[350]) );
  NANDN U8247 ( .A(n7938), .B(n7937), .Z(n7942) );
  NANDN U8248 ( .A(n7940), .B(n7939), .Z(n7941) );
  AND U8249 ( .A(n7942), .B(n7941), .Z(n8017) );
  NANDN U8250 ( .A(n7944), .B(n7943), .Z(n7948) );
  NAND U8251 ( .A(n7946), .B(n7945), .Z(n7947) );
  AND U8252 ( .A(n7948), .B(n7947), .Z(n8083) );
  NANDN U8253 ( .A(n7950), .B(n7949), .Z(n7954) );
  NANDN U8254 ( .A(n7952), .B(n7951), .Z(n7953) );
  AND U8255 ( .A(n7954), .B(n7953), .Z(n8049) );
  NAND U8256 ( .A(n19808), .B(n7955), .Z(n7957) );
  XOR U8257 ( .A(b[13]), .B(a[99]), .Z(n8035) );
  NAND U8258 ( .A(n19768), .B(n8035), .Z(n7956) );
  AND U8259 ( .A(n7957), .B(n7956), .Z(n8027) );
  AND U8260 ( .A(b[15]), .B(a[95]), .Z(n8026) );
  XNOR U8261 ( .A(n8027), .B(n8026), .Z(n8028) );
  NAND U8262 ( .A(b[0]), .B(a[111]), .Z(n7958) );
  XNOR U8263 ( .A(b[1]), .B(n7958), .Z(n7960) );
  NANDN U8264 ( .A(b[0]), .B(a[110]), .Z(n7959) );
  NAND U8265 ( .A(n7960), .B(n7959), .Z(n8029) );
  XNOR U8266 ( .A(n8028), .B(n8029), .Z(n8047) );
  NAND U8267 ( .A(n33), .B(n7961), .Z(n7963) );
  XOR U8268 ( .A(b[5]), .B(a[107]), .Z(n8038) );
  NAND U8269 ( .A(n19342), .B(n8038), .Z(n7962) );
  AND U8270 ( .A(n7963), .B(n7962), .Z(n8071) );
  NAND U8271 ( .A(n34), .B(n7964), .Z(n7966) );
  XOR U8272 ( .A(b[7]), .B(a[105]), .Z(n8041) );
  NAND U8273 ( .A(n19486), .B(n8041), .Z(n7965) );
  AND U8274 ( .A(n7966), .B(n7965), .Z(n8069) );
  NAND U8275 ( .A(n31), .B(n7967), .Z(n7969) );
  XOR U8276 ( .A(b[3]), .B(a[109]), .Z(n8044) );
  NAND U8277 ( .A(n32), .B(n8044), .Z(n7968) );
  NAND U8278 ( .A(n7969), .B(n7968), .Z(n8068) );
  XNOR U8279 ( .A(n8069), .B(n8068), .Z(n8070) );
  XOR U8280 ( .A(n8071), .B(n8070), .Z(n8048) );
  XOR U8281 ( .A(n8047), .B(n8048), .Z(n8050) );
  XOR U8282 ( .A(n8049), .B(n8050), .Z(n8021) );
  NANDN U8283 ( .A(n7971), .B(n7970), .Z(n7975) );
  OR U8284 ( .A(n7973), .B(n7972), .Z(n7974) );
  AND U8285 ( .A(n7975), .B(n7974), .Z(n8020) );
  XNOR U8286 ( .A(n8021), .B(n8020), .Z(n8023) );
  NAND U8287 ( .A(n7976), .B(n19724), .Z(n7978) );
  XOR U8288 ( .A(b[11]), .B(a[101]), .Z(n8053) );
  NAND U8289 ( .A(n19692), .B(n8053), .Z(n7977) );
  AND U8290 ( .A(n7978), .B(n7977), .Z(n8064) );
  NAND U8291 ( .A(n19838), .B(n7979), .Z(n7981) );
  XOR U8292 ( .A(b[15]), .B(a[97]), .Z(n8056) );
  NAND U8293 ( .A(n19805), .B(n8056), .Z(n7980) );
  AND U8294 ( .A(n7981), .B(n7980), .Z(n8063) );
  NAND U8295 ( .A(n35), .B(n7982), .Z(n7984) );
  XOR U8296 ( .A(b[9]), .B(a[103]), .Z(n8059) );
  NAND U8297 ( .A(n19598), .B(n8059), .Z(n7983) );
  NAND U8298 ( .A(n7984), .B(n7983), .Z(n8062) );
  XOR U8299 ( .A(n8063), .B(n8062), .Z(n8065) );
  XOR U8300 ( .A(n8064), .B(n8065), .Z(n8075) );
  NANDN U8301 ( .A(n7986), .B(n7985), .Z(n7990) );
  OR U8302 ( .A(n7988), .B(n7987), .Z(n7989) );
  AND U8303 ( .A(n7990), .B(n7989), .Z(n8074) );
  XNOR U8304 ( .A(n8075), .B(n8074), .Z(n8076) );
  NANDN U8305 ( .A(n7992), .B(n7991), .Z(n7996) );
  NANDN U8306 ( .A(n7994), .B(n7993), .Z(n7995) );
  NAND U8307 ( .A(n7996), .B(n7995), .Z(n8077) );
  XNOR U8308 ( .A(n8076), .B(n8077), .Z(n8022) );
  XOR U8309 ( .A(n8023), .B(n8022), .Z(n8081) );
  NANDN U8310 ( .A(n7998), .B(n7997), .Z(n8002) );
  NANDN U8311 ( .A(n8000), .B(n7999), .Z(n8001) );
  AND U8312 ( .A(n8002), .B(n8001), .Z(n8080) );
  XNOR U8313 ( .A(n8081), .B(n8080), .Z(n8082) );
  XOR U8314 ( .A(n8083), .B(n8082), .Z(n8015) );
  NANDN U8315 ( .A(n8004), .B(n8003), .Z(n8008) );
  NAND U8316 ( .A(n8006), .B(n8005), .Z(n8007) );
  AND U8317 ( .A(n8008), .B(n8007), .Z(n8014) );
  XNOR U8318 ( .A(n8015), .B(n8014), .Z(n8016) );
  XNOR U8319 ( .A(n8017), .B(n8016), .Z(n8086) );
  XNOR U8320 ( .A(sreg[351]), .B(n8086), .Z(n8088) );
  NANDN U8321 ( .A(sreg[350]), .B(n8009), .Z(n8013) );
  NAND U8322 ( .A(n8011), .B(n8010), .Z(n8012) );
  NAND U8323 ( .A(n8013), .B(n8012), .Z(n8087) );
  XNOR U8324 ( .A(n8088), .B(n8087), .Z(c[351]) );
  NANDN U8325 ( .A(n8015), .B(n8014), .Z(n8019) );
  NANDN U8326 ( .A(n8017), .B(n8016), .Z(n8018) );
  AND U8327 ( .A(n8019), .B(n8018), .Z(n8094) );
  NANDN U8328 ( .A(n8021), .B(n8020), .Z(n8025) );
  NAND U8329 ( .A(n8023), .B(n8022), .Z(n8024) );
  AND U8330 ( .A(n8025), .B(n8024), .Z(n8160) );
  NANDN U8331 ( .A(n8027), .B(n8026), .Z(n8031) );
  NANDN U8332 ( .A(n8029), .B(n8028), .Z(n8030) );
  AND U8333 ( .A(n8031), .B(n8030), .Z(n8126) );
  NAND U8334 ( .A(b[0]), .B(a[112]), .Z(n8032) );
  XNOR U8335 ( .A(b[1]), .B(n8032), .Z(n8034) );
  NANDN U8336 ( .A(b[0]), .B(a[111]), .Z(n8033) );
  NAND U8337 ( .A(n8034), .B(n8033), .Z(n8106) );
  NAND U8338 ( .A(n19808), .B(n8035), .Z(n8037) );
  XOR U8339 ( .A(b[13]), .B(a[100]), .Z(n8112) );
  NAND U8340 ( .A(n19768), .B(n8112), .Z(n8036) );
  AND U8341 ( .A(n8037), .B(n8036), .Z(n8104) );
  AND U8342 ( .A(b[15]), .B(a[96]), .Z(n8103) );
  XNOR U8343 ( .A(n8104), .B(n8103), .Z(n8105) );
  XNOR U8344 ( .A(n8106), .B(n8105), .Z(n8124) );
  NAND U8345 ( .A(n33), .B(n8038), .Z(n8040) );
  XOR U8346 ( .A(b[5]), .B(a[108]), .Z(n8115) );
  NAND U8347 ( .A(n19342), .B(n8115), .Z(n8039) );
  AND U8348 ( .A(n8040), .B(n8039), .Z(n8148) );
  NAND U8349 ( .A(n34), .B(n8041), .Z(n8043) );
  XOR U8350 ( .A(b[7]), .B(a[106]), .Z(n8118) );
  NAND U8351 ( .A(n19486), .B(n8118), .Z(n8042) );
  AND U8352 ( .A(n8043), .B(n8042), .Z(n8146) );
  NAND U8353 ( .A(n31), .B(n8044), .Z(n8046) );
  XOR U8354 ( .A(b[3]), .B(a[110]), .Z(n8121) );
  NAND U8355 ( .A(n32), .B(n8121), .Z(n8045) );
  NAND U8356 ( .A(n8046), .B(n8045), .Z(n8145) );
  XNOR U8357 ( .A(n8146), .B(n8145), .Z(n8147) );
  XOR U8358 ( .A(n8148), .B(n8147), .Z(n8125) );
  XOR U8359 ( .A(n8124), .B(n8125), .Z(n8127) );
  XOR U8360 ( .A(n8126), .B(n8127), .Z(n8098) );
  NANDN U8361 ( .A(n8048), .B(n8047), .Z(n8052) );
  OR U8362 ( .A(n8050), .B(n8049), .Z(n8051) );
  AND U8363 ( .A(n8052), .B(n8051), .Z(n8097) );
  XNOR U8364 ( .A(n8098), .B(n8097), .Z(n8100) );
  NAND U8365 ( .A(n8053), .B(n19724), .Z(n8055) );
  XOR U8366 ( .A(b[11]), .B(a[102]), .Z(n8130) );
  NAND U8367 ( .A(n19692), .B(n8130), .Z(n8054) );
  AND U8368 ( .A(n8055), .B(n8054), .Z(n8141) );
  NAND U8369 ( .A(n19838), .B(n8056), .Z(n8058) );
  XOR U8370 ( .A(b[15]), .B(a[98]), .Z(n8133) );
  NAND U8371 ( .A(n19805), .B(n8133), .Z(n8057) );
  AND U8372 ( .A(n8058), .B(n8057), .Z(n8140) );
  NAND U8373 ( .A(n35), .B(n8059), .Z(n8061) );
  XOR U8374 ( .A(b[9]), .B(a[104]), .Z(n8136) );
  NAND U8375 ( .A(n19598), .B(n8136), .Z(n8060) );
  NAND U8376 ( .A(n8061), .B(n8060), .Z(n8139) );
  XOR U8377 ( .A(n8140), .B(n8139), .Z(n8142) );
  XOR U8378 ( .A(n8141), .B(n8142), .Z(n8152) );
  NANDN U8379 ( .A(n8063), .B(n8062), .Z(n8067) );
  OR U8380 ( .A(n8065), .B(n8064), .Z(n8066) );
  AND U8381 ( .A(n8067), .B(n8066), .Z(n8151) );
  XNOR U8382 ( .A(n8152), .B(n8151), .Z(n8153) );
  NANDN U8383 ( .A(n8069), .B(n8068), .Z(n8073) );
  NANDN U8384 ( .A(n8071), .B(n8070), .Z(n8072) );
  NAND U8385 ( .A(n8073), .B(n8072), .Z(n8154) );
  XNOR U8386 ( .A(n8153), .B(n8154), .Z(n8099) );
  XOR U8387 ( .A(n8100), .B(n8099), .Z(n8158) );
  NANDN U8388 ( .A(n8075), .B(n8074), .Z(n8079) );
  NANDN U8389 ( .A(n8077), .B(n8076), .Z(n8078) );
  AND U8390 ( .A(n8079), .B(n8078), .Z(n8157) );
  XNOR U8391 ( .A(n8158), .B(n8157), .Z(n8159) );
  XOR U8392 ( .A(n8160), .B(n8159), .Z(n8092) );
  NANDN U8393 ( .A(n8081), .B(n8080), .Z(n8085) );
  NAND U8394 ( .A(n8083), .B(n8082), .Z(n8084) );
  AND U8395 ( .A(n8085), .B(n8084), .Z(n8091) );
  XNOR U8396 ( .A(n8092), .B(n8091), .Z(n8093) );
  XNOR U8397 ( .A(n8094), .B(n8093), .Z(n8163) );
  XNOR U8398 ( .A(sreg[352]), .B(n8163), .Z(n8165) );
  NANDN U8399 ( .A(sreg[351]), .B(n8086), .Z(n8090) );
  NAND U8400 ( .A(n8088), .B(n8087), .Z(n8089) );
  NAND U8401 ( .A(n8090), .B(n8089), .Z(n8164) );
  XNOR U8402 ( .A(n8165), .B(n8164), .Z(c[352]) );
  NANDN U8403 ( .A(n8092), .B(n8091), .Z(n8096) );
  NANDN U8404 ( .A(n8094), .B(n8093), .Z(n8095) );
  AND U8405 ( .A(n8096), .B(n8095), .Z(n8171) );
  NANDN U8406 ( .A(n8098), .B(n8097), .Z(n8102) );
  NAND U8407 ( .A(n8100), .B(n8099), .Z(n8101) );
  AND U8408 ( .A(n8102), .B(n8101), .Z(n8237) );
  NANDN U8409 ( .A(n8104), .B(n8103), .Z(n8108) );
  NANDN U8410 ( .A(n8106), .B(n8105), .Z(n8107) );
  AND U8411 ( .A(n8108), .B(n8107), .Z(n8203) );
  NAND U8412 ( .A(b[0]), .B(a[113]), .Z(n8109) );
  XNOR U8413 ( .A(b[1]), .B(n8109), .Z(n8111) );
  NANDN U8414 ( .A(b[0]), .B(a[112]), .Z(n8110) );
  NAND U8415 ( .A(n8111), .B(n8110), .Z(n8183) );
  NAND U8416 ( .A(n19808), .B(n8112), .Z(n8114) );
  XOR U8417 ( .A(b[13]), .B(a[101]), .Z(n8189) );
  NAND U8418 ( .A(n19768), .B(n8189), .Z(n8113) );
  AND U8419 ( .A(n8114), .B(n8113), .Z(n8181) );
  AND U8420 ( .A(b[15]), .B(a[97]), .Z(n8180) );
  XNOR U8421 ( .A(n8181), .B(n8180), .Z(n8182) );
  XNOR U8422 ( .A(n8183), .B(n8182), .Z(n8201) );
  NAND U8423 ( .A(n33), .B(n8115), .Z(n8117) );
  XOR U8424 ( .A(b[5]), .B(a[109]), .Z(n8192) );
  NAND U8425 ( .A(n19342), .B(n8192), .Z(n8116) );
  AND U8426 ( .A(n8117), .B(n8116), .Z(n8225) );
  NAND U8427 ( .A(n34), .B(n8118), .Z(n8120) );
  XOR U8428 ( .A(b[7]), .B(a[107]), .Z(n8195) );
  NAND U8429 ( .A(n19486), .B(n8195), .Z(n8119) );
  AND U8430 ( .A(n8120), .B(n8119), .Z(n8223) );
  NAND U8431 ( .A(n31), .B(n8121), .Z(n8123) );
  XOR U8432 ( .A(b[3]), .B(a[111]), .Z(n8198) );
  NAND U8433 ( .A(n32), .B(n8198), .Z(n8122) );
  NAND U8434 ( .A(n8123), .B(n8122), .Z(n8222) );
  XNOR U8435 ( .A(n8223), .B(n8222), .Z(n8224) );
  XOR U8436 ( .A(n8225), .B(n8224), .Z(n8202) );
  XOR U8437 ( .A(n8201), .B(n8202), .Z(n8204) );
  XOR U8438 ( .A(n8203), .B(n8204), .Z(n8175) );
  NANDN U8439 ( .A(n8125), .B(n8124), .Z(n8129) );
  OR U8440 ( .A(n8127), .B(n8126), .Z(n8128) );
  AND U8441 ( .A(n8129), .B(n8128), .Z(n8174) );
  XNOR U8442 ( .A(n8175), .B(n8174), .Z(n8177) );
  NAND U8443 ( .A(n8130), .B(n19724), .Z(n8132) );
  XOR U8444 ( .A(b[11]), .B(a[103]), .Z(n8207) );
  NAND U8445 ( .A(n19692), .B(n8207), .Z(n8131) );
  AND U8446 ( .A(n8132), .B(n8131), .Z(n8218) );
  NAND U8447 ( .A(n19838), .B(n8133), .Z(n8135) );
  XOR U8448 ( .A(b[15]), .B(a[99]), .Z(n8210) );
  NAND U8449 ( .A(n19805), .B(n8210), .Z(n8134) );
  AND U8450 ( .A(n8135), .B(n8134), .Z(n8217) );
  NAND U8451 ( .A(n35), .B(n8136), .Z(n8138) );
  XOR U8452 ( .A(b[9]), .B(a[105]), .Z(n8213) );
  NAND U8453 ( .A(n19598), .B(n8213), .Z(n8137) );
  NAND U8454 ( .A(n8138), .B(n8137), .Z(n8216) );
  XOR U8455 ( .A(n8217), .B(n8216), .Z(n8219) );
  XOR U8456 ( .A(n8218), .B(n8219), .Z(n8229) );
  NANDN U8457 ( .A(n8140), .B(n8139), .Z(n8144) );
  OR U8458 ( .A(n8142), .B(n8141), .Z(n8143) );
  AND U8459 ( .A(n8144), .B(n8143), .Z(n8228) );
  XNOR U8460 ( .A(n8229), .B(n8228), .Z(n8230) );
  NANDN U8461 ( .A(n8146), .B(n8145), .Z(n8150) );
  NANDN U8462 ( .A(n8148), .B(n8147), .Z(n8149) );
  NAND U8463 ( .A(n8150), .B(n8149), .Z(n8231) );
  XNOR U8464 ( .A(n8230), .B(n8231), .Z(n8176) );
  XOR U8465 ( .A(n8177), .B(n8176), .Z(n8235) );
  NANDN U8466 ( .A(n8152), .B(n8151), .Z(n8156) );
  NANDN U8467 ( .A(n8154), .B(n8153), .Z(n8155) );
  AND U8468 ( .A(n8156), .B(n8155), .Z(n8234) );
  XNOR U8469 ( .A(n8235), .B(n8234), .Z(n8236) );
  XOR U8470 ( .A(n8237), .B(n8236), .Z(n8169) );
  NANDN U8471 ( .A(n8158), .B(n8157), .Z(n8162) );
  NAND U8472 ( .A(n8160), .B(n8159), .Z(n8161) );
  AND U8473 ( .A(n8162), .B(n8161), .Z(n8168) );
  XNOR U8474 ( .A(n8169), .B(n8168), .Z(n8170) );
  XNOR U8475 ( .A(n8171), .B(n8170), .Z(n8240) );
  XNOR U8476 ( .A(sreg[353]), .B(n8240), .Z(n8242) );
  NANDN U8477 ( .A(sreg[352]), .B(n8163), .Z(n8167) );
  NAND U8478 ( .A(n8165), .B(n8164), .Z(n8166) );
  NAND U8479 ( .A(n8167), .B(n8166), .Z(n8241) );
  XNOR U8480 ( .A(n8242), .B(n8241), .Z(c[353]) );
  NANDN U8481 ( .A(n8169), .B(n8168), .Z(n8173) );
  NANDN U8482 ( .A(n8171), .B(n8170), .Z(n8172) );
  AND U8483 ( .A(n8173), .B(n8172), .Z(n8248) );
  NANDN U8484 ( .A(n8175), .B(n8174), .Z(n8179) );
  NAND U8485 ( .A(n8177), .B(n8176), .Z(n8178) );
  AND U8486 ( .A(n8179), .B(n8178), .Z(n8314) );
  NANDN U8487 ( .A(n8181), .B(n8180), .Z(n8185) );
  NANDN U8488 ( .A(n8183), .B(n8182), .Z(n8184) );
  AND U8489 ( .A(n8185), .B(n8184), .Z(n8280) );
  NAND U8490 ( .A(b[0]), .B(a[114]), .Z(n8186) );
  XNOR U8491 ( .A(b[1]), .B(n8186), .Z(n8188) );
  NANDN U8492 ( .A(b[0]), .B(a[113]), .Z(n8187) );
  NAND U8493 ( .A(n8188), .B(n8187), .Z(n8260) );
  NAND U8494 ( .A(n19808), .B(n8189), .Z(n8191) );
  XOR U8495 ( .A(b[13]), .B(a[102]), .Z(n8266) );
  NAND U8496 ( .A(n19768), .B(n8266), .Z(n8190) );
  AND U8497 ( .A(n8191), .B(n8190), .Z(n8258) );
  AND U8498 ( .A(b[15]), .B(a[98]), .Z(n8257) );
  XNOR U8499 ( .A(n8258), .B(n8257), .Z(n8259) );
  XNOR U8500 ( .A(n8260), .B(n8259), .Z(n8278) );
  NAND U8501 ( .A(n33), .B(n8192), .Z(n8194) );
  XOR U8502 ( .A(b[5]), .B(a[110]), .Z(n8269) );
  NAND U8503 ( .A(n19342), .B(n8269), .Z(n8193) );
  AND U8504 ( .A(n8194), .B(n8193), .Z(n8302) );
  NAND U8505 ( .A(n34), .B(n8195), .Z(n8197) );
  XOR U8506 ( .A(b[7]), .B(a[108]), .Z(n8272) );
  NAND U8507 ( .A(n19486), .B(n8272), .Z(n8196) );
  AND U8508 ( .A(n8197), .B(n8196), .Z(n8300) );
  NAND U8509 ( .A(n31), .B(n8198), .Z(n8200) );
  XOR U8510 ( .A(b[3]), .B(a[112]), .Z(n8275) );
  NAND U8511 ( .A(n32), .B(n8275), .Z(n8199) );
  NAND U8512 ( .A(n8200), .B(n8199), .Z(n8299) );
  XNOR U8513 ( .A(n8300), .B(n8299), .Z(n8301) );
  XOR U8514 ( .A(n8302), .B(n8301), .Z(n8279) );
  XOR U8515 ( .A(n8278), .B(n8279), .Z(n8281) );
  XOR U8516 ( .A(n8280), .B(n8281), .Z(n8252) );
  NANDN U8517 ( .A(n8202), .B(n8201), .Z(n8206) );
  OR U8518 ( .A(n8204), .B(n8203), .Z(n8205) );
  AND U8519 ( .A(n8206), .B(n8205), .Z(n8251) );
  XNOR U8520 ( .A(n8252), .B(n8251), .Z(n8254) );
  NAND U8521 ( .A(n8207), .B(n19724), .Z(n8209) );
  XOR U8522 ( .A(b[11]), .B(a[104]), .Z(n8284) );
  NAND U8523 ( .A(n19692), .B(n8284), .Z(n8208) );
  AND U8524 ( .A(n8209), .B(n8208), .Z(n8295) );
  NAND U8525 ( .A(n19838), .B(n8210), .Z(n8212) );
  XOR U8526 ( .A(b[15]), .B(a[100]), .Z(n8287) );
  NAND U8527 ( .A(n19805), .B(n8287), .Z(n8211) );
  AND U8528 ( .A(n8212), .B(n8211), .Z(n8294) );
  NAND U8529 ( .A(n35), .B(n8213), .Z(n8215) );
  XOR U8530 ( .A(b[9]), .B(a[106]), .Z(n8290) );
  NAND U8531 ( .A(n19598), .B(n8290), .Z(n8214) );
  NAND U8532 ( .A(n8215), .B(n8214), .Z(n8293) );
  XOR U8533 ( .A(n8294), .B(n8293), .Z(n8296) );
  XOR U8534 ( .A(n8295), .B(n8296), .Z(n8306) );
  NANDN U8535 ( .A(n8217), .B(n8216), .Z(n8221) );
  OR U8536 ( .A(n8219), .B(n8218), .Z(n8220) );
  AND U8537 ( .A(n8221), .B(n8220), .Z(n8305) );
  XNOR U8538 ( .A(n8306), .B(n8305), .Z(n8307) );
  NANDN U8539 ( .A(n8223), .B(n8222), .Z(n8227) );
  NANDN U8540 ( .A(n8225), .B(n8224), .Z(n8226) );
  NAND U8541 ( .A(n8227), .B(n8226), .Z(n8308) );
  XNOR U8542 ( .A(n8307), .B(n8308), .Z(n8253) );
  XOR U8543 ( .A(n8254), .B(n8253), .Z(n8312) );
  NANDN U8544 ( .A(n8229), .B(n8228), .Z(n8233) );
  NANDN U8545 ( .A(n8231), .B(n8230), .Z(n8232) );
  AND U8546 ( .A(n8233), .B(n8232), .Z(n8311) );
  XNOR U8547 ( .A(n8312), .B(n8311), .Z(n8313) );
  XOR U8548 ( .A(n8314), .B(n8313), .Z(n8246) );
  NANDN U8549 ( .A(n8235), .B(n8234), .Z(n8239) );
  NAND U8550 ( .A(n8237), .B(n8236), .Z(n8238) );
  AND U8551 ( .A(n8239), .B(n8238), .Z(n8245) );
  XNOR U8552 ( .A(n8246), .B(n8245), .Z(n8247) );
  XNOR U8553 ( .A(n8248), .B(n8247), .Z(n8317) );
  XNOR U8554 ( .A(sreg[354]), .B(n8317), .Z(n8319) );
  NANDN U8555 ( .A(sreg[353]), .B(n8240), .Z(n8244) );
  NAND U8556 ( .A(n8242), .B(n8241), .Z(n8243) );
  NAND U8557 ( .A(n8244), .B(n8243), .Z(n8318) );
  XNOR U8558 ( .A(n8319), .B(n8318), .Z(c[354]) );
  NANDN U8559 ( .A(n8246), .B(n8245), .Z(n8250) );
  NANDN U8560 ( .A(n8248), .B(n8247), .Z(n8249) );
  AND U8561 ( .A(n8250), .B(n8249), .Z(n8325) );
  NANDN U8562 ( .A(n8252), .B(n8251), .Z(n8256) );
  NAND U8563 ( .A(n8254), .B(n8253), .Z(n8255) );
  AND U8564 ( .A(n8256), .B(n8255), .Z(n8391) );
  NANDN U8565 ( .A(n8258), .B(n8257), .Z(n8262) );
  NANDN U8566 ( .A(n8260), .B(n8259), .Z(n8261) );
  AND U8567 ( .A(n8262), .B(n8261), .Z(n8357) );
  NAND U8568 ( .A(b[0]), .B(a[115]), .Z(n8263) );
  XNOR U8569 ( .A(b[1]), .B(n8263), .Z(n8265) );
  NANDN U8570 ( .A(b[0]), .B(a[114]), .Z(n8264) );
  NAND U8571 ( .A(n8265), .B(n8264), .Z(n8337) );
  NAND U8572 ( .A(n19808), .B(n8266), .Z(n8268) );
  XOR U8573 ( .A(b[13]), .B(a[103]), .Z(n8343) );
  NAND U8574 ( .A(n19768), .B(n8343), .Z(n8267) );
  AND U8575 ( .A(n8268), .B(n8267), .Z(n8335) );
  AND U8576 ( .A(b[15]), .B(a[99]), .Z(n8334) );
  XNOR U8577 ( .A(n8335), .B(n8334), .Z(n8336) );
  XNOR U8578 ( .A(n8337), .B(n8336), .Z(n8355) );
  NAND U8579 ( .A(n33), .B(n8269), .Z(n8271) );
  XOR U8580 ( .A(b[5]), .B(a[111]), .Z(n8346) );
  NAND U8581 ( .A(n19342), .B(n8346), .Z(n8270) );
  AND U8582 ( .A(n8271), .B(n8270), .Z(n8379) );
  NAND U8583 ( .A(n34), .B(n8272), .Z(n8274) );
  XOR U8584 ( .A(b[7]), .B(a[109]), .Z(n8349) );
  NAND U8585 ( .A(n19486), .B(n8349), .Z(n8273) );
  AND U8586 ( .A(n8274), .B(n8273), .Z(n8377) );
  NAND U8587 ( .A(n31), .B(n8275), .Z(n8277) );
  XOR U8588 ( .A(b[3]), .B(a[113]), .Z(n8352) );
  NAND U8589 ( .A(n32), .B(n8352), .Z(n8276) );
  NAND U8590 ( .A(n8277), .B(n8276), .Z(n8376) );
  XNOR U8591 ( .A(n8377), .B(n8376), .Z(n8378) );
  XOR U8592 ( .A(n8379), .B(n8378), .Z(n8356) );
  XOR U8593 ( .A(n8355), .B(n8356), .Z(n8358) );
  XOR U8594 ( .A(n8357), .B(n8358), .Z(n8329) );
  NANDN U8595 ( .A(n8279), .B(n8278), .Z(n8283) );
  OR U8596 ( .A(n8281), .B(n8280), .Z(n8282) );
  AND U8597 ( .A(n8283), .B(n8282), .Z(n8328) );
  XNOR U8598 ( .A(n8329), .B(n8328), .Z(n8331) );
  NAND U8599 ( .A(n8284), .B(n19724), .Z(n8286) );
  XOR U8600 ( .A(b[11]), .B(a[105]), .Z(n8361) );
  NAND U8601 ( .A(n19692), .B(n8361), .Z(n8285) );
  AND U8602 ( .A(n8286), .B(n8285), .Z(n8372) );
  NAND U8603 ( .A(n19838), .B(n8287), .Z(n8289) );
  XOR U8604 ( .A(b[15]), .B(a[101]), .Z(n8364) );
  NAND U8605 ( .A(n19805), .B(n8364), .Z(n8288) );
  AND U8606 ( .A(n8289), .B(n8288), .Z(n8371) );
  NAND U8607 ( .A(n35), .B(n8290), .Z(n8292) );
  XOR U8608 ( .A(b[9]), .B(a[107]), .Z(n8367) );
  NAND U8609 ( .A(n19598), .B(n8367), .Z(n8291) );
  NAND U8610 ( .A(n8292), .B(n8291), .Z(n8370) );
  XOR U8611 ( .A(n8371), .B(n8370), .Z(n8373) );
  XOR U8612 ( .A(n8372), .B(n8373), .Z(n8383) );
  NANDN U8613 ( .A(n8294), .B(n8293), .Z(n8298) );
  OR U8614 ( .A(n8296), .B(n8295), .Z(n8297) );
  AND U8615 ( .A(n8298), .B(n8297), .Z(n8382) );
  XNOR U8616 ( .A(n8383), .B(n8382), .Z(n8384) );
  NANDN U8617 ( .A(n8300), .B(n8299), .Z(n8304) );
  NANDN U8618 ( .A(n8302), .B(n8301), .Z(n8303) );
  NAND U8619 ( .A(n8304), .B(n8303), .Z(n8385) );
  XNOR U8620 ( .A(n8384), .B(n8385), .Z(n8330) );
  XOR U8621 ( .A(n8331), .B(n8330), .Z(n8389) );
  NANDN U8622 ( .A(n8306), .B(n8305), .Z(n8310) );
  NANDN U8623 ( .A(n8308), .B(n8307), .Z(n8309) );
  AND U8624 ( .A(n8310), .B(n8309), .Z(n8388) );
  XNOR U8625 ( .A(n8389), .B(n8388), .Z(n8390) );
  XOR U8626 ( .A(n8391), .B(n8390), .Z(n8323) );
  NANDN U8627 ( .A(n8312), .B(n8311), .Z(n8316) );
  NAND U8628 ( .A(n8314), .B(n8313), .Z(n8315) );
  AND U8629 ( .A(n8316), .B(n8315), .Z(n8322) );
  XNOR U8630 ( .A(n8323), .B(n8322), .Z(n8324) );
  XNOR U8631 ( .A(n8325), .B(n8324), .Z(n8394) );
  XNOR U8632 ( .A(sreg[355]), .B(n8394), .Z(n8396) );
  NANDN U8633 ( .A(sreg[354]), .B(n8317), .Z(n8321) );
  NAND U8634 ( .A(n8319), .B(n8318), .Z(n8320) );
  NAND U8635 ( .A(n8321), .B(n8320), .Z(n8395) );
  XNOR U8636 ( .A(n8396), .B(n8395), .Z(c[355]) );
  NANDN U8637 ( .A(n8323), .B(n8322), .Z(n8327) );
  NANDN U8638 ( .A(n8325), .B(n8324), .Z(n8326) );
  AND U8639 ( .A(n8327), .B(n8326), .Z(n8402) );
  NANDN U8640 ( .A(n8329), .B(n8328), .Z(n8333) );
  NAND U8641 ( .A(n8331), .B(n8330), .Z(n8332) );
  AND U8642 ( .A(n8333), .B(n8332), .Z(n8468) );
  NANDN U8643 ( .A(n8335), .B(n8334), .Z(n8339) );
  NANDN U8644 ( .A(n8337), .B(n8336), .Z(n8338) );
  AND U8645 ( .A(n8339), .B(n8338), .Z(n8434) );
  NAND U8646 ( .A(b[0]), .B(a[116]), .Z(n8340) );
  XNOR U8647 ( .A(b[1]), .B(n8340), .Z(n8342) );
  NANDN U8648 ( .A(b[0]), .B(a[115]), .Z(n8341) );
  NAND U8649 ( .A(n8342), .B(n8341), .Z(n8414) );
  NAND U8650 ( .A(n19808), .B(n8343), .Z(n8345) );
  XOR U8651 ( .A(b[13]), .B(a[104]), .Z(n8417) );
  NAND U8652 ( .A(n19768), .B(n8417), .Z(n8344) );
  AND U8653 ( .A(n8345), .B(n8344), .Z(n8412) );
  AND U8654 ( .A(b[15]), .B(a[100]), .Z(n8411) );
  XNOR U8655 ( .A(n8412), .B(n8411), .Z(n8413) );
  XNOR U8656 ( .A(n8414), .B(n8413), .Z(n8432) );
  NAND U8657 ( .A(n33), .B(n8346), .Z(n8348) );
  XOR U8658 ( .A(b[5]), .B(a[112]), .Z(n8423) );
  NAND U8659 ( .A(n19342), .B(n8423), .Z(n8347) );
  AND U8660 ( .A(n8348), .B(n8347), .Z(n8456) );
  NAND U8661 ( .A(n34), .B(n8349), .Z(n8351) );
  XOR U8662 ( .A(b[7]), .B(a[110]), .Z(n8426) );
  NAND U8663 ( .A(n19486), .B(n8426), .Z(n8350) );
  AND U8664 ( .A(n8351), .B(n8350), .Z(n8454) );
  NAND U8665 ( .A(n31), .B(n8352), .Z(n8354) );
  XOR U8666 ( .A(b[3]), .B(a[114]), .Z(n8429) );
  NAND U8667 ( .A(n32), .B(n8429), .Z(n8353) );
  NAND U8668 ( .A(n8354), .B(n8353), .Z(n8453) );
  XNOR U8669 ( .A(n8454), .B(n8453), .Z(n8455) );
  XOR U8670 ( .A(n8456), .B(n8455), .Z(n8433) );
  XOR U8671 ( .A(n8432), .B(n8433), .Z(n8435) );
  XOR U8672 ( .A(n8434), .B(n8435), .Z(n8406) );
  NANDN U8673 ( .A(n8356), .B(n8355), .Z(n8360) );
  OR U8674 ( .A(n8358), .B(n8357), .Z(n8359) );
  AND U8675 ( .A(n8360), .B(n8359), .Z(n8405) );
  XNOR U8676 ( .A(n8406), .B(n8405), .Z(n8408) );
  NAND U8677 ( .A(n8361), .B(n19724), .Z(n8363) );
  XOR U8678 ( .A(b[11]), .B(a[106]), .Z(n8438) );
  NAND U8679 ( .A(n19692), .B(n8438), .Z(n8362) );
  AND U8680 ( .A(n8363), .B(n8362), .Z(n8449) );
  NAND U8681 ( .A(n19838), .B(n8364), .Z(n8366) );
  XOR U8682 ( .A(b[15]), .B(a[102]), .Z(n8441) );
  NAND U8683 ( .A(n19805), .B(n8441), .Z(n8365) );
  AND U8684 ( .A(n8366), .B(n8365), .Z(n8448) );
  NAND U8685 ( .A(n35), .B(n8367), .Z(n8369) );
  XOR U8686 ( .A(b[9]), .B(a[108]), .Z(n8444) );
  NAND U8687 ( .A(n19598), .B(n8444), .Z(n8368) );
  NAND U8688 ( .A(n8369), .B(n8368), .Z(n8447) );
  XOR U8689 ( .A(n8448), .B(n8447), .Z(n8450) );
  XOR U8690 ( .A(n8449), .B(n8450), .Z(n8460) );
  NANDN U8691 ( .A(n8371), .B(n8370), .Z(n8375) );
  OR U8692 ( .A(n8373), .B(n8372), .Z(n8374) );
  AND U8693 ( .A(n8375), .B(n8374), .Z(n8459) );
  XNOR U8694 ( .A(n8460), .B(n8459), .Z(n8461) );
  NANDN U8695 ( .A(n8377), .B(n8376), .Z(n8381) );
  NANDN U8696 ( .A(n8379), .B(n8378), .Z(n8380) );
  NAND U8697 ( .A(n8381), .B(n8380), .Z(n8462) );
  XNOR U8698 ( .A(n8461), .B(n8462), .Z(n8407) );
  XOR U8699 ( .A(n8408), .B(n8407), .Z(n8466) );
  NANDN U8700 ( .A(n8383), .B(n8382), .Z(n8387) );
  NANDN U8701 ( .A(n8385), .B(n8384), .Z(n8386) );
  AND U8702 ( .A(n8387), .B(n8386), .Z(n8465) );
  XNOR U8703 ( .A(n8466), .B(n8465), .Z(n8467) );
  XOR U8704 ( .A(n8468), .B(n8467), .Z(n8400) );
  NANDN U8705 ( .A(n8389), .B(n8388), .Z(n8393) );
  NAND U8706 ( .A(n8391), .B(n8390), .Z(n8392) );
  AND U8707 ( .A(n8393), .B(n8392), .Z(n8399) );
  XNOR U8708 ( .A(n8400), .B(n8399), .Z(n8401) );
  XNOR U8709 ( .A(n8402), .B(n8401), .Z(n8471) );
  XNOR U8710 ( .A(sreg[356]), .B(n8471), .Z(n8473) );
  NANDN U8711 ( .A(sreg[355]), .B(n8394), .Z(n8398) );
  NAND U8712 ( .A(n8396), .B(n8395), .Z(n8397) );
  NAND U8713 ( .A(n8398), .B(n8397), .Z(n8472) );
  XNOR U8714 ( .A(n8473), .B(n8472), .Z(c[356]) );
  NANDN U8715 ( .A(n8400), .B(n8399), .Z(n8404) );
  NANDN U8716 ( .A(n8402), .B(n8401), .Z(n8403) );
  AND U8717 ( .A(n8404), .B(n8403), .Z(n8479) );
  NANDN U8718 ( .A(n8406), .B(n8405), .Z(n8410) );
  NAND U8719 ( .A(n8408), .B(n8407), .Z(n8409) );
  AND U8720 ( .A(n8410), .B(n8409), .Z(n8545) );
  NANDN U8721 ( .A(n8412), .B(n8411), .Z(n8416) );
  NANDN U8722 ( .A(n8414), .B(n8413), .Z(n8415) );
  AND U8723 ( .A(n8416), .B(n8415), .Z(n8511) );
  NAND U8724 ( .A(n19808), .B(n8417), .Z(n8419) );
  XOR U8725 ( .A(b[13]), .B(a[105]), .Z(n8497) );
  NAND U8726 ( .A(n19768), .B(n8497), .Z(n8418) );
  AND U8727 ( .A(n8419), .B(n8418), .Z(n8489) );
  AND U8728 ( .A(b[15]), .B(a[101]), .Z(n8488) );
  XNOR U8729 ( .A(n8489), .B(n8488), .Z(n8490) );
  NAND U8730 ( .A(b[0]), .B(a[117]), .Z(n8420) );
  XNOR U8731 ( .A(b[1]), .B(n8420), .Z(n8422) );
  NANDN U8732 ( .A(b[0]), .B(a[116]), .Z(n8421) );
  NAND U8733 ( .A(n8422), .B(n8421), .Z(n8491) );
  XNOR U8734 ( .A(n8490), .B(n8491), .Z(n8509) );
  NAND U8735 ( .A(n33), .B(n8423), .Z(n8425) );
  XOR U8736 ( .A(b[5]), .B(a[113]), .Z(n8500) );
  NAND U8737 ( .A(n19342), .B(n8500), .Z(n8424) );
  AND U8738 ( .A(n8425), .B(n8424), .Z(n8533) );
  NAND U8739 ( .A(n34), .B(n8426), .Z(n8428) );
  XOR U8740 ( .A(b[7]), .B(a[111]), .Z(n8503) );
  NAND U8741 ( .A(n19486), .B(n8503), .Z(n8427) );
  AND U8742 ( .A(n8428), .B(n8427), .Z(n8531) );
  NAND U8743 ( .A(n31), .B(n8429), .Z(n8431) );
  XOR U8744 ( .A(b[3]), .B(a[115]), .Z(n8506) );
  NAND U8745 ( .A(n32), .B(n8506), .Z(n8430) );
  NAND U8746 ( .A(n8431), .B(n8430), .Z(n8530) );
  XNOR U8747 ( .A(n8531), .B(n8530), .Z(n8532) );
  XOR U8748 ( .A(n8533), .B(n8532), .Z(n8510) );
  XOR U8749 ( .A(n8509), .B(n8510), .Z(n8512) );
  XOR U8750 ( .A(n8511), .B(n8512), .Z(n8483) );
  NANDN U8751 ( .A(n8433), .B(n8432), .Z(n8437) );
  OR U8752 ( .A(n8435), .B(n8434), .Z(n8436) );
  AND U8753 ( .A(n8437), .B(n8436), .Z(n8482) );
  XNOR U8754 ( .A(n8483), .B(n8482), .Z(n8485) );
  NAND U8755 ( .A(n8438), .B(n19724), .Z(n8440) );
  XOR U8756 ( .A(b[11]), .B(a[107]), .Z(n8515) );
  NAND U8757 ( .A(n19692), .B(n8515), .Z(n8439) );
  AND U8758 ( .A(n8440), .B(n8439), .Z(n8526) );
  NAND U8759 ( .A(n19838), .B(n8441), .Z(n8443) );
  XOR U8760 ( .A(b[15]), .B(a[103]), .Z(n8518) );
  NAND U8761 ( .A(n19805), .B(n8518), .Z(n8442) );
  AND U8762 ( .A(n8443), .B(n8442), .Z(n8525) );
  NAND U8763 ( .A(n35), .B(n8444), .Z(n8446) );
  XOR U8764 ( .A(b[9]), .B(a[109]), .Z(n8521) );
  NAND U8765 ( .A(n19598), .B(n8521), .Z(n8445) );
  NAND U8766 ( .A(n8446), .B(n8445), .Z(n8524) );
  XOR U8767 ( .A(n8525), .B(n8524), .Z(n8527) );
  XOR U8768 ( .A(n8526), .B(n8527), .Z(n8537) );
  NANDN U8769 ( .A(n8448), .B(n8447), .Z(n8452) );
  OR U8770 ( .A(n8450), .B(n8449), .Z(n8451) );
  AND U8771 ( .A(n8452), .B(n8451), .Z(n8536) );
  XNOR U8772 ( .A(n8537), .B(n8536), .Z(n8538) );
  NANDN U8773 ( .A(n8454), .B(n8453), .Z(n8458) );
  NANDN U8774 ( .A(n8456), .B(n8455), .Z(n8457) );
  NAND U8775 ( .A(n8458), .B(n8457), .Z(n8539) );
  XNOR U8776 ( .A(n8538), .B(n8539), .Z(n8484) );
  XOR U8777 ( .A(n8485), .B(n8484), .Z(n8543) );
  NANDN U8778 ( .A(n8460), .B(n8459), .Z(n8464) );
  NANDN U8779 ( .A(n8462), .B(n8461), .Z(n8463) );
  AND U8780 ( .A(n8464), .B(n8463), .Z(n8542) );
  XNOR U8781 ( .A(n8543), .B(n8542), .Z(n8544) );
  XOR U8782 ( .A(n8545), .B(n8544), .Z(n8477) );
  NANDN U8783 ( .A(n8466), .B(n8465), .Z(n8470) );
  NAND U8784 ( .A(n8468), .B(n8467), .Z(n8469) );
  AND U8785 ( .A(n8470), .B(n8469), .Z(n8476) );
  XNOR U8786 ( .A(n8477), .B(n8476), .Z(n8478) );
  XNOR U8787 ( .A(n8479), .B(n8478), .Z(n8548) );
  XNOR U8788 ( .A(sreg[357]), .B(n8548), .Z(n8550) );
  NANDN U8789 ( .A(sreg[356]), .B(n8471), .Z(n8475) );
  NAND U8790 ( .A(n8473), .B(n8472), .Z(n8474) );
  NAND U8791 ( .A(n8475), .B(n8474), .Z(n8549) );
  XNOR U8792 ( .A(n8550), .B(n8549), .Z(c[357]) );
  NANDN U8793 ( .A(n8477), .B(n8476), .Z(n8481) );
  NANDN U8794 ( .A(n8479), .B(n8478), .Z(n8480) );
  AND U8795 ( .A(n8481), .B(n8480), .Z(n8556) );
  NANDN U8796 ( .A(n8483), .B(n8482), .Z(n8487) );
  NAND U8797 ( .A(n8485), .B(n8484), .Z(n8486) );
  AND U8798 ( .A(n8487), .B(n8486), .Z(n8622) );
  NANDN U8799 ( .A(n8489), .B(n8488), .Z(n8493) );
  NANDN U8800 ( .A(n8491), .B(n8490), .Z(n8492) );
  AND U8801 ( .A(n8493), .B(n8492), .Z(n8609) );
  NAND U8802 ( .A(b[0]), .B(a[118]), .Z(n8494) );
  XNOR U8803 ( .A(b[1]), .B(n8494), .Z(n8496) );
  NANDN U8804 ( .A(b[0]), .B(a[117]), .Z(n8495) );
  NAND U8805 ( .A(n8496), .B(n8495), .Z(n8589) );
  NAND U8806 ( .A(n19808), .B(n8497), .Z(n8499) );
  XOR U8807 ( .A(b[13]), .B(a[106]), .Z(n8595) );
  NAND U8808 ( .A(n19768), .B(n8595), .Z(n8498) );
  AND U8809 ( .A(n8499), .B(n8498), .Z(n8587) );
  AND U8810 ( .A(b[15]), .B(a[102]), .Z(n8586) );
  XNOR U8811 ( .A(n8587), .B(n8586), .Z(n8588) );
  XNOR U8812 ( .A(n8589), .B(n8588), .Z(n8607) );
  NAND U8813 ( .A(n33), .B(n8500), .Z(n8502) );
  XOR U8814 ( .A(b[5]), .B(a[114]), .Z(n8598) );
  NAND U8815 ( .A(n19342), .B(n8598), .Z(n8501) );
  AND U8816 ( .A(n8502), .B(n8501), .Z(n8583) );
  NAND U8817 ( .A(n34), .B(n8503), .Z(n8505) );
  XOR U8818 ( .A(b[7]), .B(a[112]), .Z(n8601) );
  NAND U8819 ( .A(n19486), .B(n8601), .Z(n8504) );
  AND U8820 ( .A(n8505), .B(n8504), .Z(n8581) );
  NAND U8821 ( .A(n31), .B(n8506), .Z(n8508) );
  XOR U8822 ( .A(b[3]), .B(a[116]), .Z(n8604) );
  NAND U8823 ( .A(n32), .B(n8604), .Z(n8507) );
  NAND U8824 ( .A(n8508), .B(n8507), .Z(n8580) );
  XNOR U8825 ( .A(n8581), .B(n8580), .Z(n8582) );
  XOR U8826 ( .A(n8583), .B(n8582), .Z(n8608) );
  XOR U8827 ( .A(n8607), .B(n8608), .Z(n8610) );
  XOR U8828 ( .A(n8609), .B(n8610), .Z(n8560) );
  NANDN U8829 ( .A(n8510), .B(n8509), .Z(n8514) );
  OR U8830 ( .A(n8512), .B(n8511), .Z(n8513) );
  AND U8831 ( .A(n8514), .B(n8513), .Z(n8559) );
  XNOR U8832 ( .A(n8560), .B(n8559), .Z(n8562) );
  NAND U8833 ( .A(n8515), .B(n19724), .Z(n8517) );
  XOR U8834 ( .A(b[11]), .B(a[108]), .Z(n8565) );
  NAND U8835 ( .A(n19692), .B(n8565), .Z(n8516) );
  AND U8836 ( .A(n8517), .B(n8516), .Z(n8576) );
  NAND U8837 ( .A(n19838), .B(n8518), .Z(n8520) );
  XOR U8838 ( .A(b[15]), .B(a[104]), .Z(n8568) );
  NAND U8839 ( .A(n19805), .B(n8568), .Z(n8519) );
  AND U8840 ( .A(n8520), .B(n8519), .Z(n8575) );
  NAND U8841 ( .A(n35), .B(n8521), .Z(n8523) );
  XOR U8842 ( .A(b[9]), .B(a[110]), .Z(n8571) );
  NAND U8843 ( .A(n19598), .B(n8571), .Z(n8522) );
  NAND U8844 ( .A(n8523), .B(n8522), .Z(n8574) );
  XOR U8845 ( .A(n8575), .B(n8574), .Z(n8577) );
  XOR U8846 ( .A(n8576), .B(n8577), .Z(n8614) );
  NANDN U8847 ( .A(n8525), .B(n8524), .Z(n8529) );
  OR U8848 ( .A(n8527), .B(n8526), .Z(n8528) );
  AND U8849 ( .A(n8529), .B(n8528), .Z(n8613) );
  XNOR U8850 ( .A(n8614), .B(n8613), .Z(n8615) );
  NANDN U8851 ( .A(n8531), .B(n8530), .Z(n8535) );
  NANDN U8852 ( .A(n8533), .B(n8532), .Z(n8534) );
  NAND U8853 ( .A(n8535), .B(n8534), .Z(n8616) );
  XNOR U8854 ( .A(n8615), .B(n8616), .Z(n8561) );
  XOR U8855 ( .A(n8562), .B(n8561), .Z(n8620) );
  NANDN U8856 ( .A(n8537), .B(n8536), .Z(n8541) );
  NANDN U8857 ( .A(n8539), .B(n8538), .Z(n8540) );
  AND U8858 ( .A(n8541), .B(n8540), .Z(n8619) );
  XNOR U8859 ( .A(n8620), .B(n8619), .Z(n8621) );
  XOR U8860 ( .A(n8622), .B(n8621), .Z(n8554) );
  NANDN U8861 ( .A(n8543), .B(n8542), .Z(n8547) );
  NAND U8862 ( .A(n8545), .B(n8544), .Z(n8546) );
  AND U8863 ( .A(n8547), .B(n8546), .Z(n8553) );
  XNOR U8864 ( .A(n8554), .B(n8553), .Z(n8555) );
  XNOR U8865 ( .A(n8556), .B(n8555), .Z(n8625) );
  XNOR U8866 ( .A(sreg[358]), .B(n8625), .Z(n8627) );
  NANDN U8867 ( .A(sreg[357]), .B(n8548), .Z(n8552) );
  NAND U8868 ( .A(n8550), .B(n8549), .Z(n8551) );
  NAND U8869 ( .A(n8552), .B(n8551), .Z(n8626) );
  XNOR U8870 ( .A(n8627), .B(n8626), .Z(c[358]) );
  NANDN U8871 ( .A(n8554), .B(n8553), .Z(n8558) );
  NANDN U8872 ( .A(n8556), .B(n8555), .Z(n8557) );
  AND U8873 ( .A(n8558), .B(n8557), .Z(n8633) );
  NANDN U8874 ( .A(n8560), .B(n8559), .Z(n8564) );
  NAND U8875 ( .A(n8562), .B(n8561), .Z(n8563) );
  AND U8876 ( .A(n8564), .B(n8563), .Z(n8699) );
  NAND U8877 ( .A(n8565), .B(n19724), .Z(n8567) );
  XOR U8878 ( .A(b[11]), .B(a[109]), .Z(n8669) );
  NAND U8879 ( .A(n19692), .B(n8669), .Z(n8566) );
  AND U8880 ( .A(n8567), .B(n8566), .Z(n8680) );
  NAND U8881 ( .A(n19838), .B(n8568), .Z(n8570) );
  XOR U8882 ( .A(b[15]), .B(a[105]), .Z(n8672) );
  NAND U8883 ( .A(n19805), .B(n8672), .Z(n8569) );
  AND U8884 ( .A(n8570), .B(n8569), .Z(n8679) );
  NAND U8885 ( .A(n35), .B(n8571), .Z(n8573) );
  XOR U8886 ( .A(b[9]), .B(a[111]), .Z(n8675) );
  NAND U8887 ( .A(n19598), .B(n8675), .Z(n8572) );
  NAND U8888 ( .A(n8573), .B(n8572), .Z(n8678) );
  XOR U8889 ( .A(n8679), .B(n8678), .Z(n8681) );
  XOR U8890 ( .A(n8680), .B(n8681), .Z(n8691) );
  NANDN U8891 ( .A(n8575), .B(n8574), .Z(n8579) );
  OR U8892 ( .A(n8577), .B(n8576), .Z(n8578) );
  AND U8893 ( .A(n8579), .B(n8578), .Z(n8690) );
  XNOR U8894 ( .A(n8691), .B(n8690), .Z(n8692) );
  NANDN U8895 ( .A(n8581), .B(n8580), .Z(n8585) );
  NANDN U8896 ( .A(n8583), .B(n8582), .Z(n8584) );
  NAND U8897 ( .A(n8585), .B(n8584), .Z(n8693) );
  XNOR U8898 ( .A(n8692), .B(n8693), .Z(n8639) );
  NANDN U8899 ( .A(n8587), .B(n8586), .Z(n8591) );
  NANDN U8900 ( .A(n8589), .B(n8588), .Z(n8590) );
  AND U8901 ( .A(n8591), .B(n8590), .Z(n8665) );
  NAND U8902 ( .A(b[0]), .B(a[119]), .Z(n8592) );
  XNOR U8903 ( .A(b[1]), .B(n8592), .Z(n8594) );
  NANDN U8904 ( .A(b[0]), .B(a[118]), .Z(n8593) );
  NAND U8905 ( .A(n8594), .B(n8593), .Z(n8645) );
  NAND U8906 ( .A(n19808), .B(n8595), .Z(n8597) );
  XOR U8907 ( .A(b[13]), .B(a[107]), .Z(n8651) );
  NAND U8908 ( .A(n19768), .B(n8651), .Z(n8596) );
  AND U8909 ( .A(n8597), .B(n8596), .Z(n8643) );
  AND U8910 ( .A(b[15]), .B(a[103]), .Z(n8642) );
  XNOR U8911 ( .A(n8643), .B(n8642), .Z(n8644) );
  XNOR U8912 ( .A(n8645), .B(n8644), .Z(n8663) );
  NAND U8913 ( .A(n33), .B(n8598), .Z(n8600) );
  XOR U8914 ( .A(b[5]), .B(a[115]), .Z(n8654) );
  NAND U8915 ( .A(n19342), .B(n8654), .Z(n8599) );
  AND U8916 ( .A(n8600), .B(n8599), .Z(n8687) );
  NAND U8917 ( .A(n34), .B(n8601), .Z(n8603) );
  XOR U8918 ( .A(b[7]), .B(a[113]), .Z(n8657) );
  NAND U8919 ( .A(n19486), .B(n8657), .Z(n8602) );
  AND U8920 ( .A(n8603), .B(n8602), .Z(n8685) );
  NAND U8921 ( .A(n31), .B(n8604), .Z(n8606) );
  XOR U8922 ( .A(b[3]), .B(a[117]), .Z(n8660) );
  NAND U8923 ( .A(n32), .B(n8660), .Z(n8605) );
  NAND U8924 ( .A(n8606), .B(n8605), .Z(n8684) );
  XNOR U8925 ( .A(n8685), .B(n8684), .Z(n8686) );
  XOR U8926 ( .A(n8687), .B(n8686), .Z(n8664) );
  XOR U8927 ( .A(n8663), .B(n8664), .Z(n8666) );
  XOR U8928 ( .A(n8665), .B(n8666), .Z(n8637) );
  NANDN U8929 ( .A(n8608), .B(n8607), .Z(n8612) );
  OR U8930 ( .A(n8610), .B(n8609), .Z(n8611) );
  AND U8931 ( .A(n8612), .B(n8611), .Z(n8636) );
  XNOR U8932 ( .A(n8637), .B(n8636), .Z(n8638) );
  XOR U8933 ( .A(n8639), .B(n8638), .Z(n8697) );
  NANDN U8934 ( .A(n8614), .B(n8613), .Z(n8618) );
  NANDN U8935 ( .A(n8616), .B(n8615), .Z(n8617) );
  AND U8936 ( .A(n8618), .B(n8617), .Z(n8696) );
  XNOR U8937 ( .A(n8697), .B(n8696), .Z(n8698) );
  XOR U8938 ( .A(n8699), .B(n8698), .Z(n8631) );
  NANDN U8939 ( .A(n8620), .B(n8619), .Z(n8624) );
  NAND U8940 ( .A(n8622), .B(n8621), .Z(n8623) );
  AND U8941 ( .A(n8624), .B(n8623), .Z(n8630) );
  XNOR U8942 ( .A(n8631), .B(n8630), .Z(n8632) );
  XNOR U8943 ( .A(n8633), .B(n8632), .Z(n8702) );
  XNOR U8944 ( .A(sreg[359]), .B(n8702), .Z(n8704) );
  NANDN U8945 ( .A(sreg[358]), .B(n8625), .Z(n8629) );
  NAND U8946 ( .A(n8627), .B(n8626), .Z(n8628) );
  NAND U8947 ( .A(n8629), .B(n8628), .Z(n8703) );
  XNOR U8948 ( .A(n8704), .B(n8703), .Z(c[359]) );
  NANDN U8949 ( .A(n8631), .B(n8630), .Z(n8635) );
  NANDN U8950 ( .A(n8633), .B(n8632), .Z(n8634) );
  AND U8951 ( .A(n8635), .B(n8634), .Z(n8710) );
  NANDN U8952 ( .A(n8637), .B(n8636), .Z(n8641) );
  NAND U8953 ( .A(n8639), .B(n8638), .Z(n8640) );
  AND U8954 ( .A(n8641), .B(n8640), .Z(n8776) );
  NANDN U8955 ( .A(n8643), .B(n8642), .Z(n8647) );
  NANDN U8956 ( .A(n8645), .B(n8644), .Z(n8646) );
  AND U8957 ( .A(n8647), .B(n8646), .Z(n8742) );
  NAND U8958 ( .A(b[0]), .B(a[120]), .Z(n8648) );
  XNOR U8959 ( .A(b[1]), .B(n8648), .Z(n8650) );
  NANDN U8960 ( .A(b[0]), .B(a[119]), .Z(n8649) );
  NAND U8961 ( .A(n8650), .B(n8649), .Z(n8722) );
  NAND U8962 ( .A(n19808), .B(n8651), .Z(n8653) );
  XOR U8963 ( .A(b[13]), .B(a[108]), .Z(n8728) );
  NAND U8964 ( .A(n19768), .B(n8728), .Z(n8652) );
  AND U8965 ( .A(n8653), .B(n8652), .Z(n8720) );
  AND U8966 ( .A(b[15]), .B(a[104]), .Z(n8719) );
  XNOR U8967 ( .A(n8720), .B(n8719), .Z(n8721) );
  XNOR U8968 ( .A(n8722), .B(n8721), .Z(n8740) );
  NAND U8969 ( .A(n33), .B(n8654), .Z(n8656) );
  XOR U8970 ( .A(b[5]), .B(a[116]), .Z(n8731) );
  NAND U8971 ( .A(n19342), .B(n8731), .Z(n8655) );
  AND U8972 ( .A(n8656), .B(n8655), .Z(n8764) );
  NAND U8973 ( .A(n34), .B(n8657), .Z(n8659) );
  XOR U8974 ( .A(b[7]), .B(a[114]), .Z(n8734) );
  NAND U8975 ( .A(n19486), .B(n8734), .Z(n8658) );
  AND U8976 ( .A(n8659), .B(n8658), .Z(n8762) );
  NAND U8977 ( .A(n31), .B(n8660), .Z(n8662) );
  XOR U8978 ( .A(b[3]), .B(a[118]), .Z(n8737) );
  NAND U8979 ( .A(n32), .B(n8737), .Z(n8661) );
  NAND U8980 ( .A(n8662), .B(n8661), .Z(n8761) );
  XNOR U8981 ( .A(n8762), .B(n8761), .Z(n8763) );
  XOR U8982 ( .A(n8764), .B(n8763), .Z(n8741) );
  XOR U8983 ( .A(n8740), .B(n8741), .Z(n8743) );
  XOR U8984 ( .A(n8742), .B(n8743), .Z(n8714) );
  NANDN U8985 ( .A(n8664), .B(n8663), .Z(n8668) );
  OR U8986 ( .A(n8666), .B(n8665), .Z(n8667) );
  AND U8987 ( .A(n8668), .B(n8667), .Z(n8713) );
  XNOR U8988 ( .A(n8714), .B(n8713), .Z(n8716) );
  NAND U8989 ( .A(n8669), .B(n19724), .Z(n8671) );
  XOR U8990 ( .A(b[11]), .B(a[110]), .Z(n8746) );
  NAND U8991 ( .A(n19692), .B(n8746), .Z(n8670) );
  AND U8992 ( .A(n8671), .B(n8670), .Z(n8757) );
  NAND U8993 ( .A(n19838), .B(n8672), .Z(n8674) );
  XOR U8994 ( .A(b[15]), .B(a[106]), .Z(n8749) );
  NAND U8995 ( .A(n19805), .B(n8749), .Z(n8673) );
  AND U8996 ( .A(n8674), .B(n8673), .Z(n8756) );
  NAND U8997 ( .A(n35), .B(n8675), .Z(n8677) );
  XOR U8998 ( .A(b[9]), .B(a[112]), .Z(n8752) );
  NAND U8999 ( .A(n19598), .B(n8752), .Z(n8676) );
  NAND U9000 ( .A(n8677), .B(n8676), .Z(n8755) );
  XOR U9001 ( .A(n8756), .B(n8755), .Z(n8758) );
  XOR U9002 ( .A(n8757), .B(n8758), .Z(n8768) );
  NANDN U9003 ( .A(n8679), .B(n8678), .Z(n8683) );
  OR U9004 ( .A(n8681), .B(n8680), .Z(n8682) );
  AND U9005 ( .A(n8683), .B(n8682), .Z(n8767) );
  XNOR U9006 ( .A(n8768), .B(n8767), .Z(n8769) );
  NANDN U9007 ( .A(n8685), .B(n8684), .Z(n8689) );
  NANDN U9008 ( .A(n8687), .B(n8686), .Z(n8688) );
  NAND U9009 ( .A(n8689), .B(n8688), .Z(n8770) );
  XNOR U9010 ( .A(n8769), .B(n8770), .Z(n8715) );
  XOR U9011 ( .A(n8716), .B(n8715), .Z(n8774) );
  NANDN U9012 ( .A(n8691), .B(n8690), .Z(n8695) );
  NANDN U9013 ( .A(n8693), .B(n8692), .Z(n8694) );
  AND U9014 ( .A(n8695), .B(n8694), .Z(n8773) );
  XNOR U9015 ( .A(n8774), .B(n8773), .Z(n8775) );
  XOR U9016 ( .A(n8776), .B(n8775), .Z(n8708) );
  NANDN U9017 ( .A(n8697), .B(n8696), .Z(n8701) );
  NAND U9018 ( .A(n8699), .B(n8698), .Z(n8700) );
  AND U9019 ( .A(n8701), .B(n8700), .Z(n8707) );
  XNOR U9020 ( .A(n8708), .B(n8707), .Z(n8709) );
  XNOR U9021 ( .A(n8710), .B(n8709), .Z(n8779) );
  XNOR U9022 ( .A(sreg[360]), .B(n8779), .Z(n8781) );
  NANDN U9023 ( .A(sreg[359]), .B(n8702), .Z(n8706) );
  NAND U9024 ( .A(n8704), .B(n8703), .Z(n8705) );
  NAND U9025 ( .A(n8706), .B(n8705), .Z(n8780) );
  XNOR U9026 ( .A(n8781), .B(n8780), .Z(c[360]) );
  NANDN U9027 ( .A(n8708), .B(n8707), .Z(n8712) );
  NANDN U9028 ( .A(n8710), .B(n8709), .Z(n8711) );
  AND U9029 ( .A(n8712), .B(n8711), .Z(n8787) );
  NANDN U9030 ( .A(n8714), .B(n8713), .Z(n8718) );
  NAND U9031 ( .A(n8716), .B(n8715), .Z(n8717) );
  AND U9032 ( .A(n8718), .B(n8717), .Z(n8853) );
  NANDN U9033 ( .A(n8720), .B(n8719), .Z(n8724) );
  NANDN U9034 ( .A(n8722), .B(n8721), .Z(n8723) );
  AND U9035 ( .A(n8724), .B(n8723), .Z(n8819) );
  NAND U9036 ( .A(b[0]), .B(a[121]), .Z(n8725) );
  XNOR U9037 ( .A(b[1]), .B(n8725), .Z(n8727) );
  NANDN U9038 ( .A(b[0]), .B(a[120]), .Z(n8726) );
  NAND U9039 ( .A(n8727), .B(n8726), .Z(n8799) );
  NAND U9040 ( .A(n19808), .B(n8728), .Z(n8730) );
  XOR U9041 ( .A(b[13]), .B(a[109]), .Z(n8805) );
  NAND U9042 ( .A(n19768), .B(n8805), .Z(n8729) );
  AND U9043 ( .A(n8730), .B(n8729), .Z(n8797) );
  AND U9044 ( .A(b[15]), .B(a[105]), .Z(n8796) );
  XNOR U9045 ( .A(n8797), .B(n8796), .Z(n8798) );
  XNOR U9046 ( .A(n8799), .B(n8798), .Z(n8817) );
  NAND U9047 ( .A(n33), .B(n8731), .Z(n8733) );
  XOR U9048 ( .A(b[5]), .B(a[117]), .Z(n8808) );
  NAND U9049 ( .A(n19342), .B(n8808), .Z(n8732) );
  AND U9050 ( .A(n8733), .B(n8732), .Z(n8841) );
  NAND U9051 ( .A(n34), .B(n8734), .Z(n8736) );
  XOR U9052 ( .A(b[7]), .B(a[115]), .Z(n8811) );
  NAND U9053 ( .A(n19486), .B(n8811), .Z(n8735) );
  AND U9054 ( .A(n8736), .B(n8735), .Z(n8839) );
  NAND U9055 ( .A(n31), .B(n8737), .Z(n8739) );
  XOR U9056 ( .A(b[3]), .B(a[119]), .Z(n8814) );
  NAND U9057 ( .A(n32), .B(n8814), .Z(n8738) );
  NAND U9058 ( .A(n8739), .B(n8738), .Z(n8838) );
  XNOR U9059 ( .A(n8839), .B(n8838), .Z(n8840) );
  XOR U9060 ( .A(n8841), .B(n8840), .Z(n8818) );
  XOR U9061 ( .A(n8817), .B(n8818), .Z(n8820) );
  XOR U9062 ( .A(n8819), .B(n8820), .Z(n8791) );
  NANDN U9063 ( .A(n8741), .B(n8740), .Z(n8745) );
  OR U9064 ( .A(n8743), .B(n8742), .Z(n8744) );
  AND U9065 ( .A(n8745), .B(n8744), .Z(n8790) );
  XNOR U9066 ( .A(n8791), .B(n8790), .Z(n8793) );
  NAND U9067 ( .A(n8746), .B(n19724), .Z(n8748) );
  XOR U9068 ( .A(b[11]), .B(a[111]), .Z(n8823) );
  NAND U9069 ( .A(n19692), .B(n8823), .Z(n8747) );
  AND U9070 ( .A(n8748), .B(n8747), .Z(n8834) );
  NAND U9071 ( .A(n19838), .B(n8749), .Z(n8751) );
  XOR U9072 ( .A(b[15]), .B(a[107]), .Z(n8826) );
  NAND U9073 ( .A(n19805), .B(n8826), .Z(n8750) );
  AND U9074 ( .A(n8751), .B(n8750), .Z(n8833) );
  NAND U9075 ( .A(n35), .B(n8752), .Z(n8754) );
  XOR U9076 ( .A(b[9]), .B(a[113]), .Z(n8829) );
  NAND U9077 ( .A(n19598), .B(n8829), .Z(n8753) );
  NAND U9078 ( .A(n8754), .B(n8753), .Z(n8832) );
  XOR U9079 ( .A(n8833), .B(n8832), .Z(n8835) );
  XOR U9080 ( .A(n8834), .B(n8835), .Z(n8845) );
  NANDN U9081 ( .A(n8756), .B(n8755), .Z(n8760) );
  OR U9082 ( .A(n8758), .B(n8757), .Z(n8759) );
  AND U9083 ( .A(n8760), .B(n8759), .Z(n8844) );
  XNOR U9084 ( .A(n8845), .B(n8844), .Z(n8846) );
  NANDN U9085 ( .A(n8762), .B(n8761), .Z(n8766) );
  NANDN U9086 ( .A(n8764), .B(n8763), .Z(n8765) );
  NAND U9087 ( .A(n8766), .B(n8765), .Z(n8847) );
  XNOR U9088 ( .A(n8846), .B(n8847), .Z(n8792) );
  XOR U9089 ( .A(n8793), .B(n8792), .Z(n8851) );
  NANDN U9090 ( .A(n8768), .B(n8767), .Z(n8772) );
  NANDN U9091 ( .A(n8770), .B(n8769), .Z(n8771) );
  AND U9092 ( .A(n8772), .B(n8771), .Z(n8850) );
  XNOR U9093 ( .A(n8851), .B(n8850), .Z(n8852) );
  XOR U9094 ( .A(n8853), .B(n8852), .Z(n8785) );
  NANDN U9095 ( .A(n8774), .B(n8773), .Z(n8778) );
  NAND U9096 ( .A(n8776), .B(n8775), .Z(n8777) );
  AND U9097 ( .A(n8778), .B(n8777), .Z(n8784) );
  XNOR U9098 ( .A(n8785), .B(n8784), .Z(n8786) );
  XNOR U9099 ( .A(n8787), .B(n8786), .Z(n8856) );
  XNOR U9100 ( .A(sreg[361]), .B(n8856), .Z(n8858) );
  NANDN U9101 ( .A(sreg[360]), .B(n8779), .Z(n8783) );
  NAND U9102 ( .A(n8781), .B(n8780), .Z(n8782) );
  NAND U9103 ( .A(n8783), .B(n8782), .Z(n8857) );
  XNOR U9104 ( .A(n8858), .B(n8857), .Z(c[361]) );
  NANDN U9105 ( .A(n8785), .B(n8784), .Z(n8789) );
  NANDN U9106 ( .A(n8787), .B(n8786), .Z(n8788) );
  AND U9107 ( .A(n8789), .B(n8788), .Z(n8864) );
  NANDN U9108 ( .A(n8791), .B(n8790), .Z(n8795) );
  NAND U9109 ( .A(n8793), .B(n8792), .Z(n8794) );
  AND U9110 ( .A(n8795), .B(n8794), .Z(n8930) );
  NANDN U9111 ( .A(n8797), .B(n8796), .Z(n8801) );
  NANDN U9112 ( .A(n8799), .B(n8798), .Z(n8800) );
  AND U9113 ( .A(n8801), .B(n8800), .Z(n8896) );
  NAND U9114 ( .A(b[0]), .B(a[122]), .Z(n8802) );
  XNOR U9115 ( .A(b[1]), .B(n8802), .Z(n8804) );
  NANDN U9116 ( .A(b[0]), .B(a[121]), .Z(n8803) );
  NAND U9117 ( .A(n8804), .B(n8803), .Z(n8876) );
  NAND U9118 ( .A(n19808), .B(n8805), .Z(n8807) );
  XOR U9119 ( .A(b[13]), .B(a[110]), .Z(n8882) );
  NAND U9120 ( .A(n19768), .B(n8882), .Z(n8806) );
  AND U9121 ( .A(n8807), .B(n8806), .Z(n8874) );
  AND U9122 ( .A(b[15]), .B(a[106]), .Z(n8873) );
  XNOR U9123 ( .A(n8874), .B(n8873), .Z(n8875) );
  XNOR U9124 ( .A(n8876), .B(n8875), .Z(n8894) );
  NAND U9125 ( .A(n33), .B(n8808), .Z(n8810) );
  XOR U9126 ( .A(b[5]), .B(a[118]), .Z(n8885) );
  NAND U9127 ( .A(n19342), .B(n8885), .Z(n8809) );
  AND U9128 ( .A(n8810), .B(n8809), .Z(n8918) );
  NAND U9129 ( .A(n34), .B(n8811), .Z(n8813) );
  XOR U9130 ( .A(b[7]), .B(a[116]), .Z(n8888) );
  NAND U9131 ( .A(n19486), .B(n8888), .Z(n8812) );
  AND U9132 ( .A(n8813), .B(n8812), .Z(n8916) );
  NAND U9133 ( .A(n31), .B(n8814), .Z(n8816) );
  XOR U9134 ( .A(b[3]), .B(a[120]), .Z(n8891) );
  NAND U9135 ( .A(n32), .B(n8891), .Z(n8815) );
  NAND U9136 ( .A(n8816), .B(n8815), .Z(n8915) );
  XNOR U9137 ( .A(n8916), .B(n8915), .Z(n8917) );
  XOR U9138 ( .A(n8918), .B(n8917), .Z(n8895) );
  XOR U9139 ( .A(n8894), .B(n8895), .Z(n8897) );
  XOR U9140 ( .A(n8896), .B(n8897), .Z(n8868) );
  NANDN U9141 ( .A(n8818), .B(n8817), .Z(n8822) );
  OR U9142 ( .A(n8820), .B(n8819), .Z(n8821) );
  AND U9143 ( .A(n8822), .B(n8821), .Z(n8867) );
  XNOR U9144 ( .A(n8868), .B(n8867), .Z(n8870) );
  NAND U9145 ( .A(n8823), .B(n19724), .Z(n8825) );
  XOR U9146 ( .A(b[11]), .B(a[112]), .Z(n8900) );
  NAND U9147 ( .A(n19692), .B(n8900), .Z(n8824) );
  AND U9148 ( .A(n8825), .B(n8824), .Z(n8911) );
  NAND U9149 ( .A(n19838), .B(n8826), .Z(n8828) );
  XOR U9150 ( .A(b[15]), .B(a[108]), .Z(n8903) );
  NAND U9151 ( .A(n19805), .B(n8903), .Z(n8827) );
  AND U9152 ( .A(n8828), .B(n8827), .Z(n8910) );
  NAND U9153 ( .A(n35), .B(n8829), .Z(n8831) );
  XOR U9154 ( .A(b[9]), .B(a[114]), .Z(n8906) );
  NAND U9155 ( .A(n19598), .B(n8906), .Z(n8830) );
  NAND U9156 ( .A(n8831), .B(n8830), .Z(n8909) );
  XOR U9157 ( .A(n8910), .B(n8909), .Z(n8912) );
  XOR U9158 ( .A(n8911), .B(n8912), .Z(n8922) );
  NANDN U9159 ( .A(n8833), .B(n8832), .Z(n8837) );
  OR U9160 ( .A(n8835), .B(n8834), .Z(n8836) );
  AND U9161 ( .A(n8837), .B(n8836), .Z(n8921) );
  XNOR U9162 ( .A(n8922), .B(n8921), .Z(n8923) );
  NANDN U9163 ( .A(n8839), .B(n8838), .Z(n8843) );
  NANDN U9164 ( .A(n8841), .B(n8840), .Z(n8842) );
  NAND U9165 ( .A(n8843), .B(n8842), .Z(n8924) );
  XNOR U9166 ( .A(n8923), .B(n8924), .Z(n8869) );
  XOR U9167 ( .A(n8870), .B(n8869), .Z(n8928) );
  NANDN U9168 ( .A(n8845), .B(n8844), .Z(n8849) );
  NANDN U9169 ( .A(n8847), .B(n8846), .Z(n8848) );
  AND U9170 ( .A(n8849), .B(n8848), .Z(n8927) );
  XNOR U9171 ( .A(n8928), .B(n8927), .Z(n8929) );
  XOR U9172 ( .A(n8930), .B(n8929), .Z(n8862) );
  NANDN U9173 ( .A(n8851), .B(n8850), .Z(n8855) );
  NAND U9174 ( .A(n8853), .B(n8852), .Z(n8854) );
  AND U9175 ( .A(n8855), .B(n8854), .Z(n8861) );
  XNOR U9176 ( .A(n8862), .B(n8861), .Z(n8863) );
  XNOR U9177 ( .A(n8864), .B(n8863), .Z(n8933) );
  XNOR U9178 ( .A(sreg[362]), .B(n8933), .Z(n8935) );
  NANDN U9179 ( .A(sreg[361]), .B(n8856), .Z(n8860) );
  NAND U9180 ( .A(n8858), .B(n8857), .Z(n8859) );
  NAND U9181 ( .A(n8860), .B(n8859), .Z(n8934) );
  XNOR U9182 ( .A(n8935), .B(n8934), .Z(c[362]) );
  NANDN U9183 ( .A(n8862), .B(n8861), .Z(n8866) );
  NANDN U9184 ( .A(n8864), .B(n8863), .Z(n8865) );
  AND U9185 ( .A(n8866), .B(n8865), .Z(n8941) );
  NANDN U9186 ( .A(n8868), .B(n8867), .Z(n8872) );
  NAND U9187 ( .A(n8870), .B(n8869), .Z(n8871) );
  AND U9188 ( .A(n8872), .B(n8871), .Z(n9007) );
  NANDN U9189 ( .A(n8874), .B(n8873), .Z(n8878) );
  NANDN U9190 ( .A(n8876), .B(n8875), .Z(n8877) );
  AND U9191 ( .A(n8878), .B(n8877), .Z(n8973) );
  NAND U9192 ( .A(b[0]), .B(a[123]), .Z(n8879) );
  XNOR U9193 ( .A(b[1]), .B(n8879), .Z(n8881) );
  NANDN U9194 ( .A(b[0]), .B(a[122]), .Z(n8880) );
  NAND U9195 ( .A(n8881), .B(n8880), .Z(n8953) );
  NAND U9196 ( .A(n19808), .B(n8882), .Z(n8884) );
  XOR U9197 ( .A(b[13]), .B(a[111]), .Z(n8959) );
  NAND U9198 ( .A(n19768), .B(n8959), .Z(n8883) );
  AND U9199 ( .A(n8884), .B(n8883), .Z(n8951) );
  AND U9200 ( .A(b[15]), .B(a[107]), .Z(n8950) );
  XNOR U9201 ( .A(n8951), .B(n8950), .Z(n8952) );
  XNOR U9202 ( .A(n8953), .B(n8952), .Z(n8971) );
  NAND U9203 ( .A(n33), .B(n8885), .Z(n8887) );
  XOR U9204 ( .A(b[5]), .B(a[119]), .Z(n8962) );
  NAND U9205 ( .A(n19342), .B(n8962), .Z(n8886) );
  AND U9206 ( .A(n8887), .B(n8886), .Z(n8995) );
  NAND U9207 ( .A(n34), .B(n8888), .Z(n8890) );
  XOR U9208 ( .A(b[7]), .B(a[117]), .Z(n8965) );
  NAND U9209 ( .A(n19486), .B(n8965), .Z(n8889) );
  AND U9210 ( .A(n8890), .B(n8889), .Z(n8993) );
  NAND U9211 ( .A(n31), .B(n8891), .Z(n8893) );
  XOR U9212 ( .A(b[3]), .B(a[121]), .Z(n8968) );
  NAND U9213 ( .A(n32), .B(n8968), .Z(n8892) );
  NAND U9214 ( .A(n8893), .B(n8892), .Z(n8992) );
  XNOR U9215 ( .A(n8993), .B(n8992), .Z(n8994) );
  XOR U9216 ( .A(n8995), .B(n8994), .Z(n8972) );
  XOR U9217 ( .A(n8971), .B(n8972), .Z(n8974) );
  XOR U9218 ( .A(n8973), .B(n8974), .Z(n8945) );
  NANDN U9219 ( .A(n8895), .B(n8894), .Z(n8899) );
  OR U9220 ( .A(n8897), .B(n8896), .Z(n8898) );
  AND U9221 ( .A(n8899), .B(n8898), .Z(n8944) );
  XNOR U9222 ( .A(n8945), .B(n8944), .Z(n8947) );
  NAND U9223 ( .A(n8900), .B(n19724), .Z(n8902) );
  XOR U9224 ( .A(b[11]), .B(a[113]), .Z(n8977) );
  NAND U9225 ( .A(n19692), .B(n8977), .Z(n8901) );
  AND U9226 ( .A(n8902), .B(n8901), .Z(n8988) );
  NAND U9227 ( .A(n19838), .B(n8903), .Z(n8905) );
  XOR U9228 ( .A(b[15]), .B(a[109]), .Z(n8980) );
  NAND U9229 ( .A(n19805), .B(n8980), .Z(n8904) );
  AND U9230 ( .A(n8905), .B(n8904), .Z(n8987) );
  NAND U9231 ( .A(n35), .B(n8906), .Z(n8908) );
  XOR U9232 ( .A(b[9]), .B(a[115]), .Z(n8983) );
  NAND U9233 ( .A(n19598), .B(n8983), .Z(n8907) );
  NAND U9234 ( .A(n8908), .B(n8907), .Z(n8986) );
  XOR U9235 ( .A(n8987), .B(n8986), .Z(n8989) );
  XOR U9236 ( .A(n8988), .B(n8989), .Z(n8999) );
  NANDN U9237 ( .A(n8910), .B(n8909), .Z(n8914) );
  OR U9238 ( .A(n8912), .B(n8911), .Z(n8913) );
  AND U9239 ( .A(n8914), .B(n8913), .Z(n8998) );
  XNOR U9240 ( .A(n8999), .B(n8998), .Z(n9000) );
  NANDN U9241 ( .A(n8916), .B(n8915), .Z(n8920) );
  NANDN U9242 ( .A(n8918), .B(n8917), .Z(n8919) );
  NAND U9243 ( .A(n8920), .B(n8919), .Z(n9001) );
  XNOR U9244 ( .A(n9000), .B(n9001), .Z(n8946) );
  XOR U9245 ( .A(n8947), .B(n8946), .Z(n9005) );
  NANDN U9246 ( .A(n8922), .B(n8921), .Z(n8926) );
  NANDN U9247 ( .A(n8924), .B(n8923), .Z(n8925) );
  AND U9248 ( .A(n8926), .B(n8925), .Z(n9004) );
  XNOR U9249 ( .A(n9005), .B(n9004), .Z(n9006) );
  XOR U9250 ( .A(n9007), .B(n9006), .Z(n8939) );
  NANDN U9251 ( .A(n8928), .B(n8927), .Z(n8932) );
  NAND U9252 ( .A(n8930), .B(n8929), .Z(n8931) );
  AND U9253 ( .A(n8932), .B(n8931), .Z(n8938) );
  XNOR U9254 ( .A(n8939), .B(n8938), .Z(n8940) );
  XNOR U9255 ( .A(n8941), .B(n8940), .Z(n9010) );
  XNOR U9256 ( .A(sreg[363]), .B(n9010), .Z(n9012) );
  NANDN U9257 ( .A(sreg[362]), .B(n8933), .Z(n8937) );
  NAND U9258 ( .A(n8935), .B(n8934), .Z(n8936) );
  NAND U9259 ( .A(n8937), .B(n8936), .Z(n9011) );
  XNOR U9260 ( .A(n9012), .B(n9011), .Z(c[363]) );
  NANDN U9261 ( .A(n8939), .B(n8938), .Z(n8943) );
  NANDN U9262 ( .A(n8941), .B(n8940), .Z(n8942) );
  AND U9263 ( .A(n8943), .B(n8942), .Z(n9018) );
  NANDN U9264 ( .A(n8945), .B(n8944), .Z(n8949) );
  NAND U9265 ( .A(n8947), .B(n8946), .Z(n8948) );
  AND U9266 ( .A(n8949), .B(n8948), .Z(n9084) );
  NANDN U9267 ( .A(n8951), .B(n8950), .Z(n8955) );
  NANDN U9268 ( .A(n8953), .B(n8952), .Z(n8954) );
  AND U9269 ( .A(n8955), .B(n8954), .Z(n9050) );
  NAND U9270 ( .A(b[0]), .B(a[124]), .Z(n8956) );
  XNOR U9271 ( .A(b[1]), .B(n8956), .Z(n8958) );
  NANDN U9272 ( .A(b[0]), .B(a[123]), .Z(n8957) );
  NAND U9273 ( .A(n8958), .B(n8957), .Z(n9030) );
  NAND U9274 ( .A(n19808), .B(n8959), .Z(n8961) );
  XOR U9275 ( .A(b[13]), .B(a[112]), .Z(n9036) );
  NAND U9276 ( .A(n19768), .B(n9036), .Z(n8960) );
  AND U9277 ( .A(n8961), .B(n8960), .Z(n9028) );
  AND U9278 ( .A(b[15]), .B(a[108]), .Z(n9027) );
  XNOR U9279 ( .A(n9028), .B(n9027), .Z(n9029) );
  XNOR U9280 ( .A(n9030), .B(n9029), .Z(n9048) );
  NAND U9281 ( .A(n33), .B(n8962), .Z(n8964) );
  XOR U9282 ( .A(b[5]), .B(a[120]), .Z(n9039) );
  NAND U9283 ( .A(n19342), .B(n9039), .Z(n8963) );
  AND U9284 ( .A(n8964), .B(n8963), .Z(n9072) );
  NAND U9285 ( .A(n34), .B(n8965), .Z(n8967) );
  XOR U9286 ( .A(b[7]), .B(a[118]), .Z(n9042) );
  NAND U9287 ( .A(n19486), .B(n9042), .Z(n8966) );
  AND U9288 ( .A(n8967), .B(n8966), .Z(n9070) );
  NAND U9289 ( .A(n31), .B(n8968), .Z(n8970) );
  XOR U9290 ( .A(b[3]), .B(a[122]), .Z(n9045) );
  NAND U9291 ( .A(n32), .B(n9045), .Z(n8969) );
  NAND U9292 ( .A(n8970), .B(n8969), .Z(n9069) );
  XNOR U9293 ( .A(n9070), .B(n9069), .Z(n9071) );
  XOR U9294 ( .A(n9072), .B(n9071), .Z(n9049) );
  XOR U9295 ( .A(n9048), .B(n9049), .Z(n9051) );
  XOR U9296 ( .A(n9050), .B(n9051), .Z(n9022) );
  NANDN U9297 ( .A(n8972), .B(n8971), .Z(n8976) );
  OR U9298 ( .A(n8974), .B(n8973), .Z(n8975) );
  AND U9299 ( .A(n8976), .B(n8975), .Z(n9021) );
  XNOR U9300 ( .A(n9022), .B(n9021), .Z(n9024) );
  NAND U9301 ( .A(n8977), .B(n19724), .Z(n8979) );
  XOR U9302 ( .A(b[11]), .B(a[114]), .Z(n9054) );
  NAND U9303 ( .A(n19692), .B(n9054), .Z(n8978) );
  AND U9304 ( .A(n8979), .B(n8978), .Z(n9065) );
  NAND U9305 ( .A(n19838), .B(n8980), .Z(n8982) );
  XOR U9306 ( .A(b[15]), .B(a[110]), .Z(n9057) );
  NAND U9307 ( .A(n19805), .B(n9057), .Z(n8981) );
  AND U9308 ( .A(n8982), .B(n8981), .Z(n9064) );
  NAND U9309 ( .A(n35), .B(n8983), .Z(n8985) );
  XOR U9310 ( .A(b[9]), .B(a[116]), .Z(n9060) );
  NAND U9311 ( .A(n19598), .B(n9060), .Z(n8984) );
  NAND U9312 ( .A(n8985), .B(n8984), .Z(n9063) );
  XOR U9313 ( .A(n9064), .B(n9063), .Z(n9066) );
  XOR U9314 ( .A(n9065), .B(n9066), .Z(n9076) );
  NANDN U9315 ( .A(n8987), .B(n8986), .Z(n8991) );
  OR U9316 ( .A(n8989), .B(n8988), .Z(n8990) );
  AND U9317 ( .A(n8991), .B(n8990), .Z(n9075) );
  XNOR U9318 ( .A(n9076), .B(n9075), .Z(n9077) );
  NANDN U9319 ( .A(n8993), .B(n8992), .Z(n8997) );
  NANDN U9320 ( .A(n8995), .B(n8994), .Z(n8996) );
  NAND U9321 ( .A(n8997), .B(n8996), .Z(n9078) );
  XNOR U9322 ( .A(n9077), .B(n9078), .Z(n9023) );
  XOR U9323 ( .A(n9024), .B(n9023), .Z(n9082) );
  NANDN U9324 ( .A(n8999), .B(n8998), .Z(n9003) );
  NANDN U9325 ( .A(n9001), .B(n9000), .Z(n9002) );
  AND U9326 ( .A(n9003), .B(n9002), .Z(n9081) );
  XNOR U9327 ( .A(n9082), .B(n9081), .Z(n9083) );
  XOR U9328 ( .A(n9084), .B(n9083), .Z(n9016) );
  NANDN U9329 ( .A(n9005), .B(n9004), .Z(n9009) );
  NAND U9330 ( .A(n9007), .B(n9006), .Z(n9008) );
  AND U9331 ( .A(n9009), .B(n9008), .Z(n9015) );
  XNOR U9332 ( .A(n9016), .B(n9015), .Z(n9017) );
  XNOR U9333 ( .A(n9018), .B(n9017), .Z(n9087) );
  XNOR U9334 ( .A(sreg[364]), .B(n9087), .Z(n9089) );
  NANDN U9335 ( .A(sreg[363]), .B(n9010), .Z(n9014) );
  NAND U9336 ( .A(n9012), .B(n9011), .Z(n9013) );
  NAND U9337 ( .A(n9014), .B(n9013), .Z(n9088) );
  XNOR U9338 ( .A(n9089), .B(n9088), .Z(c[364]) );
  NANDN U9339 ( .A(n9016), .B(n9015), .Z(n9020) );
  NANDN U9340 ( .A(n9018), .B(n9017), .Z(n9019) );
  AND U9341 ( .A(n9020), .B(n9019), .Z(n9095) );
  NANDN U9342 ( .A(n9022), .B(n9021), .Z(n9026) );
  NAND U9343 ( .A(n9024), .B(n9023), .Z(n9025) );
  AND U9344 ( .A(n9026), .B(n9025), .Z(n9161) );
  NANDN U9345 ( .A(n9028), .B(n9027), .Z(n9032) );
  NANDN U9346 ( .A(n9030), .B(n9029), .Z(n9031) );
  AND U9347 ( .A(n9032), .B(n9031), .Z(n9127) );
  NAND U9348 ( .A(b[0]), .B(a[125]), .Z(n9033) );
  XNOR U9349 ( .A(b[1]), .B(n9033), .Z(n9035) );
  NANDN U9350 ( .A(b[0]), .B(a[124]), .Z(n9034) );
  NAND U9351 ( .A(n9035), .B(n9034), .Z(n9107) );
  NAND U9352 ( .A(n19808), .B(n9036), .Z(n9038) );
  XOR U9353 ( .A(b[13]), .B(a[113]), .Z(n9110) );
  NAND U9354 ( .A(n19768), .B(n9110), .Z(n9037) );
  AND U9355 ( .A(n9038), .B(n9037), .Z(n9105) );
  AND U9356 ( .A(b[15]), .B(a[109]), .Z(n9104) );
  XNOR U9357 ( .A(n9105), .B(n9104), .Z(n9106) );
  XNOR U9358 ( .A(n9107), .B(n9106), .Z(n9125) );
  NAND U9359 ( .A(n33), .B(n9039), .Z(n9041) );
  XOR U9360 ( .A(b[5]), .B(a[121]), .Z(n9116) );
  NAND U9361 ( .A(n19342), .B(n9116), .Z(n9040) );
  AND U9362 ( .A(n9041), .B(n9040), .Z(n9149) );
  NAND U9363 ( .A(n34), .B(n9042), .Z(n9044) );
  XOR U9364 ( .A(b[7]), .B(a[119]), .Z(n9119) );
  NAND U9365 ( .A(n19486), .B(n9119), .Z(n9043) );
  AND U9366 ( .A(n9044), .B(n9043), .Z(n9147) );
  NAND U9367 ( .A(n31), .B(n9045), .Z(n9047) );
  XOR U9368 ( .A(b[3]), .B(a[123]), .Z(n9122) );
  NAND U9369 ( .A(n32), .B(n9122), .Z(n9046) );
  NAND U9370 ( .A(n9047), .B(n9046), .Z(n9146) );
  XNOR U9371 ( .A(n9147), .B(n9146), .Z(n9148) );
  XOR U9372 ( .A(n9149), .B(n9148), .Z(n9126) );
  XOR U9373 ( .A(n9125), .B(n9126), .Z(n9128) );
  XOR U9374 ( .A(n9127), .B(n9128), .Z(n9099) );
  NANDN U9375 ( .A(n9049), .B(n9048), .Z(n9053) );
  OR U9376 ( .A(n9051), .B(n9050), .Z(n9052) );
  AND U9377 ( .A(n9053), .B(n9052), .Z(n9098) );
  XNOR U9378 ( .A(n9099), .B(n9098), .Z(n9101) );
  NAND U9379 ( .A(n9054), .B(n19724), .Z(n9056) );
  XOR U9380 ( .A(b[11]), .B(a[115]), .Z(n9131) );
  NAND U9381 ( .A(n19692), .B(n9131), .Z(n9055) );
  AND U9382 ( .A(n9056), .B(n9055), .Z(n9142) );
  NAND U9383 ( .A(n19838), .B(n9057), .Z(n9059) );
  XOR U9384 ( .A(b[15]), .B(a[111]), .Z(n9134) );
  NAND U9385 ( .A(n19805), .B(n9134), .Z(n9058) );
  AND U9386 ( .A(n9059), .B(n9058), .Z(n9141) );
  NAND U9387 ( .A(n35), .B(n9060), .Z(n9062) );
  XOR U9388 ( .A(b[9]), .B(a[117]), .Z(n9137) );
  NAND U9389 ( .A(n19598), .B(n9137), .Z(n9061) );
  NAND U9390 ( .A(n9062), .B(n9061), .Z(n9140) );
  XOR U9391 ( .A(n9141), .B(n9140), .Z(n9143) );
  XOR U9392 ( .A(n9142), .B(n9143), .Z(n9153) );
  NANDN U9393 ( .A(n9064), .B(n9063), .Z(n9068) );
  OR U9394 ( .A(n9066), .B(n9065), .Z(n9067) );
  AND U9395 ( .A(n9068), .B(n9067), .Z(n9152) );
  XNOR U9396 ( .A(n9153), .B(n9152), .Z(n9154) );
  NANDN U9397 ( .A(n9070), .B(n9069), .Z(n9074) );
  NANDN U9398 ( .A(n9072), .B(n9071), .Z(n9073) );
  NAND U9399 ( .A(n9074), .B(n9073), .Z(n9155) );
  XNOR U9400 ( .A(n9154), .B(n9155), .Z(n9100) );
  XOR U9401 ( .A(n9101), .B(n9100), .Z(n9159) );
  NANDN U9402 ( .A(n9076), .B(n9075), .Z(n9080) );
  NANDN U9403 ( .A(n9078), .B(n9077), .Z(n9079) );
  AND U9404 ( .A(n9080), .B(n9079), .Z(n9158) );
  XNOR U9405 ( .A(n9159), .B(n9158), .Z(n9160) );
  XOR U9406 ( .A(n9161), .B(n9160), .Z(n9093) );
  NANDN U9407 ( .A(n9082), .B(n9081), .Z(n9086) );
  NAND U9408 ( .A(n9084), .B(n9083), .Z(n9085) );
  AND U9409 ( .A(n9086), .B(n9085), .Z(n9092) );
  XNOR U9410 ( .A(n9093), .B(n9092), .Z(n9094) );
  XNOR U9411 ( .A(n9095), .B(n9094), .Z(n9164) );
  XNOR U9412 ( .A(sreg[365]), .B(n9164), .Z(n9166) );
  NANDN U9413 ( .A(sreg[364]), .B(n9087), .Z(n9091) );
  NAND U9414 ( .A(n9089), .B(n9088), .Z(n9090) );
  NAND U9415 ( .A(n9091), .B(n9090), .Z(n9165) );
  XNOR U9416 ( .A(n9166), .B(n9165), .Z(c[365]) );
  NANDN U9417 ( .A(n9093), .B(n9092), .Z(n9097) );
  NANDN U9418 ( .A(n9095), .B(n9094), .Z(n9096) );
  AND U9419 ( .A(n9097), .B(n9096), .Z(n9172) );
  NANDN U9420 ( .A(n9099), .B(n9098), .Z(n9103) );
  NAND U9421 ( .A(n9101), .B(n9100), .Z(n9102) );
  AND U9422 ( .A(n9103), .B(n9102), .Z(n9238) );
  NANDN U9423 ( .A(n9105), .B(n9104), .Z(n9109) );
  NANDN U9424 ( .A(n9107), .B(n9106), .Z(n9108) );
  AND U9425 ( .A(n9109), .B(n9108), .Z(n9225) );
  NAND U9426 ( .A(n19808), .B(n9110), .Z(n9112) );
  XOR U9427 ( .A(b[13]), .B(a[114]), .Z(n9211) );
  NAND U9428 ( .A(n19768), .B(n9211), .Z(n9111) );
  AND U9429 ( .A(n9112), .B(n9111), .Z(n9203) );
  AND U9430 ( .A(b[15]), .B(a[110]), .Z(n9202) );
  XNOR U9431 ( .A(n9203), .B(n9202), .Z(n9204) );
  NAND U9432 ( .A(b[0]), .B(a[126]), .Z(n9113) );
  XNOR U9433 ( .A(b[1]), .B(n9113), .Z(n9115) );
  NANDN U9434 ( .A(b[0]), .B(a[125]), .Z(n9114) );
  NAND U9435 ( .A(n9115), .B(n9114), .Z(n9205) );
  XNOR U9436 ( .A(n9204), .B(n9205), .Z(n9223) );
  NAND U9437 ( .A(n33), .B(n9116), .Z(n9118) );
  XOR U9438 ( .A(b[5]), .B(a[122]), .Z(n9214) );
  NAND U9439 ( .A(n19342), .B(n9214), .Z(n9117) );
  AND U9440 ( .A(n9118), .B(n9117), .Z(n9199) );
  NAND U9441 ( .A(n34), .B(n9119), .Z(n9121) );
  XOR U9442 ( .A(b[7]), .B(a[120]), .Z(n9217) );
  NAND U9443 ( .A(n19486), .B(n9217), .Z(n9120) );
  AND U9444 ( .A(n9121), .B(n9120), .Z(n9197) );
  NAND U9445 ( .A(n31), .B(n9122), .Z(n9124) );
  XOR U9446 ( .A(b[3]), .B(a[124]), .Z(n9220) );
  NAND U9447 ( .A(n32), .B(n9220), .Z(n9123) );
  NAND U9448 ( .A(n9124), .B(n9123), .Z(n9196) );
  XNOR U9449 ( .A(n9197), .B(n9196), .Z(n9198) );
  XOR U9450 ( .A(n9199), .B(n9198), .Z(n9224) );
  XOR U9451 ( .A(n9223), .B(n9224), .Z(n9226) );
  XOR U9452 ( .A(n9225), .B(n9226), .Z(n9176) );
  NANDN U9453 ( .A(n9126), .B(n9125), .Z(n9130) );
  OR U9454 ( .A(n9128), .B(n9127), .Z(n9129) );
  AND U9455 ( .A(n9130), .B(n9129), .Z(n9175) );
  XNOR U9456 ( .A(n9176), .B(n9175), .Z(n9178) );
  NAND U9457 ( .A(n9131), .B(n19724), .Z(n9133) );
  XOR U9458 ( .A(b[11]), .B(a[116]), .Z(n9181) );
  NAND U9459 ( .A(n19692), .B(n9181), .Z(n9132) );
  AND U9460 ( .A(n9133), .B(n9132), .Z(n9192) );
  NAND U9461 ( .A(n19838), .B(n9134), .Z(n9136) );
  XOR U9462 ( .A(b[15]), .B(a[112]), .Z(n9184) );
  NAND U9463 ( .A(n19805), .B(n9184), .Z(n9135) );
  AND U9464 ( .A(n9136), .B(n9135), .Z(n9191) );
  NAND U9465 ( .A(n35), .B(n9137), .Z(n9139) );
  XOR U9466 ( .A(b[9]), .B(a[118]), .Z(n9187) );
  NAND U9467 ( .A(n19598), .B(n9187), .Z(n9138) );
  NAND U9468 ( .A(n9139), .B(n9138), .Z(n9190) );
  XOR U9469 ( .A(n9191), .B(n9190), .Z(n9193) );
  XOR U9470 ( .A(n9192), .B(n9193), .Z(n9230) );
  NANDN U9471 ( .A(n9141), .B(n9140), .Z(n9145) );
  OR U9472 ( .A(n9143), .B(n9142), .Z(n9144) );
  AND U9473 ( .A(n9145), .B(n9144), .Z(n9229) );
  XNOR U9474 ( .A(n9230), .B(n9229), .Z(n9231) );
  NANDN U9475 ( .A(n9147), .B(n9146), .Z(n9151) );
  NANDN U9476 ( .A(n9149), .B(n9148), .Z(n9150) );
  NAND U9477 ( .A(n9151), .B(n9150), .Z(n9232) );
  XNOR U9478 ( .A(n9231), .B(n9232), .Z(n9177) );
  XOR U9479 ( .A(n9178), .B(n9177), .Z(n9236) );
  NANDN U9480 ( .A(n9153), .B(n9152), .Z(n9157) );
  NANDN U9481 ( .A(n9155), .B(n9154), .Z(n9156) );
  AND U9482 ( .A(n9157), .B(n9156), .Z(n9235) );
  XNOR U9483 ( .A(n9236), .B(n9235), .Z(n9237) );
  XOR U9484 ( .A(n9238), .B(n9237), .Z(n9170) );
  NANDN U9485 ( .A(n9159), .B(n9158), .Z(n9163) );
  NAND U9486 ( .A(n9161), .B(n9160), .Z(n9162) );
  AND U9487 ( .A(n9163), .B(n9162), .Z(n9169) );
  XNOR U9488 ( .A(n9170), .B(n9169), .Z(n9171) );
  XNOR U9489 ( .A(n9172), .B(n9171), .Z(n9241) );
  XNOR U9490 ( .A(sreg[366]), .B(n9241), .Z(n9243) );
  NANDN U9491 ( .A(sreg[365]), .B(n9164), .Z(n9168) );
  NAND U9492 ( .A(n9166), .B(n9165), .Z(n9167) );
  NAND U9493 ( .A(n9168), .B(n9167), .Z(n9242) );
  XNOR U9494 ( .A(n9243), .B(n9242), .Z(c[366]) );
  NANDN U9495 ( .A(n9170), .B(n9169), .Z(n9174) );
  NANDN U9496 ( .A(n9172), .B(n9171), .Z(n9173) );
  AND U9497 ( .A(n9174), .B(n9173), .Z(n9249) );
  NANDN U9498 ( .A(n9176), .B(n9175), .Z(n9180) );
  NAND U9499 ( .A(n9178), .B(n9177), .Z(n9179) );
  AND U9500 ( .A(n9180), .B(n9179), .Z(n9315) );
  NAND U9501 ( .A(n9181), .B(n19724), .Z(n9183) );
  XOR U9502 ( .A(b[11]), .B(a[117]), .Z(n9285) );
  NAND U9503 ( .A(n19692), .B(n9285), .Z(n9182) );
  AND U9504 ( .A(n9183), .B(n9182), .Z(n9296) );
  NAND U9505 ( .A(n19838), .B(n9184), .Z(n9186) );
  XOR U9506 ( .A(b[15]), .B(a[113]), .Z(n9288) );
  NAND U9507 ( .A(n19805), .B(n9288), .Z(n9185) );
  AND U9508 ( .A(n9186), .B(n9185), .Z(n9295) );
  NAND U9509 ( .A(n35), .B(n9187), .Z(n9189) );
  XOR U9510 ( .A(b[9]), .B(a[119]), .Z(n9291) );
  NAND U9511 ( .A(n19598), .B(n9291), .Z(n9188) );
  NAND U9512 ( .A(n9189), .B(n9188), .Z(n9294) );
  XOR U9513 ( .A(n9295), .B(n9294), .Z(n9297) );
  XOR U9514 ( .A(n9296), .B(n9297), .Z(n9307) );
  NANDN U9515 ( .A(n9191), .B(n9190), .Z(n9195) );
  OR U9516 ( .A(n9193), .B(n9192), .Z(n9194) );
  AND U9517 ( .A(n9195), .B(n9194), .Z(n9306) );
  XNOR U9518 ( .A(n9307), .B(n9306), .Z(n9308) );
  NANDN U9519 ( .A(n9197), .B(n9196), .Z(n9201) );
  NANDN U9520 ( .A(n9199), .B(n9198), .Z(n9200) );
  NAND U9521 ( .A(n9201), .B(n9200), .Z(n9309) );
  XNOR U9522 ( .A(n9308), .B(n9309), .Z(n9255) );
  NANDN U9523 ( .A(n9203), .B(n9202), .Z(n9207) );
  NANDN U9524 ( .A(n9205), .B(n9204), .Z(n9206) );
  AND U9525 ( .A(n9207), .B(n9206), .Z(n9281) );
  NAND U9526 ( .A(b[0]), .B(a[127]), .Z(n9208) );
  XNOR U9527 ( .A(b[1]), .B(n9208), .Z(n9210) );
  NANDN U9528 ( .A(b[0]), .B(a[126]), .Z(n9209) );
  NAND U9529 ( .A(n9210), .B(n9209), .Z(n9261) );
  NAND U9530 ( .A(n19808), .B(n9211), .Z(n9213) );
  XOR U9531 ( .A(b[13]), .B(a[115]), .Z(n9264) );
  NAND U9532 ( .A(n19768), .B(n9264), .Z(n9212) );
  AND U9533 ( .A(n9213), .B(n9212), .Z(n9259) );
  AND U9534 ( .A(b[15]), .B(a[111]), .Z(n9258) );
  XNOR U9535 ( .A(n9259), .B(n9258), .Z(n9260) );
  XNOR U9536 ( .A(n9261), .B(n9260), .Z(n9279) );
  NAND U9537 ( .A(n33), .B(n9214), .Z(n9216) );
  XOR U9538 ( .A(b[5]), .B(a[123]), .Z(n9270) );
  NAND U9539 ( .A(n19342), .B(n9270), .Z(n9215) );
  AND U9540 ( .A(n9216), .B(n9215), .Z(n9303) );
  NAND U9541 ( .A(n34), .B(n9217), .Z(n9219) );
  XOR U9542 ( .A(b[7]), .B(a[121]), .Z(n9273) );
  NAND U9543 ( .A(n19486), .B(n9273), .Z(n9218) );
  AND U9544 ( .A(n9219), .B(n9218), .Z(n9301) );
  NAND U9545 ( .A(n31), .B(n9220), .Z(n9222) );
  XOR U9546 ( .A(b[3]), .B(a[125]), .Z(n9276) );
  NAND U9547 ( .A(n32), .B(n9276), .Z(n9221) );
  NAND U9548 ( .A(n9222), .B(n9221), .Z(n9300) );
  XNOR U9549 ( .A(n9301), .B(n9300), .Z(n9302) );
  XOR U9550 ( .A(n9303), .B(n9302), .Z(n9280) );
  XOR U9551 ( .A(n9279), .B(n9280), .Z(n9282) );
  XOR U9552 ( .A(n9281), .B(n9282), .Z(n9253) );
  NANDN U9553 ( .A(n9224), .B(n9223), .Z(n9228) );
  OR U9554 ( .A(n9226), .B(n9225), .Z(n9227) );
  AND U9555 ( .A(n9228), .B(n9227), .Z(n9252) );
  XNOR U9556 ( .A(n9253), .B(n9252), .Z(n9254) );
  XOR U9557 ( .A(n9255), .B(n9254), .Z(n9313) );
  NANDN U9558 ( .A(n9230), .B(n9229), .Z(n9234) );
  NANDN U9559 ( .A(n9232), .B(n9231), .Z(n9233) );
  AND U9560 ( .A(n9234), .B(n9233), .Z(n9312) );
  XNOR U9561 ( .A(n9313), .B(n9312), .Z(n9314) );
  XOR U9562 ( .A(n9315), .B(n9314), .Z(n9247) );
  NANDN U9563 ( .A(n9236), .B(n9235), .Z(n9240) );
  NAND U9564 ( .A(n9238), .B(n9237), .Z(n9239) );
  AND U9565 ( .A(n9240), .B(n9239), .Z(n9246) );
  XNOR U9566 ( .A(n9247), .B(n9246), .Z(n9248) );
  XNOR U9567 ( .A(n9249), .B(n9248), .Z(n9318) );
  XNOR U9568 ( .A(sreg[367]), .B(n9318), .Z(n9320) );
  NANDN U9569 ( .A(sreg[366]), .B(n9241), .Z(n9245) );
  NAND U9570 ( .A(n9243), .B(n9242), .Z(n9244) );
  NAND U9571 ( .A(n9245), .B(n9244), .Z(n9319) );
  XNOR U9572 ( .A(n9320), .B(n9319), .Z(c[367]) );
  NANDN U9573 ( .A(n9247), .B(n9246), .Z(n9251) );
  NANDN U9574 ( .A(n9249), .B(n9248), .Z(n9250) );
  AND U9575 ( .A(n9251), .B(n9250), .Z(n9326) );
  NANDN U9576 ( .A(n9253), .B(n9252), .Z(n9257) );
  NAND U9577 ( .A(n9255), .B(n9254), .Z(n9256) );
  AND U9578 ( .A(n9257), .B(n9256), .Z(n9392) );
  NANDN U9579 ( .A(n9259), .B(n9258), .Z(n9263) );
  NANDN U9580 ( .A(n9261), .B(n9260), .Z(n9262) );
  AND U9581 ( .A(n9263), .B(n9262), .Z(n9358) );
  NAND U9582 ( .A(n19808), .B(n9264), .Z(n9266) );
  XOR U9583 ( .A(b[13]), .B(a[116]), .Z(n9344) );
  NAND U9584 ( .A(n19768), .B(n9344), .Z(n9265) );
  AND U9585 ( .A(n9266), .B(n9265), .Z(n9336) );
  AND U9586 ( .A(b[15]), .B(a[112]), .Z(n9335) );
  XNOR U9587 ( .A(n9336), .B(n9335), .Z(n9337) );
  NAND U9588 ( .A(b[0]), .B(a[128]), .Z(n9267) );
  XNOR U9589 ( .A(b[1]), .B(n9267), .Z(n9269) );
  NANDN U9590 ( .A(b[0]), .B(a[127]), .Z(n9268) );
  NAND U9591 ( .A(n9269), .B(n9268), .Z(n9338) );
  XNOR U9592 ( .A(n9337), .B(n9338), .Z(n9356) );
  NAND U9593 ( .A(n33), .B(n9270), .Z(n9272) );
  XOR U9594 ( .A(b[5]), .B(a[124]), .Z(n9347) );
  NAND U9595 ( .A(n19342), .B(n9347), .Z(n9271) );
  AND U9596 ( .A(n9272), .B(n9271), .Z(n9380) );
  NAND U9597 ( .A(n34), .B(n9273), .Z(n9275) );
  XOR U9598 ( .A(b[7]), .B(a[122]), .Z(n9350) );
  NAND U9599 ( .A(n19486), .B(n9350), .Z(n9274) );
  AND U9600 ( .A(n9275), .B(n9274), .Z(n9378) );
  NAND U9601 ( .A(n31), .B(n9276), .Z(n9278) );
  XOR U9602 ( .A(b[3]), .B(a[126]), .Z(n9353) );
  NAND U9603 ( .A(n32), .B(n9353), .Z(n9277) );
  NAND U9604 ( .A(n9278), .B(n9277), .Z(n9377) );
  XNOR U9605 ( .A(n9378), .B(n9377), .Z(n9379) );
  XOR U9606 ( .A(n9380), .B(n9379), .Z(n9357) );
  XOR U9607 ( .A(n9356), .B(n9357), .Z(n9359) );
  XOR U9608 ( .A(n9358), .B(n9359), .Z(n9330) );
  NANDN U9609 ( .A(n9280), .B(n9279), .Z(n9284) );
  OR U9610 ( .A(n9282), .B(n9281), .Z(n9283) );
  AND U9611 ( .A(n9284), .B(n9283), .Z(n9329) );
  XNOR U9612 ( .A(n9330), .B(n9329), .Z(n9332) );
  NAND U9613 ( .A(n9285), .B(n19724), .Z(n9287) );
  XOR U9614 ( .A(b[11]), .B(a[118]), .Z(n9362) );
  NAND U9615 ( .A(n19692), .B(n9362), .Z(n9286) );
  AND U9616 ( .A(n9287), .B(n9286), .Z(n9373) );
  NAND U9617 ( .A(n19838), .B(n9288), .Z(n9290) );
  XOR U9618 ( .A(b[15]), .B(a[114]), .Z(n9365) );
  NAND U9619 ( .A(n19805), .B(n9365), .Z(n9289) );
  AND U9620 ( .A(n9290), .B(n9289), .Z(n9372) );
  NAND U9621 ( .A(n35), .B(n9291), .Z(n9293) );
  XOR U9622 ( .A(b[9]), .B(a[120]), .Z(n9368) );
  NAND U9623 ( .A(n19598), .B(n9368), .Z(n9292) );
  NAND U9624 ( .A(n9293), .B(n9292), .Z(n9371) );
  XOR U9625 ( .A(n9372), .B(n9371), .Z(n9374) );
  XOR U9626 ( .A(n9373), .B(n9374), .Z(n9384) );
  NANDN U9627 ( .A(n9295), .B(n9294), .Z(n9299) );
  OR U9628 ( .A(n9297), .B(n9296), .Z(n9298) );
  AND U9629 ( .A(n9299), .B(n9298), .Z(n9383) );
  XNOR U9630 ( .A(n9384), .B(n9383), .Z(n9385) );
  NANDN U9631 ( .A(n9301), .B(n9300), .Z(n9305) );
  NANDN U9632 ( .A(n9303), .B(n9302), .Z(n9304) );
  NAND U9633 ( .A(n9305), .B(n9304), .Z(n9386) );
  XNOR U9634 ( .A(n9385), .B(n9386), .Z(n9331) );
  XOR U9635 ( .A(n9332), .B(n9331), .Z(n9390) );
  NANDN U9636 ( .A(n9307), .B(n9306), .Z(n9311) );
  NANDN U9637 ( .A(n9309), .B(n9308), .Z(n9310) );
  AND U9638 ( .A(n9311), .B(n9310), .Z(n9389) );
  XNOR U9639 ( .A(n9390), .B(n9389), .Z(n9391) );
  XOR U9640 ( .A(n9392), .B(n9391), .Z(n9324) );
  NANDN U9641 ( .A(n9313), .B(n9312), .Z(n9317) );
  NAND U9642 ( .A(n9315), .B(n9314), .Z(n9316) );
  AND U9643 ( .A(n9317), .B(n9316), .Z(n9323) );
  XNOR U9644 ( .A(n9324), .B(n9323), .Z(n9325) );
  XNOR U9645 ( .A(n9326), .B(n9325), .Z(n9395) );
  XNOR U9646 ( .A(sreg[368]), .B(n9395), .Z(n9397) );
  NANDN U9647 ( .A(sreg[367]), .B(n9318), .Z(n9322) );
  NAND U9648 ( .A(n9320), .B(n9319), .Z(n9321) );
  NAND U9649 ( .A(n9322), .B(n9321), .Z(n9396) );
  XNOR U9650 ( .A(n9397), .B(n9396), .Z(c[368]) );
  NANDN U9651 ( .A(n9324), .B(n9323), .Z(n9328) );
  NANDN U9652 ( .A(n9326), .B(n9325), .Z(n9327) );
  AND U9653 ( .A(n9328), .B(n9327), .Z(n9403) );
  NANDN U9654 ( .A(n9330), .B(n9329), .Z(n9334) );
  NAND U9655 ( .A(n9332), .B(n9331), .Z(n9333) );
  AND U9656 ( .A(n9334), .B(n9333), .Z(n9469) );
  NANDN U9657 ( .A(n9336), .B(n9335), .Z(n9340) );
  NANDN U9658 ( .A(n9338), .B(n9337), .Z(n9339) );
  AND U9659 ( .A(n9340), .B(n9339), .Z(n9456) );
  NAND U9660 ( .A(b[0]), .B(a[129]), .Z(n9341) );
  XNOR U9661 ( .A(b[1]), .B(n9341), .Z(n9343) );
  NANDN U9662 ( .A(b[0]), .B(a[128]), .Z(n9342) );
  NAND U9663 ( .A(n9343), .B(n9342), .Z(n9436) );
  NAND U9664 ( .A(n19808), .B(n9344), .Z(n9346) );
  XOR U9665 ( .A(b[13]), .B(a[117]), .Z(n9442) );
  NAND U9666 ( .A(n19768), .B(n9442), .Z(n9345) );
  AND U9667 ( .A(n9346), .B(n9345), .Z(n9434) );
  AND U9668 ( .A(b[15]), .B(a[113]), .Z(n9433) );
  XNOR U9669 ( .A(n9434), .B(n9433), .Z(n9435) );
  XNOR U9670 ( .A(n9436), .B(n9435), .Z(n9454) );
  NAND U9671 ( .A(n33), .B(n9347), .Z(n9349) );
  XOR U9672 ( .A(b[5]), .B(a[125]), .Z(n9445) );
  NAND U9673 ( .A(n19342), .B(n9445), .Z(n9348) );
  AND U9674 ( .A(n9349), .B(n9348), .Z(n9430) );
  NAND U9675 ( .A(n34), .B(n9350), .Z(n9352) );
  XOR U9676 ( .A(b[7]), .B(a[123]), .Z(n9448) );
  NAND U9677 ( .A(n19486), .B(n9448), .Z(n9351) );
  AND U9678 ( .A(n9352), .B(n9351), .Z(n9428) );
  NAND U9679 ( .A(n31), .B(n9353), .Z(n9355) );
  XOR U9680 ( .A(b[3]), .B(a[127]), .Z(n9451) );
  NAND U9681 ( .A(n32), .B(n9451), .Z(n9354) );
  NAND U9682 ( .A(n9355), .B(n9354), .Z(n9427) );
  XNOR U9683 ( .A(n9428), .B(n9427), .Z(n9429) );
  XOR U9684 ( .A(n9430), .B(n9429), .Z(n9455) );
  XOR U9685 ( .A(n9454), .B(n9455), .Z(n9457) );
  XOR U9686 ( .A(n9456), .B(n9457), .Z(n9407) );
  NANDN U9687 ( .A(n9357), .B(n9356), .Z(n9361) );
  OR U9688 ( .A(n9359), .B(n9358), .Z(n9360) );
  AND U9689 ( .A(n9361), .B(n9360), .Z(n9406) );
  XNOR U9690 ( .A(n9407), .B(n9406), .Z(n9409) );
  NAND U9691 ( .A(n9362), .B(n19724), .Z(n9364) );
  XOR U9692 ( .A(b[11]), .B(a[119]), .Z(n9412) );
  NAND U9693 ( .A(n19692), .B(n9412), .Z(n9363) );
  AND U9694 ( .A(n9364), .B(n9363), .Z(n9423) );
  NAND U9695 ( .A(n19838), .B(n9365), .Z(n9367) );
  XOR U9696 ( .A(b[15]), .B(a[115]), .Z(n9415) );
  NAND U9697 ( .A(n19805), .B(n9415), .Z(n9366) );
  AND U9698 ( .A(n9367), .B(n9366), .Z(n9422) );
  NAND U9699 ( .A(n35), .B(n9368), .Z(n9370) );
  XOR U9700 ( .A(b[9]), .B(a[121]), .Z(n9418) );
  NAND U9701 ( .A(n19598), .B(n9418), .Z(n9369) );
  NAND U9702 ( .A(n9370), .B(n9369), .Z(n9421) );
  XOR U9703 ( .A(n9422), .B(n9421), .Z(n9424) );
  XOR U9704 ( .A(n9423), .B(n9424), .Z(n9461) );
  NANDN U9705 ( .A(n9372), .B(n9371), .Z(n9376) );
  OR U9706 ( .A(n9374), .B(n9373), .Z(n9375) );
  AND U9707 ( .A(n9376), .B(n9375), .Z(n9460) );
  XNOR U9708 ( .A(n9461), .B(n9460), .Z(n9462) );
  NANDN U9709 ( .A(n9378), .B(n9377), .Z(n9382) );
  NANDN U9710 ( .A(n9380), .B(n9379), .Z(n9381) );
  NAND U9711 ( .A(n9382), .B(n9381), .Z(n9463) );
  XNOR U9712 ( .A(n9462), .B(n9463), .Z(n9408) );
  XOR U9713 ( .A(n9409), .B(n9408), .Z(n9467) );
  NANDN U9714 ( .A(n9384), .B(n9383), .Z(n9388) );
  NANDN U9715 ( .A(n9386), .B(n9385), .Z(n9387) );
  AND U9716 ( .A(n9388), .B(n9387), .Z(n9466) );
  XNOR U9717 ( .A(n9467), .B(n9466), .Z(n9468) );
  XOR U9718 ( .A(n9469), .B(n9468), .Z(n9401) );
  NANDN U9719 ( .A(n9390), .B(n9389), .Z(n9394) );
  NAND U9720 ( .A(n9392), .B(n9391), .Z(n9393) );
  AND U9721 ( .A(n9394), .B(n9393), .Z(n9400) );
  XNOR U9722 ( .A(n9401), .B(n9400), .Z(n9402) );
  XNOR U9723 ( .A(n9403), .B(n9402), .Z(n9472) );
  XNOR U9724 ( .A(sreg[369]), .B(n9472), .Z(n9474) );
  NANDN U9725 ( .A(sreg[368]), .B(n9395), .Z(n9399) );
  NAND U9726 ( .A(n9397), .B(n9396), .Z(n9398) );
  NAND U9727 ( .A(n9399), .B(n9398), .Z(n9473) );
  XNOR U9728 ( .A(n9474), .B(n9473), .Z(c[369]) );
  NANDN U9729 ( .A(n9401), .B(n9400), .Z(n9405) );
  NANDN U9730 ( .A(n9403), .B(n9402), .Z(n9404) );
  AND U9731 ( .A(n9405), .B(n9404), .Z(n9480) );
  NANDN U9732 ( .A(n9407), .B(n9406), .Z(n9411) );
  NAND U9733 ( .A(n9409), .B(n9408), .Z(n9410) );
  AND U9734 ( .A(n9411), .B(n9410), .Z(n9546) );
  NAND U9735 ( .A(n9412), .B(n19724), .Z(n9414) );
  XOR U9736 ( .A(b[11]), .B(a[120]), .Z(n9489) );
  NAND U9737 ( .A(n19692), .B(n9489), .Z(n9413) );
  AND U9738 ( .A(n9414), .B(n9413), .Z(n9500) );
  NAND U9739 ( .A(n19838), .B(n9415), .Z(n9417) );
  XOR U9740 ( .A(b[15]), .B(a[116]), .Z(n9492) );
  NAND U9741 ( .A(n19805), .B(n9492), .Z(n9416) );
  AND U9742 ( .A(n9417), .B(n9416), .Z(n9499) );
  NAND U9743 ( .A(n35), .B(n9418), .Z(n9420) );
  XOR U9744 ( .A(b[9]), .B(a[122]), .Z(n9495) );
  NAND U9745 ( .A(n19598), .B(n9495), .Z(n9419) );
  NAND U9746 ( .A(n9420), .B(n9419), .Z(n9498) );
  XOR U9747 ( .A(n9499), .B(n9498), .Z(n9501) );
  XOR U9748 ( .A(n9500), .B(n9501), .Z(n9538) );
  NANDN U9749 ( .A(n9422), .B(n9421), .Z(n9426) );
  OR U9750 ( .A(n9424), .B(n9423), .Z(n9425) );
  AND U9751 ( .A(n9426), .B(n9425), .Z(n9537) );
  XNOR U9752 ( .A(n9538), .B(n9537), .Z(n9539) );
  NANDN U9753 ( .A(n9428), .B(n9427), .Z(n9432) );
  NANDN U9754 ( .A(n9430), .B(n9429), .Z(n9431) );
  NAND U9755 ( .A(n9432), .B(n9431), .Z(n9540) );
  XNOR U9756 ( .A(n9539), .B(n9540), .Z(n9486) );
  NANDN U9757 ( .A(n9434), .B(n9433), .Z(n9438) );
  NANDN U9758 ( .A(n9436), .B(n9435), .Z(n9437) );
  AND U9759 ( .A(n9438), .B(n9437), .Z(n9533) );
  NAND U9760 ( .A(b[0]), .B(a[130]), .Z(n9439) );
  XNOR U9761 ( .A(b[1]), .B(n9439), .Z(n9441) );
  NANDN U9762 ( .A(b[0]), .B(a[129]), .Z(n9440) );
  NAND U9763 ( .A(n9441), .B(n9440), .Z(n9513) );
  NAND U9764 ( .A(n19808), .B(n9442), .Z(n9444) );
  XOR U9765 ( .A(b[13]), .B(a[118]), .Z(n9516) );
  NAND U9766 ( .A(n19768), .B(n9516), .Z(n9443) );
  AND U9767 ( .A(n9444), .B(n9443), .Z(n9511) );
  AND U9768 ( .A(b[15]), .B(a[114]), .Z(n9510) );
  XNOR U9769 ( .A(n9511), .B(n9510), .Z(n9512) );
  XNOR U9770 ( .A(n9513), .B(n9512), .Z(n9531) );
  NAND U9771 ( .A(n33), .B(n9445), .Z(n9447) );
  XOR U9772 ( .A(b[5]), .B(a[126]), .Z(n9522) );
  NAND U9773 ( .A(n19342), .B(n9522), .Z(n9446) );
  AND U9774 ( .A(n9447), .B(n9446), .Z(n9507) );
  NAND U9775 ( .A(n34), .B(n9448), .Z(n9450) );
  XOR U9776 ( .A(b[7]), .B(a[124]), .Z(n9525) );
  NAND U9777 ( .A(n19486), .B(n9525), .Z(n9449) );
  AND U9778 ( .A(n9450), .B(n9449), .Z(n9505) );
  NAND U9779 ( .A(n31), .B(n9451), .Z(n9453) );
  XOR U9780 ( .A(b[3]), .B(a[128]), .Z(n9528) );
  NAND U9781 ( .A(n32), .B(n9528), .Z(n9452) );
  NAND U9782 ( .A(n9453), .B(n9452), .Z(n9504) );
  XNOR U9783 ( .A(n9505), .B(n9504), .Z(n9506) );
  XOR U9784 ( .A(n9507), .B(n9506), .Z(n9532) );
  XOR U9785 ( .A(n9531), .B(n9532), .Z(n9534) );
  XOR U9786 ( .A(n9533), .B(n9534), .Z(n9484) );
  NANDN U9787 ( .A(n9455), .B(n9454), .Z(n9459) );
  OR U9788 ( .A(n9457), .B(n9456), .Z(n9458) );
  AND U9789 ( .A(n9459), .B(n9458), .Z(n9483) );
  XNOR U9790 ( .A(n9484), .B(n9483), .Z(n9485) );
  XOR U9791 ( .A(n9486), .B(n9485), .Z(n9544) );
  NANDN U9792 ( .A(n9461), .B(n9460), .Z(n9465) );
  NANDN U9793 ( .A(n9463), .B(n9462), .Z(n9464) );
  AND U9794 ( .A(n9465), .B(n9464), .Z(n9543) );
  XNOR U9795 ( .A(n9544), .B(n9543), .Z(n9545) );
  XOR U9796 ( .A(n9546), .B(n9545), .Z(n9478) );
  NANDN U9797 ( .A(n9467), .B(n9466), .Z(n9471) );
  NAND U9798 ( .A(n9469), .B(n9468), .Z(n9470) );
  AND U9799 ( .A(n9471), .B(n9470), .Z(n9477) );
  XNOR U9800 ( .A(n9478), .B(n9477), .Z(n9479) );
  XNOR U9801 ( .A(n9480), .B(n9479), .Z(n9549) );
  XNOR U9802 ( .A(sreg[370]), .B(n9549), .Z(n9551) );
  NANDN U9803 ( .A(sreg[369]), .B(n9472), .Z(n9476) );
  NAND U9804 ( .A(n9474), .B(n9473), .Z(n9475) );
  NAND U9805 ( .A(n9476), .B(n9475), .Z(n9550) );
  XNOR U9806 ( .A(n9551), .B(n9550), .Z(c[370]) );
  NANDN U9807 ( .A(n9478), .B(n9477), .Z(n9482) );
  NANDN U9808 ( .A(n9480), .B(n9479), .Z(n9481) );
  AND U9809 ( .A(n9482), .B(n9481), .Z(n9557) );
  NANDN U9810 ( .A(n9484), .B(n9483), .Z(n9488) );
  NAND U9811 ( .A(n9486), .B(n9485), .Z(n9487) );
  AND U9812 ( .A(n9488), .B(n9487), .Z(n9623) );
  NAND U9813 ( .A(n9489), .B(n19724), .Z(n9491) );
  XOR U9814 ( .A(b[11]), .B(a[121]), .Z(n9593) );
  NAND U9815 ( .A(n19692), .B(n9593), .Z(n9490) );
  AND U9816 ( .A(n9491), .B(n9490), .Z(n9604) );
  NAND U9817 ( .A(n19838), .B(n9492), .Z(n9494) );
  XOR U9818 ( .A(b[15]), .B(a[117]), .Z(n9596) );
  NAND U9819 ( .A(n19805), .B(n9596), .Z(n9493) );
  AND U9820 ( .A(n9494), .B(n9493), .Z(n9603) );
  NAND U9821 ( .A(n35), .B(n9495), .Z(n9497) );
  XOR U9822 ( .A(b[9]), .B(a[123]), .Z(n9599) );
  NAND U9823 ( .A(n19598), .B(n9599), .Z(n9496) );
  NAND U9824 ( .A(n9497), .B(n9496), .Z(n9602) );
  XOR U9825 ( .A(n9603), .B(n9602), .Z(n9605) );
  XOR U9826 ( .A(n9604), .B(n9605), .Z(n9615) );
  NANDN U9827 ( .A(n9499), .B(n9498), .Z(n9503) );
  OR U9828 ( .A(n9501), .B(n9500), .Z(n9502) );
  AND U9829 ( .A(n9503), .B(n9502), .Z(n9614) );
  XNOR U9830 ( .A(n9615), .B(n9614), .Z(n9616) );
  NANDN U9831 ( .A(n9505), .B(n9504), .Z(n9509) );
  NANDN U9832 ( .A(n9507), .B(n9506), .Z(n9508) );
  NAND U9833 ( .A(n9509), .B(n9508), .Z(n9617) );
  XNOR U9834 ( .A(n9616), .B(n9617), .Z(n9563) );
  NANDN U9835 ( .A(n9511), .B(n9510), .Z(n9515) );
  NANDN U9836 ( .A(n9513), .B(n9512), .Z(n9514) );
  AND U9837 ( .A(n9515), .B(n9514), .Z(n9589) );
  NAND U9838 ( .A(n19808), .B(n9516), .Z(n9518) );
  XOR U9839 ( .A(b[13]), .B(a[119]), .Z(n9575) );
  NAND U9840 ( .A(n19768), .B(n9575), .Z(n9517) );
  AND U9841 ( .A(n9518), .B(n9517), .Z(n9567) );
  AND U9842 ( .A(b[15]), .B(a[115]), .Z(n9566) );
  XNOR U9843 ( .A(n9567), .B(n9566), .Z(n9568) );
  NAND U9844 ( .A(b[0]), .B(a[131]), .Z(n9519) );
  XNOR U9845 ( .A(b[1]), .B(n9519), .Z(n9521) );
  NANDN U9846 ( .A(b[0]), .B(a[130]), .Z(n9520) );
  NAND U9847 ( .A(n9521), .B(n9520), .Z(n9569) );
  XNOR U9848 ( .A(n9568), .B(n9569), .Z(n9587) );
  NAND U9849 ( .A(n33), .B(n9522), .Z(n9524) );
  XOR U9850 ( .A(b[5]), .B(a[127]), .Z(n9578) );
  NAND U9851 ( .A(n19342), .B(n9578), .Z(n9523) );
  AND U9852 ( .A(n9524), .B(n9523), .Z(n9611) );
  NAND U9853 ( .A(n34), .B(n9525), .Z(n9527) );
  XOR U9854 ( .A(b[7]), .B(a[125]), .Z(n9581) );
  NAND U9855 ( .A(n19486), .B(n9581), .Z(n9526) );
  AND U9856 ( .A(n9527), .B(n9526), .Z(n9609) );
  NAND U9857 ( .A(n31), .B(n9528), .Z(n9530) );
  XOR U9858 ( .A(b[3]), .B(a[129]), .Z(n9584) );
  NAND U9859 ( .A(n32), .B(n9584), .Z(n9529) );
  NAND U9860 ( .A(n9530), .B(n9529), .Z(n9608) );
  XNOR U9861 ( .A(n9609), .B(n9608), .Z(n9610) );
  XOR U9862 ( .A(n9611), .B(n9610), .Z(n9588) );
  XOR U9863 ( .A(n9587), .B(n9588), .Z(n9590) );
  XOR U9864 ( .A(n9589), .B(n9590), .Z(n9561) );
  NANDN U9865 ( .A(n9532), .B(n9531), .Z(n9536) );
  OR U9866 ( .A(n9534), .B(n9533), .Z(n9535) );
  AND U9867 ( .A(n9536), .B(n9535), .Z(n9560) );
  XNOR U9868 ( .A(n9561), .B(n9560), .Z(n9562) );
  XOR U9869 ( .A(n9563), .B(n9562), .Z(n9621) );
  NANDN U9870 ( .A(n9538), .B(n9537), .Z(n9542) );
  NANDN U9871 ( .A(n9540), .B(n9539), .Z(n9541) );
  AND U9872 ( .A(n9542), .B(n9541), .Z(n9620) );
  XNOR U9873 ( .A(n9621), .B(n9620), .Z(n9622) );
  XOR U9874 ( .A(n9623), .B(n9622), .Z(n9555) );
  NANDN U9875 ( .A(n9544), .B(n9543), .Z(n9548) );
  NAND U9876 ( .A(n9546), .B(n9545), .Z(n9547) );
  AND U9877 ( .A(n9548), .B(n9547), .Z(n9554) );
  XNOR U9878 ( .A(n9555), .B(n9554), .Z(n9556) );
  XNOR U9879 ( .A(n9557), .B(n9556), .Z(n9626) );
  XNOR U9880 ( .A(sreg[371]), .B(n9626), .Z(n9628) );
  NANDN U9881 ( .A(sreg[370]), .B(n9549), .Z(n9553) );
  NAND U9882 ( .A(n9551), .B(n9550), .Z(n9552) );
  NAND U9883 ( .A(n9553), .B(n9552), .Z(n9627) );
  XNOR U9884 ( .A(n9628), .B(n9627), .Z(c[371]) );
  NANDN U9885 ( .A(n9555), .B(n9554), .Z(n9559) );
  NANDN U9886 ( .A(n9557), .B(n9556), .Z(n9558) );
  AND U9887 ( .A(n9559), .B(n9558), .Z(n9634) );
  NANDN U9888 ( .A(n9561), .B(n9560), .Z(n9565) );
  NAND U9889 ( .A(n9563), .B(n9562), .Z(n9564) );
  AND U9890 ( .A(n9565), .B(n9564), .Z(n9700) );
  NANDN U9891 ( .A(n9567), .B(n9566), .Z(n9571) );
  NANDN U9892 ( .A(n9569), .B(n9568), .Z(n9570) );
  AND U9893 ( .A(n9571), .B(n9570), .Z(n9666) );
  NAND U9894 ( .A(b[0]), .B(a[132]), .Z(n9572) );
  XNOR U9895 ( .A(b[1]), .B(n9572), .Z(n9574) );
  NANDN U9896 ( .A(b[0]), .B(a[131]), .Z(n9573) );
  NAND U9897 ( .A(n9574), .B(n9573), .Z(n9646) );
  NAND U9898 ( .A(n19808), .B(n9575), .Z(n9577) );
  XOR U9899 ( .A(b[13]), .B(a[120]), .Z(n9652) );
  NAND U9900 ( .A(n19768), .B(n9652), .Z(n9576) );
  AND U9901 ( .A(n9577), .B(n9576), .Z(n9644) );
  AND U9902 ( .A(b[15]), .B(a[116]), .Z(n9643) );
  XNOR U9903 ( .A(n9644), .B(n9643), .Z(n9645) );
  XNOR U9904 ( .A(n9646), .B(n9645), .Z(n9664) );
  NAND U9905 ( .A(n33), .B(n9578), .Z(n9580) );
  XOR U9906 ( .A(b[5]), .B(a[128]), .Z(n9655) );
  NAND U9907 ( .A(n19342), .B(n9655), .Z(n9579) );
  AND U9908 ( .A(n9580), .B(n9579), .Z(n9688) );
  NAND U9909 ( .A(n34), .B(n9581), .Z(n9583) );
  XOR U9910 ( .A(b[7]), .B(a[126]), .Z(n9658) );
  NAND U9911 ( .A(n19486), .B(n9658), .Z(n9582) );
  AND U9912 ( .A(n9583), .B(n9582), .Z(n9686) );
  NAND U9913 ( .A(n31), .B(n9584), .Z(n9586) );
  XOR U9914 ( .A(b[3]), .B(a[130]), .Z(n9661) );
  NAND U9915 ( .A(n32), .B(n9661), .Z(n9585) );
  NAND U9916 ( .A(n9586), .B(n9585), .Z(n9685) );
  XNOR U9917 ( .A(n9686), .B(n9685), .Z(n9687) );
  XOR U9918 ( .A(n9688), .B(n9687), .Z(n9665) );
  XOR U9919 ( .A(n9664), .B(n9665), .Z(n9667) );
  XOR U9920 ( .A(n9666), .B(n9667), .Z(n9638) );
  NANDN U9921 ( .A(n9588), .B(n9587), .Z(n9592) );
  OR U9922 ( .A(n9590), .B(n9589), .Z(n9591) );
  AND U9923 ( .A(n9592), .B(n9591), .Z(n9637) );
  XNOR U9924 ( .A(n9638), .B(n9637), .Z(n9640) );
  NAND U9925 ( .A(n9593), .B(n19724), .Z(n9595) );
  XOR U9926 ( .A(b[11]), .B(a[122]), .Z(n9670) );
  NAND U9927 ( .A(n19692), .B(n9670), .Z(n9594) );
  AND U9928 ( .A(n9595), .B(n9594), .Z(n9681) );
  NAND U9929 ( .A(n19838), .B(n9596), .Z(n9598) );
  XOR U9930 ( .A(b[15]), .B(a[118]), .Z(n9673) );
  NAND U9931 ( .A(n19805), .B(n9673), .Z(n9597) );
  AND U9932 ( .A(n9598), .B(n9597), .Z(n9680) );
  NAND U9933 ( .A(n35), .B(n9599), .Z(n9601) );
  XOR U9934 ( .A(b[9]), .B(a[124]), .Z(n9676) );
  NAND U9935 ( .A(n19598), .B(n9676), .Z(n9600) );
  NAND U9936 ( .A(n9601), .B(n9600), .Z(n9679) );
  XOR U9937 ( .A(n9680), .B(n9679), .Z(n9682) );
  XOR U9938 ( .A(n9681), .B(n9682), .Z(n9692) );
  NANDN U9939 ( .A(n9603), .B(n9602), .Z(n9607) );
  OR U9940 ( .A(n9605), .B(n9604), .Z(n9606) );
  AND U9941 ( .A(n9607), .B(n9606), .Z(n9691) );
  XNOR U9942 ( .A(n9692), .B(n9691), .Z(n9693) );
  NANDN U9943 ( .A(n9609), .B(n9608), .Z(n9613) );
  NANDN U9944 ( .A(n9611), .B(n9610), .Z(n9612) );
  NAND U9945 ( .A(n9613), .B(n9612), .Z(n9694) );
  XNOR U9946 ( .A(n9693), .B(n9694), .Z(n9639) );
  XOR U9947 ( .A(n9640), .B(n9639), .Z(n9698) );
  NANDN U9948 ( .A(n9615), .B(n9614), .Z(n9619) );
  NANDN U9949 ( .A(n9617), .B(n9616), .Z(n9618) );
  AND U9950 ( .A(n9619), .B(n9618), .Z(n9697) );
  XNOR U9951 ( .A(n9698), .B(n9697), .Z(n9699) );
  XOR U9952 ( .A(n9700), .B(n9699), .Z(n9632) );
  NANDN U9953 ( .A(n9621), .B(n9620), .Z(n9625) );
  NAND U9954 ( .A(n9623), .B(n9622), .Z(n9624) );
  AND U9955 ( .A(n9625), .B(n9624), .Z(n9631) );
  XNOR U9956 ( .A(n9632), .B(n9631), .Z(n9633) );
  XNOR U9957 ( .A(n9634), .B(n9633), .Z(n9703) );
  XNOR U9958 ( .A(sreg[372]), .B(n9703), .Z(n9705) );
  NANDN U9959 ( .A(sreg[371]), .B(n9626), .Z(n9630) );
  NAND U9960 ( .A(n9628), .B(n9627), .Z(n9629) );
  NAND U9961 ( .A(n9630), .B(n9629), .Z(n9704) );
  XNOR U9962 ( .A(n9705), .B(n9704), .Z(c[372]) );
  NANDN U9963 ( .A(n9632), .B(n9631), .Z(n9636) );
  NANDN U9964 ( .A(n9634), .B(n9633), .Z(n9635) );
  AND U9965 ( .A(n9636), .B(n9635), .Z(n9711) );
  NANDN U9966 ( .A(n9638), .B(n9637), .Z(n9642) );
  NAND U9967 ( .A(n9640), .B(n9639), .Z(n9641) );
  AND U9968 ( .A(n9642), .B(n9641), .Z(n9777) );
  NANDN U9969 ( .A(n9644), .B(n9643), .Z(n9648) );
  NANDN U9970 ( .A(n9646), .B(n9645), .Z(n9647) );
  AND U9971 ( .A(n9648), .B(n9647), .Z(n9743) );
  NAND U9972 ( .A(b[0]), .B(a[133]), .Z(n9649) );
  XNOR U9973 ( .A(b[1]), .B(n9649), .Z(n9651) );
  NANDN U9974 ( .A(b[0]), .B(a[132]), .Z(n9650) );
  NAND U9975 ( .A(n9651), .B(n9650), .Z(n9723) );
  NAND U9976 ( .A(n19808), .B(n9652), .Z(n9654) );
  XOR U9977 ( .A(b[13]), .B(a[121]), .Z(n9729) );
  NAND U9978 ( .A(n19768), .B(n9729), .Z(n9653) );
  AND U9979 ( .A(n9654), .B(n9653), .Z(n9721) );
  AND U9980 ( .A(b[15]), .B(a[117]), .Z(n9720) );
  XNOR U9981 ( .A(n9721), .B(n9720), .Z(n9722) );
  XNOR U9982 ( .A(n9723), .B(n9722), .Z(n9741) );
  NAND U9983 ( .A(n33), .B(n9655), .Z(n9657) );
  XOR U9984 ( .A(b[5]), .B(a[129]), .Z(n9732) );
  NAND U9985 ( .A(n19342), .B(n9732), .Z(n9656) );
  AND U9986 ( .A(n9657), .B(n9656), .Z(n9765) );
  NAND U9987 ( .A(n34), .B(n9658), .Z(n9660) );
  XOR U9988 ( .A(b[7]), .B(a[127]), .Z(n9735) );
  NAND U9989 ( .A(n19486), .B(n9735), .Z(n9659) );
  AND U9990 ( .A(n9660), .B(n9659), .Z(n9763) );
  NAND U9991 ( .A(n31), .B(n9661), .Z(n9663) );
  XOR U9992 ( .A(b[3]), .B(a[131]), .Z(n9738) );
  NAND U9993 ( .A(n32), .B(n9738), .Z(n9662) );
  NAND U9994 ( .A(n9663), .B(n9662), .Z(n9762) );
  XNOR U9995 ( .A(n9763), .B(n9762), .Z(n9764) );
  XOR U9996 ( .A(n9765), .B(n9764), .Z(n9742) );
  XOR U9997 ( .A(n9741), .B(n9742), .Z(n9744) );
  XOR U9998 ( .A(n9743), .B(n9744), .Z(n9715) );
  NANDN U9999 ( .A(n9665), .B(n9664), .Z(n9669) );
  OR U10000 ( .A(n9667), .B(n9666), .Z(n9668) );
  AND U10001 ( .A(n9669), .B(n9668), .Z(n9714) );
  XNOR U10002 ( .A(n9715), .B(n9714), .Z(n9717) );
  NAND U10003 ( .A(n9670), .B(n19724), .Z(n9672) );
  XOR U10004 ( .A(b[11]), .B(a[123]), .Z(n9747) );
  NAND U10005 ( .A(n19692), .B(n9747), .Z(n9671) );
  AND U10006 ( .A(n9672), .B(n9671), .Z(n9758) );
  NAND U10007 ( .A(n19838), .B(n9673), .Z(n9675) );
  XOR U10008 ( .A(b[15]), .B(a[119]), .Z(n9750) );
  NAND U10009 ( .A(n19805), .B(n9750), .Z(n9674) );
  AND U10010 ( .A(n9675), .B(n9674), .Z(n9757) );
  NAND U10011 ( .A(n35), .B(n9676), .Z(n9678) );
  XOR U10012 ( .A(b[9]), .B(a[125]), .Z(n9753) );
  NAND U10013 ( .A(n19598), .B(n9753), .Z(n9677) );
  NAND U10014 ( .A(n9678), .B(n9677), .Z(n9756) );
  XOR U10015 ( .A(n9757), .B(n9756), .Z(n9759) );
  XOR U10016 ( .A(n9758), .B(n9759), .Z(n9769) );
  NANDN U10017 ( .A(n9680), .B(n9679), .Z(n9684) );
  OR U10018 ( .A(n9682), .B(n9681), .Z(n9683) );
  AND U10019 ( .A(n9684), .B(n9683), .Z(n9768) );
  XNOR U10020 ( .A(n9769), .B(n9768), .Z(n9770) );
  NANDN U10021 ( .A(n9686), .B(n9685), .Z(n9690) );
  NANDN U10022 ( .A(n9688), .B(n9687), .Z(n9689) );
  NAND U10023 ( .A(n9690), .B(n9689), .Z(n9771) );
  XNOR U10024 ( .A(n9770), .B(n9771), .Z(n9716) );
  XOR U10025 ( .A(n9717), .B(n9716), .Z(n9775) );
  NANDN U10026 ( .A(n9692), .B(n9691), .Z(n9696) );
  NANDN U10027 ( .A(n9694), .B(n9693), .Z(n9695) );
  AND U10028 ( .A(n9696), .B(n9695), .Z(n9774) );
  XNOR U10029 ( .A(n9775), .B(n9774), .Z(n9776) );
  XOR U10030 ( .A(n9777), .B(n9776), .Z(n9709) );
  NANDN U10031 ( .A(n9698), .B(n9697), .Z(n9702) );
  NAND U10032 ( .A(n9700), .B(n9699), .Z(n9701) );
  AND U10033 ( .A(n9702), .B(n9701), .Z(n9708) );
  XNOR U10034 ( .A(n9709), .B(n9708), .Z(n9710) );
  XNOR U10035 ( .A(n9711), .B(n9710), .Z(n9780) );
  XNOR U10036 ( .A(sreg[373]), .B(n9780), .Z(n9782) );
  NANDN U10037 ( .A(sreg[372]), .B(n9703), .Z(n9707) );
  NAND U10038 ( .A(n9705), .B(n9704), .Z(n9706) );
  NAND U10039 ( .A(n9707), .B(n9706), .Z(n9781) );
  XNOR U10040 ( .A(n9782), .B(n9781), .Z(c[373]) );
  NANDN U10041 ( .A(n9709), .B(n9708), .Z(n9713) );
  NANDN U10042 ( .A(n9711), .B(n9710), .Z(n9712) );
  AND U10043 ( .A(n9713), .B(n9712), .Z(n9788) );
  NANDN U10044 ( .A(n9715), .B(n9714), .Z(n9719) );
  NAND U10045 ( .A(n9717), .B(n9716), .Z(n9718) );
  AND U10046 ( .A(n9719), .B(n9718), .Z(n9854) );
  NANDN U10047 ( .A(n9721), .B(n9720), .Z(n9725) );
  NANDN U10048 ( .A(n9723), .B(n9722), .Z(n9724) );
  AND U10049 ( .A(n9725), .B(n9724), .Z(n9820) );
  NAND U10050 ( .A(b[0]), .B(a[134]), .Z(n9726) );
  XNOR U10051 ( .A(b[1]), .B(n9726), .Z(n9728) );
  NANDN U10052 ( .A(b[0]), .B(a[133]), .Z(n9727) );
  NAND U10053 ( .A(n9728), .B(n9727), .Z(n9800) );
  NAND U10054 ( .A(n19808), .B(n9729), .Z(n9731) );
  XOR U10055 ( .A(b[13]), .B(a[122]), .Z(n9806) );
  NAND U10056 ( .A(n19768), .B(n9806), .Z(n9730) );
  AND U10057 ( .A(n9731), .B(n9730), .Z(n9798) );
  AND U10058 ( .A(b[15]), .B(a[118]), .Z(n9797) );
  XNOR U10059 ( .A(n9798), .B(n9797), .Z(n9799) );
  XNOR U10060 ( .A(n9800), .B(n9799), .Z(n9818) );
  NAND U10061 ( .A(n33), .B(n9732), .Z(n9734) );
  XOR U10062 ( .A(b[5]), .B(a[130]), .Z(n9809) );
  NAND U10063 ( .A(n19342), .B(n9809), .Z(n9733) );
  AND U10064 ( .A(n9734), .B(n9733), .Z(n9842) );
  NAND U10065 ( .A(n34), .B(n9735), .Z(n9737) );
  XOR U10066 ( .A(b[7]), .B(a[128]), .Z(n9812) );
  NAND U10067 ( .A(n19486), .B(n9812), .Z(n9736) );
  AND U10068 ( .A(n9737), .B(n9736), .Z(n9840) );
  NAND U10069 ( .A(n31), .B(n9738), .Z(n9740) );
  XOR U10070 ( .A(b[3]), .B(a[132]), .Z(n9815) );
  NAND U10071 ( .A(n32), .B(n9815), .Z(n9739) );
  NAND U10072 ( .A(n9740), .B(n9739), .Z(n9839) );
  XNOR U10073 ( .A(n9840), .B(n9839), .Z(n9841) );
  XOR U10074 ( .A(n9842), .B(n9841), .Z(n9819) );
  XOR U10075 ( .A(n9818), .B(n9819), .Z(n9821) );
  XOR U10076 ( .A(n9820), .B(n9821), .Z(n9792) );
  NANDN U10077 ( .A(n9742), .B(n9741), .Z(n9746) );
  OR U10078 ( .A(n9744), .B(n9743), .Z(n9745) );
  AND U10079 ( .A(n9746), .B(n9745), .Z(n9791) );
  XNOR U10080 ( .A(n9792), .B(n9791), .Z(n9794) );
  NAND U10081 ( .A(n9747), .B(n19724), .Z(n9749) );
  XOR U10082 ( .A(b[11]), .B(a[124]), .Z(n9824) );
  NAND U10083 ( .A(n19692), .B(n9824), .Z(n9748) );
  AND U10084 ( .A(n9749), .B(n9748), .Z(n9835) );
  NAND U10085 ( .A(n19838), .B(n9750), .Z(n9752) );
  XOR U10086 ( .A(b[15]), .B(a[120]), .Z(n9827) );
  NAND U10087 ( .A(n19805), .B(n9827), .Z(n9751) );
  AND U10088 ( .A(n9752), .B(n9751), .Z(n9834) );
  NAND U10089 ( .A(n35), .B(n9753), .Z(n9755) );
  XOR U10090 ( .A(b[9]), .B(a[126]), .Z(n9830) );
  NAND U10091 ( .A(n19598), .B(n9830), .Z(n9754) );
  NAND U10092 ( .A(n9755), .B(n9754), .Z(n9833) );
  XOR U10093 ( .A(n9834), .B(n9833), .Z(n9836) );
  XOR U10094 ( .A(n9835), .B(n9836), .Z(n9846) );
  NANDN U10095 ( .A(n9757), .B(n9756), .Z(n9761) );
  OR U10096 ( .A(n9759), .B(n9758), .Z(n9760) );
  AND U10097 ( .A(n9761), .B(n9760), .Z(n9845) );
  XNOR U10098 ( .A(n9846), .B(n9845), .Z(n9847) );
  NANDN U10099 ( .A(n9763), .B(n9762), .Z(n9767) );
  NANDN U10100 ( .A(n9765), .B(n9764), .Z(n9766) );
  NAND U10101 ( .A(n9767), .B(n9766), .Z(n9848) );
  XNOR U10102 ( .A(n9847), .B(n9848), .Z(n9793) );
  XOR U10103 ( .A(n9794), .B(n9793), .Z(n9852) );
  NANDN U10104 ( .A(n9769), .B(n9768), .Z(n9773) );
  NANDN U10105 ( .A(n9771), .B(n9770), .Z(n9772) );
  AND U10106 ( .A(n9773), .B(n9772), .Z(n9851) );
  XNOR U10107 ( .A(n9852), .B(n9851), .Z(n9853) );
  XOR U10108 ( .A(n9854), .B(n9853), .Z(n9786) );
  NANDN U10109 ( .A(n9775), .B(n9774), .Z(n9779) );
  NAND U10110 ( .A(n9777), .B(n9776), .Z(n9778) );
  AND U10111 ( .A(n9779), .B(n9778), .Z(n9785) );
  XNOR U10112 ( .A(n9786), .B(n9785), .Z(n9787) );
  XNOR U10113 ( .A(n9788), .B(n9787), .Z(n9857) );
  XNOR U10114 ( .A(sreg[374]), .B(n9857), .Z(n9859) );
  NANDN U10115 ( .A(sreg[373]), .B(n9780), .Z(n9784) );
  NAND U10116 ( .A(n9782), .B(n9781), .Z(n9783) );
  NAND U10117 ( .A(n9784), .B(n9783), .Z(n9858) );
  XNOR U10118 ( .A(n9859), .B(n9858), .Z(c[374]) );
  NANDN U10119 ( .A(n9786), .B(n9785), .Z(n9790) );
  NANDN U10120 ( .A(n9788), .B(n9787), .Z(n9789) );
  AND U10121 ( .A(n9790), .B(n9789), .Z(n9865) );
  NANDN U10122 ( .A(n9792), .B(n9791), .Z(n9796) );
  NAND U10123 ( .A(n9794), .B(n9793), .Z(n9795) );
  AND U10124 ( .A(n9796), .B(n9795), .Z(n9931) );
  NANDN U10125 ( .A(n9798), .B(n9797), .Z(n9802) );
  NANDN U10126 ( .A(n9800), .B(n9799), .Z(n9801) );
  AND U10127 ( .A(n9802), .B(n9801), .Z(n9897) );
  NAND U10128 ( .A(b[0]), .B(a[135]), .Z(n9803) );
  XNOR U10129 ( .A(b[1]), .B(n9803), .Z(n9805) );
  NANDN U10130 ( .A(b[0]), .B(a[134]), .Z(n9804) );
  NAND U10131 ( .A(n9805), .B(n9804), .Z(n9877) );
  NAND U10132 ( .A(n19808), .B(n9806), .Z(n9808) );
  XOR U10133 ( .A(b[13]), .B(a[123]), .Z(n9880) );
  NAND U10134 ( .A(n19768), .B(n9880), .Z(n9807) );
  AND U10135 ( .A(n9808), .B(n9807), .Z(n9875) );
  AND U10136 ( .A(b[15]), .B(a[119]), .Z(n9874) );
  XNOR U10137 ( .A(n9875), .B(n9874), .Z(n9876) );
  XNOR U10138 ( .A(n9877), .B(n9876), .Z(n9895) );
  NAND U10139 ( .A(n33), .B(n9809), .Z(n9811) );
  XOR U10140 ( .A(b[5]), .B(a[131]), .Z(n9886) );
  NAND U10141 ( .A(n19342), .B(n9886), .Z(n9810) );
  AND U10142 ( .A(n9811), .B(n9810), .Z(n9919) );
  NAND U10143 ( .A(n34), .B(n9812), .Z(n9814) );
  XOR U10144 ( .A(b[7]), .B(a[129]), .Z(n9889) );
  NAND U10145 ( .A(n19486), .B(n9889), .Z(n9813) );
  AND U10146 ( .A(n9814), .B(n9813), .Z(n9917) );
  NAND U10147 ( .A(n31), .B(n9815), .Z(n9817) );
  XOR U10148 ( .A(b[3]), .B(a[133]), .Z(n9892) );
  NAND U10149 ( .A(n32), .B(n9892), .Z(n9816) );
  NAND U10150 ( .A(n9817), .B(n9816), .Z(n9916) );
  XNOR U10151 ( .A(n9917), .B(n9916), .Z(n9918) );
  XOR U10152 ( .A(n9919), .B(n9918), .Z(n9896) );
  XOR U10153 ( .A(n9895), .B(n9896), .Z(n9898) );
  XOR U10154 ( .A(n9897), .B(n9898), .Z(n9869) );
  NANDN U10155 ( .A(n9819), .B(n9818), .Z(n9823) );
  OR U10156 ( .A(n9821), .B(n9820), .Z(n9822) );
  AND U10157 ( .A(n9823), .B(n9822), .Z(n9868) );
  XNOR U10158 ( .A(n9869), .B(n9868), .Z(n9871) );
  NAND U10159 ( .A(n9824), .B(n19724), .Z(n9826) );
  XOR U10160 ( .A(b[11]), .B(a[125]), .Z(n9901) );
  NAND U10161 ( .A(n19692), .B(n9901), .Z(n9825) );
  AND U10162 ( .A(n9826), .B(n9825), .Z(n9912) );
  NAND U10163 ( .A(n19838), .B(n9827), .Z(n9829) );
  XOR U10164 ( .A(b[15]), .B(a[121]), .Z(n9904) );
  NAND U10165 ( .A(n19805), .B(n9904), .Z(n9828) );
  AND U10166 ( .A(n9829), .B(n9828), .Z(n9911) );
  NAND U10167 ( .A(n35), .B(n9830), .Z(n9832) );
  XOR U10168 ( .A(b[9]), .B(a[127]), .Z(n9907) );
  NAND U10169 ( .A(n19598), .B(n9907), .Z(n9831) );
  NAND U10170 ( .A(n9832), .B(n9831), .Z(n9910) );
  XOR U10171 ( .A(n9911), .B(n9910), .Z(n9913) );
  XOR U10172 ( .A(n9912), .B(n9913), .Z(n9923) );
  NANDN U10173 ( .A(n9834), .B(n9833), .Z(n9838) );
  OR U10174 ( .A(n9836), .B(n9835), .Z(n9837) );
  AND U10175 ( .A(n9838), .B(n9837), .Z(n9922) );
  XNOR U10176 ( .A(n9923), .B(n9922), .Z(n9924) );
  NANDN U10177 ( .A(n9840), .B(n9839), .Z(n9844) );
  NANDN U10178 ( .A(n9842), .B(n9841), .Z(n9843) );
  NAND U10179 ( .A(n9844), .B(n9843), .Z(n9925) );
  XNOR U10180 ( .A(n9924), .B(n9925), .Z(n9870) );
  XOR U10181 ( .A(n9871), .B(n9870), .Z(n9929) );
  NANDN U10182 ( .A(n9846), .B(n9845), .Z(n9850) );
  NANDN U10183 ( .A(n9848), .B(n9847), .Z(n9849) );
  AND U10184 ( .A(n9850), .B(n9849), .Z(n9928) );
  XNOR U10185 ( .A(n9929), .B(n9928), .Z(n9930) );
  XOR U10186 ( .A(n9931), .B(n9930), .Z(n9863) );
  NANDN U10187 ( .A(n9852), .B(n9851), .Z(n9856) );
  NAND U10188 ( .A(n9854), .B(n9853), .Z(n9855) );
  AND U10189 ( .A(n9856), .B(n9855), .Z(n9862) );
  XNOR U10190 ( .A(n9863), .B(n9862), .Z(n9864) );
  XNOR U10191 ( .A(n9865), .B(n9864), .Z(n9934) );
  XNOR U10192 ( .A(sreg[375]), .B(n9934), .Z(n9936) );
  NANDN U10193 ( .A(sreg[374]), .B(n9857), .Z(n9861) );
  NAND U10194 ( .A(n9859), .B(n9858), .Z(n9860) );
  NAND U10195 ( .A(n9861), .B(n9860), .Z(n9935) );
  XNOR U10196 ( .A(n9936), .B(n9935), .Z(c[375]) );
  NANDN U10197 ( .A(n9863), .B(n9862), .Z(n9867) );
  NANDN U10198 ( .A(n9865), .B(n9864), .Z(n9866) );
  AND U10199 ( .A(n9867), .B(n9866), .Z(n9942) );
  NANDN U10200 ( .A(n9869), .B(n9868), .Z(n9873) );
  NAND U10201 ( .A(n9871), .B(n9870), .Z(n9872) );
  AND U10202 ( .A(n9873), .B(n9872), .Z(n10008) );
  NANDN U10203 ( .A(n9875), .B(n9874), .Z(n9879) );
  NANDN U10204 ( .A(n9877), .B(n9876), .Z(n9878) );
  AND U10205 ( .A(n9879), .B(n9878), .Z(n9974) );
  NAND U10206 ( .A(n19808), .B(n9880), .Z(n9882) );
  XOR U10207 ( .A(b[13]), .B(a[124]), .Z(n9960) );
  NAND U10208 ( .A(n19768), .B(n9960), .Z(n9881) );
  AND U10209 ( .A(n9882), .B(n9881), .Z(n9952) );
  AND U10210 ( .A(b[15]), .B(a[120]), .Z(n9951) );
  XNOR U10211 ( .A(n9952), .B(n9951), .Z(n9953) );
  NAND U10212 ( .A(b[0]), .B(a[136]), .Z(n9883) );
  XNOR U10213 ( .A(b[1]), .B(n9883), .Z(n9885) );
  NANDN U10214 ( .A(b[0]), .B(a[135]), .Z(n9884) );
  NAND U10215 ( .A(n9885), .B(n9884), .Z(n9954) );
  XNOR U10216 ( .A(n9953), .B(n9954), .Z(n9972) );
  NAND U10217 ( .A(n33), .B(n9886), .Z(n9888) );
  XOR U10218 ( .A(b[5]), .B(a[132]), .Z(n9963) );
  NAND U10219 ( .A(n19342), .B(n9963), .Z(n9887) );
  AND U10220 ( .A(n9888), .B(n9887), .Z(n9996) );
  NAND U10221 ( .A(n34), .B(n9889), .Z(n9891) );
  XOR U10222 ( .A(b[7]), .B(a[130]), .Z(n9966) );
  NAND U10223 ( .A(n19486), .B(n9966), .Z(n9890) );
  AND U10224 ( .A(n9891), .B(n9890), .Z(n9994) );
  NAND U10225 ( .A(n31), .B(n9892), .Z(n9894) );
  XOR U10226 ( .A(b[3]), .B(a[134]), .Z(n9969) );
  NAND U10227 ( .A(n32), .B(n9969), .Z(n9893) );
  NAND U10228 ( .A(n9894), .B(n9893), .Z(n9993) );
  XNOR U10229 ( .A(n9994), .B(n9993), .Z(n9995) );
  XOR U10230 ( .A(n9996), .B(n9995), .Z(n9973) );
  XOR U10231 ( .A(n9972), .B(n9973), .Z(n9975) );
  XOR U10232 ( .A(n9974), .B(n9975), .Z(n9946) );
  NANDN U10233 ( .A(n9896), .B(n9895), .Z(n9900) );
  OR U10234 ( .A(n9898), .B(n9897), .Z(n9899) );
  AND U10235 ( .A(n9900), .B(n9899), .Z(n9945) );
  XNOR U10236 ( .A(n9946), .B(n9945), .Z(n9948) );
  NAND U10237 ( .A(n9901), .B(n19724), .Z(n9903) );
  XOR U10238 ( .A(b[11]), .B(a[126]), .Z(n9978) );
  NAND U10239 ( .A(n19692), .B(n9978), .Z(n9902) );
  AND U10240 ( .A(n9903), .B(n9902), .Z(n9989) );
  NAND U10241 ( .A(n19838), .B(n9904), .Z(n9906) );
  XOR U10242 ( .A(b[15]), .B(a[122]), .Z(n9981) );
  NAND U10243 ( .A(n19805), .B(n9981), .Z(n9905) );
  AND U10244 ( .A(n9906), .B(n9905), .Z(n9988) );
  NAND U10245 ( .A(n35), .B(n9907), .Z(n9909) );
  XOR U10246 ( .A(b[9]), .B(a[128]), .Z(n9984) );
  NAND U10247 ( .A(n19598), .B(n9984), .Z(n9908) );
  NAND U10248 ( .A(n9909), .B(n9908), .Z(n9987) );
  XOR U10249 ( .A(n9988), .B(n9987), .Z(n9990) );
  XOR U10250 ( .A(n9989), .B(n9990), .Z(n10000) );
  NANDN U10251 ( .A(n9911), .B(n9910), .Z(n9915) );
  OR U10252 ( .A(n9913), .B(n9912), .Z(n9914) );
  AND U10253 ( .A(n9915), .B(n9914), .Z(n9999) );
  XNOR U10254 ( .A(n10000), .B(n9999), .Z(n10001) );
  NANDN U10255 ( .A(n9917), .B(n9916), .Z(n9921) );
  NANDN U10256 ( .A(n9919), .B(n9918), .Z(n9920) );
  NAND U10257 ( .A(n9921), .B(n9920), .Z(n10002) );
  XNOR U10258 ( .A(n10001), .B(n10002), .Z(n9947) );
  XOR U10259 ( .A(n9948), .B(n9947), .Z(n10006) );
  NANDN U10260 ( .A(n9923), .B(n9922), .Z(n9927) );
  NANDN U10261 ( .A(n9925), .B(n9924), .Z(n9926) );
  AND U10262 ( .A(n9927), .B(n9926), .Z(n10005) );
  XNOR U10263 ( .A(n10006), .B(n10005), .Z(n10007) );
  XOR U10264 ( .A(n10008), .B(n10007), .Z(n9940) );
  NANDN U10265 ( .A(n9929), .B(n9928), .Z(n9933) );
  NAND U10266 ( .A(n9931), .B(n9930), .Z(n9932) );
  AND U10267 ( .A(n9933), .B(n9932), .Z(n9939) );
  XNOR U10268 ( .A(n9940), .B(n9939), .Z(n9941) );
  XNOR U10269 ( .A(n9942), .B(n9941), .Z(n10011) );
  XNOR U10270 ( .A(sreg[376]), .B(n10011), .Z(n10013) );
  NANDN U10271 ( .A(sreg[375]), .B(n9934), .Z(n9938) );
  NAND U10272 ( .A(n9936), .B(n9935), .Z(n9937) );
  NAND U10273 ( .A(n9938), .B(n9937), .Z(n10012) );
  XNOR U10274 ( .A(n10013), .B(n10012), .Z(c[376]) );
  NANDN U10275 ( .A(n9940), .B(n9939), .Z(n9944) );
  NANDN U10276 ( .A(n9942), .B(n9941), .Z(n9943) );
  AND U10277 ( .A(n9944), .B(n9943), .Z(n10024) );
  NANDN U10278 ( .A(n9946), .B(n9945), .Z(n9950) );
  NAND U10279 ( .A(n9948), .B(n9947), .Z(n9949) );
  AND U10280 ( .A(n9950), .B(n9949), .Z(n10090) );
  NANDN U10281 ( .A(n9952), .B(n9951), .Z(n9956) );
  NANDN U10282 ( .A(n9954), .B(n9953), .Z(n9955) );
  AND U10283 ( .A(n9956), .B(n9955), .Z(n10056) );
  NAND U10284 ( .A(b[0]), .B(a[137]), .Z(n9957) );
  XNOR U10285 ( .A(b[1]), .B(n9957), .Z(n9959) );
  NANDN U10286 ( .A(b[0]), .B(a[136]), .Z(n9958) );
  NAND U10287 ( .A(n9959), .B(n9958), .Z(n10036) );
  NAND U10288 ( .A(n19808), .B(n9960), .Z(n9962) );
  XOR U10289 ( .A(b[13]), .B(a[125]), .Z(n10039) );
  NAND U10290 ( .A(n19768), .B(n10039), .Z(n9961) );
  AND U10291 ( .A(n9962), .B(n9961), .Z(n10034) );
  AND U10292 ( .A(b[15]), .B(a[121]), .Z(n10033) );
  XNOR U10293 ( .A(n10034), .B(n10033), .Z(n10035) );
  XNOR U10294 ( .A(n10036), .B(n10035), .Z(n10054) );
  NAND U10295 ( .A(n33), .B(n9963), .Z(n9965) );
  XOR U10296 ( .A(b[5]), .B(a[133]), .Z(n10045) );
  NAND U10297 ( .A(n19342), .B(n10045), .Z(n9964) );
  AND U10298 ( .A(n9965), .B(n9964), .Z(n10078) );
  NAND U10299 ( .A(n34), .B(n9966), .Z(n9968) );
  XOR U10300 ( .A(b[7]), .B(a[131]), .Z(n10048) );
  NAND U10301 ( .A(n19486), .B(n10048), .Z(n9967) );
  AND U10302 ( .A(n9968), .B(n9967), .Z(n10076) );
  NAND U10303 ( .A(n31), .B(n9969), .Z(n9971) );
  XOR U10304 ( .A(b[3]), .B(a[135]), .Z(n10051) );
  NAND U10305 ( .A(n32), .B(n10051), .Z(n9970) );
  NAND U10306 ( .A(n9971), .B(n9970), .Z(n10075) );
  XNOR U10307 ( .A(n10076), .B(n10075), .Z(n10077) );
  XOR U10308 ( .A(n10078), .B(n10077), .Z(n10055) );
  XOR U10309 ( .A(n10054), .B(n10055), .Z(n10057) );
  XOR U10310 ( .A(n10056), .B(n10057), .Z(n10028) );
  NANDN U10311 ( .A(n9973), .B(n9972), .Z(n9977) );
  OR U10312 ( .A(n9975), .B(n9974), .Z(n9976) );
  AND U10313 ( .A(n9977), .B(n9976), .Z(n10027) );
  XNOR U10314 ( .A(n10028), .B(n10027), .Z(n10030) );
  NAND U10315 ( .A(n9978), .B(n19724), .Z(n9980) );
  XOR U10316 ( .A(b[11]), .B(a[127]), .Z(n10060) );
  NAND U10317 ( .A(n19692), .B(n10060), .Z(n9979) );
  AND U10318 ( .A(n9980), .B(n9979), .Z(n10071) );
  NAND U10319 ( .A(n19838), .B(n9981), .Z(n9983) );
  XOR U10320 ( .A(b[15]), .B(a[123]), .Z(n10063) );
  NAND U10321 ( .A(n19805), .B(n10063), .Z(n9982) );
  AND U10322 ( .A(n9983), .B(n9982), .Z(n10070) );
  NAND U10323 ( .A(n35), .B(n9984), .Z(n9986) );
  XOR U10324 ( .A(b[9]), .B(a[129]), .Z(n10066) );
  NAND U10325 ( .A(n19598), .B(n10066), .Z(n9985) );
  NAND U10326 ( .A(n9986), .B(n9985), .Z(n10069) );
  XOR U10327 ( .A(n10070), .B(n10069), .Z(n10072) );
  XOR U10328 ( .A(n10071), .B(n10072), .Z(n10082) );
  NANDN U10329 ( .A(n9988), .B(n9987), .Z(n9992) );
  OR U10330 ( .A(n9990), .B(n9989), .Z(n9991) );
  AND U10331 ( .A(n9992), .B(n9991), .Z(n10081) );
  XNOR U10332 ( .A(n10082), .B(n10081), .Z(n10083) );
  NANDN U10333 ( .A(n9994), .B(n9993), .Z(n9998) );
  NANDN U10334 ( .A(n9996), .B(n9995), .Z(n9997) );
  NAND U10335 ( .A(n9998), .B(n9997), .Z(n10084) );
  XNOR U10336 ( .A(n10083), .B(n10084), .Z(n10029) );
  XOR U10337 ( .A(n10030), .B(n10029), .Z(n10088) );
  NANDN U10338 ( .A(n10000), .B(n9999), .Z(n10004) );
  NANDN U10339 ( .A(n10002), .B(n10001), .Z(n10003) );
  AND U10340 ( .A(n10004), .B(n10003), .Z(n10087) );
  XNOR U10341 ( .A(n10088), .B(n10087), .Z(n10089) );
  XOR U10342 ( .A(n10090), .B(n10089), .Z(n10022) );
  NANDN U10343 ( .A(n10006), .B(n10005), .Z(n10010) );
  NAND U10344 ( .A(n10008), .B(n10007), .Z(n10009) );
  AND U10345 ( .A(n10010), .B(n10009), .Z(n10021) );
  XNOR U10346 ( .A(n10022), .B(n10021), .Z(n10023) );
  XNOR U10347 ( .A(n10024), .B(n10023), .Z(n10016) );
  XNOR U10348 ( .A(sreg[377]), .B(n10016), .Z(n10018) );
  NANDN U10349 ( .A(sreg[376]), .B(n10011), .Z(n10015) );
  NAND U10350 ( .A(n10013), .B(n10012), .Z(n10014) );
  NAND U10351 ( .A(n10015), .B(n10014), .Z(n10017) );
  XNOR U10352 ( .A(n10018), .B(n10017), .Z(c[377]) );
  NANDN U10353 ( .A(sreg[377]), .B(n10016), .Z(n10020) );
  NAND U10354 ( .A(n10018), .B(n10017), .Z(n10019) );
  AND U10355 ( .A(n10020), .B(n10019), .Z(n10095) );
  NANDN U10356 ( .A(n10022), .B(n10021), .Z(n10026) );
  NANDN U10357 ( .A(n10024), .B(n10023), .Z(n10025) );
  AND U10358 ( .A(n10026), .B(n10025), .Z(n10100) );
  NANDN U10359 ( .A(n10028), .B(n10027), .Z(n10032) );
  NAND U10360 ( .A(n10030), .B(n10029), .Z(n10031) );
  AND U10361 ( .A(n10032), .B(n10031), .Z(n10167) );
  NANDN U10362 ( .A(n10034), .B(n10033), .Z(n10038) );
  NANDN U10363 ( .A(n10036), .B(n10035), .Z(n10037) );
  AND U10364 ( .A(n10038), .B(n10037), .Z(n10133) );
  NAND U10365 ( .A(n19808), .B(n10039), .Z(n10041) );
  XOR U10366 ( .A(b[13]), .B(a[126]), .Z(n10119) );
  NAND U10367 ( .A(n19768), .B(n10119), .Z(n10040) );
  AND U10368 ( .A(n10041), .B(n10040), .Z(n10111) );
  AND U10369 ( .A(b[15]), .B(a[122]), .Z(n10110) );
  XNOR U10370 ( .A(n10111), .B(n10110), .Z(n10112) );
  NAND U10371 ( .A(b[0]), .B(a[138]), .Z(n10042) );
  XNOR U10372 ( .A(b[1]), .B(n10042), .Z(n10044) );
  NANDN U10373 ( .A(b[0]), .B(a[137]), .Z(n10043) );
  NAND U10374 ( .A(n10044), .B(n10043), .Z(n10113) );
  XNOR U10375 ( .A(n10112), .B(n10113), .Z(n10131) );
  NAND U10376 ( .A(n33), .B(n10045), .Z(n10047) );
  XOR U10377 ( .A(b[5]), .B(a[134]), .Z(n10122) );
  NAND U10378 ( .A(n19342), .B(n10122), .Z(n10046) );
  AND U10379 ( .A(n10047), .B(n10046), .Z(n10155) );
  NAND U10380 ( .A(n34), .B(n10048), .Z(n10050) );
  XOR U10381 ( .A(b[7]), .B(a[132]), .Z(n10125) );
  NAND U10382 ( .A(n19486), .B(n10125), .Z(n10049) );
  AND U10383 ( .A(n10050), .B(n10049), .Z(n10153) );
  NAND U10384 ( .A(n31), .B(n10051), .Z(n10053) );
  XOR U10385 ( .A(b[3]), .B(a[136]), .Z(n10128) );
  NAND U10386 ( .A(n32), .B(n10128), .Z(n10052) );
  NAND U10387 ( .A(n10053), .B(n10052), .Z(n10152) );
  XNOR U10388 ( .A(n10153), .B(n10152), .Z(n10154) );
  XOR U10389 ( .A(n10155), .B(n10154), .Z(n10132) );
  XOR U10390 ( .A(n10131), .B(n10132), .Z(n10134) );
  XOR U10391 ( .A(n10133), .B(n10134), .Z(n10105) );
  NANDN U10392 ( .A(n10055), .B(n10054), .Z(n10059) );
  OR U10393 ( .A(n10057), .B(n10056), .Z(n10058) );
  AND U10394 ( .A(n10059), .B(n10058), .Z(n10104) );
  XNOR U10395 ( .A(n10105), .B(n10104), .Z(n10107) );
  NAND U10396 ( .A(n10060), .B(n19724), .Z(n10062) );
  XOR U10397 ( .A(b[11]), .B(a[128]), .Z(n10137) );
  NAND U10398 ( .A(n19692), .B(n10137), .Z(n10061) );
  AND U10399 ( .A(n10062), .B(n10061), .Z(n10148) );
  NAND U10400 ( .A(n19838), .B(n10063), .Z(n10065) );
  XOR U10401 ( .A(b[15]), .B(a[124]), .Z(n10140) );
  NAND U10402 ( .A(n19805), .B(n10140), .Z(n10064) );
  AND U10403 ( .A(n10065), .B(n10064), .Z(n10147) );
  NAND U10404 ( .A(n35), .B(n10066), .Z(n10068) );
  XOR U10405 ( .A(b[9]), .B(a[130]), .Z(n10143) );
  NAND U10406 ( .A(n19598), .B(n10143), .Z(n10067) );
  NAND U10407 ( .A(n10068), .B(n10067), .Z(n10146) );
  XOR U10408 ( .A(n10147), .B(n10146), .Z(n10149) );
  XOR U10409 ( .A(n10148), .B(n10149), .Z(n10159) );
  NANDN U10410 ( .A(n10070), .B(n10069), .Z(n10074) );
  OR U10411 ( .A(n10072), .B(n10071), .Z(n10073) );
  AND U10412 ( .A(n10074), .B(n10073), .Z(n10158) );
  XNOR U10413 ( .A(n10159), .B(n10158), .Z(n10160) );
  NANDN U10414 ( .A(n10076), .B(n10075), .Z(n10080) );
  NANDN U10415 ( .A(n10078), .B(n10077), .Z(n10079) );
  NAND U10416 ( .A(n10080), .B(n10079), .Z(n10161) );
  XNOR U10417 ( .A(n10160), .B(n10161), .Z(n10106) );
  XOR U10418 ( .A(n10107), .B(n10106), .Z(n10165) );
  NANDN U10419 ( .A(n10082), .B(n10081), .Z(n10086) );
  NANDN U10420 ( .A(n10084), .B(n10083), .Z(n10085) );
  AND U10421 ( .A(n10086), .B(n10085), .Z(n10164) );
  XNOR U10422 ( .A(n10165), .B(n10164), .Z(n10166) );
  XOR U10423 ( .A(n10167), .B(n10166), .Z(n10099) );
  NANDN U10424 ( .A(n10088), .B(n10087), .Z(n10092) );
  NAND U10425 ( .A(n10090), .B(n10089), .Z(n10091) );
  AND U10426 ( .A(n10092), .B(n10091), .Z(n10098) );
  XOR U10427 ( .A(n10099), .B(n10098), .Z(n10101) );
  XOR U10428 ( .A(n10100), .B(n10101), .Z(n10093) );
  XNOR U10429 ( .A(n10093), .B(sreg[378]), .Z(n10094) );
  XOR U10430 ( .A(n10095), .B(n10094), .Z(c[378]) );
  NANDN U10431 ( .A(n10093), .B(sreg[378]), .Z(n10097) );
  NAND U10432 ( .A(n10095), .B(n10094), .Z(n10096) );
  AND U10433 ( .A(n10097), .B(n10096), .Z(n10244) );
  NANDN U10434 ( .A(n10099), .B(n10098), .Z(n10103) );
  OR U10435 ( .A(n10101), .B(n10100), .Z(n10102) );
  AND U10436 ( .A(n10103), .B(n10102), .Z(n10173) );
  NANDN U10437 ( .A(n10105), .B(n10104), .Z(n10109) );
  NAND U10438 ( .A(n10107), .B(n10106), .Z(n10108) );
  AND U10439 ( .A(n10109), .B(n10108), .Z(n10239) );
  NANDN U10440 ( .A(n10111), .B(n10110), .Z(n10115) );
  NANDN U10441 ( .A(n10113), .B(n10112), .Z(n10114) );
  AND U10442 ( .A(n10115), .B(n10114), .Z(n10226) );
  NAND U10443 ( .A(b[0]), .B(a[139]), .Z(n10116) );
  XNOR U10444 ( .A(b[1]), .B(n10116), .Z(n10118) );
  NANDN U10445 ( .A(b[0]), .B(a[138]), .Z(n10117) );
  NAND U10446 ( .A(n10118), .B(n10117), .Z(n10206) );
  NAND U10447 ( .A(n19808), .B(n10119), .Z(n10121) );
  XOR U10448 ( .A(b[13]), .B(a[127]), .Z(n10212) );
  NAND U10449 ( .A(n19768), .B(n10212), .Z(n10120) );
  AND U10450 ( .A(n10121), .B(n10120), .Z(n10204) );
  AND U10451 ( .A(b[15]), .B(a[123]), .Z(n10203) );
  XNOR U10452 ( .A(n10204), .B(n10203), .Z(n10205) );
  XNOR U10453 ( .A(n10206), .B(n10205), .Z(n10224) );
  NAND U10454 ( .A(n33), .B(n10122), .Z(n10124) );
  XOR U10455 ( .A(b[5]), .B(a[135]), .Z(n10215) );
  NAND U10456 ( .A(n19342), .B(n10215), .Z(n10123) );
  AND U10457 ( .A(n10124), .B(n10123), .Z(n10200) );
  NAND U10458 ( .A(n34), .B(n10125), .Z(n10127) );
  XOR U10459 ( .A(b[7]), .B(a[133]), .Z(n10218) );
  NAND U10460 ( .A(n19486), .B(n10218), .Z(n10126) );
  AND U10461 ( .A(n10127), .B(n10126), .Z(n10198) );
  NAND U10462 ( .A(n31), .B(n10128), .Z(n10130) );
  XOR U10463 ( .A(b[3]), .B(a[137]), .Z(n10221) );
  NAND U10464 ( .A(n32), .B(n10221), .Z(n10129) );
  NAND U10465 ( .A(n10130), .B(n10129), .Z(n10197) );
  XNOR U10466 ( .A(n10198), .B(n10197), .Z(n10199) );
  XOR U10467 ( .A(n10200), .B(n10199), .Z(n10225) );
  XOR U10468 ( .A(n10224), .B(n10225), .Z(n10227) );
  XOR U10469 ( .A(n10226), .B(n10227), .Z(n10177) );
  NANDN U10470 ( .A(n10132), .B(n10131), .Z(n10136) );
  OR U10471 ( .A(n10134), .B(n10133), .Z(n10135) );
  AND U10472 ( .A(n10136), .B(n10135), .Z(n10176) );
  XNOR U10473 ( .A(n10177), .B(n10176), .Z(n10179) );
  NAND U10474 ( .A(n10137), .B(n19724), .Z(n10139) );
  XOR U10475 ( .A(b[11]), .B(a[129]), .Z(n10182) );
  NAND U10476 ( .A(n19692), .B(n10182), .Z(n10138) );
  AND U10477 ( .A(n10139), .B(n10138), .Z(n10193) );
  NAND U10478 ( .A(n19838), .B(n10140), .Z(n10142) );
  XOR U10479 ( .A(b[15]), .B(a[125]), .Z(n10185) );
  NAND U10480 ( .A(n19805), .B(n10185), .Z(n10141) );
  AND U10481 ( .A(n10142), .B(n10141), .Z(n10192) );
  NAND U10482 ( .A(n35), .B(n10143), .Z(n10145) );
  XOR U10483 ( .A(b[9]), .B(a[131]), .Z(n10188) );
  NAND U10484 ( .A(n19598), .B(n10188), .Z(n10144) );
  NAND U10485 ( .A(n10145), .B(n10144), .Z(n10191) );
  XOR U10486 ( .A(n10192), .B(n10191), .Z(n10194) );
  XOR U10487 ( .A(n10193), .B(n10194), .Z(n10231) );
  NANDN U10488 ( .A(n10147), .B(n10146), .Z(n10151) );
  OR U10489 ( .A(n10149), .B(n10148), .Z(n10150) );
  AND U10490 ( .A(n10151), .B(n10150), .Z(n10230) );
  XNOR U10491 ( .A(n10231), .B(n10230), .Z(n10232) );
  NANDN U10492 ( .A(n10153), .B(n10152), .Z(n10157) );
  NANDN U10493 ( .A(n10155), .B(n10154), .Z(n10156) );
  NAND U10494 ( .A(n10157), .B(n10156), .Z(n10233) );
  XNOR U10495 ( .A(n10232), .B(n10233), .Z(n10178) );
  XOR U10496 ( .A(n10179), .B(n10178), .Z(n10237) );
  NANDN U10497 ( .A(n10159), .B(n10158), .Z(n10163) );
  NANDN U10498 ( .A(n10161), .B(n10160), .Z(n10162) );
  AND U10499 ( .A(n10163), .B(n10162), .Z(n10236) );
  XNOR U10500 ( .A(n10237), .B(n10236), .Z(n10238) );
  XOR U10501 ( .A(n10239), .B(n10238), .Z(n10171) );
  NANDN U10502 ( .A(n10165), .B(n10164), .Z(n10169) );
  NAND U10503 ( .A(n10167), .B(n10166), .Z(n10168) );
  AND U10504 ( .A(n10169), .B(n10168), .Z(n10170) );
  XNOR U10505 ( .A(n10171), .B(n10170), .Z(n10172) );
  XNOR U10506 ( .A(n10173), .B(n10172), .Z(n10242) );
  XNOR U10507 ( .A(sreg[379]), .B(n10242), .Z(n10243) );
  XNOR U10508 ( .A(n10244), .B(n10243), .Z(c[379]) );
  NANDN U10509 ( .A(n10171), .B(n10170), .Z(n10175) );
  NANDN U10510 ( .A(n10173), .B(n10172), .Z(n10174) );
  AND U10511 ( .A(n10175), .B(n10174), .Z(n10250) );
  NANDN U10512 ( .A(n10177), .B(n10176), .Z(n10181) );
  NAND U10513 ( .A(n10179), .B(n10178), .Z(n10180) );
  AND U10514 ( .A(n10181), .B(n10180), .Z(n10316) );
  NAND U10515 ( .A(n10182), .B(n19724), .Z(n10184) );
  XOR U10516 ( .A(b[11]), .B(a[130]), .Z(n10286) );
  NAND U10517 ( .A(n19692), .B(n10286), .Z(n10183) );
  AND U10518 ( .A(n10184), .B(n10183), .Z(n10297) );
  NAND U10519 ( .A(n19838), .B(n10185), .Z(n10187) );
  XOR U10520 ( .A(b[15]), .B(a[126]), .Z(n10289) );
  NAND U10521 ( .A(n19805), .B(n10289), .Z(n10186) );
  AND U10522 ( .A(n10187), .B(n10186), .Z(n10296) );
  NAND U10523 ( .A(n35), .B(n10188), .Z(n10190) );
  XOR U10524 ( .A(b[9]), .B(a[132]), .Z(n10292) );
  NAND U10525 ( .A(n19598), .B(n10292), .Z(n10189) );
  NAND U10526 ( .A(n10190), .B(n10189), .Z(n10295) );
  XOR U10527 ( .A(n10296), .B(n10295), .Z(n10298) );
  XOR U10528 ( .A(n10297), .B(n10298), .Z(n10308) );
  NANDN U10529 ( .A(n10192), .B(n10191), .Z(n10196) );
  OR U10530 ( .A(n10194), .B(n10193), .Z(n10195) );
  AND U10531 ( .A(n10196), .B(n10195), .Z(n10307) );
  XNOR U10532 ( .A(n10308), .B(n10307), .Z(n10309) );
  NANDN U10533 ( .A(n10198), .B(n10197), .Z(n10202) );
  NANDN U10534 ( .A(n10200), .B(n10199), .Z(n10201) );
  NAND U10535 ( .A(n10202), .B(n10201), .Z(n10310) );
  XNOR U10536 ( .A(n10309), .B(n10310), .Z(n10256) );
  NANDN U10537 ( .A(n10204), .B(n10203), .Z(n10208) );
  NANDN U10538 ( .A(n10206), .B(n10205), .Z(n10207) );
  AND U10539 ( .A(n10208), .B(n10207), .Z(n10282) );
  NAND U10540 ( .A(b[0]), .B(a[140]), .Z(n10209) );
  XNOR U10541 ( .A(b[1]), .B(n10209), .Z(n10211) );
  NANDN U10542 ( .A(b[0]), .B(a[139]), .Z(n10210) );
  NAND U10543 ( .A(n10211), .B(n10210), .Z(n10262) );
  NAND U10544 ( .A(n19808), .B(n10212), .Z(n10214) );
  XOR U10545 ( .A(b[13]), .B(a[128]), .Z(n10268) );
  NAND U10546 ( .A(n19768), .B(n10268), .Z(n10213) );
  AND U10547 ( .A(n10214), .B(n10213), .Z(n10260) );
  AND U10548 ( .A(b[15]), .B(a[124]), .Z(n10259) );
  XNOR U10549 ( .A(n10260), .B(n10259), .Z(n10261) );
  XNOR U10550 ( .A(n10262), .B(n10261), .Z(n10280) );
  NAND U10551 ( .A(n33), .B(n10215), .Z(n10217) );
  XOR U10552 ( .A(b[5]), .B(a[136]), .Z(n10271) );
  NAND U10553 ( .A(n19342), .B(n10271), .Z(n10216) );
  AND U10554 ( .A(n10217), .B(n10216), .Z(n10304) );
  NAND U10555 ( .A(n34), .B(n10218), .Z(n10220) );
  XOR U10556 ( .A(b[7]), .B(a[134]), .Z(n10274) );
  NAND U10557 ( .A(n19486), .B(n10274), .Z(n10219) );
  AND U10558 ( .A(n10220), .B(n10219), .Z(n10302) );
  NAND U10559 ( .A(n31), .B(n10221), .Z(n10223) );
  XOR U10560 ( .A(b[3]), .B(a[138]), .Z(n10277) );
  NAND U10561 ( .A(n32), .B(n10277), .Z(n10222) );
  NAND U10562 ( .A(n10223), .B(n10222), .Z(n10301) );
  XNOR U10563 ( .A(n10302), .B(n10301), .Z(n10303) );
  XOR U10564 ( .A(n10304), .B(n10303), .Z(n10281) );
  XOR U10565 ( .A(n10280), .B(n10281), .Z(n10283) );
  XOR U10566 ( .A(n10282), .B(n10283), .Z(n10254) );
  NANDN U10567 ( .A(n10225), .B(n10224), .Z(n10229) );
  OR U10568 ( .A(n10227), .B(n10226), .Z(n10228) );
  AND U10569 ( .A(n10229), .B(n10228), .Z(n10253) );
  XNOR U10570 ( .A(n10254), .B(n10253), .Z(n10255) );
  XOR U10571 ( .A(n10256), .B(n10255), .Z(n10314) );
  NANDN U10572 ( .A(n10231), .B(n10230), .Z(n10235) );
  NANDN U10573 ( .A(n10233), .B(n10232), .Z(n10234) );
  AND U10574 ( .A(n10235), .B(n10234), .Z(n10313) );
  XNOR U10575 ( .A(n10314), .B(n10313), .Z(n10315) );
  XOR U10576 ( .A(n10316), .B(n10315), .Z(n10248) );
  NANDN U10577 ( .A(n10237), .B(n10236), .Z(n10241) );
  NAND U10578 ( .A(n10239), .B(n10238), .Z(n10240) );
  AND U10579 ( .A(n10241), .B(n10240), .Z(n10247) );
  XNOR U10580 ( .A(n10248), .B(n10247), .Z(n10249) );
  XNOR U10581 ( .A(n10250), .B(n10249), .Z(n10319) );
  XNOR U10582 ( .A(sreg[380]), .B(n10319), .Z(n10321) );
  NANDN U10583 ( .A(sreg[379]), .B(n10242), .Z(n10246) );
  NAND U10584 ( .A(n10244), .B(n10243), .Z(n10245) );
  NAND U10585 ( .A(n10246), .B(n10245), .Z(n10320) );
  XNOR U10586 ( .A(n10321), .B(n10320), .Z(c[380]) );
  NANDN U10587 ( .A(n10248), .B(n10247), .Z(n10252) );
  NANDN U10588 ( .A(n10250), .B(n10249), .Z(n10251) );
  AND U10589 ( .A(n10252), .B(n10251), .Z(n10331) );
  NANDN U10590 ( .A(n10254), .B(n10253), .Z(n10258) );
  NAND U10591 ( .A(n10256), .B(n10255), .Z(n10257) );
  AND U10592 ( .A(n10258), .B(n10257), .Z(n10398) );
  NANDN U10593 ( .A(n10260), .B(n10259), .Z(n10264) );
  NANDN U10594 ( .A(n10262), .B(n10261), .Z(n10263) );
  AND U10595 ( .A(n10264), .B(n10263), .Z(n10364) );
  NAND U10596 ( .A(b[0]), .B(a[141]), .Z(n10265) );
  XNOR U10597 ( .A(b[1]), .B(n10265), .Z(n10267) );
  NANDN U10598 ( .A(b[0]), .B(a[140]), .Z(n10266) );
  NAND U10599 ( .A(n10267), .B(n10266), .Z(n10344) );
  NAND U10600 ( .A(n19808), .B(n10268), .Z(n10270) );
  XOR U10601 ( .A(b[13]), .B(a[129]), .Z(n10347) );
  NAND U10602 ( .A(n19768), .B(n10347), .Z(n10269) );
  AND U10603 ( .A(n10270), .B(n10269), .Z(n10342) );
  AND U10604 ( .A(b[15]), .B(a[125]), .Z(n10341) );
  XNOR U10605 ( .A(n10342), .B(n10341), .Z(n10343) );
  XNOR U10606 ( .A(n10344), .B(n10343), .Z(n10362) );
  NAND U10607 ( .A(n33), .B(n10271), .Z(n10273) );
  XOR U10608 ( .A(b[5]), .B(a[137]), .Z(n10353) );
  NAND U10609 ( .A(n19342), .B(n10353), .Z(n10272) );
  AND U10610 ( .A(n10273), .B(n10272), .Z(n10386) );
  NAND U10611 ( .A(n34), .B(n10274), .Z(n10276) );
  XOR U10612 ( .A(b[7]), .B(a[135]), .Z(n10356) );
  NAND U10613 ( .A(n19486), .B(n10356), .Z(n10275) );
  AND U10614 ( .A(n10276), .B(n10275), .Z(n10384) );
  NAND U10615 ( .A(n31), .B(n10277), .Z(n10279) );
  XOR U10616 ( .A(b[3]), .B(a[139]), .Z(n10359) );
  NAND U10617 ( .A(n32), .B(n10359), .Z(n10278) );
  NAND U10618 ( .A(n10279), .B(n10278), .Z(n10383) );
  XNOR U10619 ( .A(n10384), .B(n10383), .Z(n10385) );
  XOR U10620 ( .A(n10386), .B(n10385), .Z(n10363) );
  XOR U10621 ( .A(n10362), .B(n10363), .Z(n10365) );
  XOR U10622 ( .A(n10364), .B(n10365), .Z(n10336) );
  NANDN U10623 ( .A(n10281), .B(n10280), .Z(n10285) );
  OR U10624 ( .A(n10283), .B(n10282), .Z(n10284) );
  AND U10625 ( .A(n10285), .B(n10284), .Z(n10335) );
  XNOR U10626 ( .A(n10336), .B(n10335), .Z(n10338) );
  NAND U10627 ( .A(n10286), .B(n19724), .Z(n10288) );
  XOR U10628 ( .A(b[11]), .B(a[131]), .Z(n10368) );
  NAND U10629 ( .A(n19692), .B(n10368), .Z(n10287) );
  AND U10630 ( .A(n10288), .B(n10287), .Z(n10379) );
  NAND U10631 ( .A(n19838), .B(n10289), .Z(n10291) );
  XOR U10632 ( .A(b[15]), .B(a[127]), .Z(n10371) );
  NAND U10633 ( .A(n19805), .B(n10371), .Z(n10290) );
  AND U10634 ( .A(n10291), .B(n10290), .Z(n10378) );
  NAND U10635 ( .A(n35), .B(n10292), .Z(n10294) );
  XOR U10636 ( .A(b[9]), .B(a[133]), .Z(n10374) );
  NAND U10637 ( .A(n19598), .B(n10374), .Z(n10293) );
  NAND U10638 ( .A(n10294), .B(n10293), .Z(n10377) );
  XOR U10639 ( .A(n10378), .B(n10377), .Z(n10380) );
  XOR U10640 ( .A(n10379), .B(n10380), .Z(n10390) );
  NANDN U10641 ( .A(n10296), .B(n10295), .Z(n10300) );
  OR U10642 ( .A(n10298), .B(n10297), .Z(n10299) );
  AND U10643 ( .A(n10300), .B(n10299), .Z(n10389) );
  XNOR U10644 ( .A(n10390), .B(n10389), .Z(n10391) );
  NANDN U10645 ( .A(n10302), .B(n10301), .Z(n10306) );
  NANDN U10646 ( .A(n10304), .B(n10303), .Z(n10305) );
  NAND U10647 ( .A(n10306), .B(n10305), .Z(n10392) );
  XNOR U10648 ( .A(n10391), .B(n10392), .Z(n10337) );
  XOR U10649 ( .A(n10338), .B(n10337), .Z(n10396) );
  NANDN U10650 ( .A(n10308), .B(n10307), .Z(n10312) );
  NANDN U10651 ( .A(n10310), .B(n10309), .Z(n10311) );
  AND U10652 ( .A(n10312), .B(n10311), .Z(n10395) );
  XNOR U10653 ( .A(n10396), .B(n10395), .Z(n10397) );
  XOR U10654 ( .A(n10398), .B(n10397), .Z(n10330) );
  NANDN U10655 ( .A(n10314), .B(n10313), .Z(n10318) );
  NAND U10656 ( .A(n10316), .B(n10315), .Z(n10317) );
  AND U10657 ( .A(n10318), .B(n10317), .Z(n10329) );
  XOR U10658 ( .A(n10330), .B(n10329), .Z(n10332) );
  XOR U10659 ( .A(n10331), .B(n10332), .Z(n10324) );
  XNOR U10660 ( .A(n10324), .B(sreg[381]), .Z(n10326) );
  NANDN U10661 ( .A(sreg[380]), .B(n10319), .Z(n10323) );
  NAND U10662 ( .A(n10321), .B(n10320), .Z(n10322) );
  AND U10663 ( .A(n10323), .B(n10322), .Z(n10325) );
  XOR U10664 ( .A(n10326), .B(n10325), .Z(c[381]) );
  NANDN U10665 ( .A(n10324), .B(sreg[381]), .Z(n10328) );
  NAND U10666 ( .A(n10326), .B(n10325), .Z(n10327) );
  AND U10667 ( .A(n10328), .B(n10327), .Z(n10475) );
  NANDN U10668 ( .A(n10330), .B(n10329), .Z(n10334) );
  OR U10669 ( .A(n10332), .B(n10331), .Z(n10333) );
  AND U10670 ( .A(n10334), .B(n10333), .Z(n10404) );
  NANDN U10671 ( .A(n10336), .B(n10335), .Z(n10340) );
  NAND U10672 ( .A(n10338), .B(n10337), .Z(n10339) );
  AND U10673 ( .A(n10340), .B(n10339), .Z(n10470) );
  NANDN U10674 ( .A(n10342), .B(n10341), .Z(n10346) );
  NANDN U10675 ( .A(n10344), .B(n10343), .Z(n10345) );
  AND U10676 ( .A(n10346), .B(n10345), .Z(n10436) );
  NAND U10677 ( .A(n19808), .B(n10347), .Z(n10349) );
  XOR U10678 ( .A(b[13]), .B(a[130]), .Z(n10422) );
  NAND U10679 ( .A(n19768), .B(n10422), .Z(n10348) );
  AND U10680 ( .A(n10349), .B(n10348), .Z(n10414) );
  AND U10681 ( .A(b[15]), .B(a[126]), .Z(n10413) );
  XNOR U10682 ( .A(n10414), .B(n10413), .Z(n10415) );
  NAND U10683 ( .A(b[0]), .B(a[142]), .Z(n10350) );
  XNOR U10684 ( .A(b[1]), .B(n10350), .Z(n10352) );
  NANDN U10685 ( .A(b[0]), .B(a[141]), .Z(n10351) );
  NAND U10686 ( .A(n10352), .B(n10351), .Z(n10416) );
  XNOR U10687 ( .A(n10415), .B(n10416), .Z(n10434) );
  NAND U10688 ( .A(n33), .B(n10353), .Z(n10355) );
  XOR U10689 ( .A(b[5]), .B(a[138]), .Z(n10425) );
  NAND U10690 ( .A(n19342), .B(n10425), .Z(n10354) );
  AND U10691 ( .A(n10355), .B(n10354), .Z(n10458) );
  NAND U10692 ( .A(n34), .B(n10356), .Z(n10358) );
  XOR U10693 ( .A(b[7]), .B(a[136]), .Z(n10428) );
  NAND U10694 ( .A(n19486), .B(n10428), .Z(n10357) );
  AND U10695 ( .A(n10358), .B(n10357), .Z(n10456) );
  NAND U10696 ( .A(n31), .B(n10359), .Z(n10361) );
  XOR U10697 ( .A(b[3]), .B(a[140]), .Z(n10431) );
  NAND U10698 ( .A(n32), .B(n10431), .Z(n10360) );
  NAND U10699 ( .A(n10361), .B(n10360), .Z(n10455) );
  XNOR U10700 ( .A(n10456), .B(n10455), .Z(n10457) );
  XOR U10701 ( .A(n10458), .B(n10457), .Z(n10435) );
  XOR U10702 ( .A(n10434), .B(n10435), .Z(n10437) );
  XOR U10703 ( .A(n10436), .B(n10437), .Z(n10408) );
  NANDN U10704 ( .A(n10363), .B(n10362), .Z(n10367) );
  OR U10705 ( .A(n10365), .B(n10364), .Z(n10366) );
  AND U10706 ( .A(n10367), .B(n10366), .Z(n10407) );
  XNOR U10707 ( .A(n10408), .B(n10407), .Z(n10410) );
  NAND U10708 ( .A(n10368), .B(n19724), .Z(n10370) );
  XOR U10709 ( .A(b[11]), .B(a[132]), .Z(n10440) );
  NAND U10710 ( .A(n19692), .B(n10440), .Z(n10369) );
  AND U10711 ( .A(n10370), .B(n10369), .Z(n10451) );
  NAND U10712 ( .A(n19838), .B(n10371), .Z(n10373) );
  XOR U10713 ( .A(b[15]), .B(a[128]), .Z(n10443) );
  NAND U10714 ( .A(n19805), .B(n10443), .Z(n10372) );
  AND U10715 ( .A(n10373), .B(n10372), .Z(n10450) );
  NAND U10716 ( .A(n35), .B(n10374), .Z(n10376) );
  XOR U10717 ( .A(b[9]), .B(a[134]), .Z(n10446) );
  NAND U10718 ( .A(n19598), .B(n10446), .Z(n10375) );
  NAND U10719 ( .A(n10376), .B(n10375), .Z(n10449) );
  XOR U10720 ( .A(n10450), .B(n10449), .Z(n10452) );
  XOR U10721 ( .A(n10451), .B(n10452), .Z(n10462) );
  NANDN U10722 ( .A(n10378), .B(n10377), .Z(n10382) );
  OR U10723 ( .A(n10380), .B(n10379), .Z(n10381) );
  AND U10724 ( .A(n10382), .B(n10381), .Z(n10461) );
  XNOR U10725 ( .A(n10462), .B(n10461), .Z(n10463) );
  NANDN U10726 ( .A(n10384), .B(n10383), .Z(n10388) );
  NANDN U10727 ( .A(n10386), .B(n10385), .Z(n10387) );
  NAND U10728 ( .A(n10388), .B(n10387), .Z(n10464) );
  XNOR U10729 ( .A(n10463), .B(n10464), .Z(n10409) );
  XOR U10730 ( .A(n10410), .B(n10409), .Z(n10468) );
  NANDN U10731 ( .A(n10390), .B(n10389), .Z(n10394) );
  NANDN U10732 ( .A(n10392), .B(n10391), .Z(n10393) );
  AND U10733 ( .A(n10394), .B(n10393), .Z(n10467) );
  XNOR U10734 ( .A(n10468), .B(n10467), .Z(n10469) );
  XOR U10735 ( .A(n10470), .B(n10469), .Z(n10402) );
  NANDN U10736 ( .A(n10396), .B(n10395), .Z(n10400) );
  NAND U10737 ( .A(n10398), .B(n10397), .Z(n10399) );
  AND U10738 ( .A(n10400), .B(n10399), .Z(n10401) );
  XNOR U10739 ( .A(n10402), .B(n10401), .Z(n10403) );
  XNOR U10740 ( .A(n10404), .B(n10403), .Z(n10473) );
  XNOR U10741 ( .A(sreg[382]), .B(n10473), .Z(n10474) );
  XNOR U10742 ( .A(n10475), .B(n10474), .Z(c[382]) );
  NANDN U10743 ( .A(n10402), .B(n10401), .Z(n10406) );
  NANDN U10744 ( .A(n10404), .B(n10403), .Z(n10405) );
  AND U10745 ( .A(n10406), .B(n10405), .Z(n10481) );
  NANDN U10746 ( .A(n10408), .B(n10407), .Z(n10412) );
  NAND U10747 ( .A(n10410), .B(n10409), .Z(n10411) );
  AND U10748 ( .A(n10412), .B(n10411), .Z(n10547) );
  NANDN U10749 ( .A(n10414), .B(n10413), .Z(n10418) );
  NANDN U10750 ( .A(n10416), .B(n10415), .Z(n10417) );
  AND U10751 ( .A(n10418), .B(n10417), .Z(n10513) );
  NAND U10752 ( .A(b[0]), .B(a[143]), .Z(n10419) );
  XNOR U10753 ( .A(b[1]), .B(n10419), .Z(n10421) );
  NANDN U10754 ( .A(b[0]), .B(a[142]), .Z(n10420) );
  NAND U10755 ( .A(n10421), .B(n10420), .Z(n10493) );
  NAND U10756 ( .A(n19808), .B(n10422), .Z(n10424) );
  XOR U10757 ( .A(b[13]), .B(a[131]), .Z(n10499) );
  NAND U10758 ( .A(n19768), .B(n10499), .Z(n10423) );
  AND U10759 ( .A(n10424), .B(n10423), .Z(n10491) );
  AND U10760 ( .A(b[15]), .B(a[127]), .Z(n10490) );
  XNOR U10761 ( .A(n10491), .B(n10490), .Z(n10492) );
  XNOR U10762 ( .A(n10493), .B(n10492), .Z(n10511) );
  NAND U10763 ( .A(n33), .B(n10425), .Z(n10427) );
  XOR U10764 ( .A(b[5]), .B(a[139]), .Z(n10502) );
  NAND U10765 ( .A(n19342), .B(n10502), .Z(n10426) );
  AND U10766 ( .A(n10427), .B(n10426), .Z(n10535) );
  NAND U10767 ( .A(n34), .B(n10428), .Z(n10430) );
  XOR U10768 ( .A(b[7]), .B(a[137]), .Z(n10505) );
  NAND U10769 ( .A(n19486), .B(n10505), .Z(n10429) );
  AND U10770 ( .A(n10430), .B(n10429), .Z(n10533) );
  NAND U10771 ( .A(n31), .B(n10431), .Z(n10433) );
  XOR U10772 ( .A(b[3]), .B(a[141]), .Z(n10508) );
  NAND U10773 ( .A(n32), .B(n10508), .Z(n10432) );
  NAND U10774 ( .A(n10433), .B(n10432), .Z(n10532) );
  XNOR U10775 ( .A(n10533), .B(n10532), .Z(n10534) );
  XOR U10776 ( .A(n10535), .B(n10534), .Z(n10512) );
  XOR U10777 ( .A(n10511), .B(n10512), .Z(n10514) );
  XOR U10778 ( .A(n10513), .B(n10514), .Z(n10485) );
  NANDN U10779 ( .A(n10435), .B(n10434), .Z(n10439) );
  OR U10780 ( .A(n10437), .B(n10436), .Z(n10438) );
  AND U10781 ( .A(n10439), .B(n10438), .Z(n10484) );
  XNOR U10782 ( .A(n10485), .B(n10484), .Z(n10487) );
  NAND U10783 ( .A(n10440), .B(n19724), .Z(n10442) );
  XOR U10784 ( .A(b[11]), .B(a[133]), .Z(n10517) );
  NAND U10785 ( .A(n19692), .B(n10517), .Z(n10441) );
  AND U10786 ( .A(n10442), .B(n10441), .Z(n10528) );
  NAND U10787 ( .A(n19838), .B(n10443), .Z(n10445) );
  XOR U10788 ( .A(b[15]), .B(a[129]), .Z(n10520) );
  NAND U10789 ( .A(n19805), .B(n10520), .Z(n10444) );
  AND U10790 ( .A(n10445), .B(n10444), .Z(n10527) );
  NAND U10791 ( .A(n35), .B(n10446), .Z(n10448) );
  XOR U10792 ( .A(b[9]), .B(a[135]), .Z(n10523) );
  NAND U10793 ( .A(n19598), .B(n10523), .Z(n10447) );
  NAND U10794 ( .A(n10448), .B(n10447), .Z(n10526) );
  XOR U10795 ( .A(n10527), .B(n10526), .Z(n10529) );
  XOR U10796 ( .A(n10528), .B(n10529), .Z(n10539) );
  NANDN U10797 ( .A(n10450), .B(n10449), .Z(n10454) );
  OR U10798 ( .A(n10452), .B(n10451), .Z(n10453) );
  AND U10799 ( .A(n10454), .B(n10453), .Z(n10538) );
  XNOR U10800 ( .A(n10539), .B(n10538), .Z(n10540) );
  NANDN U10801 ( .A(n10456), .B(n10455), .Z(n10460) );
  NANDN U10802 ( .A(n10458), .B(n10457), .Z(n10459) );
  NAND U10803 ( .A(n10460), .B(n10459), .Z(n10541) );
  XNOR U10804 ( .A(n10540), .B(n10541), .Z(n10486) );
  XOR U10805 ( .A(n10487), .B(n10486), .Z(n10545) );
  NANDN U10806 ( .A(n10462), .B(n10461), .Z(n10466) );
  NANDN U10807 ( .A(n10464), .B(n10463), .Z(n10465) );
  AND U10808 ( .A(n10466), .B(n10465), .Z(n10544) );
  XNOR U10809 ( .A(n10545), .B(n10544), .Z(n10546) );
  XOR U10810 ( .A(n10547), .B(n10546), .Z(n10479) );
  NANDN U10811 ( .A(n10468), .B(n10467), .Z(n10472) );
  NAND U10812 ( .A(n10470), .B(n10469), .Z(n10471) );
  AND U10813 ( .A(n10472), .B(n10471), .Z(n10478) );
  XNOR U10814 ( .A(n10479), .B(n10478), .Z(n10480) );
  XNOR U10815 ( .A(n10481), .B(n10480), .Z(n10550) );
  XNOR U10816 ( .A(sreg[383]), .B(n10550), .Z(n10552) );
  NANDN U10817 ( .A(sreg[382]), .B(n10473), .Z(n10477) );
  NAND U10818 ( .A(n10475), .B(n10474), .Z(n10476) );
  NAND U10819 ( .A(n10477), .B(n10476), .Z(n10551) );
  XNOR U10820 ( .A(n10552), .B(n10551), .Z(c[383]) );
  NANDN U10821 ( .A(n10479), .B(n10478), .Z(n10483) );
  NANDN U10822 ( .A(n10481), .B(n10480), .Z(n10482) );
  AND U10823 ( .A(n10483), .B(n10482), .Z(n10558) );
  NANDN U10824 ( .A(n10485), .B(n10484), .Z(n10489) );
  NAND U10825 ( .A(n10487), .B(n10486), .Z(n10488) );
  AND U10826 ( .A(n10489), .B(n10488), .Z(n10624) );
  NANDN U10827 ( .A(n10491), .B(n10490), .Z(n10495) );
  NANDN U10828 ( .A(n10493), .B(n10492), .Z(n10494) );
  AND U10829 ( .A(n10495), .B(n10494), .Z(n10590) );
  NAND U10830 ( .A(b[0]), .B(a[144]), .Z(n10496) );
  XNOR U10831 ( .A(b[1]), .B(n10496), .Z(n10498) );
  NANDN U10832 ( .A(b[0]), .B(a[143]), .Z(n10497) );
  NAND U10833 ( .A(n10498), .B(n10497), .Z(n10570) );
  NAND U10834 ( .A(n19808), .B(n10499), .Z(n10501) );
  XOR U10835 ( .A(b[13]), .B(a[132]), .Z(n10576) );
  NAND U10836 ( .A(n19768), .B(n10576), .Z(n10500) );
  AND U10837 ( .A(n10501), .B(n10500), .Z(n10568) );
  AND U10838 ( .A(b[15]), .B(a[128]), .Z(n10567) );
  XNOR U10839 ( .A(n10568), .B(n10567), .Z(n10569) );
  XNOR U10840 ( .A(n10570), .B(n10569), .Z(n10588) );
  NAND U10841 ( .A(n33), .B(n10502), .Z(n10504) );
  XOR U10842 ( .A(b[5]), .B(a[140]), .Z(n10579) );
  NAND U10843 ( .A(n19342), .B(n10579), .Z(n10503) );
  AND U10844 ( .A(n10504), .B(n10503), .Z(n10612) );
  NAND U10845 ( .A(n34), .B(n10505), .Z(n10507) );
  XOR U10846 ( .A(b[7]), .B(a[138]), .Z(n10582) );
  NAND U10847 ( .A(n19486), .B(n10582), .Z(n10506) );
  AND U10848 ( .A(n10507), .B(n10506), .Z(n10610) );
  NAND U10849 ( .A(n31), .B(n10508), .Z(n10510) );
  XOR U10850 ( .A(b[3]), .B(a[142]), .Z(n10585) );
  NAND U10851 ( .A(n32), .B(n10585), .Z(n10509) );
  NAND U10852 ( .A(n10510), .B(n10509), .Z(n10609) );
  XNOR U10853 ( .A(n10610), .B(n10609), .Z(n10611) );
  XOR U10854 ( .A(n10612), .B(n10611), .Z(n10589) );
  XOR U10855 ( .A(n10588), .B(n10589), .Z(n10591) );
  XOR U10856 ( .A(n10590), .B(n10591), .Z(n10562) );
  NANDN U10857 ( .A(n10512), .B(n10511), .Z(n10516) );
  OR U10858 ( .A(n10514), .B(n10513), .Z(n10515) );
  AND U10859 ( .A(n10516), .B(n10515), .Z(n10561) );
  XNOR U10860 ( .A(n10562), .B(n10561), .Z(n10564) );
  NAND U10861 ( .A(n10517), .B(n19724), .Z(n10519) );
  XOR U10862 ( .A(b[11]), .B(a[134]), .Z(n10594) );
  NAND U10863 ( .A(n19692), .B(n10594), .Z(n10518) );
  AND U10864 ( .A(n10519), .B(n10518), .Z(n10605) );
  NAND U10865 ( .A(n19838), .B(n10520), .Z(n10522) );
  XOR U10866 ( .A(b[15]), .B(a[130]), .Z(n10597) );
  NAND U10867 ( .A(n19805), .B(n10597), .Z(n10521) );
  AND U10868 ( .A(n10522), .B(n10521), .Z(n10604) );
  NAND U10869 ( .A(n35), .B(n10523), .Z(n10525) );
  XOR U10870 ( .A(b[9]), .B(a[136]), .Z(n10600) );
  NAND U10871 ( .A(n19598), .B(n10600), .Z(n10524) );
  NAND U10872 ( .A(n10525), .B(n10524), .Z(n10603) );
  XOR U10873 ( .A(n10604), .B(n10603), .Z(n10606) );
  XOR U10874 ( .A(n10605), .B(n10606), .Z(n10616) );
  NANDN U10875 ( .A(n10527), .B(n10526), .Z(n10531) );
  OR U10876 ( .A(n10529), .B(n10528), .Z(n10530) );
  AND U10877 ( .A(n10531), .B(n10530), .Z(n10615) );
  XNOR U10878 ( .A(n10616), .B(n10615), .Z(n10617) );
  NANDN U10879 ( .A(n10533), .B(n10532), .Z(n10537) );
  NANDN U10880 ( .A(n10535), .B(n10534), .Z(n10536) );
  NAND U10881 ( .A(n10537), .B(n10536), .Z(n10618) );
  XNOR U10882 ( .A(n10617), .B(n10618), .Z(n10563) );
  XOR U10883 ( .A(n10564), .B(n10563), .Z(n10622) );
  NANDN U10884 ( .A(n10539), .B(n10538), .Z(n10543) );
  NANDN U10885 ( .A(n10541), .B(n10540), .Z(n10542) );
  AND U10886 ( .A(n10543), .B(n10542), .Z(n10621) );
  XNOR U10887 ( .A(n10622), .B(n10621), .Z(n10623) );
  XOR U10888 ( .A(n10624), .B(n10623), .Z(n10556) );
  NANDN U10889 ( .A(n10545), .B(n10544), .Z(n10549) );
  NAND U10890 ( .A(n10547), .B(n10546), .Z(n10548) );
  AND U10891 ( .A(n10549), .B(n10548), .Z(n10555) );
  XNOR U10892 ( .A(n10556), .B(n10555), .Z(n10557) );
  XNOR U10893 ( .A(n10558), .B(n10557), .Z(n10627) );
  XNOR U10894 ( .A(sreg[384]), .B(n10627), .Z(n10629) );
  NANDN U10895 ( .A(sreg[383]), .B(n10550), .Z(n10554) );
  NAND U10896 ( .A(n10552), .B(n10551), .Z(n10553) );
  NAND U10897 ( .A(n10554), .B(n10553), .Z(n10628) );
  XNOR U10898 ( .A(n10629), .B(n10628), .Z(c[384]) );
  NANDN U10899 ( .A(n10556), .B(n10555), .Z(n10560) );
  NANDN U10900 ( .A(n10558), .B(n10557), .Z(n10559) );
  AND U10901 ( .A(n10560), .B(n10559), .Z(n10635) );
  NANDN U10902 ( .A(n10562), .B(n10561), .Z(n10566) );
  NAND U10903 ( .A(n10564), .B(n10563), .Z(n10565) );
  AND U10904 ( .A(n10566), .B(n10565), .Z(n10701) );
  NANDN U10905 ( .A(n10568), .B(n10567), .Z(n10572) );
  NANDN U10906 ( .A(n10570), .B(n10569), .Z(n10571) );
  AND U10907 ( .A(n10572), .B(n10571), .Z(n10667) );
  NAND U10908 ( .A(b[0]), .B(a[145]), .Z(n10573) );
  XNOR U10909 ( .A(b[1]), .B(n10573), .Z(n10575) );
  NANDN U10910 ( .A(b[0]), .B(a[144]), .Z(n10574) );
  NAND U10911 ( .A(n10575), .B(n10574), .Z(n10647) );
  NAND U10912 ( .A(n19808), .B(n10576), .Z(n10578) );
  XOR U10913 ( .A(b[13]), .B(a[133]), .Z(n10653) );
  NAND U10914 ( .A(n19768), .B(n10653), .Z(n10577) );
  AND U10915 ( .A(n10578), .B(n10577), .Z(n10645) );
  AND U10916 ( .A(b[15]), .B(a[129]), .Z(n10644) );
  XNOR U10917 ( .A(n10645), .B(n10644), .Z(n10646) );
  XNOR U10918 ( .A(n10647), .B(n10646), .Z(n10665) );
  NAND U10919 ( .A(n33), .B(n10579), .Z(n10581) );
  XOR U10920 ( .A(b[5]), .B(a[141]), .Z(n10656) );
  NAND U10921 ( .A(n19342), .B(n10656), .Z(n10580) );
  AND U10922 ( .A(n10581), .B(n10580), .Z(n10689) );
  NAND U10923 ( .A(n34), .B(n10582), .Z(n10584) );
  XOR U10924 ( .A(b[7]), .B(a[139]), .Z(n10659) );
  NAND U10925 ( .A(n19486), .B(n10659), .Z(n10583) );
  AND U10926 ( .A(n10584), .B(n10583), .Z(n10687) );
  NAND U10927 ( .A(n31), .B(n10585), .Z(n10587) );
  XOR U10928 ( .A(b[3]), .B(a[143]), .Z(n10662) );
  NAND U10929 ( .A(n32), .B(n10662), .Z(n10586) );
  NAND U10930 ( .A(n10587), .B(n10586), .Z(n10686) );
  XNOR U10931 ( .A(n10687), .B(n10686), .Z(n10688) );
  XOR U10932 ( .A(n10689), .B(n10688), .Z(n10666) );
  XOR U10933 ( .A(n10665), .B(n10666), .Z(n10668) );
  XOR U10934 ( .A(n10667), .B(n10668), .Z(n10639) );
  NANDN U10935 ( .A(n10589), .B(n10588), .Z(n10593) );
  OR U10936 ( .A(n10591), .B(n10590), .Z(n10592) );
  AND U10937 ( .A(n10593), .B(n10592), .Z(n10638) );
  XNOR U10938 ( .A(n10639), .B(n10638), .Z(n10641) );
  NAND U10939 ( .A(n10594), .B(n19724), .Z(n10596) );
  XOR U10940 ( .A(b[11]), .B(a[135]), .Z(n10671) );
  NAND U10941 ( .A(n19692), .B(n10671), .Z(n10595) );
  AND U10942 ( .A(n10596), .B(n10595), .Z(n10682) );
  NAND U10943 ( .A(n19838), .B(n10597), .Z(n10599) );
  XOR U10944 ( .A(b[15]), .B(a[131]), .Z(n10674) );
  NAND U10945 ( .A(n19805), .B(n10674), .Z(n10598) );
  AND U10946 ( .A(n10599), .B(n10598), .Z(n10681) );
  NAND U10947 ( .A(n35), .B(n10600), .Z(n10602) );
  XOR U10948 ( .A(b[9]), .B(a[137]), .Z(n10677) );
  NAND U10949 ( .A(n19598), .B(n10677), .Z(n10601) );
  NAND U10950 ( .A(n10602), .B(n10601), .Z(n10680) );
  XOR U10951 ( .A(n10681), .B(n10680), .Z(n10683) );
  XOR U10952 ( .A(n10682), .B(n10683), .Z(n10693) );
  NANDN U10953 ( .A(n10604), .B(n10603), .Z(n10608) );
  OR U10954 ( .A(n10606), .B(n10605), .Z(n10607) );
  AND U10955 ( .A(n10608), .B(n10607), .Z(n10692) );
  XNOR U10956 ( .A(n10693), .B(n10692), .Z(n10694) );
  NANDN U10957 ( .A(n10610), .B(n10609), .Z(n10614) );
  NANDN U10958 ( .A(n10612), .B(n10611), .Z(n10613) );
  NAND U10959 ( .A(n10614), .B(n10613), .Z(n10695) );
  XNOR U10960 ( .A(n10694), .B(n10695), .Z(n10640) );
  XOR U10961 ( .A(n10641), .B(n10640), .Z(n10699) );
  NANDN U10962 ( .A(n10616), .B(n10615), .Z(n10620) );
  NANDN U10963 ( .A(n10618), .B(n10617), .Z(n10619) );
  AND U10964 ( .A(n10620), .B(n10619), .Z(n10698) );
  XNOR U10965 ( .A(n10699), .B(n10698), .Z(n10700) );
  XOR U10966 ( .A(n10701), .B(n10700), .Z(n10633) );
  NANDN U10967 ( .A(n10622), .B(n10621), .Z(n10626) );
  NAND U10968 ( .A(n10624), .B(n10623), .Z(n10625) );
  AND U10969 ( .A(n10626), .B(n10625), .Z(n10632) );
  XNOR U10970 ( .A(n10633), .B(n10632), .Z(n10634) );
  XNOR U10971 ( .A(n10635), .B(n10634), .Z(n10704) );
  XNOR U10972 ( .A(sreg[385]), .B(n10704), .Z(n10706) );
  NANDN U10973 ( .A(sreg[384]), .B(n10627), .Z(n10631) );
  NAND U10974 ( .A(n10629), .B(n10628), .Z(n10630) );
  NAND U10975 ( .A(n10631), .B(n10630), .Z(n10705) );
  XNOR U10976 ( .A(n10706), .B(n10705), .Z(c[385]) );
  NANDN U10977 ( .A(n10633), .B(n10632), .Z(n10637) );
  NANDN U10978 ( .A(n10635), .B(n10634), .Z(n10636) );
  AND U10979 ( .A(n10637), .B(n10636), .Z(n10712) );
  NANDN U10980 ( .A(n10639), .B(n10638), .Z(n10643) );
  NAND U10981 ( .A(n10641), .B(n10640), .Z(n10642) );
  AND U10982 ( .A(n10643), .B(n10642), .Z(n10778) );
  NANDN U10983 ( .A(n10645), .B(n10644), .Z(n10649) );
  NANDN U10984 ( .A(n10647), .B(n10646), .Z(n10648) );
  AND U10985 ( .A(n10649), .B(n10648), .Z(n10744) );
  NAND U10986 ( .A(b[0]), .B(a[146]), .Z(n10650) );
  XNOR U10987 ( .A(b[1]), .B(n10650), .Z(n10652) );
  NANDN U10988 ( .A(b[0]), .B(a[145]), .Z(n10651) );
  NAND U10989 ( .A(n10652), .B(n10651), .Z(n10724) );
  NAND U10990 ( .A(n19808), .B(n10653), .Z(n10655) );
  XOR U10991 ( .A(b[13]), .B(a[134]), .Z(n10730) );
  NAND U10992 ( .A(n19768), .B(n10730), .Z(n10654) );
  AND U10993 ( .A(n10655), .B(n10654), .Z(n10722) );
  AND U10994 ( .A(b[15]), .B(a[130]), .Z(n10721) );
  XNOR U10995 ( .A(n10722), .B(n10721), .Z(n10723) );
  XNOR U10996 ( .A(n10724), .B(n10723), .Z(n10742) );
  NAND U10997 ( .A(n33), .B(n10656), .Z(n10658) );
  XOR U10998 ( .A(b[5]), .B(a[142]), .Z(n10733) );
  NAND U10999 ( .A(n19342), .B(n10733), .Z(n10657) );
  AND U11000 ( .A(n10658), .B(n10657), .Z(n10766) );
  NAND U11001 ( .A(n34), .B(n10659), .Z(n10661) );
  XOR U11002 ( .A(b[7]), .B(a[140]), .Z(n10736) );
  NAND U11003 ( .A(n19486), .B(n10736), .Z(n10660) );
  AND U11004 ( .A(n10661), .B(n10660), .Z(n10764) );
  NAND U11005 ( .A(n31), .B(n10662), .Z(n10664) );
  XOR U11006 ( .A(b[3]), .B(a[144]), .Z(n10739) );
  NAND U11007 ( .A(n32), .B(n10739), .Z(n10663) );
  NAND U11008 ( .A(n10664), .B(n10663), .Z(n10763) );
  XNOR U11009 ( .A(n10764), .B(n10763), .Z(n10765) );
  XOR U11010 ( .A(n10766), .B(n10765), .Z(n10743) );
  XOR U11011 ( .A(n10742), .B(n10743), .Z(n10745) );
  XOR U11012 ( .A(n10744), .B(n10745), .Z(n10716) );
  NANDN U11013 ( .A(n10666), .B(n10665), .Z(n10670) );
  OR U11014 ( .A(n10668), .B(n10667), .Z(n10669) );
  AND U11015 ( .A(n10670), .B(n10669), .Z(n10715) );
  XNOR U11016 ( .A(n10716), .B(n10715), .Z(n10718) );
  NAND U11017 ( .A(n10671), .B(n19724), .Z(n10673) );
  XOR U11018 ( .A(b[11]), .B(a[136]), .Z(n10748) );
  NAND U11019 ( .A(n19692), .B(n10748), .Z(n10672) );
  AND U11020 ( .A(n10673), .B(n10672), .Z(n10759) );
  NAND U11021 ( .A(n19838), .B(n10674), .Z(n10676) );
  XOR U11022 ( .A(b[15]), .B(a[132]), .Z(n10751) );
  NAND U11023 ( .A(n19805), .B(n10751), .Z(n10675) );
  AND U11024 ( .A(n10676), .B(n10675), .Z(n10758) );
  NAND U11025 ( .A(n35), .B(n10677), .Z(n10679) );
  XOR U11026 ( .A(b[9]), .B(a[138]), .Z(n10754) );
  NAND U11027 ( .A(n19598), .B(n10754), .Z(n10678) );
  NAND U11028 ( .A(n10679), .B(n10678), .Z(n10757) );
  XOR U11029 ( .A(n10758), .B(n10757), .Z(n10760) );
  XOR U11030 ( .A(n10759), .B(n10760), .Z(n10770) );
  NANDN U11031 ( .A(n10681), .B(n10680), .Z(n10685) );
  OR U11032 ( .A(n10683), .B(n10682), .Z(n10684) );
  AND U11033 ( .A(n10685), .B(n10684), .Z(n10769) );
  XNOR U11034 ( .A(n10770), .B(n10769), .Z(n10771) );
  NANDN U11035 ( .A(n10687), .B(n10686), .Z(n10691) );
  NANDN U11036 ( .A(n10689), .B(n10688), .Z(n10690) );
  NAND U11037 ( .A(n10691), .B(n10690), .Z(n10772) );
  XNOR U11038 ( .A(n10771), .B(n10772), .Z(n10717) );
  XOR U11039 ( .A(n10718), .B(n10717), .Z(n10776) );
  NANDN U11040 ( .A(n10693), .B(n10692), .Z(n10697) );
  NANDN U11041 ( .A(n10695), .B(n10694), .Z(n10696) );
  AND U11042 ( .A(n10697), .B(n10696), .Z(n10775) );
  XNOR U11043 ( .A(n10776), .B(n10775), .Z(n10777) );
  XOR U11044 ( .A(n10778), .B(n10777), .Z(n10710) );
  NANDN U11045 ( .A(n10699), .B(n10698), .Z(n10703) );
  NAND U11046 ( .A(n10701), .B(n10700), .Z(n10702) );
  AND U11047 ( .A(n10703), .B(n10702), .Z(n10709) );
  XNOR U11048 ( .A(n10710), .B(n10709), .Z(n10711) );
  XNOR U11049 ( .A(n10712), .B(n10711), .Z(n10781) );
  XNOR U11050 ( .A(sreg[386]), .B(n10781), .Z(n10783) );
  NANDN U11051 ( .A(sreg[385]), .B(n10704), .Z(n10708) );
  NAND U11052 ( .A(n10706), .B(n10705), .Z(n10707) );
  NAND U11053 ( .A(n10708), .B(n10707), .Z(n10782) );
  XNOR U11054 ( .A(n10783), .B(n10782), .Z(c[386]) );
  NANDN U11055 ( .A(n10710), .B(n10709), .Z(n10714) );
  NANDN U11056 ( .A(n10712), .B(n10711), .Z(n10713) );
  AND U11057 ( .A(n10714), .B(n10713), .Z(n10789) );
  NANDN U11058 ( .A(n10716), .B(n10715), .Z(n10720) );
  NAND U11059 ( .A(n10718), .B(n10717), .Z(n10719) );
  AND U11060 ( .A(n10720), .B(n10719), .Z(n10855) );
  NANDN U11061 ( .A(n10722), .B(n10721), .Z(n10726) );
  NANDN U11062 ( .A(n10724), .B(n10723), .Z(n10725) );
  AND U11063 ( .A(n10726), .B(n10725), .Z(n10821) );
  NAND U11064 ( .A(b[0]), .B(a[147]), .Z(n10727) );
  XNOR U11065 ( .A(b[1]), .B(n10727), .Z(n10729) );
  NANDN U11066 ( .A(b[0]), .B(a[146]), .Z(n10728) );
  NAND U11067 ( .A(n10729), .B(n10728), .Z(n10801) );
  NAND U11068 ( .A(n19808), .B(n10730), .Z(n10732) );
  XOR U11069 ( .A(b[13]), .B(a[135]), .Z(n10807) );
  NAND U11070 ( .A(n19768), .B(n10807), .Z(n10731) );
  AND U11071 ( .A(n10732), .B(n10731), .Z(n10799) );
  AND U11072 ( .A(b[15]), .B(a[131]), .Z(n10798) );
  XNOR U11073 ( .A(n10799), .B(n10798), .Z(n10800) );
  XNOR U11074 ( .A(n10801), .B(n10800), .Z(n10819) );
  NAND U11075 ( .A(n33), .B(n10733), .Z(n10735) );
  XOR U11076 ( .A(b[5]), .B(a[143]), .Z(n10810) );
  NAND U11077 ( .A(n19342), .B(n10810), .Z(n10734) );
  AND U11078 ( .A(n10735), .B(n10734), .Z(n10843) );
  NAND U11079 ( .A(n34), .B(n10736), .Z(n10738) );
  XOR U11080 ( .A(b[7]), .B(a[141]), .Z(n10813) );
  NAND U11081 ( .A(n19486), .B(n10813), .Z(n10737) );
  AND U11082 ( .A(n10738), .B(n10737), .Z(n10841) );
  NAND U11083 ( .A(n31), .B(n10739), .Z(n10741) );
  XOR U11084 ( .A(b[3]), .B(a[145]), .Z(n10816) );
  NAND U11085 ( .A(n32), .B(n10816), .Z(n10740) );
  NAND U11086 ( .A(n10741), .B(n10740), .Z(n10840) );
  XNOR U11087 ( .A(n10841), .B(n10840), .Z(n10842) );
  XOR U11088 ( .A(n10843), .B(n10842), .Z(n10820) );
  XOR U11089 ( .A(n10819), .B(n10820), .Z(n10822) );
  XOR U11090 ( .A(n10821), .B(n10822), .Z(n10793) );
  NANDN U11091 ( .A(n10743), .B(n10742), .Z(n10747) );
  OR U11092 ( .A(n10745), .B(n10744), .Z(n10746) );
  AND U11093 ( .A(n10747), .B(n10746), .Z(n10792) );
  XNOR U11094 ( .A(n10793), .B(n10792), .Z(n10795) );
  NAND U11095 ( .A(n10748), .B(n19724), .Z(n10750) );
  XOR U11096 ( .A(b[11]), .B(a[137]), .Z(n10825) );
  NAND U11097 ( .A(n19692), .B(n10825), .Z(n10749) );
  AND U11098 ( .A(n10750), .B(n10749), .Z(n10836) );
  NAND U11099 ( .A(n19838), .B(n10751), .Z(n10753) );
  XOR U11100 ( .A(b[15]), .B(a[133]), .Z(n10828) );
  NAND U11101 ( .A(n19805), .B(n10828), .Z(n10752) );
  AND U11102 ( .A(n10753), .B(n10752), .Z(n10835) );
  NAND U11103 ( .A(n35), .B(n10754), .Z(n10756) );
  XOR U11104 ( .A(b[9]), .B(a[139]), .Z(n10831) );
  NAND U11105 ( .A(n19598), .B(n10831), .Z(n10755) );
  NAND U11106 ( .A(n10756), .B(n10755), .Z(n10834) );
  XOR U11107 ( .A(n10835), .B(n10834), .Z(n10837) );
  XOR U11108 ( .A(n10836), .B(n10837), .Z(n10847) );
  NANDN U11109 ( .A(n10758), .B(n10757), .Z(n10762) );
  OR U11110 ( .A(n10760), .B(n10759), .Z(n10761) );
  AND U11111 ( .A(n10762), .B(n10761), .Z(n10846) );
  XNOR U11112 ( .A(n10847), .B(n10846), .Z(n10848) );
  NANDN U11113 ( .A(n10764), .B(n10763), .Z(n10768) );
  NANDN U11114 ( .A(n10766), .B(n10765), .Z(n10767) );
  NAND U11115 ( .A(n10768), .B(n10767), .Z(n10849) );
  XNOR U11116 ( .A(n10848), .B(n10849), .Z(n10794) );
  XOR U11117 ( .A(n10795), .B(n10794), .Z(n10853) );
  NANDN U11118 ( .A(n10770), .B(n10769), .Z(n10774) );
  NANDN U11119 ( .A(n10772), .B(n10771), .Z(n10773) );
  AND U11120 ( .A(n10774), .B(n10773), .Z(n10852) );
  XNOR U11121 ( .A(n10853), .B(n10852), .Z(n10854) );
  XOR U11122 ( .A(n10855), .B(n10854), .Z(n10787) );
  NANDN U11123 ( .A(n10776), .B(n10775), .Z(n10780) );
  NAND U11124 ( .A(n10778), .B(n10777), .Z(n10779) );
  AND U11125 ( .A(n10780), .B(n10779), .Z(n10786) );
  XNOR U11126 ( .A(n10787), .B(n10786), .Z(n10788) );
  XNOR U11127 ( .A(n10789), .B(n10788), .Z(n10858) );
  XNOR U11128 ( .A(sreg[387]), .B(n10858), .Z(n10860) );
  NANDN U11129 ( .A(sreg[386]), .B(n10781), .Z(n10785) );
  NAND U11130 ( .A(n10783), .B(n10782), .Z(n10784) );
  NAND U11131 ( .A(n10785), .B(n10784), .Z(n10859) );
  XNOR U11132 ( .A(n10860), .B(n10859), .Z(c[387]) );
  NANDN U11133 ( .A(n10787), .B(n10786), .Z(n10791) );
  NANDN U11134 ( .A(n10789), .B(n10788), .Z(n10790) );
  AND U11135 ( .A(n10791), .B(n10790), .Z(n10866) );
  NANDN U11136 ( .A(n10793), .B(n10792), .Z(n10797) );
  NAND U11137 ( .A(n10795), .B(n10794), .Z(n10796) );
  AND U11138 ( .A(n10797), .B(n10796), .Z(n10932) );
  NANDN U11139 ( .A(n10799), .B(n10798), .Z(n10803) );
  NANDN U11140 ( .A(n10801), .B(n10800), .Z(n10802) );
  AND U11141 ( .A(n10803), .B(n10802), .Z(n10898) );
  NAND U11142 ( .A(b[0]), .B(a[148]), .Z(n10804) );
  XNOR U11143 ( .A(b[1]), .B(n10804), .Z(n10806) );
  NANDN U11144 ( .A(b[0]), .B(a[147]), .Z(n10805) );
  NAND U11145 ( .A(n10806), .B(n10805), .Z(n10878) );
  NAND U11146 ( .A(n19808), .B(n10807), .Z(n10809) );
  XOR U11147 ( .A(b[13]), .B(a[136]), .Z(n10884) );
  NAND U11148 ( .A(n19768), .B(n10884), .Z(n10808) );
  AND U11149 ( .A(n10809), .B(n10808), .Z(n10876) );
  AND U11150 ( .A(b[15]), .B(a[132]), .Z(n10875) );
  XNOR U11151 ( .A(n10876), .B(n10875), .Z(n10877) );
  XNOR U11152 ( .A(n10878), .B(n10877), .Z(n10896) );
  NAND U11153 ( .A(n33), .B(n10810), .Z(n10812) );
  XOR U11154 ( .A(b[5]), .B(a[144]), .Z(n10887) );
  NAND U11155 ( .A(n19342), .B(n10887), .Z(n10811) );
  AND U11156 ( .A(n10812), .B(n10811), .Z(n10920) );
  NAND U11157 ( .A(n34), .B(n10813), .Z(n10815) );
  XOR U11158 ( .A(b[7]), .B(a[142]), .Z(n10890) );
  NAND U11159 ( .A(n19486), .B(n10890), .Z(n10814) );
  AND U11160 ( .A(n10815), .B(n10814), .Z(n10918) );
  NAND U11161 ( .A(n31), .B(n10816), .Z(n10818) );
  XOR U11162 ( .A(b[3]), .B(a[146]), .Z(n10893) );
  NAND U11163 ( .A(n32), .B(n10893), .Z(n10817) );
  NAND U11164 ( .A(n10818), .B(n10817), .Z(n10917) );
  XNOR U11165 ( .A(n10918), .B(n10917), .Z(n10919) );
  XOR U11166 ( .A(n10920), .B(n10919), .Z(n10897) );
  XOR U11167 ( .A(n10896), .B(n10897), .Z(n10899) );
  XOR U11168 ( .A(n10898), .B(n10899), .Z(n10870) );
  NANDN U11169 ( .A(n10820), .B(n10819), .Z(n10824) );
  OR U11170 ( .A(n10822), .B(n10821), .Z(n10823) );
  AND U11171 ( .A(n10824), .B(n10823), .Z(n10869) );
  XNOR U11172 ( .A(n10870), .B(n10869), .Z(n10872) );
  NAND U11173 ( .A(n10825), .B(n19724), .Z(n10827) );
  XOR U11174 ( .A(b[11]), .B(a[138]), .Z(n10902) );
  NAND U11175 ( .A(n19692), .B(n10902), .Z(n10826) );
  AND U11176 ( .A(n10827), .B(n10826), .Z(n10913) );
  NAND U11177 ( .A(n19838), .B(n10828), .Z(n10830) );
  XOR U11178 ( .A(b[15]), .B(a[134]), .Z(n10905) );
  NAND U11179 ( .A(n19805), .B(n10905), .Z(n10829) );
  AND U11180 ( .A(n10830), .B(n10829), .Z(n10912) );
  NAND U11181 ( .A(n35), .B(n10831), .Z(n10833) );
  XOR U11182 ( .A(b[9]), .B(a[140]), .Z(n10908) );
  NAND U11183 ( .A(n19598), .B(n10908), .Z(n10832) );
  NAND U11184 ( .A(n10833), .B(n10832), .Z(n10911) );
  XOR U11185 ( .A(n10912), .B(n10911), .Z(n10914) );
  XOR U11186 ( .A(n10913), .B(n10914), .Z(n10924) );
  NANDN U11187 ( .A(n10835), .B(n10834), .Z(n10839) );
  OR U11188 ( .A(n10837), .B(n10836), .Z(n10838) );
  AND U11189 ( .A(n10839), .B(n10838), .Z(n10923) );
  XNOR U11190 ( .A(n10924), .B(n10923), .Z(n10925) );
  NANDN U11191 ( .A(n10841), .B(n10840), .Z(n10845) );
  NANDN U11192 ( .A(n10843), .B(n10842), .Z(n10844) );
  NAND U11193 ( .A(n10845), .B(n10844), .Z(n10926) );
  XNOR U11194 ( .A(n10925), .B(n10926), .Z(n10871) );
  XOR U11195 ( .A(n10872), .B(n10871), .Z(n10930) );
  NANDN U11196 ( .A(n10847), .B(n10846), .Z(n10851) );
  NANDN U11197 ( .A(n10849), .B(n10848), .Z(n10850) );
  AND U11198 ( .A(n10851), .B(n10850), .Z(n10929) );
  XNOR U11199 ( .A(n10930), .B(n10929), .Z(n10931) );
  XOR U11200 ( .A(n10932), .B(n10931), .Z(n10864) );
  NANDN U11201 ( .A(n10853), .B(n10852), .Z(n10857) );
  NAND U11202 ( .A(n10855), .B(n10854), .Z(n10856) );
  AND U11203 ( .A(n10857), .B(n10856), .Z(n10863) );
  XNOR U11204 ( .A(n10864), .B(n10863), .Z(n10865) );
  XNOR U11205 ( .A(n10866), .B(n10865), .Z(n10935) );
  XNOR U11206 ( .A(sreg[388]), .B(n10935), .Z(n10937) );
  NANDN U11207 ( .A(sreg[387]), .B(n10858), .Z(n10862) );
  NAND U11208 ( .A(n10860), .B(n10859), .Z(n10861) );
  NAND U11209 ( .A(n10862), .B(n10861), .Z(n10936) );
  XNOR U11210 ( .A(n10937), .B(n10936), .Z(c[388]) );
  NANDN U11211 ( .A(n10864), .B(n10863), .Z(n10868) );
  NANDN U11212 ( .A(n10866), .B(n10865), .Z(n10867) );
  AND U11213 ( .A(n10868), .B(n10867), .Z(n10943) );
  NANDN U11214 ( .A(n10870), .B(n10869), .Z(n10874) );
  NAND U11215 ( .A(n10872), .B(n10871), .Z(n10873) );
  AND U11216 ( .A(n10874), .B(n10873), .Z(n11009) );
  NANDN U11217 ( .A(n10876), .B(n10875), .Z(n10880) );
  NANDN U11218 ( .A(n10878), .B(n10877), .Z(n10879) );
  AND U11219 ( .A(n10880), .B(n10879), .Z(n10975) );
  NAND U11220 ( .A(b[0]), .B(a[149]), .Z(n10881) );
  XNOR U11221 ( .A(b[1]), .B(n10881), .Z(n10883) );
  NANDN U11222 ( .A(b[0]), .B(a[148]), .Z(n10882) );
  NAND U11223 ( .A(n10883), .B(n10882), .Z(n10955) );
  NAND U11224 ( .A(n19808), .B(n10884), .Z(n10886) );
  XOR U11225 ( .A(b[13]), .B(a[137]), .Z(n10961) );
  NAND U11226 ( .A(n19768), .B(n10961), .Z(n10885) );
  AND U11227 ( .A(n10886), .B(n10885), .Z(n10953) );
  AND U11228 ( .A(b[15]), .B(a[133]), .Z(n10952) );
  XNOR U11229 ( .A(n10953), .B(n10952), .Z(n10954) );
  XNOR U11230 ( .A(n10955), .B(n10954), .Z(n10973) );
  NAND U11231 ( .A(n33), .B(n10887), .Z(n10889) );
  XOR U11232 ( .A(b[5]), .B(a[145]), .Z(n10964) );
  NAND U11233 ( .A(n19342), .B(n10964), .Z(n10888) );
  AND U11234 ( .A(n10889), .B(n10888), .Z(n10997) );
  NAND U11235 ( .A(n34), .B(n10890), .Z(n10892) );
  XOR U11236 ( .A(b[7]), .B(a[143]), .Z(n10967) );
  NAND U11237 ( .A(n19486), .B(n10967), .Z(n10891) );
  AND U11238 ( .A(n10892), .B(n10891), .Z(n10995) );
  NAND U11239 ( .A(n31), .B(n10893), .Z(n10895) );
  XOR U11240 ( .A(b[3]), .B(a[147]), .Z(n10970) );
  NAND U11241 ( .A(n32), .B(n10970), .Z(n10894) );
  NAND U11242 ( .A(n10895), .B(n10894), .Z(n10994) );
  XNOR U11243 ( .A(n10995), .B(n10994), .Z(n10996) );
  XOR U11244 ( .A(n10997), .B(n10996), .Z(n10974) );
  XOR U11245 ( .A(n10973), .B(n10974), .Z(n10976) );
  XOR U11246 ( .A(n10975), .B(n10976), .Z(n10947) );
  NANDN U11247 ( .A(n10897), .B(n10896), .Z(n10901) );
  OR U11248 ( .A(n10899), .B(n10898), .Z(n10900) );
  AND U11249 ( .A(n10901), .B(n10900), .Z(n10946) );
  XNOR U11250 ( .A(n10947), .B(n10946), .Z(n10949) );
  NAND U11251 ( .A(n10902), .B(n19724), .Z(n10904) );
  XOR U11252 ( .A(b[11]), .B(a[139]), .Z(n10979) );
  NAND U11253 ( .A(n19692), .B(n10979), .Z(n10903) );
  AND U11254 ( .A(n10904), .B(n10903), .Z(n10990) );
  NAND U11255 ( .A(n19838), .B(n10905), .Z(n10907) );
  XOR U11256 ( .A(b[15]), .B(a[135]), .Z(n10982) );
  NAND U11257 ( .A(n19805), .B(n10982), .Z(n10906) );
  AND U11258 ( .A(n10907), .B(n10906), .Z(n10989) );
  NAND U11259 ( .A(n35), .B(n10908), .Z(n10910) );
  XOR U11260 ( .A(b[9]), .B(a[141]), .Z(n10985) );
  NAND U11261 ( .A(n19598), .B(n10985), .Z(n10909) );
  NAND U11262 ( .A(n10910), .B(n10909), .Z(n10988) );
  XOR U11263 ( .A(n10989), .B(n10988), .Z(n10991) );
  XOR U11264 ( .A(n10990), .B(n10991), .Z(n11001) );
  NANDN U11265 ( .A(n10912), .B(n10911), .Z(n10916) );
  OR U11266 ( .A(n10914), .B(n10913), .Z(n10915) );
  AND U11267 ( .A(n10916), .B(n10915), .Z(n11000) );
  XNOR U11268 ( .A(n11001), .B(n11000), .Z(n11002) );
  NANDN U11269 ( .A(n10918), .B(n10917), .Z(n10922) );
  NANDN U11270 ( .A(n10920), .B(n10919), .Z(n10921) );
  NAND U11271 ( .A(n10922), .B(n10921), .Z(n11003) );
  XNOR U11272 ( .A(n11002), .B(n11003), .Z(n10948) );
  XOR U11273 ( .A(n10949), .B(n10948), .Z(n11007) );
  NANDN U11274 ( .A(n10924), .B(n10923), .Z(n10928) );
  NANDN U11275 ( .A(n10926), .B(n10925), .Z(n10927) );
  AND U11276 ( .A(n10928), .B(n10927), .Z(n11006) );
  XNOR U11277 ( .A(n11007), .B(n11006), .Z(n11008) );
  XOR U11278 ( .A(n11009), .B(n11008), .Z(n10941) );
  NANDN U11279 ( .A(n10930), .B(n10929), .Z(n10934) );
  NAND U11280 ( .A(n10932), .B(n10931), .Z(n10933) );
  AND U11281 ( .A(n10934), .B(n10933), .Z(n10940) );
  XNOR U11282 ( .A(n10941), .B(n10940), .Z(n10942) );
  XNOR U11283 ( .A(n10943), .B(n10942), .Z(n11012) );
  XNOR U11284 ( .A(sreg[389]), .B(n11012), .Z(n11014) );
  NANDN U11285 ( .A(sreg[388]), .B(n10935), .Z(n10939) );
  NAND U11286 ( .A(n10937), .B(n10936), .Z(n10938) );
  NAND U11287 ( .A(n10939), .B(n10938), .Z(n11013) );
  XNOR U11288 ( .A(n11014), .B(n11013), .Z(c[389]) );
  NANDN U11289 ( .A(n10941), .B(n10940), .Z(n10945) );
  NANDN U11290 ( .A(n10943), .B(n10942), .Z(n10944) );
  AND U11291 ( .A(n10945), .B(n10944), .Z(n11020) );
  NANDN U11292 ( .A(n10947), .B(n10946), .Z(n10951) );
  NAND U11293 ( .A(n10949), .B(n10948), .Z(n10950) );
  AND U11294 ( .A(n10951), .B(n10950), .Z(n11086) );
  NANDN U11295 ( .A(n10953), .B(n10952), .Z(n10957) );
  NANDN U11296 ( .A(n10955), .B(n10954), .Z(n10956) );
  AND U11297 ( .A(n10957), .B(n10956), .Z(n11052) );
  NAND U11298 ( .A(b[0]), .B(a[150]), .Z(n10958) );
  XNOR U11299 ( .A(b[1]), .B(n10958), .Z(n10960) );
  NANDN U11300 ( .A(b[0]), .B(a[149]), .Z(n10959) );
  NAND U11301 ( .A(n10960), .B(n10959), .Z(n11032) );
  NAND U11302 ( .A(n19808), .B(n10961), .Z(n10963) );
  XOR U11303 ( .A(b[13]), .B(a[138]), .Z(n11038) );
  NAND U11304 ( .A(n19768), .B(n11038), .Z(n10962) );
  AND U11305 ( .A(n10963), .B(n10962), .Z(n11030) );
  AND U11306 ( .A(b[15]), .B(a[134]), .Z(n11029) );
  XNOR U11307 ( .A(n11030), .B(n11029), .Z(n11031) );
  XNOR U11308 ( .A(n11032), .B(n11031), .Z(n11050) );
  NAND U11309 ( .A(n33), .B(n10964), .Z(n10966) );
  XOR U11310 ( .A(b[5]), .B(a[146]), .Z(n11041) );
  NAND U11311 ( .A(n19342), .B(n11041), .Z(n10965) );
  AND U11312 ( .A(n10966), .B(n10965), .Z(n11074) );
  NAND U11313 ( .A(n34), .B(n10967), .Z(n10969) );
  XOR U11314 ( .A(b[7]), .B(a[144]), .Z(n11044) );
  NAND U11315 ( .A(n19486), .B(n11044), .Z(n10968) );
  AND U11316 ( .A(n10969), .B(n10968), .Z(n11072) );
  NAND U11317 ( .A(n31), .B(n10970), .Z(n10972) );
  XOR U11318 ( .A(b[3]), .B(a[148]), .Z(n11047) );
  NAND U11319 ( .A(n32), .B(n11047), .Z(n10971) );
  NAND U11320 ( .A(n10972), .B(n10971), .Z(n11071) );
  XNOR U11321 ( .A(n11072), .B(n11071), .Z(n11073) );
  XOR U11322 ( .A(n11074), .B(n11073), .Z(n11051) );
  XOR U11323 ( .A(n11050), .B(n11051), .Z(n11053) );
  XOR U11324 ( .A(n11052), .B(n11053), .Z(n11024) );
  NANDN U11325 ( .A(n10974), .B(n10973), .Z(n10978) );
  OR U11326 ( .A(n10976), .B(n10975), .Z(n10977) );
  AND U11327 ( .A(n10978), .B(n10977), .Z(n11023) );
  XNOR U11328 ( .A(n11024), .B(n11023), .Z(n11026) );
  NAND U11329 ( .A(n10979), .B(n19724), .Z(n10981) );
  XOR U11330 ( .A(b[11]), .B(a[140]), .Z(n11056) );
  NAND U11331 ( .A(n19692), .B(n11056), .Z(n10980) );
  AND U11332 ( .A(n10981), .B(n10980), .Z(n11067) );
  NAND U11333 ( .A(n19838), .B(n10982), .Z(n10984) );
  XOR U11334 ( .A(b[15]), .B(a[136]), .Z(n11059) );
  NAND U11335 ( .A(n19805), .B(n11059), .Z(n10983) );
  AND U11336 ( .A(n10984), .B(n10983), .Z(n11066) );
  NAND U11337 ( .A(n35), .B(n10985), .Z(n10987) );
  XOR U11338 ( .A(b[9]), .B(a[142]), .Z(n11062) );
  NAND U11339 ( .A(n19598), .B(n11062), .Z(n10986) );
  NAND U11340 ( .A(n10987), .B(n10986), .Z(n11065) );
  XOR U11341 ( .A(n11066), .B(n11065), .Z(n11068) );
  XOR U11342 ( .A(n11067), .B(n11068), .Z(n11078) );
  NANDN U11343 ( .A(n10989), .B(n10988), .Z(n10993) );
  OR U11344 ( .A(n10991), .B(n10990), .Z(n10992) );
  AND U11345 ( .A(n10993), .B(n10992), .Z(n11077) );
  XNOR U11346 ( .A(n11078), .B(n11077), .Z(n11079) );
  NANDN U11347 ( .A(n10995), .B(n10994), .Z(n10999) );
  NANDN U11348 ( .A(n10997), .B(n10996), .Z(n10998) );
  NAND U11349 ( .A(n10999), .B(n10998), .Z(n11080) );
  XNOR U11350 ( .A(n11079), .B(n11080), .Z(n11025) );
  XOR U11351 ( .A(n11026), .B(n11025), .Z(n11084) );
  NANDN U11352 ( .A(n11001), .B(n11000), .Z(n11005) );
  NANDN U11353 ( .A(n11003), .B(n11002), .Z(n11004) );
  AND U11354 ( .A(n11005), .B(n11004), .Z(n11083) );
  XNOR U11355 ( .A(n11084), .B(n11083), .Z(n11085) );
  XOR U11356 ( .A(n11086), .B(n11085), .Z(n11018) );
  NANDN U11357 ( .A(n11007), .B(n11006), .Z(n11011) );
  NAND U11358 ( .A(n11009), .B(n11008), .Z(n11010) );
  AND U11359 ( .A(n11011), .B(n11010), .Z(n11017) );
  XNOR U11360 ( .A(n11018), .B(n11017), .Z(n11019) );
  XNOR U11361 ( .A(n11020), .B(n11019), .Z(n11089) );
  XNOR U11362 ( .A(sreg[390]), .B(n11089), .Z(n11091) );
  NANDN U11363 ( .A(sreg[389]), .B(n11012), .Z(n11016) );
  NAND U11364 ( .A(n11014), .B(n11013), .Z(n11015) );
  NAND U11365 ( .A(n11016), .B(n11015), .Z(n11090) );
  XNOR U11366 ( .A(n11091), .B(n11090), .Z(c[390]) );
  NANDN U11367 ( .A(n11018), .B(n11017), .Z(n11022) );
  NANDN U11368 ( .A(n11020), .B(n11019), .Z(n11021) );
  AND U11369 ( .A(n11022), .B(n11021), .Z(n11097) );
  NANDN U11370 ( .A(n11024), .B(n11023), .Z(n11028) );
  NAND U11371 ( .A(n11026), .B(n11025), .Z(n11027) );
  AND U11372 ( .A(n11028), .B(n11027), .Z(n11163) );
  NANDN U11373 ( .A(n11030), .B(n11029), .Z(n11034) );
  NANDN U11374 ( .A(n11032), .B(n11031), .Z(n11033) );
  AND U11375 ( .A(n11034), .B(n11033), .Z(n11150) );
  NAND U11376 ( .A(b[0]), .B(a[151]), .Z(n11035) );
  XNOR U11377 ( .A(b[1]), .B(n11035), .Z(n11037) );
  NANDN U11378 ( .A(b[0]), .B(a[150]), .Z(n11036) );
  NAND U11379 ( .A(n11037), .B(n11036), .Z(n11130) );
  NAND U11380 ( .A(n19808), .B(n11038), .Z(n11040) );
  XOR U11381 ( .A(b[13]), .B(a[139]), .Z(n11136) );
  NAND U11382 ( .A(n19768), .B(n11136), .Z(n11039) );
  AND U11383 ( .A(n11040), .B(n11039), .Z(n11128) );
  AND U11384 ( .A(b[15]), .B(a[135]), .Z(n11127) );
  XNOR U11385 ( .A(n11128), .B(n11127), .Z(n11129) );
  XNOR U11386 ( .A(n11130), .B(n11129), .Z(n11148) );
  NAND U11387 ( .A(n33), .B(n11041), .Z(n11043) );
  XOR U11388 ( .A(b[5]), .B(a[147]), .Z(n11139) );
  NAND U11389 ( .A(n19342), .B(n11139), .Z(n11042) );
  AND U11390 ( .A(n11043), .B(n11042), .Z(n11124) );
  NAND U11391 ( .A(n34), .B(n11044), .Z(n11046) );
  XOR U11392 ( .A(b[7]), .B(a[145]), .Z(n11142) );
  NAND U11393 ( .A(n19486), .B(n11142), .Z(n11045) );
  AND U11394 ( .A(n11046), .B(n11045), .Z(n11122) );
  NAND U11395 ( .A(n31), .B(n11047), .Z(n11049) );
  XOR U11396 ( .A(b[3]), .B(a[149]), .Z(n11145) );
  NAND U11397 ( .A(n32), .B(n11145), .Z(n11048) );
  NAND U11398 ( .A(n11049), .B(n11048), .Z(n11121) );
  XNOR U11399 ( .A(n11122), .B(n11121), .Z(n11123) );
  XOR U11400 ( .A(n11124), .B(n11123), .Z(n11149) );
  XOR U11401 ( .A(n11148), .B(n11149), .Z(n11151) );
  XOR U11402 ( .A(n11150), .B(n11151), .Z(n11101) );
  NANDN U11403 ( .A(n11051), .B(n11050), .Z(n11055) );
  OR U11404 ( .A(n11053), .B(n11052), .Z(n11054) );
  AND U11405 ( .A(n11055), .B(n11054), .Z(n11100) );
  XNOR U11406 ( .A(n11101), .B(n11100), .Z(n11103) );
  NAND U11407 ( .A(n11056), .B(n19724), .Z(n11058) );
  XOR U11408 ( .A(b[11]), .B(a[141]), .Z(n11106) );
  NAND U11409 ( .A(n19692), .B(n11106), .Z(n11057) );
  AND U11410 ( .A(n11058), .B(n11057), .Z(n11117) );
  NAND U11411 ( .A(n19838), .B(n11059), .Z(n11061) );
  XOR U11412 ( .A(b[15]), .B(a[137]), .Z(n11109) );
  NAND U11413 ( .A(n19805), .B(n11109), .Z(n11060) );
  AND U11414 ( .A(n11061), .B(n11060), .Z(n11116) );
  NAND U11415 ( .A(n35), .B(n11062), .Z(n11064) );
  XOR U11416 ( .A(b[9]), .B(a[143]), .Z(n11112) );
  NAND U11417 ( .A(n19598), .B(n11112), .Z(n11063) );
  NAND U11418 ( .A(n11064), .B(n11063), .Z(n11115) );
  XOR U11419 ( .A(n11116), .B(n11115), .Z(n11118) );
  XOR U11420 ( .A(n11117), .B(n11118), .Z(n11155) );
  NANDN U11421 ( .A(n11066), .B(n11065), .Z(n11070) );
  OR U11422 ( .A(n11068), .B(n11067), .Z(n11069) );
  AND U11423 ( .A(n11070), .B(n11069), .Z(n11154) );
  XNOR U11424 ( .A(n11155), .B(n11154), .Z(n11156) );
  NANDN U11425 ( .A(n11072), .B(n11071), .Z(n11076) );
  NANDN U11426 ( .A(n11074), .B(n11073), .Z(n11075) );
  NAND U11427 ( .A(n11076), .B(n11075), .Z(n11157) );
  XNOR U11428 ( .A(n11156), .B(n11157), .Z(n11102) );
  XOR U11429 ( .A(n11103), .B(n11102), .Z(n11161) );
  NANDN U11430 ( .A(n11078), .B(n11077), .Z(n11082) );
  NANDN U11431 ( .A(n11080), .B(n11079), .Z(n11081) );
  AND U11432 ( .A(n11082), .B(n11081), .Z(n11160) );
  XNOR U11433 ( .A(n11161), .B(n11160), .Z(n11162) );
  XOR U11434 ( .A(n11163), .B(n11162), .Z(n11095) );
  NANDN U11435 ( .A(n11084), .B(n11083), .Z(n11088) );
  NAND U11436 ( .A(n11086), .B(n11085), .Z(n11087) );
  AND U11437 ( .A(n11088), .B(n11087), .Z(n11094) );
  XNOR U11438 ( .A(n11095), .B(n11094), .Z(n11096) );
  XNOR U11439 ( .A(n11097), .B(n11096), .Z(n11166) );
  XNOR U11440 ( .A(sreg[391]), .B(n11166), .Z(n11168) );
  NANDN U11441 ( .A(sreg[390]), .B(n11089), .Z(n11093) );
  NAND U11442 ( .A(n11091), .B(n11090), .Z(n11092) );
  NAND U11443 ( .A(n11093), .B(n11092), .Z(n11167) );
  XNOR U11444 ( .A(n11168), .B(n11167), .Z(c[391]) );
  NANDN U11445 ( .A(n11095), .B(n11094), .Z(n11099) );
  NANDN U11446 ( .A(n11097), .B(n11096), .Z(n11098) );
  AND U11447 ( .A(n11099), .B(n11098), .Z(n11174) );
  NANDN U11448 ( .A(n11101), .B(n11100), .Z(n11105) );
  NAND U11449 ( .A(n11103), .B(n11102), .Z(n11104) );
  AND U11450 ( .A(n11105), .B(n11104), .Z(n11240) );
  NAND U11451 ( .A(n11106), .B(n19724), .Z(n11108) );
  XOR U11452 ( .A(b[11]), .B(a[142]), .Z(n11210) );
  NAND U11453 ( .A(n19692), .B(n11210), .Z(n11107) );
  AND U11454 ( .A(n11108), .B(n11107), .Z(n11221) );
  NAND U11455 ( .A(n19838), .B(n11109), .Z(n11111) );
  XOR U11456 ( .A(b[15]), .B(a[138]), .Z(n11213) );
  NAND U11457 ( .A(n19805), .B(n11213), .Z(n11110) );
  AND U11458 ( .A(n11111), .B(n11110), .Z(n11220) );
  NAND U11459 ( .A(n35), .B(n11112), .Z(n11114) );
  XOR U11460 ( .A(b[9]), .B(a[144]), .Z(n11216) );
  NAND U11461 ( .A(n19598), .B(n11216), .Z(n11113) );
  NAND U11462 ( .A(n11114), .B(n11113), .Z(n11219) );
  XOR U11463 ( .A(n11220), .B(n11219), .Z(n11222) );
  XOR U11464 ( .A(n11221), .B(n11222), .Z(n11232) );
  NANDN U11465 ( .A(n11116), .B(n11115), .Z(n11120) );
  OR U11466 ( .A(n11118), .B(n11117), .Z(n11119) );
  AND U11467 ( .A(n11120), .B(n11119), .Z(n11231) );
  XNOR U11468 ( .A(n11232), .B(n11231), .Z(n11233) );
  NANDN U11469 ( .A(n11122), .B(n11121), .Z(n11126) );
  NANDN U11470 ( .A(n11124), .B(n11123), .Z(n11125) );
  NAND U11471 ( .A(n11126), .B(n11125), .Z(n11234) );
  XNOR U11472 ( .A(n11233), .B(n11234), .Z(n11180) );
  NANDN U11473 ( .A(n11128), .B(n11127), .Z(n11132) );
  NANDN U11474 ( .A(n11130), .B(n11129), .Z(n11131) );
  AND U11475 ( .A(n11132), .B(n11131), .Z(n11206) );
  NAND U11476 ( .A(b[0]), .B(a[152]), .Z(n11133) );
  XNOR U11477 ( .A(b[1]), .B(n11133), .Z(n11135) );
  NANDN U11478 ( .A(b[0]), .B(a[151]), .Z(n11134) );
  NAND U11479 ( .A(n11135), .B(n11134), .Z(n11186) );
  NAND U11480 ( .A(n19808), .B(n11136), .Z(n11138) );
  XOR U11481 ( .A(b[13]), .B(a[140]), .Z(n11192) );
  NAND U11482 ( .A(n19768), .B(n11192), .Z(n11137) );
  AND U11483 ( .A(n11138), .B(n11137), .Z(n11184) );
  AND U11484 ( .A(b[15]), .B(a[136]), .Z(n11183) );
  XNOR U11485 ( .A(n11184), .B(n11183), .Z(n11185) );
  XNOR U11486 ( .A(n11186), .B(n11185), .Z(n11204) );
  NAND U11487 ( .A(n33), .B(n11139), .Z(n11141) );
  XOR U11488 ( .A(b[5]), .B(a[148]), .Z(n11195) );
  NAND U11489 ( .A(n19342), .B(n11195), .Z(n11140) );
  AND U11490 ( .A(n11141), .B(n11140), .Z(n11228) );
  NAND U11491 ( .A(n34), .B(n11142), .Z(n11144) );
  XOR U11492 ( .A(b[7]), .B(a[146]), .Z(n11198) );
  NAND U11493 ( .A(n19486), .B(n11198), .Z(n11143) );
  AND U11494 ( .A(n11144), .B(n11143), .Z(n11226) );
  NAND U11495 ( .A(n31), .B(n11145), .Z(n11147) );
  XOR U11496 ( .A(b[3]), .B(a[150]), .Z(n11201) );
  NAND U11497 ( .A(n32), .B(n11201), .Z(n11146) );
  NAND U11498 ( .A(n11147), .B(n11146), .Z(n11225) );
  XNOR U11499 ( .A(n11226), .B(n11225), .Z(n11227) );
  XOR U11500 ( .A(n11228), .B(n11227), .Z(n11205) );
  XOR U11501 ( .A(n11204), .B(n11205), .Z(n11207) );
  XOR U11502 ( .A(n11206), .B(n11207), .Z(n11178) );
  NANDN U11503 ( .A(n11149), .B(n11148), .Z(n11153) );
  OR U11504 ( .A(n11151), .B(n11150), .Z(n11152) );
  AND U11505 ( .A(n11153), .B(n11152), .Z(n11177) );
  XNOR U11506 ( .A(n11178), .B(n11177), .Z(n11179) );
  XOR U11507 ( .A(n11180), .B(n11179), .Z(n11238) );
  NANDN U11508 ( .A(n11155), .B(n11154), .Z(n11159) );
  NANDN U11509 ( .A(n11157), .B(n11156), .Z(n11158) );
  AND U11510 ( .A(n11159), .B(n11158), .Z(n11237) );
  XNOR U11511 ( .A(n11238), .B(n11237), .Z(n11239) );
  XOR U11512 ( .A(n11240), .B(n11239), .Z(n11172) );
  NANDN U11513 ( .A(n11161), .B(n11160), .Z(n11165) );
  NAND U11514 ( .A(n11163), .B(n11162), .Z(n11164) );
  AND U11515 ( .A(n11165), .B(n11164), .Z(n11171) );
  XNOR U11516 ( .A(n11172), .B(n11171), .Z(n11173) );
  XNOR U11517 ( .A(n11174), .B(n11173), .Z(n11243) );
  XNOR U11518 ( .A(sreg[392]), .B(n11243), .Z(n11245) );
  NANDN U11519 ( .A(sreg[391]), .B(n11166), .Z(n11170) );
  NAND U11520 ( .A(n11168), .B(n11167), .Z(n11169) );
  NAND U11521 ( .A(n11170), .B(n11169), .Z(n11244) );
  XNOR U11522 ( .A(n11245), .B(n11244), .Z(c[392]) );
  NANDN U11523 ( .A(n11172), .B(n11171), .Z(n11176) );
  NANDN U11524 ( .A(n11174), .B(n11173), .Z(n11175) );
  AND U11525 ( .A(n11176), .B(n11175), .Z(n11251) );
  NANDN U11526 ( .A(n11178), .B(n11177), .Z(n11182) );
  NAND U11527 ( .A(n11180), .B(n11179), .Z(n11181) );
  AND U11528 ( .A(n11182), .B(n11181), .Z(n11317) );
  NANDN U11529 ( .A(n11184), .B(n11183), .Z(n11188) );
  NANDN U11530 ( .A(n11186), .B(n11185), .Z(n11187) );
  AND U11531 ( .A(n11188), .B(n11187), .Z(n11283) );
  NAND U11532 ( .A(b[0]), .B(a[153]), .Z(n11189) );
  XNOR U11533 ( .A(b[1]), .B(n11189), .Z(n11191) );
  NANDN U11534 ( .A(b[0]), .B(a[152]), .Z(n11190) );
  NAND U11535 ( .A(n11191), .B(n11190), .Z(n11263) );
  NAND U11536 ( .A(n19808), .B(n11192), .Z(n11194) );
  XOR U11537 ( .A(b[13]), .B(a[141]), .Z(n11266) );
  NAND U11538 ( .A(n19768), .B(n11266), .Z(n11193) );
  AND U11539 ( .A(n11194), .B(n11193), .Z(n11261) );
  AND U11540 ( .A(b[15]), .B(a[137]), .Z(n11260) );
  XNOR U11541 ( .A(n11261), .B(n11260), .Z(n11262) );
  XNOR U11542 ( .A(n11263), .B(n11262), .Z(n11281) );
  NAND U11543 ( .A(n33), .B(n11195), .Z(n11197) );
  XOR U11544 ( .A(b[5]), .B(a[149]), .Z(n11272) );
  NAND U11545 ( .A(n19342), .B(n11272), .Z(n11196) );
  AND U11546 ( .A(n11197), .B(n11196), .Z(n11305) );
  NAND U11547 ( .A(n34), .B(n11198), .Z(n11200) );
  XOR U11548 ( .A(b[7]), .B(a[147]), .Z(n11275) );
  NAND U11549 ( .A(n19486), .B(n11275), .Z(n11199) );
  AND U11550 ( .A(n11200), .B(n11199), .Z(n11303) );
  NAND U11551 ( .A(n31), .B(n11201), .Z(n11203) );
  XOR U11552 ( .A(b[3]), .B(a[151]), .Z(n11278) );
  NAND U11553 ( .A(n32), .B(n11278), .Z(n11202) );
  NAND U11554 ( .A(n11203), .B(n11202), .Z(n11302) );
  XNOR U11555 ( .A(n11303), .B(n11302), .Z(n11304) );
  XOR U11556 ( .A(n11305), .B(n11304), .Z(n11282) );
  XOR U11557 ( .A(n11281), .B(n11282), .Z(n11284) );
  XOR U11558 ( .A(n11283), .B(n11284), .Z(n11255) );
  NANDN U11559 ( .A(n11205), .B(n11204), .Z(n11209) );
  OR U11560 ( .A(n11207), .B(n11206), .Z(n11208) );
  AND U11561 ( .A(n11209), .B(n11208), .Z(n11254) );
  XNOR U11562 ( .A(n11255), .B(n11254), .Z(n11257) );
  NAND U11563 ( .A(n11210), .B(n19724), .Z(n11212) );
  XOR U11564 ( .A(b[11]), .B(a[143]), .Z(n11287) );
  NAND U11565 ( .A(n19692), .B(n11287), .Z(n11211) );
  AND U11566 ( .A(n11212), .B(n11211), .Z(n11298) );
  NAND U11567 ( .A(n19838), .B(n11213), .Z(n11215) );
  XOR U11568 ( .A(b[15]), .B(a[139]), .Z(n11290) );
  NAND U11569 ( .A(n19805), .B(n11290), .Z(n11214) );
  AND U11570 ( .A(n11215), .B(n11214), .Z(n11297) );
  NAND U11571 ( .A(n35), .B(n11216), .Z(n11218) );
  XOR U11572 ( .A(b[9]), .B(a[145]), .Z(n11293) );
  NAND U11573 ( .A(n19598), .B(n11293), .Z(n11217) );
  NAND U11574 ( .A(n11218), .B(n11217), .Z(n11296) );
  XOR U11575 ( .A(n11297), .B(n11296), .Z(n11299) );
  XOR U11576 ( .A(n11298), .B(n11299), .Z(n11309) );
  NANDN U11577 ( .A(n11220), .B(n11219), .Z(n11224) );
  OR U11578 ( .A(n11222), .B(n11221), .Z(n11223) );
  AND U11579 ( .A(n11224), .B(n11223), .Z(n11308) );
  XNOR U11580 ( .A(n11309), .B(n11308), .Z(n11310) );
  NANDN U11581 ( .A(n11226), .B(n11225), .Z(n11230) );
  NANDN U11582 ( .A(n11228), .B(n11227), .Z(n11229) );
  NAND U11583 ( .A(n11230), .B(n11229), .Z(n11311) );
  XNOR U11584 ( .A(n11310), .B(n11311), .Z(n11256) );
  XOR U11585 ( .A(n11257), .B(n11256), .Z(n11315) );
  NANDN U11586 ( .A(n11232), .B(n11231), .Z(n11236) );
  NANDN U11587 ( .A(n11234), .B(n11233), .Z(n11235) );
  AND U11588 ( .A(n11236), .B(n11235), .Z(n11314) );
  XNOR U11589 ( .A(n11315), .B(n11314), .Z(n11316) );
  XOR U11590 ( .A(n11317), .B(n11316), .Z(n11249) );
  NANDN U11591 ( .A(n11238), .B(n11237), .Z(n11242) );
  NAND U11592 ( .A(n11240), .B(n11239), .Z(n11241) );
  AND U11593 ( .A(n11242), .B(n11241), .Z(n11248) );
  XNOR U11594 ( .A(n11249), .B(n11248), .Z(n11250) );
  XNOR U11595 ( .A(n11251), .B(n11250), .Z(n11320) );
  XNOR U11596 ( .A(sreg[393]), .B(n11320), .Z(n11322) );
  NANDN U11597 ( .A(sreg[392]), .B(n11243), .Z(n11247) );
  NAND U11598 ( .A(n11245), .B(n11244), .Z(n11246) );
  NAND U11599 ( .A(n11247), .B(n11246), .Z(n11321) );
  XNOR U11600 ( .A(n11322), .B(n11321), .Z(c[393]) );
  NANDN U11601 ( .A(n11249), .B(n11248), .Z(n11253) );
  NANDN U11602 ( .A(n11251), .B(n11250), .Z(n11252) );
  AND U11603 ( .A(n11253), .B(n11252), .Z(n11328) );
  NANDN U11604 ( .A(n11255), .B(n11254), .Z(n11259) );
  NAND U11605 ( .A(n11257), .B(n11256), .Z(n11258) );
  AND U11606 ( .A(n11259), .B(n11258), .Z(n11394) );
  NANDN U11607 ( .A(n11261), .B(n11260), .Z(n11265) );
  NANDN U11608 ( .A(n11263), .B(n11262), .Z(n11264) );
  AND U11609 ( .A(n11265), .B(n11264), .Z(n11360) );
  NAND U11610 ( .A(n19808), .B(n11266), .Z(n11268) );
  XOR U11611 ( .A(b[13]), .B(a[142]), .Z(n11346) );
  NAND U11612 ( .A(n19768), .B(n11346), .Z(n11267) );
  AND U11613 ( .A(n11268), .B(n11267), .Z(n11338) );
  AND U11614 ( .A(b[15]), .B(a[138]), .Z(n11337) );
  XNOR U11615 ( .A(n11338), .B(n11337), .Z(n11339) );
  NAND U11616 ( .A(b[0]), .B(a[154]), .Z(n11269) );
  XNOR U11617 ( .A(b[1]), .B(n11269), .Z(n11271) );
  NANDN U11618 ( .A(b[0]), .B(a[153]), .Z(n11270) );
  NAND U11619 ( .A(n11271), .B(n11270), .Z(n11340) );
  XNOR U11620 ( .A(n11339), .B(n11340), .Z(n11358) );
  NAND U11621 ( .A(n33), .B(n11272), .Z(n11274) );
  XOR U11622 ( .A(b[5]), .B(a[150]), .Z(n11349) );
  NAND U11623 ( .A(n19342), .B(n11349), .Z(n11273) );
  AND U11624 ( .A(n11274), .B(n11273), .Z(n11382) );
  NAND U11625 ( .A(n34), .B(n11275), .Z(n11277) );
  XOR U11626 ( .A(b[7]), .B(a[148]), .Z(n11352) );
  NAND U11627 ( .A(n19486), .B(n11352), .Z(n11276) );
  AND U11628 ( .A(n11277), .B(n11276), .Z(n11380) );
  NAND U11629 ( .A(n31), .B(n11278), .Z(n11280) );
  XOR U11630 ( .A(b[3]), .B(a[152]), .Z(n11355) );
  NAND U11631 ( .A(n32), .B(n11355), .Z(n11279) );
  NAND U11632 ( .A(n11280), .B(n11279), .Z(n11379) );
  XNOR U11633 ( .A(n11380), .B(n11379), .Z(n11381) );
  XOR U11634 ( .A(n11382), .B(n11381), .Z(n11359) );
  XOR U11635 ( .A(n11358), .B(n11359), .Z(n11361) );
  XOR U11636 ( .A(n11360), .B(n11361), .Z(n11332) );
  NANDN U11637 ( .A(n11282), .B(n11281), .Z(n11286) );
  OR U11638 ( .A(n11284), .B(n11283), .Z(n11285) );
  AND U11639 ( .A(n11286), .B(n11285), .Z(n11331) );
  XNOR U11640 ( .A(n11332), .B(n11331), .Z(n11334) );
  NAND U11641 ( .A(n11287), .B(n19724), .Z(n11289) );
  XOR U11642 ( .A(b[11]), .B(a[144]), .Z(n11364) );
  NAND U11643 ( .A(n19692), .B(n11364), .Z(n11288) );
  AND U11644 ( .A(n11289), .B(n11288), .Z(n11375) );
  NAND U11645 ( .A(n19838), .B(n11290), .Z(n11292) );
  XOR U11646 ( .A(b[15]), .B(a[140]), .Z(n11367) );
  NAND U11647 ( .A(n19805), .B(n11367), .Z(n11291) );
  AND U11648 ( .A(n11292), .B(n11291), .Z(n11374) );
  NAND U11649 ( .A(n35), .B(n11293), .Z(n11295) );
  XOR U11650 ( .A(b[9]), .B(a[146]), .Z(n11370) );
  NAND U11651 ( .A(n19598), .B(n11370), .Z(n11294) );
  NAND U11652 ( .A(n11295), .B(n11294), .Z(n11373) );
  XOR U11653 ( .A(n11374), .B(n11373), .Z(n11376) );
  XOR U11654 ( .A(n11375), .B(n11376), .Z(n11386) );
  NANDN U11655 ( .A(n11297), .B(n11296), .Z(n11301) );
  OR U11656 ( .A(n11299), .B(n11298), .Z(n11300) );
  AND U11657 ( .A(n11301), .B(n11300), .Z(n11385) );
  XNOR U11658 ( .A(n11386), .B(n11385), .Z(n11387) );
  NANDN U11659 ( .A(n11303), .B(n11302), .Z(n11307) );
  NANDN U11660 ( .A(n11305), .B(n11304), .Z(n11306) );
  NAND U11661 ( .A(n11307), .B(n11306), .Z(n11388) );
  XNOR U11662 ( .A(n11387), .B(n11388), .Z(n11333) );
  XOR U11663 ( .A(n11334), .B(n11333), .Z(n11392) );
  NANDN U11664 ( .A(n11309), .B(n11308), .Z(n11313) );
  NANDN U11665 ( .A(n11311), .B(n11310), .Z(n11312) );
  AND U11666 ( .A(n11313), .B(n11312), .Z(n11391) );
  XNOR U11667 ( .A(n11392), .B(n11391), .Z(n11393) );
  XOR U11668 ( .A(n11394), .B(n11393), .Z(n11326) );
  NANDN U11669 ( .A(n11315), .B(n11314), .Z(n11319) );
  NAND U11670 ( .A(n11317), .B(n11316), .Z(n11318) );
  AND U11671 ( .A(n11319), .B(n11318), .Z(n11325) );
  XNOR U11672 ( .A(n11326), .B(n11325), .Z(n11327) );
  XNOR U11673 ( .A(n11328), .B(n11327), .Z(n11397) );
  XNOR U11674 ( .A(sreg[394]), .B(n11397), .Z(n11399) );
  NANDN U11675 ( .A(sreg[393]), .B(n11320), .Z(n11324) );
  NAND U11676 ( .A(n11322), .B(n11321), .Z(n11323) );
  NAND U11677 ( .A(n11324), .B(n11323), .Z(n11398) );
  XNOR U11678 ( .A(n11399), .B(n11398), .Z(c[394]) );
  NANDN U11679 ( .A(n11326), .B(n11325), .Z(n11330) );
  NANDN U11680 ( .A(n11328), .B(n11327), .Z(n11329) );
  AND U11681 ( .A(n11330), .B(n11329), .Z(n11405) );
  NANDN U11682 ( .A(n11332), .B(n11331), .Z(n11336) );
  NAND U11683 ( .A(n11334), .B(n11333), .Z(n11335) );
  AND U11684 ( .A(n11336), .B(n11335), .Z(n11471) );
  NANDN U11685 ( .A(n11338), .B(n11337), .Z(n11342) );
  NANDN U11686 ( .A(n11340), .B(n11339), .Z(n11341) );
  AND U11687 ( .A(n11342), .B(n11341), .Z(n11437) );
  NAND U11688 ( .A(b[0]), .B(a[155]), .Z(n11343) );
  XNOR U11689 ( .A(b[1]), .B(n11343), .Z(n11345) );
  NANDN U11690 ( .A(b[0]), .B(a[154]), .Z(n11344) );
  NAND U11691 ( .A(n11345), .B(n11344), .Z(n11417) );
  NAND U11692 ( .A(n19808), .B(n11346), .Z(n11348) );
  XOR U11693 ( .A(b[13]), .B(a[143]), .Z(n11420) );
  NAND U11694 ( .A(n19768), .B(n11420), .Z(n11347) );
  AND U11695 ( .A(n11348), .B(n11347), .Z(n11415) );
  AND U11696 ( .A(b[15]), .B(a[139]), .Z(n11414) );
  XNOR U11697 ( .A(n11415), .B(n11414), .Z(n11416) );
  XNOR U11698 ( .A(n11417), .B(n11416), .Z(n11435) );
  NAND U11699 ( .A(n33), .B(n11349), .Z(n11351) );
  XOR U11700 ( .A(b[5]), .B(a[151]), .Z(n11426) );
  NAND U11701 ( .A(n19342), .B(n11426), .Z(n11350) );
  AND U11702 ( .A(n11351), .B(n11350), .Z(n11459) );
  NAND U11703 ( .A(n34), .B(n11352), .Z(n11354) );
  XOR U11704 ( .A(b[7]), .B(a[149]), .Z(n11429) );
  NAND U11705 ( .A(n19486), .B(n11429), .Z(n11353) );
  AND U11706 ( .A(n11354), .B(n11353), .Z(n11457) );
  NAND U11707 ( .A(n31), .B(n11355), .Z(n11357) );
  XOR U11708 ( .A(b[3]), .B(a[153]), .Z(n11432) );
  NAND U11709 ( .A(n32), .B(n11432), .Z(n11356) );
  NAND U11710 ( .A(n11357), .B(n11356), .Z(n11456) );
  XNOR U11711 ( .A(n11457), .B(n11456), .Z(n11458) );
  XOR U11712 ( .A(n11459), .B(n11458), .Z(n11436) );
  XOR U11713 ( .A(n11435), .B(n11436), .Z(n11438) );
  XOR U11714 ( .A(n11437), .B(n11438), .Z(n11409) );
  NANDN U11715 ( .A(n11359), .B(n11358), .Z(n11363) );
  OR U11716 ( .A(n11361), .B(n11360), .Z(n11362) );
  AND U11717 ( .A(n11363), .B(n11362), .Z(n11408) );
  XNOR U11718 ( .A(n11409), .B(n11408), .Z(n11411) );
  NAND U11719 ( .A(n11364), .B(n19724), .Z(n11366) );
  XOR U11720 ( .A(b[11]), .B(a[145]), .Z(n11441) );
  NAND U11721 ( .A(n19692), .B(n11441), .Z(n11365) );
  AND U11722 ( .A(n11366), .B(n11365), .Z(n11452) );
  NAND U11723 ( .A(n19838), .B(n11367), .Z(n11369) );
  XOR U11724 ( .A(b[15]), .B(a[141]), .Z(n11444) );
  NAND U11725 ( .A(n19805), .B(n11444), .Z(n11368) );
  AND U11726 ( .A(n11369), .B(n11368), .Z(n11451) );
  NAND U11727 ( .A(n35), .B(n11370), .Z(n11372) );
  XOR U11728 ( .A(b[9]), .B(a[147]), .Z(n11447) );
  NAND U11729 ( .A(n19598), .B(n11447), .Z(n11371) );
  NAND U11730 ( .A(n11372), .B(n11371), .Z(n11450) );
  XOR U11731 ( .A(n11451), .B(n11450), .Z(n11453) );
  XOR U11732 ( .A(n11452), .B(n11453), .Z(n11463) );
  NANDN U11733 ( .A(n11374), .B(n11373), .Z(n11378) );
  OR U11734 ( .A(n11376), .B(n11375), .Z(n11377) );
  AND U11735 ( .A(n11378), .B(n11377), .Z(n11462) );
  XNOR U11736 ( .A(n11463), .B(n11462), .Z(n11464) );
  NANDN U11737 ( .A(n11380), .B(n11379), .Z(n11384) );
  NANDN U11738 ( .A(n11382), .B(n11381), .Z(n11383) );
  NAND U11739 ( .A(n11384), .B(n11383), .Z(n11465) );
  XNOR U11740 ( .A(n11464), .B(n11465), .Z(n11410) );
  XOR U11741 ( .A(n11411), .B(n11410), .Z(n11469) );
  NANDN U11742 ( .A(n11386), .B(n11385), .Z(n11390) );
  NANDN U11743 ( .A(n11388), .B(n11387), .Z(n11389) );
  AND U11744 ( .A(n11390), .B(n11389), .Z(n11468) );
  XNOR U11745 ( .A(n11469), .B(n11468), .Z(n11470) );
  XOR U11746 ( .A(n11471), .B(n11470), .Z(n11403) );
  NANDN U11747 ( .A(n11392), .B(n11391), .Z(n11396) );
  NAND U11748 ( .A(n11394), .B(n11393), .Z(n11395) );
  AND U11749 ( .A(n11396), .B(n11395), .Z(n11402) );
  XNOR U11750 ( .A(n11403), .B(n11402), .Z(n11404) );
  XNOR U11751 ( .A(n11405), .B(n11404), .Z(n11474) );
  XNOR U11752 ( .A(sreg[395]), .B(n11474), .Z(n11476) );
  NANDN U11753 ( .A(sreg[394]), .B(n11397), .Z(n11401) );
  NAND U11754 ( .A(n11399), .B(n11398), .Z(n11400) );
  NAND U11755 ( .A(n11401), .B(n11400), .Z(n11475) );
  XNOR U11756 ( .A(n11476), .B(n11475), .Z(c[395]) );
  NANDN U11757 ( .A(n11403), .B(n11402), .Z(n11407) );
  NANDN U11758 ( .A(n11405), .B(n11404), .Z(n11406) );
  AND U11759 ( .A(n11407), .B(n11406), .Z(n11482) );
  NANDN U11760 ( .A(n11409), .B(n11408), .Z(n11413) );
  NAND U11761 ( .A(n11411), .B(n11410), .Z(n11412) );
  AND U11762 ( .A(n11413), .B(n11412), .Z(n11548) );
  NANDN U11763 ( .A(n11415), .B(n11414), .Z(n11419) );
  NANDN U11764 ( .A(n11417), .B(n11416), .Z(n11418) );
  AND U11765 ( .A(n11419), .B(n11418), .Z(n11514) );
  NAND U11766 ( .A(n19808), .B(n11420), .Z(n11422) );
  XOR U11767 ( .A(b[13]), .B(a[144]), .Z(n11500) );
  NAND U11768 ( .A(n19768), .B(n11500), .Z(n11421) );
  AND U11769 ( .A(n11422), .B(n11421), .Z(n11492) );
  AND U11770 ( .A(b[15]), .B(a[140]), .Z(n11491) );
  XNOR U11771 ( .A(n11492), .B(n11491), .Z(n11493) );
  NAND U11772 ( .A(b[0]), .B(a[156]), .Z(n11423) );
  XNOR U11773 ( .A(b[1]), .B(n11423), .Z(n11425) );
  NANDN U11774 ( .A(b[0]), .B(a[155]), .Z(n11424) );
  NAND U11775 ( .A(n11425), .B(n11424), .Z(n11494) );
  XNOR U11776 ( .A(n11493), .B(n11494), .Z(n11512) );
  NAND U11777 ( .A(n33), .B(n11426), .Z(n11428) );
  XOR U11778 ( .A(b[5]), .B(a[152]), .Z(n11503) );
  NAND U11779 ( .A(n19342), .B(n11503), .Z(n11427) );
  AND U11780 ( .A(n11428), .B(n11427), .Z(n11536) );
  NAND U11781 ( .A(n34), .B(n11429), .Z(n11431) );
  XOR U11782 ( .A(b[7]), .B(a[150]), .Z(n11506) );
  NAND U11783 ( .A(n19486), .B(n11506), .Z(n11430) );
  AND U11784 ( .A(n11431), .B(n11430), .Z(n11534) );
  NAND U11785 ( .A(n31), .B(n11432), .Z(n11434) );
  XOR U11786 ( .A(b[3]), .B(a[154]), .Z(n11509) );
  NAND U11787 ( .A(n32), .B(n11509), .Z(n11433) );
  NAND U11788 ( .A(n11434), .B(n11433), .Z(n11533) );
  XNOR U11789 ( .A(n11534), .B(n11533), .Z(n11535) );
  XOR U11790 ( .A(n11536), .B(n11535), .Z(n11513) );
  XOR U11791 ( .A(n11512), .B(n11513), .Z(n11515) );
  XOR U11792 ( .A(n11514), .B(n11515), .Z(n11486) );
  NANDN U11793 ( .A(n11436), .B(n11435), .Z(n11440) );
  OR U11794 ( .A(n11438), .B(n11437), .Z(n11439) );
  AND U11795 ( .A(n11440), .B(n11439), .Z(n11485) );
  XNOR U11796 ( .A(n11486), .B(n11485), .Z(n11488) );
  NAND U11797 ( .A(n11441), .B(n19724), .Z(n11443) );
  XOR U11798 ( .A(b[11]), .B(a[146]), .Z(n11518) );
  NAND U11799 ( .A(n19692), .B(n11518), .Z(n11442) );
  AND U11800 ( .A(n11443), .B(n11442), .Z(n11529) );
  NAND U11801 ( .A(n19838), .B(n11444), .Z(n11446) );
  XOR U11802 ( .A(b[15]), .B(a[142]), .Z(n11521) );
  NAND U11803 ( .A(n19805), .B(n11521), .Z(n11445) );
  AND U11804 ( .A(n11446), .B(n11445), .Z(n11528) );
  NAND U11805 ( .A(n35), .B(n11447), .Z(n11449) );
  XOR U11806 ( .A(b[9]), .B(a[148]), .Z(n11524) );
  NAND U11807 ( .A(n19598), .B(n11524), .Z(n11448) );
  NAND U11808 ( .A(n11449), .B(n11448), .Z(n11527) );
  XOR U11809 ( .A(n11528), .B(n11527), .Z(n11530) );
  XOR U11810 ( .A(n11529), .B(n11530), .Z(n11540) );
  NANDN U11811 ( .A(n11451), .B(n11450), .Z(n11455) );
  OR U11812 ( .A(n11453), .B(n11452), .Z(n11454) );
  AND U11813 ( .A(n11455), .B(n11454), .Z(n11539) );
  XNOR U11814 ( .A(n11540), .B(n11539), .Z(n11541) );
  NANDN U11815 ( .A(n11457), .B(n11456), .Z(n11461) );
  NANDN U11816 ( .A(n11459), .B(n11458), .Z(n11460) );
  NAND U11817 ( .A(n11461), .B(n11460), .Z(n11542) );
  XNOR U11818 ( .A(n11541), .B(n11542), .Z(n11487) );
  XOR U11819 ( .A(n11488), .B(n11487), .Z(n11546) );
  NANDN U11820 ( .A(n11463), .B(n11462), .Z(n11467) );
  NANDN U11821 ( .A(n11465), .B(n11464), .Z(n11466) );
  AND U11822 ( .A(n11467), .B(n11466), .Z(n11545) );
  XNOR U11823 ( .A(n11546), .B(n11545), .Z(n11547) );
  XOR U11824 ( .A(n11548), .B(n11547), .Z(n11480) );
  NANDN U11825 ( .A(n11469), .B(n11468), .Z(n11473) );
  NAND U11826 ( .A(n11471), .B(n11470), .Z(n11472) );
  AND U11827 ( .A(n11473), .B(n11472), .Z(n11479) );
  XNOR U11828 ( .A(n11480), .B(n11479), .Z(n11481) );
  XNOR U11829 ( .A(n11482), .B(n11481), .Z(n11551) );
  XNOR U11830 ( .A(sreg[396]), .B(n11551), .Z(n11553) );
  NANDN U11831 ( .A(sreg[395]), .B(n11474), .Z(n11478) );
  NAND U11832 ( .A(n11476), .B(n11475), .Z(n11477) );
  NAND U11833 ( .A(n11478), .B(n11477), .Z(n11552) );
  XNOR U11834 ( .A(n11553), .B(n11552), .Z(c[396]) );
  NANDN U11835 ( .A(n11480), .B(n11479), .Z(n11484) );
  NANDN U11836 ( .A(n11482), .B(n11481), .Z(n11483) );
  AND U11837 ( .A(n11484), .B(n11483), .Z(n11559) );
  NANDN U11838 ( .A(n11486), .B(n11485), .Z(n11490) );
  NAND U11839 ( .A(n11488), .B(n11487), .Z(n11489) );
  AND U11840 ( .A(n11490), .B(n11489), .Z(n11625) );
  NANDN U11841 ( .A(n11492), .B(n11491), .Z(n11496) );
  NANDN U11842 ( .A(n11494), .B(n11493), .Z(n11495) );
  AND U11843 ( .A(n11496), .B(n11495), .Z(n11591) );
  NAND U11844 ( .A(b[0]), .B(a[157]), .Z(n11497) );
  XNOR U11845 ( .A(b[1]), .B(n11497), .Z(n11499) );
  NANDN U11846 ( .A(b[0]), .B(a[156]), .Z(n11498) );
  NAND U11847 ( .A(n11499), .B(n11498), .Z(n11571) );
  NAND U11848 ( .A(n19808), .B(n11500), .Z(n11502) );
  XOR U11849 ( .A(b[13]), .B(a[145]), .Z(n11577) );
  NAND U11850 ( .A(n19768), .B(n11577), .Z(n11501) );
  AND U11851 ( .A(n11502), .B(n11501), .Z(n11569) );
  AND U11852 ( .A(b[15]), .B(a[141]), .Z(n11568) );
  XNOR U11853 ( .A(n11569), .B(n11568), .Z(n11570) );
  XNOR U11854 ( .A(n11571), .B(n11570), .Z(n11589) );
  NAND U11855 ( .A(n33), .B(n11503), .Z(n11505) );
  XOR U11856 ( .A(b[5]), .B(a[153]), .Z(n11580) );
  NAND U11857 ( .A(n19342), .B(n11580), .Z(n11504) );
  AND U11858 ( .A(n11505), .B(n11504), .Z(n11613) );
  NAND U11859 ( .A(n34), .B(n11506), .Z(n11508) );
  XOR U11860 ( .A(b[7]), .B(a[151]), .Z(n11583) );
  NAND U11861 ( .A(n19486), .B(n11583), .Z(n11507) );
  AND U11862 ( .A(n11508), .B(n11507), .Z(n11611) );
  NAND U11863 ( .A(n31), .B(n11509), .Z(n11511) );
  XOR U11864 ( .A(b[3]), .B(a[155]), .Z(n11586) );
  NAND U11865 ( .A(n32), .B(n11586), .Z(n11510) );
  NAND U11866 ( .A(n11511), .B(n11510), .Z(n11610) );
  XNOR U11867 ( .A(n11611), .B(n11610), .Z(n11612) );
  XOR U11868 ( .A(n11613), .B(n11612), .Z(n11590) );
  XOR U11869 ( .A(n11589), .B(n11590), .Z(n11592) );
  XOR U11870 ( .A(n11591), .B(n11592), .Z(n11563) );
  NANDN U11871 ( .A(n11513), .B(n11512), .Z(n11517) );
  OR U11872 ( .A(n11515), .B(n11514), .Z(n11516) );
  AND U11873 ( .A(n11517), .B(n11516), .Z(n11562) );
  XNOR U11874 ( .A(n11563), .B(n11562), .Z(n11565) );
  NAND U11875 ( .A(n11518), .B(n19724), .Z(n11520) );
  XOR U11876 ( .A(b[11]), .B(a[147]), .Z(n11595) );
  NAND U11877 ( .A(n19692), .B(n11595), .Z(n11519) );
  AND U11878 ( .A(n11520), .B(n11519), .Z(n11606) );
  NAND U11879 ( .A(n19838), .B(n11521), .Z(n11523) );
  XOR U11880 ( .A(b[15]), .B(a[143]), .Z(n11598) );
  NAND U11881 ( .A(n19805), .B(n11598), .Z(n11522) );
  AND U11882 ( .A(n11523), .B(n11522), .Z(n11605) );
  NAND U11883 ( .A(n35), .B(n11524), .Z(n11526) );
  XOR U11884 ( .A(b[9]), .B(a[149]), .Z(n11601) );
  NAND U11885 ( .A(n19598), .B(n11601), .Z(n11525) );
  NAND U11886 ( .A(n11526), .B(n11525), .Z(n11604) );
  XOR U11887 ( .A(n11605), .B(n11604), .Z(n11607) );
  XOR U11888 ( .A(n11606), .B(n11607), .Z(n11617) );
  NANDN U11889 ( .A(n11528), .B(n11527), .Z(n11532) );
  OR U11890 ( .A(n11530), .B(n11529), .Z(n11531) );
  AND U11891 ( .A(n11532), .B(n11531), .Z(n11616) );
  XNOR U11892 ( .A(n11617), .B(n11616), .Z(n11618) );
  NANDN U11893 ( .A(n11534), .B(n11533), .Z(n11538) );
  NANDN U11894 ( .A(n11536), .B(n11535), .Z(n11537) );
  NAND U11895 ( .A(n11538), .B(n11537), .Z(n11619) );
  XNOR U11896 ( .A(n11618), .B(n11619), .Z(n11564) );
  XOR U11897 ( .A(n11565), .B(n11564), .Z(n11623) );
  NANDN U11898 ( .A(n11540), .B(n11539), .Z(n11544) );
  NANDN U11899 ( .A(n11542), .B(n11541), .Z(n11543) );
  AND U11900 ( .A(n11544), .B(n11543), .Z(n11622) );
  XNOR U11901 ( .A(n11623), .B(n11622), .Z(n11624) );
  XOR U11902 ( .A(n11625), .B(n11624), .Z(n11557) );
  NANDN U11903 ( .A(n11546), .B(n11545), .Z(n11550) );
  NAND U11904 ( .A(n11548), .B(n11547), .Z(n11549) );
  AND U11905 ( .A(n11550), .B(n11549), .Z(n11556) );
  XNOR U11906 ( .A(n11557), .B(n11556), .Z(n11558) );
  XNOR U11907 ( .A(n11559), .B(n11558), .Z(n11628) );
  XNOR U11908 ( .A(sreg[397]), .B(n11628), .Z(n11630) );
  NANDN U11909 ( .A(sreg[396]), .B(n11551), .Z(n11555) );
  NAND U11910 ( .A(n11553), .B(n11552), .Z(n11554) );
  NAND U11911 ( .A(n11555), .B(n11554), .Z(n11629) );
  XNOR U11912 ( .A(n11630), .B(n11629), .Z(c[397]) );
  NANDN U11913 ( .A(n11557), .B(n11556), .Z(n11561) );
  NANDN U11914 ( .A(n11559), .B(n11558), .Z(n11560) );
  AND U11915 ( .A(n11561), .B(n11560), .Z(n11636) );
  NANDN U11916 ( .A(n11563), .B(n11562), .Z(n11567) );
  NAND U11917 ( .A(n11565), .B(n11564), .Z(n11566) );
  AND U11918 ( .A(n11567), .B(n11566), .Z(n11702) );
  NANDN U11919 ( .A(n11569), .B(n11568), .Z(n11573) );
  NANDN U11920 ( .A(n11571), .B(n11570), .Z(n11572) );
  AND U11921 ( .A(n11573), .B(n11572), .Z(n11668) );
  NAND U11922 ( .A(b[0]), .B(a[158]), .Z(n11574) );
  XNOR U11923 ( .A(b[1]), .B(n11574), .Z(n11576) );
  NANDN U11924 ( .A(b[0]), .B(a[157]), .Z(n11575) );
  NAND U11925 ( .A(n11576), .B(n11575), .Z(n11648) );
  NAND U11926 ( .A(n19808), .B(n11577), .Z(n11579) );
  XOR U11927 ( .A(b[13]), .B(a[146]), .Z(n11651) );
  NAND U11928 ( .A(n19768), .B(n11651), .Z(n11578) );
  AND U11929 ( .A(n11579), .B(n11578), .Z(n11646) );
  AND U11930 ( .A(b[15]), .B(a[142]), .Z(n11645) );
  XNOR U11931 ( .A(n11646), .B(n11645), .Z(n11647) );
  XNOR U11932 ( .A(n11648), .B(n11647), .Z(n11666) );
  NAND U11933 ( .A(n33), .B(n11580), .Z(n11582) );
  XOR U11934 ( .A(b[5]), .B(a[154]), .Z(n11657) );
  NAND U11935 ( .A(n19342), .B(n11657), .Z(n11581) );
  AND U11936 ( .A(n11582), .B(n11581), .Z(n11690) );
  NAND U11937 ( .A(n34), .B(n11583), .Z(n11585) );
  XOR U11938 ( .A(b[7]), .B(a[152]), .Z(n11660) );
  NAND U11939 ( .A(n19486), .B(n11660), .Z(n11584) );
  AND U11940 ( .A(n11585), .B(n11584), .Z(n11688) );
  NAND U11941 ( .A(n31), .B(n11586), .Z(n11588) );
  XOR U11942 ( .A(b[3]), .B(a[156]), .Z(n11663) );
  NAND U11943 ( .A(n32), .B(n11663), .Z(n11587) );
  NAND U11944 ( .A(n11588), .B(n11587), .Z(n11687) );
  XNOR U11945 ( .A(n11688), .B(n11687), .Z(n11689) );
  XOR U11946 ( .A(n11690), .B(n11689), .Z(n11667) );
  XOR U11947 ( .A(n11666), .B(n11667), .Z(n11669) );
  XOR U11948 ( .A(n11668), .B(n11669), .Z(n11640) );
  NANDN U11949 ( .A(n11590), .B(n11589), .Z(n11594) );
  OR U11950 ( .A(n11592), .B(n11591), .Z(n11593) );
  AND U11951 ( .A(n11594), .B(n11593), .Z(n11639) );
  XNOR U11952 ( .A(n11640), .B(n11639), .Z(n11642) );
  NAND U11953 ( .A(n11595), .B(n19724), .Z(n11597) );
  XOR U11954 ( .A(b[11]), .B(a[148]), .Z(n11672) );
  NAND U11955 ( .A(n19692), .B(n11672), .Z(n11596) );
  AND U11956 ( .A(n11597), .B(n11596), .Z(n11683) );
  NAND U11957 ( .A(n19838), .B(n11598), .Z(n11600) );
  XOR U11958 ( .A(b[15]), .B(a[144]), .Z(n11675) );
  NAND U11959 ( .A(n19805), .B(n11675), .Z(n11599) );
  AND U11960 ( .A(n11600), .B(n11599), .Z(n11682) );
  NAND U11961 ( .A(n35), .B(n11601), .Z(n11603) );
  XOR U11962 ( .A(b[9]), .B(a[150]), .Z(n11678) );
  NAND U11963 ( .A(n19598), .B(n11678), .Z(n11602) );
  NAND U11964 ( .A(n11603), .B(n11602), .Z(n11681) );
  XOR U11965 ( .A(n11682), .B(n11681), .Z(n11684) );
  XOR U11966 ( .A(n11683), .B(n11684), .Z(n11694) );
  NANDN U11967 ( .A(n11605), .B(n11604), .Z(n11609) );
  OR U11968 ( .A(n11607), .B(n11606), .Z(n11608) );
  AND U11969 ( .A(n11609), .B(n11608), .Z(n11693) );
  XNOR U11970 ( .A(n11694), .B(n11693), .Z(n11695) );
  NANDN U11971 ( .A(n11611), .B(n11610), .Z(n11615) );
  NANDN U11972 ( .A(n11613), .B(n11612), .Z(n11614) );
  NAND U11973 ( .A(n11615), .B(n11614), .Z(n11696) );
  XNOR U11974 ( .A(n11695), .B(n11696), .Z(n11641) );
  XOR U11975 ( .A(n11642), .B(n11641), .Z(n11700) );
  NANDN U11976 ( .A(n11617), .B(n11616), .Z(n11621) );
  NANDN U11977 ( .A(n11619), .B(n11618), .Z(n11620) );
  AND U11978 ( .A(n11621), .B(n11620), .Z(n11699) );
  XNOR U11979 ( .A(n11700), .B(n11699), .Z(n11701) );
  XOR U11980 ( .A(n11702), .B(n11701), .Z(n11634) );
  NANDN U11981 ( .A(n11623), .B(n11622), .Z(n11627) );
  NAND U11982 ( .A(n11625), .B(n11624), .Z(n11626) );
  AND U11983 ( .A(n11627), .B(n11626), .Z(n11633) );
  XNOR U11984 ( .A(n11634), .B(n11633), .Z(n11635) );
  XNOR U11985 ( .A(n11636), .B(n11635), .Z(n11705) );
  XNOR U11986 ( .A(sreg[398]), .B(n11705), .Z(n11707) );
  NANDN U11987 ( .A(sreg[397]), .B(n11628), .Z(n11632) );
  NAND U11988 ( .A(n11630), .B(n11629), .Z(n11631) );
  NAND U11989 ( .A(n11632), .B(n11631), .Z(n11706) );
  XNOR U11990 ( .A(n11707), .B(n11706), .Z(c[398]) );
  NANDN U11991 ( .A(n11634), .B(n11633), .Z(n11638) );
  NANDN U11992 ( .A(n11636), .B(n11635), .Z(n11637) );
  AND U11993 ( .A(n11638), .B(n11637), .Z(n11713) );
  NANDN U11994 ( .A(n11640), .B(n11639), .Z(n11644) );
  NAND U11995 ( .A(n11642), .B(n11641), .Z(n11643) );
  AND U11996 ( .A(n11644), .B(n11643), .Z(n11779) );
  NANDN U11997 ( .A(n11646), .B(n11645), .Z(n11650) );
  NANDN U11998 ( .A(n11648), .B(n11647), .Z(n11649) );
  AND U11999 ( .A(n11650), .B(n11649), .Z(n11745) );
  NAND U12000 ( .A(n19808), .B(n11651), .Z(n11653) );
  XOR U12001 ( .A(b[13]), .B(a[147]), .Z(n11731) );
  NAND U12002 ( .A(n19768), .B(n11731), .Z(n11652) );
  AND U12003 ( .A(n11653), .B(n11652), .Z(n11723) );
  AND U12004 ( .A(b[15]), .B(a[143]), .Z(n11722) );
  XNOR U12005 ( .A(n11723), .B(n11722), .Z(n11724) );
  NAND U12006 ( .A(b[0]), .B(a[159]), .Z(n11654) );
  XNOR U12007 ( .A(b[1]), .B(n11654), .Z(n11656) );
  NANDN U12008 ( .A(b[0]), .B(a[158]), .Z(n11655) );
  NAND U12009 ( .A(n11656), .B(n11655), .Z(n11725) );
  XNOR U12010 ( .A(n11724), .B(n11725), .Z(n11743) );
  NAND U12011 ( .A(n33), .B(n11657), .Z(n11659) );
  XOR U12012 ( .A(b[5]), .B(a[155]), .Z(n11734) );
  NAND U12013 ( .A(n19342), .B(n11734), .Z(n11658) );
  AND U12014 ( .A(n11659), .B(n11658), .Z(n11767) );
  NAND U12015 ( .A(n34), .B(n11660), .Z(n11662) );
  XOR U12016 ( .A(b[7]), .B(a[153]), .Z(n11737) );
  NAND U12017 ( .A(n19486), .B(n11737), .Z(n11661) );
  AND U12018 ( .A(n11662), .B(n11661), .Z(n11765) );
  NAND U12019 ( .A(n31), .B(n11663), .Z(n11665) );
  XOR U12020 ( .A(b[3]), .B(a[157]), .Z(n11740) );
  NAND U12021 ( .A(n32), .B(n11740), .Z(n11664) );
  NAND U12022 ( .A(n11665), .B(n11664), .Z(n11764) );
  XNOR U12023 ( .A(n11765), .B(n11764), .Z(n11766) );
  XOR U12024 ( .A(n11767), .B(n11766), .Z(n11744) );
  XOR U12025 ( .A(n11743), .B(n11744), .Z(n11746) );
  XOR U12026 ( .A(n11745), .B(n11746), .Z(n11717) );
  NANDN U12027 ( .A(n11667), .B(n11666), .Z(n11671) );
  OR U12028 ( .A(n11669), .B(n11668), .Z(n11670) );
  AND U12029 ( .A(n11671), .B(n11670), .Z(n11716) );
  XNOR U12030 ( .A(n11717), .B(n11716), .Z(n11719) );
  NAND U12031 ( .A(n11672), .B(n19724), .Z(n11674) );
  XOR U12032 ( .A(b[11]), .B(a[149]), .Z(n11749) );
  NAND U12033 ( .A(n19692), .B(n11749), .Z(n11673) );
  AND U12034 ( .A(n11674), .B(n11673), .Z(n11760) );
  NAND U12035 ( .A(n19838), .B(n11675), .Z(n11677) );
  XOR U12036 ( .A(b[15]), .B(a[145]), .Z(n11752) );
  NAND U12037 ( .A(n19805), .B(n11752), .Z(n11676) );
  AND U12038 ( .A(n11677), .B(n11676), .Z(n11759) );
  NAND U12039 ( .A(n35), .B(n11678), .Z(n11680) );
  XOR U12040 ( .A(b[9]), .B(a[151]), .Z(n11755) );
  NAND U12041 ( .A(n19598), .B(n11755), .Z(n11679) );
  NAND U12042 ( .A(n11680), .B(n11679), .Z(n11758) );
  XOR U12043 ( .A(n11759), .B(n11758), .Z(n11761) );
  XOR U12044 ( .A(n11760), .B(n11761), .Z(n11771) );
  NANDN U12045 ( .A(n11682), .B(n11681), .Z(n11686) );
  OR U12046 ( .A(n11684), .B(n11683), .Z(n11685) );
  AND U12047 ( .A(n11686), .B(n11685), .Z(n11770) );
  XNOR U12048 ( .A(n11771), .B(n11770), .Z(n11772) );
  NANDN U12049 ( .A(n11688), .B(n11687), .Z(n11692) );
  NANDN U12050 ( .A(n11690), .B(n11689), .Z(n11691) );
  NAND U12051 ( .A(n11692), .B(n11691), .Z(n11773) );
  XNOR U12052 ( .A(n11772), .B(n11773), .Z(n11718) );
  XOR U12053 ( .A(n11719), .B(n11718), .Z(n11777) );
  NANDN U12054 ( .A(n11694), .B(n11693), .Z(n11698) );
  NANDN U12055 ( .A(n11696), .B(n11695), .Z(n11697) );
  AND U12056 ( .A(n11698), .B(n11697), .Z(n11776) );
  XNOR U12057 ( .A(n11777), .B(n11776), .Z(n11778) );
  XOR U12058 ( .A(n11779), .B(n11778), .Z(n11711) );
  NANDN U12059 ( .A(n11700), .B(n11699), .Z(n11704) );
  NAND U12060 ( .A(n11702), .B(n11701), .Z(n11703) );
  AND U12061 ( .A(n11704), .B(n11703), .Z(n11710) );
  XNOR U12062 ( .A(n11711), .B(n11710), .Z(n11712) );
  XNOR U12063 ( .A(n11713), .B(n11712), .Z(n11782) );
  XNOR U12064 ( .A(sreg[399]), .B(n11782), .Z(n11784) );
  NANDN U12065 ( .A(sreg[398]), .B(n11705), .Z(n11709) );
  NAND U12066 ( .A(n11707), .B(n11706), .Z(n11708) );
  NAND U12067 ( .A(n11709), .B(n11708), .Z(n11783) );
  XNOR U12068 ( .A(n11784), .B(n11783), .Z(c[399]) );
  NANDN U12069 ( .A(n11711), .B(n11710), .Z(n11715) );
  NANDN U12070 ( .A(n11713), .B(n11712), .Z(n11714) );
  AND U12071 ( .A(n11715), .B(n11714), .Z(n11790) );
  NANDN U12072 ( .A(n11717), .B(n11716), .Z(n11721) );
  NAND U12073 ( .A(n11719), .B(n11718), .Z(n11720) );
  AND U12074 ( .A(n11721), .B(n11720), .Z(n11856) );
  NANDN U12075 ( .A(n11723), .B(n11722), .Z(n11727) );
  NANDN U12076 ( .A(n11725), .B(n11724), .Z(n11726) );
  AND U12077 ( .A(n11727), .B(n11726), .Z(n11822) );
  NAND U12078 ( .A(b[0]), .B(a[160]), .Z(n11728) );
  XNOR U12079 ( .A(b[1]), .B(n11728), .Z(n11730) );
  NANDN U12080 ( .A(b[0]), .B(a[159]), .Z(n11729) );
  NAND U12081 ( .A(n11730), .B(n11729), .Z(n11802) );
  NAND U12082 ( .A(n19808), .B(n11731), .Z(n11733) );
  XOR U12083 ( .A(b[13]), .B(a[148]), .Z(n11805) );
  NAND U12084 ( .A(n19768), .B(n11805), .Z(n11732) );
  AND U12085 ( .A(n11733), .B(n11732), .Z(n11800) );
  AND U12086 ( .A(b[15]), .B(a[144]), .Z(n11799) );
  XNOR U12087 ( .A(n11800), .B(n11799), .Z(n11801) );
  XNOR U12088 ( .A(n11802), .B(n11801), .Z(n11820) );
  NAND U12089 ( .A(n33), .B(n11734), .Z(n11736) );
  XOR U12090 ( .A(b[5]), .B(a[156]), .Z(n11811) );
  NAND U12091 ( .A(n19342), .B(n11811), .Z(n11735) );
  AND U12092 ( .A(n11736), .B(n11735), .Z(n11844) );
  NAND U12093 ( .A(n34), .B(n11737), .Z(n11739) );
  XOR U12094 ( .A(b[7]), .B(a[154]), .Z(n11814) );
  NAND U12095 ( .A(n19486), .B(n11814), .Z(n11738) );
  AND U12096 ( .A(n11739), .B(n11738), .Z(n11842) );
  NAND U12097 ( .A(n31), .B(n11740), .Z(n11742) );
  XOR U12098 ( .A(b[3]), .B(a[158]), .Z(n11817) );
  NAND U12099 ( .A(n32), .B(n11817), .Z(n11741) );
  NAND U12100 ( .A(n11742), .B(n11741), .Z(n11841) );
  XNOR U12101 ( .A(n11842), .B(n11841), .Z(n11843) );
  XOR U12102 ( .A(n11844), .B(n11843), .Z(n11821) );
  XOR U12103 ( .A(n11820), .B(n11821), .Z(n11823) );
  XOR U12104 ( .A(n11822), .B(n11823), .Z(n11794) );
  NANDN U12105 ( .A(n11744), .B(n11743), .Z(n11748) );
  OR U12106 ( .A(n11746), .B(n11745), .Z(n11747) );
  AND U12107 ( .A(n11748), .B(n11747), .Z(n11793) );
  XNOR U12108 ( .A(n11794), .B(n11793), .Z(n11796) );
  NAND U12109 ( .A(n11749), .B(n19724), .Z(n11751) );
  XOR U12110 ( .A(b[11]), .B(a[150]), .Z(n11826) );
  NAND U12111 ( .A(n19692), .B(n11826), .Z(n11750) );
  AND U12112 ( .A(n11751), .B(n11750), .Z(n11837) );
  NAND U12113 ( .A(n19838), .B(n11752), .Z(n11754) );
  XOR U12114 ( .A(b[15]), .B(a[146]), .Z(n11829) );
  NAND U12115 ( .A(n19805), .B(n11829), .Z(n11753) );
  AND U12116 ( .A(n11754), .B(n11753), .Z(n11836) );
  NAND U12117 ( .A(n35), .B(n11755), .Z(n11757) );
  XOR U12118 ( .A(b[9]), .B(a[152]), .Z(n11832) );
  NAND U12119 ( .A(n19598), .B(n11832), .Z(n11756) );
  NAND U12120 ( .A(n11757), .B(n11756), .Z(n11835) );
  XOR U12121 ( .A(n11836), .B(n11835), .Z(n11838) );
  XOR U12122 ( .A(n11837), .B(n11838), .Z(n11848) );
  NANDN U12123 ( .A(n11759), .B(n11758), .Z(n11763) );
  OR U12124 ( .A(n11761), .B(n11760), .Z(n11762) );
  AND U12125 ( .A(n11763), .B(n11762), .Z(n11847) );
  XNOR U12126 ( .A(n11848), .B(n11847), .Z(n11849) );
  NANDN U12127 ( .A(n11765), .B(n11764), .Z(n11769) );
  NANDN U12128 ( .A(n11767), .B(n11766), .Z(n11768) );
  NAND U12129 ( .A(n11769), .B(n11768), .Z(n11850) );
  XNOR U12130 ( .A(n11849), .B(n11850), .Z(n11795) );
  XOR U12131 ( .A(n11796), .B(n11795), .Z(n11854) );
  NANDN U12132 ( .A(n11771), .B(n11770), .Z(n11775) );
  NANDN U12133 ( .A(n11773), .B(n11772), .Z(n11774) );
  AND U12134 ( .A(n11775), .B(n11774), .Z(n11853) );
  XNOR U12135 ( .A(n11854), .B(n11853), .Z(n11855) );
  XOR U12136 ( .A(n11856), .B(n11855), .Z(n11788) );
  NANDN U12137 ( .A(n11777), .B(n11776), .Z(n11781) );
  NAND U12138 ( .A(n11779), .B(n11778), .Z(n11780) );
  AND U12139 ( .A(n11781), .B(n11780), .Z(n11787) );
  XNOR U12140 ( .A(n11788), .B(n11787), .Z(n11789) );
  XNOR U12141 ( .A(n11790), .B(n11789), .Z(n11859) );
  XNOR U12142 ( .A(sreg[400]), .B(n11859), .Z(n11861) );
  NANDN U12143 ( .A(sreg[399]), .B(n11782), .Z(n11786) );
  NAND U12144 ( .A(n11784), .B(n11783), .Z(n11785) );
  NAND U12145 ( .A(n11786), .B(n11785), .Z(n11860) );
  XNOR U12146 ( .A(n11861), .B(n11860), .Z(c[400]) );
  NANDN U12147 ( .A(n11788), .B(n11787), .Z(n11792) );
  NANDN U12148 ( .A(n11790), .B(n11789), .Z(n11791) );
  AND U12149 ( .A(n11792), .B(n11791), .Z(n11867) );
  NANDN U12150 ( .A(n11794), .B(n11793), .Z(n11798) );
  NAND U12151 ( .A(n11796), .B(n11795), .Z(n11797) );
  AND U12152 ( .A(n11798), .B(n11797), .Z(n11933) );
  NANDN U12153 ( .A(n11800), .B(n11799), .Z(n11804) );
  NANDN U12154 ( .A(n11802), .B(n11801), .Z(n11803) );
  AND U12155 ( .A(n11804), .B(n11803), .Z(n11899) );
  NAND U12156 ( .A(n19808), .B(n11805), .Z(n11807) );
  XOR U12157 ( .A(b[13]), .B(a[149]), .Z(n11885) );
  NAND U12158 ( .A(n19768), .B(n11885), .Z(n11806) );
  AND U12159 ( .A(n11807), .B(n11806), .Z(n11877) );
  AND U12160 ( .A(b[15]), .B(a[145]), .Z(n11876) );
  XNOR U12161 ( .A(n11877), .B(n11876), .Z(n11878) );
  NAND U12162 ( .A(b[0]), .B(a[161]), .Z(n11808) );
  XNOR U12163 ( .A(b[1]), .B(n11808), .Z(n11810) );
  NANDN U12164 ( .A(b[0]), .B(a[160]), .Z(n11809) );
  NAND U12165 ( .A(n11810), .B(n11809), .Z(n11879) );
  XNOR U12166 ( .A(n11878), .B(n11879), .Z(n11897) );
  NAND U12167 ( .A(n33), .B(n11811), .Z(n11813) );
  XOR U12168 ( .A(b[5]), .B(a[157]), .Z(n11888) );
  NAND U12169 ( .A(n19342), .B(n11888), .Z(n11812) );
  AND U12170 ( .A(n11813), .B(n11812), .Z(n11921) );
  NAND U12171 ( .A(n34), .B(n11814), .Z(n11816) );
  XOR U12172 ( .A(b[7]), .B(a[155]), .Z(n11891) );
  NAND U12173 ( .A(n19486), .B(n11891), .Z(n11815) );
  AND U12174 ( .A(n11816), .B(n11815), .Z(n11919) );
  NAND U12175 ( .A(n31), .B(n11817), .Z(n11819) );
  XOR U12176 ( .A(b[3]), .B(a[159]), .Z(n11894) );
  NAND U12177 ( .A(n32), .B(n11894), .Z(n11818) );
  NAND U12178 ( .A(n11819), .B(n11818), .Z(n11918) );
  XNOR U12179 ( .A(n11919), .B(n11918), .Z(n11920) );
  XOR U12180 ( .A(n11921), .B(n11920), .Z(n11898) );
  XOR U12181 ( .A(n11897), .B(n11898), .Z(n11900) );
  XOR U12182 ( .A(n11899), .B(n11900), .Z(n11871) );
  NANDN U12183 ( .A(n11821), .B(n11820), .Z(n11825) );
  OR U12184 ( .A(n11823), .B(n11822), .Z(n11824) );
  AND U12185 ( .A(n11825), .B(n11824), .Z(n11870) );
  XNOR U12186 ( .A(n11871), .B(n11870), .Z(n11873) );
  NAND U12187 ( .A(n11826), .B(n19724), .Z(n11828) );
  XOR U12188 ( .A(b[11]), .B(a[151]), .Z(n11903) );
  NAND U12189 ( .A(n19692), .B(n11903), .Z(n11827) );
  AND U12190 ( .A(n11828), .B(n11827), .Z(n11914) );
  NAND U12191 ( .A(n19838), .B(n11829), .Z(n11831) );
  XOR U12192 ( .A(b[15]), .B(a[147]), .Z(n11906) );
  NAND U12193 ( .A(n19805), .B(n11906), .Z(n11830) );
  AND U12194 ( .A(n11831), .B(n11830), .Z(n11913) );
  NAND U12195 ( .A(n35), .B(n11832), .Z(n11834) );
  XOR U12196 ( .A(b[9]), .B(a[153]), .Z(n11909) );
  NAND U12197 ( .A(n19598), .B(n11909), .Z(n11833) );
  NAND U12198 ( .A(n11834), .B(n11833), .Z(n11912) );
  XOR U12199 ( .A(n11913), .B(n11912), .Z(n11915) );
  XOR U12200 ( .A(n11914), .B(n11915), .Z(n11925) );
  NANDN U12201 ( .A(n11836), .B(n11835), .Z(n11840) );
  OR U12202 ( .A(n11838), .B(n11837), .Z(n11839) );
  AND U12203 ( .A(n11840), .B(n11839), .Z(n11924) );
  XNOR U12204 ( .A(n11925), .B(n11924), .Z(n11926) );
  NANDN U12205 ( .A(n11842), .B(n11841), .Z(n11846) );
  NANDN U12206 ( .A(n11844), .B(n11843), .Z(n11845) );
  NAND U12207 ( .A(n11846), .B(n11845), .Z(n11927) );
  XNOR U12208 ( .A(n11926), .B(n11927), .Z(n11872) );
  XOR U12209 ( .A(n11873), .B(n11872), .Z(n11931) );
  NANDN U12210 ( .A(n11848), .B(n11847), .Z(n11852) );
  NANDN U12211 ( .A(n11850), .B(n11849), .Z(n11851) );
  AND U12212 ( .A(n11852), .B(n11851), .Z(n11930) );
  XNOR U12213 ( .A(n11931), .B(n11930), .Z(n11932) );
  XOR U12214 ( .A(n11933), .B(n11932), .Z(n11865) );
  NANDN U12215 ( .A(n11854), .B(n11853), .Z(n11858) );
  NAND U12216 ( .A(n11856), .B(n11855), .Z(n11857) );
  AND U12217 ( .A(n11858), .B(n11857), .Z(n11864) );
  XNOR U12218 ( .A(n11865), .B(n11864), .Z(n11866) );
  XNOR U12219 ( .A(n11867), .B(n11866), .Z(n11936) );
  XNOR U12220 ( .A(sreg[401]), .B(n11936), .Z(n11938) );
  NANDN U12221 ( .A(sreg[400]), .B(n11859), .Z(n11863) );
  NAND U12222 ( .A(n11861), .B(n11860), .Z(n11862) );
  NAND U12223 ( .A(n11863), .B(n11862), .Z(n11937) );
  XNOR U12224 ( .A(n11938), .B(n11937), .Z(c[401]) );
  NANDN U12225 ( .A(n11865), .B(n11864), .Z(n11869) );
  NANDN U12226 ( .A(n11867), .B(n11866), .Z(n11868) );
  AND U12227 ( .A(n11869), .B(n11868), .Z(n11944) );
  NANDN U12228 ( .A(n11871), .B(n11870), .Z(n11875) );
  NAND U12229 ( .A(n11873), .B(n11872), .Z(n11874) );
  AND U12230 ( .A(n11875), .B(n11874), .Z(n12010) );
  NANDN U12231 ( .A(n11877), .B(n11876), .Z(n11881) );
  NANDN U12232 ( .A(n11879), .B(n11878), .Z(n11880) );
  AND U12233 ( .A(n11881), .B(n11880), .Z(n11997) );
  NAND U12234 ( .A(b[0]), .B(a[162]), .Z(n11882) );
  XNOR U12235 ( .A(b[1]), .B(n11882), .Z(n11884) );
  NANDN U12236 ( .A(b[0]), .B(a[161]), .Z(n11883) );
  NAND U12237 ( .A(n11884), .B(n11883), .Z(n11977) );
  NAND U12238 ( .A(n19808), .B(n11885), .Z(n11887) );
  XOR U12239 ( .A(b[13]), .B(a[150]), .Z(n11983) );
  NAND U12240 ( .A(n19768), .B(n11983), .Z(n11886) );
  AND U12241 ( .A(n11887), .B(n11886), .Z(n11975) );
  AND U12242 ( .A(b[15]), .B(a[146]), .Z(n11974) );
  XNOR U12243 ( .A(n11975), .B(n11974), .Z(n11976) );
  XNOR U12244 ( .A(n11977), .B(n11976), .Z(n11995) );
  NAND U12245 ( .A(n33), .B(n11888), .Z(n11890) );
  XOR U12246 ( .A(b[5]), .B(a[158]), .Z(n11986) );
  NAND U12247 ( .A(n19342), .B(n11986), .Z(n11889) );
  AND U12248 ( .A(n11890), .B(n11889), .Z(n11971) );
  NAND U12249 ( .A(n34), .B(n11891), .Z(n11893) );
  XOR U12250 ( .A(b[7]), .B(a[156]), .Z(n11989) );
  NAND U12251 ( .A(n19486), .B(n11989), .Z(n11892) );
  AND U12252 ( .A(n11893), .B(n11892), .Z(n11969) );
  NAND U12253 ( .A(n31), .B(n11894), .Z(n11896) );
  XOR U12254 ( .A(b[3]), .B(a[160]), .Z(n11992) );
  NAND U12255 ( .A(n32), .B(n11992), .Z(n11895) );
  NAND U12256 ( .A(n11896), .B(n11895), .Z(n11968) );
  XNOR U12257 ( .A(n11969), .B(n11968), .Z(n11970) );
  XOR U12258 ( .A(n11971), .B(n11970), .Z(n11996) );
  XOR U12259 ( .A(n11995), .B(n11996), .Z(n11998) );
  XOR U12260 ( .A(n11997), .B(n11998), .Z(n11948) );
  NANDN U12261 ( .A(n11898), .B(n11897), .Z(n11902) );
  OR U12262 ( .A(n11900), .B(n11899), .Z(n11901) );
  AND U12263 ( .A(n11902), .B(n11901), .Z(n11947) );
  XNOR U12264 ( .A(n11948), .B(n11947), .Z(n11950) );
  NAND U12265 ( .A(n11903), .B(n19724), .Z(n11905) );
  XOR U12266 ( .A(b[11]), .B(a[152]), .Z(n11953) );
  NAND U12267 ( .A(n19692), .B(n11953), .Z(n11904) );
  AND U12268 ( .A(n11905), .B(n11904), .Z(n11964) );
  NAND U12269 ( .A(n19838), .B(n11906), .Z(n11908) );
  XOR U12270 ( .A(b[15]), .B(a[148]), .Z(n11956) );
  NAND U12271 ( .A(n19805), .B(n11956), .Z(n11907) );
  AND U12272 ( .A(n11908), .B(n11907), .Z(n11963) );
  NAND U12273 ( .A(n35), .B(n11909), .Z(n11911) );
  XOR U12274 ( .A(b[9]), .B(a[154]), .Z(n11959) );
  NAND U12275 ( .A(n19598), .B(n11959), .Z(n11910) );
  NAND U12276 ( .A(n11911), .B(n11910), .Z(n11962) );
  XOR U12277 ( .A(n11963), .B(n11962), .Z(n11965) );
  XOR U12278 ( .A(n11964), .B(n11965), .Z(n12002) );
  NANDN U12279 ( .A(n11913), .B(n11912), .Z(n11917) );
  OR U12280 ( .A(n11915), .B(n11914), .Z(n11916) );
  AND U12281 ( .A(n11917), .B(n11916), .Z(n12001) );
  XNOR U12282 ( .A(n12002), .B(n12001), .Z(n12003) );
  NANDN U12283 ( .A(n11919), .B(n11918), .Z(n11923) );
  NANDN U12284 ( .A(n11921), .B(n11920), .Z(n11922) );
  NAND U12285 ( .A(n11923), .B(n11922), .Z(n12004) );
  XNOR U12286 ( .A(n12003), .B(n12004), .Z(n11949) );
  XOR U12287 ( .A(n11950), .B(n11949), .Z(n12008) );
  NANDN U12288 ( .A(n11925), .B(n11924), .Z(n11929) );
  NANDN U12289 ( .A(n11927), .B(n11926), .Z(n11928) );
  AND U12290 ( .A(n11929), .B(n11928), .Z(n12007) );
  XNOR U12291 ( .A(n12008), .B(n12007), .Z(n12009) );
  XOR U12292 ( .A(n12010), .B(n12009), .Z(n11942) );
  NANDN U12293 ( .A(n11931), .B(n11930), .Z(n11935) );
  NAND U12294 ( .A(n11933), .B(n11932), .Z(n11934) );
  AND U12295 ( .A(n11935), .B(n11934), .Z(n11941) );
  XNOR U12296 ( .A(n11942), .B(n11941), .Z(n11943) );
  XNOR U12297 ( .A(n11944), .B(n11943), .Z(n12013) );
  XNOR U12298 ( .A(sreg[402]), .B(n12013), .Z(n12015) );
  NANDN U12299 ( .A(sreg[401]), .B(n11936), .Z(n11940) );
  NAND U12300 ( .A(n11938), .B(n11937), .Z(n11939) );
  NAND U12301 ( .A(n11940), .B(n11939), .Z(n12014) );
  XNOR U12302 ( .A(n12015), .B(n12014), .Z(c[402]) );
  NANDN U12303 ( .A(n11942), .B(n11941), .Z(n11946) );
  NANDN U12304 ( .A(n11944), .B(n11943), .Z(n11945) );
  AND U12305 ( .A(n11946), .B(n11945), .Z(n12021) );
  NANDN U12306 ( .A(n11948), .B(n11947), .Z(n11952) );
  NAND U12307 ( .A(n11950), .B(n11949), .Z(n11951) );
  AND U12308 ( .A(n11952), .B(n11951), .Z(n12087) );
  NAND U12309 ( .A(n11953), .B(n19724), .Z(n11955) );
  XOR U12310 ( .A(b[11]), .B(a[153]), .Z(n12057) );
  NAND U12311 ( .A(n19692), .B(n12057), .Z(n11954) );
  AND U12312 ( .A(n11955), .B(n11954), .Z(n12068) );
  NAND U12313 ( .A(n19838), .B(n11956), .Z(n11958) );
  XOR U12314 ( .A(b[15]), .B(a[149]), .Z(n12060) );
  NAND U12315 ( .A(n19805), .B(n12060), .Z(n11957) );
  AND U12316 ( .A(n11958), .B(n11957), .Z(n12067) );
  NAND U12317 ( .A(n35), .B(n11959), .Z(n11961) );
  XOR U12318 ( .A(b[9]), .B(a[155]), .Z(n12063) );
  NAND U12319 ( .A(n19598), .B(n12063), .Z(n11960) );
  NAND U12320 ( .A(n11961), .B(n11960), .Z(n12066) );
  XOR U12321 ( .A(n12067), .B(n12066), .Z(n12069) );
  XOR U12322 ( .A(n12068), .B(n12069), .Z(n12079) );
  NANDN U12323 ( .A(n11963), .B(n11962), .Z(n11967) );
  OR U12324 ( .A(n11965), .B(n11964), .Z(n11966) );
  AND U12325 ( .A(n11967), .B(n11966), .Z(n12078) );
  XNOR U12326 ( .A(n12079), .B(n12078), .Z(n12080) );
  NANDN U12327 ( .A(n11969), .B(n11968), .Z(n11973) );
  NANDN U12328 ( .A(n11971), .B(n11970), .Z(n11972) );
  NAND U12329 ( .A(n11973), .B(n11972), .Z(n12081) );
  XNOR U12330 ( .A(n12080), .B(n12081), .Z(n12027) );
  NANDN U12331 ( .A(n11975), .B(n11974), .Z(n11979) );
  NANDN U12332 ( .A(n11977), .B(n11976), .Z(n11978) );
  AND U12333 ( .A(n11979), .B(n11978), .Z(n12053) );
  NAND U12334 ( .A(b[0]), .B(a[163]), .Z(n11980) );
  XNOR U12335 ( .A(b[1]), .B(n11980), .Z(n11982) );
  NANDN U12336 ( .A(b[0]), .B(a[162]), .Z(n11981) );
  NAND U12337 ( .A(n11982), .B(n11981), .Z(n12033) );
  NAND U12338 ( .A(n19808), .B(n11983), .Z(n11985) );
  XOR U12339 ( .A(b[13]), .B(a[151]), .Z(n12039) );
  NAND U12340 ( .A(n19768), .B(n12039), .Z(n11984) );
  AND U12341 ( .A(n11985), .B(n11984), .Z(n12031) );
  AND U12342 ( .A(b[15]), .B(a[147]), .Z(n12030) );
  XNOR U12343 ( .A(n12031), .B(n12030), .Z(n12032) );
  XNOR U12344 ( .A(n12033), .B(n12032), .Z(n12051) );
  NAND U12345 ( .A(n33), .B(n11986), .Z(n11988) );
  XOR U12346 ( .A(b[5]), .B(a[159]), .Z(n12042) );
  NAND U12347 ( .A(n19342), .B(n12042), .Z(n11987) );
  AND U12348 ( .A(n11988), .B(n11987), .Z(n12075) );
  NAND U12349 ( .A(n34), .B(n11989), .Z(n11991) );
  XOR U12350 ( .A(b[7]), .B(a[157]), .Z(n12045) );
  NAND U12351 ( .A(n19486), .B(n12045), .Z(n11990) );
  AND U12352 ( .A(n11991), .B(n11990), .Z(n12073) );
  NAND U12353 ( .A(n31), .B(n11992), .Z(n11994) );
  XOR U12354 ( .A(b[3]), .B(a[161]), .Z(n12048) );
  NAND U12355 ( .A(n32), .B(n12048), .Z(n11993) );
  NAND U12356 ( .A(n11994), .B(n11993), .Z(n12072) );
  XNOR U12357 ( .A(n12073), .B(n12072), .Z(n12074) );
  XOR U12358 ( .A(n12075), .B(n12074), .Z(n12052) );
  XOR U12359 ( .A(n12051), .B(n12052), .Z(n12054) );
  XOR U12360 ( .A(n12053), .B(n12054), .Z(n12025) );
  NANDN U12361 ( .A(n11996), .B(n11995), .Z(n12000) );
  OR U12362 ( .A(n11998), .B(n11997), .Z(n11999) );
  AND U12363 ( .A(n12000), .B(n11999), .Z(n12024) );
  XNOR U12364 ( .A(n12025), .B(n12024), .Z(n12026) );
  XOR U12365 ( .A(n12027), .B(n12026), .Z(n12085) );
  NANDN U12366 ( .A(n12002), .B(n12001), .Z(n12006) );
  NANDN U12367 ( .A(n12004), .B(n12003), .Z(n12005) );
  AND U12368 ( .A(n12006), .B(n12005), .Z(n12084) );
  XNOR U12369 ( .A(n12085), .B(n12084), .Z(n12086) );
  XOR U12370 ( .A(n12087), .B(n12086), .Z(n12019) );
  NANDN U12371 ( .A(n12008), .B(n12007), .Z(n12012) );
  NAND U12372 ( .A(n12010), .B(n12009), .Z(n12011) );
  AND U12373 ( .A(n12012), .B(n12011), .Z(n12018) );
  XNOR U12374 ( .A(n12019), .B(n12018), .Z(n12020) );
  XNOR U12375 ( .A(n12021), .B(n12020), .Z(n12090) );
  XNOR U12376 ( .A(sreg[403]), .B(n12090), .Z(n12092) );
  NANDN U12377 ( .A(sreg[402]), .B(n12013), .Z(n12017) );
  NAND U12378 ( .A(n12015), .B(n12014), .Z(n12016) );
  NAND U12379 ( .A(n12017), .B(n12016), .Z(n12091) );
  XNOR U12380 ( .A(n12092), .B(n12091), .Z(c[403]) );
  NANDN U12381 ( .A(n12019), .B(n12018), .Z(n12023) );
  NANDN U12382 ( .A(n12021), .B(n12020), .Z(n12022) );
  AND U12383 ( .A(n12023), .B(n12022), .Z(n12098) );
  NANDN U12384 ( .A(n12025), .B(n12024), .Z(n12029) );
  NAND U12385 ( .A(n12027), .B(n12026), .Z(n12028) );
  AND U12386 ( .A(n12029), .B(n12028), .Z(n12164) );
  NANDN U12387 ( .A(n12031), .B(n12030), .Z(n12035) );
  NANDN U12388 ( .A(n12033), .B(n12032), .Z(n12034) );
  AND U12389 ( .A(n12035), .B(n12034), .Z(n12130) );
  NAND U12390 ( .A(b[0]), .B(a[164]), .Z(n12036) );
  XNOR U12391 ( .A(b[1]), .B(n12036), .Z(n12038) );
  NANDN U12392 ( .A(b[0]), .B(a[163]), .Z(n12037) );
  NAND U12393 ( .A(n12038), .B(n12037), .Z(n12110) );
  NAND U12394 ( .A(n19808), .B(n12039), .Z(n12041) );
  XOR U12395 ( .A(b[13]), .B(a[152]), .Z(n12116) );
  NAND U12396 ( .A(n19768), .B(n12116), .Z(n12040) );
  AND U12397 ( .A(n12041), .B(n12040), .Z(n12108) );
  AND U12398 ( .A(b[15]), .B(a[148]), .Z(n12107) );
  XNOR U12399 ( .A(n12108), .B(n12107), .Z(n12109) );
  XNOR U12400 ( .A(n12110), .B(n12109), .Z(n12128) );
  NAND U12401 ( .A(n33), .B(n12042), .Z(n12044) );
  XOR U12402 ( .A(b[5]), .B(a[160]), .Z(n12119) );
  NAND U12403 ( .A(n19342), .B(n12119), .Z(n12043) );
  AND U12404 ( .A(n12044), .B(n12043), .Z(n12152) );
  NAND U12405 ( .A(n34), .B(n12045), .Z(n12047) );
  XOR U12406 ( .A(b[7]), .B(a[158]), .Z(n12122) );
  NAND U12407 ( .A(n19486), .B(n12122), .Z(n12046) );
  AND U12408 ( .A(n12047), .B(n12046), .Z(n12150) );
  NAND U12409 ( .A(n31), .B(n12048), .Z(n12050) );
  XOR U12410 ( .A(b[3]), .B(a[162]), .Z(n12125) );
  NAND U12411 ( .A(n32), .B(n12125), .Z(n12049) );
  NAND U12412 ( .A(n12050), .B(n12049), .Z(n12149) );
  XNOR U12413 ( .A(n12150), .B(n12149), .Z(n12151) );
  XOR U12414 ( .A(n12152), .B(n12151), .Z(n12129) );
  XOR U12415 ( .A(n12128), .B(n12129), .Z(n12131) );
  XOR U12416 ( .A(n12130), .B(n12131), .Z(n12102) );
  NANDN U12417 ( .A(n12052), .B(n12051), .Z(n12056) );
  OR U12418 ( .A(n12054), .B(n12053), .Z(n12055) );
  AND U12419 ( .A(n12056), .B(n12055), .Z(n12101) );
  XNOR U12420 ( .A(n12102), .B(n12101), .Z(n12104) );
  NAND U12421 ( .A(n12057), .B(n19724), .Z(n12059) );
  XOR U12422 ( .A(b[11]), .B(a[154]), .Z(n12134) );
  NAND U12423 ( .A(n19692), .B(n12134), .Z(n12058) );
  AND U12424 ( .A(n12059), .B(n12058), .Z(n12145) );
  NAND U12425 ( .A(n19838), .B(n12060), .Z(n12062) );
  XOR U12426 ( .A(b[15]), .B(a[150]), .Z(n12137) );
  NAND U12427 ( .A(n19805), .B(n12137), .Z(n12061) );
  AND U12428 ( .A(n12062), .B(n12061), .Z(n12144) );
  NAND U12429 ( .A(n35), .B(n12063), .Z(n12065) );
  XOR U12430 ( .A(b[9]), .B(a[156]), .Z(n12140) );
  NAND U12431 ( .A(n19598), .B(n12140), .Z(n12064) );
  NAND U12432 ( .A(n12065), .B(n12064), .Z(n12143) );
  XOR U12433 ( .A(n12144), .B(n12143), .Z(n12146) );
  XOR U12434 ( .A(n12145), .B(n12146), .Z(n12156) );
  NANDN U12435 ( .A(n12067), .B(n12066), .Z(n12071) );
  OR U12436 ( .A(n12069), .B(n12068), .Z(n12070) );
  AND U12437 ( .A(n12071), .B(n12070), .Z(n12155) );
  XNOR U12438 ( .A(n12156), .B(n12155), .Z(n12157) );
  NANDN U12439 ( .A(n12073), .B(n12072), .Z(n12077) );
  NANDN U12440 ( .A(n12075), .B(n12074), .Z(n12076) );
  NAND U12441 ( .A(n12077), .B(n12076), .Z(n12158) );
  XNOR U12442 ( .A(n12157), .B(n12158), .Z(n12103) );
  XOR U12443 ( .A(n12104), .B(n12103), .Z(n12162) );
  NANDN U12444 ( .A(n12079), .B(n12078), .Z(n12083) );
  NANDN U12445 ( .A(n12081), .B(n12080), .Z(n12082) );
  AND U12446 ( .A(n12083), .B(n12082), .Z(n12161) );
  XNOR U12447 ( .A(n12162), .B(n12161), .Z(n12163) );
  XOR U12448 ( .A(n12164), .B(n12163), .Z(n12096) );
  NANDN U12449 ( .A(n12085), .B(n12084), .Z(n12089) );
  NAND U12450 ( .A(n12087), .B(n12086), .Z(n12088) );
  AND U12451 ( .A(n12089), .B(n12088), .Z(n12095) );
  XNOR U12452 ( .A(n12096), .B(n12095), .Z(n12097) );
  XNOR U12453 ( .A(n12098), .B(n12097), .Z(n12167) );
  XNOR U12454 ( .A(sreg[404]), .B(n12167), .Z(n12169) );
  NANDN U12455 ( .A(sreg[403]), .B(n12090), .Z(n12094) );
  NAND U12456 ( .A(n12092), .B(n12091), .Z(n12093) );
  NAND U12457 ( .A(n12094), .B(n12093), .Z(n12168) );
  XNOR U12458 ( .A(n12169), .B(n12168), .Z(c[404]) );
  NANDN U12459 ( .A(n12096), .B(n12095), .Z(n12100) );
  NANDN U12460 ( .A(n12098), .B(n12097), .Z(n12099) );
  AND U12461 ( .A(n12100), .B(n12099), .Z(n12175) );
  NANDN U12462 ( .A(n12102), .B(n12101), .Z(n12106) );
  NAND U12463 ( .A(n12104), .B(n12103), .Z(n12105) );
  AND U12464 ( .A(n12106), .B(n12105), .Z(n12241) );
  NANDN U12465 ( .A(n12108), .B(n12107), .Z(n12112) );
  NANDN U12466 ( .A(n12110), .B(n12109), .Z(n12111) );
  AND U12467 ( .A(n12112), .B(n12111), .Z(n12207) );
  NAND U12468 ( .A(b[0]), .B(a[165]), .Z(n12113) );
  XNOR U12469 ( .A(b[1]), .B(n12113), .Z(n12115) );
  NANDN U12470 ( .A(b[0]), .B(a[164]), .Z(n12114) );
  NAND U12471 ( .A(n12115), .B(n12114), .Z(n12187) );
  NAND U12472 ( .A(n19808), .B(n12116), .Z(n12118) );
  XOR U12473 ( .A(b[13]), .B(a[153]), .Z(n12193) );
  NAND U12474 ( .A(n19768), .B(n12193), .Z(n12117) );
  AND U12475 ( .A(n12118), .B(n12117), .Z(n12185) );
  AND U12476 ( .A(b[15]), .B(a[149]), .Z(n12184) );
  XNOR U12477 ( .A(n12185), .B(n12184), .Z(n12186) );
  XNOR U12478 ( .A(n12187), .B(n12186), .Z(n12205) );
  NAND U12479 ( .A(n33), .B(n12119), .Z(n12121) );
  XOR U12480 ( .A(b[5]), .B(a[161]), .Z(n12196) );
  NAND U12481 ( .A(n19342), .B(n12196), .Z(n12120) );
  AND U12482 ( .A(n12121), .B(n12120), .Z(n12229) );
  NAND U12483 ( .A(n34), .B(n12122), .Z(n12124) );
  XOR U12484 ( .A(b[7]), .B(a[159]), .Z(n12199) );
  NAND U12485 ( .A(n19486), .B(n12199), .Z(n12123) );
  AND U12486 ( .A(n12124), .B(n12123), .Z(n12227) );
  NAND U12487 ( .A(n31), .B(n12125), .Z(n12127) );
  XOR U12488 ( .A(b[3]), .B(a[163]), .Z(n12202) );
  NAND U12489 ( .A(n32), .B(n12202), .Z(n12126) );
  NAND U12490 ( .A(n12127), .B(n12126), .Z(n12226) );
  XNOR U12491 ( .A(n12227), .B(n12226), .Z(n12228) );
  XOR U12492 ( .A(n12229), .B(n12228), .Z(n12206) );
  XOR U12493 ( .A(n12205), .B(n12206), .Z(n12208) );
  XOR U12494 ( .A(n12207), .B(n12208), .Z(n12179) );
  NANDN U12495 ( .A(n12129), .B(n12128), .Z(n12133) );
  OR U12496 ( .A(n12131), .B(n12130), .Z(n12132) );
  AND U12497 ( .A(n12133), .B(n12132), .Z(n12178) );
  XNOR U12498 ( .A(n12179), .B(n12178), .Z(n12181) );
  NAND U12499 ( .A(n12134), .B(n19724), .Z(n12136) );
  XOR U12500 ( .A(b[11]), .B(a[155]), .Z(n12211) );
  NAND U12501 ( .A(n19692), .B(n12211), .Z(n12135) );
  AND U12502 ( .A(n12136), .B(n12135), .Z(n12222) );
  NAND U12503 ( .A(n19838), .B(n12137), .Z(n12139) );
  XOR U12504 ( .A(b[15]), .B(a[151]), .Z(n12214) );
  NAND U12505 ( .A(n19805), .B(n12214), .Z(n12138) );
  AND U12506 ( .A(n12139), .B(n12138), .Z(n12221) );
  NAND U12507 ( .A(n35), .B(n12140), .Z(n12142) );
  XOR U12508 ( .A(b[9]), .B(a[157]), .Z(n12217) );
  NAND U12509 ( .A(n19598), .B(n12217), .Z(n12141) );
  NAND U12510 ( .A(n12142), .B(n12141), .Z(n12220) );
  XOR U12511 ( .A(n12221), .B(n12220), .Z(n12223) );
  XOR U12512 ( .A(n12222), .B(n12223), .Z(n12233) );
  NANDN U12513 ( .A(n12144), .B(n12143), .Z(n12148) );
  OR U12514 ( .A(n12146), .B(n12145), .Z(n12147) );
  AND U12515 ( .A(n12148), .B(n12147), .Z(n12232) );
  XNOR U12516 ( .A(n12233), .B(n12232), .Z(n12234) );
  NANDN U12517 ( .A(n12150), .B(n12149), .Z(n12154) );
  NANDN U12518 ( .A(n12152), .B(n12151), .Z(n12153) );
  NAND U12519 ( .A(n12154), .B(n12153), .Z(n12235) );
  XNOR U12520 ( .A(n12234), .B(n12235), .Z(n12180) );
  XOR U12521 ( .A(n12181), .B(n12180), .Z(n12239) );
  NANDN U12522 ( .A(n12156), .B(n12155), .Z(n12160) );
  NANDN U12523 ( .A(n12158), .B(n12157), .Z(n12159) );
  AND U12524 ( .A(n12160), .B(n12159), .Z(n12238) );
  XNOR U12525 ( .A(n12239), .B(n12238), .Z(n12240) );
  XOR U12526 ( .A(n12241), .B(n12240), .Z(n12173) );
  NANDN U12527 ( .A(n12162), .B(n12161), .Z(n12166) );
  NAND U12528 ( .A(n12164), .B(n12163), .Z(n12165) );
  AND U12529 ( .A(n12166), .B(n12165), .Z(n12172) );
  XNOR U12530 ( .A(n12173), .B(n12172), .Z(n12174) );
  XNOR U12531 ( .A(n12175), .B(n12174), .Z(n12244) );
  XNOR U12532 ( .A(sreg[405]), .B(n12244), .Z(n12246) );
  NANDN U12533 ( .A(sreg[404]), .B(n12167), .Z(n12171) );
  NAND U12534 ( .A(n12169), .B(n12168), .Z(n12170) );
  NAND U12535 ( .A(n12171), .B(n12170), .Z(n12245) );
  XNOR U12536 ( .A(n12246), .B(n12245), .Z(c[405]) );
  NANDN U12537 ( .A(n12173), .B(n12172), .Z(n12177) );
  NANDN U12538 ( .A(n12175), .B(n12174), .Z(n12176) );
  AND U12539 ( .A(n12177), .B(n12176), .Z(n12252) );
  NANDN U12540 ( .A(n12179), .B(n12178), .Z(n12183) );
  NAND U12541 ( .A(n12181), .B(n12180), .Z(n12182) );
  AND U12542 ( .A(n12183), .B(n12182), .Z(n12318) );
  NANDN U12543 ( .A(n12185), .B(n12184), .Z(n12189) );
  NANDN U12544 ( .A(n12187), .B(n12186), .Z(n12188) );
  AND U12545 ( .A(n12189), .B(n12188), .Z(n12284) );
  NAND U12546 ( .A(b[0]), .B(a[166]), .Z(n12190) );
  XNOR U12547 ( .A(b[1]), .B(n12190), .Z(n12192) );
  NANDN U12548 ( .A(b[0]), .B(a[165]), .Z(n12191) );
  NAND U12549 ( .A(n12192), .B(n12191), .Z(n12264) );
  NAND U12550 ( .A(n19808), .B(n12193), .Z(n12195) );
  XOR U12551 ( .A(b[13]), .B(a[154]), .Z(n12270) );
  NAND U12552 ( .A(n19768), .B(n12270), .Z(n12194) );
  AND U12553 ( .A(n12195), .B(n12194), .Z(n12262) );
  AND U12554 ( .A(b[15]), .B(a[150]), .Z(n12261) );
  XNOR U12555 ( .A(n12262), .B(n12261), .Z(n12263) );
  XNOR U12556 ( .A(n12264), .B(n12263), .Z(n12282) );
  NAND U12557 ( .A(n33), .B(n12196), .Z(n12198) );
  XOR U12558 ( .A(b[5]), .B(a[162]), .Z(n12273) );
  NAND U12559 ( .A(n19342), .B(n12273), .Z(n12197) );
  AND U12560 ( .A(n12198), .B(n12197), .Z(n12306) );
  NAND U12561 ( .A(n34), .B(n12199), .Z(n12201) );
  XOR U12562 ( .A(b[7]), .B(a[160]), .Z(n12276) );
  NAND U12563 ( .A(n19486), .B(n12276), .Z(n12200) );
  AND U12564 ( .A(n12201), .B(n12200), .Z(n12304) );
  NAND U12565 ( .A(n31), .B(n12202), .Z(n12204) );
  XOR U12566 ( .A(b[3]), .B(a[164]), .Z(n12279) );
  NAND U12567 ( .A(n32), .B(n12279), .Z(n12203) );
  NAND U12568 ( .A(n12204), .B(n12203), .Z(n12303) );
  XNOR U12569 ( .A(n12304), .B(n12303), .Z(n12305) );
  XOR U12570 ( .A(n12306), .B(n12305), .Z(n12283) );
  XOR U12571 ( .A(n12282), .B(n12283), .Z(n12285) );
  XOR U12572 ( .A(n12284), .B(n12285), .Z(n12256) );
  NANDN U12573 ( .A(n12206), .B(n12205), .Z(n12210) );
  OR U12574 ( .A(n12208), .B(n12207), .Z(n12209) );
  AND U12575 ( .A(n12210), .B(n12209), .Z(n12255) );
  XNOR U12576 ( .A(n12256), .B(n12255), .Z(n12258) );
  NAND U12577 ( .A(n12211), .B(n19724), .Z(n12213) );
  XOR U12578 ( .A(b[11]), .B(a[156]), .Z(n12288) );
  NAND U12579 ( .A(n19692), .B(n12288), .Z(n12212) );
  AND U12580 ( .A(n12213), .B(n12212), .Z(n12299) );
  NAND U12581 ( .A(n19838), .B(n12214), .Z(n12216) );
  XOR U12582 ( .A(b[15]), .B(a[152]), .Z(n12291) );
  NAND U12583 ( .A(n19805), .B(n12291), .Z(n12215) );
  AND U12584 ( .A(n12216), .B(n12215), .Z(n12298) );
  NAND U12585 ( .A(n35), .B(n12217), .Z(n12219) );
  XOR U12586 ( .A(b[9]), .B(a[158]), .Z(n12294) );
  NAND U12587 ( .A(n19598), .B(n12294), .Z(n12218) );
  NAND U12588 ( .A(n12219), .B(n12218), .Z(n12297) );
  XOR U12589 ( .A(n12298), .B(n12297), .Z(n12300) );
  XOR U12590 ( .A(n12299), .B(n12300), .Z(n12310) );
  NANDN U12591 ( .A(n12221), .B(n12220), .Z(n12225) );
  OR U12592 ( .A(n12223), .B(n12222), .Z(n12224) );
  AND U12593 ( .A(n12225), .B(n12224), .Z(n12309) );
  XNOR U12594 ( .A(n12310), .B(n12309), .Z(n12311) );
  NANDN U12595 ( .A(n12227), .B(n12226), .Z(n12231) );
  NANDN U12596 ( .A(n12229), .B(n12228), .Z(n12230) );
  NAND U12597 ( .A(n12231), .B(n12230), .Z(n12312) );
  XNOR U12598 ( .A(n12311), .B(n12312), .Z(n12257) );
  XOR U12599 ( .A(n12258), .B(n12257), .Z(n12316) );
  NANDN U12600 ( .A(n12233), .B(n12232), .Z(n12237) );
  NANDN U12601 ( .A(n12235), .B(n12234), .Z(n12236) );
  AND U12602 ( .A(n12237), .B(n12236), .Z(n12315) );
  XNOR U12603 ( .A(n12316), .B(n12315), .Z(n12317) );
  XOR U12604 ( .A(n12318), .B(n12317), .Z(n12250) );
  NANDN U12605 ( .A(n12239), .B(n12238), .Z(n12243) );
  NAND U12606 ( .A(n12241), .B(n12240), .Z(n12242) );
  AND U12607 ( .A(n12243), .B(n12242), .Z(n12249) );
  XNOR U12608 ( .A(n12250), .B(n12249), .Z(n12251) );
  XNOR U12609 ( .A(n12252), .B(n12251), .Z(n12321) );
  XNOR U12610 ( .A(sreg[406]), .B(n12321), .Z(n12323) );
  NANDN U12611 ( .A(sreg[405]), .B(n12244), .Z(n12248) );
  NAND U12612 ( .A(n12246), .B(n12245), .Z(n12247) );
  NAND U12613 ( .A(n12248), .B(n12247), .Z(n12322) );
  XNOR U12614 ( .A(n12323), .B(n12322), .Z(c[406]) );
  NANDN U12615 ( .A(n12250), .B(n12249), .Z(n12254) );
  NANDN U12616 ( .A(n12252), .B(n12251), .Z(n12253) );
  AND U12617 ( .A(n12254), .B(n12253), .Z(n12329) );
  NANDN U12618 ( .A(n12256), .B(n12255), .Z(n12260) );
  NAND U12619 ( .A(n12258), .B(n12257), .Z(n12259) );
  AND U12620 ( .A(n12260), .B(n12259), .Z(n12395) );
  NANDN U12621 ( .A(n12262), .B(n12261), .Z(n12266) );
  NANDN U12622 ( .A(n12264), .B(n12263), .Z(n12265) );
  AND U12623 ( .A(n12266), .B(n12265), .Z(n12361) );
  NAND U12624 ( .A(b[0]), .B(a[167]), .Z(n12267) );
  XNOR U12625 ( .A(b[1]), .B(n12267), .Z(n12269) );
  NANDN U12626 ( .A(b[0]), .B(a[166]), .Z(n12268) );
  NAND U12627 ( .A(n12269), .B(n12268), .Z(n12341) );
  NAND U12628 ( .A(n19808), .B(n12270), .Z(n12272) );
  XOR U12629 ( .A(b[13]), .B(a[155]), .Z(n12347) );
  NAND U12630 ( .A(n19768), .B(n12347), .Z(n12271) );
  AND U12631 ( .A(n12272), .B(n12271), .Z(n12339) );
  AND U12632 ( .A(b[15]), .B(a[151]), .Z(n12338) );
  XNOR U12633 ( .A(n12339), .B(n12338), .Z(n12340) );
  XNOR U12634 ( .A(n12341), .B(n12340), .Z(n12359) );
  NAND U12635 ( .A(n33), .B(n12273), .Z(n12275) );
  XOR U12636 ( .A(b[5]), .B(a[163]), .Z(n12350) );
  NAND U12637 ( .A(n19342), .B(n12350), .Z(n12274) );
  AND U12638 ( .A(n12275), .B(n12274), .Z(n12383) );
  NAND U12639 ( .A(n34), .B(n12276), .Z(n12278) );
  XOR U12640 ( .A(b[7]), .B(a[161]), .Z(n12353) );
  NAND U12641 ( .A(n19486), .B(n12353), .Z(n12277) );
  AND U12642 ( .A(n12278), .B(n12277), .Z(n12381) );
  NAND U12643 ( .A(n31), .B(n12279), .Z(n12281) );
  XOR U12644 ( .A(b[3]), .B(a[165]), .Z(n12356) );
  NAND U12645 ( .A(n32), .B(n12356), .Z(n12280) );
  NAND U12646 ( .A(n12281), .B(n12280), .Z(n12380) );
  XNOR U12647 ( .A(n12381), .B(n12380), .Z(n12382) );
  XOR U12648 ( .A(n12383), .B(n12382), .Z(n12360) );
  XOR U12649 ( .A(n12359), .B(n12360), .Z(n12362) );
  XOR U12650 ( .A(n12361), .B(n12362), .Z(n12333) );
  NANDN U12651 ( .A(n12283), .B(n12282), .Z(n12287) );
  OR U12652 ( .A(n12285), .B(n12284), .Z(n12286) );
  AND U12653 ( .A(n12287), .B(n12286), .Z(n12332) );
  XNOR U12654 ( .A(n12333), .B(n12332), .Z(n12335) );
  NAND U12655 ( .A(n12288), .B(n19724), .Z(n12290) );
  XOR U12656 ( .A(b[11]), .B(a[157]), .Z(n12365) );
  NAND U12657 ( .A(n19692), .B(n12365), .Z(n12289) );
  AND U12658 ( .A(n12290), .B(n12289), .Z(n12376) );
  NAND U12659 ( .A(n19838), .B(n12291), .Z(n12293) );
  XOR U12660 ( .A(b[15]), .B(a[153]), .Z(n12368) );
  NAND U12661 ( .A(n19805), .B(n12368), .Z(n12292) );
  AND U12662 ( .A(n12293), .B(n12292), .Z(n12375) );
  NAND U12663 ( .A(n35), .B(n12294), .Z(n12296) );
  XOR U12664 ( .A(b[9]), .B(a[159]), .Z(n12371) );
  NAND U12665 ( .A(n19598), .B(n12371), .Z(n12295) );
  NAND U12666 ( .A(n12296), .B(n12295), .Z(n12374) );
  XOR U12667 ( .A(n12375), .B(n12374), .Z(n12377) );
  XOR U12668 ( .A(n12376), .B(n12377), .Z(n12387) );
  NANDN U12669 ( .A(n12298), .B(n12297), .Z(n12302) );
  OR U12670 ( .A(n12300), .B(n12299), .Z(n12301) );
  AND U12671 ( .A(n12302), .B(n12301), .Z(n12386) );
  XNOR U12672 ( .A(n12387), .B(n12386), .Z(n12388) );
  NANDN U12673 ( .A(n12304), .B(n12303), .Z(n12308) );
  NANDN U12674 ( .A(n12306), .B(n12305), .Z(n12307) );
  NAND U12675 ( .A(n12308), .B(n12307), .Z(n12389) );
  XNOR U12676 ( .A(n12388), .B(n12389), .Z(n12334) );
  XOR U12677 ( .A(n12335), .B(n12334), .Z(n12393) );
  NANDN U12678 ( .A(n12310), .B(n12309), .Z(n12314) );
  NANDN U12679 ( .A(n12312), .B(n12311), .Z(n12313) );
  AND U12680 ( .A(n12314), .B(n12313), .Z(n12392) );
  XNOR U12681 ( .A(n12393), .B(n12392), .Z(n12394) );
  XOR U12682 ( .A(n12395), .B(n12394), .Z(n12327) );
  NANDN U12683 ( .A(n12316), .B(n12315), .Z(n12320) );
  NAND U12684 ( .A(n12318), .B(n12317), .Z(n12319) );
  AND U12685 ( .A(n12320), .B(n12319), .Z(n12326) );
  XNOR U12686 ( .A(n12327), .B(n12326), .Z(n12328) );
  XNOR U12687 ( .A(n12329), .B(n12328), .Z(n12398) );
  XNOR U12688 ( .A(sreg[407]), .B(n12398), .Z(n12400) );
  NANDN U12689 ( .A(sreg[406]), .B(n12321), .Z(n12325) );
  NAND U12690 ( .A(n12323), .B(n12322), .Z(n12324) );
  NAND U12691 ( .A(n12325), .B(n12324), .Z(n12399) );
  XNOR U12692 ( .A(n12400), .B(n12399), .Z(c[407]) );
  NANDN U12693 ( .A(n12327), .B(n12326), .Z(n12331) );
  NANDN U12694 ( .A(n12329), .B(n12328), .Z(n12330) );
  AND U12695 ( .A(n12331), .B(n12330), .Z(n12406) );
  NANDN U12696 ( .A(n12333), .B(n12332), .Z(n12337) );
  NAND U12697 ( .A(n12335), .B(n12334), .Z(n12336) );
  AND U12698 ( .A(n12337), .B(n12336), .Z(n12472) );
  NANDN U12699 ( .A(n12339), .B(n12338), .Z(n12343) );
  NANDN U12700 ( .A(n12341), .B(n12340), .Z(n12342) );
  AND U12701 ( .A(n12343), .B(n12342), .Z(n12438) );
  NAND U12702 ( .A(b[0]), .B(a[168]), .Z(n12344) );
  XNOR U12703 ( .A(b[1]), .B(n12344), .Z(n12346) );
  NANDN U12704 ( .A(b[0]), .B(a[167]), .Z(n12345) );
  NAND U12705 ( .A(n12346), .B(n12345), .Z(n12418) );
  NAND U12706 ( .A(n19808), .B(n12347), .Z(n12349) );
  XOR U12707 ( .A(b[13]), .B(a[156]), .Z(n12421) );
  NAND U12708 ( .A(n19768), .B(n12421), .Z(n12348) );
  AND U12709 ( .A(n12349), .B(n12348), .Z(n12416) );
  AND U12710 ( .A(b[15]), .B(a[152]), .Z(n12415) );
  XNOR U12711 ( .A(n12416), .B(n12415), .Z(n12417) );
  XNOR U12712 ( .A(n12418), .B(n12417), .Z(n12436) );
  NAND U12713 ( .A(n33), .B(n12350), .Z(n12352) );
  XOR U12714 ( .A(b[5]), .B(a[164]), .Z(n12427) );
  NAND U12715 ( .A(n19342), .B(n12427), .Z(n12351) );
  AND U12716 ( .A(n12352), .B(n12351), .Z(n12460) );
  NAND U12717 ( .A(n34), .B(n12353), .Z(n12355) );
  XOR U12718 ( .A(b[7]), .B(a[162]), .Z(n12430) );
  NAND U12719 ( .A(n19486), .B(n12430), .Z(n12354) );
  AND U12720 ( .A(n12355), .B(n12354), .Z(n12458) );
  NAND U12721 ( .A(n31), .B(n12356), .Z(n12358) );
  XOR U12722 ( .A(b[3]), .B(a[166]), .Z(n12433) );
  NAND U12723 ( .A(n32), .B(n12433), .Z(n12357) );
  NAND U12724 ( .A(n12358), .B(n12357), .Z(n12457) );
  XNOR U12725 ( .A(n12458), .B(n12457), .Z(n12459) );
  XOR U12726 ( .A(n12460), .B(n12459), .Z(n12437) );
  XOR U12727 ( .A(n12436), .B(n12437), .Z(n12439) );
  XOR U12728 ( .A(n12438), .B(n12439), .Z(n12410) );
  NANDN U12729 ( .A(n12360), .B(n12359), .Z(n12364) );
  OR U12730 ( .A(n12362), .B(n12361), .Z(n12363) );
  AND U12731 ( .A(n12364), .B(n12363), .Z(n12409) );
  XNOR U12732 ( .A(n12410), .B(n12409), .Z(n12412) );
  NAND U12733 ( .A(n12365), .B(n19724), .Z(n12367) );
  XOR U12734 ( .A(b[11]), .B(a[158]), .Z(n12442) );
  NAND U12735 ( .A(n19692), .B(n12442), .Z(n12366) );
  AND U12736 ( .A(n12367), .B(n12366), .Z(n12453) );
  NAND U12737 ( .A(n19838), .B(n12368), .Z(n12370) );
  XOR U12738 ( .A(b[15]), .B(a[154]), .Z(n12445) );
  NAND U12739 ( .A(n19805), .B(n12445), .Z(n12369) );
  AND U12740 ( .A(n12370), .B(n12369), .Z(n12452) );
  NAND U12741 ( .A(n35), .B(n12371), .Z(n12373) );
  XOR U12742 ( .A(b[9]), .B(a[160]), .Z(n12448) );
  NAND U12743 ( .A(n19598), .B(n12448), .Z(n12372) );
  NAND U12744 ( .A(n12373), .B(n12372), .Z(n12451) );
  XOR U12745 ( .A(n12452), .B(n12451), .Z(n12454) );
  XOR U12746 ( .A(n12453), .B(n12454), .Z(n12464) );
  NANDN U12747 ( .A(n12375), .B(n12374), .Z(n12379) );
  OR U12748 ( .A(n12377), .B(n12376), .Z(n12378) );
  AND U12749 ( .A(n12379), .B(n12378), .Z(n12463) );
  XNOR U12750 ( .A(n12464), .B(n12463), .Z(n12465) );
  NANDN U12751 ( .A(n12381), .B(n12380), .Z(n12385) );
  NANDN U12752 ( .A(n12383), .B(n12382), .Z(n12384) );
  NAND U12753 ( .A(n12385), .B(n12384), .Z(n12466) );
  XNOR U12754 ( .A(n12465), .B(n12466), .Z(n12411) );
  XOR U12755 ( .A(n12412), .B(n12411), .Z(n12470) );
  NANDN U12756 ( .A(n12387), .B(n12386), .Z(n12391) );
  NANDN U12757 ( .A(n12389), .B(n12388), .Z(n12390) );
  AND U12758 ( .A(n12391), .B(n12390), .Z(n12469) );
  XNOR U12759 ( .A(n12470), .B(n12469), .Z(n12471) );
  XOR U12760 ( .A(n12472), .B(n12471), .Z(n12404) );
  NANDN U12761 ( .A(n12393), .B(n12392), .Z(n12397) );
  NAND U12762 ( .A(n12395), .B(n12394), .Z(n12396) );
  AND U12763 ( .A(n12397), .B(n12396), .Z(n12403) );
  XNOR U12764 ( .A(n12404), .B(n12403), .Z(n12405) );
  XNOR U12765 ( .A(n12406), .B(n12405), .Z(n12475) );
  XNOR U12766 ( .A(sreg[408]), .B(n12475), .Z(n12477) );
  NANDN U12767 ( .A(sreg[407]), .B(n12398), .Z(n12402) );
  NAND U12768 ( .A(n12400), .B(n12399), .Z(n12401) );
  NAND U12769 ( .A(n12402), .B(n12401), .Z(n12476) );
  XNOR U12770 ( .A(n12477), .B(n12476), .Z(c[408]) );
  NANDN U12771 ( .A(n12404), .B(n12403), .Z(n12408) );
  NANDN U12772 ( .A(n12406), .B(n12405), .Z(n12407) );
  AND U12773 ( .A(n12408), .B(n12407), .Z(n12483) );
  NANDN U12774 ( .A(n12410), .B(n12409), .Z(n12414) );
  NAND U12775 ( .A(n12412), .B(n12411), .Z(n12413) );
  AND U12776 ( .A(n12414), .B(n12413), .Z(n12549) );
  NANDN U12777 ( .A(n12416), .B(n12415), .Z(n12420) );
  NANDN U12778 ( .A(n12418), .B(n12417), .Z(n12419) );
  AND U12779 ( .A(n12420), .B(n12419), .Z(n12515) );
  NAND U12780 ( .A(n19808), .B(n12421), .Z(n12423) );
  XOR U12781 ( .A(b[13]), .B(a[157]), .Z(n12498) );
  NAND U12782 ( .A(n19768), .B(n12498), .Z(n12422) );
  AND U12783 ( .A(n12423), .B(n12422), .Z(n12493) );
  AND U12784 ( .A(b[15]), .B(a[153]), .Z(n12492) );
  XNOR U12785 ( .A(n12493), .B(n12492), .Z(n12494) );
  NAND U12786 ( .A(b[0]), .B(a[169]), .Z(n12424) );
  XNOR U12787 ( .A(b[1]), .B(n12424), .Z(n12426) );
  NANDN U12788 ( .A(b[0]), .B(a[168]), .Z(n12425) );
  NAND U12789 ( .A(n12426), .B(n12425), .Z(n12495) );
  XNOR U12790 ( .A(n12494), .B(n12495), .Z(n12513) );
  NAND U12791 ( .A(n33), .B(n12427), .Z(n12429) );
  XOR U12792 ( .A(b[5]), .B(a[165]), .Z(n12504) );
  NAND U12793 ( .A(n19342), .B(n12504), .Z(n12428) );
  AND U12794 ( .A(n12429), .B(n12428), .Z(n12537) );
  NAND U12795 ( .A(n34), .B(n12430), .Z(n12432) );
  XOR U12796 ( .A(b[7]), .B(a[163]), .Z(n12507) );
  NAND U12797 ( .A(n19486), .B(n12507), .Z(n12431) );
  AND U12798 ( .A(n12432), .B(n12431), .Z(n12535) );
  NAND U12799 ( .A(n31), .B(n12433), .Z(n12435) );
  XOR U12800 ( .A(b[3]), .B(a[167]), .Z(n12510) );
  NAND U12801 ( .A(n32), .B(n12510), .Z(n12434) );
  NAND U12802 ( .A(n12435), .B(n12434), .Z(n12534) );
  XNOR U12803 ( .A(n12535), .B(n12534), .Z(n12536) );
  XOR U12804 ( .A(n12537), .B(n12536), .Z(n12514) );
  XOR U12805 ( .A(n12513), .B(n12514), .Z(n12516) );
  XOR U12806 ( .A(n12515), .B(n12516), .Z(n12487) );
  NANDN U12807 ( .A(n12437), .B(n12436), .Z(n12441) );
  OR U12808 ( .A(n12439), .B(n12438), .Z(n12440) );
  AND U12809 ( .A(n12441), .B(n12440), .Z(n12486) );
  XNOR U12810 ( .A(n12487), .B(n12486), .Z(n12489) );
  NAND U12811 ( .A(n12442), .B(n19724), .Z(n12444) );
  XOR U12812 ( .A(b[11]), .B(a[159]), .Z(n12519) );
  NAND U12813 ( .A(n19692), .B(n12519), .Z(n12443) );
  AND U12814 ( .A(n12444), .B(n12443), .Z(n12530) );
  NAND U12815 ( .A(n19838), .B(n12445), .Z(n12447) );
  XOR U12816 ( .A(b[15]), .B(a[155]), .Z(n12522) );
  NAND U12817 ( .A(n19805), .B(n12522), .Z(n12446) );
  AND U12818 ( .A(n12447), .B(n12446), .Z(n12529) );
  NAND U12819 ( .A(n35), .B(n12448), .Z(n12450) );
  XOR U12820 ( .A(b[9]), .B(a[161]), .Z(n12525) );
  NAND U12821 ( .A(n19598), .B(n12525), .Z(n12449) );
  NAND U12822 ( .A(n12450), .B(n12449), .Z(n12528) );
  XOR U12823 ( .A(n12529), .B(n12528), .Z(n12531) );
  XOR U12824 ( .A(n12530), .B(n12531), .Z(n12541) );
  NANDN U12825 ( .A(n12452), .B(n12451), .Z(n12456) );
  OR U12826 ( .A(n12454), .B(n12453), .Z(n12455) );
  AND U12827 ( .A(n12456), .B(n12455), .Z(n12540) );
  XNOR U12828 ( .A(n12541), .B(n12540), .Z(n12542) );
  NANDN U12829 ( .A(n12458), .B(n12457), .Z(n12462) );
  NANDN U12830 ( .A(n12460), .B(n12459), .Z(n12461) );
  NAND U12831 ( .A(n12462), .B(n12461), .Z(n12543) );
  XNOR U12832 ( .A(n12542), .B(n12543), .Z(n12488) );
  XOR U12833 ( .A(n12489), .B(n12488), .Z(n12547) );
  NANDN U12834 ( .A(n12464), .B(n12463), .Z(n12468) );
  NANDN U12835 ( .A(n12466), .B(n12465), .Z(n12467) );
  AND U12836 ( .A(n12468), .B(n12467), .Z(n12546) );
  XNOR U12837 ( .A(n12547), .B(n12546), .Z(n12548) );
  XOR U12838 ( .A(n12549), .B(n12548), .Z(n12481) );
  NANDN U12839 ( .A(n12470), .B(n12469), .Z(n12474) );
  NAND U12840 ( .A(n12472), .B(n12471), .Z(n12473) );
  AND U12841 ( .A(n12474), .B(n12473), .Z(n12480) );
  XNOR U12842 ( .A(n12481), .B(n12480), .Z(n12482) );
  XNOR U12843 ( .A(n12483), .B(n12482), .Z(n12552) );
  XNOR U12844 ( .A(sreg[409]), .B(n12552), .Z(n12554) );
  NANDN U12845 ( .A(sreg[408]), .B(n12475), .Z(n12479) );
  NAND U12846 ( .A(n12477), .B(n12476), .Z(n12478) );
  NAND U12847 ( .A(n12479), .B(n12478), .Z(n12553) );
  XNOR U12848 ( .A(n12554), .B(n12553), .Z(c[409]) );
  NANDN U12849 ( .A(n12481), .B(n12480), .Z(n12485) );
  NANDN U12850 ( .A(n12483), .B(n12482), .Z(n12484) );
  AND U12851 ( .A(n12485), .B(n12484), .Z(n12560) );
  NANDN U12852 ( .A(n12487), .B(n12486), .Z(n12491) );
  NAND U12853 ( .A(n12489), .B(n12488), .Z(n12490) );
  AND U12854 ( .A(n12491), .B(n12490), .Z(n12626) );
  NANDN U12855 ( .A(n12493), .B(n12492), .Z(n12497) );
  NANDN U12856 ( .A(n12495), .B(n12494), .Z(n12496) );
  AND U12857 ( .A(n12497), .B(n12496), .Z(n12592) );
  NAND U12858 ( .A(n19808), .B(n12498), .Z(n12500) );
  XOR U12859 ( .A(b[13]), .B(a[158]), .Z(n12578) );
  NAND U12860 ( .A(n19768), .B(n12578), .Z(n12499) );
  AND U12861 ( .A(n12500), .B(n12499), .Z(n12570) );
  AND U12862 ( .A(b[15]), .B(a[154]), .Z(n12569) );
  XNOR U12863 ( .A(n12570), .B(n12569), .Z(n12571) );
  NAND U12864 ( .A(b[0]), .B(a[170]), .Z(n12501) );
  XNOR U12865 ( .A(b[1]), .B(n12501), .Z(n12503) );
  NANDN U12866 ( .A(b[0]), .B(a[169]), .Z(n12502) );
  NAND U12867 ( .A(n12503), .B(n12502), .Z(n12572) );
  XNOR U12868 ( .A(n12571), .B(n12572), .Z(n12590) );
  NAND U12869 ( .A(n33), .B(n12504), .Z(n12506) );
  XOR U12870 ( .A(b[5]), .B(a[166]), .Z(n12581) );
  NAND U12871 ( .A(n19342), .B(n12581), .Z(n12505) );
  AND U12872 ( .A(n12506), .B(n12505), .Z(n12614) );
  NAND U12873 ( .A(n34), .B(n12507), .Z(n12509) );
  XOR U12874 ( .A(b[7]), .B(a[164]), .Z(n12584) );
  NAND U12875 ( .A(n19486), .B(n12584), .Z(n12508) );
  AND U12876 ( .A(n12509), .B(n12508), .Z(n12612) );
  NAND U12877 ( .A(n31), .B(n12510), .Z(n12512) );
  XOR U12878 ( .A(b[3]), .B(a[168]), .Z(n12587) );
  NAND U12879 ( .A(n32), .B(n12587), .Z(n12511) );
  NAND U12880 ( .A(n12512), .B(n12511), .Z(n12611) );
  XNOR U12881 ( .A(n12612), .B(n12611), .Z(n12613) );
  XOR U12882 ( .A(n12614), .B(n12613), .Z(n12591) );
  XOR U12883 ( .A(n12590), .B(n12591), .Z(n12593) );
  XOR U12884 ( .A(n12592), .B(n12593), .Z(n12564) );
  NANDN U12885 ( .A(n12514), .B(n12513), .Z(n12518) );
  OR U12886 ( .A(n12516), .B(n12515), .Z(n12517) );
  AND U12887 ( .A(n12518), .B(n12517), .Z(n12563) );
  XNOR U12888 ( .A(n12564), .B(n12563), .Z(n12566) );
  NAND U12889 ( .A(n12519), .B(n19724), .Z(n12521) );
  XOR U12890 ( .A(b[11]), .B(a[160]), .Z(n12596) );
  NAND U12891 ( .A(n19692), .B(n12596), .Z(n12520) );
  AND U12892 ( .A(n12521), .B(n12520), .Z(n12607) );
  NAND U12893 ( .A(n19838), .B(n12522), .Z(n12524) );
  XOR U12894 ( .A(b[15]), .B(a[156]), .Z(n12599) );
  NAND U12895 ( .A(n19805), .B(n12599), .Z(n12523) );
  AND U12896 ( .A(n12524), .B(n12523), .Z(n12606) );
  NAND U12897 ( .A(n35), .B(n12525), .Z(n12527) );
  XOR U12898 ( .A(b[9]), .B(a[162]), .Z(n12602) );
  NAND U12899 ( .A(n19598), .B(n12602), .Z(n12526) );
  NAND U12900 ( .A(n12527), .B(n12526), .Z(n12605) );
  XOR U12901 ( .A(n12606), .B(n12605), .Z(n12608) );
  XOR U12902 ( .A(n12607), .B(n12608), .Z(n12618) );
  NANDN U12903 ( .A(n12529), .B(n12528), .Z(n12533) );
  OR U12904 ( .A(n12531), .B(n12530), .Z(n12532) );
  AND U12905 ( .A(n12533), .B(n12532), .Z(n12617) );
  XNOR U12906 ( .A(n12618), .B(n12617), .Z(n12619) );
  NANDN U12907 ( .A(n12535), .B(n12534), .Z(n12539) );
  NANDN U12908 ( .A(n12537), .B(n12536), .Z(n12538) );
  NAND U12909 ( .A(n12539), .B(n12538), .Z(n12620) );
  XNOR U12910 ( .A(n12619), .B(n12620), .Z(n12565) );
  XOR U12911 ( .A(n12566), .B(n12565), .Z(n12624) );
  NANDN U12912 ( .A(n12541), .B(n12540), .Z(n12545) );
  NANDN U12913 ( .A(n12543), .B(n12542), .Z(n12544) );
  AND U12914 ( .A(n12545), .B(n12544), .Z(n12623) );
  XNOR U12915 ( .A(n12624), .B(n12623), .Z(n12625) );
  XOR U12916 ( .A(n12626), .B(n12625), .Z(n12558) );
  NANDN U12917 ( .A(n12547), .B(n12546), .Z(n12551) );
  NAND U12918 ( .A(n12549), .B(n12548), .Z(n12550) );
  AND U12919 ( .A(n12551), .B(n12550), .Z(n12557) );
  XNOR U12920 ( .A(n12558), .B(n12557), .Z(n12559) );
  XNOR U12921 ( .A(n12560), .B(n12559), .Z(n12629) );
  XNOR U12922 ( .A(sreg[410]), .B(n12629), .Z(n12631) );
  NANDN U12923 ( .A(sreg[409]), .B(n12552), .Z(n12556) );
  NAND U12924 ( .A(n12554), .B(n12553), .Z(n12555) );
  NAND U12925 ( .A(n12556), .B(n12555), .Z(n12630) );
  XNOR U12926 ( .A(n12631), .B(n12630), .Z(c[410]) );
  NANDN U12927 ( .A(n12558), .B(n12557), .Z(n12562) );
  NANDN U12928 ( .A(n12560), .B(n12559), .Z(n12561) );
  AND U12929 ( .A(n12562), .B(n12561), .Z(n12637) );
  NANDN U12930 ( .A(n12564), .B(n12563), .Z(n12568) );
  NAND U12931 ( .A(n12566), .B(n12565), .Z(n12567) );
  AND U12932 ( .A(n12568), .B(n12567), .Z(n12703) );
  NANDN U12933 ( .A(n12570), .B(n12569), .Z(n12574) );
  NANDN U12934 ( .A(n12572), .B(n12571), .Z(n12573) );
  AND U12935 ( .A(n12574), .B(n12573), .Z(n12690) );
  NAND U12936 ( .A(b[0]), .B(a[171]), .Z(n12575) );
  XNOR U12937 ( .A(b[1]), .B(n12575), .Z(n12577) );
  NANDN U12938 ( .A(b[0]), .B(a[170]), .Z(n12576) );
  NAND U12939 ( .A(n12577), .B(n12576), .Z(n12670) );
  NAND U12940 ( .A(n19808), .B(n12578), .Z(n12580) );
  XOR U12941 ( .A(b[13]), .B(a[159]), .Z(n12673) );
  NAND U12942 ( .A(n19768), .B(n12673), .Z(n12579) );
  AND U12943 ( .A(n12580), .B(n12579), .Z(n12668) );
  AND U12944 ( .A(b[15]), .B(a[155]), .Z(n12667) );
  XNOR U12945 ( .A(n12668), .B(n12667), .Z(n12669) );
  XNOR U12946 ( .A(n12670), .B(n12669), .Z(n12688) );
  NAND U12947 ( .A(n33), .B(n12581), .Z(n12583) );
  XOR U12948 ( .A(b[5]), .B(a[167]), .Z(n12679) );
  NAND U12949 ( .A(n19342), .B(n12679), .Z(n12582) );
  AND U12950 ( .A(n12583), .B(n12582), .Z(n12664) );
  NAND U12951 ( .A(n34), .B(n12584), .Z(n12586) );
  XOR U12952 ( .A(b[7]), .B(a[165]), .Z(n12682) );
  NAND U12953 ( .A(n19486), .B(n12682), .Z(n12585) );
  AND U12954 ( .A(n12586), .B(n12585), .Z(n12662) );
  NAND U12955 ( .A(n31), .B(n12587), .Z(n12589) );
  XOR U12956 ( .A(b[3]), .B(a[169]), .Z(n12685) );
  NAND U12957 ( .A(n32), .B(n12685), .Z(n12588) );
  NAND U12958 ( .A(n12589), .B(n12588), .Z(n12661) );
  XNOR U12959 ( .A(n12662), .B(n12661), .Z(n12663) );
  XOR U12960 ( .A(n12664), .B(n12663), .Z(n12689) );
  XOR U12961 ( .A(n12688), .B(n12689), .Z(n12691) );
  XOR U12962 ( .A(n12690), .B(n12691), .Z(n12641) );
  NANDN U12963 ( .A(n12591), .B(n12590), .Z(n12595) );
  OR U12964 ( .A(n12593), .B(n12592), .Z(n12594) );
  AND U12965 ( .A(n12595), .B(n12594), .Z(n12640) );
  XNOR U12966 ( .A(n12641), .B(n12640), .Z(n12643) );
  NAND U12967 ( .A(n12596), .B(n19724), .Z(n12598) );
  XOR U12968 ( .A(b[11]), .B(a[161]), .Z(n12646) );
  NAND U12969 ( .A(n19692), .B(n12646), .Z(n12597) );
  AND U12970 ( .A(n12598), .B(n12597), .Z(n12657) );
  NAND U12971 ( .A(n19838), .B(n12599), .Z(n12601) );
  XOR U12972 ( .A(b[15]), .B(a[157]), .Z(n12649) );
  NAND U12973 ( .A(n19805), .B(n12649), .Z(n12600) );
  AND U12974 ( .A(n12601), .B(n12600), .Z(n12656) );
  NAND U12975 ( .A(n35), .B(n12602), .Z(n12604) );
  XOR U12976 ( .A(b[9]), .B(a[163]), .Z(n12652) );
  NAND U12977 ( .A(n19598), .B(n12652), .Z(n12603) );
  NAND U12978 ( .A(n12604), .B(n12603), .Z(n12655) );
  XOR U12979 ( .A(n12656), .B(n12655), .Z(n12658) );
  XOR U12980 ( .A(n12657), .B(n12658), .Z(n12695) );
  NANDN U12981 ( .A(n12606), .B(n12605), .Z(n12610) );
  OR U12982 ( .A(n12608), .B(n12607), .Z(n12609) );
  AND U12983 ( .A(n12610), .B(n12609), .Z(n12694) );
  XNOR U12984 ( .A(n12695), .B(n12694), .Z(n12696) );
  NANDN U12985 ( .A(n12612), .B(n12611), .Z(n12616) );
  NANDN U12986 ( .A(n12614), .B(n12613), .Z(n12615) );
  NAND U12987 ( .A(n12616), .B(n12615), .Z(n12697) );
  XNOR U12988 ( .A(n12696), .B(n12697), .Z(n12642) );
  XOR U12989 ( .A(n12643), .B(n12642), .Z(n12701) );
  NANDN U12990 ( .A(n12618), .B(n12617), .Z(n12622) );
  NANDN U12991 ( .A(n12620), .B(n12619), .Z(n12621) );
  AND U12992 ( .A(n12622), .B(n12621), .Z(n12700) );
  XNOR U12993 ( .A(n12701), .B(n12700), .Z(n12702) );
  XOR U12994 ( .A(n12703), .B(n12702), .Z(n12635) );
  NANDN U12995 ( .A(n12624), .B(n12623), .Z(n12628) );
  NAND U12996 ( .A(n12626), .B(n12625), .Z(n12627) );
  AND U12997 ( .A(n12628), .B(n12627), .Z(n12634) );
  XNOR U12998 ( .A(n12635), .B(n12634), .Z(n12636) );
  XNOR U12999 ( .A(n12637), .B(n12636), .Z(n12706) );
  XNOR U13000 ( .A(sreg[411]), .B(n12706), .Z(n12708) );
  NANDN U13001 ( .A(sreg[410]), .B(n12629), .Z(n12633) );
  NAND U13002 ( .A(n12631), .B(n12630), .Z(n12632) );
  NAND U13003 ( .A(n12633), .B(n12632), .Z(n12707) );
  XNOR U13004 ( .A(n12708), .B(n12707), .Z(c[411]) );
  NANDN U13005 ( .A(n12635), .B(n12634), .Z(n12639) );
  NANDN U13006 ( .A(n12637), .B(n12636), .Z(n12638) );
  AND U13007 ( .A(n12639), .B(n12638), .Z(n12714) );
  NANDN U13008 ( .A(n12641), .B(n12640), .Z(n12645) );
  NAND U13009 ( .A(n12643), .B(n12642), .Z(n12644) );
  AND U13010 ( .A(n12645), .B(n12644), .Z(n12780) );
  NAND U13011 ( .A(n12646), .B(n19724), .Z(n12648) );
  XOR U13012 ( .A(b[11]), .B(a[162]), .Z(n12750) );
  NAND U13013 ( .A(n19692), .B(n12750), .Z(n12647) );
  AND U13014 ( .A(n12648), .B(n12647), .Z(n12761) );
  NAND U13015 ( .A(n19838), .B(n12649), .Z(n12651) );
  XOR U13016 ( .A(b[15]), .B(a[158]), .Z(n12753) );
  NAND U13017 ( .A(n19805), .B(n12753), .Z(n12650) );
  AND U13018 ( .A(n12651), .B(n12650), .Z(n12760) );
  NAND U13019 ( .A(n35), .B(n12652), .Z(n12654) );
  XOR U13020 ( .A(b[9]), .B(a[164]), .Z(n12756) );
  NAND U13021 ( .A(n19598), .B(n12756), .Z(n12653) );
  NAND U13022 ( .A(n12654), .B(n12653), .Z(n12759) );
  XOR U13023 ( .A(n12760), .B(n12759), .Z(n12762) );
  XOR U13024 ( .A(n12761), .B(n12762), .Z(n12772) );
  NANDN U13025 ( .A(n12656), .B(n12655), .Z(n12660) );
  OR U13026 ( .A(n12658), .B(n12657), .Z(n12659) );
  AND U13027 ( .A(n12660), .B(n12659), .Z(n12771) );
  XNOR U13028 ( .A(n12772), .B(n12771), .Z(n12773) );
  NANDN U13029 ( .A(n12662), .B(n12661), .Z(n12666) );
  NANDN U13030 ( .A(n12664), .B(n12663), .Z(n12665) );
  NAND U13031 ( .A(n12666), .B(n12665), .Z(n12774) );
  XNOR U13032 ( .A(n12773), .B(n12774), .Z(n12720) );
  NANDN U13033 ( .A(n12668), .B(n12667), .Z(n12672) );
  NANDN U13034 ( .A(n12670), .B(n12669), .Z(n12671) );
  AND U13035 ( .A(n12672), .B(n12671), .Z(n12746) );
  NAND U13036 ( .A(n19808), .B(n12673), .Z(n12675) );
  XOR U13037 ( .A(b[13]), .B(a[160]), .Z(n12732) );
  NAND U13038 ( .A(n19768), .B(n12732), .Z(n12674) );
  AND U13039 ( .A(n12675), .B(n12674), .Z(n12724) );
  AND U13040 ( .A(b[15]), .B(a[156]), .Z(n12723) );
  XNOR U13041 ( .A(n12724), .B(n12723), .Z(n12725) );
  NAND U13042 ( .A(b[0]), .B(a[172]), .Z(n12676) );
  XNOR U13043 ( .A(b[1]), .B(n12676), .Z(n12678) );
  NANDN U13044 ( .A(b[0]), .B(a[171]), .Z(n12677) );
  NAND U13045 ( .A(n12678), .B(n12677), .Z(n12726) );
  XNOR U13046 ( .A(n12725), .B(n12726), .Z(n12744) );
  NAND U13047 ( .A(n33), .B(n12679), .Z(n12681) );
  XOR U13048 ( .A(b[5]), .B(a[168]), .Z(n12735) );
  NAND U13049 ( .A(n19342), .B(n12735), .Z(n12680) );
  AND U13050 ( .A(n12681), .B(n12680), .Z(n12768) );
  NAND U13051 ( .A(n34), .B(n12682), .Z(n12684) );
  XOR U13052 ( .A(b[7]), .B(a[166]), .Z(n12738) );
  NAND U13053 ( .A(n19486), .B(n12738), .Z(n12683) );
  AND U13054 ( .A(n12684), .B(n12683), .Z(n12766) );
  NAND U13055 ( .A(n31), .B(n12685), .Z(n12687) );
  XOR U13056 ( .A(b[3]), .B(a[170]), .Z(n12741) );
  NAND U13057 ( .A(n32), .B(n12741), .Z(n12686) );
  NAND U13058 ( .A(n12687), .B(n12686), .Z(n12765) );
  XNOR U13059 ( .A(n12766), .B(n12765), .Z(n12767) );
  XOR U13060 ( .A(n12768), .B(n12767), .Z(n12745) );
  XOR U13061 ( .A(n12744), .B(n12745), .Z(n12747) );
  XOR U13062 ( .A(n12746), .B(n12747), .Z(n12718) );
  NANDN U13063 ( .A(n12689), .B(n12688), .Z(n12693) );
  OR U13064 ( .A(n12691), .B(n12690), .Z(n12692) );
  AND U13065 ( .A(n12693), .B(n12692), .Z(n12717) );
  XNOR U13066 ( .A(n12718), .B(n12717), .Z(n12719) );
  XOR U13067 ( .A(n12720), .B(n12719), .Z(n12778) );
  NANDN U13068 ( .A(n12695), .B(n12694), .Z(n12699) );
  NANDN U13069 ( .A(n12697), .B(n12696), .Z(n12698) );
  AND U13070 ( .A(n12699), .B(n12698), .Z(n12777) );
  XNOR U13071 ( .A(n12778), .B(n12777), .Z(n12779) );
  XOR U13072 ( .A(n12780), .B(n12779), .Z(n12712) );
  NANDN U13073 ( .A(n12701), .B(n12700), .Z(n12705) );
  NAND U13074 ( .A(n12703), .B(n12702), .Z(n12704) );
  AND U13075 ( .A(n12705), .B(n12704), .Z(n12711) );
  XNOR U13076 ( .A(n12712), .B(n12711), .Z(n12713) );
  XNOR U13077 ( .A(n12714), .B(n12713), .Z(n12783) );
  XNOR U13078 ( .A(sreg[412]), .B(n12783), .Z(n12785) );
  NANDN U13079 ( .A(sreg[411]), .B(n12706), .Z(n12710) );
  NAND U13080 ( .A(n12708), .B(n12707), .Z(n12709) );
  NAND U13081 ( .A(n12710), .B(n12709), .Z(n12784) );
  XNOR U13082 ( .A(n12785), .B(n12784), .Z(c[412]) );
  NANDN U13083 ( .A(n12712), .B(n12711), .Z(n12716) );
  NANDN U13084 ( .A(n12714), .B(n12713), .Z(n12715) );
  AND U13085 ( .A(n12716), .B(n12715), .Z(n12791) );
  NANDN U13086 ( .A(n12718), .B(n12717), .Z(n12722) );
  NAND U13087 ( .A(n12720), .B(n12719), .Z(n12721) );
  AND U13088 ( .A(n12722), .B(n12721), .Z(n12857) );
  NANDN U13089 ( .A(n12724), .B(n12723), .Z(n12728) );
  NANDN U13090 ( .A(n12726), .B(n12725), .Z(n12727) );
  AND U13091 ( .A(n12728), .B(n12727), .Z(n12823) );
  NAND U13092 ( .A(b[0]), .B(a[173]), .Z(n12729) );
  XNOR U13093 ( .A(b[1]), .B(n12729), .Z(n12731) );
  NANDN U13094 ( .A(b[0]), .B(a[172]), .Z(n12730) );
  NAND U13095 ( .A(n12731), .B(n12730), .Z(n12803) );
  NAND U13096 ( .A(n19808), .B(n12732), .Z(n12734) );
  XOR U13097 ( .A(b[13]), .B(a[161]), .Z(n12809) );
  NAND U13098 ( .A(n19768), .B(n12809), .Z(n12733) );
  AND U13099 ( .A(n12734), .B(n12733), .Z(n12801) );
  AND U13100 ( .A(b[15]), .B(a[157]), .Z(n12800) );
  XNOR U13101 ( .A(n12801), .B(n12800), .Z(n12802) );
  XNOR U13102 ( .A(n12803), .B(n12802), .Z(n12821) );
  NAND U13103 ( .A(n33), .B(n12735), .Z(n12737) );
  XOR U13104 ( .A(b[5]), .B(a[169]), .Z(n12812) );
  NAND U13105 ( .A(n19342), .B(n12812), .Z(n12736) );
  AND U13106 ( .A(n12737), .B(n12736), .Z(n12845) );
  NAND U13107 ( .A(n34), .B(n12738), .Z(n12740) );
  XOR U13108 ( .A(b[7]), .B(a[167]), .Z(n12815) );
  NAND U13109 ( .A(n19486), .B(n12815), .Z(n12739) );
  AND U13110 ( .A(n12740), .B(n12739), .Z(n12843) );
  NAND U13111 ( .A(n31), .B(n12741), .Z(n12743) );
  XOR U13112 ( .A(b[3]), .B(a[171]), .Z(n12818) );
  NAND U13113 ( .A(n32), .B(n12818), .Z(n12742) );
  NAND U13114 ( .A(n12743), .B(n12742), .Z(n12842) );
  XNOR U13115 ( .A(n12843), .B(n12842), .Z(n12844) );
  XOR U13116 ( .A(n12845), .B(n12844), .Z(n12822) );
  XOR U13117 ( .A(n12821), .B(n12822), .Z(n12824) );
  XOR U13118 ( .A(n12823), .B(n12824), .Z(n12795) );
  NANDN U13119 ( .A(n12745), .B(n12744), .Z(n12749) );
  OR U13120 ( .A(n12747), .B(n12746), .Z(n12748) );
  AND U13121 ( .A(n12749), .B(n12748), .Z(n12794) );
  XNOR U13122 ( .A(n12795), .B(n12794), .Z(n12797) );
  NAND U13123 ( .A(n12750), .B(n19724), .Z(n12752) );
  XOR U13124 ( .A(b[11]), .B(a[163]), .Z(n12827) );
  NAND U13125 ( .A(n19692), .B(n12827), .Z(n12751) );
  AND U13126 ( .A(n12752), .B(n12751), .Z(n12838) );
  NAND U13127 ( .A(n19838), .B(n12753), .Z(n12755) );
  XOR U13128 ( .A(b[15]), .B(a[159]), .Z(n12830) );
  NAND U13129 ( .A(n19805), .B(n12830), .Z(n12754) );
  AND U13130 ( .A(n12755), .B(n12754), .Z(n12837) );
  NAND U13131 ( .A(n35), .B(n12756), .Z(n12758) );
  XOR U13132 ( .A(b[9]), .B(a[165]), .Z(n12833) );
  NAND U13133 ( .A(n19598), .B(n12833), .Z(n12757) );
  NAND U13134 ( .A(n12758), .B(n12757), .Z(n12836) );
  XOR U13135 ( .A(n12837), .B(n12836), .Z(n12839) );
  XOR U13136 ( .A(n12838), .B(n12839), .Z(n12849) );
  NANDN U13137 ( .A(n12760), .B(n12759), .Z(n12764) );
  OR U13138 ( .A(n12762), .B(n12761), .Z(n12763) );
  AND U13139 ( .A(n12764), .B(n12763), .Z(n12848) );
  XNOR U13140 ( .A(n12849), .B(n12848), .Z(n12850) );
  NANDN U13141 ( .A(n12766), .B(n12765), .Z(n12770) );
  NANDN U13142 ( .A(n12768), .B(n12767), .Z(n12769) );
  NAND U13143 ( .A(n12770), .B(n12769), .Z(n12851) );
  XNOR U13144 ( .A(n12850), .B(n12851), .Z(n12796) );
  XOR U13145 ( .A(n12797), .B(n12796), .Z(n12855) );
  NANDN U13146 ( .A(n12772), .B(n12771), .Z(n12776) );
  NANDN U13147 ( .A(n12774), .B(n12773), .Z(n12775) );
  AND U13148 ( .A(n12776), .B(n12775), .Z(n12854) );
  XNOR U13149 ( .A(n12855), .B(n12854), .Z(n12856) );
  XOR U13150 ( .A(n12857), .B(n12856), .Z(n12789) );
  NANDN U13151 ( .A(n12778), .B(n12777), .Z(n12782) );
  NAND U13152 ( .A(n12780), .B(n12779), .Z(n12781) );
  AND U13153 ( .A(n12782), .B(n12781), .Z(n12788) );
  XNOR U13154 ( .A(n12789), .B(n12788), .Z(n12790) );
  XNOR U13155 ( .A(n12791), .B(n12790), .Z(n12860) );
  XNOR U13156 ( .A(sreg[413]), .B(n12860), .Z(n12862) );
  NANDN U13157 ( .A(sreg[412]), .B(n12783), .Z(n12787) );
  NAND U13158 ( .A(n12785), .B(n12784), .Z(n12786) );
  NAND U13159 ( .A(n12787), .B(n12786), .Z(n12861) );
  XNOR U13160 ( .A(n12862), .B(n12861), .Z(c[413]) );
  NANDN U13161 ( .A(n12789), .B(n12788), .Z(n12793) );
  NANDN U13162 ( .A(n12791), .B(n12790), .Z(n12792) );
  AND U13163 ( .A(n12793), .B(n12792), .Z(n12868) );
  NANDN U13164 ( .A(n12795), .B(n12794), .Z(n12799) );
  NAND U13165 ( .A(n12797), .B(n12796), .Z(n12798) );
  AND U13166 ( .A(n12799), .B(n12798), .Z(n12934) );
  NANDN U13167 ( .A(n12801), .B(n12800), .Z(n12805) );
  NANDN U13168 ( .A(n12803), .B(n12802), .Z(n12804) );
  AND U13169 ( .A(n12805), .B(n12804), .Z(n12900) );
  NAND U13170 ( .A(b[0]), .B(a[174]), .Z(n12806) );
  XNOR U13171 ( .A(b[1]), .B(n12806), .Z(n12808) );
  NANDN U13172 ( .A(b[0]), .B(a[173]), .Z(n12807) );
  NAND U13173 ( .A(n12808), .B(n12807), .Z(n12880) );
  NAND U13174 ( .A(n19808), .B(n12809), .Z(n12811) );
  XOR U13175 ( .A(b[13]), .B(a[162]), .Z(n12883) );
  NAND U13176 ( .A(n19768), .B(n12883), .Z(n12810) );
  AND U13177 ( .A(n12811), .B(n12810), .Z(n12878) );
  AND U13178 ( .A(b[15]), .B(a[158]), .Z(n12877) );
  XNOR U13179 ( .A(n12878), .B(n12877), .Z(n12879) );
  XNOR U13180 ( .A(n12880), .B(n12879), .Z(n12898) );
  NAND U13181 ( .A(n33), .B(n12812), .Z(n12814) );
  XOR U13182 ( .A(b[5]), .B(a[170]), .Z(n12889) );
  NAND U13183 ( .A(n19342), .B(n12889), .Z(n12813) );
  AND U13184 ( .A(n12814), .B(n12813), .Z(n12922) );
  NAND U13185 ( .A(n34), .B(n12815), .Z(n12817) );
  XOR U13186 ( .A(b[7]), .B(a[168]), .Z(n12892) );
  NAND U13187 ( .A(n19486), .B(n12892), .Z(n12816) );
  AND U13188 ( .A(n12817), .B(n12816), .Z(n12920) );
  NAND U13189 ( .A(n31), .B(n12818), .Z(n12820) );
  XOR U13190 ( .A(b[3]), .B(a[172]), .Z(n12895) );
  NAND U13191 ( .A(n32), .B(n12895), .Z(n12819) );
  NAND U13192 ( .A(n12820), .B(n12819), .Z(n12919) );
  XNOR U13193 ( .A(n12920), .B(n12919), .Z(n12921) );
  XOR U13194 ( .A(n12922), .B(n12921), .Z(n12899) );
  XOR U13195 ( .A(n12898), .B(n12899), .Z(n12901) );
  XOR U13196 ( .A(n12900), .B(n12901), .Z(n12872) );
  NANDN U13197 ( .A(n12822), .B(n12821), .Z(n12826) );
  OR U13198 ( .A(n12824), .B(n12823), .Z(n12825) );
  AND U13199 ( .A(n12826), .B(n12825), .Z(n12871) );
  XNOR U13200 ( .A(n12872), .B(n12871), .Z(n12874) );
  NAND U13201 ( .A(n12827), .B(n19724), .Z(n12829) );
  XOR U13202 ( .A(b[11]), .B(a[164]), .Z(n12904) );
  NAND U13203 ( .A(n19692), .B(n12904), .Z(n12828) );
  AND U13204 ( .A(n12829), .B(n12828), .Z(n12915) );
  NAND U13205 ( .A(n19838), .B(n12830), .Z(n12832) );
  XOR U13206 ( .A(b[15]), .B(a[160]), .Z(n12907) );
  NAND U13207 ( .A(n19805), .B(n12907), .Z(n12831) );
  AND U13208 ( .A(n12832), .B(n12831), .Z(n12914) );
  NAND U13209 ( .A(n35), .B(n12833), .Z(n12835) );
  XOR U13210 ( .A(b[9]), .B(a[166]), .Z(n12910) );
  NAND U13211 ( .A(n19598), .B(n12910), .Z(n12834) );
  NAND U13212 ( .A(n12835), .B(n12834), .Z(n12913) );
  XOR U13213 ( .A(n12914), .B(n12913), .Z(n12916) );
  XOR U13214 ( .A(n12915), .B(n12916), .Z(n12926) );
  NANDN U13215 ( .A(n12837), .B(n12836), .Z(n12841) );
  OR U13216 ( .A(n12839), .B(n12838), .Z(n12840) );
  AND U13217 ( .A(n12841), .B(n12840), .Z(n12925) );
  XNOR U13218 ( .A(n12926), .B(n12925), .Z(n12927) );
  NANDN U13219 ( .A(n12843), .B(n12842), .Z(n12847) );
  NANDN U13220 ( .A(n12845), .B(n12844), .Z(n12846) );
  NAND U13221 ( .A(n12847), .B(n12846), .Z(n12928) );
  XNOR U13222 ( .A(n12927), .B(n12928), .Z(n12873) );
  XOR U13223 ( .A(n12874), .B(n12873), .Z(n12932) );
  NANDN U13224 ( .A(n12849), .B(n12848), .Z(n12853) );
  NANDN U13225 ( .A(n12851), .B(n12850), .Z(n12852) );
  AND U13226 ( .A(n12853), .B(n12852), .Z(n12931) );
  XNOR U13227 ( .A(n12932), .B(n12931), .Z(n12933) );
  XOR U13228 ( .A(n12934), .B(n12933), .Z(n12866) );
  NANDN U13229 ( .A(n12855), .B(n12854), .Z(n12859) );
  NAND U13230 ( .A(n12857), .B(n12856), .Z(n12858) );
  AND U13231 ( .A(n12859), .B(n12858), .Z(n12865) );
  XNOR U13232 ( .A(n12866), .B(n12865), .Z(n12867) );
  XNOR U13233 ( .A(n12868), .B(n12867), .Z(n12937) );
  XNOR U13234 ( .A(sreg[414]), .B(n12937), .Z(n12939) );
  NANDN U13235 ( .A(sreg[413]), .B(n12860), .Z(n12864) );
  NAND U13236 ( .A(n12862), .B(n12861), .Z(n12863) );
  NAND U13237 ( .A(n12864), .B(n12863), .Z(n12938) );
  XNOR U13238 ( .A(n12939), .B(n12938), .Z(c[414]) );
  NANDN U13239 ( .A(n12866), .B(n12865), .Z(n12870) );
  NANDN U13240 ( .A(n12868), .B(n12867), .Z(n12869) );
  AND U13241 ( .A(n12870), .B(n12869), .Z(n12945) );
  NANDN U13242 ( .A(n12872), .B(n12871), .Z(n12876) );
  NAND U13243 ( .A(n12874), .B(n12873), .Z(n12875) );
  AND U13244 ( .A(n12876), .B(n12875), .Z(n13011) );
  NANDN U13245 ( .A(n12878), .B(n12877), .Z(n12882) );
  NANDN U13246 ( .A(n12880), .B(n12879), .Z(n12881) );
  AND U13247 ( .A(n12882), .B(n12881), .Z(n12977) );
  NAND U13248 ( .A(n19808), .B(n12883), .Z(n12885) );
  XOR U13249 ( .A(b[13]), .B(a[163]), .Z(n12963) );
  NAND U13250 ( .A(n19768), .B(n12963), .Z(n12884) );
  AND U13251 ( .A(n12885), .B(n12884), .Z(n12955) );
  AND U13252 ( .A(b[15]), .B(a[159]), .Z(n12954) );
  XNOR U13253 ( .A(n12955), .B(n12954), .Z(n12956) );
  NAND U13254 ( .A(b[0]), .B(a[175]), .Z(n12886) );
  XNOR U13255 ( .A(b[1]), .B(n12886), .Z(n12888) );
  NANDN U13256 ( .A(b[0]), .B(a[174]), .Z(n12887) );
  NAND U13257 ( .A(n12888), .B(n12887), .Z(n12957) );
  XNOR U13258 ( .A(n12956), .B(n12957), .Z(n12975) );
  NAND U13259 ( .A(n33), .B(n12889), .Z(n12891) );
  XOR U13260 ( .A(b[5]), .B(a[171]), .Z(n12966) );
  NAND U13261 ( .A(n19342), .B(n12966), .Z(n12890) );
  AND U13262 ( .A(n12891), .B(n12890), .Z(n12999) );
  NAND U13263 ( .A(n34), .B(n12892), .Z(n12894) );
  XOR U13264 ( .A(b[7]), .B(a[169]), .Z(n12969) );
  NAND U13265 ( .A(n19486), .B(n12969), .Z(n12893) );
  AND U13266 ( .A(n12894), .B(n12893), .Z(n12997) );
  NAND U13267 ( .A(n31), .B(n12895), .Z(n12897) );
  XOR U13268 ( .A(b[3]), .B(a[173]), .Z(n12972) );
  NAND U13269 ( .A(n32), .B(n12972), .Z(n12896) );
  NAND U13270 ( .A(n12897), .B(n12896), .Z(n12996) );
  XNOR U13271 ( .A(n12997), .B(n12996), .Z(n12998) );
  XOR U13272 ( .A(n12999), .B(n12998), .Z(n12976) );
  XOR U13273 ( .A(n12975), .B(n12976), .Z(n12978) );
  XOR U13274 ( .A(n12977), .B(n12978), .Z(n12949) );
  NANDN U13275 ( .A(n12899), .B(n12898), .Z(n12903) );
  OR U13276 ( .A(n12901), .B(n12900), .Z(n12902) );
  AND U13277 ( .A(n12903), .B(n12902), .Z(n12948) );
  XNOR U13278 ( .A(n12949), .B(n12948), .Z(n12951) );
  NAND U13279 ( .A(n12904), .B(n19724), .Z(n12906) );
  XOR U13280 ( .A(b[11]), .B(a[165]), .Z(n12981) );
  NAND U13281 ( .A(n19692), .B(n12981), .Z(n12905) );
  AND U13282 ( .A(n12906), .B(n12905), .Z(n12992) );
  NAND U13283 ( .A(n19838), .B(n12907), .Z(n12909) );
  XOR U13284 ( .A(b[15]), .B(a[161]), .Z(n12984) );
  NAND U13285 ( .A(n19805), .B(n12984), .Z(n12908) );
  AND U13286 ( .A(n12909), .B(n12908), .Z(n12991) );
  NAND U13287 ( .A(n35), .B(n12910), .Z(n12912) );
  XOR U13288 ( .A(b[9]), .B(a[167]), .Z(n12987) );
  NAND U13289 ( .A(n19598), .B(n12987), .Z(n12911) );
  NAND U13290 ( .A(n12912), .B(n12911), .Z(n12990) );
  XOR U13291 ( .A(n12991), .B(n12990), .Z(n12993) );
  XOR U13292 ( .A(n12992), .B(n12993), .Z(n13003) );
  NANDN U13293 ( .A(n12914), .B(n12913), .Z(n12918) );
  OR U13294 ( .A(n12916), .B(n12915), .Z(n12917) );
  AND U13295 ( .A(n12918), .B(n12917), .Z(n13002) );
  XNOR U13296 ( .A(n13003), .B(n13002), .Z(n13004) );
  NANDN U13297 ( .A(n12920), .B(n12919), .Z(n12924) );
  NANDN U13298 ( .A(n12922), .B(n12921), .Z(n12923) );
  NAND U13299 ( .A(n12924), .B(n12923), .Z(n13005) );
  XNOR U13300 ( .A(n13004), .B(n13005), .Z(n12950) );
  XOR U13301 ( .A(n12951), .B(n12950), .Z(n13009) );
  NANDN U13302 ( .A(n12926), .B(n12925), .Z(n12930) );
  NANDN U13303 ( .A(n12928), .B(n12927), .Z(n12929) );
  AND U13304 ( .A(n12930), .B(n12929), .Z(n13008) );
  XNOR U13305 ( .A(n13009), .B(n13008), .Z(n13010) );
  XOR U13306 ( .A(n13011), .B(n13010), .Z(n12943) );
  NANDN U13307 ( .A(n12932), .B(n12931), .Z(n12936) );
  NAND U13308 ( .A(n12934), .B(n12933), .Z(n12935) );
  AND U13309 ( .A(n12936), .B(n12935), .Z(n12942) );
  XNOR U13310 ( .A(n12943), .B(n12942), .Z(n12944) );
  XNOR U13311 ( .A(n12945), .B(n12944), .Z(n13014) );
  XNOR U13312 ( .A(sreg[415]), .B(n13014), .Z(n13016) );
  NANDN U13313 ( .A(sreg[414]), .B(n12937), .Z(n12941) );
  NAND U13314 ( .A(n12939), .B(n12938), .Z(n12940) );
  NAND U13315 ( .A(n12941), .B(n12940), .Z(n13015) );
  XNOR U13316 ( .A(n13016), .B(n13015), .Z(c[415]) );
  NANDN U13317 ( .A(n12943), .B(n12942), .Z(n12947) );
  NANDN U13318 ( .A(n12945), .B(n12944), .Z(n12946) );
  AND U13319 ( .A(n12947), .B(n12946), .Z(n13022) );
  NANDN U13320 ( .A(n12949), .B(n12948), .Z(n12953) );
  NAND U13321 ( .A(n12951), .B(n12950), .Z(n12952) );
  AND U13322 ( .A(n12953), .B(n12952), .Z(n13088) );
  NANDN U13323 ( .A(n12955), .B(n12954), .Z(n12959) );
  NANDN U13324 ( .A(n12957), .B(n12956), .Z(n12958) );
  AND U13325 ( .A(n12959), .B(n12958), .Z(n13075) );
  NAND U13326 ( .A(b[0]), .B(a[176]), .Z(n12960) );
  XNOR U13327 ( .A(b[1]), .B(n12960), .Z(n12962) );
  NANDN U13328 ( .A(b[0]), .B(a[175]), .Z(n12961) );
  NAND U13329 ( .A(n12962), .B(n12961), .Z(n13055) );
  NAND U13330 ( .A(n19808), .B(n12963), .Z(n12965) );
  XOR U13331 ( .A(b[13]), .B(a[164]), .Z(n13058) );
  NAND U13332 ( .A(n19768), .B(n13058), .Z(n12964) );
  AND U13333 ( .A(n12965), .B(n12964), .Z(n13053) );
  AND U13334 ( .A(b[15]), .B(a[160]), .Z(n13052) );
  XNOR U13335 ( .A(n13053), .B(n13052), .Z(n13054) );
  XNOR U13336 ( .A(n13055), .B(n13054), .Z(n13073) );
  NAND U13337 ( .A(n33), .B(n12966), .Z(n12968) );
  XOR U13338 ( .A(b[5]), .B(a[172]), .Z(n13064) );
  NAND U13339 ( .A(n19342), .B(n13064), .Z(n12967) );
  AND U13340 ( .A(n12968), .B(n12967), .Z(n13049) );
  NAND U13341 ( .A(n34), .B(n12969), .Z(n12971) );
  XOR U13342 ( .A(b[7]), .B(a[170]), .Z(n13067) );
  NAND U13343 ( .A(n19486), .B(n13067), .Z(n12970) );
  AND U13344 ( .A(n12971), .B(n12970), .Z(n13047) );
  NAND U13345 ( .A(n31), .B(n12972), .Z(n12974) );
  XOR U13346 ( .A(b[3]), .B(a[174]), .Z(n13070) );
  NAND U13347 ( .A(n32), .B(n13070), .Z(n12973) );
  NAND U13348 ( .A(n12974), .B(n12973), .Z(n13046) );
  XNOR U13349 ( .A(n13047), .B(n13046), .Z(n13048) );
  XOR U13350 ( .A(n13049), .B(n13048), .Z(n13074) );
  XOR U13351 ( .A(n13073), .B(n13074), .Z(n13076) );
  XOR U13352 ( .A(n13075), .B(n13076), .Z(n13026) );
  NANDN U13353 ( .A(n12976), .B(n12975), .Z(n12980) );
  OR U13354 ( .A(n12978), .B(n12977), .Z(n12979) );
  AND U13355 ( .A(n12980), .B(n12979), .Z(n13025) );
  XNOR U13356 ( .A(n13026), .B(n13025), .Z(n13028) );
  NAND U13357 ( .A(n12981), .B(n19724), .Z(n12983) );
  XOR U13358 ( .A(b[11]), .B(a[166]), .Z(n13031) );
  NAND U13359 ( .A(n19692), .B(n13031), .Z(n12982) );
  AND U13360 ( .A(n12983), .B(n12982), .Z(n13042) );
  NAND U13361 ( .A(n19838), .B(n12984), .Z(n12986) );
  XOR U13362 ( .A(b[15]), .B(a[162]), .Z(n13034) );
  NAND U13363 ( .A(n19805), .B(n13034), .Z(n12985) );
  AND U13364 ( .A(n12986), .B(n12985), .Z(n13041) );
  NAND U13365 ( .A(n35), .B(n12987), .Z(n12989) );
  XOR U13366 ( .A(b[9]), .B(a[168]), .Z(n13037) );
  NAND U13367 ( .A(n19598), .B(n13037), .Z(n12988) );
  NAND U13368 ( .A(n12989), .B(n12988), .Z(n13040) );
  XOR U13369 ( .A(n13041), .B(n13040), .Z(n13043) );
  XOR U13370 ( .A(n13042), .B(n13043), .Z(n13080) );
  NANDN U13371 ( .A(n12991), .B(n12990), .Z(n12995) );
  OR U13372 ( .A(n12993), .B(n12992), .Z(n12994) );
  AND U13373 ( .A(n12995), .B(n12994), .Z(n13079) );
  XNOR U13374 ( .A(n13080), .B(n13079), .Z(n13081) );
  NANDN U13375 ( .A(n12997), .B(n12996), .Z(n13001) );
  NANDN U13376 ( .A(n12999), .B(n12998), .Z(n13000) );
  NAND U13377 ( .A(n13001), .B(n13000), .Z(n13082) );
  XNOR U13378 ( .A(n13081), .B(n13082), .Z(n13027) );
  XOR U13379 ( .A(n13028), .B(n13027), .Z(n13086) );
  NANDN U13380 ( .A(n13003), .B(n13002), .Z(n13007) );
  NANDN U13381 ( .A(n13005), .B(n13004), .Z(n13006) );
  AND U13382 ( .A(n13007), .B(n13006), .Z(n13085) );
  XNOR U13383 ( .A(n13086), .B(n13085), .Z(n13087) );
  XOR U13384 ( .A(n13088), .B(n13087), .Z(n13020) );
  NANDN U13385 ( .A(n13009), .B(n13008), .Z(n13013) );
  NAND U13386 ( .A(n13011), .B(n13010), .Z(n13012) );
  AND U13387 ( .A(n13013), .B(n13012), .Z(n13019) );
  XNOR U13388 ( .A(n13020), .B(n13019), .Z(n13021) );
  XNOR U13389 ( .A(n13022), .B(n13021), .Z(n13091) );
  XNOR U13390 ( .A(sreg[416]), .B(n13091), .Z(n13093) );
  NANDN U13391 ( .A(sreg[415]), .B(n13014), .Z(n13018) );
  NAND U13392 ( .A(n13016), .B(n13015), .Z(n13017) );
  NAND U13393 ( .A(n13018), .B(n13017), .Z(n13092) );
  XNOR U13394 ( .A(n13093), .B(n13092), .Z(c[416]) );
  NANDN U13395 ( .A(n13020), .B(n13019), .Z(n13024) );
  NANDN U13396 ( .A(n13022), .B(n13021), .Z(n13023) );
  AND U13397 ( .A(n13024), .B(n13023), .Z(n13099) );
  NANDN U13398 ( .A(n13026), .B(n13025), .Z(n13030) );
  NAND U13399 ( .A(n13028), .B(n13027), .Z(n13029) );
  AND U13400 ( .A(n13030), .B(n13029), .Z(n13165) );
  NAND U13401 ( .A(n13031), .B(n19724), .Z(n13033) );
  XOR U13402 ( .A(b[11]), .B(a[167]), .Z(n13135) );
  NAND U13403 ( .A(n19692), .B(n13135), .Z(n13032) );
  AND U13404 ( .A(n13033), .B(n13032), .Z(n13146) );
  NAND U13405 ( .A(n19838), .B(n13034), .Z(n13036) );
  XOR U13406 ( .A(b[15]), .B(a[163]), .Z(n13138) );
  NAND U13407 ( .A(n19805), .B(n13138), .Z(n13035) );
  AND U13408 ( .A(n13036), .B(n13035), .Z(n13145) );
  NAND U13409 ( .A(n35), .B(n13037), .Z(n13039) );
  XOR U13410 ( .A(b[9]), .B(a[169]), .Z(n13141) );
  NAND U13411 ( .A(n19598), .B(n13141), .Z(n13038) );
  NAND U13412 ( .A(n13039), .B(n13038), .Z(n13144) );
  XOR U13413 ( .A(n13145), .B(n13144), .Z(n13147) );
  XOR U13414 ( .A(n13146), .B(n13147), .Z(n13157) );
  NANDN U13415 ( .A(n13041), .B(n13040), .Z(n13045) );
  OR U13416 ( .A(n13043), .B(n13042), .Z(n13044) );
  AND U13417 ( .A(n13045), .B(n13044), .Z(n13156) );
  XNOR U13418 ( .A(n13157), .B(n13156), .Z(n13158) );
  NANDN U13419 ( .A(n13047), .B(n13046), .Z(n13051) );
  NANDN U13420 ( .A(n13049), .B(n13048), .Z(n13050) );
  NAND U13421 ( .A(n13051), .B(n13050), .Z(n13159) );
  XNOR U13422 ( .A(n13158), .B(n13159), .Z(n13105) );
  NANDN U13423 ( .A(n13053), .B(n13052), .Z(n13057) );
  NANDN U13424 ( .A(n13055), .B(n13054), .Z(n13056) );
  AND U13425 ( .A(n13057), .B(n13056), .Z(n13131) );
  NAND U13426 ( .A(n19808), .B(n13058), .Z(n13060) );
  XOR U13427 ( .A(b[13]), .B(a[165]), .Z(n13114) );
  NAND U13428 ( .A(n19768), .B(n13114), .Z(n13059) );
  AND U13429 ( .A(n13060), .B(n13059), .Z(n13109) );
  AND U13430 ( .A(b[15]), .B(a[161]), .Z(n13108) );
  XNOR U13431 ( .A(n13109), .B(n13108), .Z(n13110) );
  NAND U13432 ( .A(b[0]), .B(a[177]), .Z(n13061) );
  XNOR U13433 ( .A(b[1]), .B(n13061), .Z(n13063) );
  NANDN U13434 ( .A(b[0]), .B(a[176]), .Z(n13062) );
  NAND U13435 ( .A(n13063), .B(n13062), .Z(n13111) );
  XNOR U13436 ( .A(n13110), .B(n13111), .Z(n13129) );
  NAND U13437 ( .A(n33), .B(n13064), .Z(n13066) );
  XOR U13438 ( .A(b[5]), .B(a[173]), .Z(n13120) );
  NAND U13439 ( .A(n19342), .B(n13120), .Z(n13065) );
  AND U13440 ( .A(n13066), .B(n13065), .Z(n13153) );
  NAND U13441 ( .A(n34), .B(n13067), .Z(n13069) );
  XOR U13442 ( .A(b[7]), .B(a[171]), .Z(n13123) );
  NAND U13443 ( .A(n19486), .B(n13123), .Z(n13068) );
  AND U13444 ( .A(n13069), .B(n13068), .Z(n13151) );
  NAND U13445 ( .A(n31), .B(n13070), .Z(n13072) );
  XOR U13446 ( .A(b[3]), .B(a[175]), .Z(n13126) );
  NAND U13447 ( .A(n32), .B(n13126), .Z(n13071) );
  NAND U13448 ( .A(n13072), .B(n13071), .Z(n13150) );
  XNOR U13449 ( .A(n13151), .B(n13150), .Z(n13152) );
  XOR U13450 ( .A(n13153), .B(n13152), .Z(n13130) );
  XOR U13451 ( .A(n13129), .B(n13130), .Z(n13132) );
  XOR U13452 ( .A(n13131), .B(n13132), .Z(n13103) );
  NANDN U13453 ( .A(n13074), .B(n13073), .Z(n13078) );
  OR U13454 ( .A(n13076), .B(n13075), .Z(n13077) );
  AND U13455 ( .A(n13078), .B(n13077), .Z(n13102) );
  XNOR U13456 ( .A(n13103), .B(n13102), .Z(n13104) );
  XOR U13457 ( .A(n13105), .B(n13104), .Z(n13163) );
  NANDN U13458 ( .A(n13080), .B(n13079), .Z(n13084) );
  NANDN U13459 ( .A(n13082), .B(n13081), .Z(n13083) );
  AND U13460 ( .A(n13084), .B(n13083), .Z(n13162) );
  XNOR U13461 ( .A(n13163), .B(n13162), .Z(n13164) );
  XOR U13462 ( .A(n13165), .B(n13164), .Z(n13097) );
  NANDN U13463 ( .A(n13086), .B(n13085), .Z(n13090) );
  NAND U13464 ( .A(n13088), .B(n13087), .Z(n13089) );
  AND U13465 ( .A(n13090), .B(n13089), .Z(n13096) );
  XNOR U13466 ( .A(n13097), .B(n13096), .Z(n13098) );
  XNOR U13467 ( .A(n13099), .B(n13098), .Z(n13168) );
  XNOR U13468 ( .A(sreg[417]), .B(n13168), .Z(n13170) );
  NANDN U13469 ( .A(sreg[416]), .B(n13091), .Z(n13095) );
  NAND U13470 ( .A(n13093), .B(n13092), .Z(n13094) );
  NAND U13471 ( .A(n13095), .B(n13094), .Z(n13169) );
  XNOR U13472 ( .A(n13170), .B(n13169), .Z(c[417]) );
  NANDN U13473 ( .A(n13097), .B(n13096), .Z(n13101) );
  NANDN U13474 ( .A(n13099), .B(n13098), .Z(n13100) );
  AND U13475 ( .A(n13101), .B(n13100), .Z(n13176) );
  NANDN U13476 ( .A(n13103), .B(n13102), .Z(n13107) );
  NAND U13477 ( .A(n13105), .B(n13104), .Z(n13106) );
  AND U13478 ( .A(n13107), .B(n13106), .Z(n13242) );
  NANDN U13479 ( .A(n13109), .B(n13108), .Z(n13113) );
  NANDN U13480 ( .A(n13111), .B(n13110), .Z(n13112) );
  AND U13481 ( .A(n13113), .B(n13112), .Z(n13208) );
  NAND U13482 ( .A(n19808), .B(n13114), .Z(n13116) );
  XOR U13483 ( .A(b[13]), .B(a[166]), .Z(n13194) );
  NAND U13484 ( .A(n19768), .B(n13194), .Z(n13115) );
  AND U13485 ( .A(n13116), .B(n13115), .Z(n13186) );
  AND U13486 ( .A(b[15]), .B(a[162]), .Z(n13185) );
  XNOR U13487 ( .A(n13186), .B(n13185), .Z(n13187) );
  NAND U13488 ( .A(b[0]), .B(a[178]), .Z(n13117) );
  XNOR U13489 ( .A(b[1]), .B(n13117), .Z(n13119) );
  NANDN U13490 ( .A(b[0]), .B(a[177]), .Z(n13118) );
  NAND U13491 ( .A(n13119), .B(n13118), .Z(n13188) );
  XNOR U13492 ( .A(n13187), .B(n13188), .Z(n13206) );
  NAND U13493 ( .A(n33), .B(n13120), .Z(n13122) );
  XOR U13494 ( .A(b[5]), .B(a[174]), .Z(n13197) );
  NAND U13495 ( .A(n19342), .B(n13197), .Z(n13121) );
  AND U13496 ( .A(n13122), .B(n13121), .Z(n13230) );
  NAND U13497 ( .A(n34), .B(n13123), .Z(n13125) );
  XOR U13498 ( .A(b[7]), .B(a[172]), .Z(n13200) );
  NAND U13499 ( .A(n19486), .B(n13200), .Z(n13124) );
  AND U13500 ( .A(n13125), .B(n13124), .Z(n13228) );
  NAND U13501 ( .A(n31), .B(n13126), .Z(n13128) );
  XOR U13502 ( .A(b[3]), .B(a[176]), .Z(n13203) );
  NAND U13503 ( .A(n32), .B(n13203), .Z(n13127) );
  NAND U13504 ( .A(n13128), .B(n13127), .Z(n13227) );
  XNOR U13505 ( .A(n13228), .B(n13227), .Z(n13229) );
  XOR U13506 ( .A(n13230), .B(n13229), .Z(n13207) );
  XOR U13507 ( .A(n13206), .B(n13207), .Z(n13209) );
  XOR U13508 ( .A(n13208), .B(n13209), .Z(n13180) );
  NANDN U13509 ( .A(n13130), .B(n13129), .Z(n13134) );
  OR U13510 ( .A(n13132), .B(n13131), .Z(n13133) );
  AND U13511 ( .A(n13134), .B(n13133), .Z(n13179) );
  XNOR U13512 ( .A(n13180), .B(n13179), .Z(n13182) );
  NAND U13513 ( .A(n13135), .B(n19724), .Z(n13137) );
  XOR U13514 ( .A(b[11]), .B(a[168]), .Z(n13212) );
  NAND U13515 ( .A(n19692), .B(n13212), .Z(n13136) );
  AND U13516 ( .A(n13137), .B(n13136), .Z(n13223) );
  NAND U13517 ( .A(n19838), .B(n13138), .Z(n13140) );
  XOR U13518 ( .A(b[15]), .B(a[164]), .Z(n13215) );
  NAND U13519 ( .A(n19805), .B(n13215), .Z(n13139) );
  AND U13520 ( .A(n13140), .B(n13139), .Z(n13222) );
  NAND U13521 ( .A(n35), .B(n13141), .Z(n13143) );
  XOR U13522 ( .A(b[9]), .B(a[170]), .Z(n13218) );
  NAND U13523 ( .A(n19598), .B(n13218), .Z(n13142) );
  NAND U13524 ( .A(n13143), .B(n13142), .Z(n13221) );
  XOR U13525 ( .A(n13222), .B(n13221), .Z(n13224) );
  XOR U13526 ( .A(n13223), .B(n13224), .Z(n13234) );
  NANDN U13527 ( .A(n13145), .B(n13144), .Z(n13149) );
  OR U13528 ( .A(n13147), .B(n13146), .Z(n13148) );
  AND U13529 ( .A(n13149), .B(n13148), .Z(n13233) );
  XNOR U13530 ( .A(n13234), .B(n13233), .Z(n13235) );
  NANDN U13531 ( .A(n13151), .B(n13150), .Z(n13155) );
  NANDN U13532 ( .A(n13153), .B(n13152), .Z(n13154) );
  NAND U13533 ( .A(n13155), .B(n13154), .Z(n13236) );
  XNOR U13534 ( .A(n13235), .B(n13236), .Z(n13181) );
  XOR U13535 ( .A(n13182), .B(n13181), .Z(n13240) );
  NANDN U13536 ( .A(n13157), .B(n13156), .Z(n13161) );
  NANDN U13537 ( .A(n13159), .B(n13158), .Z(n13160) );
  AND U13538 ( .A(n13161), .B(n13160), .Z(n13239) );
  XNOR U13539 ( .A(n13240), .B(n13239), .Z(n13241) );
  XOR U13540 ( .A(n13242), .B(n13241), .Z(n13174) );
  NANDN U13541 ( .A(n13163), .B(n13162), .Z(n13167) );
  NAND U13542 ( .A(n13165), .B(n13164), .Z(n13166) );
  AND U13543 ( .A(n13167), .B(n13166), .Z(n13173) );
  XNOR U13544 ( .A(n13174), .B(n13173), .Z(n13175) );
  XNOR U13545 ( .A(n13176), .B(n13175), .Z(n13245) );
  XNOR U13546 ( .A(sreg[418]), .B(n13245), .Z(n13247) );
  NANDN U13547 ( .A(sreg[417]), .B(n13168), .Z(n13172) );
  NAND U13548 ( .A(n13170), .B(n13169), .Z(n13171) );
  NAND U13549 ( .A(n13172), .B(n13171), .Z(n13246) );
  XNOR U13550 ( .A(n13247), .B(n13246), .Z(c[418]) );
  NANDN U13551 ( .A(n13174), .B(n13173), .Z(n13178) );
  NANDN U13552 ( .A(n13176), .B(n13175), .Z(n13177) );
  AND U13553 ( .A(n13178), .B(n13177), .Z(n13253) );
  NANDN U13554 ( .A(n13180), .B(n13179), .Z(n13184) );
  NAND U13555 ( .A(n13182), .B(n13181), .Z(n13183) );
  AND U13556 ( .A(n13184), .B(n13183), .Z(n13319) );
  NANDN U13557 ( .A(n13186), .B(n13185), .Z(n13190) );
  NANDN U13558 ( .A(n13188), .B(n13187), .Z(n13189) );
  AND U13559 ( .A(n13190), .B(n13189), .Z(n13285) );
  NAND U13560 ( .A(b[0]), .B(a[179]), .Z(n13191) );
  XNOR U13561 ( .A(b[1]), .B(n13191), .Z(n13193) );
  NANDN U13562 ( .A(b[0]), .B(a[178]), .Z(n13192) );
  NAND U13563 ( .A(n13193), .B(n13192), .Z(n13265) );
  NAND U13564 ( .A(n19808), .B(n13194), .Z(n13196) );
  XOR U13565 ( .A(b[13]), .B(a[167]), .Z(n13271) );
  NAND U13566 ( .A(n19768), .B(n13271), .Z(n13195) );
  AND U13567 ( .A(n13196), .B(n13195), .Z(n13263) );
  AND U13568 ( .A(b[15]), .B(a[163]), .Z(n13262) );
  XNOR U13569 ( .A(n13263), .B(n13262), .Z(n13264) );
  XNOR U13570 ( .A(n13265), .B(n13264), .Z(n13283) );
  NAND U13571 ( .A(n33), .B(n13197), .Z(n13199) );
  XOR U13572 ( .A(b[5]), .B(a[175]), .Z(n13274) );
  NAND U13573 ( .A(n19342), .B(n13274), .Z(n13198) );
  AND U13574 ( .A(n13199), .B(n13198), .Z(n13307) );
  NAND U13575 ( .A(n34), .B(n13200), .Z(n13202) );
  XOR U13576 ( .A(b[7]), .B(a[173]), .Z(n13277) );
  NAND U13577 ( .A(n19486), .B(n13277), .Z(n13201) );
  AND U13578 ( .A(n13202), .B(n13201), .Z(n13305) );
  NAND U13579 ( .A(n31), .B(n13203), .Z(n13205) );
  XOR U13580 ( .A(b[3]), .B(a[177]), .Z(n13280) );
  NAND U13581 ( .A(n32), .B(n13280), .Z(n13204) );
  NAND U13582 ( .A(n13205), .B(n13204), .Z(n13304) );
  XNOR U13583 ( .A(n13305), .B(n13304), .Z(n13306) );
  XOR U13584 ( .A(n13307), .B(n13306), .Z(n13284) );
  XOR U13585 ( .A(n13283), .B(n13284), .Z(n13286) );
  XOR U13586 ( .A(n13285), .B(n13286), .Z(n13257) );
  NANDN U13587 ( .A(n13207), .B(n13206), .Z(n13211) );
  OR U13588 ( .A(n13209), .B(n13208), .Z(n13210) );
  AND U13589 ( .A(n13211), .B(n13210), .Z(n13256) );
  XNOR U13590 ( .A(n13257), .B(n13256), .Z(n13259) );
  NAND U13591 ( .A(n13212), .B(n19724), .Z(n13214) );
  XOR U13592 ( .A(b[11]), .B(a[169]), .Z(n13289) );
  NAND U13593 ( .A(n19692), .B(n13289), .Z(n13213) );
  AND U13594 ( .A(n13214), .B(n13213), .Z(n13300) );
  NAND U13595 ( .A(n19838), .B(n13215), .Z(n13217) );
  XOR U13596 ( .A(b[15]), .B(a[165]), .Z(n13292) );
  NAND U13597 ( .A(n19805), .B(n13292), .Z(n13216) );
  AND U13598 ( .A(n13217), .B(n13216), .Z(n13299) );
  NAND U13599 ( .A(n35), .B(n13218), .Z(n13220) );
  XOR U13600 ( .A(b[9]), .B(a[171]), .Z(n13295) );
  NAND U13601 ( .A(n19598), .B(n13295), .Z(n13219) );
  NAND U13602 ( .A(n13220), .B(n13219), .Z(n13298) );
  XOR U13603 ( .A(n13299), .B(n13298), .Z(n13301) );
  XOR U13604 ( .A(n13300), .B(n13301), .Z(n13311) );
  NANDN U13605 ( .A(n13222), .B(n13221), .Z(n13226) );
  OR U13606 ( .A(n13224), .B(n13223), .Z(n13225) );
  AND U13607 ( .A(n13226), .B(n13225), .Z(n13310) );
  XNOR U13608 ( .A(n13311), .B(n13310), .Z(n13312) );
  NANDN U13609 ( .A(n13228), .B(n13227), .Z(n13232) );
  NANDN U13610 ( .A(n13230), .B(n13229), .Z(n13231) );
  NAND U13611 ( .A(n13232), .B(n13231), .Z(n13313) );
  XNOR U13612 ( .A(n13312), .B(n13313), .Z(n13258) );
  XOR U13613 ( .A(n13259), .B(n13258), .Z(n13317) );
  NANDN U13614 ( .A(n13234), .B(n13233), .Z(n13238) );
  NANDN U13615 ( .A(n13236), .B(n13235), .Z(n13237) );
  AND U13616 ( .A(n13238), .B(n13237), .Z(n13316) );
  XNOR U13617 ( .A(n13317), .B(n13316), .Z(n13318) );
  XOR U13618 ( .A(n13319), .B(n13318), .Z(n13251) );
  NANDN U13619 ( .A(n13240), .B(n13239), .Z(n13244) );
  NAND U13620 ( .A(n13242), .B(n13241), .Z(n13243) );
  AND U13621 ( .A(n13244), .B(n13243), .Z(n13250) );
  XNOR U13622 ( .A(n13251), .B(n13250), .Z(n13252) );
  XNOR U13623 ( .A(n13253), .B(n13252), .Z(n13322) );
  XNOR U13624 ( .A(sreg[419]), .B(n13322), .Z(n13324) );
  NANDN U13625 ( .A(sreg[418]), .B(n13245), .Z(n13249) );
  NAND U13626 ( .A(n13247), .B(n13246), .Z(n13248) );
  NAND U13627 ( .A(n13249), .B(n13248), .Z(n13323) );
  XNOR U13628 ( .A(n13324), .B(n13323), .Z(c[419]) );
  NANDN U13629 ( .A(n13251), .B(n13250), .Z(n13255) );
  NANDN U13630 ( .A(n13253), .B(n13252), .Z(n13254) );
  AND U13631 ( .A(n13255), .B(n13254), .Z(n13330) );
  NANDN U13632 ( .A(n13257), .B(n13256), .Z(n13261) );
  NAND U13633 ( .A(n13259), .B(n13258), .Z(n13260) );
  AND U13634 ( .A(n13261), .B(n13260), .Z(n13396) );
  NANDN U13635 ( .A(n13263), .B(n13262), .Z(n13267) );
  NANDN U13636 ( .A(n13265), .B(n13264), .Z(n13266) );
  AND U13637 ( .A(n13267), .B(n13266), .Z(n13362) );
  NAND U13638 ( .A(b[0]), .B(a[180]), .Z(n13268) );
  XNOR U13639 ( .A(b[1]), .B(n13268), .Z(n13270) );
  NANDN U13640 ( .A(b[0]), .B(a[179]), .Z(n13269) );
  NAND U13641 ( .A(n13270), .B(n13269), .Z(n13342) );
  NAND U13642 ( .A(n19808), .B(n13271), .Z(n13273) );
  XOR U13643 ( .A(b[13]), .B(a[168]), .Z(n13348) );
  NAND U13644 ( .A(n19768), .B(n13348), .Z(n13272) );
  AND U13645 ( .A(n13273), .B(n13272), .Z(n13340) );
  AND U13646 ( .A(b[15]), .B(a[164]), .Z(n13339) );
  XNOR U13647 ( .A(n13340), .B(n13339), .Z(n13341) );
  XNOR U13648 ( .A(n13342), .B(n13341), .Z(n13360) );
  NAND U13649 ( .A(n33), .B(n13274), .Z(n13276) );
  XOR U13650 ( .A(b[5]), .B(a[176]), .Z(n13351) );
  NAND U13651 ( .A(n19342), .B(n13351), .Z(n13275) );
  AND U13652 ( .A(n13276), .B(n13275), .Z(n13384) );
  NAND U13653 ( .A(n34), .B(n13277), .Z(n13279) );
  XOR U13654 ( .A(b[7]), .B(a[174]), .Z(n13354) );
  NAND U13655 ( .A(n19486), .B(n13354), .Z(n13278) );
  AND U13656 ( .A(n13279), .B(n13278), .Z(n13382) );
  NAND U13657 ( .A(n31), .B(n13280), .Z(n13282) );
  XOR U13658 ( .A(b[3]), .B(a[178]), .Z(n13357) );
  NAND U13659 ( .A(n32), .B(n13357), .Z(n13281) );
  NAND U13660 ( .A(n13282), .B(n13281), .Z(n13381) );
  XNOR U13661 ( .A(n13382), .B(n13381), .Z(n13383) );
  XOR U13662 ( .A(n13384), .B(n13383), .Z(n13361) );
  XOR U13663 ( .A(n13360), .B(n13361), .Z(n13363) );
  XOR U13664 ( .A(n13362), .B(n13363), .Z(n13334) );
  NANDN U13665 ( .A(n13284), .B(n13283), .Z(n13288) );
  OR U13666 ( .A(n13286), .B(n13285), .Z(n13287) );
  AND U13667 ( .A(n13288), .B(n13287), .Z(n13333) );
  XNOR U13668 ( .A(n13334), .B(n13333), .Z(n13336) );
  NAND U13669 ( .A(n13289), .B(n19724), .Z(n13291) );
  XOR U13670 ( .A(b[11]), .B(a[170]), .Z(n13366) );
  NAND U13671 ( .A(n19692), .B(n13366), .Z(n13290) );
  AND U13672 ( .A(n13291), .B(n13290), .Z(n13377) );
  NAND U13673 ( .A(n19838), .B(n13292), .Z(n13294) );
  XOR U13674 ( .A(b[15]), .B(a[166]), .Z(n13369) );
  NAND U13675 ( .A(n19805), .B(n13369), .Z(n13293) );
  AND U13676 ( .A(n13294), .B(n13293), .Z(n13376) );
  NAND U13677 ( .A(n35), .B(n13295), .Z(n13297) );
  XOR U13678 ( .A(b[9]), .B(a[172]), .Z(n13372) );
  NAND U13679 ( .A(n19598), .B(n13372), .Z(n13296) );
  NAND U13680 ( .A(n13297), .B(n13296), .Z(n13375) );
  XOR U13681 ( .A(n13376), .B(n13375), .Z(n13378) );
  XOR U13682 ( .A(n13377), .B(n13378), .Z(n13388) );
  NANDN U13683 ( .A(n13299), .B(n13298), .Z(n13303) );
  OR U13684 ( .A(n13301), .B(n13300), .Z(n13302) );
  AND U13685 ( .A(n13303), .B(n13302), .Z(n13387) );
  XNOR U13686 ( .A(n13388), .B(n13387), .Z(n13389) );
  NANDN U13687 ( .A(n13305), .B(n13304), .Z(n13309) );
  NANDN U13688 ( .A(n13307), .B(n13306), .Z(n13308) );
  NAND U13689 ( .A(n13309), .B(n13308), .Z(n13390) );
  XNOR U13690 ( .A(n13389), .B(n13390), .Z(n13335) );
  XOR U13691 ( .A(n13336), .B(n13335), .Z(n13394) );
  NANDN U13692 ( .A(n13311), .B(n13310), .Z(n13315) );
  NANDN U13693 ( .A(n13313), .B(n13312), .Z(n13314) );
  AND U13694 ( .A(n13315), .B(n13314), .Z(n13393) );
  XNOR U13695 ( .A(n13394), .B(n13393), .Z(n13395) );
  XOR U13696 ( .A(n13396), .B(n13395), .Z(n13328) );
  NANDN U13697 ( .A(n13317), .B(n13316), .Z(n13321) );
  NAND U13698 ( .A(n13319), .B(n13318), .Z(n13320) );
  AND U13699 ( .A(n13321), .B(n13320), .Z(n13327) );
  XNOR U13700 ( .A(n13328), .B(n13327), .Z(n13329) );
  XNOR U13701 ( .A(n13330), .B(n13329), .Z(n13399) );
  XNOR U13702 ( .A(sreg[420]), .B(n13399), .Z(n13401) );
  NANDN U13703 ( .A(sreg[419]), .B(n13322), .Z(n13326) );
  NAND U13704 ( .A(n13324), .B(n13323), .Z(n13325) );
  NAND U13705 ( .A(n13326), .B(n13325), .Z(n13400) );
  XNOR U13706 ( .A(n13401), .B(n13400), .Z(c[420]) );
  NANDN U13707 ( .A(n13328), .B(n13327), .Z(n13332) );
  NANDN U13708 ( .A(n13330), .B(n13329), .Z(n13331) );
  AND U13709 ( .A(n13332), .B(n13331), .Z(n13407) );
  NANDN U13710 ( .A(n13334), .B(n13333), .Z(n13338) );
  NAND U13711 ( .A(n13336), .B(n13335), .Z(n13337) );
  AND U13712 ( .A(n13338), .B(n13337), .Z(n13473) );
  NANDN U13713 ( .A(n13340), .B(n13339), .Z(n13344) );
  NANDN U13714 ( .A(n13342), .B(n13341), .Z(n13343) );
  AND U13715 ( .A(n13344), .B(n13343), .Z(n13439) );
  NAND U13716 ( .A(b[0]), .B(a[181]), .Z(n13345) );
  XNOR U13717 ( .A(b[1]), .B(n13345), .Z(n13347) );
  NANDN U13718 ( .A(b[0]), .B(a[180]), .Z(n13346) );
  NAND U13719 ( .A(n13347), .B(n13346), .Z(n13419) );
  NAND U13720 ( .A(n19808), .B(n13348), .Z(n13350) );
  XOR U13721 ( .A(b[13]), .B(a[169]), .Z(n13425) );
  NAND U13722 ( .A(n19768), .B(n13425), .Z(n13349) );
  AND U13723 ( .A(n13350), .B(n13349), .Z(n13417) );
  AND U13724 ( .A(b[15]), .B(a[165]), .Z(n13416) );
  XNOR U13725 ( .A(n13417), .B(n13416), .Z(n13418) );
  XNOR U13726 ( .A(n13419), .B(n13418), .Z(n13437) );
  NAND U13727 ( .A(n33), .B(n13351), .Z(n13353) );
  XOR U13728 ( .A(b[5]), .B(a[177]), .Z(n13428) );
  NAND U13729 ( .A(n19342), .B(n13428), .Z(n13352) );
  AND U13730 ( .A(n13353), .B(n13352), .Z(n13461) );
  NAND U13731 ( .A(n34), .B(n13354), .Z(n13356) );
  XOR U13732 ( .A(b[7]), .B(a[175]), .Z(n13431) );
  NAND U13733 ( .A(n19486), .B(n13431), .Z(n13355) );
  AND U13734 ( .A(n13356), .B(n13355), .Z(n13459) );
  NAND U13735 ( .A(n31), .B(n13357), .Z(n13359) );
  XOR U13736 ( .A(b[3]), .B(a[179]), .Z(n13434) );
  NAND U13737 ( .A(n32), .B(n13434), .Z(n13358) );
  NAND U13738 ( .A(n13359), .B(n13358), .Z(n13458) );
  XNOR U13739 ( .A(n13459), .B(n13458), .Z(n13460) );
  XOR U13740 ( .A(n13461), .B(n13460), .Z(n13438) );
  XOR U13741 ( .A(n13437), .B(n13438), .Z(n13440) );
  XOR U13742 ( .A(n13439), .B(n13440), .Z(n13411) );
  NANDN U13743 ( .A(n13361), .B(n13360), .Z(n13365) );
  OR U13744 ( .A(n13363), .B(n13362), .Z(n13364) );
  AND U13745 ( .A(n13365), .B(n13364), .Z(n13410) );
  XNOR U13746 ( .A(n13411), .B(n13410), .Z(n13413) );
  NAND U13747 ( .A(n13366), .B(n19724), .Z(n13368) );
  XOR U13748 ( .A(b[11]), .B(a[171]), .Z(n13443) );
  NAND U13749 ( .A(n19692), .B(n13443), .Z(n13367) );
  AND U13750 ( .A(n13368), .B(n13367), .Z(n13454) );
  NAND U13751 ( .A(n19838), .B(n13369), .Z(n13371) );
  XOR U13752 ( .A(b[15]), .B(a[167]), .Z(n13446) );
  NAND U13753 ( .A(n19805), .B(n13446), .Z(n13370) );
  AND U13754 ( .A(n13371), .B(n13370), .Z(n13453) );
  NAND U13755 ( .A(n35), .B(n13372), .Z(n13374) );
  XOR U13756 ( .A(b[9]), .B(a[173]), .Z(n13449) );
  NAND U13757 ( .A(n19598), .B(n13449), .Z(n13373) );
  NAND U13758 ( .A(n13374), .B(n13373), .Z(n13452) );
  XOR U13759 ( .A(n13453), .B(n13452), .Z(n13455) );
  XOR U13760 ( .A(n13454), .B(n13455), .Z(n13465) );
  NANDN U13761 ( .A(n13376), .B(n13375), .Z(n13380) );
  OR U13762 ( .A(n13378), .B(n13377), .Z(n13379) );
  AND U13763 ( .A(n13380), .B(n13379), .Z(n13464) );
  XNOR U13764 ( .A(n13465), .B(n13464), .Z(n13466) );
  NANDN U13765 ( .A(n13382), .B(n13381), .Z(n13386) );
  NANDN U13766 ( .A(n13384), .B(n13383), .Z(n13385) );
  NAND U13767 ( .A(n13386), .B(n13385), .Z(n13467) );
  XNOR U13768 ( .A(n13466), .B(n13467), .Z(n13412) );
  XOR U13769 ( .A(n13413), .B(n13412), .Z(n13471) );
  NANDN U13770 ( .A(n13388), .B(n13387), .Z(n13392) );
  NANDN U13771 ( .A(n13390), .B(n13389), .Z(n13391) );
  AND U13772 ( .A(n13392), .B(n13391), .Z(n13470) );
  XNOR U13773 ( .A(n13471), .B(n13470), .Z(n13472) );
  XOR U13774 ( .A(n13473), .B(n13472), .Z(n13405) );
  NANDN U13775 ( .A(n13394), .B(n13393), .Z(n13398) );
  NAND U13776 ( .A(n13396), .B(n13395), .Z(n13397) );
  AND U13777 ( .A(n13398), .B(n13397), .Z(n13404) );
  XNOR U13778 ( .A(n13405), .B(n13404), .Z(n13406) );
  XNOR U13779 ( .A(n13407), .B(n13406), .Z(n13476) );
  XNOR U13780 ( .A(sreg[421]), .B(n13476), .Z(n13478) );
  NANDN U13781 ( .A(sreg[420]), .B(n13399), .Z(n13403) );
  NAND U13782 ( .A(n13401), .B(n13400), .Z(n13402) );
  NAND U13783 ( .A(n13403), .B(n13402), .Z(n13477) );
  XNOR U13784 ( .A(n13478), .B(n13477), .Z(c[421]) );
  NANDN U13785 ( .A(n13405), .B(n13404), .Z(n13409) );
  NANDN U13786 ( .A(n13407), .B(n13406), .Z(n13408) );
  AND U13787 ( .A(n13409), .B(n13408), .Z(n13484) );
  NANDN U13788 ( .A(n13411), .B(n13410), .Z(n13415) );
  NAND U13789 ( .A(n13413), .B(n13412), .Z(n13414) );
  AND U13790 ( .A(n13415), .B(n13414), .Z(n13550) );
  NANDN U13791 ( .A(n13417), .B(n13416), .Z(n13421) );
  NANDN U13792 ( .A(n13419), .B(n13418), .Z(n13420) );
  AND U13793 ( .A(n13421), .B(n13420), .Z(n13516) );
  NAND U13794 ( .A(b[0]), .B(a[182]), .Z(n13422) );
  XNOR U13795 ( .A(b[1]), .B(n13422), .Z(n13424) );
  NANDN U13796 ( .A(b[0]), .B(a[181]), .Z(n13423) );
  NAND U13797 ( .A(n13424), .B(n13423), .Z(n13496) );
  NAND U13798 ( .A(n19808), .B(n13425), .Z(n13427) );
  XOR U13799 ( .A(b[13]), .B(a[170]), .Z(n13502) );
  NAND U13800 ( .A(n19768), .B(n13502), .Z(n13426) );
  AND U13801 ( .A(n13427), .B(n13426), .Z(n13494) );
  AND U13802 ( .A(b[15]), .B(a[166]), .Z(n13493) );
  XNOR U13803 ( .A(n13494), .B(n13493), .Z(n13495) );
  XNOR U13804 ( .A(n13496), .B(n13495), .Z(n13514) );
  NAND U13805 ( .A(n33), .B(n13428), .Z(n13430) );
  XOR U13806 ( .A(b[5]), .B(a[178]), .Z(n13505) );
  NAND U13807 ( .A(n19342), .B(n13505), .Z(n13429) );
  AND U13808 ( .A(n13430), .B(n13429), .Z(n13538) );
  NAND U13809 ( .A(n34), .B(n13431), .Z(n13433) );
  XOR U13810 ( .A(b[7]), .B(a[176]), .Z(n13508) );
  NAND U13811 ( .A(n19486), .B(n13508), .Z(n13432) );
  AND U13812 ( .A(n13433), .B(n13432), .Z(n13536) );
  NAND U13813 ( .A(n31), .B(n13434), .Z(n13436) );
  XOR U13814 ( .A(b[3]), .B(a[180]), .Z(n13511) );
  NAND U13815 ( .A(n32), .B(n13511), .Z(n13435) );
  NAND U13816 ( .A(n13436), .B(n13435), .Z(n13535) );
  XNOR U13817 ( .A(n13536), .B(n13535), .Z(n13537) );
  XOR U13818 ( .A(n13538), .B(n13537), .Z(n13515) );
  XOR U13819 ( .A(n13514), .B(n13515), .Z(n13517) );
  XOR U13820 ( .A(n13516), .B(n13517), .Z(n13488) );
  NANDN U13821 ( .A(n13438), .B(n13437), .Z(n13442) );
  OR U13822 ( .A(n13440), .B(n13439), .Z(n13441) );
  AND U13823 ( .A(n13442), .B(n13441), .Z(n13487) );
  XNOR U13824 ( .A(n13488), .B(n13487), .Z(n13490) );
  NAND U13825 ( .A(n13443), .B(n19724), .Z(n13445) );
  XOR U13826 ( .A(b[11]), .B(a[172]), .Z(n13520) );
  NAND U13827 ( .A(n19692), .B(n13520), .Z(n13444) );
  AND U13828 ( .A(n13445), .B(n13444), .Z(n13531) );
  NAND U13829 ( .A(n19838), .B(n13446), .Z(n13448) );
  XOR U13830 ( .A(b[15]), .B(a[168]), .Z(n13523) );
  NAND U13831 ( .A(n19805), .B(n13523), .Z(n13447) );
  AND U13832 ( .A(n13448), .B(n13447), .Z(n13530) );
  NAND U13833 ( .A(n35), .B(n13449), .Z(n13451) );
  XOR U13834 ( .A(b[9]), .B(a[174]), .Z(n13526) );
  NAND U13835 ( .A(n19598), .B(n13526), .Z(n13450) );
  NAND U13836 ( .A(n13451), .B(n13450), .Z(n13529) );
  XOR U13837 ( .A(n13530), .B(n13529), .Z(n13532) );
  XOR U13838 ( .A(n13531), .B(n13532), .Z(n13542) );
  NANDN U13839 ( .A(n13453), .B(n13452), .Z(n13457) );
  OR U13840 ( .A(n13455), .B(n13454), .Z(n13456) );
  AND U13841 ( .A(n13457), .B(n13456), .Z(n13541) );
  XNOR U13842 ( .A(n13542), .B(n13541), .Z(n13543) );
  NANDN U13843 ( .A(n13459), .B(n13458), .Z(n13463) );
  NANDN U13844 ( .A(n13461), .B(n13460), .Z(n13462) );
  NAND U13845 ( .A(n13463), .B(n13462), .Z(n13544) );
  XNOR U13846 ( .A(n13543), .B(n13544), .Z(n13489) );
  XOR U13847 ( .A(n13490), .B(n13489), .Z(n13548) );
  NANDN U13848 ( .A(n13465), .B(n13464), .Z(n13469) );
  NANDN U13849 ( .A(n13467), .B(n13466), .Z(n13468) );
  AND U13850 ( .A(n13469), .B(n13468), .Z(n13547) );
  XNOR U13851 ( .A(n13548), .B(n13547), .Z(n13549) );
  XOR U13852 ( .A(n13550), .B(n13549), .Z(n13482) );
  NANDN U13853 ( .A(n13471), .B(n13470), .Z(n13475) );
  NAND U13854 ( .A(n13473), .B(n13472), .Z(n13474) );
  AND U13855 ( .A(n13475), .B(n13474), .Z(n13481) );
  XNOR U13856 ( .A(n13482), .B(n13481), .Z(n13483) );
  XNOR U13857 ( .A(n13484), .B(n13483), .Z(n13553) );
  XNOR U13858 ( .A(sreg[422]), .B(n13553), .Z(n13555) );
  NANDN U13859 ( .A(sreg[421]), .B(n13476), .Z(n13480) );
  NAND U13860 ( .A(n13478), .B(n13477), .Z(n13479) );
  NAND U13861 ( .A(n13480), .B(n13479), .Z(n13554) );
  XNOR U13862 ( .A(n13555), .B(n13554), .Z(c[422]) );
  NANDN U13863 ( .A(n13482), .B(n13481), .Z(n13486) );
  NANDN U13864 ( .A(n13484), .B(n13483), .Z(n13485) );
  AND U13865 ( .A(n13486), .B(n13485), .Z(n13561) );
  NANDN U13866 ( .A(n13488), .B(n13487), .Z(n13492) );
  NAND U13867 ( .A(n13490), .B(n13489), .Z(n13491) );
  AND U13868 ( .A(n13492), .B(n13491), .Z(n13627) );
  NANDN U13869 ( .A(n13494), .B(n13493), .Z(n13498) );
  NANDN U13870 ( .A(n13496), .B(n13495), .Z(n13497) );
  AND U13871 ( .A(n13498), .B(n13497), .Z(n13593) );
  NAND U13872 ( .A(b[0]), .B(a[183]), .Z(n13499) );
  XNOR U13873 ( .A(b[1]), .B(n13499), .Z(n13501) );
  NANDN U13874 ( .A(b[0]), .B(a[182]), .Z(n13500) );
  NAND U13875 ( .A(n13501), .B(n13500), .Z(n13573) );
  NAND U13876 ( .A(n19808), .B(n13502), .Z(n13504) );
  XOR U13877 ( .A(b[13]), .B(a[171]), .Z(n13579) );
  NAND U13878 ( .A(n19768), .B(n13579), .Z(n13503) );
  AND U13879 ( .A(n13504), .B(n13503), .Z(n13571) );
  AND U13880 ( .A(b[15]), .B(a[167]), .Z(n13570) );
  XNOR U13881 ( .A(n13571), .B(n13570), .Z(n13572) );
  XNOR U13882 ( .A(n13573), .B(n13572), .Z(n13591) );
  NAND U13883 ( .A(n33), .B(n13505), .Z(n13507) );
  XOR U13884 ( .A(b[5]), .B(a[179]), .Z(n13582) );
  NAND U13885 ( .A(n19342), .B(n13582), .Z(n13506) );
  AND U13886 ( .A(n13507), .B(n13506), .Z(n13615) );
  NAND U13887 ( .A(n34), .B(n13508), .Z(n13510) );
  XOR U13888 ( .A(b[7]), .B(a[177]), .Z(n13585) );
  NAND U13889 ( .A(n19486), .B(n13585), .Z(n13509) );
  AND U13890 ( .A(n13510), .B(n13509), .Z(n13613) );
  NAND U13891 ( .A(n31), .B(n13511), .Z(n13513) );
  XOR U13892 ( .A(b[3]), .B(a[181]), .Z(n13588) );
  NAND U13893 ( .A(n32), .B(n13588), .Z(n13512) );
  NAND U13894 ( .A(n13513), .B(n13512), .Z(n13612) );
  XNOR U13895 ( .A(n13613), .B(n13612), .Z(n13614) );
  XOR U13896 ( .A(n13615), .B(n13614), .Z(n13592) );
  XOR U13897 ( .A(n13591), .B(n13592), .Z(n13594) );
  XOR U13898 ( .A(n13593), .B(n13594), .Z(n13565) );
  NANDN U13899 ( .A(n13515), .B(n13514), .Z(n13519) );
  OR U13900 ( .A(n13517), .B(n13516), .Z(n13518) );
  AND U13901 ( .A(n13519), .B(n13518), .Z(n13564) );
  XNOR U13902 ( .A(n13565), .B(n13564), .Z(n13567) );
  NAND U13903 ( .A(n13520), .B(n19724), .Z(n13522) );
  XOR U13904 ( .A(b[11]), .B(a[173]), .Z(n13597) );
  NAND U13905 ( .A(n19692), .B(n13597), .Z(n13521) );
  AND U13906 ( .A(n13522), .B(n13521), .Z(n13608) );
  NAND U13907 ( .A(n19838), .B(n13523), .Z(n13525) );
  XOR U13908 ( .A(b[15]), .B(a[169]), .Z(n13600) );
  NAND U13909 ( .A(n19805), .B(n13600), .Z(n13524) );
  AND U13910 ( .A(n13525), .B(n13524), .Z(n13607) );
  NAND U13911 ( .A(n35), .B(n13526), .Z(n13528) );
  XOR U13912 ( .A(b[9]), .B(a[175]), .Z(n13603) );
  NAND U13913 ( .A(n19598), .B(n13603), .Z(n13527) );
  NAND U13914 ( .A(n13528), .B(n13527), .Z(n13606) );
  XOR U13915 ( .A(n13607), .B(n13606), .Z(n13609) );
  XOR U13916 ( .A(n13608), .B(n13609), .Z(n13619) );
  NANDN U13917 ( .A(n13530), .B(n13529), .Z(n13534) );
  OR U13918 ( .A(n13532), .B(n13531), .Z(n13533) );
  AND U13919 ( .A(n13534), .B(n13533), .Z(n13618) );
  XNOR U13920 ( .A(n13619), .B(n13618), .Z(n13620) );
  NANDN U13921 ( .A(n13536), .B(n13535), .Z(n13540) );
  NANDN U13922 ( .A(n13538), .B(n13537), .Z(n13539) );
  NAND U13923 ( .A(n13540), .B(n13539), .Z(n13621) );
  XNOR U13924 ( .A(n13620), .B(n13621), .Z(n13566) );
  XOR U13925 ( .A(n13567), .B(n13566), .Z(n13625) );
  NANDN U13926 ( .A(n13542), .B(n13541), .Z(n13546) );
  NANDN U13927 ( .A(n13544), .B(n13543), .Z(n13545) );
  AND U13928 ( .A(n13546), .B(n13545), .Z(n13624) );
  XNOR U13929 ( .A(n13625), .B(n13624), .Z(n13626) );
  XOR U13930 ( .A(n13627), .B(n13626), .Z(n13559) );
  NANDN U13931 ( .A(n13548), .B(n13547), .Z(n13552) );
  NAND U13932 ( .A(n13550), .B(n13549), .Z(n13551) );
  AND U13933 ( .A(n13552), .B(n13551), .Z(n13558) );
  XNOR U13934 ( .A(n13559), .B(n13558), .Z(n13560) );
  XNOR U13935 ( .A(n13561), .B(n13560), .Z(n13630) );
  XNOR U13936 ( .A(sreg[423]), .B(n13630), .Z(n13632) );
  NANDN U13937 ( .A(sreg[422]), .B(n13553), .Z(n13557) );
  NAND U13938 ( .A(n13555), .B(n13554), .Z(n13556) );
  NAND U13939 ( .A(n13557), .B(n13556), .Z(n13631) );
  XNOR U13940 ( .A(n13632), .B(n13631), .Z(c[423]) );
  NANDN U13941 ( .A(n13559), .B(n13558), .Z(n13563) );
  NANDN U13942 ( .A(n13561), .B(n13560), .Z(n13562) );
  AND U13943 ( .A(n13563), .B(n13562), .Z(n13638) );
  NANDN U13944 ( .A(n13565), .B(n13564), .Z(n13569) );
  NAND U13945 ( .A(n13567), .B(n13566), .Z(n13568) );
  AND U13946 ( .A(n13569), .B(n13568), .Z(n13704) );
  NANDN U13947 ( .A(n13571), .B(n13570), .Z(n13575) );
  NANDN U13948 ( .A(n13573), .B(n13572), .Z(n13574) );
  AND U13949 ( .A(n13575), .B(n13574), .Z(n13670) );
  NAND U13950 ( .A(b[0]), .B(a[184]), .Z(n13576) );
  XNOR U13951 ( .A(b[1]), .B(n13576), .Z(n13578) );
  NANDN U13952 ( .A(b[0]), .B(a[183]), .Z(n13577) );
  NAND U13953 ( .A(n13578), .B(n13577), .Z(n13650) );
  NAND U13954 ( .A(n19808), .B(n13579), .Z(n13581) );
  XOR U13955 ( .A(b[13]), .B(a[172]), .Z(n13656) );
  NAND U13956 ( .A(n19768), .B(n13656), .Z(n13580) );
  AND U13957 ( .A(n13581), .B(n13580), .Z(n13648) );
  AND U13958 ( .A(b[15]), .B(a[168]), .Z(n13647) );
  XNOR U13959 ( .A(n13648), .B(n13647), .Z(n13649) );
  XNOR U13960 ( .A(n13650), .B(n13649), .Z(n13668) );
  NAND U13961 ( .A(n33), .B(n13582), .Z(n13584) );
  XOR U13962 ( .A(b[5]), .B(a[180]), .Z(n13659) );
  NAND U13963 ( .A(n19342), .B(n13659), .Z(n13583) );
  AND U13964 ( .A(n13584), .B(n13583), .Z(n13692) );
  NAND U13965 ( .A(n34), .B(n13585), .Z(n13587) );
  XOR U13966 ( .A(b[7]), .B(a[178]), .Z(n13662) );
  NAND U13967 ( .A(n19486), .B(n13662), .Z(n13586) );
  AND U13968 ( .A(n13587), .B(n13586), .Z(n13690) );
  NAND U13969 ( .A(n31), .B(n13588), .Z(n13590) );
  XOR U13970 ( .A(b[3]), .B(a[182]), .Z(n13665) );
  NAND U13971 ( .A(n32), .B(n13665), .Z(n13589) );
  NAND U13972 ( .A(n13590), .B(n13589), .Z(n13689) );
  XNOR U13973 ( .A(n13690), .B(n13689), .Z(n13691) );
  XOR U13974 ( .A(n13692), .B(n13691), .Z(n13669) );
  XOR U13975 ( .A(n13668), .B(n13669), .Z(n13671) );
  XOR U13976 ( .A(n13670), .B(n13671), .Z(n13642) );
  NANDN U13977 ( .A(n13592), .B(n13591), .Z(n13596) );
  OR U13978 ( .A(n13594), .B(n13593), .Z(n13595) );
  AND U13979 ( .A(n13596), .B(n13595), .Z(n13641) );
  XNOR U13980 ( .A(n13642), .B(n13641), .Z(n13644) );
  NAND U13981 ( .A(n13597), .B(n19724), .Z(n13599) );
  XOR U13982 ( .A(b[11]), .B(a[174]), .Z(n13674) );
  NAND U13983 ( .A(n19692), .B(n13674), .Z(n13598) );
  AND U13984 ( .A(n13599), .B(n13598), .Z(n13685) );
  NAND U13985 ( .A(n19838), .B(n13600), .Z(n13602) );
  XOR U13986 ( .A(b[15]), .B(a[170]), .Z(n13677) );
  NAND U13987 ( .A(n19805), .B(n13677), .Z(n13601) );
  AND U13988 ( .A(n13602), .B(n13601), .Z(n13684) );
  NAND U13989 ( .A(n35), .B(n13603), .Z(n13605) );
  XOR U13990 ( .A(b[9]), .B(a[176]), .Z(n13680) );
  NAND U13991 ( .A(n19598), .B(n13680), .Z(n13604) );
  NAND U13992 ( .A(n13605), .B(n13604), .Z(n13683) );
  XOR U13993 ( .A(n13684), .B(n13683), .Z(n13686) );
  XOR U13994 ( .A(n13685), .B(n13686), .Z(n13696) );
  NANDN U13995 ( .A(n13607), .B(n13606), .Z(n13611) );
  OR U13996 ( .A(n13609), .B(n13608), .Z(n13610) );
  AND U13997 ( .A(n13611), .B(n13610), .Z(n13695) );
  XNOR U13998 ( .A(n13696), .B(n13695), .Z(n13697) );
  NANDN U13999 ( .A(n13613), .B(n13612), .Z(n13617) );
  NANDN U14000 ( .A(n13615), .B(n13614), .Z(n13616) );
  NAND U14001 ( .A(n13617), .B(n13616), .Z(n13698) );
  XNOR U14002 ( .A(n13697), .B(n13698), .Z(n13643) );
  XOR U14003 ( .A(n13644), .B(n13643), .Z(n13702) );
  NANDN U14004 ( .A(n13619), .B(n13618), .Z(n13623) );
  NANDN U14005 ( .A(n13621), .B(n13620), .Z(n13622) );
  AND U14006 ( .A(n13623), .B(n13622), .Z(n13701) );
  XNOR U14007 ( .A(n13702), .B(n13701), .Z(n13703) );
  XOR U14008 ( .A(n13704), .B(n13703), .Z(n13636) );
  NANDN U14009 ( .A(n13625), .B(n13624), .Z(n13629) );
  NAND U14010 ( .A(n13627), .B(n13626), .Z(n13628) );
  AND U14011 ( .A(n13629), .B(n13628), .Z(n13635) );
  XNOR U14012 ( .A(n13636), .B(n13635), .Z(n13637) );
  XNOR U14013 ( .A(n13638), .B(n13637), .Z(n13707) );
  XNOR U14014 ( .A(sreg[424]), .B(n13707), .Z(n13709) );
  NANDN U14015 ( .A(sreg[423]), .B(n13630), .Z(n13634) );
  NAND U14016 ( .A(n13632), .B(n13631), .Z(n13633) );
  NAND U14017 ( .A(n13634), .B(n13633), .Z(n13708) );
  XNOR U14018 ( .A(n13709), .B(n13708), .Z(c[424]) );
  NANDN U14019 ( .A(n13636), .B(n13635), .Z(n13640) );
  NANDN U14020 ( .A(n13638), .B(n13637), .Z(n13639) );
  AND U14021 ( .A(n13640), .B(n13639), .Z(n13715) );
  NANDN U14022 ( .A(n13642), .B(n13641), .Z(n13646) );
  NAND U14023 ( .A(n13644), .B(n13643), .Z(n13645) );
  AND U14024 ( .A(n13646), .B(n13645), .Z(n13781) );
  NANDN U14025 ( .A(n13648), .B(n13647), .Z(n13652) );
  NANDN U14026 ( .A(n13650), .B(n13649), .Z(n13651) );
  AND U14027 ( .A(n13652), .B(n13651), .Z(n13747) );
  NAND U14028 ( .A(b[0]), .B(a[185]), .Z(n13653) );
  XNOR U14029 ( .A(b[1]), .B(n13653), .Z(n13655) );
  NANDN U14030 ( .A(b[0]), .B(a[184]), .Z(n13654) );
  NAND U14031 ( .A(n13655), .B(n13654), .Z(n13727) );
  NAND U14032 ( .A(n19808), .B(n13656), .Z(n13658) );
  XOR U14033 ( .A(b[13]), .B(a[173]), .Z(n13733) );
  NAND U14034 ( .A(n19768), .B(n13733), .Z(n13657) );
  AND U14035 ( .A(n13658), .B(n13657), .Z(n13725) );
  AND U14036 ( .A(b[15]), .B(a[169]), .Z(n13724) );
  XNOR U14037 ( .A(n13725), .B(n13724), .Z(n13726) );
  XNOR U14038 ( .A(n13727), .B(n13726), .Z(n13745) );
  NAND U14039 ( .A(n33), .B(n13659), .Z(n13661) );
  XOR U14040 ( .A(b[5]), .B(a[181]), .Z(n13736) );
  NAND U14041 ( .A(n19342), .B(n13736), .Z(n13660) );
  AND U14042 ( .A(n13661), .B(n13660), .Z(n13769) );
  NAND U14043 ( .A(n34), .B(n13662), .Z(n13664) );
  XOR U14044 ( .A(b[7]), .B(a[179]), .Z(n13739) );
  NAND U14045 ( .A(n19486), .B(n13739), .Z(n13663) );
  AND U14046 ( .A(n13664), .B(n13663), .Z(n13767) );
  NAND U14047 ( .A(n31), .B(n13665), .Z(n13667) );
  XOR U14048 ( .A(b[3]), .B(a[183]), .Z(n13742) );
  NAND U14049 ( .A(n32), .B(n13742), .Z(n13666) );
  NAND U14050 ( .A(n13667), .B(n13666), .Z(n13766) );
  XNOR U14051 ( .A(n13767), .B(n13766), .Z(n13768) );
  XOR U14052 ( .A(n13769), .B(n13768), .Z(n13746) );
  XOR U14053 ( .A(n13745), .B(n13746), .Z(n13748) );
  XOR U14054 ( .A(n13747), .B(n13748), .Z(n13719) );
  NANDN U14055 ( .A(n13669), .B(n13668), .Z(n13673) );
  OR U14056 ( .A(n13671), .B(n13670), .Z(n13672) );
  AND U14057 ( .A(n13673), .B(n13672), .Z(n13718) );
  XNOR U14058 ( .A(n13719), .B(n13718), .Z(n13721) );
  NAND U14059 ( .A(n13674), .B(n19724), .Z(n13676) );
  XOR U14060 ( .A(b[11]), .B(a[175]), .Z(n13751) );
  NAND U14061 ( .A(n19692), .B(n13751), .Z(n13675) );
  AND U14062 ( .A(n13676), .B(n13675), .Z(n13762) );
  NAND U14063 ( .A(n19838), .B(n13677), .Z(n13679) );
  XOR U14064 ( .A(b[15]), .B(a[171]), .Z(n13754) );
  NAND U14065 ( .A(n19805), .B(n13754), .Z(n13678) );
  AND U14066 ( .A(n13679), .B(n13678), .Z(n13761) );
  NAND U14067 ( .A(n35), .B(n13680), .Z(n13682) );
  XOR U14068 ( .A(b[9]), .B(a[177]), .Z(n13757) );
  NAND U14069 ( .A(n19598), .B(n13757), .Z(n13681) );
  NAND U14070 ( .A(n13682), .B(n13681), .Z(n13760) );
  XOR U14071 ( .A(n13761), .B(n13760), .Z(n13763) );
  XOR U14072 ( .A(n13762), .B(n13763), .Z(n13773) );
  NANDN U14073 ( .A(n13684), .B(n13683), .Z(n13688) );
  OR U14074 ( .A(n13686), .B(n13685), .Z(n13687) );
  AND U14075 ( .A(n13688), .B(n13687), .Z(n13772) );
  XNOR U14076 ( .A(n13773), .B(n13772), .Z(n13774) );
  NANDN U14077 ( .A(n13690), .B(n13689), .Z(n13694) );
  NANDN U14078 ( .A(n13692), .B(n13691), .Z(n13693) );
  NAND U14079 ( .A(n13694), .B(n13693), .Z(n13775) );
  XNOR U14080 ( .A(n13774), .B(n13775), .Z(n13720) );
  XOR U14081 ( .A(n13721), .B(n13720), .Z(n13779) );
  NANDN U14082 ( .A(n13696), .B(n13695), .Z(n13700) );
  NANDN U14083 ( .A(n13698), .B(n13697), .Z(n13699) );
  AND U14084 ( .A(n13700), .B(n13699), .Z(n13778) );
  XNOR U14085 ( .A(n13779), .B(n13778), .Z(n13780) );
  XOR U14086 ( .A(n13781), .B(n13780), .Z(n13713) );
  NANDN U14087 ( .A(n13702), .B(n13701), .Z(n13706) );
  NAND U14088 ( .A(n13704), .B(n13703), .Z(n13705) );
  AND U14089 ( .A(n13706), .B(n13705), .Z(n13712) );
  XNOR U14090 ( .A(n13713), .B(n13712), .Z(n13714) );
  XNOR U14091 ( .A(n13715), .B(n13714), .Z(n13784) );
  XNOR U14092 ( .A(sreg[425]), .B(n13784), .Z(n13786) );
  NANDN U14093 ( .A(sreg[424]), .B(n13707), .Z(n13711) );
  NAND U14094 ( .A(n13709), .B(n13708), .Z(n13710) );
  NAND U14095 ( .A(n13711), .B(n13710), .Z(n13785) );
  XNOR U14096 ( .A(n13786), .B(n13785), .Z(c[425]) );
  NANDN U14097 ( .A(n13713), .B(n13712), .Z(n13717) );
  NANDN U14098 ( .A(n13715), .B(n13714), .Z(n13716) );
  AND U14099 ( .A(n13717), .B(n13716), .Z(n13792) );
  NANDN U14100 ( .A(n13719), .B(n13718), .Z(n13723) );
  NAND U14101 ( .A(n13721), .B(n13720), .Z(n13722) );
  AND U14102 ( .A(n13723), .B(n13722), .Z(n13858) );
  NANDN U14103 ( .A(n13725), .B(n13724), .Z(n13729) );
  NANDN U14104 ( .A(n13727), .B(n13726), .Z(n13728) );
  AND U14105 ( .A(n13729), .B(n13728), .Z(n13824) );
  NAND U14106 ( .A(b[0]), .B(a[186]), .Z(n13730) );
  XNOR U14107 ( .A(b[1]), .B(n13730), .Z(n13732) );
  NANDN U14108 ( .A(b[0]), .B(a[185]), .Z(n13731) );
  NAND U14109 ( .A(n13732), .B(n13731), .Z(n13804) );
  NAND U14110 ( .A(n19808), .B(n13733), .Z(n13735) );
  XOR U14111 ( .A(b[13]), .B(a[174]), .Z(n13807) );
  NAND U14112 ( .A(n19768), .B(n13807), .Z(n13734) );
  AND U14113 ( .A(n13735), .B(n13734), .Z(n13802) );
  AND U14114 ( .A(b[15]), .B(a[170]), .Z(n13801) );
  XNOR U14115 ( .A(n13802), .B(n13801), .Z(n13803) );
  XNOR U14116 ( .A(n13804), .B(n13803), .Z(n13822) );
  NAND U14117 ( .A(n33), .B(n13736), .Z(n13738) );
  XOR U14118 ( .A(b[5]), .B(a[182]), .Z(n13813) );
  NAND U14119 ( .A(n19342), .B(n13813), .Z(n13737) );
  AND U14120 ( .A(n13738), .B(n13737), .Z(n13846) );
  NAND U14121 ( .A(n34), .B(n13739), .Z(n13741) );
  XOR U14122 ( .A(b[7]), .B(a[180]), .Z(n13816) );
  NAND U14123 ( .A(n19486), .B(n13816), .Z(n13740) );
  AND U14124 ( .A(n13741), .B(n13740), .Z(n13844) );
  NAND U14125 ( .A(n31), .B(n13742), .Z(n13744) );
  XOR U14126 ( .A(b[3]), .B(a[184]), .Z(n13819) );
  NAND U14127 ( .A(n32), .B(n13819), .Z(n13743) );
  NAND U14128 ( .A(n13744), .B(n13743), .Z(n13843) );
  XNOR U14129 ( .A(n13844), .B(n13843), .Z(n13845) );
  XOR U14130 ( .A(n13846), .B(n13845), .Z(n13823) );
  XOR U14131 ( .A(n13822), .B(n13823), .Z(n13825) );
  XOR U14132 ( .A(n13824), .B(n13825), .Z(n13796) );
  NANDN U14133 ( .A(n13746), .B(n13745), .Z(n13750) );
  OR U14134 ( .A(n13748), .B(n13747), .Z(n13749) );
  AND U14135 ( .A(n13750), .B(n13749), .Z(n13795) );
  XNOR U14136 ( .A(n13796), .B(n13795), .Z(n13798) );
  NAND U14137 ( .A(n13751), .B(n19724), .Z(n13753) );
  XOR U14138 ( .A(b[11]), .B(a[176]), .Z(n13828) );
  NAND U14139 ( .A(n19692), .B(n13828), .Z(n13752) );
  AND U14140 ( .A(n13753), .B(n13752), .Z(n13839) );
  NAND U14141 ( .A(n19838), .B(n13754), .Z(n13756) );
  XOR U14142 ( .A(b[15]), .B(a[172]), .Z(n13831) );
  NAND U14143 ( .A(n19805), .B(n13831), .Z(n13755) );
  AND U14144 ( .A(n13756), .B(n13755), .Z(n13838) );
  NAND U14145 ( .A(n35), .B(n13757), .Z(n13759) );
  XOR U14146 ( .A(b[9]), .B(a[178]), .Z(n13834) );
  NAND U14147 ( .A(n19598), .B(n13834), .Z(n13758) );
  NAND U14148 ( .A(n13759), .B(n13758), .Z(n13837) );
  XOR U14149 ( .A(n13838), .B(n13837), .Z(n13840) );
  XOR U14150 ( .A(n13839), .B(n13840), .Z(n13850) );
  NANDN U14151 ( .A(n13761), .B(n13760), .Z(n13765) );
  OR U14152 ( .A(n13763), .B(n13762), .Z(n13764) );
  AND U14153 ( .A(n13765), .B(n13764), .Z(n13849) );
  XNOR U14154 ( .A(n13850), .B(n13849), .Z(n13851) );
  NANDN U14155 ( .A(n13767), .B(n13766), .Z(n13771) );
  NANDN U14156 ( .A(n13769), .B(n13768), .Z(n13770) );
  NAND U14157 ( .A(n13771), .B(n13770), .Z(n13852) );
  XNOR U14158 ( .A(n13851), .B(n13852), .Z(n13797) );
  XOR U14159 ( .A(n13798), .B(n13797), .Z(n13856) );
  NANDN U14160 ( .A(n13773), .B(n13772), .Z(n13777) );
  NANDN U14161 ( .A(n13775), .B(n13774), .Z(n13776) );
  AND U14162 ( .A(n13777), .B(n13776), .Z(n13855) );
  XNOR U14163 ( .A(n13856), .B(n13855), .Z(n13857) );
  XOR U14164 ( .A(n13858), .B(n13857), .Z(n13790) );
  NANDN U14165 ( .A(n13779), .B(n13778), .Z(n13783) );
  NAND U14166 ( .A(n13781), .B(n13780), .Z(n13782) );
  AND U14167 ( .A(n13783), .B(n13782), .Z(n13789) );
  XNOR U14168 ( .A(n13790), .B(n13789), .Z(n13791) );
  XNOR U14169 ( .A(n13792), .B(n13791), .Z(n13861) );
  XNOR U14170 ( .A(sreg[426]), .B(n13861), .Z(n13863) );
  NANDN U14171 ( .A(sreg[425]), .B(n13784), .Z(n13788) );
  NAND U14172 ( .A(n13786), .B(n13785), .Z(n13787) );
  NAND U14173 ( .A(n13788), .B(n13787), .Z(n13862) );
  XNOR U14174 ( .A(n13863), .B(n13862), .Z(c[426]) );
  NANDN U14175 ( .A(n13790), .B(n13789), .Z(n13794) );
  NANDN U14176 ( .A(n13792), .B(n13791), .Z(n13793) );
  AND U14177 ( .A(n13794), .B(n13793), .Z(n13869) );
  NANDN U14178 ( .A(n13796), .B(n13795), .Z(n13800) );
  NAND U14179 ( .A(n13798), .B(n13797), .Z(n13799) );
  AND U14180 ( .A(n13800), .B(n13799), .Z(n13935) );
  NANDN U14181 ( .A(n13802), .B(n13801), .Z(n13806) );
  NANDN U14182 ( .A(n13804), .B(n13803), .Z(n13805) );
  AND U14183 ( .A(n13806), .B(n13805), .Z(n13901) );
  NAND U14184 ( .A(n19808), .B(n13807), .Z(n13809) );
  XOR U14185 ( .A(b[13]), .B(a[175]), .Z(n13887) );
  NAND U14186 ( .A(n19768), .B(n13887), .Z(n13808) );
  AND U14187 ( .A(n13809), .B(n13808), .Z(n13879) );
  AND U14188 ( .A(b[15]), .B(a[171]), .Z(n13878) );
  XNOR U14189 ( .A(n13879), .B(n13878), .Z(n13880) );
  NAND U14190 ( .A(b[0]), .B(a[187]), .Z(n13810) );
  XNOR U14191 ( .A(b[1]), .B(n13810), .Z(n13812) );
  NANDN U14192 ( .A(b[0]), .B(a[186]), .Z(n13811) );
  NAND U14193 ( .A(n13812), .B(n13811), .Z(n13881) );
  XNOR U14194 ( .A(n13880), .B(n13881), .Z(n13899) );
  NAND U14195 ( .A(n33), .B(n13813), .Z(n13815) );
  XOR U14196 ( .A(b[5]), .B(a[183]), .Z(n13890) );
  NAND U14197 ( .A(n19342), .B(n13890), .Z(n13814) );
  AND U14198 ( .A(n13815), .B(n13814), .Z(n13923) );
  NAND U14199 ( .A(n34), .B(n13816), .Z(n13818) );
  XOR U14200 ( .A(b[7]), .B(a[181]), .Z(n13893) );
  NAND U14201 ( .A(n19486), .B(n13893), .Z(n13817) );
  AND U14202 ( .A(n13818), .B(n13817), .Z(n13921) );
  NAND U14203 ( .A(n31), .B(n13819), .Z(n13821) );
  XOR U14204 ( .A(b[3]), .B(a[185]), .Z(n13896) );
  NAND U14205 ( .A(n32), .B(n13896), .Z(n13820) );
  NAND U14206 ( .A(n13821), .B(n13820), .Z(n13920) );
  XNOR U14207 ( .A(n13921), .B(n13920), .Z(n13922) );
  XOR U14208 ( .A(n13923), .B(n13922), .Z(n13900) );
  XOR U14209 ( .A(n13899), .B(n13900), .Z(n13902) );
  XOR U14210 ( .A(n13901), .B(n13902), .Z(n13873) );
  NANDN U14211 ( .A(n13823), .B(n13822), .Z(n13827) );
  OR U14212 ( .A(n13825), .B(n13824), .Z(n13826) );
  AND U14213 ( .A(n13827), .B(n13826), .Z(n13872) );
  XNOR U14214 ( .A(n13873), .B(n13872), .Z(n13875) );
  NAND U14215 ( .A(n13828), .B(n19724), .Z(n13830) );
  XOR U14216 ( .A(b[11]), .B(a[177]), .Z(n13905) );
  NAND U14217 ( .A(n19692), .B(n13905), .Z(n13829) );
  AND U14218 ( .A(n13830), .B(n13829), .Z(n13916) );
  NAND U14219 ( .A(n19838), .B(n13831), .Z(n13833) );
  XOR U14220 ( .A(b[15]), .B(a[173]), .Z(n13908) );
  NAND U14221 ( .A(n19805), .B(n13908), .Z(n13832) );
  AND U14222 ( .A(n13833), .B(n13832), .Z(n13915) );
  NAND U14223 ( .A(n35), .B(n13834), .Z(n13836) );
  XOR U14224 ( .A(b[9]), .B(a[179]), .Z(n13911) );
  NAND U14225 ( .A(n19598), .B(n13911), .Z(n13835) );
  NAND U14226 ( .A(n13836), .B(n13835), .Z(n13914) );
  XOR U14227 ( .A(n13915), .B(n13914), .Z(n13917) );
  XOR U14228 ( .A(n13916), .B(n13917), .Z(n13927) );
  NANDN U14229 ( .A(n13838), .B(n13837), .Z(n13842) );
  OR U14230 ( .A(n13840), .B(n13839), .Z(n13841) );
  AND U14231 ( .A(n13842), .B(n13841), .Z(n13926) );
  XNOR U14232 ( .A(n13927), .B(n13926), .Z(n13928) );
  NANDN U14233 ( .A(n13844), .B(n13843), .Z(n13848) );
  NANDN U14234 ( .A(n13846), .B(n13845), .Z(n13847) );
  NAND U14235 ( .A(n13848), .B(n13847), .Z(n13929) );
  XNOR U14236 ( .A(n13928), .B(n13929), .Z(n13874) );
  XOR U14237 ( .A(n13875), .B(n13874), .Z(n13933) );
  NANDN U14238 ( .A(n13850), .B(n13849), .Z(n13854) );
  NANDN U14239 ( .A(n13852), .B(n13851), .Z(n13853) );
  AND U14240 ( .A(n13854), .B(n13853), .Z(n13932) );
  XNOR U14241 ( .A(n13933), .B(n13932), .Z(n13934) );
  XOR U14242 ( .A(n13935), .B(n13934), .Z(n13867) );
  NANDN U14243 ( .A(n13856), .B(n13855), .Z(n13860) );
  NAND U14244 ( .A(n13858), .B(n13857), .Z(n13859) );
  AND U14245 ( .A(n13860), .B(n13859), .Z(n13866) );
  XNOR U14246 ( .A(n13867), .B(n13866), .Z(n13868) );
  XNOR U14247 ( .A(n13869), .B(n13868), .Z(n13938) );
  XNOR U14248 ( .A(sreg[427]), .B(n13938), .Z(n13940) );
  NANDN U14249 ( .A(sreg[426]), .B(n13861), .Z(n13865) );
  NAND U14250 ( .A(n13863), .B(n13862), .Z(n13864) );
  NAND U14251 ( .A(n13865), .B(n13864), .Z(n13939) );
  XNOR U14252 ( .A(n13940), .B(n13939), .Z(c[427]) );
  NANDN U14253 ( .A(n13867), .B(n13866), .Z(n13871) );
  NANDN U14254 ( .A(n13869), .B(n13868), .Z(n13870) );
  AND U14255 ( .A(n13871), .B(n13870), .Z(n13946) );
  NANDN U14256 ( .A(n13873), .B(n13872), .Z(n13877) );
  NAND U14257 ( .A(n13875), .B(n13874), .Z(n13876) );
  AND U14258 ( .A(n13877), .B(n13876), .Z(n14012) );
  NANDN U14259 ( .A(n13879), .B(n13878), .Z(n13883) );
  NANDN U14260 ( .A(n13881), .B(n13880), .Z(n13882) );
  AND U14261 ( .A(n13883), .B(n13882), .Z(n13978) );
  NAND U14262 ( .A(b[0]), .B(a[188]), .Z(n13884) );
  XNOR U14263 ( .A(b[1]), .B(n13884), .Z(n13886) );
  NANDN U14264 ( .A(b[0]), .B(a[187]), .Z(n13885) );
  NAND U14265 ( .A(n13886), .B(n13885), .Z(n13958) );
  NAND U14266 ( .A(n19808), .B(n13887), .Z(n13889) );
  XOR U14267 ( .A(b[13]), .B(a[176]), .Z(n13961) );
  NAND U14268 ( .A(n19768), .B(n13961), .Z(n13888) );
  AND U14269 ( .A(n13889), .B(n13888), .Z(n13956) );
  AND U14270 ( .A(b[15]), .B(a[172]), .Z(n13955) );
  XNOR U14271 ( .A(n13956), .B(n13955), .Z(n13957) );
  XNOR U14272 ( .A(n13958), .B(n13957), .Z(n13976) );
  NAND U14273 ( .A(n33), .B(n13890), .Z(n13892) );
  XOR U14274 ( .A(b[5]), .B(a[184]), .Z(n13967) );
  NAND U14275 ( .A(n19342), .B(n13967), .Z(n13891) );
  AND U14276 ( .A(n13892), .B(n13891), .Z(n14000) );
  NAND U14277 ( .A(n34), .B(n13893), .Z(n13895) );
  XOR U14278 ( .A(b[7]), .B(a[182]), .Z(n13970) );
  NAND U14279 ( .A(n19486), .B(n13970), .Z(n13894) );
  AND U14280 ( .A(n13895), .B(n13894), .Z(n13998) );
  NAND U14281 ( .A(n31), .B(n13896), .Z(n13898) );
  XOR U14282 ( .A(b[3]), .B(a[186]), .Z(n13973) );
  NAND U14283 ( .A(n32), .B(n13973), .Z(n13897) );
  NAND U14284 ( .A(n13898), .B(n13897), .Z(n13997) );
  XNOR U14285 ( .A(n13998), .B(n13997), .Z(n13999) );
  XOR U14286 ( .A(n14000), .B(n13999), .Z(n13977) );
  XOR U14287 ( .A(n13976), .B(n13977), .Z(n13979) );
  XOR U14288 ( .A(n13978), .B(n13979), .Z(n13950) );
  NANDN U14289 ( .A(n13900), .B(n13899), .Z(n13904) );
  OR U14290 ( .A(n13902), .B(n13901), .Z(n13903) );
  AND U14291 ( .A(n13904), .B(n13903), .Z(n13949) );
  XNOR U14292 ( .A(n13950), .B(n13949), .Z(n13952) );
  NAND U14293 ( .A(n13905), .B(n19724), .Z(n13907) );
  XOR U14294 ( .A(b[11]), .B(a[178]), .Z(n13982) );
  NAND U14295 ( .A(n19692), .B(n13982), .Z(n13906) );
  AND U14296 ( .A(n13907), .B(n13906), .Z(n13993) );
  NAND U14297 ( .A(n19838), .B(n13908), .Z(n13910) );
  XOR U14298 ( .A(b[15]), .B(a[174]), .Z(n13985) );
  NAND U14299 ( .A(n19805), .B(n13985), .Z(n13909) );
  AND U14300 ( .A(n13910), .B(n13909), .Z(n13992) );
  NAND U14301 ( .A(n35), .B(n13911), .Z(n13913) );
  XOR U14302 ( .A(b[9]), .B(a[180]), .Z(n13988) );
  NAND U14303 ( .A(n19598), .B(n13988), .Z(n13912) );
  NAND U14304 ( .A(n13913), .B(n13912), .Z(n13991) );
  XOR U14305 ( .A(n13992), .B(n13991), .Z(n13994) );
  XOR U14306 ( .A(n13993), .B(n13994), .Z(n14004) );
  NANDN U14307 ( .A(n13915), .B(n13914), .Z(n13919) );
  OR U14308 ( .A(n13917), .B(n13916), .Z(n13918) );
  AND U14309 ( .A(n13919), .B(n13918), .Z(n14003) );
  XNOR U14310 ( .A(n14004), .B(n14003), .Z(n14005) );
  NANDN U14311 ( .A(n13921), .B(n13920), .Z(n13925) );
  NANDN U14312 ( .A(n13923), .B(n13922), .Z(n13924) );
  NAND U14313 ( .A(n13925), .B(n13924), .Z(n14006) );
  XNOR U14314 ( .A(n14005), .B(n14006), .Z(n13951) );
  XOR U14315 ( .A(n13952), .B(n13951), .Z(n14010) );
  NANDN U14316 ( .A(n13927), .B(n13926), .Z(n13931) );
  NANDN U14317 ( .A(n13929), .B(n13928), .Z(n13930) );
  AND U14318 ( .A(n13931), .B(n13930), .Z(n14009) );
  XNOR U14319 ( .A(n14010), .B(n14009), .Z(n14011) );
  XOR U14320 ( .A(n14012), .B(n14011), .Z(n13944) );
  NANDN U14321 ( .A(n13933), .B(n13932), .Z(n13937) );
  NAND U14322 ( .A(n13935), .B(n13934), .Z(n13936) );
  AND U14323 ( .A(n13937), .B(n13936), .Z(n13943) );
  XNOR U14324 ( .A(n13944), .B(n13943), .Z(n13945) );
  XNOR U14325 ( .A(n13946), .B(n13945), .Z(n14015) );
  XNOR U14326 ( .A(sreg[428]), .B(n14015), .Z(n14017) );
  NANDN U14327 ( .A(sreg[427]), .B(n13938), .Z(n13942) );
  NAND U14328 ( .A(n13940), .B(n13939), .Z(n13941) );
  NAND U14329 ( .A(n13942), .B(n13941), .Z(n14016) );
  XNOR U14330 ( .A(n14017), .B(n14016), .Z(c[428]) );
  NANDN U14331 ( .A(n13944), .B(n13943), .Z(n13948) );
  NANDN U14332 ( .A(n13946), .B(n13945), .Z(n13947) );
  AND U14333 ( .A(n13948), .B(n13947), .Z(n14023) );
  NANDN U14334 ( .A(n13950), .B(n13949), .Z(n13954) );
  NAND U14335 ( .A(n13952), .B(n13951), .Z(n13953) );
  AND U14336 ( .A(n13954), .B(n13953), .Z(n14089) );
  NANDN U14337 ( .A(n13956), .B(n13955), .Z(n13960) );
  NANDN U14338 ( .A(n13958), .B(n13957), .Z(n13959) );
  AND U14339 ( .A(n13960), .B(n13959), .Z(n14055) );
  NAND U14340 ( .A(n19808), .B(n13961), .Z(n13963) );
  XOR U14341 ( .A(b[13]), .B(a[177]), .Z(n14041) );
  NAND U14342 ( .A(n19768), .B(n14041), .Z(n13962) );
  AND U14343 ( .A(n13963), .B(n13962), .Z(n14033) );
  AND U14344 ( .A(b[15]), .B(a[173]), .Z(n14032) );
  XNOR U14345 ( .A(n14033), .B(n14032), .Z(n14034) );
  NAND U14346 ( .A(b[0]), .B(a[189]), .Z(n13964) );
  XNOR U14347 ( .A(b[1]), .B(n13964), .Z(n13966) );
  NANDN U14348 ( .A(b[0]), .B(a[188]), .Z(n13965) );
  NAND U14349 ( .A(n13966), .B(n13965), .Z(n14035) );
  XNOR U14350 ( .A(n14034), .B(n14035), .Z(n14053) );
  NAND U14351 ( .A(n33), .B(n13967), .Z(n13969) );
  XOR U14352 ( .A(b[5]), .B(a[185]), .Z(n14044) );
  NAND U14353 ( .A(n19342), .B(n14044), .Z(n13968) );
  AND U14354 ( .A(n13969), .B(n13968), .Z(n14077) );
  NAND U14355 ( .A(n34), .B(n13970), .Z(n13972) );
  XOR U14356 ( .A(b[7]), .B(a[183]), .Z(n14047) );
  NAND U14357 ( .A(n19486), .B(n14047), .Z(n13971) );
  AND U14358 ( .A(n13972), .B(n13971), .Z(n14075) );
  NAND U14359 ( .A(n31), .B(n13973), .Z(n13975) );
  XOR U14360 ( .A(b[3]), .B(a[187]), .Z(n14050) );
  NAND U14361 ( .A(n32), .B(n14050), .Z(n13974) );
  NAND U14362 ( .A(n13975), .B(n13974), .Z(n14074) );
  XNOR U14363 ( .A(n14075), .B(n14074), .Z(n14076) );
  XOR U14364 ( .A(n14077), .B(n14076), .Z(n14054) );
  XOR U14365 ( .A(n14053), .B(n14054), .Z(n14056) );
  XOR U14366 ( .A(n14055), .B(n14056), .Z(n14027) );
  NANDN U14367 ( .A(n13977), .B(n13976), .Z(n13981) );
  OR U14368 ( .A(n13979), .B(n13978), .Z(n13980) );
  AND U14369 ( .A(n13981), .B(n13980), .Z(n14026) );
  XNOR U14370 ( .A(n14027), .B(n14026), .Z(n14029) );
  NAND U14371 ( .A(n13982), .B(n19724), .Z(n13984) );
  XOR U14372 ( .A(b[11]), .B(a[179]), .Z(n14059) );
  NAND U14373 ( .A(n19692), .B(n14059), .Z(n13983) );
  AND U14374 ( .A(n13984), .B(n13983), .Z(n14070) );
  NAND U14375 ( .A(n19838), .B(n13985), .Z(n13987) );
  XOR U14376 ( .A(b[15]), .B(a[175]), .Z(n14062) );
  NAND U14377 ( .A(n19805), .B(n14062), .Z(n13986) );
  AND U14378 ( .A(n13987), .B(n13986), .Z(n14069) );
  NAND U14379 ( .A(n35), .B(n13988), .Z(n13990) );
  XOR U14380 ( .A(b[9]), .B(a[181]), .Z(n14065) );
  NAND U14381 ( .A(n19598), .B(n14065), .Z(n13989) );
  NAND U14382 ( .A(n13990), .B(n13989), .Z(n14068) );
  XOR U14383 ( .A(n14069), .B(n14068), .Z(n14071) );
  XOR U14384 ( .A(n14070), .B(n14071), .Z(n14081) );
  NANDN U14385 ( .A(n13992), .B(n13991), .Z(n13996) );
  OR U14386 ( .A(n13994), .B(n13993), .Z(n13995) );
  AND U14387 ( .A(n13996), .B(n13995), .Z(n14080) );
  XNOR U14388 ( .A(n14081), .B(n14080), .Z(n14082) );
  NANDN U14389 ( .A(n13998), .B(n13997), .Z(n14002) );
  NANDN U14390 ( .A(n14000), .B(n13999), .Z(n14001) );
  NAND U14391 ( .A(n14002), .B(n14001), .Z(n14083) );
  XNOR U14392 ( .A(n14082), .B(n14083), .Z(n14028) );
  XOR U14393 ( .A(n14029), .B(n14028), .Z(n14087) );
  NANDN U14394 ( .A(n14004), .B(n14003), .Z(n14008) );
  NANDN U14395 ( .A(n14006), .B(n14005), .Z(n14007) );
  AND U14396 ( .A(n14008), .B(n14007), .Z(n14086) );
  XNOR U14397 ( .A(n14087), .B(n14086), .Z(n14088) );
  XOR U14398 ( .A(n14089), .B(n14088), .Z(n14021) );
  NANDN U14399 ( .A(n14010), .B(n14009), .Z(n14014) );
  NAND U14400 ( .A(n14012), .B(n14011), .Z(n14013) );
  AND U14401 ( .A(n14014), .B(n14013), .Z(n14020) );
  XNOR U14402 ( .A(n14021), .B(n14020), .Z(n14022) );
  XNOR U14403 ( .A(n14023), .B(n14022), .Z(n14092) );
  XNOR U14404 ( .A(sreg[429]), .B(n14092), .Z(n14094) );
  NANDN U14405 ( .A(sreg[428]), .B(n14015), .Z(n14019) );
  NAND U14406 ( .A(n14017), .B(n14016), .Z(n14018) );
  NAND U14407 ( .A(n14019), .B(n14018), .Z(n14093) );
  XNOR U14408 ( .A(n14094), .B(n14093), .Z(c[429]) );
  NANDN U14409 ( .A(n14021), .B(n14020), .Z(n14025) );
  NANDN U14410 ( .A(n14023), .B(n14022), .Z(n14024) );
  AND U14411 ( .A(n14025), .B(n14024), .Z(n14100) );
  NANDN U14412 ( .A(n14027), .B(n14026), .Z(n14031) );
  NAND U14413 ( .A(n14029), .B(n14028), .Z(n14030) );
  AND U14414 ( .A(n14031), .B(n14030), .Z(n14166) );
  NANDN U14415 ( .A(n14033), .B(n14032), .Z(n14037) );
  NANDN U14416 ( .A(n14035), .B(n14034), .Z(n14036) );
  AND U14417 ( .A(n14037), .B(n14036), .Z(n14132) );
  NAND U14418 ( .A(b[0]), .B(a[190]), .Z(n14038) );
  XNOR U14419 ( .A(b[1]), .B(n14038), .Z(n14040) );
  NANDN U14420 ( .A(b[0]), .B(a[189]), .Z(n14039) );
  NAND U14421 ( .A(n14040), .B(n14039), .Z(n14112) );
  NAND U14422 ( .A(n19808), .B(n14041), .Z(n14043) );
  XOR U14423 ( .A(b[13]), .B(a[178]), .Z(n14118) );
  NAND U14424 ( .A(n19768), .B(n14118), .Z(n14042) );
  AND U14425 ( .A(n14043), .B(n14042), .Z(n14110) );
  AND U14426 ( .A(b[15]), .B(a[174]), .Z(n14109) );
  XNOR U14427 ( .A(n14110), .B(n14109), .Z(n14111) );
  XNOR U14428 ( .A(n14112), .B(n14111), .Z(n14130) );
  NAND U14429 ( .A(n33), .B(n14044), .Z(n14046) );
  XOR U14430 ( .A(b[5]), .B(a[186]), .Z(n14121) );
  NAND U14431 ( .A(n19342), .B(n14121), .Z(n14045) );
  AND U14432 ( .A(n14046), .B(n14045), .Z(n14154) );
  NAND U14433 ( .A(n34), .B(n14047), .Z(n14049) );
  XOR U14434 ( .A(b[7]), .B(a[184]), .Z(n14124) );
  NAND U14435 ( .A(n19486), .B(n14124), .Z(n14048) );
  AND U14436 ( .A(n14049), .B(n14048), .Z(n14152) );
  NAND U14437 ( .A(n31), .B(n14050), .Z(n14052) );
  XOR U14438 ( .A(b[3]), .B(a[188]), .Z(n14127) );
  NAND U14439 ( .A(n32), .B(n14127), .Z(n14051) );
  NAND U14440 ( .A(n14052), .B(n14051), .Z(n14151) );
  XNOR U14441 ( .A(n14152), .B(n14151), .Z(n14153) );
  XOR U14442 ( .A(n14154), .B(n14153), .Z(n14131) );
  XOR U14443 ( .A(n14130), .B(n14131), .Z(n14133) );
  XOR U14444 ( .A(n14132), .B(n14133), .Z(n14104) );
  NANDN U14445 ( .A(n14054), .B(n14053), .Z(n14058) );
  OR U14446 ( .A(n14056), .B(n14055), .Z(n14057) );
  AND U14447 ( .A(n14058), .B(n14057), .Z(n14103) );
  XNOR U14448 ( .A(n14104), .B(n14103), .Z(n14106) );
  NAND U14449 ( .A(n14059), .B(n19724), .Z(n14061) );
  XOR U14450 ( .A(b[11]), .B(a[180]), .Z(n14136) );
  NAND U14451 ( .A(n19692), .B(n14136), .Z(n14060) );
  AND U14452 ( .A(n14061), .B(n14060), .Z(n14147) );
  NAND U14453 ( .A(n19838), .B(n14062), .Z(n14064) );
  XOR U14454 ( .A(b[15]), .B(a[176]), .Z(n14139) );
  NAND U14455 ( .A(n19805), .B(n14139), .Z(n14063) );
  AND U14456 ( .A(n14064), .B(n14063), .Z(n14146) );
  NAND U14457 ( .A(n35), .B(n14065), .Z(n14067) );
  XOR U14458 ( .A(b[9]), .B(a[182]), .Z(n14142) );
  NAND U14459 ( .A(n19598), .B(n14142), .Z(n14066) );
  NAND U14460 ( .A(n14067), .B(n14066), .Z(n14145) );
  XOR U14461 ( .A(n14146), .B(n14145), .Z(n14148) );
  XOR U14462 ( .A(n14147), .B(n14148), .Z(n14158) );
  NANDN U14463 ( .A(n14069), .B(n14068), .Z(n14073) );
  OR U14464 ( .A(n14071), .B(n14070), .Z(n14072) );
  AND U14465 ( .A(n14073), .B(n14072), .Z(n14157) );
  XNOR U14466 ( .A(n14158), .B(n14157), .Z(n14159) );
  NANDN U14467 ( .A(n14075), .B(n14074), .Z(n14079) );
  NANDN U14468 ( .A(n14077), .B(n14076), .Z(n14078) );
  NAND U14469 ( .A(n14079), .B(n14078), .Z(n14160) );
  XNOR U14470 ( .A(n14159), .B(n14160), .Z(n14105) );
  XOR U14471 ( .A(n14106), .B(n14105), .Z(n14164) );
  NANDN U14472 ( .A(n14081), .B(n14080), .Z(n14085) );
  NANDN U14473 ( .A(n14083), .B(n14082), .Z(n14084) );
  AND U14474 ( .A(n14085), .B(n14084), .Z(n14163) );
  XNOR U14475 ( .A(n14164), .B(n14163), .Z(n14165) );
  XOR U14476 ( .A(n14166), .B(n14165), .Z(n14098) );
  NANDN U14477 ( .A(n14087), .B(n14086), .Z(n14091) );
  NAND U14478 ( .A(n14089), .B(n14088), .Z(n14090) );
  AND U14479 ( .A(n14091), .B(n14090), .Z(n14097) );
  XNOR U14480 ( .A(n14098), .B(n14097), .Z(n14099) );
  XNOR U14481 ( .A(n14100), .B(n14099), .Z(n14169) );
  XNOR U14482 ( .A(sreg[430]), .B(n14169), .Z(n14171) );
  NANDN U14483 ( .A(sreg[429]), .B(n14092), .Z(n14096) );
  NAND U14484 ( .A(n14094), .B(n14093), .Z(n14095) );
  NAND U14485 ( .A(n14096), .B(n14095), .Z(n14170) );
  XNOR U14486 ( .A(n14171), .B(n14170), .Z(c[430]) );
  NANDN U14487 ( .A(n14098), .B(n14097), .Z(n14102) );
  NANDN U14488 ( .A(n14100), .B(n14099), .Z(n14101) );
  AND U14489 ( .A(n14102), .B(n14101), .Z(n14177) );
  NANDN U14490 ( .A(n14104), .B(n14103), .Z(n14108) );
  NAND U14491 ( .A(n14106), .B(n14105), .Z(n14107) );
  AND U14492 ( .A(n14108), .B(n14107), .Z(n14243) );
  NANDN U14493 ( .A(n14110), .B(n14109), .Z(n14114) );
  NANDN U14494 ( .A(n14112), .B(n14111), .Z(n14113) );
  AND U14495 ( .A(n14114), .B(n14113), .Z(n14209) );
  NAND U14496 ( .A(b[0]), .B(a[191]), .Z(n14115) );
  XNOR U14497 ( .A(b[1]), .B(n14115), .Z(n14117) );
  NANDN U14498 ( .A(b[0]), .B(a[190]), .Z(n14116) );
  NAND U14499 ( .A(n14117), .B(n14116), .Z(n14189) );
  NAND U14500 ( .A(n19808), .B(n14118), .Z(n14120) );
  XOR U14501 ( .A(b[13]), .B(a[179]), .Z(n14192) );
  NAND U14502 ( .A(n19768), .B(n14192), .Z(n14119) );
  AND U14503 ( .A(n14120), .B(n14119), .Z(n14187) );
  AND U14504 ( .A(b[15]), .B(a[175]), .Z(n14186) );
  XNOR U14505 ( .A(n14187), .B(n14186), .Z(n14188) );
  XNOR U14506 ( .A(n14189), .B(n14188), .Z(n14207) );
  NAND U14507 ( .A(n33), .B(n14121), .Z(n14123) );
  XOR U14508 ( .A(b[5]), .B(a[187]), .Z(n14198) );
  NAND U14509 ( .A(n19342), .B(n14198), .Z(n14122) );
  AND U14510 ( .A(n14123), .B(n14122), .Z(n14231) );
  NAND U14511 ( .A(n34), .B(n14124), .Z(n14126) );
  XOR U14512 ( .A(b[7]), .B(a[185]), .Z(n14201) );
  NAND U14513 ( .A(n19486), .B(n14201), .Z(n14125) );
  AND U14514 ( .A(n14126), .B(n14125), .Z(n14229) );
  NAND U14515 ( .A(n31), .B(n14127), .Z(n14129) );
  XOR U14516 ( .A(b[3]), .B(a[189]), .Z(n14204) );
  NAND U14517 ( .A(n32), .B(n14204), .Z(n14128) );
  NAND U14518 ( .A(n14129), .B(n14128), .Z(n14228) );
  XNOR U14519 ( .A(n14229), .B(n14228), .Z(n14230) );
  XOR U14520 ( .A(n14231), .B(n14230), .Z(n14208) );
  XOR U14521 ( .A(n14207), .B(n14208), .Z(n14210) );
  XOR U14522 ( .A(n14209), .B(n14210), .Z(n14181) );
  NANDN U14523 ( .A(n14131), .B(n14130), .Z(n14135) );
  OR U14524 ( .A(n14133), .B(n14132), .Z(n14134) );
  AND U14525 ( .A(n14135), .B(n14134), .Z(n14180) );
  XNOR U14526 ( .A(n14181), .B(n14180), .Z(n14183) );
  NAND U14527 ( .A(n14136), .B(n19724), .Z(n14138) );
  XOR U14528 ( .A(b[11]), .B(a[181]), .Z(n14213) );
  NAND U14529 ( .A(n19692), .B(n14213), .Z(n14137) );
  AND U14530 ( .A(n14138), .B(n14137), .Z(n14224) );
  NAND U14531 ( .A(n19838), .B(n14139), .Z(n14141) );
  XOR U14532 ( .A(b[15]), .B(a[177]), .Z(n14216) );
  NAND U14533 ( .A(n19805), .B(n14216), .Z(n14140) );
  AND U14534 ( .A(n14141), .B(n14140), .Z(n14223) );
  NAND U14535 ( .A(n35), .B(n14142), .Z(n14144) );
  XOR U14536 ( .A(b[9]), .B(a[183]), .Z(n14219) );
  NAND U14537 ( .A(n19598), .B(n14219), .Z(n14143) );
  NAND U14538 ( .A(n14144), .B(n14143), .Z(n14222) );
  XOR U14539 ( .A(n14223), .B(n14222), .Z(n14225) );
  XOR U14540 ( .A(n14224), .B(n14225), .Z(n14235) );
  NANDN U14541 ( .A(n14146), .B(n14145), .Z(n14150) );
  OR U14542 ( .A(n14148), .B(n14147), .Z(n14149) );
  AND U14543 ( .A(n14150), .B(n14149), .Z(n14234) );
  XNOR U14544 ( .A(n14235), .B(n14234), .Z(n14236) );
  NANDN U14545 ( .A(n14152), .B(n14151), .Z(n14156) );
  NANDN U14546 ( .A(n14154), .B(n14153), .Z(n14155) );
  NAND U14547 ( .A(n14156), .B(n14155), .Z(n14237) );
  XNOR U14548 ( .A(n14236), .B(n14237), .Z(n14182) );
  XOR U14549 ( .A(n14183), .B(n14182), .Z(n14241) );
  NANDN U14550 ( .A(n14158), .B(n14157), .Z(n14162) );
  NANDN U14551 ( .A(n14160), .B(n14159), .Z(n14161) );
  AND U14552 ( .A(n14162), .B(n14161), .Z(n14240) );
  XNOR U14553 ( .A(n14241), .B(n14240), .Z(n14242) );
  XOR U14554 ( .A(n14243), .B(n14242), .Z(n14175) );
  NANDN U14555 ( .A(n14164), .B(n14163), .Z(n14168) );
  NAND U14556 ( .A(n14166), .B(n14165), .Z(n14167) );
  AND U14557 ( .A(n14168), .B(n14167), .Z(n14174) );
  XNOR U14558 ( .A(n14175), .B(n14174), .Z(n14176) );
  XNOR U14559 ( .A(n14177), .B(n14176), .Z(n14246) );
  XNOR U14560 ( .A(sreg[431]), .B(n14246), .Z(n14248) );
  NANDN U14561 ( .A(sreg[430]), .B(n14169), .Z(n14173) );
  NAND U14562 ( .A(n14171), .B(n14170), .Z(n14172) );
  NAND U14563 ( .A(n14173), .B(n14172), .Z(n14247) );
  XNOR U14564 ( .A(n14248), .B(n14247), .Z(c[431]) );
  NANDN U14565 ( .A(n14175), .B(n14174), .Z(n14179) );
  NANDN U14566 ( .A(n14177), .B(n14176), .Z(n14178) );
  AND U14567 ( .A(n14179), .B(n14178), .Z(n14254) );
  NANDN U14568 ( .A(n14181), .B(n14180), .Z(n14185) );
  NAND U14569 ( .A(n14183), .B(n14182), .Z(n14184) );
  AND U14570 ( .A(n14185), .B(n14184), .Z(n14320) );
  NANDN U14571 ( .A(n14187), .B(n14186), .Z(n14191) );
  NANDN U14572 ( .A(n14189), .B(n14188), .Z(n14190) );
  AND U14573 ( .A(n14191), .B(n14190), .Z(n14286) );
  NAND U14574 ( .A(n19808), .B(n14192), .Z(n14194) );
  XOR U14575 ( .A(b[13]), .B(a[180]), .Z(n14272) );
  NAND U14576 ( .A(n19768), .B(n14272), .Z(n14193) );
  AND U14577 ( .A(n14194), .B(n14193), .Z(n14264) );
  AND U14578 ( .A(b[15]), .B(a[176]), .Z(n14263) );
  XNOR U14579 ( .A(n14264), .B(n14263), .Z(n14265) );
  NAND U14580 ( .A(b[0]), .B(a[192]), .Z(n14195) );
  XNOR U14581 ( .A(b[1]), .B(n14195), .Z(n14197) );
  NANDN U14582 ( .A(b[0]), .B(a[191]), .Z(n14196) );
  NAND U14583 ( .A(n14197), .B(n14196), .Z(n14266) );
  XNOR U14584 ( .A(n14265), .B(n14266), .Z(n14284) );
  NAND U14585 ( .A(n33), .B(n14198), .Z(n14200) );
  XOR U14586 ( .A(b[5]), .B(a[188]), .Z(n14275) );
  NAND U14587 ( .A(n19342), .B(n14275), .Z(n14199) );
  AND U14588 ( .A(n14200), .B(n14199), .Z(n14308) );
  NAND U14589 ( .A(n34), .B(n14201), .Z(n14203) );
  XOR U14590 ( .A(b[7]), .B(a[186]), .Z(n14278) );
  NAND U14591 ( .A(n19486), .B(n14278), .Z(n14202) );
  AND U14592 ( .A(n14203), .B(n14202), .Z(n14306) );
  NAND U14593 ( .A(n31), .B(n14204), .Z(n14206) );
  XOR U14594 ( .A(b[3]), .B(a[190]), .Z(n14281) );
  NAND U14595 ( .A(n32), .B(n14281), .Z(n14205) );
  NAND U14596 ( .A(n14206), .B(n14205), .Z(n14305) );
  XNOR U14597 ( .A(n14306), .B(n14305), .Z(n14307) );
  XOR U14598 ( .A(n14308), .B(n14307), .Z(n14285) );
  XOR U14599 ( .A(n14284), .B(n14285), .Z(n14287) );
  XOR U14600 ( .A(n14286), .B(n14287), .Z(n14258) );
  NANDN U14601 ( .A(n14208), .B(n14207), .Z(n14212) );
  OR U14602 ( .A(n14210), .B(n14209), .Z(n14211) );
  AND U14603 ( .A(n14212), .B(n14211), .Z(n14257) );
  XNOR U14604 ( .A(n14258), .B(n14257), .Z(n14260) );
  NAND U14605 ( .A(n14213), .B(n19724), .Z(n14215) );
  XOR U14606 ( .A(b[11]), .B(a[182]), .Z(n14290) );
  NAND U14607 ( .A(n19692), .B(n14290), .Z(n14214) );
  AND U14608 ( .A(n14215), .B(n14214), .Z(n14301) );
  NAND U14609 ( .A(n19838), .B(n14216), .Z(n14218) );
  XOR U14610 ( .A(b[15]), .B(a[178]), .Z(n14293) );
  NAND U14611 ( .A(n19805), .B(n14293), .Z(n14217) );
  AND U14612 ( .A(n14218), .B(n14217), .Z(n14300) );
  NAND U14613 ( .A(n35), .B(n14219), .Z(n14221) );
  XOR U14614 ( .A(b[9]), .B(a[184]), .Z(n14296) );
  NAND U14615 ( .A(n19598), .B(n14296), .Z(n14220) );
  NAND U14616 ( .A(n14221), .B(n14220), .Z(n14299) );
  XOR U14617 ( .A(n14300), .B(n14299), .Z(n14302) );
  XOR U14618 ( .A(n14301), .B(n14302), .Z(n14312) );
  NANDN U14619 ( .A(n14223), .B(n14222), .Z(n14227) );
  OR U14620 ( .A(n14225), .B(n14224), .Z(n14226) );
  AND U14621 ( .A(n14227), .B(n14226), .Z(n14311) );
  XNOR U14622 ( .A(n14312), .B(n14311), .Z(n14313) );
  NANDN U14623 ( .A(n14229), .B(n14228), .Z(n14233) );
  NANDN U14624 ( .A(n14231), .B(n14230), .Z(n14232) );
  NAND U14625 ( .A(n14233), .B(n14232), .Z(n14314) );
  XNOR U14626 ( .A(n14313), .B(n14314), .Z(n14259) );
  XOR U14627 ( .A(n14260), .B(n14259), .Z(n14318) );
  NANDN U14628 ( .A(n14235), .B(n14234), .Z(n14239) );
  NANDN U14629 ( .A(n14237), .B(n14236), .Z(n14238) );
  AND U14630 ( .A(n14239), .B(n14238), .Z(n14317) );
  XNOR U14631 ( .A(n14318), .B(n14317), .Z(n14319) );
  XOR U14632 ( .A(n14320), .B(n14319), .Z(n14252) );
  NANDN U14633 ( .A(n14241), .B(n14240), .Z(n14245) );
  NAND U14634 ( .A(n14243), .B(n14242), .Z(n14244) );
  AND U14635 ( .A(n14245), .B(n14244), .Z(n14251) );
  XNOR U14636 ( .A(n14252), .B(n14251), .Z(n14253) );
  XNOR U14637 ( .A(n14254), .B(n14253), .Z(n14323) );
  XNOR U14638 ( .A(sreg[432]), .B(n14323), .Z(n14325) );
  NANDN U14639 ( .A(sreg[431]), .B(n14246), .Z(n14250) );
  NAND U14640 ( .A(n14248), .B(n14247), .Z(n14249) );
  NAND U14641 ( .A(n14250), .B(n14249), .Z(n14324) );
  XNOR U14642 ( .A(n14325), .B(n14324), .Z(c[432]) );
  NANDN U14643 ( .A(n14252), .B(n14251), .Z(n14256) );
  NANDN U14644 ( .A(n14254), .B(n14253), .Z(n14255) );
  AND U14645 ( .A(n14256), .B(n14255), .Z(n14331) );
  NANDN U14646 ( .A(n14258), .B(n14257), .Z(n14262) );
  NAND U14647 ( .A(n14260), .B(n14259), .Z(n14261) );
  AND U14648 ( .A(n14262), .B(n14261), .Z(n14397) );
  NANDN U14649 ( .A(n14264), .B(n14263), .Z(n14268) );
  NANDN U14650 ( .A(n14266), .B(n14265), .Z(n14267) );
  AND U14651 ( .A(n14268), .B(n14267), .Z(n14363) );
  NAND U14652 ( .A(b[0]), .B(a[193]), .Z(n14269) );
  XNOR U14653 ( .A(b[1]), .B(n14269), .Z(n14271) );
  NANDN U14654 ( .A(b[0]), .B(a[192]), .Z(n14270) );
  NAND U14655 ( .A(n14271), .B(n14270), .Z(n14343) );
  NAND U14656 ( .A(n19808), .B(n14272), .Z(n14274) );
  XOR U14657 ( .A(b[13]), .B(a[181]), .Z(n14349) );
  NAND U14658 ( .A(n19768), .B(n14349), .Z(n14273) );
  AND U14659 ( .A(n14274), .B(n14273), .Z(n14341) );
  AND U14660 ( .A(b[15]), .B(a[177]), .Z(n14340) );
  XNOR U14661 ( .A(n14341), .B(n14340), .Z(n14342) );
  XNOR U14662 ( .A(n14343), .B(n14342), .Z(n14361) );
  NAND U14663 ( .A(n33), .B(n14275), .Z(n14277) );
  XOR U14664 ( .A(b[5]), .B(a[189]), .Z(n14352) );
  NAND U14665 ( .A(n19342), .B(n14352), .Z(n14276) );
  AND U14666 ( .A(n14277), .B(n14276), .Z(n14385) );
  NAND U14667 ( .A(n34), .B(n14278), .Z(n14280) );
  XOR U14668 ( .A(b[7]), .B(a[187]), .Z(n14355) );
  NAND U14669 ( .A(n19486), .B(n14355), .Z(n14279) );
  AND U14670 ( .A(n14280), .B(n14279), .Z(n14383) );
  NAND U14671 ( .A(n31), .B(n14281), .Z(n14283) );
  XOR U14672 ( .A(b[3]), .B(a[191]), .Z(n14358) );
  NAND U14673 ( .A(n32), .B(n14358), .Z(n14282) );
  NAND U14674 ( .A(n14283), .B(n14282), .Z(n14382) );
  XNOR U14675 ( .A(n14383), .B(n14382), .Z(n14384) );
  XOR U14676 ( .A(n14385), .B(n14384), .Z(n14362) );
  XOR U14677 ( .A(n14361), .B(n14362), .Z(n14364) );
  XOR U14678 ( .A(n14363), .B(n14364), .Z(n14335) );
  NANDN U14679 ( .A(n14285), .B(n14284), .Z(n14289) );
  OR U14680 ( .A(n14287), .B(n14286), .Z(n14288) );
  AND U14681 ( .A(n14289), .B(n14288), .Z(n14334) );
  XNOR U14682 ( .A(n14335), .B(n14334), .Z(n14337) );
  NAND U14683 ( .A(n14290), .B(n19724), .Z(n14292) );
  XOR U14684 ( .A(b[11]), .B(a[183]), .Z(n14367) );
  NAND U14685 ( .A(n19692), .B(n14367), .Z(n14291) );
  AND U14686 ( .A(n14292), .B(n14291), .Z(n14378) );
  NAND U14687 ( .A(n19838), .B(n14293), .Z(n14295) );
  XOR U14688 ( .A(b[15]), .B(a[179]), .Z(n14370) );
  NAND U14689 ( .A(n19805), .B(n14370), .Z(n14294) );
  AND U14690 ( .A(n14295), .B(n14294), .Z(n14377) );
  NAND U14691 ( .A(n35), .B(n14296), .Z(n14298) );
  XOR U14692 ( .A(b[9]), .B(a[185]), .Z(n14373) );
  NAND U14693 ( .A(n19598), .B(n14373), .Z(n14297) );
  NAND U14694 ( .A(n14298), .B(n14297), .Z(n14376) );
  XOR U14695 ( .A(n14377), .B(n14376), .Z(n14379) );
  XOR U14696 ( .A(n14378), .B(n14379), .Z(n14389) );
  NANDN U14697 ( .A(n14300), .B(n14299), .Z(n14304) );
  OR U14698 ( .A(n14302), .B(n14301), .Z(n14303) );
  AND U14699 ( .A(n14304), .B(n14303), .Z(n14388) );
  XNOR U14700 ( .A(n14389), .B(n14388), .Z(n14390) );
  NANDN U14701 ( .A(n14306), .B(n14305), .Z(n14310) );
  NANDN U14702 ( .A(n14308), .B(n14307), .Z(n14309) );
  NAND U14703 ( .A(n14310), .B(n14309), .Z(n14391) );
  XNOR U14704 ( .A(n14390), .B(n14391), .Z(n14336) );
  XOR U14705 ( .A(n14337), .B(n14336), .Z(n14395) );
  NANDN U14706 ( .A(n14312), .B(n14311), .Z(n14316) );
  NANDN U14707 ( .A(n14314), .B(n14313), .Z(n14315) );
  AND U14708 ( .A(n14316), .B(n14315), .Z(n14394) );
  XNOR U14709 ( .A(n14395), .B(n14394), .Z(n14396) );
  XOR U14710 ( .A(n14397), .B(n14396), .Z(n14329) );
  NANDN U14711 ( .A(n14318), .B(n14317), .Z(n14322) );
  NAND U14712 ( .A(n14320), .B(n14319), .Z(n14321) );
  AND U14713 ( .A(n14322), .B(n14321), .Z(n14328) );
  XNOR U14714 ( .A(n14329), .B(n14328), .Z(n14330) );
  XNOR U14715 ( .A(n14331), .B(n14330), .Z(n14400) );
  XNOR U14716 ( .A(sreg[433]), .B(n14400), .Z(n14402) );
  NANDN U14717 ( .A(sreg[432]), .B(n14323), .Z(n14327) );
  NAND U14718 ( .A(n14325), .B(n14324), .Z(n14326) );
  NAND U14719 ( .A(n14327), .B(n14326), .Z(n14401) );
  XNOR U14720 ( .A(n14402), .B(n14401), .Z(c[433]) );
  NANDN U14721 ( .A(n14329), .B(n14328), .Z(n14333) );
  NANDN U14722 ( .A(n14331), .B(n14330), .Z(n14332) );
  AND U14723 ( .A(n14333), .B(n14332), .Z(n14408) );
  NANDN U14724 ( .A(n14335), .B(n14334), .Z(n14339) );
  NAND U14725 ( .A(n14337), .B(n14336), .Z(n14338) );
  AND U14726 ( .A(n14339), .B(n14338), .Z(n14474) );
  NANDN U14727 ( .A(n14341), .B(n14340), .Z(n14345) );
  NANDN U14728 ( .A(n14343), .B(n14342), .Z(n14344) );
  AND U14729 ( .A(n14345), .B(n14344), .Z(n14440) );
  NAND U14730 ( .A(b[0]), .B(a[194]), .Z(n14346) );
  XNOR U14731 ( .A(b[1]), .B(n14346), .Z(n14348) );
  NANDN U14732 ( .A(b[0]), .B(a[193]), .Z(n14347) );
  NAND U14733 ( .A(n14348), .B(n14347), .Z(n14420) );
  NAND U14734 ( .A(n19808), .B(n14349), .Z(n14351) );
  XOR U14735 ( .A(b[13]), .B(a[182]), .Z(n14426) );
  NAND U14736 ( .A(n19768), .B(n14426), .Z(n14350) );
  AND U14737 ( .A(n14351), .B(n14350), .Z(n14418) );
  AND U14738 ( .A(b[15]), .B(a[178]), .Z(n14417) );
  XNOR U14739 ( .A(n14418), .B(n14417), .Z(n14419) );
  XNOR U14740 ( .A(n14420), .B(n14419), .Z(n14438) );
  NAND U14741 ( .A(n33), .B(n14352), .Z(n14354) );
  XOR U14742 ( .A(b[5]), .B(a[190]), .Z(n14429) );
  NAND U14743 ( .A(n19342), .B(n14429), .Z(n14353) );
  AND U14744 ( .A(n14354), .B(n14353), .Z(n14462) );
  NAND U14745 ( .A(n34), .B(n14355), .Z(n14357) );
  XOR U14746 ( .A(b[7]), .B(a[188]), .Z(n14432) );
  NAND U14747 ( .A(n19486), .B(n14432), .Z(n14356) );
  AND U14748 ( .A(n14357), .B(n14356), .Z(n14460) );
  NAND U14749 ( .A(n31), .B(n14358), .Z(n14360) );
  XOR U14750 ( .A(b[3]), .B(a[192]), .Z(n14435) );
  NAND U14751 ( .A(n32), .B(n14435), .Z(n14359) );
  NAND U14752 ( .A(n14360), .B(n14359), .Z(n14459) );
  XNOR U14753 ( .A(n14460), .B(n14459), .Z(n14461) );
  XOR U14754 ( .A(n14462), .B(n14461), .Z(n14439) );
  XOR U14755 ( .A(n14438), .B(n14439), .Z(n14441) );
  XOR U14756 ( .A(n14440), .B(n14441), .Z(n14412) );
  NANDN U14757 ( .A(n14362), .B(n14361), .Z(n14366) );
  OR U14758 ( .A(n14364), .B(n14363), .Z(n14365) );
  AND U14759 ( .A(n14366), .B(n14365), .Z(n14411) );
  XNOR U14760 ( .A(n14412), .B(n14411), .Z(n14414) );
  NAND U14761 ( .A(n14367), .B(n19724), .Z(n14369) );
  XOR U14762 ( .A(b[11]), .B(a[184]), .Z(n14444) );
  NAND U14763 ( .A(n19692), .B(n14444), .Z(n14368) );
  AND U14764 ( .A(n14369), .B(n14368), .Z(n14455) );
  NAND U14765 ( .A(n19838), .B(n14370), .Z(n14372) );
  XOR U14766 ( .A(b[15]), .B(a[180]), .Z(n14447) );
  NAND U14767 ( .A(n19805), .B(n14447), .Z(n14371) );
  AND U14768 ( .A(n14372), .B(n14371), .Z(n14454) );
  NAND U14769 ( .A(n35), .B(n14373), .Z(n14375) );
  XOR U14770 ( .A(b[9]), .B(a[186]), .Z(n14450) );
  NAND U14771 ( .A(n19598), .B(n14450), .Z(n14374) );
  NAND U14772 ( .A(n14375), .B(n14374), .Z(n14453) );
  XOR U14773 ( .A(n14454), .B(n14453), .Z(n14456) );
  XOR U14774 ( .A(n14455), .B(n14456), .Z(n14466) );
  NANDN U14775 ( .A(n14377), .B(n14376), .Z(n14381) );
  OR U14776 ( .A(n14379), .B(n14378), .Z(n14380) );
  AND U14777 ( .A(n14381), .B(n14380), .Z(n14465) );
  XNOR U14778 ( .A(n14466), .B(n14465), .Z(n14467) );
  NANDN U14779 ( .A(n14383), .B(n14382), .Z(n14387) );
  NANDN U14780 ( .A(n14385), .B(n14384), .Z(n14386) );
  NAND U14781 ( .A(n14387), .B(n14386), .Z(n14468) );
  XNOR U14782 ( .A(n14467), .B(n14468), .Z(n14413) );
  XOR U14783 ( .A(n14414), .B(n14413), .Z(n14472) );
  NANDN U14784 ( .A(n14389), .B(n14388), .Z(n14393) );
  NANDN U14785 ( .A(n14391), .B(n14390), .Z(n14392) );
  AND U14786 ( .A(n14393), .B(n14392), .Z(n14471) );
  XNOR U14787 ( .A(n14472), .B(n14471), .Z(n14473) );
  XOR U14788 ( .A(n14474), .B(n14473), .Z(n14406) );
  NANDN U14789 ( .A(n14395), .B(n14394), .Z(n14399) );
  NAND U14790 ( .A(n14397), .B(n14396), .Z(n14398) );
  AND U14791 ( .A(n14399), .B(n14398), .Z(n14405) );
  XNOR U14792 ( .A(n14406), .B(n14405), .Z(n14407) );
  XNOR U14793 ( .A(n14408), .B(n14407), .Z(n14477) );
  XNOR U14794 ( .A(sreg[434]), .B(n14477), .Z(n14479) );
  NANDN U14795 ( .A(sreg[433]), .B(n14400), .Z(n14404) );
  NAND U14796 ( .A(n14402), .B(n14401), .Z(n14403) );
  NAND U14797 ( .A(n14404), .B(n14403), .Z(n14478) );
  XNOR U14798 ( .A(n14479), .B(n14478), .Z(c[434]) );
  NANDN U14799 ( .A(n14406), .B(n14405), .Z(n14410) );
  NANDN U14800 ( .A(n14408), .B(n14407), .Z(n14409) );
  AND U14801 ( .A(n14410), .B(n14409), .Z(n14485) );
  NANDN U14802 ( .A(n14412), .B(n14411), .Z(n14416) );
  NAND U14803 ( .A(n14414), .B(n14413), .Z(n14415) );
  AND U14804 ( .A(n14416), .B(n14415), .Z(n14551) );
  NANDN U14805 ( .A(n14418), .B(n14417), .Z(n14422) );
  NANDN U14806 ( .A(n14420), .B(n14419), .Z(n14421) );
  AND U14807 ( .A(n14422), .B(n14421), .Z(n14517) );
  NAND U14808 ( .A(b[0]), .B(a[195]), .Z(n14423) );
  XNOR U14809 ( .A(b[1]), .B(n14423), .Z(n14425) );
  NANDN U14810 ( .A(b[0]), .B(a[194]), .Z(n14424) );
  NAND U14811 ( .A(n14425), .B(n14424), .Z(n14497) );
  NAND U14812 ( .A(n19808), .B(n14426), .Z(n14428) );
  XOR U14813 ( .A(b[13]), .B(a[183]), .Z(n14500) );
  NAND U14814 ( .A(n19768), .B(n14500), .Z(n14427) );
  AND U14815 ( .A(n14428), .B(n14427), .Z(n14495) );
  AND U14816 ( .A(b[15]), .B(a[179]), .Z(n14494) );
  XNOR U14817 ( .A(n14495), .B(n14494), .Z(n14496) );
  XNOR U14818 ( .A(n14497), .B(n14496), .Z(n14515) );
  NAND U14819 ( .A(n33), .B(n14429), .Z(n14431) );
  XOR U14820 ( .A(b[5]), .B(a[191]), .Z(n14506) );
  NAND U14821 ( .A(n19342), .B(n14506), .Z(n14430) );
  AND U14822 ( .A(n14431), .B(n14430), .Z(n14539) );
  NAND U14823 ( .A(n34), .B(n14432), .Z(n14434) );
  XOR U14824 ( .A(b[7]), .B(a[189]), .Z(n14509) );
  NAND U14825 ( .A(n19486), .B(n14509), .Z(n14433) );
  AND U14826 ( .A(n14434), .B(n14433), .Z(n14537) );
  NAND U14827 ( .A(n31), .B(n14435), .Z(n14437) );
  XOR U14828 ( .A(b[3]), .B(a[193]), .Z(n14512) );
  NAND U14829 ( .A(n32), .B(n14512), .Z(n14436) );
  NAND U14830 ( .A(n14437), .B(n14436), .Z(n14536) );
  XNOR U14831 ( .A(n14537), .B(n14536), .Z(n14538) );
  XOR U14832 ( .A(n14539), .B(n14538), .Z(n14516) );
  XOR U14833 ( .A(n14515), .B(n14516), .Z(n14518) );
  XOR U14834 ( .A(n14517), .B(n14518), .Z(n14489) );
  NANDN U14835 ( .A(n14439), .B(n14438), .Z(n14443) );
  OR U14836 ( .A(n14441), .B(n14440), .Z(n14442) );
  AND U14837 ( .A(n14443), .B(n14442), .Z(n14488) );
  XNOR U14838 ( .A(n14489), .B(n14488), .Z(n14491) );
  NAND U14839 ( .A(n14444), .B(n19724), .Z(n14446) );
  XOR U14840 ( .A(b[11]), .B(a[185]), .Z(n14521) );
  NAND U14841 ( .A(n19692), .B(n14521), .Z(n14445) );
  AND U14842 ( .A(n14446), .B(n14445), .Z(n14532) );
  NAND U14843 ( .A(n19838), .B(n14447), .Z(n14449) );
  XOR U14844 ( .A(b[15]), .B(a[181]), .Z(n14524) );
  NAND U14845 ( .A(n19805), .B(n14524), .Z(n14448) );
  AND U14846 ( .A(n14449), .B(n14448), .Z(n14531) );
  NAND U14847 ( .A(n35), .B(n14450), .Z(n14452) );
  XOR U14848 ( .A(b[9]), .B(a[187]), .Z(n14527) );
  NAND U14849 ( .A(n19598), .B(n14527), .Z(n14451) );
  NAND U14850 ( .A(n14452), .B(n14451), .Z(n14530) );
  XOR U14851 ( .A(n14531), .B(n14530), .Z(n14533) );
  XOR U14852 ( .A(n14532), .B(n14533), .Z(n14543) );
  NANDN U14853 ( .A(n14454), .B(n14453), .Z(n14458) );
  OR U14854 ( .A(n14456), .B(n14455), .Z(n14457) );
  AND U14855 ( .A(n14458), .B(n14457), .Z(n14542) );
  XNOR U14856 ( .A(n14543), .B(n14542), .Z(n14544) );
  NANDN U14857 ( .A(n14460), .B(n14459), .Z(n14464) );
  NANDN U14858 ( .A(n14462), .B(n14461), .Z(n14463) );
  NAND U14859 ( .A(n14464), .B(n14463), .Z(n14545) );
  XNOR U14860 ( .A(n14544), .B(n14545), .Z(n14490) );
  XOR U14861 ( .A(n14491), .B(n14490), .Z(n14549) );
  NANDN U14862 ( .A(n14466), .B(n14465), .Z(n14470) );
  NANDN U14863 ( .A(n14468), .B(n14467), .Z(n14469) );
  AND U14864 ( .A(n14470), .B(n14469), .Z(n14548) );
  XNOR U14865 ( .A(n14549), .B(n14548), .Z(n14550) );
  XOR U14866 ( .A(n14551), .B(n14550), .Z(n14483) );
  NANDN U14867 ( .A(n14472), .B(n14471), .Z(n14476) );
  NAND U14868 ( .A(n14474), .B(n14473), .Z(n14475) );
  AND U14869 ( .A(n14476), .B(n14475), .Z(n14482) );
  XNOR U14870 ( .A(n14483), .B(n14482), .Z(n14484) );
  XNOR U14871 ( .A(n14485), .B(n14484), .Z(n14554) );
  XNOR U14872 ( .A(sreg[435]), .B(n14554), .Z(n14556) );
  NANDN U14873 ( .A(sreg[434]), .B(n14477), .Z(n14481) );
  NAND U14874 ( .A(n14479), .B(n14478), .Z(n14480) );
  NAND U14875 ( .A(n14481), .B(n14480), .Z(n14555) );
  XNOR U14876 ( .A(n14556), .B(n14555), .Z(c[435]) );
  NANDN U14877 ( .A(n14483), .B(n14482), .Z(n14487) );
  NANDN U14878 ( .A(n14485), .B(n14484), .Z(n14486) );
  AND U14879 ( .A(n14487), .B(n14486), .Z(n14562) );
  NANDN U14880 ( .A(n14489), .B(n14488), .Z(n14493) );
  NAND U14881 ( .A(n14491), .B(n14490), .Z(n14492) );
  AND U14882 ( .A(n14493), .B(n14492), .Z(n14628) );
  NANDN U14883 ( .A(n14495), .B(n14494), .Z(n14499) );
  NANDN U14884 ( .A(n14497), .B(n14496), .Z(n14498) );
  AND U14885 ( .A(n14499), .B(n14498), .Z(n14594) );
  NAND U14886 ( .A(n19808), .B(n14500), .Z(n14502) );
  XOR U14887 ( .A(b[13]), .B(a[184]), .Z(n14580) );
  NAND U14888 ( .A(n19768), .B(n14580), .Z(n14501) );
  AND U14889 ( .A(n14502), .B(n14501), .Z(n14572) );
  AND U14890 ( .A(b[15]), .B(a[180]), .Z(n14571) );
  XNOR U14891 ( .A(n14572), .B(n14571), .Z(n14573) );
  NAND U14892 ( .A(b[0]), .B(a[196]), .Z(n14503) );
  XNOR U14893 ( .A(b[1]), .B(n14503), .Z(n14505) );
  NANDN U14894 ( .A(b[0]), .B(a[195]), .Z(n14504) );
  NAND U14895 ( .A(n14505), .B(n14504), .Z(n14574) );
  XNOR U14896 ( .A(n14573), .B(n14574), .Z(n14592) );
  NAND U14897 ( .A(n33), .B(n14506), .Z(n14508) );
  XOR U14898 ( .A(b[5]), .B(a[192]), .Z(n14583) );
  NAND U14899 ( .A(n19342), .B(n14583), .Z(n14507) );
  AND U14900 ( .A(n14508), .B(n14507), .Z(n14616) );
  NAND U14901 ( .A(n34), .B(n14509), .Z(n14511) );
  XOR U14902 ( .A(b[7]), .B(a[190]), .Z(n14586) );
  NAND U14903 ( .A(n19486), .B(n14586), .Z(n14510) );
  AND U14904 ( .A(n14511), .B(n14510), .Z(n14614) );
  NAND U14905 ( .A(n31), .B(n14512), .Z(n14514) );
  XOR U14906 ( .A(b[3]), .B(a[194]), .Z(n14589) );
  NAND U14907 ( .A(n32), .B(n14589), .Z(n14513) );
  NAND U14908 ( .A(n14514), .B(n14513), .Z(n14613) );
  XNOR U14909 ( .A(n14614), .B(n14613), .Z(n14615) );
  XOR U14910 ( .A(n14616), .B(n14615), .Z(n14593) );
  XOR U14911 ( .A(n14592), .B(n14593), .Z(n14595) );
  XOR U14912 ( .A(n14594), .B(n14595), .Z(n14566) );
  NANDN U14913 ( .A(n14516), .B(n14515), .Z(n14520) );
  OR U14914 ( .A(n14518), .B(n14517), .Z(n14519) );
  AND U14915 ( .A(n14520), .B(n14519), .Z(n14565) );
  XNOR U14916 ( .A(n14566), .B(n14565), .Z(n14568) );
  NAND U14917 ( .A(n14521), .B(n19724), .Z(n14523) );
  XOR U14918 ( .A(b[11]), .B(a[186]), .Z(n14598) );
  NAND U14919 ( .A(n19692), .B(n14598), .Z(n14522) );
  AND U14920 ( .A(n14523), .B(n14522), .Z(n14609) );
  NAND U14921 ( .A(n19838), .B(n14524), .Z(n14526) );
  XOR U14922 ( .A(b[15]), .B(a[182]), .Z(n14601) );
  NAND U14923 ( .A(n19805), .B(n14601), .Z(n14525) );
  AND U14924 ( .A(n14526), .B(n14525), .Z(n14608) );
  NAND U14925 ( .A(n35), .B(n14527), .Z(n14529) );
  XOR U14926 ( .A(b[9]), .B(a[188]), .Z(n14604) );
  NAND U14927 ( .A(n19598), .B(n14604), .Z(n14528) );
  NAND U14928 ( .A(n14529), .B(n14528), .Z(n14607) );
  XOR U14929 ( .A(n14608), .B(n14607), .Z(n14610) );
  XOR U14930 ( .A(n14609), .B(n14610), .Z(n14620) );
  NANDN U14931 ( .A(n14531), .B(n14530), .Z(n14535) );
  OR U14932 ( .A(n14533), .B(n14532), .Z(n14534) );
  AND U14933 ( .A(n14535), .B(n14534), .Z(n14619) );
  XNOR U14934 ( .A(n14620), .B(n14619), .Z(n14621) );
  NANDN U14935 ( .A(n14537), .B(n14536), .Z(n14541) );
  NANDN U14936 ( .A(n14539), .B(n14538), .Z(n14540) );
  NAND U14937 ( .A(n14541), .B(n14540), .Z(n14622) );
  XNOR U14938 ( .A(n14621), .B(n14622), .Z(n14567) );
  XOR U14939 ( .A(n14568), .B(n14567), .Z(n14626) );
  NANDN U14940 ( .A(n14543), .B(n14542), .Z(n14547) );
  NANDN U14941 ( .A(n14545), .B(n14544), .Z(n14546) );
  AND U14942 ( .A(n14547), .B(n14546), .Z(n14625) );
  XNOR U14943 ( .A(n14626), .B(n14625), .Z(n14627) );
  XOR U14944 ( .A(n14628), .B(n14627), .Z(n14560) );
  NANDN U14945 ( .A(n14549), .B(n14548), .Z(n14553) );
  NAND U14946 ( .A(n14551), .B(n14550), .Z(n14552) );
  AND U14947 ( .A(n14553), .B(n14552), .Z(n14559) );
  XNOR U14948 ( .A(n14560), .B(n14559), .Z(n14561) );
  XNOR U14949 ( .A(n14562), .B(n14561), .Z(n14631) );
  XNOR U14950 ( .A(sreg[436]), .B(n14631), .Z(n14633) );
  NANDN U14951 ( .A(sreg[435]), .B(n14554), .Z(n14558) );
  NAND U14952 ( .A(n14556), .B(n14555), .Z(n14557) );
  NAND U14953 ( .A(n14558), .B(n14557), .Z(n14632) );
  XNOR U14954 ( .A(n14633), .B(n14632), .Z(c[436]) );
  NANDN U14955 ( .A(n14560), .B(n14559), .Z(n14564) );
  NANDN U14956 ( .A(n14562), .B(n14561), .Z(n14563) );
  AND U14957 ( .A(n14564), .B(n14563), .Z(n14639) );
  NANDN U14958 ( .A(n14566), .B(n14565), .Z(n14570) );
  NAND U14959 ( .A(n14568), .B(n14567), .Z(n14569) );
  AND U14960 ( .A(n14570), .B(n14569), .Z(n14705) );
  NANDN U14961 ( .A(n14572), .B(n14571), .Z(n14576) );
  NANDN U14962 ( .A(n14574), .B(n14573), .Z(n14575) );
  AND U14963 ( .A(n14576), .B(n14575), .Z(n14671) );
  NAND U14964 ( .A(b[0]), .B(a[197]), .Z(n14577) );
  XNOR U14965 ( .A(b[1]), .B(n14577), .Z(n14579) );
  NANDN U14966 ( .A(b[0]), .B(a[196]), .Z(n14578) );
  NAND U14967 ( .A(n14579), .B(n14578), .Z(n14651) );
  NAND U14968 ( .A(n19808), .B(n14580), .Z(n14582) );
  XOR U14969 ( .A(b[13]), .B(a[185]), .Z(n14657) );
  NAND U14970 ( .A(n19768), .B(n14657), .Z(n14581) );
  AND U14971 ( .A(n14582), .B(n14581), .Z(n14649) );
  AND U14972 ( .A(b[15]), .B(a[181]), .Z(n14648) );
  XNOR U14973 ( .A(n14649), .B(n14648), .Z(n14650) );
  XNOR U14974 ( .A(n14651), .B(n14650), .Z(n14669) );
  NAND U14975 ( .A(n33), .B(n14583), .Z(n14585) );
  XOR U14976 ( .A(b[5]), .B(a[193]), .Z(n14660) );
  NAND U14977 ( .A(n19342), .B(n14660), .Z(n14584) );
  AND U14978 ( .A(n14585), .B(n14584), .Z(n14693) );
  NAND U14979 ( .A(n34), .B(n14586), .Z(n14588) );
  XOR U14980 ( .A(b[7]), .B(a[191]), .Z(n14663) );
  NAND U14981 ( .A(n19486), .B(n14663), .Z(n14587) );
  AND U14982 ( .A(n14588), .B(n14587), .Z(n14691) );
  NAND U14983 ( .A(n31), .B(n14589), .Z(n14591) );
  XOR U14984 ( .A(b[3]), .B(a[195]), .Z(n14666) );
  NAND U14985 ( .A(n32), .B(n14666), .Z(n14590) );
  NAND U14986 ( .A(n14591), .B(n14590), .Z(n14690) );
  XNOR U14987 ( .A(n14691), .B(n14690), .Z(n14692) );
  XOR U14988 ( .A(n14693), .B(n14692), .Z(n14670) );
  XOR U14989 ( .A(n14669), .B(n14670), .Z(n14672) );
  XOR U14990 ( .A(n14671), .B(n14672), .Z(n14643) );
  NANDN U14991 ( .A(n14593), .B(n14592), .Z(n14597) );
  OR U14992 ( .A(n14595), .B(n14594), .Z(n14596) );
  AND U14993 ( .A(n14597), .B(n14596), .Z(n14642) );
  XNOR U14994 ( .A(n14643), .B(n14642), .Z(n14645) );
  NAND U14995 ( .A(n14598), .B(n19724), .Z(n14600) );
  XOR U14996 ( .A(b[11]), .B(a[187]), .Z(n14675) );
  NAND U14997 ( .A(n19692), .B(n14675), .Z(n14599) );
  AND U14998 ( .A(n14600), .B(n14599), .Z(n14686) );
  NAND U14999 ( .A(n19838), .B(n14601), .Z(n14603) );
  XOR U15000 ( .A(b[15]), .B(a[183]), .Z(n14678) );
  NAND U15001 ( .A(n19805), .B(n14678), .Z(n14602) );
  AND U15002 ( .A(n14603), .B(n14602), .Z(n14685) );
  NAND U15003 ( .A(n35), .B(n14604), .Z(n14606) );
  XOR U15004 ( .A(b[9]), .B(a[189]), .Z(n14681) );
  NAND U15005 ( .A(n19598), .B(n14681), .Z(n14605) );
  NAND U15006 ( .A(n14606), .B(n14605), .Z(n14684) );
  XOR U15007 ( .A(n14685), .B(n14684), .Z(n14687) );
  XOR U15008 ( .A(n14686), .B(n14687), .Z(n14697) );
  NANDN U15009 ( .A(n14608), .B(n14607), .Z(n14612) );
  OR U15010 ( .A(n14610), .B(n14609), .Z(n14611) );
  AND U15011 ( .A(n14612), .B(n14611), .Z(n14696) );
  XNOR U15012 ( .A(n14697), .B(n14696), .Z(n14698) );
  NANDN U15013 ( .A(n14614), .B(n14613), .Z(n14618) );
  NANDN U15014 ( .A(n14616), .B(n14615), .Z(n14617) );
  NAND U15015 ( .A(n14618), .B(n14617), .Z(n14699) );
  XNOR U15016 ( .A(n14698), .B(n14699), .Z(n14644) );
  XOR U15017 ( .A(n14645), .B(n14644), .Z(n14703) );
  NANDN U15018 ( .A(n14620), .B(n14619), .Z(n14624) );
  NANDN U15019 ( .A(n14622), .B(n14621), .Z(n14623) );
  AND U15020 ( .A(n14624), .B(n14623), .Z(n14702) );
  XNOR U15021 ( .A(n14703), .B(n14702), .Z(n14704) );
  XOR U15022 ( .A(n14705), .B(n14704), .Z(n14637) );
  NANDN U15023 ( .A(n14626), .B(n14625), .Z(n14630) );
  NAND U15024 ( .A(n14628), .B(n14627), .Z(n14629) );
  AND U15025 ( .A(n14630), .B(n14629), .Z(n14636) );
  XNOR U15026 ( .A(n14637), .B(n14636), .Z(n14638) );
  XNOR U15027 ( .A(n14639), .B(n14638), .Z(n14708) );
  XNOR U15028 ( .A(sreg[437]), .B(n14708), .Z(n14710) );
  NANDN U15029 ( .A(sreg[436]), .B(n14631), .Z(n14635) );
  NAND U15030 ( .A(n14633), .B(n14632), .Z(n14634) );
  NAND U15031 ( .A(n14635), .B(n14634), .Z(n14709) );
  XNOR U15032 ( .A(n14710), .B(n14709), .Z(c[437]) );
  NANDN U15033 ( .A(n14637), .B(n14636), .Z(n14641) );
  NANDN U15034 ( .A(n14639), .B(n14638), .Z(n14640) );
  AND U15035 ( .A(n14641), .B(n14640), .Z(n14716) );
  NANDN U15036 ( .A(n14643), .B(n14642), .Z(n14647) );
  NAND U15037 ( .A(n14645), .B(n14644), .Z(n14646) );
  AND U15038 ( .A(n14647), .B(n14646), .Z(n14782) );
  NANDN U15039 ( .A(n14649), .B(n14648), .Z(n14653) );
  NANDN U15040 ( .A(n14651), .B(n14650), .Z(n14652) );
  AND U15041 ( .A(n14653), .B(n14652), .Z(n14748) );
  NAND U15042 ( .A(b[0]), .B(a[198]), .Z(n14654) );
  XNOR U15043 ( .A(b[1]), .B(n14654), .Z(n14656) );
  NANDN U15044 ( .A(b[0]), .B(a[197]), .Z(n14655) );
  NAND U15045 ( .A(n14656), .B(n14655), .Z(n14728) );
  NAND U15046 ( .A(n19808), .B(n14657), .Z(n14659) );
  XOR U15047 ( .A(b[13]), .B(a[186]), .Z(n14734) );
  NAND U15048 ( .A(n19768), .B(n14734), .Z(n14658) );
  AND U15049 ( .A(n14659), .B(n14658), .Z(n14726) );
  AND U15050 ( .A(b[15]), .B(a[182]), .Z(n14725) );
  XNOR U15051 ( .A(n14726), .B(n14725), .Z(n14727) );
  XNOR U15052 ( .A(n14728), .B(n14727), .Z(n14746) );
  NAND U15053 ( .A(n33), .B(n14660), .Z(n14662) );
  XOR U15054 ( .A(b[5]), .B(a[194]), .Z(n14737) );
  NAND U15055 ( .A(n19342), .B(n14737), .Z(n14661) );
  AND U15056 ( .A(n14662), .B(n14661), .Z(n14770) );
  NAND U15057 ( .A(n34), .B(n14663), .Z(n14665) );
  XOR U15058 ( .A(b[7]), .B(a[192]), .Z(n14740) );
  NAND U15059 ( .A(n19486), .B(n14740), .Z(n14664) );
  AND U15060 ( .A(n14665), .B(n14664), .Z(n14768) );
  NAND U15061 ( .A(n31), .B(n14666), .Z(n14668) );
  XOR U15062 ( .A(b[3]), .B(a[196]), .Z(n14743) );
  NAND U15063 ( .A(n32), .B(n14743), .Z(n14667) );
  NAND U15064 ( .A(n14668), .B(n14667), .Z(n14767) );
  XNOR U15065 ( .A(n14768), .B(n14767), .Z(n14769) );
  XOR U15066 ( .A(n14770), .B(n14769), .Z(n14747) );
  XOR U15067 ( .A(n14746), .B(n14747), .Z(n14749) );
  XOR U15068 ( .A(n14748), .B(n14749), .Z(n14720) );
  NANDN U15069 ( .A(n14670), .B(n14669), .Z(n14674) );
  OR U15070 ( .A(n14672), .B(n14671), .Z(n14673) );
  AND U15071 ( .A(n14674), .B(n14673), .Z(n14719) );
  XNOR U15072 ( .A(n14720), .B(n14719), .Z(n14722) );
  NAND U15073 ( .A(n14675), .B(n19724), .Z(n14677) );
  XOR U15074 ( .A(b[11]), .B(a[188]), .Z(n14752) );
  NAND U15075 ( .A(n19692), .B(n14752), .Z(n14676) );
  AND U15076 ( .A(n14677), .B(n14676), .Z(n14763) );
  NAND U15077 ( .A(n19838), .B(n14678), .Z(n14680) );
  XOR U15078 ( .A(b[15]), .B(a[184]), .Z(n14755) );
  NAND U15079 ( .A(n19805), .B(n14755), .Z(n14679) );
  AND U15080 ( .A(n14680), .B(n14679), .Z(n14762) );
  NAND U15081 ( .A(n35), .B(n14681), .Z(n14683) );
  XOR U15082 ( .A(b[9]), .B(a[190]), .Z(n14758) );
  NAND U15083 ( .A(n19598), .B(n14758), .Z(n14682) );
  NAND U15084 ( .A(n14683), .B(n14682), .Z(n14761) );
  XOR U15085 ( .A(n14762), .B(n14761), .Z(n14764) );
  XOR U15086 ( .A(n14763), .B(n14764), .Z(n14774) );
  NANDN U15087 ( .A(n14685), .B(n14684), .Z(n14689) );
  OR U15088 ( .A(n14687), .B(n14686), .Z(n14688) );
  AND U15089 ( .A(n14689), .B(n14688), .Z(n14773) );
  XNOR U15090 ( .A(n14774), .B(n14773), .Z(n14775) );
  NANDN U15091 ( .A(n14691), .B(n14690), .Z(n14695) );
  NANDN U15092 ( .A(n14693), .B(n14692), .Z(n14694) );
  NAND U15093 ( .A(n14695), .B(n14694), .Z(n14776) );
  XNOR U15094 ( .A(n14775), .B(n14776), .Z(n14721) );
  XOR U15095 ( .A(n14722), .B(n14721), .Z(n14780) );
  NANDN U15096 ( .A(n14697), .B(n14696), .Z(n14701) );
  NANDN U15097 ( .A(n14699), .B(n14698), .Z(n14700) );
  AND U15098 ( .A(n14701), .B(n14700), .Z(n14779) );
  XNOR U15099 ( .A(n14780), .B(n14779), .Z(n14781) );
  XOR U15100 ( .A(n14782), .B(n14781), .Z(n14714) );
  NANDN U15101 ( .A(n14703), .B(n14702), .Z(n14707) );
  NAND U15102 ( .A(n14705), .B(n14704), .Z(n14706) );
  AND U15103 ( .A(n14707), .B(n14706), .Z(n14713) );
  XNOR U15104 ( .A(n14714), .B(n14713), .Z(n14715) );
  XNOR U15105 ( .A(n14716), .B(n14715), .Z(n14785) );
  XNOR U15106 ( .A(sreg[438]), .B(n14785), .Z(n14787) );
  NANDN U15107 ( .A(sreg[437]), .B(n14708), .Z(n14712) );
  NAND U15108 ( .A(n14710), .B(n14709), .Z(n14711) );
  NAND U15109 ( .A(n14712), .B(n14711), .Z(n14786) );
  XNOR U15110 ( .A(n14787), .B(n14786), .Z(c[438]) );
  NANDN U15111 ( .A(n14714), .B(n14713), .Z(n14718) );
  NANDN U15112 ( .A(n14716), .B(n14715), .Z(n14717) );
  AND U15113 ( .A(n14718), .B(n14717), .Z(n14793) );
  NANDN U15114 ( .A(n14720), .B(n14719), .Z(n14724) );
  NAND U15115 ( .A(n14722), .B(n14721), .Z(n14723) );
  AND U15116 ( .A(n14724), .B(n14723), .Z(n14859) );
  NANDN U15117 ( .A(n14726), .B(n14725), .Z(n14730) );
  NANDN U15118 ( .A(n14728), .B(n14727), .Z(n14729) );
  AND U15119 ( .A(n14730), .B(n14729), .Z(n14825) );
  NAND U15120 ( .A(b[0]), .B(a[199]), .Z(n14731) );
  XNOR U15121 ( .A(b[1]), .B(n14731), .Z(n14733) );
  NANDN U15122 ( .A(b[0]), .B(a[198]), .Z(n14732) );
  NAND U15123 ( .A(n14733), .B(n14732), .Z(n14805) );
  NAND U15124 ( .A(n19808), .B(n14734), .Z(n14736) );
  XOR U15125 ( .A(b[13]), .B(a[187]), .Z(n14808) );
  NAND U15126 ( .A(n19768), .B(n14808), .Z(n14735) );
  AND U15127 ( .A(n14736), .B(n14735), .Z(n14803) );
  AND U15128 ( .A(b[15]), .B(a[183]), .Z(n14802) );
  XNOR U15129 ( .A(n14803), .B(n14802), .Z(n14804) );
  XNOR U15130 ( .A(n14805), .B(n14804), .Z(n14823) );
  NAND U15131 ( .A(n33), .B(n14737), .Z(n14739) );
  XOR U15132 ( .A(b[5]), .B(a[195]), .Z(n14814) );
  NAND U15133 ( .A(n19342), .B(n14814), .Z(n14738) );
  AND U15134 ( .A(n14739), .B(n14738), .Z(n14847) );
  NAND U15135 ( .A(n34), .B(n14740), .Z(n14742) );
  XOR U15136 ( .A(b[7]), .B(a[193]), .Z(n14817) );
  NAND U15137 ( .A(n19486), .B(n14817), .Z(n14741) );
  AND U15138 ( .A(n14742), .B(n14741), .Z(n14845) );
  NAND U15139 ( .A(n31), .B(n14743), .Z(n14745) );
  XOR U15140 ( .A(b[3]), .B(a[197]), .Z(n14820) );
  NAND U15141 ( .A(n32), .B(n14820), .Z(n14744) );
  NAND U15142 ( .A(n14745), .B(n14744), .Z(n14844) );
  XNOR U15143 ( .A(n14845), .B(n14844), .Z(n14846) );
  XOR U15144 ( .A(n14847), .B(n14846), .Z(n14824) );
  XOR U15145 ( .A(n14823), .B(n14824), .Z(n14826) );
  XOR U15146 ( .A(n14825), .B(n14826), .Z(n14797) );
  NANDN U15147 ( .A(n14747), .B(n14746), .Z(n14751) );
  OR U15148 ( .A(n14749), .B(n14748), .Z(n14750) );
  AND U15149 ( .A(n14751), .B(n14750), .Z(n14796) );
  XNOR U15150 ( .A(n14797), .B(n14796), .Z(n14799) );
  NAND U15151 ( .A(n14752), .B(n19724), .Z(n14754) );
  XOR U15152 ( .A(b[11]), .B(a[189]), .Z(n14829) );
  NAND U15153 ( .A(n19692), .B(n14829), .Z(n14753) );
  AND U15154 ( .A(n14754), .B(n14753), .Z(n14840) );
  NAND U15155 ( .A(n19838), .B(n14755), .Z(n14757) );
  XOR U15156 ( .A(b[15]), .B(a[185]), .Z(n14832) );
  NAND U15157 ( .A(n19805), .B(n14832), .Z(n14756) );
  AND U15158 ( .A(n14757), .B(n14756), .Z(n14839) );
  NAND U15159 ( .A(n35), .B(n14758), .Z(n14760) );
  XOR U15160 ( .A(b[9]), .B(a[191]), .Z(n14835) );
  NAND U15161 ( .A(n19598), .B(n14835), .Z(n14759) );
  NAND U15162 ( .A(n14760), .B(n14759), .Z(n14838) );
  XOR U15163 ( .A(n14839), .B(n14838), .Z(n14841) );
  XOR U15164 ( .A(n14840), .B(n14841), .Z(n14851) );
  NANDN U15165 ( .A(n14762), .B(n14761), .Z(n14766) );
  OR U15166 ( .A(n14764), .B(n14763), .Z(n14765) );
  AND U15167 ( .A(n14766), .B(n14765), .Z(n14850) );
  XNOR U15168 ( .A(n14851), .B(n14850), .Z(n14852) );
  NANDN U15169 ( .A(n14768), .B(n14767), .Z(n14772) );
  NANDN U15170 ( .A(n14770), .B(n14769), .Z(n14771) );
  NAND U15171 ( .A(n14772), .B(n14771), .Z(n14853) );
  XNOR U15172 ( .A(n14852), .B(n14853), .Z(n14798) );
  XOR U15173 ( .A(n14799), .B(n14798), .Z(n14857) );
  NANDN U15174 ( .A(n14774), .B(n14773), .Z(n14778) );
  NANDN U15175 ( .A(n14776), .B(n14775), .Z(n14777) );
  AND U15176 ( .A(n14778), .B(n14777), .Z(n14856) );
  XNOR U15177 ( .A(n14857), .B(n14856), .Z(n14858) );
  XOR U15178 ( .A(n14859), .B(n14858), .Z(n14791) );
  NANDN U15179 ( .A(n14780), .B(n14779), .Z(n14784) );
  NAND U15180 ( .A(n14782), .B(n14781), .Z(n14783) );
  AND U15181 ( .A(n14784), .B(n14783), .Z(n14790) );
  XNOR U15182 ( .A(n14791), .B(n14790), .Z(n14792) );
  XNOR U15183 ( .A(n14793), .B(n14792), .Z(n14862) );
  XNOR U15184 ( .A(sreg[439]), .B(n14862), .Z(n14864) );
  NANDN U15185 ( .A(sreg[438]), .B(n14785), .Z(n14789) );
  NAND U15186 ( .A(n14787), .B(n14786), .Z(n14788) );
  NAND U15187 ( .A(n14789), .B(n14788), .Z(n14863) );
  XNOR U15188 ( .A(n14864), .B(n14863), .Z(c[439]) );
  NANDN U15189 ( .A(n14791), .B(n14790), .Z(n14795) );
  NANDN U15190 ( .A(n14793), .B(n14792), .Z(n14794) );
  AND U15191 ( .A(n14795), .B(n14794), .Z(n14870) );
  NANDN U15192 ( .A(n14797), .B(n14796), .Z(n14801) );
  NAND U15193 ( .A(n14799), .B(n14798), .Z(n14800) );
  AND U15194 ( .A(n14801), .B(n14800), .Z(n14936) );
  NANDN U15195 ( .A(n14803), .B(n14802), .Z(n14807) );
  NANDN U15196 ( .A(n14805), .B(n14804), .Z(n14806) );
  AND U15197 ( .A(n14807), .B(n14806), .Z(n14923) );
  NAND U15198 ( .A(n19808), .B(n14808), .Z(n14810) );
  XOR U15199 ( .A(b[13]), .B(a[188]), .Z(n14909) );
  NAND U15200 ( .A(n19768), .B(n14909), .Z(n14809) );
  AND U15201 ( .A(n14810), .B(n14809), .Z(n14901) );
  AND U15202 ( .A(b[15]), .B(a[184]), .Z(n14900) );
  XNOR U15203 ( .A(n14901), .B(n14900), .Z(n14902) );
  NAND U15204 ( .A(b[0]), .B(a[200]), .Z(n14811) );
  XNOR U15205 ( .A(b[1]), .B(n14811), .Z(n14813) );
  NANDN U15206 ( .A(b[0]), .B(a[199]), .Z(n14812) );
  NAND U15207 ( .A(n14813), .B(n14812), .Z(n14903) );
  XNOR U15208 ( .A(n14902), .B(n14903), .Z(n14921) );
  NAND U15209 ( .A(n33), .B(n14814), .Z(n14816) );
  XOR U15210 ( .A(b[5]), .B(a[196]), .Z(n14912) );
  NAND U15211 ( .A(n19342), .B(n14912), .Z(n14815) );
  AND U15212 ( .A(n14816), .B(n14815), .Z(n14897) );
  NAND U15213 ( .A(n34), .B(n14817), .Z(n14819) );
  XOR U15214 ( .A(b[7]), .B(a[194]), .Z(n14915) );
  NAND U15215 ( .A(n19486), .B(n14915), .Z(n14818) );
  AND U15216 ( .A(n14819), .B(n14818), .Z(n14895) );
  NAND U15217 ( .A(n31), .B(n14820), .Z(n14822) );
  XOR U15218 ( .A(b[3]), .B(a[198]), .Z(n14918) );
  NAND U15219 ( .A(n32), .B(n14918), .Z(n14821) );
  NAND U15220 ( .A(n14822), .B(n14821), .Z(n14894) );
  XNOR U15221 ( .A(n14895), .B(n14894), .Z(n14896) );
  XOR U15222 ( .A(n14897), .B(n14896), .Z(n14922) );
  XOR U15223 ( .A(n14921), .B(n14922), .Z(n14924) );
  XOR U15224 ( .A(n14923), .B(n14924), .Z(n14874) );
  NANDN U15225 ( .A(n14824), .B(n14823), .Z(n14828) );
  OR U15226 ( .A(n14826), .B(n14825), .Z(n14827) );
  AND U15227 ( .A(n14828), .B(n14827), .Z(n14873) );
  XNOR U15228 ( .A(n14874), .B(n14873), .Z(n14876) );
  NAND U15229 ( .A(n14829), .B(n19724), .Z(n14831) );
  XOR U15230 ( .A(b[11]), .B(a[190]), .Z(n14879) );
  NAND U15231 ( .A(n19692), .B(n14879), .Z(n14830) );
  AND U15232 ( .A(n14831), .B(n14830), .Z(n14890) );
  NAND U15233 ( .A(n19838), .B(n14832), .Z(n14834) );
  XOR U15234 ( .A(b[15]), .B(a[186]), .Z(n14882) );
  NAND U15235 ( .A(n19805), .B(n14882), .Z(n14833) );
  AND U15236 ( .A(n14834), .B(n14833), .Z(n14889) );
  NAND U15237 ( .A(n35), .B(n14835), .Z(n14837) );
  XOR U15238 ( .A(b[9]), .B(a[192]), .Z(n14885) );
  NAND U15239 ( .A(n19598), .B(n14885), .Z(n14836) );
  NAND U15240 ( .A(n14837), .B(n14836), .Z(n14888) );
  XOR U15241 ( .A(n14889), .B(n14888), .Z(n14891) );
  XOR U15242 ( .A(n14890), .B(n14891), .Z(n14928) );
  NANDN U15243 ( .A(n14839), .B(n14838), .Z(n14843) );
  OR U15244 ( .A(n14841), .B(n14840), .Z(n14842) );
  AND U15245 ( .A(n14843), .B(n14842), .Z(n14927) );
  XNOR U15246 ( .A(n14928), .B(n14927), .Z(n14929) );
  NANDN U15247 ( .A(n14845), .B(n14844), .Z(n14849) );
  NANDN U15248 ( .A(n14847), .B(n14846), .Z(n14848) );
  NAND U15249 ( .A(n14849), .B(n14848), .Z(n14930) );
  XNOR U15250 ( .A(n14929), .B(n14930), .Z(n14875) );
  XOR U15251 ( .A(n14876), .B(n14875), .Z(n14934) );
  NANDN U15252 ( .A(n14851), .B(n14850), .Z(n14855) );
  NANDN U15253 ( .A(n14853), .B(n14852), .Z(n14854) );
  AND U15254 ( .A(n14855), .B(n14854), .Z(n14933) );
  XNOR U15255 ( .A(n14934), .B(n14933), .Z(n14935) );
  XOR U15256 ( .A(n14936), .B(n14935), .Z(n14868) );
  NANDN U15257 ( .A(n14857), .B(n14856), .Z(n14861) );
  NAND U15258 ( .A(n14859), .B(n14858), .Z(n14860) );
  AND U15259 ( .A(n14861), .B(n14860), .Z(n14867) );
  XNOR U15260 ( .A(n14868), .B(n14867), .Z(n14869) );
  XNOR U15261 ( .A(n14870), .B(n14869), .Z(n14939) );
  XNOR U15262 ( .A(sreg[440]), .B(n14939), .Z(n14941) );
  NANDN U15263 ( .A(sreg[439]), .B(n14862), .Z(n14866) );
  NAND U15264 ( .A(n14864), .B(n14863), .Z(n14865) );
  NAND U15265 ( .A(n14866), .B(n14865), .Z(n14940) );
  XNOR U15266 ( .A(n14941), .B(n14940), .Z(c[440]) );
  NANDN U15267 ( .A(n14868), .B(n14867), .Z(n14872) );
  NANDN U15268 ( .A(n14870), .B(n14869), .Z(n14871) );
  AND U15269 ( .A(n14872), .B(n14871), .Z(n14947) );
  NANDN U15270 ( .A(n14874), .B(n14873), .Z(n14878) );
  NAND U15271 ( .A(n14876), .B(n14875), .Z(n14877) );
  AND U15272 ( .A(n14878), .B(n14877), .Z(n15013) );
  NAND U15273 ( .A(n14879), .B(n19724), .Z(n14881) );
  XOR U15274 ( .A(b[11]), .B(a[191]), .Z(n14983) );
  NAND U15275 ( .A(n19692), .B(n14983), .Z(n14880) );
  AND U15276 ( .A(n14881), .B(n14880), .Z(n14994) );
  NAND U15277 ( .A(n19838), .B(n14882), .Z(n14884) );
  XOR U15278 ( .A(b[15]), .B(a[187]), .Z(n14986) );
  NAND U15279 ( .A(n19805), .B(n14986), .Z(n14883) );
  AND U15280 ( .A(n14884), .B(n14883), .Z(n14993) );
  NAND U15281 ( .A(n35), .B(n14885), .Z(n14887) );
  XOR U15282 ( .A(b[9]), .B(a[193]), .Z(n14989) );
  NAND U15283 ( .A(n19598), .B(n14989), .Z(n14886) );
  NAND U15284 ( .A(n14887), .B(n14886), .Z(n14992) );
  XOR U15285 ( .A(n14993), .B(n14992), .Z(n14995) );
  XOR U15286 ( .A(n14994), .B(n14995), .Z(n15005) );
  NANDN U15287 ( .A(n14889), .B(n14888), .Z(n14893) );
  OR U15288 ( .A(n14891), .B(n14890), .Z(n14892) );
  AND U15289 ( .A(n14893), .B(n14892), .Z(n15004) );
  XNOR U15290 ( .A(n15005), .B(n15004), .Z(n15006) );
  NANDN U15291 ( .A(n14895), .B(n14894), .Z(n14899) );
  NANDN U15292 ( .A(n14897), .B(n14896), .Z(n14898) );
  NAND U15293 ( .A(n14899), .B(n14898), .Z(n15007) );
  XNOR U15294 ( .A(n15006), .B(n15007), .Z(n14953) );
  NANDN U15295 ( .A(n14901), .B(n14900), .Z(n14905) );
  NANDN U15296 ( .A(n14903), .B(n14902), .Z(n14904) );
  AND U15297 ( .A(n14905), .B(n14904), .Z(n14979) );
  NAND U15298 ( .A(b[0]), .B(a[201]), .Z(n14906) );
  XNOR U15299 ( .A(b[1]), .B(n14906), .Z(n14908) );
  NANDN U15300 ( .A(b[0]), .B(a[200]), .Z(n14907) );
  NAND U15301 ( .A(n14908), .B(n14907), .Z(n14959) );
  NAND U15302 ( .A(n19808), .B(n14909), .Z(n14911) );
  XOR U15303 ( .A(b[13]), .B(a[189]), .Z(n14965) );
  NAND U15304 ( .A(n19768), .B(n14965), .Z(n14910) );
  AND U15305 ( .A(n14911), .B(n14910), .Z(n14957) );
  AND U15306 ( .A(b[15]), .B(a[185]), .Z(n14956) );
  XNOR U15307 ( .A(n14957), .B(n14956), .Z(n14958) );
  XNOR U15308 ( .A(n14959), .B(n14958), .Z(n14977) );
  NAND U15309 ( .A(n33), .B(n14912), .Z(n14914) );
  XOR U15310 ( .A(b[5]), .B(a[197]), .Z(n14968) );
  NAND U15311 ( .A(n19342), .B(n14968), .Z(n14913) );
  AND U15312 ( .A(n14914), .B(n14913), .Z(n15001) );
  NAND U15313 ( .A(n34), .B(n14915), .Z(n14917) );
  XOR U15314 ( .A(b[7]), .B(a[195]), .Z(n14971) );
  NAND U15315 ( .A(n19486), .B(n14971), .Z(n14916) );
  AND U15316 ( .A(n14917), .B(n14916), .Z(n14999) );
  NAND U15317 ( .A(n31), .B(n14918), .Z(n14920) );
  XOR U15318 ( .A(b[3]), .B(a[199]), .Z(n14974) );
  NAND U15319 ( .A(n32), .B(n14974), .Z(n14919) );
  NAND U15320 ( .A(n14920), .B(n14919), .Z(n14998) );
  XNOR U15321 ( .A(n14999), .B(n14998), .Z(n15000) );
  XOR U15322 ( .A(n15001), .B(n15000), .Z(n14978) );
  XOR U15323 ( .A(n14977), .B(n14978), .Z(n14980) );
  XOR U15324 ( .A(n14979), .B(n14980), .Z(n14951) );
  NANDN U15325 ( .A(n14922), .B(n14921), .Z(n14926) );
  OR U15326 ( .A(n14924), .B(n14923), .Z(n14925) );
  AND U15327 ( .A(n14926), .B(n14925), .Z(n14950) );
  XNOR U15328 ( .A(n14951), .B(n14950), .Z(n14952) );
  XOR U15329 ( .A(n14953), .B(n14952), .Z(n15011) );
  NANDN U15330 ( .A(n14928), .B(n14927), .Z(n14932) );
  NANDN U15331 ( .A(n14930), .B(n14929), .Z(n14931) );
  AND U15332 ( .A(n14932), .B(n14931), .Z(n15010) );
  XNOR U15333 ( .A(n15011), .B(n15010), .Z(n15012) );
  XOR U15334 ( .A(n15013), .B(n15012), .Z(n14945) );
  NANDN U15335 ( .A(n14934), .B(n14933), .Z(n14938) );
  NAND U15336 ( .A(n14936), .B(n14935), .Z(n14937) );
  AND U15337 ( .A(n14938), .B(n14937), .Z(n14944) );
  XNOR U15338 ( .A(n14945), .B(n14944), .Z(n14946) );
  XNOR U15339 ( .A(n14947), .B(n14946), .Z(n15016) );
  XNOR U15340 ( .A(sreg[441]), .B(n15016), .Z(n15018) );
  NANDN U15341 ( .A(sreg[440]), .B(n14939), .Z(n14943) );
  NAND U15342 ( .A(n14941), .B(n14940), .Z(n14942) );
  NAND U15343 ( .A(n14943), .B(n14942), .Z(n15017) );
  XNOR U15344 ( .A(n15018), .B(n15017), .Z(c[441]) );
  NANDN U15345 ( .A(n14945), .B(n14944), .Z(n14949) );
  NANDN U15346 ( .A(n14947), .B(n14946), .Z(n14948) );
  AND U15347 ( .A(n14949), .B(n14948), .Z(n15024) );
  NANDN U15348 ( .A(n14951), .B(n14950), .Z(n14955) );
  NAND U15349 ( .A(n14953), .B(n14952), .Z(n14954) );
  AND U15350 ( .A(n14955), .B(n14954), .Z(n15090) );
  NANDN U15351 ( .A(n14957), .B(n14956), .Z(n14961) );
  NANDN U15352 ( .A(n14959), .B(n14958), .Z(n14960) );
  AND U15353 ( .A(n14961), .B(n14960), .Z(n15056) );
  NAND U15354 ( .A(b[0]), .B(a[202]), .Z(n14962) );
  XNOR U15355 ( .A(b[1]), .B(n14962), .Z(n14964) );
  NANDN U15356 ( .A(b[0]), .B(a[201]), .Z(n14963) );
  NAND U15357 ( .A(n14964), .B(n14963), .Z(n15036) );
  NAND U15358 ( .A(n19808), .B(n14965), .Z(n14967) );
  XOR U15359 ( .A(b[13]), .B(a[190]), .Z(n15039) );
  NAND U15360 ( .A(n19768), .B(n15039), .Z(n14966) );
  AND U15361 ( .A(n14967), .B(n14966), .Z(n15034) );
  AND U15362 ( .A(b[15]), .B(a[186]), .Z(n15033) );
  XNOR U15363 ( .A(n15034), .B(n15033), .Z(n15035) );
  XNOR U15364 ( .A(n15036), .B(n15035), .Z(n15054) );
  NAND U15365 ( .A(n33), .B(n14968), .Z(n14970) );
  XOR U15366 ( .A(b[5]), .B(a[198]), .Z(n15045) );
  NAND U15367 ( .A(n19342), .B(n15045), .Z(n14969) );
  AND U15368 ( .A(n14970), .B(n14969), .Z(n15078) );
  NAND U15369 ( .A(n34), .B(n14971), .Z(n14973) );
  XOR U15370 ( .A(b[7]), .B(a[196]), .Z(n15048) );
  NAND U15371 ( .A(n19486), .B(n15048), .Z(n14972) );
  AND U15372 ( .A(n14973), .B(n14972), .Z(n15076) );
  NAND U15373 ( .A(n31), .B(n14974), .Z(n14976) );
  XOR U15374 ( .A(b[3]), .B(a[200]), .Z(n15051) );
  NAND U15375 ( .A(n32), .B(n15051), .Z(n14975) );
  NAND U15376 ( .A(n14976), .B(n14975), .Z(n15075) );
  XNOR U15377 ( .A(n15076), .B(n15075), .Z(n15077) );
  XOR U15378 ( .A(n15078), .B(n15077), .Z(n15055) );
  XOR U15379 ( .A(n15054), .B(n15055), .Z(n15057) );
  XOR U15380 ( .A(n15056), .B(n15057), .Z(n15028) );
  NANDN U15381 ( .A(n14978), .B(n14977), .Z(n14982) );
  OR U15382 ( .A(n14980), .B(n14979), .Z(n14981) );
  AND U15383 ( .A(n14982), .B(n14981), .Z(n15027) );
  XNOR U15384 ( .A(n15028), .B(n15027), .Z(n15030) );
  NAND U15385 ( .A(n14983), .B(n19724), .Z(n14985) );
  XOR U15386 ( .A(b[11]), .B(a[192]), .Z(n15060) );
  NAND U15387 ( .A(n19692), .B(n15060), .Z(n14984) );
  AND U15388 ( .A(n14985), .B(n14984), .Z(n15071) );
  NAND U15389 ( .A(n19838), .B(n14986), .Z(n14988) );
  XOR U15390 ( .A(b[15]), .B(a[188]), .Z(n15063) );
  NAND U15391 ( .A(n19805), .B(n15063), .Z(n14987) );
  AND U15392 ( .A(n14988), .B(n14987), .Z(n15070) );
  NAND U15393 ( .A(n35), .B(n14989), .Z(n14991) );
  XOR U15394 ( .A(b[9]), .B(a[194]), .Z(n15066) );
  NAND U15395 ( .A(n19598), .B(n15066), .Z(n14990) );
  NAND U15396 ( .A(n14991), .B(n14990), .Z(n15069) );
  XOR U15397 ( .A(n15070), .B(n15069), .Z(n15072) );
  XOR U15398 ( .A(n15071), .B(n15072), .Z(n15082) );
  NANDN U15399 ( .A(n14993), .B(n14992), .Z(n14997) );
  OR U15400 ( .A(n14995), .B(n14994), .Z(n14996) );
  AND U15401 ( .A(n14997), .B(n14996), .Z(n15081) );
  XNOR U15402 ( .A(n15082), .B(n15081), .Z(n15083) );
  NANDN U15403 ( .A(n14999), .B(n14998), .Z(n15003) );
  NANDN U15404 ( .A(n15001), .B(n15000), .Z(n15002) );
  NAND U15405 ( .A(n15003), .B(n15002), .Z(n15084) );
  XNOR U15406 ( .A(n15083), .B(n15084), .Z(n15029) );
  XOR U15407 ( .A(n15030), .B(n15029), .Z(n15088) );
  NANDN U15408 ( .A(n15005), .B(n15004), .Z(n15009) );
  NANDN U15409 ( .A(n15007), .B(n15006), .Z(n15008) );
  AND U15410 ( .A(n15009), .B(n15008), .Z(n15087) );
  XNOR U15411 ( .A(n15088), .B(n15087), .Z(n15089) );
  XOR U15412 ( .A(n15090), .B(n15089), .Z(n15022) );
  NANDN U15413 ( .A(n15011), .B(n15010), .Z(n15015) );
  NAND U15414 ( .A(n15013), .B(n15012), .Z(n15014) );
  AND U15415 ( .A(n15015), .B(n15014), .Z(n15021) );
  XNOR U15416 ( .A(n15022), .B(n15021), .Z(n15023) );
  XNOR U15417 ( .A(n15024), .B(n15023), .Z(n15093) );
  XNOR U15418 ( .A(sreg[442]), .B(n15093), .Z(n15095) );
  NANDN U15419 ( .A(sreg[441]), .B(n15016), .Z(n15020) );
  NAND U15420 ( .A(n15018), .B(n15017), .Z(n15019) );
  NAND U15421 ( .A(n15020), .B(n15019), .Z(n15094) );
  XNOR U15422 ( .A(n15095), .B(n15094), .Z(c[442]) );
  NANDN U15423 ( .A(n15022), .B(n15021), .Z(n15026) );
  NANDN U15424 ( .A(n15024), .B(n15023), .Z(n15025) );
  AND U15425 ( .A(n15026), .B(n15025), .Z(n15101) );
  NANDN U15426 ( .A(n15028), .B(n15027), .Z(n15032) );
  NAND U15427 ( .A(n15030), .B(n15029), .Z(n15031) );
  AND U15428 ( .A(n15032), .B(n15031), .Z(n15167) );
  NANDN U15429 ( .A(n15034), .B(n15033), .Z(n15038) );
  NANDN U15430 ( .A(n15036), .B(n15035), .Z(n15037) );
  AND U15431 ( .A(n15038), .B(n15037), .Z(n15133) );
  NAND U15432 ( .A(n19808), .B(n15039), .Z(n15041) );
  XOR U15433 ( .A(b[13]), .B(a[191]), .Z(n15119) );
  NAND U15434 ( .A(n19768), .B(n15119), .Z(n15040) );
  AND U15435 ( .A(n15041), .B(n15040), .Z(n15111) );
  AND U15436 ( .A(b[15]), .B(a[187]), .Z(n15110) );
  XNOR U15437 ( .A(n15111), .B(n15110), .Z(n15112) );
  NAND U15438 ( .A(b[0]), .B(a[203]), .Z(n15042) );
  XNOR U15439 ( .A(b[1]), .B(n15042), .Z(n15044) );
  NANDN U15440 ( .A(b[0]), .B(a[202]), .Z(n15043) );
  NAND U15441 ( .A(n15044), .B(n15043), .Z(n15113) );
  XNOR U15442 ( .A(n15112), .B(n15113), .Z(n15131) );
  NAND U15443 ( .A(n33), .B(n15045), .Z(n15047) );
  XOR U15444 ( .A(b[5]), .B(a[199]), .Z(n15122) );
  NAND U15445 ( .A(n19342), .B(n15122), .Z(n15046) );
  AND U15446 ( .A(n15047), .B(n15046), .Z(n15155) );
  NAND U15447 ( .A(n34), .B(n15048), .Z(n15050) );
  XOR U15448 ( .A(b[7]), .B(a[197]), .Z(n15125) );
  NAND U15449 ( .A(n19486), .B(n15125), .Z(n15049) );
  AND U15450 ( .A(n15050), .B(n15049), .Z(n15153) );
  NAND U15451 ( .A(n31), .B(n15051), .Z(n15053) );
  XOR U15452 ( .A(b[3]), .B(a[201]), .Z(n15128) );
  NAND U15453 ( .A(n32), .B(n15128), .Z(n15052) );
  NAND U15454 ( .A(n15053), .B(n15052), .Z(n15152) );
  XNOR U15455 ( .A(n15153), .B(n15152), .Z(n15154) );
  XOR U15456 ( .A(n15155), .B(n15154), .Z(n15132) );
  XOR U15457 ( .A(n15131), .B(n15132), .Z(n15134) );
  XOR U15458 ( .A(n15133), .B(n15134), .Z(n15105) );
  NANDN U15459 ( .A(n15055), .B(n15054), .Z(n15059) );
  OR U15460 ( .A(n15057), .B(n15056), .Z(n15058) );
  AND U15461 ( .A(n15059), .B(n15058), .Z(n15104) );
  XNOR U15462 ( .A(n15105), .B(n15104), .Z(n15107) );
  NAND U15463 ( .A(n15060), .B(n19724), .Z(n15062) );
  XOR U15464 ( .A(b[11]), .B(a[193]), .Z(n15137) );
  NAND U15465 ( .A(n19692), .B(n15137), .Z(n15061) );
  AND U15466 ( .A(n15062), .B(n15061), .Z(n15148) );
  NAND U15467 ( .A(n19838), .B(n15063), .Z(n15065) );
  XOR U15468 ( .A(b[15]), .B(a[189]), .Z(n15140) );
  NAND U15469 ( .A(n19805), .B(n15140), .Z(n15064) );
  AND U15470 ( .A(n15065), .B(n15064), .Z(n15147) );
  NAND U15471 ( .A(n35), .B(n15066), .Z(n15068) );
  XOR U15472 ( .A(b[9]), .B(a[195]), .Z(n15143) );
  NAND U15473 ( .A(n19598), .B(n15143), .Z(n15067) );
  NAND U15474 ( .A(n15068), .B(n15067), .Z(n15146) );
  XOR U15475 ( .A(n15147), .B(n15146), .Z(n15149) );
  XOR U15476 ( .A(n15148), .B(n15149), .Z(n15159) );
  NANDN U15477 ( .A(n15070), .B(n15069), .Z(n15074) );
  OR U15478 ( .A(n15072), .B(n15071), .Z(n15073) );
  AND U15479 ( .A(n15074), .B(n15073), .Z(n15158) );
  XNOR U15480 ( .A(n15159), .B(n15158), .Z(n15160) );
  NANDN U15481 ( .A(n15076), .B(n15075), .Z(n15080) );
  NANDN U15482 ( .A(n15078), .B(n15077), .Z(n15079) );
  NAND U15483 ( .A(n15080), .B(n15079), .Z(n15161) );
  XNOR U15484 ( .A(n15160), .B(n15161), .Z(n15106) );
  XOR U15485 ( .A(n15107), .B(n15106), .Z(n15165) );
  NANDN U15486 ( .A(n15082), .B(n15081), .Z(n15086) );
  NANDN U15487 ( .A(n15084), .B(n15083), .Z(n15085) );
  AND U15488 ( .A(n15086), .B(n15085), .Z(n15164) );
  XNOR U15489 ( .A(n15165), .B(n15164), .Z(n15166) );
  XOR U15490 ( .A(n15167), .B(n15166), .Z(n15099) );
  NANDN U15491 ( .A(n15088), .B(n15087), .Z(n15092) );
  NAND U15492 ( .A(n15090), .B(n15089), .Z(n15091) );
  AND U15493 ( .A(n15092), .B(n15091), .Z(n15098) );
  XNOR U15494 ( .A(n15099), .B(n15098), .Z(n15100) );
  XNOR U15495 ( .A(n15101), .B(n15100), .Z(n15170) );
  XNOR U15496 ( .A(sreg[443]), .B(n15170), .Z(n15172) );
  NANDN U15497 ( .A(sreg[442]), .B(n15093), .Z(n15097) );
  NAND U15498 ( .A(n15095), .B(n15094), .Z(n15096) );
  NAND U15499 ( .A(n15097), .B(n15096), .Z(n15171) );
  XNOR U15500 ( .A(n15172), .B(n15171), .Z(c[443]) );
  NANDN U15501 ( .A(n15099), .B(n15098), .Z(n15103) );
  NANDN U15502 ( .A(n15101), .B(n15100), .Z(n15102) );
  AND U15503 ( .A(n15103), .B(n15102), .Z(n15178) );
  NANDN U15504 ( .A(n15105), .B(n15104), .Z(n15109) );
  NAND U15505 ( .A(n15107), .B(n15106), .Z(n15108) );
  AND U15506 ( .A(n15109), .B(n15108), .Z(n15244) );
  NANDN U15507 ( .A(n15111), .B(n15110), .Z(n15115) );
  NANDN U15508 ( .A(n15113), .B(n15112), .Z(n15114) );
  AND U15509 ( .A(n15115), .B(n15114), .Z(n15210) );
  NAND U15510 ( .A(b[0]), .B(a[204]), .Z(n15116) );
  XNOR U15511 ( .A(b[1]), .B(n15116), .Z(n15118) );
  NANDN U15512 ( .A(b[0]), .B(a[203]), .Z(n15117) );
  NAND U15513 ( .A(n15118), .B(n15117), .Z(n15190) );
  NAND U15514 ( .A(n19808), .B(n15119), .Z(n15121) );
  XOR U15515 ( .A(b[13]), .B(a[192]), .Z(n15196) );
  NAND U15516 ( .A(n19768), .B(n15196), .Z(n15120) );
  AND U15517 ( .A(n15121), .B(n15120), .Z(n15188) );
  AND U15518 ( .A(b[15]), .B(a[188]), .Z(n15187) );
  XNOR U15519 ( .A(n15188), .B(n15187), .Z(n15189) );
  XNOR U15520 ( .A(n15190), .B(n15189), .Z(n15208) );
  NAND U15521 ( .A(n33), .B(n15122), .Z(n15124) );
  XOR U15522 ( .A(b[5]), .B(a[200]), .Z(n15199) );
  NAND U15523 ( .A(n19342), .B(n15199), .Z(n15123) );
  AND U15524 ( .A(n15124), .B(n15123), .Z(n15232) );
  NAND U15525 ( .A(n34), .B(n15125), .Z(n15127) );
  XOR U15526 ( .A(b[7]), .B(a[198]), .Z(n15202) );
  NAND U15527 ( .A(n19486), .B(n15202), .Z(n15126) );
  AND U15528 ( .A(n15127), .B(n15126), .Z(n15230) );
  NAND U15529 ( .A(n31), .B(n15128), .Z(n15130) );
  XOR U15530 ( .A(b[3]), .B(a[202]), .Z(n15205) );
  NAND U15531 ( .A(n32), .B(n15205), .Z(n15129) );
  NAND U15532 ( .A(n15130), .B(n15129), .Z(n15229) );
  XNOR U15533 ( .A(n15230), .B(n15229), .Z(n15231) );
  XOR U15534 ( .A(n15232), .B(n15231), .Z(n15209) );
  XOR U15535 ( .A(n15208), .B(n15209), .Z(n15211) );
  XOR U15536 ( .A(n15210), .B(n15211), .Z(n15182) );
  NANDN U15537 ( .A(n15132), .B(n15131), .Z(n15136) );
  OR U15538 ( .A(n15134), .B(n15133), .Z(n15135) );
  AND U15539 ( .A(n15136), .B(n15135), .Z(n15181) );
  XNOR U15540 ( .A(n15182), .B(n15181), .Z(n15184) );
  NAND U15541 ( .A(n15137), .B(n19724), .Z(n15139) );
  XOR U15542 ( .A(b[11]), .B(a[194]), .Z(n15214) );
  NAND U15543 ( .A(n19692), .B(n15214), .Z(n15138) );
  AND U15544 ( .A(n15139), .B(n15138), .Z(n15225) );
  NAND U15545 ( .A(n19838), .B(n15140), .Z(n15142) );
  XOR U15546 ( .A(b[15]), .B(a[190]), .Z(n15217) );
  NAND U15547 ( .A(n19805), .B(n15217), .Z(n15141) );
  AND U15548 ( .A(n15142), .B(n15141), .Z(n15224) );
  NAND U15549 ( .A(n35), .B(n15143), .Z(n15145) );
  XOR U15550 ( .A(b[9]), .B(a[196]), .Z(n15220) );
  NAND U15551 ( .A(n19598), .B(n15220), .Z(n15144) );
  NAND U15552 ( .A(n15145), .B(n15144), .Z(n15223) );
  XOR U15553 ( .A(n15224), .B(n15223), .Z(n15226) );
  XOR U15554 ( .A(n15225), .B(n15226), .Z(n15236) );
  NANDN U15555 ( .A(n15147), .B(n15146), .Z(n15151) );
  OR U15556 ( .A(n15149), .B(n15148), .Z(n15150) );
  AND U15557 ( .A(n15151), .B(n15150), .Z(n15235) );
  XNOR U15558 ( .A(n15236), .B(n15235), .Z(n15237) );
  NANDN U15559 ( .A(n15153), .B(n15152), .Z(n15157) );
  NANDN U15560 ( .A(n15155), .B(n15154), .Z(n15156) );
  NAND U15561 ( .A(n15157), .B(n15156), .Z(n15238) );
  XNOR U15562 ( .A(n15237), .B(n15238), .Z(n15183) );
  XOR U15563 ( .A(n15184), .B(n15183), .Z(n15242) );
  NANDN U15564 ( .A(n15159), .B(n15158), .Z(n15163) );
  NANDN U15565 ( .A(n15161), .B(n15160), .Z(n15162) );
  AND U15566 ( .A(n15163), .B(n15162), .Z(n15241) );
  XNOR U15567 ( .A(n15242), .B(n15241), .Z(n15243) );
  XOR U15568 ( .A(n15244), .B(n15243), .Z(n15176) );
  NANDN U15569 ( .A(n15165), .B(n15164), .Z(n15169) );
  NAND U15570 ( .A(n15167), .B(n15166), .Z(n15168) );
  AND U15571 ( .A(n15169), .B(n15168), .Z(n15175) );
  XNOR U15572 ( .A(n15176), .B(n15175), .Z(n15177) );
  XNOR U15573 ( .A(n15178), .B(n15177), .Z(n15247) );
  XNOR U15574 ( .A(sreg[444]), .B(n15247), .Z(n15249) );
  NANDN U15575 ( .A(sreg[443]), .B(n15170), .Z(n15174) );
  NAND U15576 ( .A(n15172), .B(n15171), .Z(n15173) );
  NAND U15577 ( .A(n15174), .B(n15173), .Z(n15248) );
  XNOR U15578 ( .A(n15249), .B(n15248), .Z(c[444]) );
  NANDN U15579 ( .A(n15176), .B(n15175), .Z(n15180) );
  NANDN U15580 ( .A(n15178), .B(n15177), .Z(n15179) );
  AND U15581 ( .A(n15180), .B(n15179), .Z(n15255) );
  NANDN U15582 ( .A(n15182), .B(n15181), .Z(n15186) );
  NAND U15583 ( .A(n15184), .B(n15183), .Z(n15185) );
  AND U15584 ( .A(n15186), .B(n15185), .Z(n15321) );
  NANDN U15585 ( .A(n15188), .B(n15187), .Z(n15192) );
  NANDN U15586 ( .A(n15190), .B(n15189), .Z(n15191) );
  AND U15587 ( .A(n15192), .B(n15191), .Z(n15287) );
  NAND U15588 ( .A(b[0]), .B(a[205]), .Z(n15193) );
  XNOR U15589 ( .A(b[1]), .B(n15193), .Z(n15195) );
  NANDN U15590 ( .A(b[0]), .B(a[204]), .Z(n15194) );
  NAND U15591 ( .A(n15195), .B(n15194), .Z(n15267) );
  NAND U15592 ( .A(n19808), .B(n15196), .Z(n15198) );
  XOR U15593 ( .A(b[13]), .B(a[193]), .Z(n15273) );
  NAND U15594 ( .A(n19768), .B(n15273), .Z(n15197) );
  AND U15595 ( .A(n15198), .B(n15197), .Z(n15265) );
  AND U15596 ( .A(b[15]), .B(a[189]), .Z(n15264) );
  XNOR U15597 ( .A(n15265), .B(n15264), .Z(n15266) );
  XNOR U15598 ( .A(n15267), .B(n15266), .Z(n15285) );
  NAND U15599 ( .A(n33), .B(n15199), .Z(n15201) );
  XOR U15600 ( .A(b[5]), .B(a[201]), .Z(n15276) );
  NAND U15601 ( .A(n19342), .B(n15276), .Z(n15200) );
  AND U15602 ( .A(n15201), .B(n15200), .Z(n15309) );
  NAND U15603 ( .A(n34), .B(n15202), .Z(n15204) );
  XOR U15604 ( .A(b[7]), .B(a[199]), .Z(n15279) );
  NAND U15605 ( .A(n19486), .B(n15279), .Z(n15203) );
  AND U15606 ( .A(n15204), .B(n15203), .Z(n15307) );
  NAND U15607 ( .A(n31), .B(n15205), .Z(n15207) );
  XOR U15608 ( .A(b[3]), .B(a[203]), .Z(n15282) );
  NAND U15609 ( .A(n32), .B(n15282), .Z(n15206) );
  NAND U15610 ( .A(n15207), .B(n15206), .Z(n15306) );
  XNOR U15611 ( .A(n15307), .B(n15306), .Z(n15308) );
  XOR U15612 ( .A(n15309), .B(n15308), .Z(n15286) );
  XOR U15613 ( .A(n15285), .B(n15286), .Z(n15288) );
  XOR U15614 ( .A(n15287), .B(n15288), .Z(n15259) );
  NANDN U15615 ( .A(n15209), .B(n15208), .Z(n15213) );
  OR U15616 ( .A(n15211), .B(n15210), .Z(n15212) );
  AND U15617 ( .A(n15213), .B(n15212), .Z(n15258) );
  XNOR U15618 ( .A(n15259), .B(n15258), .Z(n15261) );
  NAND U15619 ( .A(n15214), .B(n19724), .Z(n15216) );
  XOR U15620 ( .A(b[11]), .B(a[195]), .Z(n15291) );
  NAND U15621 ( .A(n19692), .B(n15291), .Z(n15215) );
  AND U15622 ( .A(n15216), .B(n15215), .Z(n15302) );
  NAND U15623 ( .A(n19838), .B(n15217), .Z(n15219) );
  XOR U15624 ( .A(b[15]), .B(a[191]), .Z(n15294) );
  NAND U15625 ( .A(n19805), .B(n15294), .Z(n15218) );
  AND U15626 ( .A(n15219), .B(n15218), .Z(n15301) );
  NAND U15627 ( .A(n35), .B(n15220), .Z(n15222) );
  XOR U15628 ( .A(b[9]), .B(a[197]), .Z(n15297) );
  NAND U15629 ( .A(n19598), .B(n15297), .Z(n15221) );
  NAND U15630 ( .A(n15222), .B(n15221), .Z(n15300) );
  XOR U15631 ( .A(n15301), .B(n15300), .Z(n15303) );
  XOR U15632 ( .A(n15302), .B(n15303), .Z(n15313) );
  NANDN U15633 ( .A(n15224), .B(n15223), .Z(n15228) );
  OR U15634 ( .A(n15226), .B(n15225), .Z(n15227) );
  AND U15635 ( .A(n15228), .B(n15227), .Z(n15312) );
  XNOR U15636 ( .A(n15313), .B(n15312), .Z(n15314) );
  NANDN U15637 ( .A(n15230), .B(n15229), .Z(n15234) );
  NANDN U15638 ( .A(n15232), .B(n15231), .Z(n15233) );
  NAND U15639 ( .A(n15234), .B(n15233), .Z(n15315) );
  XNOR U15640 ( .A(n15314), .B(n15315), .Z(n15260) );
  XOR U15641 ( .A(n15261), .B(n15260), .Z(n15319) );
  NANDN U15642 ( .A(n15236), .B(n15235), .Z(n15240) );
  NANDN U15643 ( .A(n15238), .B(n15237), .Z(n15239) );
  AND U15644 ( .A(n15240), .B(n15239), .Z(n15318) );
  XNOR U15645 ( .A(n15319), .B(n15318), .Z(n15320) );
  XOR U15646 ( .A(n15321), .B(n15320), .Z(n15253) );
  NANDN U15647 ( .A(n15242), .B(n15241), .Z(n15246) );
  NAND U15648 ( .A(n15244), .B(n15243), .Z(n15245) );
  AND U15649 ( .A(n15246), .B(n15245), .Z(n15252) );
  XNOR U15650 ( .A(n15253), .B(n15252), .Z(n15254) );
  XNOR U15651 ( .A(n15255), .B(n15254), .Z(n15324) );
  XNOR U15652 ( .A(sreg[445]), .B(n15324), .Z(n15326) );
  NANDN U15653 ( .A(sreg[444]), .B(n15247), .Z(n15251) );
  NAND U15654 ( .A(n15249), .B(n15248), .Z(n15250) );
  NAND U15655 ( .A(n15251), .B(n15250), .Z(n15325) );
  XNOR U15656 ( .A(n15326), .B(n15325), .Z(c[445]) );
  NANDN U15657 ( .A(n15253), .B(n15252), .Z(n15257) );
  NANDN U15658 ( .A(n15255), .B(n15254), .Z(n15256) );
  AND U15659 ( .A(n15257), .B(n15256), .Z(n15332) );
  NANDN U15660 ( .A(n15259), .B(n15258), .Z(n15263) );
  NAND U15661 ( .A(n15261), .B(n15260), .Z(n15262) );
  AND U15662 ( .A(n15263), .B(n15262), .Z(n15398) );
  NANDN U15663 ( .A(n15265), .B(n15264), .Z(n15269) );
  NANDN U15664 ( .A(n15267), .B(n15266), .Z(n15268) );
  AND U15665 ( .A(n15269), .B(n15268), .Z(n15364) );
  NAND U15666 ( .A(b[0]), .B(a[206]), .Z(n15270) );
  XNOR U15667 ( .A(b[1]), .B(n15270), .Z(n15272) );
  NANDN U15668 ( .A(b[0]), .B(a[205]), .Z(n15271) );
  NAND U15669 ( .A(n15272), .B(n15271), .Z(n15344) );
  NAND U15670 ( .A(n19808), .B(n15273), .Z(n15275) );
  XOR U15671 ( .A(b[13]), .B(a[194]), .Z(n15350) );
  NAND U15672 ( .A(n19768), .B(n15350), .Z(n15274) );
  AND U15673 ( .A(n15275), .B(n15274), .Z(n15342) );
  AND U15674 ( .A(b[15]), .B(a[190]), .Z(n15341) );
  XNOR U15675 ( .A(n15342), .B(n15341), .Z(n15343) );
  XNOR U15676 ( .A(n15344), .B(n15343), .Z(n15362) );
  NAND U15677 ( .A(n33), .B(n15276), .Z(n15278) );
  XOR U15678 ( .A(b[5]), .B(a[202]), .Z(n15353) );
  NAND U15679 ( .A(n19342), .B(n15353), .Z(n15277) );
  AND U15680 ( .A(n15278), .B(n15277), .Z(n15386) );
  NAND U15681 ( .A(n34), .B(n15279), .Z(n15281) );
  XOR U15682 ( .A(b[7]), .B(a[200]), .Z(n15356) );
  NAND U15683 ( .A(n19486), .B(n15356), .Z(n15280) );
  AND U15684 ( .A(n15281), .B(n15280), .Z(n15384) );
  NAND U15685 ( .A(n31), .B(n15282), .Z(n15284) );
  XOR U15686 ( .A(b[3]), .B(a[204]), .Z(n15359) );
  NAND U15687 ( .A(n32), .B(n15359), .Z(n15283) );
  NAND U15688 ( .A(n15284), .B(n15283), .Z(n15383) );
  XNOR U15689 ( .A(n15384), .B(n15383), .Z(n15385) );
  XOR U15690 ( .A(n15386), .B(n15385), .Z(n15363) );
  XOR U15691 ( .A(n15362), .B(n15363), .Z(n15365) );
  XOR U15692 ( .A(n15364), .B(n15365), .Z(n15336) );
  NANDN U15693 ( .A(n15286), .B(n15285), .Z(n15290) );
  OR U15694 ( .A(n15288), .B(n15287), .Z(n15289) );
  AND U15695 ( .A(n15290), .B(n15289), .Z(n15335) );
  XNOR U15696 ( .A(n15336), .B(n15335), .Z(n15338) );
  NAND U15697 ( .A(n15291), .B(n19724), .Z(n15293) );
  XOR U15698 ( .A(b[11]), .B(a[196]), .Z(n15368) );
  NAND U15699 ( .A(n19692), .B(n15368), .Z(n15292) );
  AND U15700 ( .A(n15293), .B(n15292), .Z(n15379) );
  NAND U15701 ( .A(n19838), .B(n15294), .Z(n15296) );
  XOR U15702 ( .A(b[15]), .B(a[192]), .Z(n15371) );
  NAND U15703 ( .A(n19805), .B(n15371), .Z(n15295) );
  AND U15704 ( .A(n15296), .B(n15295), .Z(n15378) );
  NAND U15705 ( .A(n35), .B(n15297), .Z(n15299) );
  XOR U15706 ( .A(b[9]), .B(a[198]), .Z(n15374) );
  NAND U15707 ( .A(n19598), .B(n15374), .Z(n15298) );
  NAND U15708 ( .A(n15299), .B(n15298), .Z(n15377) );
  XOR U15709 ( .A(n15378), .B(n15377), .Z(n15380) );
  XOR U15710 ( .A(n15379), .B(n15380), .Z(n15390) );
  NANDN U15711 ( .A(n15301), .B(n15300), .Z(n15305) );
  OR U15712 ( .A(n15303), .B(n15302), .Z(n15304) );
  AND U15713 ( .A(n15305), .B(n15304), .Z(n15389) );
  XNOR U15714 ( .A(n15390), .B(n15389), .Z(n15391) );
  NANDN U15715 ( .A(n15307), .B(n15306), .Z(n15311) );
  NANDN U15716 ( .A(n15309), .B(n15308), .Z(n15310) );
  NAND U15717 ( .A(n15311), .B(n15310), .Z(n15392) );
  XNOR U15718 ( .A(n15391), .B(n15392), .Z(n15337) );
  XOR U15719 ( .A(n15338), .B(n15337), .Z(n15396) );
  NANDN U15720 ( .A(n15313), .B(n15312), .Z(n15317) );
  NANDN U15721 ( .A(n15315), .B(n15314), .Z(n15316) );
  AND U15722 ( .A(n15317), .B(n15316), .Z(n15395) );
  XNOR U15723 ( .A(n15396), .B(n15395), .Z(n15397) );
  XOR U15724 ( .A(n15398), .B(n15397), .Z(n15330) );
  NANDN U15725 ( .A(n15319), .B(n15318), .Z(n15323) );
  NAND U15726 ( .A(n15321), .B(n15320), .Z(n15322) );
  AND U15727 ( .A(n15323), .B(n15322), .Z(n15329) );
  XNOR U15728 ( .A(n15330), .B(n15329), .Z(n15331) );
  XNOR U15729 ( .A(n15332), .B(n15331), .Z(n15401) );
  XNOR U15730 ( .A(sreg[446]), .B(n15401), .Z(n15403) );
  NANDN U15731 ( .A(sreg[445]), .B(n15324), .Z(n15328) );
  NAND U15732 ( .A(n15326), .B(n15325), .Z(n15327) );
  NAND U15733 ( .A(n15328), .B(n15327), .Z(n15402) );
  XNOR U15734 ( .A(n15403), .B(n15402), .Z(c[446]) );
  NANDN U15735 ( .A(n15330), .B(n15329), .Z(n15334) );
  NANDN U15736 ( .A(n15332), .B(n15331), .Z(n15333) );
  AND U15737 ( .A(n15334), .B(n15333), .Z(n15409) );
  NANDN U15738 ( .A(n15336), .B(n15335), .Z(n15340) );
  NAND U15739 ( .A(n15338), .B(n15337), .Z(n15339) );
  AND U15740 ( .A(n15340), .B(n15339), .Z(n15475) );
  NANDN U15741 ( .A(n15342), .B(n15341), .Z(n15346) );
  NANDN U15742 ( .A(n15344), .B(n15343), .Z(n15345) );
  AND U15743 ( .A(n15346), .B(n15345), .Z(n15441) );
  NAND U15744 ( .A(b[0]), .B(a[207]), .Z(n15347) );
  XNOR U15745 ( .A(b[1]), .B(n15347), .Z(n15349) );
  NANDN U15746 ( .A(b[0]), .B(a[206]), .Z(n15348) );
  NAND U15747 ( .A(n15349), .B(n15348), .Z(n15421) );
  NAND U15748 ( .A(n19808), .B(n15350), .Z(n15352) );
  XOR U15749 ( .A(b[13]), .B(a[195]), .Z(n15427) );
  NAND U15750 ( .A(n19768), .B(n15427), .Z(n15351) );
  AND U15751 ( .A(n15352), .B(n15351), .Z(n15419) );
  AND U15752 ( .A(b[15]), .B(a[191]), .Z(n15418) );
  XNOR U15753 ( .A(n15419), .B(n15418), .Z(n15420) );
  XNOR U15754 ( .A(n15421), .B(n15420), .Z(n15439) );
  NAND U15755 ( .A(n33), .B(n15353), .Z(n15355) );
  XOR U15756 ( .A(b[5]), .B(a[203]), .Z(n15430) );
  NAND U15757 ( .A(n19342), .B(n15430), .Z(n15354) );
  AND U15758 ( .A(n15355), .B(n15354), .Z(n15463) );
  NAND U15759 ( .A(n34), .B(n15356), .Z(n15358) );
  XOR U15760 ( .A(b[7]), .B(a[201]), .Z(n15433) );
  NAND U15761 ( .A(n19486), .B(n15433), .Z(n15357) );
  AND U15762 ( .A(n15358), .B(n15357), .Z(n15461) );
  NAND U15763 ( .A(n31), .B(n15359), .Z(n15361) );
  XOR U15764 ( .A(b[3]), .B(a[205]), .Z(n15436) );
  NAND U15765 ( .A(n32), .B(n15436), .Z(n15360) );
  NAND U15766 ( .A(n15361), .B(n15360), .Z(n15460) );
  XNOR U15767 ( .A(n15461), .B(n15460), .Z(n15462) );
  XOR U15768 ( .A(n15463), .B(n15462), .Z(n15440) );
  XOR U15769 ( .A(n15439), .B(n15440), .Z(n15442) );
  XOR U15770 ( .A(n15441), .B(n15442), .Z(n15413) );
  NANDN U15771 ( .A(n15363), .B(n15362), .Z(n15367) );
  OR U15772 ( .A(n15365), .B(n15364), .Z(n15366) );
  AND U15773 ( .A(n15367), .B(n15366), .Z(n15412) );
  XNOR U15774 ( .A(n15413), .B(n15412), .Z(n15415) );
  NAND U15775 ( .A(n15368), .B(n19724), .Z(n15370) );
  XOR U15776 ( .A(b[11]), .B(a[197]), .Z(n15445) );
  NAND U15777 ( .A(n19692), .B(n15445), .Z(n15369) );
  AND U15778 ( .A(n15370), .B(n15369), .Z(n15456) );
  NAND U15779 ( .A(n19838), .B(n15371), .Z(n15373) );
  XOR U15780 ( .A(b[15]), .B(a[193]), .Z(n15448) );
  NAND U15781 ( .A(n19805), .B(n15448), .Z(n15372) );
  AND U15782 ( .A(n15373), .B(n15372), .Z(n15455) );
  NAND U15783 ( .A(n35), .B(n15374), .Z(n15376) );
  XOR U15784 ( .A(b[9]), .B(a[199]), .Z(n15451) );
  NAND U15785 ( .A(n19598), .B(n15451), .Z(n15375) );
  NAND U15786 ( .A(n15376), .B(n15375), .Z(n15454) );
  XOR U15787 ( .A(n15455), .B(n15454), .Z(n15457) );
  XOR U15788 ( .A(n15456), .B(n15457), .Z(n15467) );
  NANDN U15789 ( .A(n15378), .B(n15377), .Z(n15382) );
  OR U15790 ( .A(n15380), .B(n15379), .Z(n15381) );
  AND U15791 ( .A(n15382), .B(n15381), .Z(n15466) );
  XNOR U15792 ( .A(n15467), .B(n15466), .Z(n15468) );
  NANDN U15793 ( .A(n15384), .B(n15383), .Z(n15388) );
  NANDN U15794 ( .A(n15386), .B(n15385), .Z(n15387) );
  NAND U15795 ( .A(n15388), .B(n15387), .Z(n15469) );
  XNOR U15796 ( .A(n15468), .B(n15469), .Z(n15414) );
  XOR U15797 ( .A(n15415), .B(n15414), .Z(n15473) );
  NANDN U15798 ( .A(n15390), .B(n15389), .Z(n15394) );
  NANDN U15799 ( .A(n15392), .B(n15391), .Z(n15393) );
  AND U15800 ( .A(n15394), .B(n15393), .Z(n15472) );
  XNOR U15801 ( .A(n15473), .B(n15472), .Z(n15474) );
  XOR U15802 ( .A(n15475), .B(n15474), .Z(n15407) );
  NANDN U15803 ( .A(n15396), .B(n15395), .Z(n15400) );
  NAND U15804 ( .A(n15398), .B(n15397), .Z(n15399) );
  AND U15805 ( .A(n15400), .B(n15399), .Z(n15406) );
  XNOR U15806 ( .A(n15407), .B(n15406), .Z(n15408) );
  XNOR U15807 ( .A(n15409), .B(n15408), .Z(n15478) );
  XNOR U15808 ( .A(sreg[447]), .B(n15478), .Z(n15480) );
  NANDN U15809 ( .A(sreg[446]), .B(n15401), .Z(n15405) );
  NAND U15810 ( .A(n15403), .B(n15402), .Z(n15404) );
  NAND U15811 ( .A(n15405), .B(n15404), .Z(n15479) );
  XNOR U15812 ( .A(n15480), .B(n15479), .Z(c[447]) );
  NANDN U15813 ( .A(n15407), .B(n15406), .Z(n15411) );
  NANDN U15814 ( .A(n15409), .B(n15408), .Z(n15410) );
  AND U15815 ( .A(n15411), .B(n15410), .Z(n15486) );
  NANDN U15816 ( .A(n15413), .B(n15412), .Z(n15417) );
  NAND U15817 ( .A(n15415), .B(n15414), .Z(n15416) );
  AND U15818 ( .A(n15417), .B(n15416), .Z(n15552) );
  NANDN U15819 ( .A(n15419), .B(n15418), .Z(n15423) );
  NANDN U15820 ( .A(n15421), .B(n15420), .Z(n15422) );
  AND U15821 ( .A(n15423), .B(n15422), .Z(n15539) );
  NAND U15822 ( .A(b[0]), .B(a[208]), .Z(n15424) );
  XNOR U15823 ( .A(b[1]), .B(n15424), .Z(n15426) );
  NANDN U15824 ( .A(b[0]), .B(a[207]), .Z(n15425) );
  NAND U15825 ( .A(n15426), .B(n15425), .Z(n15519) );
  NAND U15826 ( .A(n19808), .B(n15427), .Z(n15429) );
  XOR U15827 ( .A(b[13]), .B(a[196]), .Z(n15522) );
  NAND U15828 ( .A(n19768), .B(n15522), .Z(n15428) );
  AND U15829 ( .A(n15429), .B(n15428), .Z(n15517) );
  AND U15830 ( .A(b[15]), .B(a[192]), .Z(n15516) );
  XNOR U15831 ( .A(n15517), .B(n15516), .Z(n15518) );
  XNOR U15832 ( .A(n15519), .B(n15518), .Z(n15537) );
  NAND U15833 ( .A(n33), .B(n15430), .Z(n15432) );
  XOR U15834 ( .A(b[5]), .B(a[204]), .Z(n15528) );
  NAND U15835 ( .A(n19342), .B(n15528), .Z(n15431) );
  AND U15836 ( .A(n15432), .B(n15431), .Z(n15513) );
  NAND U15837 ( .A(n34), .B(n15433), .Z(n15435) );
  XOR U15838 ( .A(b[7]), .B(a[202]), .Z(n15531) );
  NAND U15839 ( .A(n19486), .B(n15531), .Z(n15434) );
  AND U15840 ( .A(n15435), .B(n15434), .Z(n15511) );
  NAND U15841 ( .A(n31), .B(n15436), .Z(n15438) );
  XOR U15842 ( .A(b[3]), .B(a[206]), .Z(n15534) );
  NAND U15843 ( .A(n32), .B(n15534), .Z(n15437) );
  NAND U15844 ( .A(n15438), .B(n15437), .Z(n15510) );
  XNOR U15845 ( .A(n15511), .B(n15510), .Z(n15512) );
  XOR U15846 ( .A(n15513), .B(n15512), .Z(n15538) );
  XOR U15847 ( .A(n15537), .B(n15538), .Z(n15540) );
  XOR U15848 ( .A(n15539), .B(n15540), .Z(n15490) );
  NANDN U15849 ( .A(n15440), .B(n15439), .Z(n15444) );
  OR U15850 ( .A(n15442), .B(n15441), .Z(n15443) );
  AND U15851 ( .A(n15444), .B(n15443), .Z(n15489) );
  XNOR U15852 ( .A(n15490), .B(n15489), .Z(n15492) );
  NAND U15853 ( .A(n15445), .B(n19724), .Z(n15447) );
  XOR U15854 ( .A(b[11]), .B(a[198]), .Z(n15495) );
  NAND U15855 ( .A(n19692), .B(n15495), .Z(n15446) );
  AND U15856 ( .A(n15447), .B(n15446), .Z(n15506) );
  NAND U15857 ( .A(n19838), .B(n15448), .Z(n15450) );
  XOR U15858 ( .A(b[15]), .B(a[194]), .Z(n15498) );
  NAND U15859 ( .A(n19805), .B(n15498), .Z(n15449) );
  AND U15860 ( .A(n15450), .B(n15449), .Z(n15505) );
  NAND U15861 ( .A(n35), .B(n15451), .Z(n15453) );
  XOR U15862 ( .A(b[9]), .B(a[200]), .Z(n15501) );
  NAND U15863 ( .A(n19598), .B(n15501), .Z(n15452) );
  NAND U15864 ( .A(n15453), .B(n15452), .Z(n15504) );
  XOR U15865 ( .A(n15505), .B(n15504), .Z(n15507) );
  XOR U15866 ( .A(n15506), .B(n15507), .Z(n15544) );
  NANDN U15867 ( .A(n15455), .B(n15454), .Z(n15459) );
  OR U15868 ( .A(n15457), .B(n15456), .Z(n15458) );
  AND U15869 ( .A(n15459), .B(n15458), .Z(n15543) );
  XNOR U15870 ( .A(n15544), .B(n15543), .Z(n15545) );
  NANDN U15871 ( .A(n15461), .B(n15460), .Z(n15465) );
  NANDN U15872 ( .A(n15463), .B(n15462), .Z(n15464) );
  NAND U15873 ( .A(n15465), .B(n15464), .Z(n15546) );
  XNOR U15874 ( .A(n15545), .B(n15546), .Z(n15491) );
  XOR U15875 ( .A(n15492), .B(n15491), .Z(n15550) );
  NANDN U15876 ( .A(n15467), .B(n15466), .Z(n15471) );
  NANDN U15877 ( .A(n15469), .B(n15468), .Z(n15470) );
  AND U15878 ( .A(n15471), .B(n15470), .Z(n15549) );
  XNOR U15879 ( .A(n15550), .B(n15549), .Z(n15551) );
  XOR U15880 ( .A(n15552), .B(n15551), .Z(n15484) );
  NANDN U15881 ( .A(n15473), .B(n15472), .Z(n15477) );
  NAND U15882 ( .A(n15475), .B(n15474), .Z(n15476) );
  AND U15883 ( .A(n15477), .B(n15476), .Z(n15483) );
  XNOR U15884 ( .A(n15484), .B(n15483), .Z(n15485) );
  XNOR U15885 ( .A(n15486), .B(n15485), .Z(n15555) );
  XNOR U15886 ( .A(sreg[448]), .B(n15555), .Z(n15557) );
  NANDN U15887 ( .A(sreg[447]), .B(n15478), .Z(n15482) );
  NAND U15888 ( .A(n15480), .B(n15479), .Z(n15481) );
  NAND U15889 ( .A(n15482), .B(n15481), .Z(n15556) );
  XNOR U15890 ( .A(n15557), .B(n15556), .Z(c[448]) );
  NANDN U15891 ( .A(n15484), .B(n15483), .Z(n15488) );
  NANDN U15892 ( .A(n15486), .B(n15485), .Z(n15487) );
  AND U15893 ( .A(n15488), .B(n15487), .Z(n15563) );
  NANDN U15894 ( .A(n15490), .B(n15489), .Z(n15494) );
  NAND U15895 ( .A(n15492), .B(n15491), .Z(n15493) );
  AND U15896 ( .A(n15494), .B(n15493), .Z(n15629) );
  NAND U15897 ( .A(n15495), .B(n19724), .Z(n15497) );
  XOR U15898 ( .A(b[11]), .B(a[199]), .Z(n15599) );
  NAND U15899 ( .A(n19692), .B(n15599), .Z(n15496) );
  AND U15900 ( .A(n15497), .B(n15496), .Z(n15610) );
  NAND U15901 ( .A(n19838), .B(n15498), .Z(n15500) );
  XOR U15902 ( .A(b[15]), .B(a[195]), .Z(n15602) );
  NAND U15903 ( .A(n19805), .B(n15602), .Z(n15499) );
  AND U15904 ( .A(n15500), .B(n15499), .Z(n15609) );
  NAND U15905 ( .A(n35), .B(n15501), .Z(n15503) );
  XOR U15906 ( .A(b[9]), .B(a[201]), .Z(n15605) );
  NAND U15907 ( .A(n19598), .B(n15605), .Z(n15502) );
  NAND U15908 ( .A(n15503), .B(n15502), .Z(n15608) );
  XOR U15909 ( .A(n15609), .B(n15608), .Z(n15611) );
  XOR U15910 ( .A(n15610), .B(n15611), .Z(n15621) );
  NANDN U15911 ( .A(n15505), .B(n15504), .Z(n15509) );
  OR U15912 ( .A(n15507), .B(n15506), .Z(n15508) );
  AND U15913 ( .A(n15509), .B(n15508), .Z(n15620) );
  XNOR U15914 ( .A(n15621), .B(n15620), .Z(n15622) );
  NANDN U15915 ( .A(n15511), .B(n15510), .Z(n15515) );
  NANDN U15916 ( .A(n15513), .B(n15512), .Z(n15514) );
  NAND U15917 ( .A(n15515), .B(n15514), .Z(n15623) );
  XNOR U15918 ( .A(n15622), .B(n15623), .Z(n15569) );
  NANDN U15919 ( .A(n15517), .B(n15516), .Z(n15521) );
  NANDN U15920 ( .A(n15519), .B(n15518), .Z(n15520) );
  AND U15921 ( .A(n15521), .B(n15520), .Z(n15595) );
  NAND U15922 ( .A(n19808), .B(n15522), .Z(n15524) );
  XOR U15923 ( .A(b[13]), .B(a[197]), .Z(n15581) );
  NAND U15924 ( .A(n19768), .B(n15581), .Z(n15523) );
  AND U15925 ( .A(n15524), .B(n15523), .Z(n15573) );
  AND U15926 ( .A(b[15]), .B(a[193]), .Z(n15572) );
  XNOR U15927 ( .A(n15573), .B(n15572), .Z(n15574) );
  NAND U15928 ( .A(b[0]), .B(a[209]), .Z(n15525) );
  XNOR U15929 ( .A(b[1]), .B(n15525), .Z(n15527) );
  NANDN U15930 ( .A(b[0]), .B(a[208]), .Z(n15526) );
  NAND U15931 ( .A(n15527), .B(n15526), .Z(n15575) );
  XNOR U15932 ( .A(n15574), .B(n15575), .Z(n15593) );
  NAND U15933 ( .A(n33), .B(n15528), .Z(n15530) );
  XOR U15934 ( .A(b[5]), .B(a[205]), .Z(n15584) );
  NAND U15935 ( .A(n19342), .B(n15584), .Z(n15529) );
  AND U15936 ( .A(n15530), .B(n15529), .Z(n15617) );
  NAND U15937 ( .A(n34), .B(n15531), .Z(n15533) );
  XOR U15938 ( .A(b[7]), .B(a[203]), .Z(n15587) );
  NAND U15939 ( .A(n19486), .B(n15587), .Z(n15532) );
  AND U15940 ( .A(n15533), .B(n15532), .Z(n15615) );
  NAND U15941 ( .A(n31), .B(n15534), .Z(n15536) );
  XOR U15942 ( .A(b[3]), .B(a[207]), .Z(n15590) );
  NAND U15943 ( .A(n32), .B(n15590), .Z(n15535) );
  NAND U15944 ( .A(n15536), .B(n15535), .Z(n15614) );
  XNOR U15945 ( .A(n15615), .B(n15614), .Z(n15616) );
  XOR U15946 ( .A(n15617), .B(n15616), .Z(n15594) );
  XOR U15947 ( .A(n15593), .B(n15594), .Z(n15596) );
  XOR U15948 ( .A(n15595), .B(n15596), .Z(n15567) );
  NANDN U15949 ( .A(n15538), .B(n15537), .Z(n15542) );
  OR U15950 ( .A(n15540), .B(n15539), .Z(n15541) );
  AND U15951 ( .A(n15542), .B(n15541), .Z(n15566) );
  XNOR U15952 ( .A(n15567), .B(n15566), .Z(n15568) );
  XOR U15953 ( .A(n15569), .B(n15568), .Z(n15627) );
  NANDN U15954 ( .A(n15544), .B(n15543), .Z(n15548) );
  NANDN U15955 ( .A(n15546), .B(n15545), .Z(n15547) );
  AND U15956 ( .A(n15548), .B(n15547), .Z(n15626) );
  XNOR U15957 ( .A(n15627), .B(n15626), .Z(n15628) );
  XOR U15958 ( .A(n15629), .B(n15628), .Z(n15561) );
  NANDN U15959 ( .A(n15550), .B(n15549), .Z(n15554) );
  NAND U15960 ( .A(n15552), .B(n15551), .Z(n15553) );
  AND U15961 ( .A(n15554), .B(n15553), .Z(n15560) );
  XNOR U15962 ( .A(n15561), .B(n15560), .Z(n15562) );
  XNOR U15963 ( .A(n15563), .B(n15562), .Z(n15632) );
  XNOR U15964 ( .A(sreg[449]), .B(n15632), .Z(n15634) );
  NANDN U15965 ( .A(sreg[448]), .B(n15555), .Z(n15559) );
  NAND U15966 ( .A(n15557), .B(n15556), .Z(n15558) );
  NAND U15967 ( .A(n15559), .B(n15558), .Z(n15633) );
  XNOR U15968 ( .A(n15634), .B(n15633), .Z(c[449]) );
  NANDN U15969 ( .A(n15561), .B(n15560), .Z(n15565) );
  NANDN U15970 ( .A(n15563), .B(n15562), .Z(n15564) );
  AND U15971 ( .A(n15565), .B(n15564), .Z(n15640) );
  NANDN U15972 ( .A(n15567), .B(n15566), .Z(n15571) );
  NAND U15973 ( .A(n15569), .B(n15568), .Z(n15570) );
  AND U15974 ( .A(n15571), .B(n15570), .Z(n15706) );
  NANDN U15975 ( .A(n15573), .B(n15572), .Z(n15577) );
  NANDN U15976 ( .A(n15575), .B(n15574), .Z(n15576) );
  AND U15977 ( .A(n15577), .B(n15576), .Z(n15672) );
  NAND U15978 ( .A(b[0]), .B(a[210]), .Z(n15578) );
  XNOR U15979 ( .A(b[1]), .B(n15578), .Z(n15580) );
  NANDN U15980 ( .A(b[0]), .B(a[209]), .Z(n15579) );
  NAND U15981 ( .A(n15580), .B(n15579), .Z(n15652) );
  NAND U15982 ( .A(n19808), .B(n15581), .Z(n15583) );
  XOR U15983 ( .A(b[13]), .B(a[198]), .Z(n15658) );
  NAND U15984 ( .A(n19768), .B(n15658), .Z(n15582) );
  AND U15985 ( .A(n15583), .B(n15582), .Z(n15650) );
  AND U15986 ( .A(b[15]), .B(a[194]), .Z(n15649) );
  XNOR U15987 ( .A(n15650), .B(n15649), .Z(n15651) );
  XNOR U15988 ( .A(n15652), .B(n15651), .Z(n15670) );
  NAND U15989 ( .A(n33), .B(n15584), .Z(n15586) );
  XOR U15990 ( .A(b[5]), .B(a[206]), .Z(n15661) );
  NAND U15991 ( .A(n19342), .B(n15661), .Z(n15585) );
  AND U15992 ( .A(n15586), .B(n15585), .Z(n15694) );
  NAND U15993 ( .A(n34), .B(n15587), .Z(n15589) );
  XOR U15994 ( .A(b[7]), .B(a[204]), .Z(n15664) );
  NAND U15995 ( .A(n19486), .B(n15664), .Z(n15588) );
  AND U15996 ( .A(n15589), .B(n15588), .Z(n15692) );
  NAND U15997 ( .A(n31), .B(n15590), .Z(n15592) );
  XOR U15998 ( .A(b[3]), .B(a[208]), .Z(n15667) );
  NAND U15999 ( .A(n32), .B(n15667), .Z(n15591) );
  NAND U16000 ( .A(n15592), .B(n15591), .Z(n15691) );
  XNOR U16001 ( .A(n15692), .B(n15691), .Z(n15693) );
  XOR U16002 ( .A(n15694), .B(n15693), .Z(n15671) );
  XOR U16003 ( .A(n15670), .B(n15671), .Z(n15673) );
  XOR U16004 ( .A(n15672), .B(n15673), .Z(n15644) );
  NANDN U16005 ( .A(n15594), .B(n15593), .Z(n15598) );
  OR U16006 ( .A(n15596), .B(n15595), .Z(n15597) );
  AND U16007 ( .A(n15598), .B(n15597), .Z(n15643) );
  XNOR U16008 ( .A(n15644), .B(n15643), .Z(n15646) );
  NAND U16009 ( .A(n15599), .B(n19724), .Z(n15601) );
  XOR U16010 ( .A(b[11]), .B(a[200]), .Z(n15676) );
  NAND U16011 ( .A(n19692), .B(n15676), .Z(n15600) );
  AND U16012 ( .A(n15601), .B(n15600), .Z(n15687) );
  NAND U16013 ( .A(n19838), .B(n15602), .Z(n15604) );
  XOR U16014 ( .A(b[15]), .B(a[196]), .Z(n15679) );
  NAND U16015 ( .A(n19805), .B(n15679), .Z(n15603) );
  AND U16016 ( .A(n15604), .B(n15603), .Z(n15686) );
  NAND U16017 ( .A(n35), .B(n15605), .Z(n15607) );
  XOR U16018 ( .A(b[9]), .B(a[202]), .Z(n15682) );
  NAND U16019 ( .A(n19598), .B(n15682), .Z(n15606) );
  NAND U16020 ( .A(n15607), .B(n15606), .Z(n15685) );
  XOR U16021 ( .A(n15686), .B(n15685), .Z(n15688) );
  XOR U16022 ( .A(n15687), .B(n15688), .Z(n15698) );
  NANDN U16023 ( .A(n15609), .B(n15608), .Z(n15613) );
  OR U16024 ( .A(n15611), .B(n15610), .Z(n15612) );
  AND U16025 ( .A(n15613), .B(n15612), .Z(n15697) );
  XNOR U16026 ( .A(n15698), .B(n15697), .Z(n15699) );
  NANDN U16027 ( .A(n15615), .B(n15614), .Z(n15619) );
  NANDN U16028 ( .A(n15617), .B(n15616), .Z(n15618) );
  NAND U16029 ( .A(n15619), .B(n15618), .Z(n15700) );
  XNOR U16030 ( .A(n15699), .B(n15700), .Z(n15645) );
  XOR U16031 ( .A(n15646), .B(n15645), .Z(n15704) );
  NANDN U16032 ( .A(n15621), .B(n15620), .Z(n15625) );
  NANDN U16033 ( .A(n15623), .B(n15622), .Z(n15624) );
  AND U16034 ( .A(n15625), .B(n15624), .Z(n15703) );
  XNOR U16035 ( .A(n15704), .B(n15703), .Z(n15705) );
  XOR U16036 ( .A(n15706), .B(n15705), .Z(n15638) );
  NANDN U16037 ( .A(n15627), .B(n15626), .Z(n15631) );
  NAND U16038 ( .A(n15629), .B(n15628), .Z(n15630) );
  AND U16039 ( .A(n15631), .B(n15630), .Z(n15637) );
  XNOR U16040 ( .A(n15638), .B(n15637), .Z(n15639) );
  XNOR U16041 ( .A(n15640), .B(n15639), .Z(n15709) );
  XNOR U16042 ( .A(sreg[450]), .B(n15709), .Z(n15711) );
  NANDN U16043 ( .A(sreg[449]), .B(n15632), .Z(n15636) );
  NAND U16044 ( .A(n15634), .B(n15633), .Z(n15635) );
  NAND U16045 ( .A(n15636), .B(n15635), .Z(n15710) );
  XNOR U16046 ( .A(n15711), .B(n15710), .Z(c[450]) );
  NANDN U16047 ( .A(n15638), .B(n15637), .Z(n15642) );
  NANDN U16048 ( .A(n15640), .B(n15639), .Z(n15641) );
  AND U16049 ( .A(n15642), .B(n15641), .Z(n15717) );
  NANDN U16050 ( .A(n15644), .B(n15643), .Z(n15648) );
  NAND U16051 ( .A(n15646), .B(n15645), .Z(n15647) );
  AND U16052 ( .A(n15648), .B(n15647), .Z(n15783) );
  NANDN U16053 ( .A(n15650), .B(n15649), .Z(n15654) );
  NANDN U16054 ( .A(n15652), .B(n15651), .Z(n15653) );
  AND U16055 ( .A(n15654), .B(n15653), .Z(n15749) );
  NAND U16056 ( .A(b[0]), .B(a[211]), .Z(n15655) );
  XNOR U16057 ( .A(b[1]), .B(n15655), .Z(n15657) );
  NANDN U16058 ( .A(b[0]), .B(a[210]), .Z(n15656) );
  NAND U16059 ( .A(n15657), .B(n15656), .Z(n15729) );
  NAND U16060 ( .A(n19808), .B(n15658), .Z(n15660) );
  XOR U16061 ( .A(b[13]), .B(a[199]), .Z(n15735) );
  NAND U16062 ( .A(n19768), .B(n15735), .Z(n15659) );
  AND U16063 ( .A(n15660), .B(n15659), .Z(n15727) );
  AND U16064 ( .A(b[15]), .B(a[195]), .Z(n15726) );
  XNOR U16065 ( .A(n15727), .B(n15726), .Z(n15728) );
  XNOR U16066 ( .A(n15729), .B(n15728), .Z(n15747) );
  NAND U16067 ( .A(n33), .B(n15661), .Z(n15663) );
  XOR U16068 ( .A(b[5]), .B(a[207]), .Z(n15738) );
  NAND U16069 ( .A(n19342), .B(n15738), .Z(n15662) );
  AND U16070 ( .A(n15663), .B(n15662), .Z(n15771) );
  NAND U16071 ( .A(n34), .B(n15664), .Z(n15666) );
  XOR U16072 ( .A(b[7]), .B(a[205]), .Z(n15741) );
  NAND U16073 ( .A(n19486), .B(n15741), .Z(n15665) );
  AND U16074 ( .A(n15666), .B(n15665), .Z(n15769) );
  NAND U16075 ( .A(n31), .B(n15667), .Z(n15669) );
  XOR U16076 ( .A(b[3]), .B(a[209]), .Z(n15744) );
  NAND U16077 ( .A(n32), .B(n15744), .Z(n15668) );
  NAND U16078 ( .A(n15669), .B(n15668), .Z(n15768) );
  XNOR U16079 ( .A(n15769), .B(n15768), .Z(n15770) );
  XOR U16080 ( .A(n15771), .B(n15770), .Z(n15748) );
  XOR U16081 ( .A(n15747), .B(n15748), .Z(n15750) );
  XOR U16082 ( .A(n15749), .B(n15750), .Z(n15721) );
  NANDN U16083 ( .A(n15671), .B(n15670), .Z(n15675) );
  OR U16084 ( .A(n15673), .B(n15672), .Z(n15674) );
  AND U16085 ( .A(n15675), .B(n15674), .Z(n15720) );
  XNOR U16086 ( .A(n15721), .B(n15720), .Z(n15723) );
  NAND U16087 ( .A(n15676), .B(n19724), .Z(n15678) );
  XOR U16088 ( .A(b[11]), .B(a[201]), .Z(n15753) );
  NAND U16089 ( .A(n19692), .B(n15753), .Z(n15677) );
  AND U16090 ( .A(n15678), .B(n15677), .Z(n15764) );
  NAND U16091 ( .A(n19838), .B(n15679), .Z(n15681) );
  XOR U16092 ( .A(b[15]), .B(a[197]), .Z(n15756) );
  NAND U16093 ( .A(n19805), .B(n15756), .Z(n15680) );
  AND U16094 ( .A(n15681), .B(n15680), .Z(n15763) );
  NAND U16095 ( .A(n35), .B(n15682), .Z(n15684) );
  XOR U16096 ( .A(b[9]), .B(a[203]), .Z(n15759) );
  NAND U16097 ( .A(n19598), .B(n15759), .Z(n15683) );
  NAND U16098 ( .A(n15684), .B(n15683), .Z(n15762) );
  XOR U16099 ( .A(n15763), .B(n15762), .Z(n15765) );
  XOR U16100 ( .A(n15764), .B(n15765), .Z(n15775) );
  NANDN U16101 ( .A(n15686), .B(n15685), .Z(n15690) );
  OR U16102 ( .A(n15688), .B(n15687), .Z(n15689) );
  AND U16103 ( .A(n15690), .B(n15689), .Z(n15774) );
  XNOR U16104 ( .A(n15775), .B(n15774), .Z(n15776) );
  NANDN U16105 ( .A(n15692), .B(n15691), .Z(n15696) );
  NANDN U16106 ( .A(n15694), .B(n15693), .Z(n15695) );
  NAND U16107 ( .A(n15696), .B(n15695), .Z(n15777) );
  XNOR U16108 ( .A(n15776), .B(n15777), .Z(n15722) );
  XOR U16109 ( .A(n15723), .B(n15722), .Z(n15781) );
  NANDN U16110 ( .A(n15698), .B(n15697), .Z(n15702) );
  NANDN U16111 ( .A(n15700), .B(n15699), .Z(n15701) );
  AND U16112 ( .A(n15702), .B(n15701), .Z(n15780) );
  XNOR U16113 ( .A(n15781), .B(n15780), .Z(n15782) );
  XOR U16114 ( .A(n15783), .B(n15782), .Z(n15715) );
  NANDN U16115 ( .A(n15704), .B(n15703), .Z(n15708) );
  NAND U16116 ( .A(n15706), .B(n15705), .Z(n15707) );
  AND U16117 ( .A(n15708), .B(n15707), .Z(n15714) );
  XNOR U16118 ( .A(n15715), .B(n15714), .Z(n15716) );
  XNOR U16119 ( .A(n15717), .B(n15716), .Z(n15786) );
  XNOR U16120 ( .A(sreg[451]), .B(n15786), .Z(n15788) );
  NANDN U16121 ( .A(sreg[450]), .B(n15709), .Z(n15713) );
  NAND U16122 ( .A(n15711), .B(n15710), .Z(n15712) );
  NAND U16123 ( .A(n15713), .B(n15712), .Z(n15787) );
  XNOR U16124 ( .A(n15788), .B(n15787), .Z(c[451]) );
  NANDN U16125 ( .A(n15715), .B(n15714), .Z(n15719) );
  NANDN U16126 ( .A(n15717), .B(n15716), .Z(n15718) );
  AND U16127 ( .A(n15719), .B(n15718), .Z(n15794) );
  NANDN U16128 ( .A(n15721), .B(n15720), .Z(n15725) );
  NAND U16129 ( .A(n15723), .B(n15722), .Z(n15724) );
  AND U16130 ( .A(n15725), .B(n15724), .Z(n15860) );
  NANDN U16131 ( .A(n15727), .B(n15726), .Z(n15731) );
  NANDN U16132 ( .A(n15729), .B(n15728), .Z(n15730) );
  AND U16133 ( .A(n15731), .B(n15730), .Z(n15826) );
  NAND U16134 ( .A(b[0]), .B(a[212]), .Z(n15732) );
  XNOR U16135 ( .A(b[1]), .B(n15732), .Z(n15734) );
  NANDN U16136 ( .A(b[0]), .B(a[211]), .Z(n15733) );
  NAND U16137 ( .A(n15734), .B(n15733), .Z(n15806) );
  NAND U16138 ( .A(n19808), .B(n15735), .Z(n15737) );
  XOR U16139 ( .A(b[13]), .B(a[200]), .Z(n15809) );
  NAND U16140 ( .A(n19768), .B(n15809), .Z(n15736) );
  AND U16141 ( .A(n15737), .B(n15736), .Z(n15804) );
  AND U16142 ( .A(b[15]), .B(a[196]), .Z(n15803) );
  XNOR U16143 ( .A(n15804), .B(n15803), .Z(n15805) );
  XNOR U16144 ( .A(n15806), .B(n15805), .Z(n15824) );
  NAND U16145 ( .A(n33), .B(n15738), .Z(n15740) );
  XOR U16146 ( .A(b[5]), .B(a[208]), .Z(n15815) );
  NAND U16147 ( .A(n19342), .B(n15815), .Z(n15739) );
  AND U16148 ( .A(n15740), .B(n15739), .Z(n15848) );
  NAND U16149 ( .A(n34), .B(n15741), .Z(n15743) );
  XOR U16150 ( .A(b[7]), .B(a[206]), .Z(n15818) );
  NAND U16151 ( .A(n19486), .B(n15818), .Z(n15742) );
  AND U16152 ( .A(n15743), .B(n15742), .Z(n15846) );
  NAND U16153 ( .A(n31), .B(n15744), .Z(n15746) );
  XOR U16154 ( .A(b[3]), .B(a[210]), .Z(n15821) );
  NAND U16155 ( .A(n32), .B(n15821), .Z(n15745) );
  NAND U16156 ( .A(n15746), .B(n15745), .Z(n15845) );
  XNOR U16157 ( .A(n15846), .B(n15845), .Z(n15847) );
  XOR U16158 ( .A(n15848), .B(n15847), .Z(n15825) );
  XOR U16159 ( .A(n15824), .B(n15825), .Z(n15827) );
  XOR U16160 ( .A(n15826), .B(n15827), .Z(n15798) );
  NANDN U16161 ( .A(n15748), .B(n15747), .Z(n15752) );
  OR U16162 ( .A(n15750), .B(n15749), .Z(n15751) );
  AND U16163 ( .A(n15752), .B(n15751), .Z(n15797) );
  XNOR U16164 ( .A(n15798), .B(n15797), .Z(n15800) );
  NAND U16165 ( .A(n15753), .B(n19724), .Z(n15755) );
  XOR U16166 ( .A(b[11]), .B(a[202]), .Z(n15830) );
  NAND U16167 ( .A(n19692), .B(n15830), .Z(n15754) );
  AND U16168 ( .A(n15755), .B(n15754), .Z(n15841) );
  NAND U16169 ( .A(n19838), .B(n15756), .Z(n15758) );
  XOR U16170 ( .A(b[15]), .B(a[198]), .Z(n15833) );
  NAND U16171 ( .A(n19805), .B(n15833), .Z(n15757) );
  AND U16172 ( .A(n15758), .B(n15757), .Z(n15840) );
  NAND U16173 ( .A(n35), .B(n15759), .Z(n15761) );
  XOR U16174 ( .A(b[9]), .B(a[204]), .Z(n15836) );
  NAND U16175 ( .A(n19598), .B(n15836), .Z(n15760) );
  NAND U16176 ( .A(n15761), .B(n15760), .Z(n15839) );
  XOR U16177 ( .A(n15840), .B(n15839), .Z(n15842) );
  XOR U16178 ( .A(n15841), .B(n15842), .Z(n15852) );
  NANDN U16179 ( .A(n15763), .B(n15762), .Z(n15767) );
  OR U16180 ( .A(n15765), .B(n15764), .Z(n15766) );
  AND U16181 ( .A(n15767), .B(n15766), .Z(n15851) );
  XNOR U16182 ( .A(n15852), .B(n15851), .Z(n15853) );
  NANDN U16183 ( .A(n15769), .B(n15768), .Z(n15773) );
  NANDN U16184 ( .A(n15771), .B(n15770), .Z(n15772) );
  NAND U16185 ( .A(n15773), .B(n15772), .Z(n15854) );
  XNOR U16186 ( .A(n15853), .B(n15854), .Z(n15799) );
  XOR U16187 ( .A(n15800), .B(n15799), .Z(n15858) );
  NANDN U16188 ( .A(n15775), .B(n15774), .Z(n15779) );
  NANDN U16189 ( .A(n15777), .B(n15776), .Z(n15778) );
  AND U16190 ( .A(n15779), .B(n15778), .Z(n15857) );
  XNOR U16191 ( .A(n15858), .B(n15857), .Z(n15859) );
  XOR U16192 ( .A(n15860), .B(n15859), .Z(n15792) );
  NANDN U16193 ( .A(n15781), .B(n15780), .Z(n15785) );
  NAND U16194 ( .A(n15783), .B(n15782), .Z(n15784) );
  AND U16195 ( .A(n15785), .B(n15784), .Z(n15791) );
  XNOR U16196 ( .A(n15792), .B(n15791), .Z(n15793) );
  XNOR U16197 ( .A(n15794), .B(n15793), .Z(n15863) );
  XNOR U16198 ( .A(sreg[452]), .B(n15863), .Z(n15865) );
  NANDN U16199 ( .A(sreg[451]), .B(n15786), .Z(n15790) );
  NAND U16200 ( .A(n15788), .B(n15787), .Z(n15789) );
  NAND U16201 ( .A(n15790), .B(n15789), .Z(n15864) );
  XNOR U16202 ( .A(n15865), .B(n15864), .Z(c[452]) );
  NANDN U16203 ( .A(n15792), .B(n15791), .Z(n15796) );
  NANDN U16204 ( .A(n15794), .B(n15793), .Z(n15795) );
  AND U16205 ( .A(n15796), .B(n15795), .Z(n15871) );
  NANDN U16206 ( .A(n15798), .B(n15797), .Z(n15802) );
  NAND U16207 ( .A(n15800), .B(n15799), .Z(n15801) );
  AND U16208 ( .A(n15802), .B(n15801), .Z(n15937) );
  NANDN U16209 ( .A(n15804), .B(n15803), .Z(n15808) );
  NANDN U16210 ( .A(n15806), .B(n15805), .Z(n15807) );
  AND U16211 ( .A(n15808), .B(n15807), .Z(n15903) );
  NAND U16212 ( .A(n19808), .B(n15809), .Z(n15811) );
  XOR U16213 ( .A(b[13]), .B(a[201]), .Z(n15889) );
  NAND U16214 ( .A(n19768), .B(n15889), .Z(n15810) );
  AND U16215 ( .A(n15811), .B(n15810), .Z(n15881) );
  AND U16216 ( .A(b[15]), .B(a[197]), .Z(n15880) );
  XNOR U16217 ( .A(n15881), .B(n15880), .Z(n15882) );
  NAND U16218 ( .A(b[0]), .B(a[213]), .Z(n15812) );
  XNOR U16219 ( .A(b[1]), .B(n15812), .Z(n15814) );
  NANDN U16220 ( .A(b[0]), .B(a[212]), .Z(n15813) );
  NAND U16221 ( .A(n15814), .B(n15813), .Z(n15883) );
  XNOR U16222 ( .A(n15882), .B(n15883), .Z(n15901) );
  NAND U16223 ( .A(n33), .B(n15815), .Z(n15817) );
  XOR U16224 ( .A(b[5]), .B(a[209]), .Z(n15892) );
  NAND U16225 ( .A(n19342), .B(n15892), .Z(n15816) );
  AND U16226 ( .A(n15817), .B(n15816), .Z(n15925) );
  NAND U16227 ( .A(n34), .B(n15818), .Z(n15820) );
  XOR U16228 ( .A(b[7]), .B(a[207]), .Z(n15895) );
  NAND U16229 ( .A(n19486), .B(n15895), .Z(n15819) );
  AND U16230 ( .A(n15820), .B(n15819), .Z(n15923) );
  NAND U16231 ( .A(n31), .B(n15821), .Z(n15823) );
  XOR U16232 ( .A(b[3]), .B(a[211]), .Z(n15898) );
  NAND U16233 ( .A(n32), .B(n15898), .Z(n15822) );
  NAND U16234 ( .A(n15823), .B(n15822), .Z(n15922) );
  XNOR U16235 ( .A(n15923), .B(n15922), .Z(n15924) );
  XOR U16236 ( .A(n15925), .B(n15924), .Z(n15902) );
  XOR U16237 ( .A(n15901), .B(n15902), .Z(n15904) );
  XOR U16238 ( .A(n15903), .B(n15904), .Z(n15875) );
  NANDN U16239 ( .A(n15825), .B(n15824), .Z(n15829) );
  OR U16240 ( .A(n15827), .B(n15826), .Z(n15828) );
  AND U16241 ( .A(n15829), .B(n15828), .Z(n15874) );
  XNOR U16242 ( .A(n15875), .B(n15874), .Z(n15877) );
  NAND U16243 ( .A(n15830), .B(n19724), .Z(n15832) );
  XOR U16244 ( .A(b[11]), .B(a[203]), .Z(n15907) );
  NAND U16245 ( .A(n19692), .B(n15907), .Z(n15831) );
  AND U16246 ( .A(n15832), .B(n15831), .Z(n15918) );
  NAND U16247 ( .A(n19838), .B(n15833), .Z(n15835) );
  XOR U16248 ( .A(b[15]), .B(a[199]), .Z(n15910) );
  NAND U16249 ( .A(n19805), .B(n15910), .Z(n15834) );
  AND U16250 ( .A(n15835), .B(n15834), .Z(n15917) );
  NAND U16251 ( .A(n35), .B(n15836), .Z(n15838) );
  XOR U16252 ( .A(b[9]), .B(a[205]), .Z(n15913) );
  NAND U16253 ( .A(n19598), .B(n15913), .Z(n15837) );
  NAND U16254 ( .A(n15838), .B(n15837), .Z(n15916) );
  XOR U16255 ( .A(n15917), .B(n15916), .Z(n15919) );
  XOR U16256 ( .A(n15918), .B(n15919), .Z(n15929) );
  NANDN U16257 ( .A(n15840), .B(n15839), .Z(n15844) );
  OR U16258 ( .A(n15842), .B(n15841), .Z(n15843) );
  AND U16259 ( .A(n15844), .B(n15843), .Z(n15928) );
  XNOR U16260 ( .A(n15929), .B(n15928), .Z(n15930) );
  NANDN U16261 ( .A(n15846), .B(n15845), .Z(n15850) );
  NANDN U16262 ( .A(n15848), .B(n15847), .Z(n15849) );
  NAND U16263 ( .A(n15850), .B(n15849), .Z(n15931) );
  XNOR U16264 ( .A(n15930), .B(n15931), .Z(n15876) );
  XOR U16265 ( .A(n15877), .B(n15876), .Z(n15935) );
  NANDN U16266 ( .A(n15852), .B(n15851), .Z(n15856) );
  NANDN U16267 ( .A(n15854), .B(n15853), .Z(n15855) );
  AND U16268 ( .A(n15856), .B(n15855), .Z(n15934) );
  XNOR U16269 ( .A(n15935), .B(n15934), .Z(n15936) );
  XOR U16270 ( .A(n15937), .B(n15936), .Z(n15869) );
  NANDN U16271 ( .A(n15858), .B(n15857), .Z(n15862) );
  NAND U16272 ( .A(n15860), .B(n15859), .Z(n15861) );
  AND U16273 ( .A(n15862), .B(n15861), .Z(n15868) );
  XNOR U16274 ( .A(n15869), .B(n15868), .Z(n15870) );
  XNOR U16275 ( .A(n15871), .B(n15870), .Z(n15940) );
  XNOR U16276 ( .A(sreg[453]), .B(n15940), .Z(n15942) );
  NANDN U16277 ( .A(sreg[452]), .B(n15863), .Z(n15867) );
  NAND U16278 ( .A(n15865), .B(n15864), .Z(n15866) );
  NAND U16279 ( .A(n15867), .B(n15866), .Z(n15941) );
  XNOR U16280 ( .A(n15942), .B(n15941), .Z(c[453]) );
  NANDN U16281 ( .A(n15869), .B(n15868), .Z(n15873) );
  NANDN U16282 ( .A(n15871), .B(n15870), .Z(n15872) );
  AND U16283 ( .A(n15873), .B(n15872), .Z(n15948) );
  NANDN U16284 ( .A(n15875), .B(n15874), .Z(n15879) );
  NAND U16285 ( .A(n15877), .B(n15876), .Z(n15878) );
  AND U16286 ( .A(n15879), .B(n15878), .Z(n16014) );
  NANDN U16287 ( .A(n15881), .B(n15880), .Z(n15885) );
  NANDN U16288 ( .A(n15883), .B(n15882), .Z(n15884) );
  AND U16289 ( .A(n15885), .B(n15884), .Z(n16001) );
  NAND U16290 ( .A(b[0]), .B(a[214]), .Z(n15886) );
  XNOR U16291 ( .A(b[1]), .B(n15886), .Z(n15888) );
  NANDN U16292 ( .A(b[0]), .B(a[213]), .Z(n15887) );
  NAND U16293 ( .A(n15888), .B(n15887), .Z(n15981) );
  NAND U16294 ( .A(n19808), .B(n15889), .Z(n15891) );
  XOR U16295 ( .A(b[13]), .B(a[202]), .Z(n15987) );
  NAND U16296 ( .A(n19768), .B(n15987), .Z(n15890) );
  AND U16297 ( .A(n15891), .B(n15890), .Z(n15979) );
  AND U16298 ( .A(b[15]), .B(a[198]), .Z(n15978) );
  XNOR U16299 ( .A(n15979), .B(n15978), .Z(n15980) );
  XNOR U16300 ( .A(n15981), .B(n15980), .Z(n15999) );
  NAND U16301 ( .A(n33), .B(n15892), .Z(n15894) );
  XOR U16302 ( .A(b[5]), .B(a[210]), .Z(n15990) );
  NAND U16303 ( .A(n19342), .B(n15990), .Z(n15893) );
  AND U16304 ( .A(n15894), .B(n15893), .Z(n15975) );
  NAND U16305 ( .A(n34), .B(n15895), .Z(n15897) );
  XOR U16306 ( .A(b[7]), .B(a[208]), .Z(n15993) );
  NAND U16307 ( .A(n19486), .B(n15993), .Z(n15896) );
  AND U16308 ( .A(n15897), .B(n15896), .Z(n15973) );
  NAND U16309 ( .A(n31), .B(n15898), .Z(n15900) );
  XOR U16310 ( .A(b[3]), .B(a[212]), .Z(n15996) );
  NAND U16311 ( .A(n32), .B(n15996), .Z(n15899) );
  NAND U16312 ( .A(n15900), .B(n15899), .Z(n15972) );
  XNOR U16313 ( .A(n15973), .B(n15972), .Z(n15974) );
  XOR U16314 ( .A(n15975), .B(n15974), .Z(n16000) );
  XOR U16315 ( .A(n15999), .B(n16000), .Z(n16002) );
  XOR U16316 ( .A(n16001), .B(n16002), .Z(n15952) );
  NANDN U16317 ( .A(n15902), .B(n15901), .Z(n15906) );
  OR U16318 ( .A(n15904), .B(n15903), .Z(n15905) );
  AND U16319 ( .A(n15906), .B(n15905), .Z(n15951) );
  XNOR U16320 ( .A(n15952), .B(n15951), .Z(n15954) );
  NAND U16321 ( .A(n15907), .B(n19724), .Z(n15909) );
  XOR U16322 ( .A(b[11]), .B(a[204]), .Z(n15957) );
  NAND U16323 ( .A(n19692), .B(n15957), .Z(n15908) );
  AND U16324 ( .A(n15909), .B(n15908), .Z(n15968) );
  NAND U16325 ( .A(n19838), .B(n15910), .Z(n15912) );
  XOR U16326 ( .A(b[15]), .B(a[200]), .Z(n15960) );
  NAND U16327 ( .A(n19805), .B(n15960), .Z(n15911) );
  AND U16328 ( .A(n15912), .B(n15911), .Z(n15967) );
  NAND U16329 ( .A(n35), .B(n15913), .Z(n15915) );
  XOR U16330 ( .A(b[9]), .B(a[206]), .Z(n15963) );
  NAND U16331 ( .A(n19598), .B(n15963), .Z(n15914) );
  NAND U16332 ( .A(n15915), .B(n15914), .Z(n15966) );
  XOR U16333 ( .A(n15967), .B(n15966), .Z(n15969) );
  XOR U16334 ( .A(n15968), .B(n15969), .Z(n16006) );
  NANDN U16335 ( .A(n15917), .B(n15916), .Z(n15921) );
  OR U16336 ( .A(n15919), .B(n15918), .Z(n15920) );
  AND U16337 ( .A(n15921), .B(n15920), .Z(n16005) );
  XNOR U16338 ( .A(n16006), .B(n16005), .Z(n16007) );
  NANDN U16339 ( .A(n15923), .B(n15922), .Z(n15927) );
  NANDN U16340 ( .A(n15925), .B(n15924), .Z(n15926) );
  NAND U16341 ( .A(n15927), .B(n15926), .Z(n16008) );
  XNOR U16342 ( .A(n16007), .B(n16008), .Z(n15953) );
  XOR U16343 ( .A(n15954), .B(n15953), .Z(n16012) );
  NANDN U16344 ( .A(n15929), .B(n15928), .Z(n15933) );
  NANDN U16345 ( .A(n15931), .B(n15930), .Z(n15932) );
  AND U16346 ( .A(n15933), .B(n15932), .Z(n16011) );
  XNOR U16347 ( .A(n16012), .B(n16011), .Z(n16013) );
  XOR U16348 ( .A(n16014), .B(n16013), .Z(n15946) );
  NANDN U16349 ( .A(n15935), .B(n15934), .Z(n15939) );
  NAND U16350 ( .A(n15937), .B(n15936), .Z(n15938) );
  AND U16351 ( .A(n15939), .B(n15938), .Z(n15945) );
  XNOR U16352 ( .A(n15946), .B(n15945), .Z(n15947) );
  XNOR U16353 ( .A(n15948), .B(n15947), .Z(n16017) );
  XNOR U16354 ( .A(sreg[454]), .B(n16017), .Z(n16019) );
  NANDN U16355 ( .A(sreg[453]), .B(n15940), .Z(n15944) );
  NAND U16356 ( .A(n15942), .B(n15941), .Z(n15943) );
  NAND U16357 ( .A(n15944), .B(n15943), .Z(n16018) );
  XNOR U16358 ( .A(n16019), .B(n16018), .Z(c[454]) );
  NANDN U16359 ( .A(n15946), .B(n15945), .Z(n15950) );
  NANDN U16360 ( .A(n15948), .B(n15947), .Z(n15949) );
  AND U16361 ( .A(n15950), .B(n15949), .Z(n16025) );
  NANDN U16362 ( .A(n15952), .B(n15951), .Z(n15956) );
  NAND U16363 ( .A(n15954), .B(n15953), .Z(n15955) );
  AND U16364 ( .A(n15956), .B(n15955), .Z(n16091) );
  NAND U16365 ( .A(n15957), .B(n19724), .Z(n15959) );
  XOR U16366 ( .A(b[11]), .B(a[205]), .Z(n16034) );
  NAND U16367 ( .A(n19692), .B(n16034), .Z(n15958) );
  AND U16368 ( .A(n15959), .B(n15958), .Z(n16045) );
  NAND U16369 ( .A(n19838), .B(n15960), .Z(n15962) );
  XOR U16370 ( .A(b[15]), .B(a[201]), .Z(n16037) );
  NAND U16371 ( .A(n19805), .B(n16037), .Z(n15961) );
  AND U16372 ( .A(n15962), .B(n15961), .Z(n16044) );
  NAND U16373 ( .A(n35), .B(n15963), .Z(n15965) );
  XOR U16374 ( .A(b[9]), .B(a[207]), .Z(n16040) );
  NAND U16375 ( .A(n19598), .B(n16040), .Z(n15964) );
  NAND U16376 ( .A(n15965), .B(n15964), .Z(n16043) );
  XOR U16377 ( .A(n16044), .B(n16043), .Z(n16046) );
  XOR U16378 ( .A(n16045), .B(n16046), .Z(n16083) );
  NANDN U16379 ( .A(n15967), .B(n15966), .Z(n15971) );
  OR U16380 ( .A(n15969), .B(n15968), .Z(n15970) );
  AND U16381 ( .A(n15971), .B(n15970), .Z(n16082) );
  XNOR U16382 ( .A(n16083), .B(n16082), .Z(n16084) );
  NANDN U16383 ( .A(n15973), .B(n15972), .Z(n15977) );
  NANDN U16384 ( .A(n15975), .B(n15974), .Z(n15976) );
  NAND U16385 ( .A(n15977), .B(n15976), .Z(n16085) );
  XNOR U16386 ( .A(n16084), .B(n16085), .Z(n16031) );
  NANDN U16387 ( .A(n15979), .B(n15978), .Z(n15983) );
  NANDN U16388 ( .A(n15981), .B(n15980), .Z(n15982) );
  AND U16389 ( .A(n15983), .B(n15982), .Z(n16078) );
  NAND U16390 ( .A(b[0]), .B(a[215]), .Z(n15984) );
  XNOR U16391 ( .A(b[1]), .B(n15984), .Z(n15986) );
  NANDN U16392 ( .A(b[0]), .B(a[214]), .Z(n15985) );
  NAND U16393 ( .A(n15986), .B(n15985), .Z(n16058) );
  NAND U16394 ( .A(n19808), .B(n15987), .Z(n15989) );
  XOR U16395 ( .A(b[13]), .B(a[203]), .Z(n16064) );
  NAND U16396 ( .A(n19768), .B(n16064), .Z(n15988) );
  AND U16397 ( .A(n15989), .B(n15988), .Z(n16056) );
  AND U16398 ( .A(b[15]), .B(a[199]), .Z(n16055) );
  XNOR U16399 ( .A(n16056), .B(n16055), .Z(n16057) );
  XNOR U16400 ( .A(n16058), .B(n16057), .Z(n16076) );
  NAND U16401 ( .A(n33), .B(n15990), .Z(n15992) );
  XOR U16402 ( .A(b[5]), .B(a[211]), .Z(n16067) );
  NAND U16403 ( .A(n19342), .B(n16067), .Z(n15991) );
  AND U16404 ( .A(n15992), .B(n15991), .Z(n16052) );
  NAND U16405 ( .A(n34), .B(n15993), .Z(n15995) );
  XOR U16406 ( .A(b[7]), .B(a[209]), .Z(n16070) );
  NAND U16407 ( .A(n19486), .B(n16070), .Z(n15994) );
  AND U16408 ( .A(n15995), .B(n15994), .Z(n16050) );
  NAND U16409 ( .A(n31), .B(n15996), .Z(n15998) );
  XOR U16410 ( .A(b[3]), .B(a[213]), .Z(n16073) );
  NAND U16411 ( .A(n32), .B(n16073), .Z(n15997) );
  NAND U16412 ( .A(n15998), .B(n15997), .Z(n16049) );
  XNOR U16413 ( .A(n16050), .B(n16049), .Z(n16051) );
  XOR U16414 ( .A(n16052), .B(n16051), .Z(n16077) );
  XOR U16415 ( .A(n16076), .B(n16077), .Z(n16079) );
  XOR U16416 ( .A(n16078), .B(n16079), .Z(n16029) );
  NANDN U16417 ( .A(n16000), .B(n15999), .Z(n16004) );
  OR U16418 ( .A(n16002), .B(n16001), .Z(n16003) );
  AND U16419 ( .A(n16004), .B(n16003), .Z(n16028) );
  XNOR U16420 ( .A(n16029), .B(n16028), .Z(n16030) );
  XOR U16421 ( .A(n16031), .B(n16030), .Z(n16089) );
  NANDN U16422 ( .A(n16006), .B(n16005), .Z(n16010) );
  NANDN U16423 ( .A(n16008), .B(n16007), .Z(n16009) );
  AND U16424 ( .A(n16010), .B(n16009), .Z(n16088) );
  XNOR U16425 ( .A(n16089), .B(n16088), .Z(n16090) );
  XOR U16426 ( .A(n16091), .B(n16090), .Z(n16023) );
  NANDN U16427 ( .A(n16012), .B(n16011), .Z(n16016) );
  NAND U16428 ( .A(n16014), .B(n16013), .Z(n16015) );
  AND U16429 ( .A(n16016), .B(n16015), .Z(n16022) );
  XNOR U16430 ( .A(n16023), .B(n16022), .Z(n16024) );
  XNOR U16431 ( .A(n16025), .B(n16024), .Z(n16094) );
  XNOR U16432 ( .A(sreg[455]), .B(n16094), .Z(n16096) );
  NANDN U16433 ( .A(sreg[454]), .B(n16017), .Z(n16021) );
  NAND U16434 ( .A(n16019), .B(n16018), .Z(n16020) );
  NAND U16435 ( .A(n16021), .B(n16020), .Z(n16095) );
  XNOR U16436 ( .A(n16096), .B(n16095), .Z(c[455]) );
  NANDN U16437 ( .A(n16023), .B(n16022), .Z(n16027) );
  NANDN U16438 ( .A(n16025), .B(n16024), .Z(n16026) );
  AND U16439 ( .A(n16027), .B(n16026), .Z(n16102) );
  NANDN U16440 ( .A(n16029), .B(n16028), .Z(n16033) );
  NAND U16441 ( .A(n16031), .B(n16030), .Z(n16032) );
  AND U16442 ( .A(n16033), .B(n16032), .Z(n16168) );
  NAND U16443 ( .A(n16034), .B(n19724), .Z(n16036) );
  XOR U16444 ( .A(b[11]), .B(a[206]), .Z(n16138) );
  NAND U16445 ( .A(n19692), .B(n16138), .Z(n16035) );
  AND U16446 ( .A(n16036), .B(n16035), .Z(n16149) );
  NAND U16447 ( .A(n19838), .B(n16037), .Z(n16039) );
  XOR U16448 ( .A(b[15]), .B(a[202]), .Z(n16141) );
  NAND U16449 ( .A(n19805), .B(n16141), .Z(n16038) );
  AND U16450 ( .A(n16039), .B(n16038), .Z(n16148) );
  NAND U16451 ( .A(n35), .B(n16040), .Z(n16042) );
  XOR U16452 ( .A(b[9]), .B(a[208]), .Z(n16144) );
  NAND U16453 ( .A(n19598), .B(n16144), .Z(n16041) );
  NAND U16454 ( .A(n16042), .B(n16041), .Z(n16147) );
  XOR U16455 ( .A(n16148), .B(n16147), .Z(n16150) );
  XOR U16456 ( .A(n16149), .B(n16150), .Z(n16160) );
  NANDN U16457 ( .A(n16044), .B(n16043), .Z(n16048) );
  OR U16458 ( .A(n16046), .B(n16045), .Z(n16047) );
  AND U16459 ( .A(n16048), .B(n16047), .Z(n16159) );
  XNOR U16460 ( .A(n16160), .B(n16159), .Z(n16161) );
  NANDN U16461 ( .A(n16050), .B(n16049), .Z(n16054) );
  NANDN U16462 ( .A(n16052), .B(n16051), .Z(n16053) );
  NAND U16463 ( .A(n16054), .B(n16053), .Z(n16162) );
  XNOR U16464 ( .A(n16161), .B(n16162), .Z(n16108) );
  NANDN U16465 ( .A(n16056), .B(n16055), .Z(n16060) );
  NANDN U16466 ( .A(n16058), .B(n16057), .Z(n16059) );
  AND U16467 ( .A(n16060), .B(n16059), .Z(n16134) );
  NAND U16468 ( .A(b[0]), .B(a[216]), .Z(n16061) );
  XNOR U16469 ( .A(b[1]), .B(n16061), .Z(n16063) );
  NANDN U16470 ( .A(b[0]), .B(a[215]), .Z(n16062) );
  NAND U16471 ( .A(n16063), .B(n16062), .Z(n16114) );
  NAND U16472 ( .A(n19808), .B(n16064), .Z(n16066) );
  XOR U16473 ( .A(b[13]), .B(a[204]), .Z(n16120) );
  NAND U16474 ( .A(n19768), .B(n16120), .Z(n16065) );
  AND U16475 ( .A(n16066), .B(n16065), .Z(n16112) );
  AND U16476 ( .A(b[15]), .B(a[200]), .Z(n16111) );
  XNOR U16477 ( .A(n16112), .B(n16111), .Z(n16113) );
  XNOR U16478 ( .A(n16114), .B(n16113), .Z(n16132) );
  NAND U16479 ( .A(n33), .B(n16067), .Z(n16069) );
  XOR U16480 ( .A(b[5]), .B(a[212]), .Z(n16123) );
  NAND U16481 ( .A(n19342), .B(n16123), .Z(n16068) );
  AND U16482 ( .A(n16069), .B(n16068), .Z(n16156) );
  NAND U16483 ( .A(n34), .B(n16070), .Z(n16072) );
  XOR U16484 ( .A(b[7]), .B(a[210]), .Z(n16126) );
  NAND U16485 ( .A(n19486), .B(n16126), .Z(n16071) );
  AND U16486 ( .A(n16072), .B(n16071), .Z(n16154) );
  NAND U16487 ( .A(n31), .B(n16073), .Z(n16075) );
  XOR U16488 ( .A(b[3]), .B(a[214]), .Z(n16129) );
  NAND U16489 ( .A(n32), .B(n16129), .Z(n16074) );
  NAND U16490 ( .A(n16075), .B(n16074), .Z(n16153) );
  XNOR U16491 ( .A(n16154), .B(n16153), .Z(n16155) );
  XOR U16492 ( .A(n16156), .B(n16155), .Z(n16133) );
  XOR U16493 ( .A(n16132), .B(n16133), .Z(n16135) );
  XOR U16494 ( .A(n16134), .B(n16135), .Z(n16106) );
  NANDN U16495 ( .A(n16077), .B(n16076), .Z(n16081) );
  OR U16496 ( .A(n16079), .B(n16078), .Z(n16080) );
  AND U16497 ( .A(n16081), .B(n16080), .Z(n16105) );
  XNOR U16498 ( .A(n16106), .B(n16105), .Z(n16107) );
  XOR U16499 ( .A(n16108), .B(n16107), .Z(n16166) );
  NANDN U16500 ( .A(n16083), .B(n16082), .Z(n16087) );
  NANDN U16501 ( .A(n16085), .B(n16084), .Z(n16086) );
  AND U16502 ( .A(n16087), .B(n16086), .Z(n16165) );
  XNOR U16503 ( .A(n16166), .B(n16165), .Z(n16167) );
  XOR U16504 ( .A(n16168), .B(n16167), .Z(n16100) );
  NANDN U16505 ( .A(n16089), .B(n16088), .Z(n16093) );
  NAND U16506 ( .A(n16091), .B(n16090), .Z(n16092) );
  AND U16507 ( .A(n16093), .B(n16092), .Z(n16099) );
  XNOR U16508 ( .A(n16100), .B(n16099), .Z(n16101) );
  XNOR U16509 ( .A(n16102), .B(n16101), .Z(n16171) );
  XNOR U16510 ( .A(sreg[456]), .B(n16171), .Z(n16173) );
  NANDN U16511 ( .A(sreg[455]), .B(n16094), .Z(n16098) );
  NAND U16512 ( .A(n16096), .B(n16095), .Z(n16097) );
  NAND U16513 ( .A(n16098), .B(n16097), .Z(n16172) );
  XNOR U16514 ( .A(n16173), .B(n16172), .Z(c[456]) );
  NANDN U16515 ( .A(n16100), .B(n16099), .Z(n16104) );
  NANDN U16516 ( .A(n16102), .B(n16101), .Z(n16103) );
  AND U16517 ( .A(n16104), .B(n16103), .Z(n16179) );
  NANDN U16518 ( .A(n16106), .B(n16105), .Z(n16110) );
  NAND U16519 ( .A(n16108), .B(n16107), .Z(n16109) );
  AND U16520 ( .A(n16110), .B(n16109), .Z(n16245) );
  NANDN U16521 ( .A(n16112), .B(n16111), .Z(n16116) );
  NANDN U16522 ( .A(n16114), .B(n16113), .Z(n16115) );
  AND U16523 ( .A(n16116), .B(n16115), .Z(n16211) );
  NAND U16524 ( .A(b[0]), .B(a[217]), .Z(n16117) );
  XNOR U16525 ( .A(b[1]), .B(n16117), .Z(n16119) );
  NANDN U16526 ( .A(b[0]), .B(a[216]), .Z(n16118) );
  NAND U16527 ( .A(n16119), .B(n16118), .Z(n16191) );
  NAND U16528 ( .A(n19808), .B(n16120), .Z(n16122) );
  XOR U16529 ( .A(b[13]), .B(a[205]), .Z(n16194) );
  NAND U16530 ( .A(n19768), .B(n16194), .Z(n16121) );
  AND U16531 ( .A(n16122), .B(n16121), .Z(n16189) );
  AND U16532 ( .A(b[15]), .B(a[201]), .Z(n16188) );
  XNOR U16533 ( .A(n16189), .B(n16188), .Z(n16190) );
  XNOR U16534 ( .A(n16191), .B(n16190), .Z(n16209) );
  NAND U16535 ( .A(n33), .B(n16123), .Z(n16125) );
  XOR U16536 ( .A(b[5]), .B(a[213]), .Z(n16200) );
  NAND U16537 ( .A(n19342), .B(n16200), .Z(n16124) );
  AND U16538 ( .A(n16125), .B(n16124), .Z(n16233) );
  NAND U16539 ( .A(n34), .B(n16126), .Z(n16128) );
  XOR U16540 ( .A(b[7]), .B(a[211]), .Z(n16203) );
  NAND U16541 ( .A(n19486), .B(n16203), .Z(n16127) );
  AND U16542 ( .A(n16128), .B(n16127), .Z(n16231) );
  NAND U16543 ( .A(n31), .B(n16129), .Z(n16131) );
  XOR U16544 ( .A(b[3]), .B(a[215]), .Z(n16206) );
  NAND U16545 ( .A(n32), .B(n16206), .Z(n16130) );
  NAND U16546 ( .A(n16131), .B(n16130), .Z(n16230) );
  XNOR U16547 ( .A(n16231), .B(n16230), .Z(n16232) );
  XOR U16548 ( .A(n16233), .B(n16232), .Z(n16210) );
  XOR U16549 ( .A(n16209), .B(n16210), .Z(n16212) );
  XOR U16550 ( .A(n16211), .B(n16212), .Z(n16183) );
  NANDN U16551 ( .A(n16133), .B(n16132), .Z(n16137) );
  OR U16552 ( .A(n16135), .B(n16134), .Z(n16136) );
  AND U16553 ( .A(n16137), .B(n16136), .Z(n16182) );
  XNOR U16554 ( .A(n16183), .B(n16182), .Z(n16185) );
  NAND U16555 ( .A(n16138), .B(n19724), .Z(n16140) );
  XOR U16556 ( .A(b[11]), .B(a[207]), .Z(n16215) );
  NAND U16557 ( .A(n19692), .B(n16215), .Z(n16139) );
  AND U16558 ( .A(n16140), .B(n16139), .Z(n16226) );
  NAND U16559 ( .A(n19838), .B(n16141), .Z(n16143) );
  XOR U16560 ( .A(b[15]), .B(a[203]), .Z(n16218) );
  NAND U16561 ( .A(n19805), .B(n16218), .Z(n16142) );
  AND U16562 ( .A(n16143), .B(n16142), .Z(n16225) );
  NAND U16563 ( .A(n35), .B(n16144), .Z(n16146) );
  XOR U16564 ( .A(b[9]), .B(a[209]), .Z(n16221) );
  NAND U16565 ( .A(n19598), .B(n16221), .Z(n16145) );
  NAND U16566 ( .A(n16146), .B(n16145), .Z(n16224) );
  XOR U16567 ( .A(n16225), .B(n16224), .Z(n16227) );
  XOR U16568 ( .A(n16226), .B(n16227), .Z(n16237) );
  NANDN U16569 ( .A(n16148), .B(n16147), .Z(n16152) );
  OR U16570 ( .A(n16150), .B(n16149), .Z(n16151) );
  AND U16571 ( .A(n16152), .B(n16151), .Z(n16236) );
  XNOR U16572 ( .A(n16237), .B(n16236), .Z(n16238) );
  NANDN U16573 ( .A(n16154), .B(n16153), .Z(n16158) );
  NANDN U16574 ( .A(n16156), .B(n16155), .Z(n16157) );
  NAND U16575 ( .A(n16158), .B(n16157), .Z(n16239) );
  XNOR U16576 ( .A(n16238), .B(n16239), .Z(n16184) );
  XOR U16577 ( .A(n16185), .B(n16184), .Z(n16243) );
  NANDN U16578 ( .A(n16160), .B(n16159), .Z(n16164) );
  NANDN U16579 ( .A(n16162), .B(n16161), .Z(n16163) );
  AND U16580 ( .A(n16164), .B(n16163), .Z(n16242) );
  XNOR U16581 ( .A(n16243), .B(n16242), .Z(n16244) );
  XOR U16582 ( .A(n16245), .B(n16244), .Z(n16177) );
  NANDN U16583 ( .A(n16166), .B(n16165), .Z(n16170) );
  NAND U16584 ( .A(n16168), .B(n16167), .Z(n16169) );
  AND U16585 ( .A(n16170), .B(n16169), .Z(n16176) );
  XNOR U16586 ( .A(n16177), .B(n16176), .Z(n16178) );
  XNOR U16587 ( .A(n16179), .B(n16178), .Z(n16248) );
  XNOR U16588 ( .A(sreg[457]), .B(n16248), .Z(n16250) );
  NANDN U16589 ( .A(sreg[456]), .B(n16171), .Z(n16175) );
  NAND U16590 ( .A(n16173), .B(n16172), .Z(n16174) );
  NAND U16591 ( .A(n16175), .B(n16174), .Z(n16249) );
  XNOR U16592 ( .A(n16250), .B(n16249), .Z(c[457]) );
  NANDN U16593 ( .A(n16177), .B(n16176), .Z(n16181) );
  NANDN U16594 ( .A(n16179), .B(n16178), .Z(n16180) );
  AND U16595 ( .A(n16181), .B(n16180), .Z(n16256) );
  NANDN U16596 ( .A(n16183), .B(n16182), .Z(n16187) );
  NAND U16597 ( .A(n16185), .B(n16184), .Z(n16186) );
  AND U16598 ( .A(n16187), .B(n16186), .Z(n16322) );
  NANDN U16599 ( .A(n16189), .B(n16188), .Z(n16193) );
  NANDN U16600 ( .A(n16191), .B(n16190), .Z(n16192) );
  AND U16601 ( .A(n16193), .B(n16192), .Z(n16288) );
  NAND U16602 ( .A(n19808), .B(n16194), .Z(n16196) );
  XOR U16603 ( .A(b[13]), .B(a[206]), .Z(n16271) );
  NAND U16604 ( .A(n19768), .B(n16271), .Z(n16195) );
  AND U16605 ( .A(n16196), .B(n16195), .Z(n16266) );
  AND U16606 ( .A(b[15]), .B(a[202]), .Z(n16265) );
  XNOR U16607 ( .A(n16266), .B(n16265), .Z(n16267) );
  NAND U16608 ( .A(b[0]), .B(a[218]), .Z(n16197) );
  XNOR U16609 ( .A(b[1]), .B(n16197), .Z(n16199) );
  NANDN U16610 ( .A(b[0]), .B(a[217]), .Z(n16198) );
  NAND U16611 ( .A(n16199), .B(n16198), .Z(n16268) );
  XNOR U16612 ( .A(n16267), .B(n16268), .Z(n16286) );
  NAND U16613 ( .A(n33), .B(n16200), .Z(n16202) );
  XOR U16614 ( .A(b[5]), .B(a[214]), .Z(n16277) );
  NAND U16615 ( .A(n19342), .B(n16277), .Z(n16201) );
  AND U16616 ( .A(n16202), .B(n16201), .Z(n16310) );
  NAND U16617 ( .A(n34), .B(n16203), .Z(n16205) );
  XOR U16618 ( .A(b[7]), .B(a[212]), .Z(n16280) );
  NAND U16619 ( .A(n19486), .B(n16280), .Z(n16204) );
  AND U16620 ( .A(n16205), .B(n16204), .Z(n16308) );
  NAND U16621 ( .A(n31), .B(n16206), .Z(n16208) );
  XOR U16622 ( .A(b[3]), .B(a[216]), .Z(n16283) );
  NAND U16623 ( .A(n32), .B(n16283), .Z(n16207) );
  NAND U16624 ( .A(n16208), .B(n16207), .Z(n16307) );
  XNOR U16625 ( .A(n16308), .B(n16307), .Z(n16309) );
  XOR U16626 ( .A(n16310), .B(n16309), .Z(n16287) );
  XOR U16627 ( .A(n16286), .B(n16287), .Z(n16289) );
  XOR U16628 ( .A(n16288), .B(n16289), .Z(n16260) );
  NANDN U16629 ( .A(n16210), .B(n16209), .Z(n16214) );
  OR U16630 ( .A(n16212), .B(n16211), .Z(n16213) );
  AND U16631 ( .A(n16214), .B(n16213), .Z(n16259) );
  XNOR U16632 ( .A(n16260), .B(n16259), .Z(n16262) );
  NAND U16633 ( .A(n16215), .B(n19724), .Z(n16217) );
  XOR U16634 ( .A(b[11]), .B(a[208]), .Z(n16292) );
  NAND U16635 ( .A(n19692), .B(n16292), .Z(n16216) );
  AND U16636 ( .A(n16217), .B(n16216), .Z(n16303) );
  NAND U16637 ( .A(n19838), .B(n16218), .Z(n16220) );
  XOR U16638 ( .A(b[15]), .B(a[204]), .Z(n16295) );
  NAND U16639 ( .A(n19805), .B(n16295), .Z(n16219) );
  AND U16640 ( .A(n16220), .B(n16219), .Z(n16302) );
  NAND U16641 ( .A(n35), .B(n16221), .Z(n16223) );
  XOR U16642 ( .A(b[9]), .B(a[210]), .Z(n16298) );
  NAND U16643 ( .A(n19598), .B(n16298), .Z(n16222) );
  NAND U16644 ( .A(n16223), .B(n16222), .Z(n16301) );
  XOR U16645 ( .A(n16302), .B(n16301), .Z(n16304) );
  XOR U16646 ( .A(n16303), .B(n16304), .Z(n16314) );
  NANDN U16647 ( .A(n16225), .B(n16224), .Z(n16229) );
  OR U16648 ( .A(n16227), .B(n16226), .Z(n16228) );
  AND U16649 ( .A(n16229), .B(n16228), .Z(n16313) );
  XNOR U16650 ( .A(n16314), .B(n16313), .Z(n16315) );
  NANDN U16651 ( .A(n16231), .B(n16230), .Z(n16235) );
  NANDN U16652 ( .A(n16233), .B(n16232), .Z(n16234) );
  NAND U16653 ( .A(n16235), .B(n16234), .Z(n16316) );
  XNOR U16654 ( .A(n16315), .B(n16316), .Z(n16261) );
  XOR U16655 ( .A(n16262), .B(n16261), .Z(n16320) );
  NANDN U16656 ( .A(n16237), .B(n16236), .Z(n16241) );
  NANDN U16657 ( .A(n16239), .B(n16238), .Z(n16240) );
  AND U16658 ( .A(n16241), .B(n16240), .Z(n16319) );
  XNOR U16659 ( .A(n16320), .B(n16319), .Z(n16321) );
  XOR U16660 ( .A(n16322), .B(n16321), .Z(n16254) );
  NANDN U16661 ( .A(n16243), .B(n16242), .Z(n16247) );
  NAND U16662 ( .A(n16245), .B(n16244), .Z(n16246) );
  AND U16663 ( .A(n16247), .B(n16246), .Z(n16253) );
  XNOR U16664 ( .A(n16254), .B(n16253), .Z(n16255) );
  XNOR U16665 ( .A(n16256), .B(n16255), .Z(n16325) );
  XNOR U16666 ( .A(sreg[458]), .B(n16325), .Z(n16327) );
  NANDN U16667 ( .A(sreg[457]), .B(n16248), .Z(n16252) );
  NAND U16668 ( .A(n16250), .B(n16249), .Z(n16251) );
  NAND U16669 ( .A(n16252), .B(n16251), .Z(n16326) );
  XNOR U16670 ( .A(n16327), .B(n16326), .Z(c[458]) );
  NANDN U16671 ( .A(n16254), .B(n16253), .Z(n16258) );
  NANDN U16672 ( .A(n16256), .B(n16255), .Z(n16257) );
  AND U16673 ( .A(n16258), .B(n16257), .Z(n16333) );
  NANDN U16674 ( .A(n16260), .B(n16259), .Z(n16264) );
  NAND U16675 ( .A(n16262), .B(n16261), .Z(n16263) );
  AND U16676 ( .A(n16264), .B(n16263), .Z(n16399) );
  NANDN U16677 ( .A(n16266), .B(n16265), .Z(n16270) );
  NANDN U16678 ( .A(n16268), .B(n16267), .Z(n16269) );
  AND U16679 ( .A(n16270), .B(n16269), .Z(n16365) );
  NAND U16680 ( .A(n19808), .B(n16271), .Z(n16273) );
  XOR U16681 ( .A(b[13]), .B(a[207]), .Z(n16351) );
  NAND U16682 ( .A(n19768), .B(n16351), .Z(n16272) );
  AND U16683 ( .A(n16273), .B(n16272), .Z(n16343) );
  AND U16684 ( .A(b[15]), .B(a[203]), .Z(n16342) );
  XNOR U16685 ( .A(n16343), .B(n16342), .Z(n16344) );
  NAND U16686 ( .A(b[0]), .B(a[219]), .Z(n16274) );
  XNOR U16687 ( .A(b[1]), .B(n16274), .Z(n16276) );
  NANDN U16688 ( .A(b[0]), .B(a[218]), .Z(n16275) );
  NAND U16689 ( .A(n16276), .B(n16275), .Z(n16345) );
  XNOR U16690 ( .A(n16344), .B(n16345), .Z(n16363) );
  NAND U16691 ( .A(n33), .B(n16277), .Z(n16279) );
  XOR U16692 ( .A(b[5]), .B(a[215]), .Z(n16354) );
  NAND U16693 ( .A(n19342), .B(n16354), .Z(n16278) );
  AND U16694 ( .A(n16279), .B(n16278), .Z(n16387) );
  NAND U16695 ( .A(n34), .B(n16280), .Z(n16282) );
  XOR U16696 ( .A(b[7]), .B(a[213]), .Z(n16357) );
  NAND U16697 ( .A(n19486), .B(n16357), .Z(n16281) );
  AND U16698 ( .A(n16282), .B(n16281), .Z(n16385) );
  NAND U16699 ( .A(n31), .B(n16283), .Z(n16285) );
  XOR U16700 ( .A(b[3]), .B(a[217]), .Z(n16360) );
  NAND U16701 ( .A(n32), .B(n16360), .Z(n16284) );
  NAND U16702 ( .A(n16285), .B(n16284), .Z(n16384) );
  XNOR U16703 ( .A(n16385), .B(n16384), .Z(n16386) );
  XOR U16704 ( .A(n16387), .B(n16386), .Z(n16364) );
  XOR U16705 ( .A(n16363), .B(n16364), .Z(n16366) );
  XOR U16706 ( .A(n16365), .B(n16366), .Z(n16337) );
  NANDN U16707 ( .A(n16287), .B(n16286), .Z(n16291) );
  OR U16708 ( .A(n16289), .B(n16288), .Z(n16290) );
  AND U16709 ( .A(n16291), .B(n16290), .Z(n16336) );
  XNOR U16710 ( .A(n16337), .B(n16336), .Z(n16339) );
  NAND U16711 ( .A(n16292), .B(n19724), .Z(n16294) );
  XOR U16712 ( .A(b[11]), .B(a[209]), .Z(n16369) );
  NAND U16713 ( .A(n19692), .B(n16369), .Z(n16293) );
  AND U16714 ( .A(n16294), .B(n16293), .Z(n16380) );
  NAND U16715 ( .A(n19838), .B(n16295), .Z(n16297) );
  XOR U16716 ( .A(b[15]), .B(a[205]), .Z(n16372) );
  NAND U16717 ( .A(n19805), .B(n16372), .Z(n16296) );
  AND U16718 ( .A(n16297), .B(n16296), .Z(n16379) );
  NAND U16719 ( .A(n35), .B(n16298), .Z(n16300) );
  XOR U16720 ( .A(b[9]), .B(a[211]), .Z(n16375) );
  NAND U16721 ( .A(n19598), .B(n16375), .Z(n16299) );
  NAND U16722 ( .A(n16300), .B(n16299), .Z(n16378) );
  XOR U16723 ( .A(n16379), .B(n16378), .Z(n16381) );
  XOR U16724 ( .A(n16380), .B(n16381), .Z(n16391) );
  NANDN U16725 ( .A(n16302), .B(n16301), .Z(n16306) );
  OR U16726 ( .A(n16304), .B(n16303), .Z(n16305) );
  AND U16727 ( .A(n16306), .B(n16305), .Z(n16390) );
  XNOR U16728 ( .A(n16391), .B(n16390), .Z(n16392) );
  NANDN U16729 ( .A(n16308), .B(n16307), .Z(n16312) );
  NANDN U16730 ( .A(n16310), .B(n16309), .Z(n16311) );
  NAND U16731 ( .A(n16312), .B(n16311), .Z(n16393) );
  XNOR U16732 ( .A(n16392), .B(n16393), .Z(n16338) );
  XOR U16733 ( .A(n16339), .B(n16338), .Z(n16397) );
  NANDN U16734 ( .A(n16314), .B(n16313), .Z(n16318) );
  NANDN U16735 ( .A(n16316), .B(n16315), .Z(n16317) );
  AND U16736 ( .A(n16318), .B(n16317), .Z(n16396) );
  XNOR U16737 ( .A(n16397), .B(n16396), .Z(n16398) );
  XOR U16738 ( .A(n16399), .B(n16398), .Z(n16331) );
  NANDN U16739 ( .A(n16320), .B(n16319), .Z(n16324) );
  NAND U16740 ( .A(n16322), .B(n16321), .Z(n16323) );
  AND U16741 ( .A(n16324), .B(n16323), .Z(n16330) );
  XNOR U16742 ( .A(n16331), .B(n16330), .Z(n16332) );
  XNOR U16743 ( .A(n16333), .B(n16332), .Z(n16402) );
  XNOR U16744 ( .A(sreg[459]), .B(n16402), .Z(n16404) );
  NANDN U16745 ( .A(sreg[458]), .B(n16325), .Z(n16329) );
  NAND U16746 ( .A(n16327), .B(n16326), .Z(n16328) );
  NAND U16747 ( .A(n16329), .B(n16328), .Z(n16403) );
  XNOR U16748 ( .A(n16404), .B(n16403), .Z(c[459]) );
  NANDN U16749 ( .A(n16331), .B(n16330), .Z(n16335) );
  NANDN U16750 ( .A(n16333), .B(n16332), .Z(n16334) );
  AND U16751 ( .A(n16335), .B(n16334), .Z(n16410) );
  NANDN U16752 ( .A(n16337), .B(n16336), .Z(n16341) );
  NAND U16753 ( .A(n16339), .B(n16338), .Z(n16340) );
  AND U16754 ( .A(n16341), .B(n16340), .Z(n16476) );
  NANDN U16755 ( .A(n16343), .B(n16342), .Z(n16347) );
  NANDN U16756 ( .A(n16345), .B(n16344), .Z(n16346) );
  AND U16757 ( .A(n16347), .B(n16346), .Z(n16442) );
  NAND U16758 ( .A(b[0]), .B(a[220]), .Z(n16348) );
  XNOR U16759 ( .A(b[1]), .B(n16348), .Z(n16350) );
  NANDN U16760 ( .A(b[0]), .B(a[219]), .Z(n16349) );
  NAND U16761 ( .A(n16350), .B(n16349), .Z(n16422) );
  NAND U16762 ( .A(n19808), .B(n16351), .Z(n16353) );
  XOR U16763 ( .A(b[13]), .B(a[208]), .Z(n16425) );
  NAND U16764 ( .A(n19768), .B(n16425), .Z(n16352) );
  AND U16765 ( .A(n16353), .B(n16352), .Z(n16420) );
  AND U16766 ( .A(b[15]), .B(a[204]), .Z(n16419) );
  XNOR U16767 ( .A(n16420), .B(n16419), .Z(n16421) );
  XNOR U16768 ( .A(n16422), .B(n16421), .Z(n16440) );
  NAND U16769 ( .A(n33), .B(n16354), .Z(n16356) );
  XOR U16770 ( .A(b[5]), .B(a[216]), .Z(n16431) );
  NAND U16771 ( .A(n19342), .B(n16431), .Z(n16355) );
  AND U16772 ( .A(n16356), .B(n16355), .Z(n16464) );
  NAND U16773 ( .A(n34), .B(n16357), .Z(n16359) );
  XOR U16774 ( .A(b[7]), .B(a[214]), .Z(n16434) );
  NAND U16775 ( .A(n19486), .B(n16434), .Z(n16358) );
  AND U16776 ( .A(n16359), .B(n16358), .Z(n16462) );
  NAND U16777 ( .A(n31), .B(n16360), .Z(n16362) );
  XOR U16778 ( .A(b[3]), .B(a[218]), .Z(n16437) );
  NAND U16779 ( .A(n32), .B(n16437), .Z(n16361) );
  NAND U16780 ( .A(n16362), .B(n16361), .Z(n16461) );
  XNOR U16781 ( .A(n16462), .B(n16461), .Z(n16463) );
  XOR U16782 ( .A(n16464), .B(n16463), .Z(n16441) );
  XOR U16783 ( .A(n16440), .B(n16441), .Z(n16443) );
  XOR U16784 ( .A(n16442), .B(n16443), .Z(n16414) );
  NANDN U16785 ( .A(n16364), .B(n16363), .Z(n16368) );
  OR U16786 ( .A(n16366), .B(n16365), .Z(n16367) );
  AND U16787 ( .A(n16368), .B(n16367), .Z(n16413) );
  XNOR U16788 ( .A(n16414), .B(n16413), .Z(n16416) );
  NAND U16789 ( .A(n16369), .B(n19724), .Z(n16371) );
  XOR U16790 ( .A(b[11]), .B(a[210]), .Z(n16446) );
  NAND U16791 ( .A(n19692), .B(n16446), .Z(n16370) );
  AND U16792 ( .A(n16371), .B(n16370), .Z(n16457) );
  NAND U16793 ( .A(n19838), .B(n16372), .Z(n16374) );
  XOR U16794 ( .A(b[15]), .B(a[206]), .Z(n16449) );
  NAND U16795 ( .A(n19805), .B(n16449), .Z(n16373) );
  AND U16796 ( .A(n16374), .B(n16373), .Z(n16456) );
  NAND U16797 ( .A(n35), .B(n16375), .Z(n16377) );
  XOR U16798 ( .A(b[9]), .B(a[212]), .Z(n16452) );
  NAND U16799 ( .A(n19598), .B(n16452), .Z(n16376) );
  NAND U16800 ( .A(n16377), .B(n16376), .Z(n16455) );
  XOR U16801 ( .A(n16456), .B(n16455), .Z(n16458) );
  XOR U16802 ( .A(n16457), .B(n16458), .Z(n16468) );
  NANDN U16803 ( .A(n16379), .B(n16378), .Z(n16383) );
  OR U16804 ( .A(n16381), .B(n16380), .Z(n16382) );
  AND U16805 ( .A(n16383), .B(n16382), .Z(n16467) );
  XNOR U16806 ( .A(n16468), .B(n16467), .Z(n16469) );
  NANDN U16807 ( .A(n16385), .B(n16384), .Z(n16389) );
  NANDN U16808 ( .A(n16387), .B(n16386), .Z(n16388) );
  NAND U16809 ( .A(n16389), .B(n16388), .Z(n16470) );
  XNOR U16810 ( .A(n16469), .B(n16470), .Z(n16415) );
  XOR U16811 ( .A(n16416), .B(n16415), .Z(n16474) );
  NANDN U16812 ( .A(n16391), .B(n16390), .Z(n16395) );
  NANDN U16813 ( .A(n16393), .B(n16392), .Z(n16394) );
  AND U16814 ( .A(n16395), .B(n16394), .Z(n16473) );
  XNOR U16815 ( .A(n16474), .B(n16473), .Z(n16475) );
  XOR U16816 ( .A(n16476), .B(n16475), .Z(n16408) );
  NANDN U16817 ( .A(n16397), .B(n16396), .Z(n16401) );
  NAND U16818 ( .A(n16399), .B(n16398), .Z(n16400) );
  AND U16819 ( .A(n16401), .B(n16400), .Z(n16407) );
  XNOR U16820 ( .A(n16408), .B(n16407), .Z(n16409) );
  XNOR U16821 ( .A(n16410), .B(n16409), .Z(n16479) );
  XNOR U16822 ( .A(sreg[460]), .B(n16479), .Z(n16481) );
  NANDN U16823 ( .A(sreg[459]), .B(n16402), .Z(n16406) );
  NAND U16824 ( .A(n16404), .B(n16403), .Z(n16405) );
  NAND U16825 ( .A(n16406), .B(n16405), .Z(n16480) );
  XNOR U16826 ( .A(n16481), .B(n16480), .Z(c[460]) );
  NANDN U16827 ( .A(n16408), .B(n16407), .Z(n16412) );
  NANDN U16828 ( .A(n16410), .B(n16409), .Z(n16411) );
  AND U16829 ( .A(n16412), .B(n16411), .Z(n16487) );
  NANDN U16830 ( .A(n16414), .B(n16413), .Z(n16418) );
  NAND U16831 ( .A(n16416), .B(n16415), .Z(n16417) );
  AND U16832 ( .A(n16418), .B(n16417), .Z(n16553) );
  NANDN U16833 ( .A(n16420), .B(n16419), .Z(n16424) );
  NANDN U16834 ( .A(n16422), .B(n16421), .Z(n16423) );
  AND U16835 ( .A(n16424), .B(n16423), .Z(n16519) );
  NAND U16836 ( .A(n19808), .B(n16425), .Z(n16427) );
  XOR U16837 ( .A(b[13]), .B(a[209]), .Z(n16505) );
  NAND U16838 ( .A(n19768), .B(n16505), .Z(n16426) );
  AND U16839 ( .A(n16427), .B(n16426), .Z(n16497) );
  AND U16840 ( .A(b[15]), .B(a[205]), .Z(n16496) );
  XNOR U16841 ( .A(n16497), .B(n16496), .Z(n16498) );
  NAND U16842 ( .A(b[0]), .B(a[221]), .Z(n16428) );
  XNOR U16843 ( .A(b[1]), .B(n16428), .Z(n16430) );
  NANDN U16844 ( .A(b[0]), .B(a[220]), .Z(n16429) );
  NAND U16845 ( .A(n16430), .B(n16429), .Z(n16499) );
  XNOR U16846 ( .A(n16498), .B(n16499), .Z(n16517) );
  NAND U16847 ( .A(n33), .B(n16431), .Z(n16433) );
  XOR U16848 ( .A(b[5]), .B(a[217]), .Z(n16508) );
  NAND U16849 ( .A(n19342), .B(n16508), .Z(n16432) );
  AND U16850 ( .A(n16433), .B(n16432), .Z(n16541) );
  NAND U16851 ( .A(n34), .B(n16434), .Z(n16436) );
  XOR U16852 ( .A(b[7]), .B(a[215]), .Z(n16511) );
  NAND U16853 ( .A(n19486), .B(n16511), .Z(n16435) );
  AND U16854 ( .A(n16436), .B(n16435), .Z(n16539) );
  NAND U16855 ( .A(n31), .B(n16437), .Z(n16439) );
  XOR U16856 ( .A(b[3]), .B(a[219]), .Z(n16514) );
  NAND U16857 ( .A(n32), .B(n16514), .Z(n16438) );
  NAND U16858 ( .A(n16439), .B(n16438), .Z(n16538) );
  XNOR U16859 ( .A(n16539), .B(n16538), .Z(n16540) );
  XOR U16860 ( .A(n16541), .B(n16540), .Z(n16518) );
  XOR U16861 ( .A(n16517), .B(n16518), .Z(n16520) );
  XOR U16862 ( .A(n16519), .B(n16520), .Z(n16491) );
  NANDN U16863 ( .A(n16441), .B(n16440), .Z(n16445) );
  OR U16864 ( .A(n16443), .B(n16442), .Z(n16444) );
  AND U16865 ( .A(n16445), .B(n16444), .Z(n16490) );
  XNOR U16866 ( .A(n16491), .B(n16490), .Z(n16493) );
  NAND U16867 ( .A(n16446), .B(n19724), .Z(n16448) );
  XOR U16868 ( .A(b[11]), .B(a[211]), .Z(n16523) );
  NAND U16869 ( .A(n19692), .B(n16523), .Z(n16447) );
  AND U16870 ( .A(n16448), .B(n16447), .Z(n16534) );
  NAND U16871 ( .A(n19838), .B(n16449), .Z(n16451) );
  XOR U16872 ( .A(b[15]), .B(a[207]), .Z(n16526) );
  NAND U16873 ( .A(n19805), .B(n16526), .Z(n16450) );
  AND U16874 ( .A(n16451), .B(n16450), .Z(n16533) );
  NAND U16875 ( .A(n35), .B(n16452), .Z(n16454) );
  XOR U16876 ( .A(b[9]), .B(a[213]), .Z(n16529) );
  NAND U16877 ( .A(n19598), .B(n16529), .Z(n16453) );
  NAND U16878 ( .A(n16454), .B(n16453), .Z(n16532) );
  XOR U16879 ( .A(n16533), .B(n16532), .Z(n16535) );
  XOR U16880 ( .A(n16534), .B(n16535), .Z(n16545) );
  NANDN U16881 ( .A(n16456), .B(n16455), .Z(n16460) );
  OR U16882 ( .A(n16458), .B(n16457), .Z(n16459) );
  AND U16883 ( .A(n16460), .B(n16459), .Z(n16544) );
  XNOR U16884 ( .A(n16545), .B(n16544), .Z(n16546) );
  NANDN U16885 ( .A(n16462), .B(n16461), .Z(n16466) );
  NANDN U16886 ( .A(n16464), .B(n16463), .Z(n16465) );
  NAND U16887 ( .A(n16466), .B(n16465), .Z(n16547) );
  XNOR U16888 ( .A(n16546), .B(n16547), .Z(n16492) );
  XOR U16889 ( .A(n16493), .B(n16492), .Z(n16551) );
  NANDN U16890 ( .A(n16468), .B(n16467), .Z(n16472) );
  NANDN U16891 ( .A(n16470), .B(n16469), .Z(n16471) );
  AND U16892 ( .A(n16472), .B(n16471), .Z(n16550) );
  XNOR U16893 ( .A(n16551), .B(n16550), .Z(n16552) );
  XOR U16894 ( .A(n16553), .B(n16552), .Z(n16485) );
  NANDN U16895 ( .A(n16474), .B(n16473), .Z(n16478) );
  NAND U16896 ( .A(n16476), .B(n16475), .Z(n16477) );
  AND U16897 ( .A(n16478), .B(n16477), .Z(n16484) );
  XNOR U16898 ( .A(n16485), .B(n16484), .Z(n16486) );
  XNOR U16899 ( .A(n16487), .B(n16486), .Z(n16556) );
  XNOR U16900 ( .A(sreg[461]), .B(n16556), .Z(n16558) );
  NANDN U16901 ( .A(sreg[460]), .B(n16479), .Z(n16483) );
  NAND U16902 ( .A(n16481), .B(n16480), .Z(n16482) );
  NAND U16903 ( .A(n16483), .B(n16482), .Z(n16557) );
  XNOR U16904 ( .A(n16558), .B(n16557), .Z(c[461]) );
  NANDN U16905 ( .A(n16485), .B(n16484), .Z(n16489) );
  NANDN U16906 ( .A(n16487), .B(n16486), .Z(n16488) );
  AND U16907 ( .A(n16489), .B(n16488), .Z(n16564) );
  NANDN U16908 ( .A(n16491), .B(n16490), .Z(n16495) );
  NAND U16909 ( .A(n16493), .B(n16492), .Z(n16494) );
  AND U16910 ( .A(n16495), .B(n16494), .Z(n16630) );
  NANDN U16911 ( .A(n16497), .B(n16496), .Z(n16501) );
  NANDN U16912 ( .A(n16499), .B(n16498), .Z(n16500) );
  AND U16913 ( .A(n16501), .B(n16500), .Z(n16596) );
  NAND U16914 ( .A(b[0]), .B(a[222]), .Z(n16502) );
  XNOR U16915 ( .A(b[1]), .B(n16502), .Z(n16504) );
  NANDN U16916 ( .A(b[0]), .B(a[221]), .Z(n16503) );
  NAND U16917 ( .A(n16504), .B(n16503), .Z(n16576) );
  NAND U16918 ( .A(n19808), .B(n16505), .Z(n16507) );
  XOR U16919 ( .A(b[13]), .B(a[210]), .Z(n16579) );
  NAND U16920 ( .A(n19768), .B(n16579), .Z(n16506) );
  AND U16921 ( .A(n16507), .B(n16506), .Z(n16574) );
  AND U16922 ( .A(b[15]), .B(a[206]), .Z(n16573) );
  XNOR U16923 ( .A(n16574), .B(n16573), .Z(n16575) );
  XNOR U16924 ( .A(n16576), .B(n16575), .Z(n16594) );
  NAND U16925 ( .A(n33), .B(n16508), .Z(n16510) );
  XOR U16926 ( .A(b[5]), .B(a[218]), .Z(n16585) );
  NAND U16927 ( .A(n19342), .B(n16585), .Z(n16509) );
  AND U16928 ( .A(n16510), .B(n16509), .Z(n16618) );
  NAND U16929 ( .A(n34), .B(n16511), .Z(n16513) );
  XOR U16930 ( .A(b[7]), .B(a[216]), .Z(n16588) );
  NAND U16931 ( .A(n19486), .B(n16588), .Z(n16512) );
  AND U16932 ( .A(n16513), .B(n16512), .Z(n16616) );
  NAND U16933 ( .A(n31), .B(n16514), .Z(n16516) );
  XOR U16934 ( .A(b[3]), .B(a[220]), .Z(n16591) );
  NAND U16935 ( .A(n32), .B(n16591), .Z(n16515) );
  NAND U16936 ( .A(n16516), .B(n16515), .Z(n16615) );
  XNOR U16937 ( .A(n16616), .B(n16615), .Z(n16617) );
  XOR U16938 ( .A(n16618), .B(n16617), .Z(n16595) );
  XOR U16939 ( .A(n16594), .B(n16595), .Z(n16597) );
  XOR U16940 ( .A(n16596), .B(n16597), .Z(n16568) );
  NANDN U16941 ( .A(n16518), .B(n16517), .Z(n16522) );
  OR U16942 ( .A(n16520), .B(n16519), .Z(n16521) );
  AND U16943 ( .A(n16522), .B(n16521), .Z(n16567) );
  XNOR U16944 ( .A(n16568), .B(n16567), .Z(n16570) );
  NAND U16945 ( .A(n16523), .B(n19724), .Z(n16525) );
  XOR U16946 ( .A(b[11]), .B(a[212]), .Z(n16600) );
  NAND U16947 ( .A(n19692), .B(n16600), .Z(n16524) );
  AND U16948 ( .A(n16525), .B(n16524), .Z(n16611) );
  NAND U16949 ( .A(n19838), .B(n16526), .Z(n16528) );
  XOR U16950 ( .A(b[15]), .B(a[208]), .Z(n16603) );
  NAND U16951 ( .A(n19805), .B(n16603), .Z(n16527) );
  AND U16952 ( .A(n16528), .B(n16527), .Z(n16610) );
  NAND U16953 ( .A(n35), .B(n16529), .Z(n16531) );
  XOR U16954 ( .A(b[9]), .B(a[214]), .Z(n16606) );
  NAND U16955 ( .A(n19598), .B(n16606), .Z(n16530) );
  NAND U16956 ( .A(n16531), .B(n16530), .Z(n16609) );
  XOR U16957 ( .A(n16610), .B(n16609), .Z(n16612) );
  XOR U16958 ( .A(n16611), .B(n16612), .Z(n16622) );
  NANDN U16959 ( .A(n16533), .B(n16532), .Z(n16537) );
  OR U16960 ( .A(n16535), .B(n16534), .Z(n16536) );
  AND U16961 ( .A(n16537), .B(n16536), .Z(n16621) );
  XNOR U16962 ( .A(n16622), .B(n16621), .Z(n16623) );
  NANDN U16963 ( .A(n16539), .B(n16538), .Z(n16543) );
  NANDN U16964 ( .A(n16541), .B(n16540), .Z(n16542) );
  NAND U16965 ( .A(n16543), .B(n16542), .Z(n16624) );
  XNOR U16966 ( .A(n16623), .B(n16624), .Z(n16569) );
  XOR U16967 ( .A(n16570), .B(n16569), .Z(n16628) );
  NANDN U16968 ( .A(n16545), .B(n16544), .Z(n16549) );
  NANDN U16969 ( .A(n16547), .B(n16546), .Z(n16548) );
  AND U16970 ( .A(n16549), .B(n16548), .Z(n16627) );
  XNOR U16971 ( .A(n16628), .B(n16627), .Z(n16629) );
  XOR U16972 ( .A(n16630), .B(n16629), .Z(n16562) );
  NANDN U16973 ( .A(n16551), .B(n16550), .Z(n16555) );
  NAND U16974 ( .A(n16553), .B(n16552), .Z(n16554) );
  AND U16975 ( .A(n16555), .B(n16554), .Z(n16561) );
  XNOR U16976 ( .A(n16562), .B(n16561), .Z(n16563) );
  XNOR U16977 ( .A(n16564), .B(n16563), .Z(n16633) );
  XNOR U16978 ( .A(sreg[462]), .B(n16633), .Z(n16635) );
  NANDN U16979 ( .A(sreg[461]), .B(n16556), .Z(n16560) );
  NAND U16980 ( .A(n16558), .B(n16557), .Z(n16559) );
  NAND U16981 ( .A(n16560), .B(n16559), .Z(n16634) );
  XNOR U16982 ( .A(n16635), .B(n16634), .Z(c[462]) );
  NANDN U16983 ( .A(n16562), .B(n16561), .Z(n16566) );
  NANDN U16984 ( .A(n16564), .B(n16563), .Z(n16565) );
  AND U16985 ( .A(n16566), .B(n16565), .Z(n16641) );
  NANDN U16986 ( .A(n16568), .B(n16567), .Z(n16572) );
  NAND U16987 ( .A(n16570), .B(n16569), .Z(n16571) );
  AND U16988 ( .A(n16572), .B(n16571), .Z(n16707) );
  NANDN U16989 ( .A(n16574), .B(n16573), .Z(n16578) );
  NANDN U16990 ( .A(n16576), .B(n16575), .Z(n16577) );
  AND U16991 ( .A(n16578), .B(n16577), .Z(n16694) );
  NAND U16992 ( .A(n19808), .B(n16579), .Z(n16581) );
  XOR U16993 ( .A(b[13]), .B(a[211]), .Z(n16680) );
  NAND U16994 ( .A(n19768), .B(n16680), .Z(n16580) );
  AND U16995 ( .A(n16581), .B(n16580), .Z(n16672) );
  AND U16996 ( .A(b[15]), .B(a[207]), .Z(n16671) );
  XNOR U16997 ( .A(n16672), .B(n16671), .Z(n16673) );
  NAND U16998 ( .A(b[0]), .B(a[223]), .Z(n16582) );
  XNOR U16999 ( .A(b[1]), .B(n16582), .Z(n16584) );
  NANDN U17000 ( .A(b[0]), .B(a[222]), .Z(n16583) );
  NAND U17001 ( .A(n16584), .B(n16583), .Z(n16674) );
  XNOR U17002 ( .A(n16673), .B(n16674), .Z(n16692) );
  NAND U17003 ( .A(n33), .B(n16585), .Z(n16587) );
  XOR U17004 ( .A(b[5]), .B(a[219]), .Z(n16683) );
  NAND U17005 ( .A(n19342), .B(n16683), .Z(n16586) );
  AND U17006 ( .A(n16587), .B(n16586), .Z(n16668) );
  NAND U17007 ( .A(n34), .B(n16588), .Z(n16590) );
  XOR U17008 ( .A(b[7]), .B(a[217]), .Z(n16686) );
  NAND U17009 ( .A(n19486), .B(n16686), .Z(n16589) );
  AND U17010 ( .A(n16590), .B(n16589), .Z(n16666) );
  NAND U17011 ( .A(n31), .B(n16591), .Z(n16593) );
  XOR U17012 ( .A(b[3]), .B(a[221]), .Z(n16689) );
  NAND U17013 ( .A(n32), .B(n16689), .Z(n16592) );
  NAND U17014 ( .A(n16593), .B(n16592), .Z(n16665) );
  XNOR U17015 ( .A(n16666), .B(n16665), .Z(n16667) );
  XOR U17016 ( .A(n16668), .B(n16667), .Z(n16693) );
  XOR U17017 ( .A(n16692), .B(n16693), .Z(n16695) );
  XOR U17018 ( .A(n16694), .B(n16695), .Z(n16645) );
  NANDN U17019 ( .A(n16595), .B(n16594), .Z(n16599) );
  OR U17020 ( .A(n16597), .B(n16596), .Z(n16598) );
  AND U17021 ( .A(n16599), .B(n16598), .Z(n16644) );
  XNOR U17022 ( .A(n16645), .B(n16644), .Z(n16647) );
  NAND U17023 ( .A(n16600), .B(n19724), .Z(n16602) );
  XOR U17024 ( .A(b[11]), .B(a[213]), .Z(n16650) );
  NAND U17025 ( .A(n19692), .B(n16650), .Z(n16601) );
  AND U17026 ( .A(n16602), .B(n16601), .Z(n16661) );
  NAND U17027 ( .A(n19838), .B(n16603), .Z(n16605) );
  XOR U17028 ( .A(b[15]), .B(a[209]), .Z(n16653) );
  NAND U17029 ( .A(n19805), .B(n16653), .Z(n16604) );
  AND U17030 ( .A(n16605), .B(n16604), .Z(n16660) );
  NAND U17031 ( .A(n35), .B(n16606), .Z(n16608) );
  XOR U17032 ( .A(b[9]), .B(a[215]), .Z(n16656) );
  NAND U17033 ( .A(n19598), .B(n16656), .Z(n16607) );
  NAND U17034 ( .A(n16608), .B(n16607), .Z(n16659) );
  XOR U17035 ( .A(n16660), .B(n16659), .Z(n16662) );
  XOR U17036 ( .A(n16661), .B(n16662), .Z(n16699) );
  NANDN U17037 ( .A(n16610), .B(n16609), .Z(n16614) );
  OR U17038 ( .A(n16612), .B(n16611), .Z(n16613) );
  AND U17039 ( .A(n16614), .B(n16613), .Z(n16698) );
  XNOR U17040 ( .A(n16699), .B(n16698), .Z(n16700) );
  NANDN U17041 ( .A(n16616), .B(n16615), .Z(n16620) );
  NANDN U17042 ( .A(n16618), .B(n16617), .Z(n16619) );
  NAND U17043 ( .A(n16620), .B(n16619), .Z(n16701) );
  XNOR U17044 ( .A(n16700), .B(n16701), .Z(n16646) );
  XOR U17045 ( .A(n16647), .B(n16646), .Z(n16705) );
  NANDN U17046 ( .A(n16622), .B(n16621), .Z(n16626) );
  NANDN U17047 ( .A(n16624), .B(n16623), .Z(n16625) );
  AND U17048 ( .A(n16626), .B(n16625), .Z(n16704) );
  XNOR U17049 ( .A(n16705), .B(n16704), .Z(n16706) );
  XOR U17050 ( .A(n16707), .B(n16706), .Z(n16639) );
  NANDN U17051 ( .A(n16628), .B(n16627), .Z(n16632) );
  NAND U17052 ( .A(n16630), .B(n16629), .Z(n16631) );
  AND U17053 ( .A(n16632), .B(n16631), .Z(n16638) );
  XNOR U17054 ( .A(n16639), .B(n16638), .Z(n16640) );
  XNOR U17055 ( .A(n16641), .B(n16640), .Z(n16710) );
  XNOR U17056 ( .A(sreg[463]), .B(n16710), .Z(n16712) );
  NANDN U17057 ( .A(sreg[462]), .B(n16633), .Z(n16637) );
  NAND U17058 ( .A(n16635), .B(n16634), .Z(n16636) );
  NAND U17059 ( .A(n16637), .B(n16636), .Z(n16711) );
  XNOR U17060 ( .A(n16712), .B(n16711), .Z(c[463]) );
  NANDN U17061 ( .A(n16639), .B(n16638), .Z(n16643) );
  NANDN U17062 ( .A(n16641), .B(n16640), .Z(n16642) );
  AND U17063 ( .A(n16643), .B(n16642), .Z(n16718) );
  NANDN U17064 ( .A(n16645), .B(n16644), .Z(n16649) );
  NAND U17065 ( .A(n16647), .B(n16646), .Z(n16648) );
  AND U17066 ( .A(n16649), .B(n16648), .Z(n16784) );
  NAND U17067 ( .A(n16650), .B(n19724), .Z(n16652) );
  XOR U17068 ( .A(b[11]), .B(a[214]), .Z(n16754) );
  NAND U17069 ( .A(n19692), .B(n16754), .Z(n16651) );
  AND U17070 ( .A(n16652), .B(n16651), .Z(n16765) );
  NAND U17071 ( .A(n19838), .B(n16653), .Z(n16655) );
  XOR U17072 ( .A(b[15]), .B(a[210]), .Z(n16757) );
  NAND U17073 ( .A(n19805), .B(n16757), .Z(n16654) );
  AND U17074 ( .A(n16655), .B(n16654), .Z(n16764) );
  NAND U17075 ( .A(n35), .B(n16656), .Z(n16658) );
  XOR U17076 ( .A(b[9]), .B(a[216]), .Z(n16760) );
  NAND U17077 ( .A(n19598), .B(n16760), .Z(n16657) );
  NAND U17078 ( .A(n16658), .B(n16657), .Z(n16763) );
  XOR U17079 ( .A(n16764), .B(n16763), .Z(n16766) );
  XOR U17080 ( .A(n16765), .B(n16766), .Z(n16776) );
  NANDN U17081 ( .A(n16660), .B(n16659), .Z(n16664) );
  OR U17082 ( .A(n16662), .B(n16661), .Z(n16663) );
  AND U17083 ( .A(n16664), .B(n16663), .Z(n16775) );
  XNOR U17084 ( .A(n16776), .B(n16775), .Z(n16777) );
  NANDN U17085 ( .A(n16666), .B(n16665), .Z(n16670) );
  NANDN U17086 ( .A(n16668), .B(n16667), .Z(n16669) );
  NAND U17087 ( .A(n16670), .B(n16669), .Z(n16778) );
  XNOR U17088 ( .A(n16777), .B(n16778), .Z(n16724) );
  NANDN U17089 ( .A(n16672), .B(n16671), .Z(n16676) );
  NANDN U17090 ( .A(n16674), .B(n16673), .Z(n16675) );
  AND U17091 ( .A(n16676), .B(n16675), .Z(n16750) );
  NAND U17092 ( .A(b[0]), .B(a[224]), .Z(n16677) );
  XNOR U17093 ( .A(b[1]), .B(n16677), .Z(n16679) );
  NANDN U17094 ( .A(b[0]), .B(a[223]), .Z(n16678) );
  NAND U17095 ( .A(n16679), .B(n16678), .Z(n16730) );
  NAND U17096 ( .A(n19808), .B(n16680), .Z(n16682) );
  XOR U17097 ( .A(b[13]), .B(a[212]), .Z(n16733) );
  NAND U17098 ( .A(n19768), .B(n16733), .Z(n16681) );
  AND U17099 ( .A(n16682), .B(n16681), .Z(n16728) );
  AND U17100 ( .A(b[15]), .B(a[208]), .Z(n16727) );
  XNOR U17101 ( .A(n16728), .B(n16727), .Z(n16729) );
  XNOR U17102 ( .A(n16730), .B(n16729), .Z(n16748) );
  NAND U17103 ( .A(n33), .B(n16683), .Z(n16685) );
  XOR U17104 ( .A(b[5]), .B(a[220]), .Z(n16739) );
  NAND U17105 ( .A(n19342), .B(n16739), .Z(n16684) );
  AND U17106 ( .A(n16685), .B(n16684), .Z(n16772) );
  NAND U17107 ( .A(n34), .B(n16686), .Z(n16688) );
  XOR U17108 ( .A(b[7]), .B(a[218]), .Z(n16742) );
  NAND U17109 ( .A(n19486), .B(n16742), .Z(n16687) );
  AND U17110 ( .A(n16688), .B(n16687), .Z(n16770) );
  NAND U17111 ( .A(n31), .B(n16689), .Z(n16691) );
  XOR U17112 ( .A(b[3]), .B(a[222]), .Z(n16745) );
  NAND U17113 ( .A(n32), .B(n16745), .Z(n16690) );
  NAND U17114 ( .A(n16691), .B(n16690), .Z(n16769) );
  XNOR U17115 ( .A(n16770), .B(n16769), .Z(n16771) );
  XOR U17116 ( .A(n16772), .B(n16771), .Z(n16749) );
  XOR U17117 ( .A(n16748), .B(n16749), .Z(n16751) );
  XOR U17118 ( .A(n16750), .B(n16751), .Z(n16722) );
  NANDN U17119 ( .A(n16693), .B(n16692), .Z(n16697) );
  OR U17120 ( .A(n16695), .B(n16694), .Z(n16696) );
  AND U17121 ( .A(n16697), .B(n16696), .Z(n16721) );
  XNOR U17122 ( .A(n16722), .B(n16721), .Z(n16723) );
  XOR U17123 ( .A(n16724), .B(n16723), .Z(n16782) );
  NANDN U17124 ( .A(n16699), .B(n16698), .Z(n16703) );
  NANDN U17125 ( .A(n16701), .B(n16700), .Z(n16702) );
  AND U17126 ( .A(n16703), .B(n16702), .Z(n16781) );
  XNOR U17127 ( .A(n16782), .B(n16781), .Z(n16783) );
  XOR U17128 ( .A(n16784), .B(n16783), .Z(n16716) );
  NANDN U17129 ( .A(n16705), .B(n16704), .Z(n16709) );
  NAND U17130 ( .A(n16707), .B(n16706), .Z(n16708) );
  AND U17131 ( .A(n16709), .B(n16708), .Z(n16715) );
  XNOR U17132 ( .A(n16716), .B(n16715), .Z(n16717) );
  XNOR U17133 ( .A(n16718), .B(n16717), .Z(n16787) );
  XNOR U17134 ( .A(sreg[464]), .B(n16787), .Z(n16789) );
  NANDN U17135 ( .A(sreg[463]), .B(n16710), .Z(n16714) );
  NAND U17136 ( .A(n16712), .B(n16711), .Z(n16713) );
  NAND U17137 ( .A(n16714), .B(n16713), .Z(n16788) );
  XNOR U17138 ( .A(n16789), .B(n16788), .Z(c[464]) );
  NANDN U17139 ( .A(n16716), .B(n16715), .Z(n16720) );
  NANDN U17140 ( .A(n16718), .B(n16717), .Z(n16719) );
  AND U17141 ( .A(n16720), .B(n16719), .Z(n16795) );
  NANDN U17142 ( .A(n16722), .B(n16721), .Z(n16726) );
  NAND U17143 ( .A(n16724), .B(n16723), .Z(n16725) );
  AND U17144 ( .A(n16726), .B(n16725), .Z(n16861) );
  NANDN U17145 ( .A(n16728), .B(n16727), .Z(n16732) );
  NANDN U17146 ( .A(n16730), .B(n16729), .Z(n16731) );
  AND U17147 ( .A(n16732), .B(n16731), .Z(n16848) );
  NAND U17148 ( .A(n19808), .B(n16733), .Z(n16735) );
  XOR U17149 ( .A(b[13]), .B(a[213]), .Z(n16831) );
  NAND U17150 ( .A(n19768), .B(n16831), .Z(n16734) );
  AND U17151 ( .A(n16735), .B(n16734), .Z(n16826) );
  AND U17152 ( .A(b[15]), .B(a[209]), .Z(n16825) );
  XNOR U17153 ( .A(n16826), .B(n16825), .Z(n16827) );
  NAND U17154 ( .A(b[0]), .B(a[225]), .Z(n16736) );
  XNOR U17155 ( .A(b[1]), .B(n16736), .Z(n16738) );
  NANDN U17156 ( .A(b[0]), .B(a[224]), .Z(n16737) );
  NAND U17157 ( .A(n16738), .B(n16737), .Z(n16828) );
  XNOR U17158 ( .A(n16827), .B(n16828), .Z(n16846) );
  NAND U17159 ( .A(n33), .B(n16739), .Z(n16741) );
  XOR U17160 ( .A(b[5]), .B(a[221]), .Z(n16837) );
  NAND U17161 ( .A(n19342), .B(n16837), .Z(n16740) );
  AND U17162 ( .A(n16741), .B(n16740), .Z(n16822) );
  NAND U17163 ( .A(n34), .B(n16742), .Z(n16744) );
  XOR U17164 ( .A(b[7]), .B(a[219]), .Z(n16840) );
  NAND U17165 ( .A(n19486), .B(n16840), .Z(n16743) );
  AND U17166 ( .A(n16744), .B(n16743), .Z(n16820) );
  NAND U17167 ( .A(n31), .B(n16745), .Z(n16747) );
  XOR U17168 ( .A(b[3]), .B(a[223]), .Z(n16843) );
  NAND U17169 ( .A(n32), .B(n16843), .Z(n16746) );
  NAND U17170 ( .A(n16747), .B(n16746), .Z(n16819) );
  XNOR U17171 ( .A(n16820), .B(n16819), .Z(n16821) );
  XOR U17172 ( .A(n16822), .B(n16821), .Z(n16847) );
  XOR U17173 ( .A(n16846), .B(n16847), .Z(n16849) );
  XOR U17174 ( .A(n16848), .B(n16849), .Z(n16799) );
  NANDN U17175 ( .A(n16749), .B(n16748), .Z(n16753) );
  OR U17176 ( .A(n16751), .B(n16750), .Z(n16752) );
  AND U17177 ( .A(n16753), .B(n16752), .Z(n16798) );
  XNOR U17178 ( .A(n16799), .B(n16798), .Z(n16801) );
  NAND U17179 ( .A(n16754), .B(n19724), .Z(n16756) );
  XOR U17180 ( .A(b[11]), .B(a[215]), .Z(n16804) );
  NAND U17181 ( .A(n19692), .B(n16804), .Z(n16755) );
  AND U17182 ( .A(n16756), .B(n16755), .Z(n16815) );
  NAND U17183 ( .A(n19838), .B(n16757), .Z(n16759) );
  XOR U17184 ( .A(b[15]), .B(a[211]), .Z(n16807) );
  NAND U17185 ( .A(n19805), .B(n16807), .Z(n16758) );
  AND U17186 ( .A(n16759), .B(n16758), .Z(n16814) );
  NAND U17187 ( .A(n35), .B(n16760), .Z(n16762) );
  XOR U17188 ( .A(b[9]), .B(a[217]), .Z(n16810) );
  NAND U17189 ( .A(n19598), .B(n16810), .Z(n16761) );
  NAND U17190 ( .A(n16762), .B(n16761), .Z(n16813) );
  XOR U17191 ( .A(n16814), .B(n16813), .Z(n16816) );
  XOR U17192 ( .A(n16815), .B(n16816), .Z(n16853) );
  NANDN U17193 ( .A(n16764), .B(n16763), .Z(n16768) );
  OR U17194 ( .A(n16766), .B(n16765), .Z(n16767) );
  AND U17195 ( .A(n16768), .B(n16767), .Z(n16852) );
  XNOR U17196 ( .A(n16853), .B(n16852), .Z(n16854) );
  NANDN U17197 ( .A(n16770), .B(n16769), .Z(n16774) );
  NANDN U17198 ( .A(n16772), .B(n16771), .Z(n16773) );
  NAND U17199 ( .A(n16774), .B(n16773), .Z(n16855) );
  XNOR U17200 ( .A(n16854), .B(n16855), .Z(n16800) );
  XOR U17201 ( .A(n16801), .B(n16800), .Z(n16859) );
  NANDN U17202 ( .A(n16776), .B(n16775), .Z(n16780) );
  NANDN U17203 ( .A(n16778), .B(n16777), .Z(n16779) );
  AND U17204 ( .A(n16780), .B(n16779), .Z(n16858) );
  XNOR U17205 ( .A(n16859), .B(n16858), .Z(n16860) );
  XOR U17206 ( .A(n16861), .B(n16860), .Z(n16793) );
  NANDN U17207 ( .A(n16782), .B(n16781), .Z(n16786) );
  NAND U17208 ( .A(n16784), .B(n16783), .Z(n16785) );
  AND U17209 ( .A(n16786), .B(n16785), .Z(n16792) );
  XNOR U17210 ( .A(n16793), .B(n16792), .Z(n16794) );
  XNOR U17211 ( .A(n16795), .B(n16794), .Z(n16864) );
  XNOR U17212 ( .A(sreg[465]), .B(n16864), .Z(n16866) );
  NANDN U17213 ( .A(sreg[464]), .B(n16787), .Z(n16791) );
  NAND U17214 ( .A(n16789), .B(n16788), .Z(n16790) );
  NAND U17215 ( .A(n16791), .B(n16790), .Z(n16865) );
  XNOR U17216 ( .A(n16866), .B(n16865), .Z(c[465]) );
  NANDN U17217 ( .A(n16793), .B(n16792), .Z(n16797) );
  NANDN U17218 ( .A(n16795), .B(n16794), .Z(n16796) );
  AND U17219 ( .A(n16797), .B(n16796), .Z(n16872) );
  NANDN U17220 ( .A(n16799), .B(n16798), .Z(n16803) );
  NAND U17221 ( .A(n16801), .B(n16800), .Z(n16802) );
  AND U17222 ( .A(n16803), .B(n16802), .Z(n16938) );
  NAND U17223 ( .A(n16804), .B(n19724), .Z(n16806) );
  XOR U17224 ( .A(b[11]), .B(a[216]), .Z(n16908) );
  NAND U17225 ( .A(n19692), .B(n16908), .Z(n16805) );
  AND U17226 ( .A(n16806), .B(n16805), .Z(n16919) );
  NAND U17227 ( .A(n19838), .B(n16807), .Z(n16809) );
  XOR U17228 ( .A(b[15]), .B(a[212]), .Z(n16911) );
  NAND U17229 ( .A(n19805), .B(n16911), .Z(n16808) );
  AND U17230 ( .A(n16809), .B(n16808), .Z(n16918) );
  NAND U17231 ( .A(n35), .B(n16810), .Z(n16812) );
  XOR U17232 ( .A(b[9]), .B(a[218]), .Z(n16914) );
  NAND U17233 ( .A(n19598), .B(n16914), .Z(n16811) );
  NAND U17234 ( .A(n16812), .B(n16811), .Z(n16917) );
  XOR U17235 ( .A(n16918), .B(n16917), .Z(n16920) );
  XOR U17236 ( .A(n16919), .B(n16920), .Z(n16930) );
  NANDN U17237 ( .A(n16814), .B(n16813), .Z(n16818) );
  OR U17238 ( .A(n16816), .B(n16815), .Z(n16817) );
  AND U17239 ( .A(n16818), .B(n16817), .Z(n16929) );
  XNOR U17240 ( .A(n16930), .B(n16929), .Z(n16931) );
  NANDN U17241 ( .A(n16820), .B(n16819), .Z(n16824) );
  NANDN U17242 ( .A(n16822), .B(n16821), .Z(n16823) );
  NAND U17243 ( .A(n16824), .B(n16823), .Z(n16932) );
  XNOR U17244 ( .A(n16931), .B(n16932), .Z(n16878) );
  NANDN U17245 ( .A(n16826), .B(n16825), .Z(n16830) );
  NANDN U17246 ( .A(n16828), .B(n16827), .Z(n16829) );
  AND U17247 ( .A(n16830), .B(n16829), .Z(n16904) );
  NAND U17248 ( .A(n19808), .B(n16831), .Z(n16833) );
  XOR U17249 ( .A(b[13]), .B(a[214]), .Z(n16890) );
  NAND U17250 ( .A(n19768), .B(n16890), .Z(n16832) );
  AND U17251 ( .A(n16833), .B(n16832), .Z(n16882) );
  AND U17252 ( .A(b[15]), .B(a[210]), .Z(n16881) );
  XNOR U17253 ( .A(n16882), .B(n16881), .Z(n16883) );
  NAND U17254 ( .A(b[0]), .B(a[226]), .Z(n16834) );
  XNOR U17255 ( .A(b[1]), .B(n16834), .Z(n16836) );
  NANDN U17256 ( .A(b[0]), .B(a[225]), .Z(n16835) );
  NAND U17257 ( .A(n16836), .B(n16835), .Z(n16884) );
  XNOR U17258 ( .A(n16883), .B(n16884), .Z(n16902) );
  NAND U17259 ( .A(n33), .B(n16837), .Z(n16839) );
  XOR U17260 ( .A(b[5]), .B(a[222]), .Z(n16893) );
  NAND U17261 ( .A(n19342), .B(n16893), .Z(n16838) );
  AND U17262 ( .A(n16839), .B(n16838), .Z(n16926) );
  NAND U17263 ( .A(n34), .B(n16840), .Z(n16842) );
  XOR U17264 ( .A(b[7]), .B(a[220]), .Z(n16896) );
  NAND U17265 ( .A(n19486), .B(n16896), .Z(n16841) );
  AND U17266 ( .A(n16842), .B(n16841), .Z(n16924) );
  NAND U17267 ( .A(n31), .B(n16843), .Z(n16845) );
  XOR U17268 ( .A(b[3]), .B(a[224]), .Z(n16899) );
  NAND U17269 ( .A(n32), .B(n16899), .Z(n16844) );
  NAND U17270 ( .A(n16845), .B(n16844), .Z(n16923) );
  XNOR U17271 ( .A(n16924), .B(n16923), .Z(n16925) );
  XOR U17272 ( .A(n16926), .B(n16925), .Z(n16903) );
  XOR U17273 ( .A(n16902), .B(n16903), .Z(n16905) );
  XOR U17274 ( .A(n16904), .B(n16905), .Z(n16876) );
  NANDN U17275 ( .A(n16847), .B(n16846), .Z(n16851) );
  OR U17276 ( .A(n16849), .B(n16848), .Z(n16850) );
  AND U17277 ( .A(n16851), .B(n16850), .Z(n16875) );
  XNOR U17278 ( .A(n16876), .B(n16875), .Z(n16877) );
  XOR U17279 ( .A(n16878), .B(n16877), .Z(n16936) );
  NANDN U17280 ( .A(n16853), .B(n16852), .Z(n16857) );
  NANDN U17281 ( .A(n16855), .B(n16854), .Z(n16856) );
  AND U17282 ( .A(n16857), .B(n16856), .Z(n16935) );
  XNOR U17283 ( .A(n16936), .B(n16935), .Z(n16937) );
  XOR U17284 ( .A(n16938), .B(n16937), .Z(n16870) );
  NANDN U17285 ( .A(n16859), .B(n16858), .Z(n16863) );
  NAND U17286 ( .A(n16861), .B(n16860), .Z(n16862) );
  AND U17287 ( .A(n16863), .B(n16862), .Z(n16869) );
  XNOR U17288 ( .A(n16870), .B(n16869), .Z(n16871) );
  XNOR U17289 ( .A(n16872), .B(n16871), .Z(n16941) );
  XNOR U17290 ( .A(sreg[466]), .B(n16941), .Z(n16943) );
  NANDN U17291 ( .A(sreg[465]), .B(n16864), .Z(n16868) );
  NAND U17292 ( .A(n16866), .B(n16865), .Z(n16867) );
  NAND U17293 ( .A(n16868), .B(n16867), .Z(n16942) );
  XNOR U17294 ( .A(n16943), .B(n16942), .Z(c[466]) );
  NANDN U17295 ( .A(n16870), .B(n16869), .Z(n16874) );
  NANDN U17296 ( .A(n16872), .B(n16871), .Z(n16873) );
  AND U17297 ( .A(n16874), .B(n16873), .Z(n16949) );
  NANDN U17298 ( .A(n16876), .B(n16875), .Z(n16880) );
  NAND U17299 ( .A(n16878), .B(n16877), .Z(n16879) );
  AND U17300 ( .A(n16880), .B(n16879), .Z(n17015) );
  NANDN U17301 ( .A(n16882), .B(n16881), .Z(n16886) );
  NANDN U17302 ( .A(n16884), .B(n16883), .Z(n16885) );
  AND U17303 ( .A(n16886), .B(n16885), .Z(n16981) );
  NAND U17304 ( .A(b[0]), .B(a[227]), .Z(n16887) );
  XNOR U17305 ( .A(b[1]), .B(n16887), .Z(n16889) );
  NANDN U17306 ( .A(b[0]), .B(a[226]), .Z(n16888) );
  NAND U17307 ( .A(n16889), .B(n16888), .Z(n16961) );
  NAND U17308 ( .A(n19808), .B(n16890), .Z(n16892) );
  XOR U17309 ( .A(b[13]), .B(a[215]), .Z(n16967) );
  NAND U17310 ( .A(n19768), .B(n16967), .Z(n16891) );
  AND U17311 ( .A(n16892), .B(n16891), .Z(n16959) );
  AND U17312 ( .A(b[15]), .B(a[211]), .Z(n16958) );
  XNOR U17313 ( .A(n16959), .B(n16958), .Z(n16960) );
  XNOR U17314 ( .A(n16961), .B(n16960), .Z(n16979) );
  NAND U17315 ( .A(n33), .B(n16893), .Z(n16895) );
  XOR U17316 ( .A(b[5]), .B(a[223]), .Z(n16970) );
  NAND U17317 ( .A(n19342), .B(n16970), .Z(n16894) );
  AND U17318 ( .A(n16895), .B(n16894), .Z(n17003) );
  NAND U17319 ( .A(n34), .B(n16896), .Z(n16898) );
  XOR U17320 ( .A(b[7]), .B(a[221]), .Z(n16973) );
  NAND U17321 ( .A(n19486), .B(n16973), .Z(n16897) );
  AND U17322 ( .A(n16898), .B(n16897), .Z(n17001) );
  NAND U17323 ( .A(n31), .B(n16899), .Z(n16901) );
  XOR U17324 ( .A(b[3]), .B(a[225]), .Z(n16976) );
  NAND U17325 ( .A(n32), .B(n16976), .Z(n16900) );
  NAND U17326 ( .A(n16901), .B(n16900), .Z(n17000) );
  XNOR U17327 ( .A(n17001), .B(n17000), .Z(n17002) );
  XOR U17328 ( .A(n17003), .B(n17002), .Z(n16980) );
  XOR U17329 ( .A(n16979), .B(n16980), .Z(n16982) );
  XOR U17330 ( .A(n16981), .B(n16982), .Z(n16953) );
  NANDN U17331 ( .A(n16903), .B(n16902), .Z(n16907) );
  OR U17332 ( .A(n16905), .B(n16904), .Z(n16906) );
  AND U17333 ( .A(n16907), .B(n16906), .Z(n16952) );
  XNOR U17334 ( .A(n16953), .B(n16952), .Z(n16955) );
  NAND U17335 ( .A(n16908), .B(n19724), .Z(n16910) );
  XOR U17336 ( .A(b[11]), .B(a[217]), .Z(n16985) );
  NAND U17337 ( .A(n19692), .B(n16985), .Z(n16909) );
  AND U17338 ( .A(n16910), .B(n16909), .Z(n16996) );
  NAND U17339 ( .A(n19838), .B(n16911), .Z(n16913) );
  XOR U17340 ( .A(b[15]), .B(a[213]), .Z(n16988) );
  NAND U17341 ( .A(n19805), .B(n16988), .Z(n16912) );
  AND U17342 ( .A(n16913), .B(n16912), .Z(n16995) );
  NAND U17343 ( .A(n35), .B(n16914), .Z(n16916) );
  XOR U17344 ( .A(b[9]), .B(a[219]), .Z(n16991) );
  NAND U17345 ( .A(n19598), .B(n16991), .Z(n16915) );
  NAND U17346 ( .A(n16916), .B(n16915), .Z(n16994) );
  XOR U17347 ( .A(n16995), .B(n16994), .Z(n16997) );
  XOR U17348 ( .A(n16996), .B(n16997), .Z(n17007) );
  NANDN U17349 ( .A(n16918), .B(n16917), .Z(n16922) );
  OR U17350 ( .A(n16920), .B(n16919), .Z(n16921) );
  AND U17351 ( .A(n16922), .B(n16921), .Z(n17006) );
  XNOR U17352 ( .A(n17007), .B(n17006), .Z(n17008) );
  NANDN U17353 ( .A(n16924), .B(n16923), .Z(n16928) );
  NANDN U17354 ( .A(n16926), .B(n16925), .Z(n16927) );
  NAND U17355 ( .A(n16928), .B(n16927), .Z(n17009) );
  XNOR U17356 ( .A(n17008), .B(n17009), .Z(n16954) );
  XOR U17357 ( .A(n16955), .B(n16954), .Z(n17013) );
  NANDN U17358 ( .A(n16930), .B(n16929), .Z(n16934) );
  NANDN U17359 ( .A(n16932), .B(n16931), .Z(n16933) );
  AND U17360 ( .A(n16934), .B(n16933), .Z(n17012) );
  XNOR U17361 ( .A(n17013), .B(n17012), .Z(n17014) );
  XOR U17362 ( .A(n17015), .B(n17014), .Z(n16947) );
  NANDN U17363 ( .A(n16936), .B(n16935), .Z(n16940) );
  NAND U17364 ( .A(n16938), .B(n16937), .Z(n16939) );
  AND U17365 ( .A(n16940), .B(n16939), .Z(n16946) );
  XNOR U17366 ( .A(n16947), .B(n16946), .Z(n16948) );
  XNOR U17367 ( .A(n16949), .B(n16948), .Z(n17018) );
  XNOR U17368 ( .A(sreg[467]), .B(n17018), .Z(n17020) );
  NANDN U17369 ( .A(sreg[466]), .B(n16941), .Z(n16945) );
  NAND U17370 ( .A(n16943), .B(n16942), .Z(n16944) );
  NAND U17371 ( .A(n16945), .B(n16944), .Z(n17019) );
  XNOR U17372 ( .A(n17020), .B(n17019), .Z(c[467]) );
  NANDN U17373 ( .A(n16947), .B(n16946), .Z(n16951) );
  NANDN U17374 ( .A(n16949), .B(n16948), .Z(n16950) );
  AND U17375 ( .A(n16951), .B(n16950), .Z(n17026) );
  NANDN U17376 ( .A(n16953), .B(n16952), .Z(n16957) );
  NAND U17377 ( .A(n16955), .B(n16954), .Z(n16956) );
  AND U17378 ( .A(n16957), .B(n16956), .Z(n17092) );
  NANDN U17379 ( .A(n16959), .B(n16958), .Z(n16963) );
  NANDN U17380 ( .A(n16961), .B(n16960), .Z(n16962) );
  AND U17381 ( .A(n16963), .B(n16962), .Z(n17058) );
  NAND U17382 ( .A(b[0]), .B(a[228]), .Z(n16964) );
  XNOR U17383 ( .A(b[1]), .B(n16964), .Z(n16966) );
  NANDN U17384 ( .A(b[0]), .B(a[227]), .Z(n16965) );
  NAND U17385 ( .A(n16966), .B(n16965), .Z(n17038) );
  NAND U17386 ( .A(n19808), .B(n16967), .Z(n16969) );
  XOR U17387 ( .A(b[13]), .B(a[216]), .Z(n17041) );
  NAND U17388 ( .A(n19768), .B(n17041), .Z(n16968) );
  AND U17389 ( .A(n16969), .B(n16968), .Z(n17036) );
  AND U17390 ( .A(b[15]), .B(a[212]), .Z(n17035) );
  XNOR U17391 ( .A(n17036), .B(n17035), .Z(n17037) );
  XNOR U17392 ( .A(n17038), .B(n17037), .Z(n17056) );
  NAND U17393 ( .A(n33), .B(n16970), .Z(n16972) );
  XOR U17394 ( .A(b[5]), .B(a[224]), .Z(n17047) );
  NAND U17395 ( .A(n19342), .B(n17047), .Z(n16971) );
  AND U17396 ( .A(n16972), .B(n16971), .Z(n17080) );
  NAND U17397 ( .A(n34), .B(n16973), .Z(n16975) );
  XOR U17398 ( .A(b[7]), .B(a[222]), .Z(n17050) );
  NAND U17399 ( .A(n19486), .B(n17050), .Z(n16974) );
  AND U17400 ( .A(n16975), .B(n16974), .Z(n17078) );
  NAND U17401 ( .A(n31), .B(n16976), .Z(n16978) );
  XOR U17402 ( .A(b[3]), .B(a[226]), .Z(n17053) );
  NAND U17403 ( .A(n32), .B(n17053), .Z(n16977) );
  NAND U17404 ( .A(n16978), .B(n16977), .Z(n17077) );
  XNOR U17405 ( .A(n17078), .B(n17077), .Z(n17079) );
  XOR U17406 ( .A(n17080), .B(n17079), .Z(n17057) );
  XOR U17407 ( .A(n17056), .B(n17057), .Z(n17059) );
  XOR U17408 ( .A(n17058), .B(n17059), .Z(n17030) );
  NANDN U17409 ( .A(n16980), .B(n16979), .Z(n16984) );
  OR U17410 ( .A(n16982), .B(n16981), .Z(n16983) );
  AND U17411 ( .A(n16984), .B(n16983), .Z(n17029) );
  XNOR U17412 ( .A(n17030), .B(n17029), .Z(n17032) );
  NAND U17413 ( .A(n16985), .B(n19724), .Z(n16987) );
  XOR U17414 ( .A(b[11]), .B(a[218]), .Z(n17062) );
  NAND U17415 ( .A(n19692), .B(n17062), .Z(n16986) );
  AND U17416 ( .A(n16987), .B(n16986), .Z(n17073) );
  NAND U17417 ( .A(n19838), .B(n16988), .Z(n16990) );
  XOR U17418 ( .A(b[15]), .B(a[214]), .Z(n17065) );
  NAND U17419 ( .A(n19805), .B(n17065), .Z(n16989) );
  AND U17420 ( .A(n16990), .B(n16989), .Z(n17072) );
  NAND U17421 ( .A(n35), .B(n16991), .Z(n16993) );
  XOR U17422 ( .A(b[9]), .B(a[220]), .Z(n17068) );
  NAND U17423 ( .A(n19598), .B(n17068), .Z(n16992) );
  NAND U17424 ( .A(n16993), .B(n16992), .Z(n17071) );
  XOR U17425 ( .A(n17072), .B(n17071), .Z(n17074) );
  XOR U17426 ( .A(n17073), .B(n17074), .Z(n17084) );
  NANDN U17427 ( .A(n16995), .B(n16994), .Z(n16999) );
  OR U17428 ( .A(n16997), .B(n16996), .Z(n16998) );
  AND U17429 ( .A(n16999), .B(n16998), .Z(n17083) );
  XNOR U17430 ( .A(n17084), .B(n17083), .Z(n17085) );
  NANDN U17431 ( .A(n17001), .B(n17000), .Z(n17005) );
  NANDN U17432 ( .A(n17003), .B(n17002), .Z(n17004) );
  NAND U17433 ( .A(n17005), .B(n17004), .Z(n17086) );
  XNOR U17434 ( .A(n17085), .B(n17086), .Z(n17031) );
  XOR U17435 ( .A(n17032), .B(n17031), .Z(n17090) );
  NANDN U17436 ( .A(n17007), .B(n17006), .Z(n17011) );
  NANDN U17437 ( .A(n17009), .B(n17008), .Z(n17010) );
  AND U17438 ( .A(n17011), .B(n17010), .Z(n17089) );
  XNOR U17439 ( .A(n17090), .B(n17089), .Z(n17091) );
  XOR U17440 ( .A(n17092), .B(n17091), .Z(n17024) );
  NANDN U17441 ( .A(n17013), .B(n17012), .Z(n17017) );
  NAND U17442 ( .A(n17015), .B(n17014), .Z(n17016) );
  AND U17443 ( .A(n17017), .B(n17016), .Z(n17023) );
  XNOR U17444 ( .A(n17024), .B(n17023), .Z(n17025) );
  XNOR U17445 ( .A(n17026), .B(n17025), .Z(n17095) );
  XNOR U17446 ( .A(sreg[468]), .B(n17095), .Z(n17097) );
  NANDN U17447 ( .A(sreg[467]), .B(n17018), .Z(n17022) );
  NAND U17448 ( .A(n17020), .B(n17019), .Z(n17021) );
  NAND U17449 ( .A(n17022), .B(n17021), .Z(n17096) );
  XNOR U17450 ( .A(n17097), .B(n17096), .Z(c[468]) );
  NANDN U17451 ( .A(n17024), .B(n17023), .Z(n17028) );
  NANDN U17452 ( .A(n17026), .B(n17025), .Z(n17027) );
  AND U17453 ( .A(n17028), .B(n17027), .Z(n17103) );
  NANDN U17454 ( .A(n17030), .B(n17029), .Z(n17034) );
  NAND U17455 ( .A(n17032), .B(n17031), .Z(n17033) );
  AND U17456 ( .A(n17034), .B(n17033), .Z(n17169) );
  NANDN U17457 ( .A(n17036), .B(n17035), .Z(n17040) );
  NANDN U17458 ( .A(n17038), .B(n17037), .Z(n17039) );
  AND U17459 ( .A(n17040), .B(n17039), .Z(n17135) );
  NAND U17460 ( .A(n19808), .B(n17041), .Z(n17043) );
  XOR U17461 ( .A(b[13]), .B(a[217]), .Z(n17121) );
  NAND U17462 ( .A(n19768), .B(n17121), .Z(n17042) );
  AND U17463 ( .A(n17043), .B(n17042), .Z(n17113) );
  AND U17464 ( .A(b[15]), .B(a[213]), .Z(n17112) );
  XNOR U17465 ( .A(n17113), .B(n17112), .Z(n17114) );
  NAND U17466 ( .A(b[0]), .B(a[229]), .Z(n17044) );
  XNOR U17467 ( .A(b[1]), .B(n17044), .Z(n17046) );
  NANDN U17468 ( .A(b[0]), .B(a[228]), .Z(n17045) );
  NAND U17469 ( .A(n17046), .B(n17045), .Z(n17115) );
  XNOR U17470 ( .A(n17114), .B(n17115), .Z(n17133) );
  NAND U17471 ( .A(n33), .B(n17047), .Z(n17049) );
  XOR U17472 ( .A(b[5]), .B(a[225]), .Z(n17124) );
  NAND U17473 ( .A(n19342), .B(n17124), .Z(n17048) );
  AND U17474 ( .A(n17049), .B(n17048), .Z(n17157) );
  NAND U17475 ( .A(n34), .B(n17050), .Z(n17052) );
  XOR U17476 ( .A(b[7]), .B(a[223]), .Z(n17127) );
  NAND U17477 ( .A(n19486), .B(n17127), .Z(n17051) );
  AND U17478 ( .A(n17052), .B(n17051), .Z(n17155) );
  NAND U17479 ( .A(n31), .B(n17053), .Z(n17055) );
  XOR U17480 ( .A(b[3]), .B(a[227]), .Z(n17130) );
  NAND U17481 ( .A(n32), .B(n17130), .Z(n17054) );
  NAND U17482 ( .A(n17055), .B(n17054), .Z(n17154) );
  XNOR U17483 ( .A(n17155), .B(n17154), .Z(n17156) );
  XOR U17484 ( .A(n17157), .B(n17156), .Z(n17134) );
  XOR U17485 ( .A(n17133), .B(n17134), .Z(n17136) );
  XOR U17486 ( .A(n17135), .B(n17136), .Z(n17107) );
  NANDN U17487 ( .A(n17057), .B(n17056), .Z(n17061) );
  OR U17488 ( .A(n17059), .B(n17058), .Z(n17060) );
  AND U17489 ( .A(n17061), .B(n17060), .Z(n17106) );
  XNOR U17490 ( .A(n17107), .B(n17106), .Z(n17109) );
  NAND U17491 ( .A(n17062), .B(n19724), .Z(n17064) );
  XOR U17492 ( .A(b[11]), .B(a[219]), .Z(n17139) );
  NAND U17493 ( .A(n19692), .B(n17139), .Z(n17063) );
  AND U17494 ( .A(n17064), .B(n17063), .Z(n17150) );
  NAND U17495 ( .A(n19838), .B(n17065), .Z(n17067) );
  XOR U17496 ( .A(b[15]), .B(a[215]), .Z(n17142) );
  NAND U17497 ( .A(n19805), .B(n17142), .Z(n17066) );
  AND U17498 ( .A(n17067), .B(n17066), .Z(n17149) );
  NAND U17499 ( .A(n35), .B(n17068), .Z(n17070) );
  XOR U17500 ( .A(b[9]), .B(a[221]), .Z(n17145) );
  NAND U17501 ( .A(n19598), .B(n17145), .Z(n17069) );
  NAND U17502 ( .A(n17070), .B(n17069), .Z(n17148) );
  XOR U17503 ( .A(n17149), .B(n17148), .Z(n17151) );
  XOR U17504 ( .A(n17150), .B(n17151), .Z(n17161) );
  NANDN U17505 ( .A(n17072), .B(n17071), .Z(n17076) );
  OR U17506 ( .A(n17074), .B(n17073), .Z(n17075) );
  AND U17507 ( .A(n17076), .B(n17075), .Z(n17160) );
  XNOR U17508 ( .A(n17161), .B(n17160), .Z(n17162) );
  NANDN U17509 ( .A(n17078), .B(n17077), .Z(n17082) );
  NANDN U17510 ( .A(n17080), .B(n17079), .Z(n17081) );
  NAND U17511 ( .A(n17082), .B(n17081), .Z(n17163) );
  XNOR U17512 ( .A(n17162), .B(n17163), .Z(n17108) );
  XOR U17513 ( .A(n17109), .B(n17108), .Z(n17167) );
  NANDN U17514 ( .A(n17084), .B(n17083), .Z(n17088) );
  NANDN U17515 ( .A(n17086), .B(n17085), .Z(n17087) );
  AND U17516 ( .A(n17088), .B(n17087), .Z(n17166) );
  XNOR U17517 ( .A(n17167), .B(n17166), .Z(n17168) );
  XOR U17518 ( .A(n17169), .B(n17168), .Z(n17101) );
  NANDN U17519 ( .A(n17090), .B(n17089), .Z(n17094) );
  NAND U17520 ( .A(n17092), .B(n17091), .Z(n17093) );
  AND U17521 ( .A(n17094), .B(n17093), .Z(n17100) );
  XNOR U17522 ( .A(n17101), .B(n17100), .Z(n17102) );
  XNOR U17523 ( .A(n17103), .B(n17102), .Z(n17172) );
  XNOR U17524 ( .A(sreg[469]), .B(n17172), .Z(n17174) );
  NANDN U17525 ( .A(sreg[468]), .B(n17095), .Z(n17099) );
  NAND U17526 ( .A(n17097), .B(n17096), .Z(n17098) );
  NAND U17527 ( .A(n17099), .B(n17098), .Z(n17173) );
  XNOR U17528 ( .A(n17174), .B(n17173), .Z(c[469]) );
  NANDN U17529 ( .A(n17101), .B(n17100), .Z(n17105) );
  NANDN U17530 ( .A(n17103), .B(n17102), .Z(n17104) );
  AND U17531 ( .A(n17105), .B(n17104), .Z(n17180) );
  NANDN U17532 ( .A(n17107), .B(n17106), .Z(n17111) );
  NAND U17533 ( .A(n17109), .B(n17108), .Z(n17110) );
  AND U17534 ( .A(n17111), .B(n17110), .Z(n17246) );
  NANDN U17535 ( .A(n17113), .B(n17112), .Z(n17117) );
  NANDN U17536 ( .A(n17115), .B(n17114), .Z(n17116) );
  AND U17537 ( .A(n17117), .B(n17116), .Z(n17212) );
  NAND U17538 ( .A(b[0]), .B(a[230]), .Z(n17118) );
  XNOR U17539 ( .A(b[1]), .B(n17118), .Z(n17120) );
  NANDN U17540 ( .A(b[0]), .B(a[229]), .Z(n17119) );
  NAND U17541 ( .A(n17120), .B(n17119), .Z(n17192) );
  NAND U17542 ( .A(n19808), .B(n17121), .Z(n17123) );
  XOR U17543 ( .A(b[13]), .B(a[218]), .Z(n17198) );
  NAND U17544 ( .A(n19768), .B(n17198), .Z(n17122) );
  AND U17545 ( .A(n17123), .B(n17122), .Z(n17190) );
  AND U17546 ( .A(b[15]), .B(a[214]), .Z(n17189) );
  XNOR U17547 ( .A(n17190), .B(n17189), .Z(n17191) );
  XNOR U17548 ( .A(n17192), .B(n17191), .Z(n17210) );
  NAND U17549 ( .A(n33), .B(n17124), .Z(n17126) );
  XOR U17550 ( .A(b[5]), .B(a[226]), .Z(n17201) );
  NAND U17551 ( .A(n19342), .B(n17201), .Z(n17125) );
  AND U17552 ( .A(n17126), .B(n17125), .Z(n17234) );
  NAND U17553 ( .A(n34), .B(n17127), .Z(n17129) );
  XOR U17554 ( .A(b[7]), .B(a[224]), .Z(n17204) );
  NAND U17555 ( .A(n19486), .B(n17204), .Z(n17128) );
  AND U17556 ( .A(n17129), .B(n17128), .Z(n17232) );
  NAND U17557 ( .A(n31), .B(n17130), .Z(n17132) );
  XOR U17558 ( .A(b[3]), .B(a[228]), .Z(n17207) );
  NAND U17559 ( .A(n32), .B(n17207), .Z(n17131) );
  NAND U17560 ( .A(n17132), .B(n17131), .Z(n17231) );
  XNOR U17561 ( .A(n17232), .B(n17231), .Z(n17233) );
  XOR U17562 ( .A(n17234), .B(n17233), .Z(n17211) );
  XOR U17563 ( .A(n17210), .B(n17211), .Z(n17213) );
  XOR U17564 ( .A(n17212), .B(n17213), .Z(n17184) );
  NANDN U17565 ( .A(n17134), .B(n17133), .Z(n17138) );
  OR U17566 ( .A(n17136), .B(n17135), .Z(n17137) );
  AND U17567 ( .A(n17138), .B(n17137), .Z(n17183) );
  XNOR U17568 ( .A(n17184), .B(n17183), .Z(n17186) );
  NAND U17569 ( .A(n17139), .B(n19724), .Z(n17141) );
  XOR U17570 ( .A(b[11]), .B(a[220]), .Z(n17216) );
  NAND U17571 ( .A(n19692), .B(n17216), .Z(n17140) );
  AND U17572 ( .A(n17141), .B(n17140), .Z(n17227) );
  NAND U17573 ( .A(n19838), .B(n17142), .Z(n17144) );
  XOR U17574 ( .A(b[15]), .B(a[216]), .Z(n17219) );
  NAND U17575 ( .A(n19805), .B(n17219), .Z(n17143) );
  AND U17576 ( .A(n17144), .B(n17143), .Z(n17226) );
  NAND U17577 ( .A(n35), .B(n17145), .Z(n17147) );
  XOR U17578 ( .A(b[9]), .B(a[222]), .Z(n17222) );
  NAND U17579 ( .A(n19598), .B(n17222), .Z(n17146) );
  NAND U17580 ( .A(n17147), .B(n17146), .Z(n17225) );
  XOR U17581 ( .A(n17226), .B(n17225), .Z(n17228) );
  XOR U17582 ( .A(n17227), .B(n17228), .Z(n17238) );
  NANDN U17583 ( .A(n17149), .B(n17148), .Z(n17153) );
  OR U17584 ( .A(n17151), .B(n17150), .Z(n17152) );
  AND U17585 ( .A(n17153), .B(n17152), .Z(n17237) );
  XNOR U17586 ( .A(n17238), .B(n17237), .Z(n17239) );
  NANDN U17587 ( .A(n17155), .B(n17154), .Z(n17159) );
  NANDN U17588 ( .A(n17157), .B(n17156), .Z(n17158) );
  NAND U17589 ( .A(n17159), .B(n17158), .Z(n17240) );
  XNOR U17590 ( .A(n17239), .B(n17240), .Z(n17185) );
  XOR U17591 ( .A(n17186), .B(n17185), .Z(n17244) );
  NANDN U17592 ( .A(n17161), .B(n17160), .Z(n17165) );
  NANDN U17593 ( .A(n17163), .B(n17162), .Z(n17164) );
  AND U17594 ( .A(n17165), .B(n17164), .Z(n17243) );
  XNOR U17595 ( .A(n17244), .B(n17243), .Z(n17245) );
  XOR U17596 ( .A(n17246), .B(n17245), .Z(n17178) );
  NANDN U17597 ( .A(n17167), .B(n17166), .Z(n17171) );
  NAND U17598 ( .A(n17169), .B(n17168), .Z(n17170) );
  AND U17599 ( .A(n17171), .B(n17170), .Z(n17177) );
  XNOR U17600 ( .A(n17178), .B(n17177), .Z(n17179) );
  XNOR U17601 ( .A(n17180), .B(n17179), .Z(n17249) );
  XNOR U17602 ( .A(sreg[470]), .B(n17249), .Z(n17251) );
  NANDN U17603 ( .A(sreg[469]), .B(n17172), .Z(n17176) );
  NAND U17604 ( .A(n17174), .B(n17173), .Z(n17175) );
  NAND U17605 ( .A(n17176), .B(n17175), .Z(n17250) );
  XNOR U17606 ( .A(n17251), .B(n17250), .Z(c[470]) );
  NANDN U17607 ( .A(n17178), .B(n17177), .Z(n17182) );
  NANDN U17608 ( .A(n17180), .B(n17179), .Z(n17181) );
  AND U17609 ( .A(n17182), .B(n17181), .Z(n17257) );
  NANDN U17610 ( .A(n17184), .B(n17183), .Z(n17188) );
  NAND U17611 ( .A(n17186), .B(n17185), .Z(n17187) );
  AND U17612 ( .A(n17188), .B(n17187), .Z(n17323) );
  NANDN U17613 ( .A(n17190), .B(n17189), .Z(n17194) );
  NANDN U17614 ( .A(n17192), .B(n17191), .Z(n17193) );
  AND U17615 ( .A(n17194), .B(n17193), .Z(n17289) );
  NAND U17616 ( .A(b[0]), .B(a[231]), .Z(n17195) );
  XNOR U17617 ( .A(b[1]), .B(n17195), .Z(n17197) );
  NANDN U17618 ( .A(b[0]), .B(a[230]), .Z(n17196) );
  NAND U17619 ( .A(n17197), .B(n17196), .Z(n17269) );
  NAND U17620 ( .A(n19808), .B(n17198), .Z(n17200) );
  XOR U17621 ( .A(b[13]), .B(a[219]), .Z(n17272) );
  NAND U17622 ( .A(n19768), .B(n17272), .Z(n17199) );
  AND U17623 ( .A(n17200), .B(n17199), .Z(n17267) );
  AND U17624 ( .A(b[15]), .B(a[215]), .Z(n17266) );
  XNOR U17625 ( .A(n17267), .B(n17266), .Z(n17268) );
  XNOR U17626 ( .A(n17269), .B(n17268), .Z(n17287) );
  NAND U17627 ( .A(n33), .B(n17201), .Z(n17203) );
  XOR U17628 ( .A(b[5]), .B(a[227]), .Z(n17278) );
  NAND U17629 ( .A(n19342), .B(n17278), .Z(n17202) );
  AND U17630 ( .A(n17203), .B(n17202), .Z(n17311) );
  NAND U17631 ( .A(n34), .B(n17204), .Z(n17206) );
  XOR U17632 ( .A(b[7]), .B(a[225]), .Z(n17281) );
  NAND U17633 ( .A(n19486), .B(n17281), .Z(n17205) );
  AND U17634 ( .A(n17206), .B(n17205), .Z(n17309) );
  NAND U17635 ( .A(n31), .B(n17207), .Z(n17209) );
  XOR U17636 ( .A(b[3]), .B(a[229]), .Z(n17284) );
  NAND U17637 ( .A(n32), .B(n17284), .Z(n17208) );
  NAND U17638 ( .A(n17209), .B(n17208), .Z(n17308) );
  XNOR U17639 ( .A(n17309), .B(n17308), .Z(n17310) );
  XOR U17640 ( .A(n17311), .B(n17310), .Z(n17288) );
  XOR U17641 ( .A(n17287), .B(n17288), .Z(n17290) );
  XOR U17642 ( .A(n17289), .B(n17290), .Z(n17261) );
  NANDN U17643 ( .A(n17211), .B(n17210), .Z(n17215) );
  OR U17644 ( .A(n17213), .B(n17212), .Z(n17214) );
  AND U17645 ( .A(n17215), .B(n17214), .Z(n17260) );
  XNOR U17646 ( .A(n17261), .B(n17260), .Z(n17263) );
  NAND U17647 ( .A(n17216), .B(n19724), .Z(n17218) );
  XOR U17648 ( .A(b[11]), .B(a[221]), .Z(n17293) );
  NAND U17649 ( .A(n19692), .B(n17293), .Z(n17217) );
  AND U17650 ( .A(n17218), .B(n17217), .Z(n17304) );
  NAND U17651 ( .A(n19838), .B(n17219), .Z(n17221) );
  XOR U17652 ( .A(b[15]), .B(a[217]), .Z(n17296) );
  NAND U17653 ( .A(n19805), .B(n17296), .Z(n17220) );
  AND U17654 ( .A(n17221), .B(n17220), .Z(n17303) );
  NAND U17655 ( .A(n35), .B(n17222), .Z(n17224) );
  XOR U17656 ( .A(b[9]), .B(a[223]), .Z(n17299) );
  NAND U17657 ( .A(n19598), .B(n17299), .Z(n17223) );
  NAND U17658 ( .A(n17224), .B(n17223), .Z(n17302) );
  XOR U17659 ( .A(n17303), .B(n17302), .Z(n17305) );
  XOR U17660 ( .A(n17304), .B(n17305), .Z(n17315) );
  NANDN U17661 ( .A(n17226), .B(n17225), .Z(n17230) );
  OR U17662 ( .A(n17228), .B(n17227), .Z(n17229) );
  AND U17663 ( .A(n17230), .B(n17229), .Z(n17314) );
  XNOR U17664 ( .A(n17315), .B(n17314), .Z(n17316) );
  NANDN U17665 ( .A(n17232), .B(n17231), .Z(n17236) );
  NANDN U17666 ( .A(n17234), .B(n17233), .Z(n17235) );
  NAND U17667 ( .A(n17236), .B(n17235), .Z(n17317) );
  XNOR U17668 ( .A(n17316), .B(n17317), .Z(n17262) );
  XOR U17669 ( .A(n17263), .B(n17262), .Z(n17321) );
  NANDN U17670 ( .A(n17238), .B(n17237), .Z(n17242) );
  NANDN U17671 ( .A(n17240), .B(n17239), .Z(n17241) );
  AND U17672 ( .A(n17242), .B(n17241), .Z(n17320) );
  XNOR U17673 ( .A(n17321), .B(n17320), .Z(n17322) );
  XOR U17674 ( .A(n17323), .B(n17322), .Z(n17255) );
  NANDN U17675 ( .A(n17244), .B(n17243), .Z(n17248) );
  NAND U17676 ( .A(n17246), .B(n17245), .Z(n17247) );
  AND U17677 ( .A(n17248), .B(n17247), .Z(n17254) );
  XNOR U17678 ( .A(n17255), .B(n17254), .Z(n17256) );
  XNOR U17679 ( .A(n17257), .B(n17256), .Z(n17326) );
  XNOR U17680 ( .A(sreg[471]), .B(n17326), .Z(n17328) );
  NANDN U17681 ( .A(sreg[470]), .B(n17249), .Z(n17253) );
  NAND U17682 ( .A(n17251), .B(n17250), .Z(n17252) );
  NAND U17683 ( .A(n17253), .B(n17252), .Z(n17327) );
  XNOR U17684 ( .A(n17328), .B(n17327), .Z(c[471]) );
  NANDN U17685 ( .A(n17255), .B(n17254), .Z(n17259) );
  NANDN U17686 ( .A(n17257), .B(n17256), .Z(n17258) );
  AND U17687 ( .A(n17259), .B(n17258), .Z(n17334) );
  NANDN U17688 ( .A(n17261), .B(n17260), .Z(n17265) );
  NAND U17689 ( .A(n17263), .B(n17262), .Z(n17264) );
  AND U17690 ( .A(n17265), .B(n17264), .Z(n17400) );
  NANDN U17691 ( .A(n17267), .B(n17266), .Z(n17271) );
  NANDN U17692 ( .A(n17269), .B(n17268), .Z(n17270) );
  AND U17693 ( .A(n17271), .B(n17270), .Z(n17366) );
  NAND U17694 ( .A(n19808), .B(n17272), .Z(n17274) );
  XOR U17695 ( .A(b[13]), .B(a[220]), .Z(n17352) );
  NAND U17696 ( .A(n19768), .B(n17352), .Z(n17273) );
  AND U17697 ( .A(n17274), .B(n17273), .Z(n17344) );
  AND U17698 ( .A(b[15]), .B(a[216]), .Z(n17343) );
  XNOR U17699 ( .A(n17344), .B(n17343), .Z(n17345) );
  NAND U17700 ( .A(b[0]), .B(a[232]), .Z(n17275) );
  XNOR U17701 ( .A(b[1]), .B(n17275), .Z(n17277) );
  NANDN U17702 ( .A(b[0]), .B(a[231]), .Z(n17276) );
  NAND U17703 ( .A(n17277), .B(n17276), .Z(n17346) );
  XNOR U17704 ( .A(n17345), .B(n17346), .Z(n17364) );
  NAND U17705 ( .A(n33), .B(n17278), .Z(n17280) );
  XOR U17706 ( .A(b[5]), .B(a[228]), .Z(n17355) );
  NAND U17707 ( .A(n19342), .B(n17355), .Z(n17279) );
  AND U17708 ( .A(n17280), .B(n17279), .Z(n17388) );
  NAND U17709 ( .A(n34), .B(n17281), .Z(n17283) );
  XOR U17710 ( .A(b[7]), .B(a[226]), .Z(n17358) );
  NAND U17711 ( .A(n19486), .B(n17358), .Z(n17282) );
  AND U17712 ( .A(n17283), .B(n17282), .Z(n17386) );
  NAND U17713 ( .A(n31), .B(n17284), .Z(n17286) );
  XOR U17714 ( .A(b[3]), .B(a[230]), .Z(n17361) );
  NAND U17715 ( .A(n32), .B(n17361), .Z(n17285) );
  NAND U17716 ( .A(n17286), .B(n17285), .Z(n17385) );
  XNOR U17717 ( .A(n17386), .B(n17385), .Z(n17387) );
  XOR U17718 ( .A(n17388), .B(n17387), .Z(n17365) );
  XOR U17719 ( .A(n17364), .B(n17365), .Z(n17367) );
  XOR U17720 ( .A(n17366), .B(n17367), .Z(n17338) );
  NANDN U17721 ( .A(n17288), .B(n17287), .Z(n17292) );
  OR U17722 ( .A(n17290), .B(n17289), .Z(n17291) );
  AND U17723 ( .A(n17292), .B(n17291), .Z(n17337) );
  XNOR U17724 ( .A(n17338), .B(n17337), .Z(n17340) );
  NAND U17725 ( .A(n17293), .B(n19724), .Z(n17295) );
  XOR U17726 ( .A(b[11]), .B(a[222]), .Z(n17370) );
  NAND U17727 ( .A(n19692), .B(n17370), .Z(n17294) );
  AND U17728 ( .A(n17295), .B(n17294), .Z(n17381) );
  NAND U17729 ( .A(n19838), .B(n17296), .Z(n17298) );
  XOR U17730 ( .A(b[15]), .B(a[218]), .Z(n17373) );
  NAND U17731 ( .A(n19805), .B(n17373), .Z(n17297) );
  AND U17732 ( .A(n17298), .B(n17297), .Z(n17380) );
  NAND U17733 ( .A(n35), .B(n17299), .Z(n17301) );
  XOR U17734 ( .A(b[9]), .B(a[224]), .Z(n17376) );
  NAND U17735 ( .A(n19598), .B(n17376), .Z(n17300) );
  NAND U17736 ( .A(n17301), .B(n17300), .Z(n17379) );
  XOR U17737 ( .A(n17380), .B(n17379), .Z(n17382) );
  XOR U17738 ( .A(n17381), .B(n17382), .Z(n17392) );
  NANDN U17739 ( .A(n17303), .B(n17302), .Z(n17307) );
  OR U17740 ( .A(n17305), .B(n17304), .Z(n17306) );
  AND U17741 ( .A(n17307), .B(n17306), .Z(n17391) );
  XNOR U17742 ( .A(n17392), .B(n17391), .Z(n17393) );
  NANDN U17743 ( .A(n17309), .B(n17308), .Z(n17313) );
  NANDN U17744 ( .A(n17311), .B(n17310), .Z(n17312) );
  NAND U17745 ( .A(n17313), .B(n17312), .Z(n17394) );
  XNOR U17746 ( .A(n17393), .B(n17394), .Z(n17339) );
  XOR U17747 ( .A(n17340), .B(n17339), .Z(n17398) );
  NANDN U17748 ( .A(n17315), .B(n17314), .Z(n17319) );
  NANDN U17749 ( .A(n17317), .B(n17316), .Z(n17318) );
  AND U17750 ( .A(n17319), .B(n17318), .Z(n17397) );
  XNOR U17751 ( .A(n17398), .B(n17397), .Z(n17399) );
  XOR U17752 ( .A(n17400), .B(n17399), .Z(n17332) );
  NANDN U17753 ( .A(n17321), .B(n17320), .Z(n17325) );
  NAND U17754 ( .A(n17323), .B(n17322), .Z(n17324) );
  AND U17755 ( .A(n17325), .B(n17324), .Z(n17331) );
  XNOR U17756 ( .A(n17332), .B(n17331), .Z(n17333) );
  XNOR U17757 ( .A(n17334), .B(n17333), .Z(n17403) );
  XNOR U17758 ( .A(sreg[472]), .B(n17403), .Z(n17405) );
  NANDN U17759 ( .A(sreg[471]), .B(n17326), .Z(n17330) );
  NAND U17760 ( .A(n17328), .B(n17327), .Z(n17329) );
  NAND U17761 ( .A(n17330), .B(n17329), .Z(n17404) );
  XNOR U17762 ( .A(n17405), .B(n17404), .Z(c[472]) );
  NANDN U17763 ( .A(n17332), .B(n17331), .Z(n17336) );
  NANDN U17764 ( .A(n17334), .B(n17333), .Z(n17335) );
  AND U17765 ( .A(n17336), .B(n17335), .Z(n17411) );
  NANDN U17766 ( .A(n17338), .B(n17337), .Z(n17342) );
  NAND U17767 ( .A(n17340), .B(n17339), .Z(n17341) );
  AND U17768 ( .A(n17342), .B(n17341), .Z(n17474) );
  NANDN U17769 ( .A(n17344), .B(n17343), .Z(n17348) );
  NANDN U17770 ( .A(n17346), .B(n17345), .Z(n17347) );
  AND U17771 ( .A(n17348), .B(n17347), .Z(n17440) );
  NAND U17772 ( .A(b[0]), .B(a[233]), .Z(n17349) );
  XNOR U17773 ( .A(b[1]), .B(n17349), .Z(n17351) );
  NANDN U17774 ( .A(b[0]), .B(a[232]), .Z(n17350) );
  NAND U17775 ( .A(n17351), .B(n17350), .Z(n17423) );
  NAND U17776 ( .A(n19808), .B(n17352), .Z(n17354) );
  XOR U17777 ( .A(b[13]), .B(a[221]), .Z(n17426) );
  NAND U17778 ( .A(n19768), .B(n17426), .Z(n17353) );
  AND U17779 ( .A(n17354), .B(n17353), .Z(n17421) );
  AND U17780 ( .A(b[15]), .B(a[217]), .Z(n17420) );
  XNOR U17781 ( .A(n17421), .B(n17420), .Z(n17422) );
  XNOR U17782 ( .A(n17423), .B(n17422), .Z(n17438) );
  NAND U17783 ( .A(n33), .B(n17355), .Z(n17357) );
  XOR U17784 ( .A(b[5]), .B(a[229]), .Z(n17429) );
  NAND U17785 ( .A(n19342), .B(n17429), .Z(n17356) );
  AND U17786 ( .A(n17357), .B(n17356), .Z(n17462) );
  NAND U17787 ( .A(n34), .B(n17358), .Z(n17360) );
  XOR U17788 ( .A(b[7]), .B(a[227]), .Z(n17432) );
  NAND U17789 ( .A(n19486), .B(n17432), .Z(n17359) );
  AND U17790 ( .A(n17360), .B(n17359), .Z(n17460) );
  NAND U17791 ( .A(n31), .B(n17361), .Z(n17363) );
  XOR U17792 ( .A(b[3]), .B(a[231]), .Z(n17435) );
  NAND U17793 ( .A(n32), .B(n17435), .Z(n17362) );
  NAND U17794 ( .A(n17363), .B(n17362), .Z(n17459) );
  XNOR U17795 ( .A(n17460), .B(n17459), .Z(n17461) );
  XOR U17796 ( .A(n17462), .B(n17461), .Z(n17439) );
  XOR U17797 ( .A(n17438), .B(n17439), .Z(n17441) );
  XOR U17798 ( .A(n17440), .B(n17441), .Z(n17415) );
  NANDN U17799 ( .A(n17365), .B(n17364), .Z(n17369) );
  OR U17800 ( .A(n17367), .B(n17366), .Z(n17368) );
  AND U17801 ( .A(n17369), .B(n17368), .Z(n17414) );
  XNOR U17802 ( .A(n17415), .B(n17414), .Z(n17417) );
  NAND U17803 ( .A(n17370), .B(n19724), .Z(n17372) );
  XOR U17804 ( .A(b[11]), .B(a[223]), .Z(n17444) );
  NAND U17805 ( .A(n19692), .B(n17444), .Z(n17371) );
  AND U17806 ( .A(n17372), .B(n17371), .Z(n17455) );
  NAND U17807 ( .A(n19838), .B(n17373), .Z(n17375) );
  XOR U17808 ( .A(b[15]), .B(a[219]), .Z(n17447) );
  NAND U17809 ( .A(n19805), .B(n17447), .Z(n17374) );
  AND U17810 ( .A(n17375), .B(n17374), .Z(n17454) );
  NAND U17811 ( .A(n35), .B(n17376), .Z(n17378) );
  XOR U17812 ( .A(b[9]), .B(a[225]), .Z(n17450) );
  NAND U17813 ( .A(n19598), .B(n17450), .Z(n17377) );
  NAND U17814 ( .A(n17378), .B(n17377), .Z(n17453) );
  XOR U17815 ( .A(n17454), .B(n17453), .Z(n17456) );
  XOR U17816 ( .A(n17455), .B(n17456), .Z(n17466) );
  NANDN U17817 ( .A(n17380), .B(n17379), .Z(n17384) );
  OR U17818 ( .A(n17382), .B(n17381), .Z(n17383) );
  AND U17819 ( .A(n17384), .B(n17383), .Z(n17465) );
  XNOR U17820 ( .A(n17466), .B(n17465), .Z(n17467) );
  NANDN U17821 ( .A(n17386), .B(n17385), .Z(n17390) );
  NANDN U17822 ( .A(n17388), .B(n17387), .Z(n17389) );
  NAND U17823 ( .A(n17390), .B(n17389), .Z(n17468) );
  XNOR U17824 ( .A(n17467), .B(n17468), .Z(n17416) );
  XOR U17825 ( .A(n17417), .B(n17416), .Z(n17472) );
  NANDN U17826 ( .A(n17392), .B(n17391), .Z(n17396) );
  NANDN U17827 ( .A(n17394), .B(n17393), .Z(n17395) );
  AND U17828 ( .A(n17396), .B(n17395), .Z(n17471) );
  XNOR U17829 ( .A(n17472), .B(n17471), .Z(n17473) );
  XOR U17830 ( .A(n17474), .B(n17473), .Z(n17409) );
  NANDN U17831 ( .A(n17398), .B(n17397), .Z(n17402) );
  NAND U17832 ( .A(n17400), .B(n17399), .Z(n17401) );
  AND U17833 ( .A(n17402), .B(n17401), .Z(n17408) );
  XNOR U17834 ( .A(n17409), .B(n17408), .Z(n17410) );
  XNOR U17835 ( .A(n17411), .B(n17410), .Z(n17477) );
  XNOR U17836 ( .A(sreg[473]), .B(n17477), .Z(n17479) );
  NANDN U17837 ( .A(sreg[472]), .B(n17403), .Z(n17407) );
  NAND U17838 ( .A(n17405), .B(n17404), .Z(n17406) );
  NAND U17839 ( .A(n17407), .B(n17406), .Z(n17478) );
  XNOR U17840 ( .A(n17479), .B(n17478), .Z(c[473]) );
  NANDN U17841 ( .A(n17409), .B(n17408), .Z(n17413) );
  NANDN U17842 ( .A(n17411), .B(n17410), .Z(n17412) );
  AND U17843 ( .A(n17413), .B(n17412), .Z(n17485) );
  NANDN U17844 ( .A(n17415), .B(n17414), .Z(n17419) );
  NAND U17845 ( .A(n17417), .B(n17416), .Z(n17418) );
  AND U17846 ( .A(n17419), .B(n17418), .Z(n17551) );
  NANDN U17847 ( .A(n17421), .B(n17420), .Z(n17425) );
  NANDN U17848 ( .A(n17423), .B(n17422), .Z(n17424) );
  AND U17849 ( .A(n17425), .B(n17424), .Z(n17517) );
  NAND U17850 ( .A(n19808), .B(n17426), .Z(n17428) );
  XOR U17851 ( .A(b[13]), .B(a[222]), .Z(n17503) );
  NAND U17852 ( .A(n19768), .B(n17503), .Z(n17427) );
  AND U17853 ( .A(n17428), .B(n17427), .Z(n17495) );
  AND U17854 ( .A(b[15]), .B(a[218]), .Z(n17494) );
  XOR U17855 ( .A(n17495), .B(n17494), .Z(n17497) );
  XNOR U17856 ( .A(n17496), .B(n17497), .Z(n17515) );
  NAND U17857 ( .A(n33), .B(n17429), .Z(n17431) );
  XOR U17858 ( .A(b[5]), .B(a[230]), .Z(n17506) );
  NAND U17859 ( .A(n19342), .B(n17506), .Z(n17430) );
  AND U17860 ( .A(n17431), .B(n17430), .Z(n17539) );
  NAND U17861 ( .A(n34), .B(n17432), .Z(n17434) );
  XOR U17862 ( .A(b[7]), .B(a[228]), .Z(n17509) );
  NAND U17863 ( .A(n19486), .B(n17509), .Z(n17433) );
  AND U17864 ( .A(n17434), .B(n17433), .Z(n17537) );
  NAND U17865 ( .A(n31), .B(n17435), .Z(n17437) );
  XOR U17866 ( .A(b[3]), .B(a[232]), .Z(n17512) );
  NAND U17867 ( .A(n32), .B(n17512), .Z(n17436) );
  NAND U17868 ( .A(n17437), .B(n17436), .Z(n17536) );
  XNOR U17869 ( .A(n17537), .B(n17536), .Z(n17538) );
  XOR U17870 ( .A(n17539), .B(n17538), .Z(n17516) );
  XOR U17871 ( .A(n17515), .B(n17516), .Z(n17518) );
  XOR U17872 ( .A(n17517), .B(n17518), .Z(n17489) );
  NANDN U17873 ( .A(n17439), .B(n17438), .Z(n17443) );
  OR U17874 ( .A(n17441), .B(n17440), .Z(n17442) );
  AND U17875 ( .A(n17443), .B(n17442), .Z(n17488) );
  XNOR U17876 ( .A(n17489), .B(n17488), .Z(n17491) );
  NAND U17877 ( .A(n17444), .B(n19724), .Z(n17446) );
  XOR U17878 ( .A(b[11]), .B(a[224]), .Z(n17521) );
  NAND U17879 ( .A(n19692), .B(n17521), .Z(n17445) );
  AND U17880 ( .A(n17446), .B(n17445), .Z(n17532) );
  NAND U17881 ( .A(n19838), .B(n17447), .Z(n17449) );
  XOR U17882 ( .A(b[15]), .B(a[220]), .Z(n17524) );
  NAND U17883 ( .A(n19805), .B(n17524), .Z(n17448) );
  AND U17884 ( .A(n17449), .B(n17448), .Z(n17531) );
  NAND U17885 ( .A(n35), .B(n17450), .Z(n17452) );
  XOR U17886 ( .A(b[9]), .B(a[226]), .Z(n17527) );
  NAND U17887 ( .A(n19598), .B(n17527), .Z(n17451) );
  NAND U17888 ( .A(n17452), .B(n17451), .Z(n17530) );
  XOR U17889 ( .A(n17531), .B(n17530), .Z(n17533) );
  XOR U17890 ( .A(n17532), .B(n17533), .Z(n17543) );
  NANDN U17891 ( .A(n17454), .B(n17453), .Z(n17458) );
  OR U17892 ( .A(n17456), .B(n17455), .Z(n17457) );
  AND U17893 ( .A(n17458), .B(n17457), .Z(n17542) );
  XNOR U17894 ( .A(n17543), .B(n17542), .Z(n17544) );
  NANDN U17895 ( .A(n17460), .B(n17459), .Z(n17464) );
  NANDN U17896 ( .A(n17462), .B(n17461), .Z(n17463) );
  NAND U17897 ( .A(n17464), .B(n17463), .Z(n17545) );
  XNOR U17898 ( .A(n17544), .B(n17545), .Z(n17490) );
  XOR U17899 ( .A(n17491), .B(n17490), .Z(n17549) );
  NANDN U17900 ( .A(n17466), .B(n17465), .Z(n17470) );
  NANDN U17901 ( .A(n17468), .B(n17467), .Z(n17469) );
  AND U17902 ( .A(n17470), .B(n17469), .Z(n17548) );
  XNOR U17903 ( .A(n17549), .B(n17548), .Z(n17550) );
  XOR U17904 ( .A(n17551), .B(n17550), .Z(n17483) );
  NANDN U17905 ( .A(n17472), .B(n17471), .Z(n17476) );
  NAND U17906 ( .A(n17474), .B(n17473), .Z(n17475) );
  AND U17907 ( .A(n17476), .B(n17475), .Z(n17482) );
  XNOR U17908 ( .A(n17483), .B(n17482), .Z(n17484) );
  XNOR U17909 ( .A(n17485), .B(n17484), .Z(n17554) );
  XNOR U17910 ( .A(sreg[474]), .B(n17554), .Z(n17556) );
  NANDN U17911 ( .A(sreg[473]), .B(n17477), .Z(n17481) );
  NAND U17912 ( .A(n17479), .B(n17478), .Z(n17480) );
  NAND U17913 ( .A(n17481), .B(n17480), .Z(n17555) );
  XNOR U17914 ( .A(n17556), .B(n17555), .Z(c[474]) );
  NANDN U17915 ( .A(n17483), .B(n17482), .Z(n17487) );
  NANDN U17916 ( .A(n17485), .B(n17484), .Z(n17486) );
  AND U17917 ( .A(n17487), .B(n17486), .Z(n17562) );
  NANDN U17918 ( .A(n17489), .B(n17488), .Z(n17493) );
  NAND U17919 ( .A(n17491), .B(n17490), .Z(n17492) );
  AND U17920 ( .A(n17493), .B(n17492), .Z(n17628) );
  NANDN U17921 ( .A(n17495), .B(n17494), .Z(n17499) );
  NANDN U17922 ( .A(n17497), .B(n17496), .Z(n17498) );
  AND U17923 ( .A(n17499), .B(n17498), .Z(n17594) );
  NAND U17924 ( .A(b[0]), .B(a[235]), .Z(n17500) );
  XNOR U17925 ( .A(b[1]), .B(n17500), .Z(n17502) );
  NANDN U17926 ( .A(b[0]), .B(a[234]), .Z(n17501) );
  NAND U17927 ( .A(n17502), .B(n17501), .Z(n17574) );
  NAND U17928 ( .A(n19808), .B(n17503), .Z(n17505) );
  XOR U17929 ( .A(b[13]), .B(a[223]), .Z(n17577) );
  NAND U17930 ( .A(n19768), .B(n17577), .Z(n17504) );
  AND U17931 ( .A(n17505), .B(n17504), .Z(n17572) );
  AND U17932 ( .A(b[15]), .B(a[219]), .Z(n17571) );
  XNOR U17933 ( .A(n17572), .B(n17571), .Z(n17573) );
  XNOR U17934 ( .A(n17574), .B(n17573), .Z(n17592) );
  NAND U17935 ( .A(n33), .B(n17506), .Z(n17508) );
  XOR U17936 ( .A(b[5]), .B(a[231]), .Z(n17583) );
  NAND U17937 ( .A(n19342), .B(n17583), .Z(n17507) );
  AND U17938 ( .A(n17508), .B(n17507), .Z(n17616) );
  NAND U17939 ( .A(n34), .B(n17509), .Z(n17511) );
  XOR U17940 ( .A(b[7]), .B(a[229]), .Z(n17586) );
  NAND U17941 ( .A(n19486), .B(n17586), .Z(n17510) );
  AND U17942 ( .A(n17511), .B(n17510), .Z(n17614) );
  NAND U17943 ( .A(n31), .B(n17512), .Z(n17514) );
  XOR U17944 ( .A(b[3]), .B(a[233]), .Z(n17589) );
  NAND U17945 ( .A(n32), .B(n17589), .Z(n17513) );
  NAND U17946 ( .A(n17514), .B(n17513), .Z(n17613) );
  XNOR U17947 ( .A(n17614), .B(n17613), .Z(n17615) );
  XOR U17948 ( .A(n17616), .B(n17615), .Z(n17593) );
  XOR U17949 ( .A(n17592), .B(n17593), .Z(n17595) );
  XOR U17950 ( .A(n17594), .B(n17595), .Z(n17566) );
  NANDN U17951 ( .A(n17516), .B(n17515), .Z(n17520) );
  OR U17952 ( .A(n17518), .B(n17517), .Z(n17519) );
  AND U17953 ( .A(n17520), .B(n17519), .Z(n17565) );
  XNOR U17954 ( .A(n17566), .B(n17565), .Z(n17568) );
  NAND U17955 ( .A(n17521), .B(n19724), .Z(n17523) );
  XOR U17956 ( .A(b[11]), .B(a[225]), .Z(n17598) );
  NAND U17957 ( .A(n19692), .B(n17598), .Z(n17522) );
  AND U17958 ( .A(n17523), .B(n17522), .Z(n17609) );
  NAND U17959 ( .A(n19838), .B(n17524), .Z(n17526) );
  XOR U17960 ( .A(b[15]), .B(a[221]), .Z(n17601) );
  NAND U17961 ( .A(n19805), .B(n17601), .Z(n17525) );
  AND U17962 ( .A(n17526), .B(n17525), .Z(n17608) );
  NAND U17963 ( .A(n35), .B(n17527), .Z(n17529) );
  XOR U17964 ( .A(b[9]), .B(a[227]), .Z(n17604) );
  NAND U17965 ( .A(n19598), .B(n17604), .Z(n17528) );
  NAND U17966 ( .A(n17529), .B(n17528), .Z(n17607) );
  XOR U17967 ( .A(n17608), .B(n17607), .Z(n17610) );
  XOR U17968 ( .A(n17609), .B(n17610), .Z(n17620) );
  NANDN U17969 ( .A(n17531), .B(n17530), .Z(n17535) );
  OR U17970 ( .A(n17533), .B(n17532), .Z(n17534) );
  AND U17971 ( .A(n17535), .B(n17534), .Z(n17619) );
  XNOR U17972 ( .A(n17620), .B(n17619), .Z(n17621) );
  NANDN U17973 ( .A(n17537), .B(n17536), .Z(n17541) );
  NANDN U17974 ( .A(n17539), .B(n17538), .Z(n17540) );
  NAND U17975 ( .A(n17541), .B(n17540), .Z(n17622) );
  XNOR U17976 ( .A(n17621), .B(n17622), .Z(n17567) );
  XOR U17977 ( .A(n17568), .B(n17567), .Z(n17626) );
  NANDN U17978 ( .A(n17543), .B(n17542), .Z(n17547) );
  NANDN U17979 ( .A(n17545), .B(n17544), .Z(n17546) );
  AND U17980 ( .A(n17547), .B(n17546), .Z(n17625) );
  XNOR U17981 ( .A(n17626), .B(n17625), .Z(n17627) );
  XOR U17982 ( .A(n17628), .B(n17627), .Z(n17560) );
  NANDN U17983 ( .A(n17549), .B(n17548), .Z(n17553) );
  NAND U17984 ( .A(n17551), .B(n17550), .Z(n17552) );
  AND U17985 ( .A(n17553), .B(n17552), .Z(n17559) );
  XNOR U17986 ( .A(n17560), .B(n17559), .Z(n17561) );
  XNOR U17987 ( .A(n17562), .B(n17561), .Z(n17631) );
  XNOR U17988 ( .A(sreg[475]), .B(n17631), .Z(n17633) );
  NANDN U17989 ( .A(sreg[474]), .B(n17554), .Z(n17558) );
  NAND U17990 ( .A(n17556), .B(n17555), .Z(n17557) );
  NAND U17991 ( .A(n17558), .B(n17557), .Z(n17632) );
  XNOR U17992 ( .A(n17633), .B(n17632), .Z(c[475]) );
  NANDN U17993 ( .A(n17560), .B(n17559), .Z(n17564) );
  NANDN U17994 ( .A(n17562), .B(n17561), .Z(n17563) );
  AND U17995 ( .A(n17564), .B(n17563), .Z(n17639) );
  NANDN U17996 ( .A(n17566), .B(n17565), .Z(n17570) );
  NAND U17997 ( .A(n17568), .B(n17567), .Z(n17569) );
  AND U17998 ( .A(n17570), .B(n17569), .Z(n17705) );
  NANDN U17999 ( .A(n17572), .B(n17571), .Z(n17576) );
  NANDN U18000 ( .A(n17574), .B(n17573), .Z(n17575) );
  AND U18001 ( .A(n17576), .B(n17575), .Z(n17671) );
  NAND U18002 ( .A(n19808), .B(n17577), .Z(n17579) );
  XOR U18003 ( .A(b[13]), .B(a[224]), .Z(n17657) );
  NAND U18004 ( .A(n19768), .B(n17657), .Z(n17578) );
  AND U18005 ( .A(n17579), .B(n17578), .Z(n17649) );
  AND U18006 ( .A(b[15]), .B(a[220]), .Z(n17648) );
  XNOR U18007 ( .A(n17649), .B(n17648), .Z(n17650) );
  NAND U18008 ( .A(b[0]), .B(a[236]), .Z(n17580) );
  XNOR U18009 ( .A(b[1]), .B(n17580), .Z(n17582) );
  NANDN U18010 ( .A(b[0]), .B(a[235]), .Z(n17581) );
  NAND U18011 ( .A(n17582), .B(n17581), .Z(n17651) );
  XNOR U18012 ( .A(n17650), .B(n17651), .Z(n17669) );
  NAND U18013 ( .A(n33), .B(n17583), .Z(n17585) );
  XOR U18014 ( .A(b[5]), .B(a[232]), .Z(n17660) );
  NAND U18015 ( .A(n19342), .B(n17660), .Z(n17584) );
  AND U18016 ( .A(n17585), .B(n17584), .Z(n17693) );
  NAND U18017 ( .A(n34), .B(n17586), .Z(n17588) );
  XOR U18018 ( .A(b[7]), .B(a[230]), .Z(n17663) );
  NAND U18019 ( .A(n19486), .B(n17663), .Z(n17587) );
  AND U18020 ( .A(n17588), .B(n17587), .Z(n17691) );
  NAND U18021 ( .A(n31), .B(n17589), .Z(n17591) );
  XOR U18022 ( .A(b[3]), .B(a[234]), .Z(n17666) );
  NAND U18023 ( .A(n32), .B(n17666), .Z(n17590) );
  NAND U18024 ( .A(n17591), .B(n17590), .Z(n17690) );
  XNOR U18025 ( .A(n17691), .B(n17690), .Z(n17692) );
  XOR U18026 ( .A(n17693), .B(n17692), .Z(n17670) );
  XOR U18027 ( .A(n17669), .B(n17670), .Z(n17672) );
  XOR U18028 ( .A(n17671), .B(n17672), .Z(n17643) );
  NANDN U18029 ( .A(n17593), .B(n17592), .Z(n17597) );
  OR U18030 ( .A(n17595), .B(n17594), .Z(n17596) );
  AND U18031 ( .A(n17597), .B(n17596), .Z(n17642) );
  XNOR U18032 ( .A(n17643), .B(n17642), .Z(n17645) );
  NAND U18033 ( .A(n17598), .B(n19724), .Z(n17600) );
  XOR U18034 ( .A(b[11]), .B(a[226]), .Z(n17675) );
  NAND U18035 ( .A(n19692), .B(n17675), .Z(n17599) );
  AND U18036 ( .A(n17600), .B(n17599), .Z(n17686) );
  NAND U18037 ( .A(n19838), .B(n17601), .Z(n17603) );
  XOR U18038 ( .A(b[15]), .B(a[222]), .Z(n17678) );
  NAND U18039 ( .A(n19805), .B(n17678), .Z(n17602) );
  AND U18040 ( .A(n17603), .B(n17602), .Z(n17685) );
  NAND U18041 ( .A(n35), .B(n17604), .Z(n17606) );
  XOR U18042 ( .A(b[9]), .B(a[228]), .Z(n17681) );
  NAND U18043 ( .A(n19598), .B(n17681), .Z(n17605) );
  NAND U18044 ( .A(n17606), .B(n17605), .Z(n17684) );
  XOR U18045 ( .A(n17685), .B(n17684), .Z(n17687) );
  XOR U18046 ( .A(n17686), .B(n17687), .Z(n17697) );
  NANDN U18047 ( .A(n17608), .B(n17607), .Z(n17612) );
  OR U18048 ( .A(n17610), .B(n17609), .Z(n17611) );
  AND U18049 ( .A(n17612), .B(n17611), .Z(n17696) );
  XNOR U18050 ( .A(n17697), .B(n17696), .Z(n17698) );
  NANDN U18051 ( .A(n17614), .B(n17613), .Z(n17618) );
  NANDN U18052 ( .A(n17616), .B(n17615), .Z(n17617) );
  NAND U18053 ( .A(n17618), .B(n17617), .Z(n17699) );
  XNOR U18054 ( .A(n17698), .B(n17699), .Z(n17644) );
  XOR U18055 ( .A(n17645), .B(n17644), .Z(n17703) );
  NANDN U18056 ( .A(n17620), .B(n17619), .Z(n17624) );
  NANDN U18057 ( .A(n17622), .B(n17621), .Z(n17623) );
  AND U18058 ( .A(n17624), .B(n17623), .Z(n17702) );
  XNOR U18059 ( .A(n17703), .B(n17702), .Z(n17704) );
  XOR U18060 ( .A(n17705), .B(n17704), .Z(n17637) );
  NANDN U18061 ( .A(n17626), .B(n17625), .Z(n17630) );
  NAND U18062 ( .A(n17628), .B(n17627), .Z(n17629) );
  AND U18063 ( .A(n17630), .B(n17629), .Z(n17636) );
  XNOR U18064 ( .A(n17637), .B(n17636), .Z(n17638) );
  XNOR U18065 ( .A(n17639), .B(n17638), .Z(n17708) );
  XNOR U18066 ( .A(sreg[476]), .B(n17708), .Z(n17710) );
  NANDN U18067 ( .A(sreg[475]), .B(n17631), .Z(n17635) );
  NAND U18068 ( .A(n17633), .B(n17632), .Z(n17634) );
  NAND U18069 ( .A(n17635), .B(n17634), .Z(n17709) );
  XNOR U18070 ( .A(n17710), .B(n17709), .Z(c[476]) );
  NANDN U18071 ( .A(n17637), .B(n17636), .Z(n17641) );
  NANDN U18072 ( .A(n17639), .B(n17638), .Z(n17640) );
  AND U18073 ( .A(n17641), .B(n17640), .Z(n17716) );
  NANDN U18074 ( .A(n17643), .B(n17642), .Z(n17647) );
  NAND U18075 ( .A(n17645), .B(n17644), .Z(n17646) );
  AND U18076 ( .A(n17647), .B(n17646), .Z(n17782) );
  NANDN U18077 ( .A(n17649), .B(n17648), .Z(n17653) );
  NANDN U18078 ( .A(n17651), .B(n17650), .Z(n17652) );
  AND U18079 ( .A(n17653), .B(n17652), .Z(n17748) );
  NAND U18080 ( .A(b[0]), .B(a[237]), .Z(n17654) );
  XNOR U18081 ( .A(b[1]), .B(n17654), .Z(n17656) );
  NANDN U18082 ( .A(b[0]), .B(a[236]), .Z(n17655) );
  NAND U18083 ( .A(n17656), .B(n17655), .Z(n17728) );
  NAND U18084 ( .A(n19808), .B(n17657), .Z(n17659) );
  XOR U18085 ( .A(b[13]), .B(a[225]), .Z(n17734) );
  NAND U18086 ( .A(n19768), .B(n17734), .Z(n17658) );
  AND U18087 ( .A(n17659), .B(n17658), .Z(n17726) );
  AND U18088 ( .A(b[15]), .B(a[221]), .Z(n17725) );
  XNOR U18089 ( .A(n17726), .B(n17725), .Z(n17727) );
  XNOR U18090 ( .A(n17728), .B(n17727), .Z(n17746) );
  NAND U18091 ( .A(n33), .B(n17660), .Z(n17662) );
  XOR U18092 ( .A(b[5]), .B(a[233]), .Z(n17737) );
  NAND U18093 ( .A(n19342), .B(n17737), .Z(n17661) );
  AND U18094 ( .A(n17662), .B(n17661), .Z(n17770) );
  NAND U18095 ( .A(n34), .B(n17663), .Z(n17665) );
  XOR U18096 ( .A(b[7]), .B(a[231]), .Z(n17740) );
  NAND U18097 ( .A(n19486), .B(n17740), .Z(n17664) );
  AND U18098 ( .A(n17665), .B(n17664), .Z(n17768) );
  NAND U18099 ( .A(n31), .B(n17666), .Z(n17668) );
  XOR U18100 ( .A(b[3]), .B(a[235]), .Z(n17743) );
  NAND U18101 ( .A(n32), .B(n17743), .Z(n17667) );
  NAND U18102 ( .A(n17668), .B(n17667), .Z(n17767) );
  XNOR U18103 ( .A(n17768), .B(n17767), .Z(n17769) );
  XOR U18104 ( .A(n17770), .B(n17769), .Z(n17747) );
  XOR U18105 ( .A(n17746), .B(n17747), .Z(n17749) );
  XOR U18106 ( .A(n17748), .B(n17749), .Z(n17720) );
  NANDN U18107 ( .A(n17670), .B(n17669), .Z(n17674) );
  OR U18108 ( .A(n17672), .B(n17671), .Z(n17673) );
  AND U18109 ( .A(n17674), .B(n17673), .Z(n17719) );
  XNOR U18110 ( .A(n17720), .B(n17719), .Z(n17722) );
  NAND U18111 ( .A(n17675), .B(n19724), .Z(n17677) );
  XOR U18112 ( .A(b[11]), .B(a[227]), .Z(n17752) );
  NAND U18113 ( .A(n19692), .B(n17752), .Z(n17676) );
  AND U18114 ( .A(n17677), .B(n17676), .Z(n17763) );
  NAND U18115 ( .A(n19838), .B(n17678), .Z(n17680) );
  XOR U18116 ( .A(b[15]), .B(a[223]), .Z(n17755) );
  NAND U18117 ( .A(n19805), .B(n17755), .Z(n17679) );
  AND U18118 ( .A(n17680), .B(n17679), .Z(n17762) );
  NAND U18119 ( .A(n35), .B(n17681), .Z(n17683) );
  XOR U18120 ( .A(b[9]), .B(a[229]), .Z(n17758) );
  NAND U18121 ( .A(n19598), .B(n17758), .Z(n17682) );
  NAND U18122 ( .A(n17683), .B(n17682), .Z(n17761) );
  XOR U18123 ( .A(n17762), .B(n17761), .Z(n17764) );
  XOR U18124 ( .A(n17763), .B(n17764), .Z(n17774) );
  NANDN U18125 ( .A(n17685), .B(n17684), .Z(n17689) );
  OR U18126 ( .A(n17687), .B(n17686), .Z(n17688) );
  AND U18127 ( .A(n17689), .B(n17688), .Z(n17773) );
  XNOR U18128 ( .A(n17774), .B(n17773), .Z(n17775) );
  NANDN U18129 ( .A(n17691), .B(n17690), .Z(n17695) );
  NANDN U18130 ( .A(n17693), .B(n17692), .Z(n17694) );
  NAND U18131 ( .A(n17695), .B(n17694), .Z(n17776) );
  XNOR U18132 ( .A(n17775), .B(n17776), .Z(n17721) );
  XOR U18133 ( .A(n17722), .B(n17721), .Z(n17780) );
  NANDN U18134 ( .A(n17697), .B(n17696), .Z(n17701) );
  NANDN U18135 ( .A(n17699), .B(n17698), .Z(n17700) );
  AND U18136 ( .A(n17701), .B(n17700), .Z(n17779) );
  XNOR U18137 ( .A(n17780), .B(n17779), .Z(n17781) );
  XOR U18138 ( .A(n17782), .B(n17781), .Z(n17714) );
  NANDN U18139 ( .A(n17703), .B(n17702), .Z(n17707) );
  NAND U18140 ( .A(n17705), .B(n17704), .Z(n17706) );
  AND U18141 ( .A(n17707), .B(n17706), .Z(n17713) );
  XNOR U18142 ( .A(n17714), .B(n17713), .Z(n17715) );
  XNOR U18143 ( .A(n17716), .B(n17715), .Z(n17785) );
  XNOR U18144 ( .A(sreg[477]), .B(n17785), .Z(n17787) );
  NANDN U18145 ( .A(sreg[476]), .B(n17708), .Z(n17712) );
  NAND U18146 ( .A(n17710), .B(n17709), .Z(n17711) );
  NAND U18147 ( .A(n17712), .B(n17711), .Z(n17786) );
  XNOR U18148 ( .A(n17787), .B(n17786), .Z(c[477]) );
  NANDN U18149 ( .A(n17714), .B(n17713), .Z(n17718) );
  NANDN U18150 ( .A(n17716), .B(n17715), .Z(n17717) );
  AND U18151 ( .A(n17718), .B(n17717), .Z(n17793) );
  NANDN U18152 ( .A(n17720), .B(n17719), .Z(n17724) );
  NAND U18153 ( .A(n17722), .B(n17721), .Z(n17723) );
  AND U18154 ( .A(n17724), .B(n17723), .Z(n17859) );
  NANDN U18155 ( .A(n17726), .B(n17725), .Z(n17730) );
  NANDN U18156 ( .A(n17728), .B(n17727), .Z(n17729) );
  AND U18157 ( .A(n17730), .B(n17729), .Z(n17825) );
  NAND U18158 ( .A(b[0]), .B(a[238]), .Z(n17731) );
  XNOR U18159 ( .A(b[1]), .B(n17731), .Z(n17733) );
  NANDN U18160 ( .A(b[0]), .B(a[237]), .Z(n17732) );
  NAND U18161 ( .A(n17733), .B(n17732), .Z(n17805) );
  NAND U18162 ( .A(n19808), .B(n17734), .Z(n17736) );
  XOR U18163 ( .A(b[13]), .B(a[226]), .Z(n17811) );
  NAND U18164 ( .A(n19768), .B(n17811), .Z(n17735) );
  AND U18165 ( .A(n17736), .B(n17735), .Z(n17803) );
  AND U18166 ( .A(b[15]), .B(a[222]), .Z(n17802) );
  XNOR U18167 ( .A(n17803), .B(n17802), .Z(n17804) );
  XNOR U18168 ( .A(n17805), .B(n17804), .Z(n17823) );
  NAND U18169 ( .A(n33), .B(n17737), .Z(n17739) );
  XOR U18170 ( .A(b[5]), .B(a[234]), .Z(n17814) );
  NAND U18171 ( .A(n19342), .B(n17814), .Z(n17738) );
  AND U18172 ( .A(n17739), .B(n17738), .Z(n17847) );
  NAND U18173 ( .A(n34), .B(n17740), .Z(n17742) );
  XOR U18174 ( .A(b[7]), .B(a[232]), .Z(n17817) );
  NAND U18175 ( .A(n19486), .B(n17817), .Z(n17741) );
  AND U18176 ( .A(n17742), .B(n17741), .Z(n17845) );
  NAND U18177 ( .A(n31), .B(n17743), .Z(n17745) );
  XOR U18178 ( .A(b[3]), .B(a[236]), .Z(n17820) );
  NAND U18179 ( .A(n32), .B(n17820), .Z(n17744) );
  NAND U18180 ( .A(n17745), .B(n17744), .Z(n17844) );
  XNOR U18181 ( .A(n17845), .B(n17844), .Z(n17846) );
  XOR U18182 ( .A(n17847), .B(n17846), .Z(n17824) );
  XOR U18183 ( .A(n17823), .B(n17824), .Z(n17826) );
  XOR U18184 ( .A(n17825), .B(n17826), .Z(n17797) );
  NANDN U18185 ( .A(n17747), .B(n17746), .Z(n17751) );
  OR U18186 ( .A(n17749), .B(n17748), .Z(n17750) );
  AND U18187 ( .A(n17751), .B(n17750), .Z(n17796) );
  XNOR U18188 ( .A(n17797), .B(n17796), .Z(n17799) );
  NAND U18189 ( .A(n17752), .B(n19724), .Z(n17754) );
  XOR U18190 ( .A(b[11]), .B(a[228]), .Z(n17829) );
  NAND U18191 ( .A(n19692), .B(n17829), .Z(n17753) );
  AND U18192 ( .A(n17754), .B(n17753), .Z(n17840) );
  NAND U18193 ( .A(n19838), .B(n17755), .Z(n17757) );
  XOR U18194 ( .A(b[15]), .B(a[224]), .Z(n17832) );
  NAND U18195 ( .A(n19805), .B(n17832), .Z(n17756) );
  AND U18196 ( .A(n17757), .B(n17756), .Z(n17839) );
  NAND U18197 ( .A(n35), .B(n17758), .Z(n17760) );
  XOR U18198 ( .A(b[9]), .B(a[230]), .Z(n17835) );
  NAND U18199 ( .A(n19598), .B(n17835), .Z(n17759) );
  NAND U18200 ( .A(n17760), .B(n17759), .Z(n17838) );
  XOR U18201 ( .A(n17839), .B(n17838), .Z(n17841) );
  XOR U18202 ( .A(n17840), .B(n17841), .Z(n17851) );
  NANDN U18203 ( .A(n17762), .B(n17761), .Z(n17766) );
  OR U18204 ( .A(n17764), .B(n17763), .Z(n17765) );
  AND U18205 ( .A(n17766), .B(n17765), .Z(n17850) );
  XNOR U18206 ( .A(n17851), .B(n17850), .Z(n17852) );
  NANDN U18207 ( .A(n17768), .B(n17767), .Z(n17772) );
  NANDN U18208 ( .A(n17770), .B(n17769), .Z(n17771) );
  NAND U18209 ( .A(n17772), .B(n17771), .Z(n17853) );
  XNOR U18210 ( .A(n17852), .B(n17853), .Z(n17798) );
  XOR U18211 ( .A(n17799), .B(n17798), .Z(n17857) );
  NANDN U18212 ( .A(n17774), .B(n17773), .Z(n17778) );
  NANDN U18213 ( .A(n17776), .B(n17775), .Z(n17777) );
  AND U18214 ( .A(n17778), .B(n17777), .Z(n17856) );
  XNOR U18215 ( .A(n17857), .B(n17856), .Z(n17858) );
  XOR U18216 ( .A(n17859), .B(n17858), .Z(n17791) );
  NANDN U18217 ( .A(n17780), .B(n17779), .Z(n17784) );
  NAND U18218 ( .A(n17782), .B(n17781), .Z(n17783) );
  AND U18219 ( .A(n17784), .B(n17783), .Z(n17790) );
  XNOR U18220 ( .A(n17791), .B(n17790), .Z(n17792) );
  XNOR U18221 ( .A(n17793), .B(n17792), .Z(n17862) );
  XNOR U18222 ( .A(sreg[478]), .B(n17862), .Z(n17864) );
  NANDN U18223 ( .A(sreg[477]), .B(n17785), .Z(n17789) );
  NAND U18224 ( .A(n17787), .B(n17786), .Z(n17788) );
  NAND U18225 ( .A(n17789), .B(n17788), .Z(n17863) );
  XNOR U18226 ( .A(n17864), .B(n17863), .Z(c[478]) );
  NANDN U18227 ( .A(n17791), .B(n17790), .Z(n17795) );
  NANDN U18228 ( .A(n17793), .B(n17792), .Z(n17794) );
  AND U18229 ( .A(n17795), .B(n17794), .Z(n17870) );
  NANDN U18230 ( .A(n17797), .B(n17796), .Z(n17801) );
  NAND U18231 ( .A(n17799), .B(n17798), .Z(n17800) );
  AND U18232 ( .A(n17801), .B(n17800), .Z(n17936) );
  NANDN U18233 ( .A(n17803), .B(n17802), .Z(n17807) );
  NANDN U18234 ( .A(n17805), .B(n17804), .Z(n17806) );
  AND U18235 ( .A(n17807), .B(n17806), .Z(n17902) );
  NAND U18236 ( .A(b[0]), .B(a[239]), .Z(n17808) );
  XNOR U18237 ( .A(b[1]), .B(n17808), .Z(n17810) );
  NANDN U18238 ( .A(b[0]), .B(a[238]), .Z(n17809) );
  NAND U18239 ( .A(n17810), .B(n17809), .Z(n17882) );
  NAND U18240 ( .A(n19808), .B(n17811), .Z(n17813) );
  XOR U18241 ( .A(b[13]), .B(a[227]), .Z(n17885) );
  NAND U18242 ( .A(n19768), .B(n17885), .Z(n17812) );
  AND U18243 ( .A(n17813), .B(n17812), .Z(n17880) );
  AND U18244 ( .A(b[15]), .B(a[223]), .Z(n17879) );
  XNOR U18245 ( .A(n17880), .B(n17879), .Z(n17881) );
  XNOR U18246 ( .A(n17882), .B(n17881), .Z(n17900) );
  NAND U18247 ( .A(n33), .B(n17814), .Z(n17816) );
  XOR U18248 ( .A(b[5]), .B(a[235]), .Z(n17891) );
  NAND U18249 ( .A(n19342), .B(n17891), .Z(n17815) );
  AND U18250 ( .A(n17816), .B(n17815), .Z(n17924) );
  NAND U18251 ( .A(n34), .B(n17817), .Z(n17819) );
  XOR U18252 ( .A(b[7]), .B(a[233]), .Z(n17894) );
  NAND U18253 ( .A(n19486), .B(n17894), .Z(n17818) );
  AND U18254 ( .A(n17819), .B(n17818), .Z(n17922) );
  NAND U18255 ( .A(n31), .B(n17820), .Z(n17822) );
  XOR U18256 ( .A(b[3]), .B(a[237]), .Z(n17897) );
  NAND U18257 ( .A(n32), .B(n17897), .Z(n17821) );
  NAND U18258 ( .A(n17822), .B(n17821), .Z(n17921) );
  XNOR U18259 ( .A(n17922), .B(n17921), .Z(n17923) );
  XOR U18260 ( .A(n17924), .B(n17923), .Z(n17901) );
  XOR U18261 ( .A(n17900), .B(n17901), .Z(n17903) );
  XOR U18262 ( .A(n17902), .B(n17903), .Z(n17874) );
  NANDN U18263 ( .A(n17824), .B(n17823), .Z(n17828) );
  OR U18264 ( .A(n17826), .B(n17825), .Z(n17827) );
  AND U18265 ( .A(n17828), .B(n17827), .Z(n17873) );
  XNOR U18266 ( .A(n17874), .B(n17873), .Z(n17876) );
  NAND U18267 ( .A(n17829), .B(n19724), .Z(n17831) );
  XOR U18268 ( .A(b[11]), .B(a[229]), .Z(n17906) );
  NAND U18269 ( .A(n19692), .B(n17906), .Z(n17830) );
  AND U18270 ( .A(n17831), .B(n17830), .Z(n17917) );
  NAND U18271 ( .A(n19838), .B(n17832), .Z(n17834) );
  XOR U18272 ( .A(b[15]), .B(a[225]), .Z(n17909) );
  NAND U18273 ( .A(n19805), .B(n17909), .Z(n17833) );
  AND U18274 ( .A(n17834), .B(n17833), .Z(n17916) );
  NAND U18275 ( .A(n35), .B(n17835), .Z(n17837) );
  XOR U18276 ( .A(b[9]), .B(a[231]), .Z(n17912) );
  NAND U18277 ( .A(n19598), .B(n17912), .Z(n17836) );
  NAND U18278 ( .A(n17837), .B(n17836), .Z(n17915) );
  XOR U18279 ( .A(n17916), .B(n17915), .Z(n17918) );
  XOR U18280 ( .A(n17917), .B(n17918), .Z(n17928) );
  NANDN U18281 ( .A(n17839), .B(n17838), .Z(n17843) );
  OR U18282 ( .A(n17841), .B(n17840), .Z(n17842) );
  AND U18283 ( .A(n17843), .B(n17842), .Z(n17927) );
  XNOR U18284 ( .A(n17928), .B(n17927), .Z(n17929) );
  NANDN U18285 ( .A(n17845), .B(n17844), .Z(n17849) );
  NANDN U18286 ( .A(n17847), .B(n17846), .Z(n17848) );
  NAND U18287 ( .A(n17849), .B(n17848), .Z(n17930) );
  XNOR U18288 ( .A(n17929), .B(n17930), .Z(n17875) );
  XOR U18289 ( .A(n17876), .B(n17875), .Z(n17934) );
  NANDN U18290 ( .A(n17851), .B(n17850), .Z(n17855) );
  NANDN U18291 ( .A(n17853), .B(n17852), .Z(n17854) );
  AND U18292 ( .A(n17855), .B(n17854), .Z(n17933) );
  XNOR U18293 ( .A(n17934), .B(n17933), .Z(n17935) );
  XOR U18294 ( .A(n17936), .B(n17935), .Z(n17868) );
  NANDN U18295 ( .A(n17857), .B(n17856), .Z(n17861) );
  NAND U18296 ( .A(n17859), .B(n17858), .Z(n17860) );
  AND U18297 ( .A(n17861), .B(n17860), .Z(n17867) );
  XNOR U18298 ( .A(n17868), .B(n17867), .Z(n17869) );
  XNOR U18299 ( .A(n17870), .B(n17869), .Z(n17939) );
  XNOR U18300 ( .A(sreg[479]), .B(n17939), .Z(n17941) );
  NANDN U18301 ( .A(sreg[478]), .B(n17862), .Z(n17866) );
  NAND U18302 ( .A(n17864), .B(n17863), .Z(n17865) );
  NAND U18303 ( .A(n17866), .B(n17865), .Z(n17940) );
  XNOR U18304 ( .A(n17941), .B(n17940), .Z(c[479]) );
  NANDN U18305 ( .A(n17868), .B(n17867), .Z(n17872) );
  NANDN U18306 ( .A(n17870), .B(n17869), .Z(n17871) );
  AND U18307 ( .A(n17872), .B(n17871), .Z(n17947) );
  NANDN U18308 ( .A(n17874), .B(n17873), .Z(n17878) );
  NAND U18309 ( .A(n17876), .B(n17875), .Z(n17877) );
  AND U18310 ( .A(n17878), .B(n17877), .Z(n18013) );
  NANDN U18311 ( .A(n17880), .B(n17879), .Z(n17884) );
  NANDN U18312 ( .A(n17882), .B(n17881), .Z(n17883) );
  AND U18313 ( .A(n17884), .B(n17883), .Z(n17979) );
  NAND U18314 ( .A(n19808), .B(n17885), .Z(n17887) );
  XOR U18315 ( .A(b[13]), .B(a[228]), .Z(n17965) );
  NAND U18316 ( .A(n19768), .B(n17965), .Z(n17886) );
  AND U18317 ( .A(n17887), .B(n17886), .Z(n17957) );
  AND U18318 ( .A(b[15]), .B(a[224]), .Z(n17956) );
  XNOR U18319 ( .A(n17957), .B(n17956), .Z(n17958) );
  NAND U18320 ( .A(b[0]), .B(a[240]), .Z(n17888) );
  XNOR U18321 ( .A(b[1]), .B(n17888), .Z(n17890) );
  NANDN U18322 ( .A(b[0]), .B(a[239]), .Z(n17889) );
  NAND U18323 ( .A(n17890), .B(n17889), .Z(n17959) );
  XNOR U18324 ( .A(n17958), .B(n17959), .Z(n17977) );
  NAND U18325 ( .A(n33), .B(n17891), .Z(n17893) );
  XOR U18326 ( .A(b[5]), .B(a[236]), .Z(n17968) );
  NAND U18327 ( .A(n19342), .B(n17968), .Z(n17892) );
  AND U18328 ( .A(n17893), .B(n17892), .Z(n18001) );
  NAND U18329 ( .A(n34), .B(n17894), .Z(n17896) );
  XOR U18330 ( .A(b[7]), .B(a[234]), .Z(n17971) );
  NAND U18331 ( .A(n19486), .B(n17971), .Z(n17895) );
  AND U18332 ( .A(n17896), .B(n17895), .Z(n17999) );
  NAND U18333 ( .A(n31), .B(n17897), .Z(n17899) );
  XOR U18334 ( .A(b[3]), .B(a[238]), .Z(n17974) );
  NAND U18335 ( .A(n32), .B(n17974), .Z(n17898) );
  NAND U18336 ( .A(n17899), .B(n17898), .Z(n17998) );
  XNOR U18337 ( .A(n17999), .B(n17998), .Z(n18000) );
  XOR U18338 ( .A(n18001), .B(n18000), .Z(n17978) );
  XOR U18339 ( .A(n17977), .B(n17978), .Z(n17980) );
  XOR U18340 ( .A(n17979), .B(n17980), .Z(n17951) );
  NANDN U18341 ( .A(n17901), .B(n17900), .Z(n17905) );
  OR U18342 ( .A(n17903), .B(n17902), .Z(n17904) );
  AND U18343 ( .A(n17905), .B(n17904), .Z(n17950) );
  XNOR U18344 ( .A(n17951), .B(n17950), .Z(n17953) );
  NAND U18345 ( .A(n17906), .B(n19724), .Z(n17908) );
  XOR U18346 ( .A(b[11]), .B(a[230]), .Z(n17983) );
  NAND U18347 ( .A(n19692), .B(n17983), .Z(n17907) );
  AND U18348 ( .A(n17908), .B(n17907), .Z(n17994) );
  NAND U18349 ( .A(n19838), .B(n17909), .Z(n17911) );
  XOR U18350 ( .A(b[15]), .B(a[226]), .Z(n17986) );
  NAND U18351 ( .A(n19805), .B(n17986), .Z(n17910) );
  AND U18352 ( .A(n17911), .B(n17910), .Z(n17993) );
  NAND U18353 ( .A(n35), .B(n17912), .Z(n17914) );
  XOR U18354 ( .A(b[9]), .B(a[232]), .Z(n17989) );
  NAND U18355 ( .A(n19598), .B(n17989), .Z(n17913) );
  NAND U18356 ( .A(n17914), .B(n17913), .Z(n17992) );
  XOR U18357 ( .A(n17993), .B(n17992), .Z(n17995) );
  XOR U18358 ( .A(n17994), .B(n17995), .Z(n18005) );
  NANDN U18359 ( .A(n17916), .B(n17915), .Z(n17920) );
  OR U18360 ( .A(n17918), .B(n17917), .Z(n17919) );
  AND U18361 ( .A(n17920), .B(n17919), .Z(n18004) );
  XNOR U18362 ( .A(n18005), .B(n18004), .Z(n18006) );
  NANDN U18363 ( .A(n17922), .B(n17921), .Z(n17926) );
  NANDN U18364 ( .A(n17924), .B(n17923), .Z(n17925) );
  NAND U18365 ( .A(n17926), .B(n17925), .Z(n18007) );
  XNOR U18366 ( .A(n18006), .B(n18007), .Z(n17952) );
  XOR U18367 ( .A(n17953), .B(n17952), .Z(n18011) );
  NANDN U18368 ( .A(n17928), .B(n17927), .Z(n17932) );
  NANDN U18369 ( .A(n17930), .B(n17929), .Z(n17931) );
  AND U18370 ( .A(n17932), .B(n17931), .Z(n18010) );
  XNOR U18371 ( .A(n18011), .B(n18010), .Z(n18012) );
  XOR U18372 ( .A(n18013), .B(n18012), .Z(n17945) );
  NANDN U18373 ( .A(n17934), .B(n17933), .Z(n17938) );
  NAND U18374 ( .A(n17936), .B(n17935), .Z(n17937) );
  AND U18375 ( .A(n17938), .B(n17937), .Z(n17944) );
  XNOR U18376 ( .A(n17945), .B(n17944), .Z(n17946) );
  XNOR U18377 ( .A(n17947), .B(n17946), .Z(n18016) );
  XNOR U18378 ( .A(sreg[480]), .B(n18016), .Z(n18018) );
  NANDN U18379 ( .A(sreg[479]), .B(n17939), .Z(n17943) );
  NAND U18380 ( .A(n17941), .B(n17940), .Z(n17942) );
  NAND U18381 ( .A(n17943), .B(n17942), .Z(n18017) );
  XNOR U18382 ( .A(n18018), .B(n18017), .Z(c[480]) );
  NANDN U18383 ( .A(n17945), .B(n17944), .Z(n17949) );
  NANDN U18384 ( .A(n17947), .B(n17946), .Z(n17948) );
  AND U18385 ( .A(n17949), .B(n17948), .Z(n18024) );
  NANDN U18386 ( .A(n17951), .B(n17950), .Z(n17955) );
  NAND U18387 ( .A(n17953), .B(n17952), .Z(n17954) );
  AND U18388 ( .A(n17955), .B(n17954), .Z(n18090) );
  NANDN U18389 ( .A(n17957), .B(n17956), .Z(n17961) );
  NANDN U18390 ( .A(n17959), .B(n17958), .Z(n17960) );
  AND U18391 ( .A(n17961), .B(n17960), .Z(n18077) );
  NAND U18392 ( .A(b[0]), .B(a[241]), .Z(n17962) );
  XNOR U18393 ( .A(b[1]), .B(n17962), .Z(n17964) );
  NANDN U18394 ( .A(b[0]), .B(a[240]), .Z(n17963) );
  NAND U18395 ( .A(n17964), .B(n17963), .Z(n18057) );
  NAND U18396 ( .A(n19808), .B(n17965), .Z(n17967) );
  XOR U18397 ( .A(b[13]), .B(a[229]), .Z(n18060) );
  NAND U18398 ( .A(n19768), .B(n18060), .Z(n17966) );
  AND U18399 ( .A(n17967), .B(n17966), .Z(n18055) );
  AND U18400 ( .A(b[15]), .B(a[225]), .Z(n18054) );
  XNOR U18401 ( .A(n18055), .B(n18054), .Z(n18056) );
  XNOR U18402 ( .A(n18057), .B(n18056), .Z(n18075) );
  NAND U18403 ( .A(n33), .B(n17968), .Z(n17970) );
  XOR U18404 ( .A(b[5]), .B(a[237]), .Z(n18066) );
  NAND U18405 ( .A(n19342), .B(n18066), .Z(n17969) );
  AND U18406 ( .A(n17970), .B(n17969), .Z(n18051) );
  NAND U18407 ( .A(n34), .B(n17971), .Z(n17973) );
  XOR U18408 ( .A(b[7]), .B(a[235]), .Z(n18069) );
  NAND U18409 ( .A(n19486), .B(n18069), .Z(n17972) );
  AND U18410 ( .A(n17973), .B(n17972), .Z(n18049) );
  NAND U18411 ( .A(n31), .B(n17974), .Z(n17976) );
  XOR U18412 ( .A(b[3]), .B(a[239]), .Z(n18072) );
  NAND U18413 ( .A(n32), .B(n18072), .Z(n17975) );
  NAND U18414 ( .A(n17976), .B(n17975), .Z(n18048) );
  XNOR U18415 ( .A(n18049), .B(n18048), .Z(n18050) );
  XOR U18416 ( .A(n18051), .B(n18050), .Z(n18076) );
  XOR U18417 ( .A(n18075), .B(n18076), .Z(n18078) );
  XOR U18418 ( .A(n18077), .B(n18078), .Z(n18028) );
  NANDN U18419 ( .A(n17978), .B(n17977), .Z(n17982) );
  OR U18420 ( .A(n17980), .B(n17979), .Z(n17981) );
  AND U18421 ( .A(n17982), .B(n17981), .Z(n18027) );
  XNOR U18422 ( .A(n18028), .B(n18027), .Z(n18030) );
  NAND U18423 ( .A(n17983), .B(n19724), .Z(n17985) );
  XOR U18424 ( .A(b[11]), .B(a[231]), .Z(n18033) );
  NAND U18425 ( .A(n19692), .B(n18033), .Z(n17984) );
  AND U18426 ( .A(n17985), .B(n17984), .Z(n18044) );
  NAND U18427 ( .A(n19838), .B(n17986), .Z(n17988) );
  XOR U18428 ( .A(b[15]), .B(a[227]), .Z(n18036) );
  NAND U18429 ( .A(n19805), .B(n18036), .Z(n17987) );
  AND U18430 ( .A(n17988), .B(n17987), .Z(n18043) );
  NAND U18431 ( .A(n35), .B(n17989), .Z(n17991) );
  XOR U18432 ( .A(b[9]), .B(a[233]), .Z(n18039) );
  NAND U18433 ( .A(n19598), .B(n18039), .Z(n17990) );
  NAND U18434 ( .A(n17991), .B(n17990), .Z(n18042) );
  XOR U18435 ( .A(n18043), .B(n18042), .Z(n18045) );
  XOR U18436 ( .A(n18044), .B(n18045), .Z(n18082) );
  NANDN U18437 ( .A(n17993), .B(n17992), .Z(n17997) );
  OR U18438 ( .A(n17995), .B(n17994), .Z(n17996) );
  AND U18439 ( .A(n17997), .B(n17996), .Z(n18081) );
  XNOR U18440 ( .A(n18082), .B(n18081), .Z(n18083) );
  NANDN U18441 ( .A(n17999), .B(n17998), .Z(n18003) );
  NANDN U18442 ( .A(n18001), .B(n18000), .Z(n18002) );
  NAND U18443 ( .A(n18003), .B(n18002), .Z(n18084) );
  XNOR U18444 ( .A(n18083), .B(n18084), .Z(n18029) );
  XOR U18445 ( .A(n18030), .B(n18029), .Z(n18088) );
  NANDN U18446 ( .A(n18005), .B(n18004), .Z(n18009) );
  NANDN U18447 ( .A(n18007), .B(n18006), .Z(n18008) );
  AND U18448 ( .A(n18009), .B(n18008), .Z(n18087) );
  XNOR U18449 ( .A(n18088), .B(n18087), .Z(n18089) );
  XOR U18450 ( .A(n18090), .B(n18089), .Z(n18022) );
  NANDN U18451 ( .A(n18011), .B(n18010), .Z(n18015) );
  NAND U18452 ( .A(n18013), .B(n18012), .Z(n18014) );
  AND U18453 ( .A(n18015), .B(n18014), .Z(n18021) );
  XNOR U18454 ( .A(n18022), .B(n18021), .Z(n18023) );
  XNOR U18455 ( .A(n18024), .B(n18023), .Z(n18093) );
  XNOR U18456 ( .A(sreg[481]), .B(n18093), .Z(n18095) );
  NANDN U18457 ( .A(sreg[480]), .B(n18016), .Z(n18020) );
  NAND U18458 ( .A(n18018), .B(n18017), .Z(n18019) );
  NAND U18459 ( .A(n18020), .B(n18019), .Z(n18094) );
  XNOR U18460 ( .A(n18095), .B(n18094), .Z(c[481]) );
  NANDN U18461 ( .A(n18022), .B(n18021), .Z(n18026) );
  NANDN U18462 ( .A(n18024), .B(n18023), .Z(n18025) );
  AND U18463 ( .A(n18026), .B(n18025), .Z(n18101) );
  NANDN U18464 ( .A(n18028), .B(n18027), .Z(n18032) );
  NAND U18465 ( .A(n18030), .B(n18029), .Z(n18031) );
  AND U18466 ( .A(n18032), .B(n18031), .Z(n18167) );
  NAND U18467 ( .A(n18033), .B(n19724), .Z(n18035) );
  XOR U18468 ( .A(b[11]), .B(a[232]), .Z(n18137) );
  NAND U18469 ( .A(n19692), .B(n18137), .Z(n18034) );
  AND U18470 ( .A(n18035), .B(n18034), .Z(n18148) );
  NAND U18471 ( .A(n19838), .B(n18036), .Z(n18038) );
  XOR U18472 ( .A(b[15]), .B(a[228]), .Z(n18140) );
  NAND U18473 ( .A(n19805), .B(n18140), .Z(n18037) );
  AND U18474 ( .A(n18038), .B(n18037), .Z(n18147) );
  NAND U18475 ( .A(n35), .B(n18039), .Z(n18041) );
  XOR U18476 ( .A(b[9]), .B(a[234]), .Z(n18143) );
  NAND U18477 ( .A(n19598), .B(n18143), .Z(n18040) );
  NAND U18478 ( .A(n18041), .B(n18040), .Z(n18146) );
  XOR U18479 ( .A(n18147), .B(n18146), .Z(n18149) );
  XOR U18480 ( .A(n18148), .B(n18149), .Z(n18159) );
  NANDN U18481 ( .A(n18043), .B(n18042), .Z(n18047) );
  OR U18482 ( .A(n18045), .B(n18044), .Z(n18046) );
  AND U18483 ( .A(n18047), .B(n18046), .Z(n18158) );
  XNOR U18484 ( .A(n18159), .B(n18158), .Z(n18160) );
  NANDN U18485 ( .A(n18049), .B(n18048), .Z(n18053) );
  NANDN U18486 ( .A(n18051), .B(n18050), .Z(n18052) );
  NAND U18487 ( .A(n18053), .B(n18052), .Z(n18161) );
  XNOR U18488 ( .A(n18160), .B(n18161), .Z(n18107) );
  NANDN U18489 ( .A(n18055), .B(n18054), .Z(n18059) );
  NANDN U18490 ( .A(n18057), .B(n18056), .Z(n18058) );
  AND U18491 ( .A(n18059), .B(n18058), .Z(n18133) );
  NAND U18492 ( .A(n19808), .B(n18060), .Z(n18062) );
  XOR U18493 ( .A(b[13]), .B(a[230]), .Z(n18119) );
  NAND U18494 ( .A(n19768), .B(n18119), .Z(n18061) );
  AND U18495 ( .A(n18062), .B(n18061), .Z(n18111) );
  AND U18496 ( .A(b[15]), .B(a[226]), .Z(n18110) );
  XNOR U18497 ( .A(n18111), .B(n18110), .Z(n18112) );
  NAND U18498 ( .A(b[0]), .B(a[242]), .Z(n18063) );
  XNOR U18499 ( .A(b[1]), .B(n18063), .Z(n18065) );
  NANDN U18500 ( .A(b[0]), .B(a[241]), .Z(n18064) );
  NAND U18501 ( .A(n18065), .B(n18064), .Z(n18113) );
  XNOR U18502 ( .A(n18112), .B(n18113), .Z(n18131) );
  NAND U18503 ( .A(n33), .B(n18066), .Z(n18068) );
  XOR U18504 ( .A(b[5]), .B(a[238]), .Z(n18122) );
  NAND U18505 ( .A(n19342), .B(n18122), .Z(n18067) );
  AND U18506 ( .A(n18068), .B(n18067), .Z(n18155) );
  NAND U18507 ( .A(n34), .B(n18069), .Z(n18071) );
  XOR U18508 ( .A(b[7]), .B(a[236]), .Z(n18125) );
  NAND U18509 ( .A(n19486), .B(n18125), .Z(n18070) );
  AND U18510 ( .A(n18071), .B(n18070), .Z(n18153) );
  NAND U18511 ( .A(n31), .B(n18072), .Z(n18074) );
  XOR U18512 ( .A(b[3]), .B(a[240]), .Z(n18128) );
  NAND U18513 ( .A(n32), .B(n18128), .Z(n18073) );
  NAND U18514 ( .A(n18074), .B(n18073), .Z(n18152) );
  XNOR U18515 ( .A(n18153), .B(n18152), .Z(n18154) );
  XOR U18516 ( .A(n18155), .B(n18154), .Z(n18132) );
  XOR U18517 ( .A(n18131), .B(n18132), .Z(n18134) );
  XOR U18518 ( .A(n18133), .B(n18134), .Z(n18105) );
  NANDN U18519 ( .A(n18076), .B(n18075), .Z(n18080) );
  OR U18520 ( .A(n18078), .B(n18077), .Z(n18079) );
  AND U18521 ( .A(n18080), .B(n18079), .Z(n18104) );
  XNOR U18522 ( .A(n18105), .B(n18104), .Z(n18106) );
  XOR U18523 ( .A(n18107), .B(n18106), .Z(n18165) );
  NANDN U18524 ( .A(n18082), .B(n18081), .Z(n18086) );
  NANDN U18525 ( .A(n18084), .B(n18083), .Z(n18085) );
  AND U18526 ( .A(n18086), .B(n18085), .Z(n18164) );
  XNOR U18527 ( .A(n18165), .B(n18164), .Z(n18166) );
  XOR U18528 ( .A(n18167), .B(n18166), .Z(n18099) );
  NANDN U18529 ( .A(n18088), .B(n18087), .Z(n18092) );
  NAND U18530 ( .A(n18090), .B(n18089), .Z(n18091) );
  AND U18531 ( .A(n18092), .B(n18091), .Z(n18098) );
  XNOR U18532 ( .A(n18099), .B(n18098), .Z(n18100) );
  XNOR U18533 ( .A(n18101), .B(n18100), .Z(n18170) );
  XNOR U18534 ( .A(sreg[482]), .B(n18170), .Z(n18172) );
  NANDN U18535 ( .A(sreg[481]), .B(n18093), .Z(n18097) );
  NAND U18536 ( .A(n18095), .B(n18094), .Z(n18096) );
  NAND U18537 ( .A(n18097), .B(n18096), .Z(n18171) );
  XNOR U18538 ( .A(n18172), .B(n18171), .Z(c[482]) );
  NANDN U18539 ( .A(n18099), .B(n18098), .Z(n18103) );
  NANDN U18540 ( .A(n18101), .B(n18100), .Z(n18102) );
  AND U18541 ( .A(n18103), .B(n18102), .Z(n18178) );
  NANDN U18542 ( .A(n18105), .B(n18104), .Z(n18109) );
  NAND U18543 ( .A(n18107), .B(n18106), .Z(n18108) );
  AND U18544 ( .A(n18109), .B(n18108), .Z(n18244) );
  NANDN U18545 ( .A(n18111), .B(n18110), .Z(n18115) );
  NANDN U18546 ( .A(n18113), .B(n18112), .Z(n18114) );
  AND U18547 ( .A(n18115), .B(n18114), .Z(n18210) );
  NAND U18548 ( .A(b[0]), .B(a[243]), .Z(n18116) );
  XNOR U18549 ( .A(b[1]), .B(n18116), .Z(n18118) );
  NANDN U18550 ( .A(b[0]), .B(a[242]), .Z(n18117) );
  NAND U18551 ( .A(n18118), .B(n18117), .Z(n18190) );
  NAND U18552 ( .A(n19808), .B(n18119), .Z(n18121) );
  XOR U18553 ( .A(b[13]), .B(a[231]), .Z(n18196) );
  NAND U18554 ( .A(n19768), .B(n18196), .Z(n18120) );
  AND U18555 ( .A(n18121), .B(n18120), .Z(n18188) );
  AND U18556 ( .A(b[15]), .B(a[227]), .Z(n18187) );
  XNOR U18557 ( .A(n18188), .B(n18187), .Z(n18189) );
  XNOR U18558 ( .A(n18190), .B(n18189), .Z(n18208) );
  NAND U18559 ( .A(n33), .B(n18122), .Z(n18124) );
  XOR U18560 ( .A(b[5]), .B(a[239]), .Z(n18199) );
  NAND U18561 ( .A(n19342), .B(n18199), .Z(n18123) );
  AND U18562 ( .A(n18124), .B(n18123), .Z(n18232) );
  NAND U18563 ( .A(n34), .B(n18125), .Z(n18127) );
  XOR U18564 ( .A(b[7]), .B(a[237]), .Z(n18202) );
  NAND U18565 ( .A(n19486), .B(n18202), .Z(n18126) );
  AND U18566 ( .A(n18127), .B(n18126), .Z(n18230) );
  NAND U18567 ( .A(n31), .B(n18128), .Z(n18130) );
  XOR U18568 ( .A(b[3]), .B(a[241]), .Z(n18205) );
  NAND U18569 ( .A(n32), .B(n18205), .Z(n18129) );
  NAND U18570 ( .A(n18130), .B(n18129), .Z(n18229) );
  XNOR U18571 ( .A(n18230), .B(n18229), .Z(n18231) );
  XOR U18572 ( .A(n18232), .B(n18231), .Z(n18209) );
  XOR U18573 ( .A(n18208), .B(n18209), .Z(n18211) );
  XOR U18574 ( .A(n18210), .B(n18211), .Z(n18182) );
  NANDN U18575 ( .A(n18132), .B(n18131), .Z(n18136) );
  OR U18576 ( .A(n18134), .B(n18133), .Z(n18135) );
  AND U18577 ( .A(n18136), .B(n18135), .Z(n18181) );
  XNOR U18578 ( .A(n18182), .B(n18181), .Z(n18184) );
  NAND U18579 ( .A(n18137), .B(n19724), .Z(n18139) );
  XOR U18580 ( .A(b[11]), .B(a[233]), .Z(n18214) );
  NAND U18581 ( .A(n19692), .B(n18214), .Z(n18138) );
  AND U18582 ( .A(n18139), .B(n18138), .Z(n18225) );
  NAND U18583 ( .A(n19838), .B(n18140), .Z(n18142) );
  XOR U18584 ( .A(b[15]), .B(a[229]), .Z(n18217) );
  NAND U18585 ( .A(n19805), .B(n18217), .Z(n18141) );
  AND U18586 ( .A(n18142), .B(n18141), .Z(n18224) );
  NAND U18587 ( .A(n35), .B(n18143), .Z(n18145) );
  XOR U18588 ( .A(b[9]), .B(a[235]), .Z(n18220) );
  NAND U18589 ( .A(n19598), .B(n18220), .Z(n18144) );
  NAND U18590 ( .A(n18145), .B(n18144), .Z(n18223) );
  XOR U18591 ( .A(n18224), .B(n18223), .Z(n18226) );
  XOR U18592 ( .A(n18225), .B(n18226), .Z(n18236) );
  NANDN U18593 ( .A(n18147), .B(n18146), .Z(n18151) );
  OR U18594 ( .A(n18149), .B(n18148), .Z(n18150) );
  AND U18595 ( .A(n18151), .B(n18150), .Z(n18235) );
  XNOR U18596 ( .A(n18236), .B(n18235), .Z(n18237) );
  NANDN U18597 ( .A(n18153), .B(n18152), .Z(n18157) );
  NANDN U18598 ( .A(n18155), .B(n18154), .Z(n18156) );
  NAND U18599 ( .A(n18157), .B(n18156), .Z(n18238) );
  XNOR U18600 ( .A(n18237), .B(n18238), .Z(n18183) );
  XOR U18601 ( .A(n18184), .B(n18183), .Z(n18242) );
  NANDN U18602 ( .A(n18159), .B(n18158), .Z(n18163) );
  NANDN U18603 ( .A(n18161), .B(n18160), .Z(n18162) );
  AND U18604 ( .A(n18163), .B(n18162), .Z(n18241) );
  XNOR U18605 ( .A(n18242), .B(n18241), .Z(n18243) );
  XOR U18606 ( .A(n18244), .B(n18243), .Z(n18176) );
  NANDN U18607 ( .A(n18165), .B(n18164), .Z(n18169) );
  NAND U18608 ( .A(n18167), .B(n18166), .Z(n18168) );
  AND U18609 ( .A(n18169), .B(n18168), .Z(n18175) );
  XNOR U18610 ( .A(n18176), .B(n18175), .Z(n18177) );
  XNOR U18611 ( .A(n18178), .B(n18177), .Z(n18247) );
  XNOR U18612 ( .A(sreg[483]), .B(n18247), .Z(n18249) );
  NANDN U18613 ( .A(sreg[482]), .B(n18170), .Z(n18174) );
  NAND U18614 ( .A(n18172), .B(n18171), .Z(n18173) );
  NAND U18615 ( .A(n18174), .B(n18173), .Z(n18248) );
  XNOR U18616 ( .A(n18249), .B(n18248), .Z(c[483]) );
  NANDN U18617 ( .A(n18176), .B(n18175), .Z(n18180) );
  NANDN U18618 ( .A(n18178), .B(n18177), .Z(n18179) );
  AND U18619 ( .A(n18180), .B(n18179), .Z(n18255) );
  NANDN U18620 ( .A(n18182), .B(n18181), .Z(n18186) );
  NAND U18621 ( .A(n18184), .B(n18183), .Z(n18185) );
  AND U18622 ( .A(n18186), .B(n18185), .Z(n18321) );
  NANDN U18623 ( .A(n18188), .B(n18187), .Z(n18192) );
  NANDN U18624 ( .A(n18190), .B(n18189), .Z(n18191) );
  AND U18625 ( .A(n18192), .B(n18191), .Z(n18287) );
  NAND U18626 ( .A(b[0]), .B(a[244]), .Z(n18193) );
  XNOR U18627 ( .A(b[1]), .B(n18193), .Z(n18195) );
  NANDN U18628 ( .A(b[0]), .B(a[243]), .Z(n18194) );
  NAND U18629 ( .A(n18195), .B(n18194), .Z(n18267) );
  NAND U18630 ( .A(n19808), .B(n18196), .Z(n18198) );
  XOR U18631 ( .A(b[13]), .B(a[232]), .Z(n18270) );
  NAND U18632 ( .A(n19768), .B(n18270), .Z(n18197) );
  AND U18633 ( .A(n18198), .B(n18197), .Z(n18265) );
  AND U18634 ( .A(b[15]), .B(a[228]), .Z(n18264) );
  XNOR U18635 ( .A(n18265), .B(n18264), .Z(n18266) );
  XNOR U18636 ( .A(n18267), .B(n18266), .Z(n18285) );
  NAND U18637 ( .A(n33), .B(n18199), .Z(n18201) );
  XOR U18638 ( .A(b[5]), .B(a[240]), .Z(n18276) );
  NAND U18639 ( .A(n19342), .B(n18276), .Z(n18200) );
  AND U18640 ( .A(n18201), .B(n18200), .Z(n18309) );
  NAND U18641 ( .A(n34), .B(n18202), .Z(n18204) );
  XOR U18642 ( .A(b[7]), .B(a[238]), .Z(n18279) );
  NAND U18643 ( .A(n19486), .B(n18279), .Z(n18203) );
  AND U18644 ( .A(n18204), .B(n18203), .Z(n18307) );
  NAND U18645 ( .A(n31), .B(n18205), .Z(n18207) );
  XOR U18646 ( .A(b[3]), .B(a[242]), .Z(n18282) );
  NAND U18647 ( .A(n32), .B(n18282), .Z(n18206) );
  NAND U18648 ( .A(n18207), .B(n18206), .Z(n18306) );
  XNOR U18649 ( .A(n18307), .B(n18306), .Z(n18308) );
  XOR U18650 ( .A(n18309), .B(n18308), .Z(n18286) );
  XOR U18651 ( .A(n18285), .B(n18286), .Z(n18288) );
  XOR U18652 ( .A(n18287), .B(n18288), .Z(n18259) );
  NANDN U18653 ( .A(n18209), .B(n18208), .Z(n18213) );
  OR U18654 ( .A(n18211), .B(n18210), .Z(n18212) );
  AND U18655 ( .A(n18213), .B(n18212), .Z(n18258) );
  XNOR U18656 ( .A(n18259), .B(n18258), .Z(n18261) );
  NAND U18657 ( .A(n18214), .B(n19724), .Z(n18216) );
  XOR U18658 ( .A(b[11]), .B(a[234]), .Z(n18291) );
  NAND U18659 ( .A(n19692), .B(n18291), .Z(n18215) );
  AND U18660 ( .A(n18216), .B(n18215), .Z(n18302) );
  NAND U18661 ( .A(n19838), .B(n18217), .Z(n18219) );
  XOR U18662 ( .A(b[15]), .B(a[230]), .Z(n18294) );
  NAND U18663 ( .A(n19805), .B(n18294), .Z(n18218) );
  AND U18664 ( .A(n18219), .B(n18218), .Z(n18301) );
  NAND U18665 ( .A(n35), .B(n18220), .Z(n18222) );
  XOR U18666 ( .A(b[9]), .B(a[236]), .Z(n18297) );
  NAND U18667 ( .A(n19598), .B(n18297), .Z(n18221) );
  NAND U18668 ( .A(n18222), .B(n18221), .Z(n18300) );
  XOR U18669 ( .A(n18301), .B(n18300), .Z(n18303) );
  XOR U18670 ( .A(n18302), .B(n18303), .Z(n18313) );
  NANDN U18671 ( .A(n18224), .B(n18223), .Z(n18228) );
  OR U18672 ( .A(n18226), .B(n18225), .Z(n18227) );
  AND U18673 ( .A(n18228), .B(n18227), .Z(n18312) );
  XNOR U18674 ( .A(n18313), .B(n18312), .Z(n18314) );
  NANDN U18675 ( .A(n18230), .B(n18229), .Z(n18234) );
  NANDN U18676 ( .A(n18232), .B(n18231), .Z(n18233) );
  NAND U18677 ( .A(n18234), .B(n18233), .Z(n18315) );
  XNOR U18678 ( .A(n18314), .B(n18315), .Z(n18260) );
  XOR U18679 ( .A(n18261), .B(n18260), .Z(n18319) );
  NANDN U18680 ( .A(n18236), .B(n18235), .Z(n18240) );
  NANDN U18681 ( .A(n18238), .B(n18237), .Z(n18239) );
  AND U18682 ( .A(n18240), .B(n18239), .Z(n18318) );
  XNOR U18683 ( .A(n18319), .B(n18318), .Z(n18320) );
  XOR U18684 ( .A(n18321), .B(n18320), .Z(n18253) );
  NANDN U18685 ( .A(n18242), .B(n18241), .Z(n18246) );
  NAND U18686 ( .A(n18244), .B(n18243), .Z(n18245) );
  AND U18687 ( .A(n18246), .B(n18245), .Z(n18252) );
  XNOR U18688 ( .A(n18253), .B(n18252), .Z(n18254) );
  XNOR U18689 ( .A(n18255), .B(n18254), .Z(n18324) );
  XNOR U18690 ( .A(sreg[484]), .B(n18324), .Z(n18326) );
  NANDN U18691 ( .A(sreg[483]), .B(n18247), .Z(n18251) );
  NAND U18692 ( .A(n18249), .B(n18248), .Z(n18250) );
  NAND U18693 ( .A(n18251), .B(n18250), .Z(n18325) );
  XNOR U18694 ( .A(n18326), .B(n18325), .Z(c[484]) );
  NANDN U18695 ( .A(n18253), .B(n18252), .Z(n18257) );
  NANDN U18696 ( .A(n18255), .B(n18254), .Z(n18256) );
  AND U18697 ( .A(n18257), .B(n18256), .Z(n18332) );
  NANDN U18698 ( .A(n18259), .B(n18258), .Z(n18263) );
  NAND U18699 ( .A(n18261), .B(n18260), .Z(n18262) );
  AND U18700 ( .A(n18263), .B(n18262), .Z(n18398) );
  NANDN U18701 ( .A(n18265), .B(n18264), .Z(n18269) );
  NANDN U18702 ( .A(n18267), .B(n18266), .Z(n18268) );
  AND U18703 ( .A(n18269), .B(n18268), .Z(n18364) );
  NAND U18704 ( .A(n19808), .B(n18270), .Z(n18272) );
  XOR U18705 ( .A(b[13]), .B(a[233]), .Z(n18350) );
  NAND U18706 ( .A(n19768), .B(n18350), .Z(n18271) );
  AND U18707 ( .A(n18272), .B(n18271), .Z(n18342) );
  AND U18708 ( .A(b[15]), .B(a[229]), .Z(n18341) );
  XNOR U18709 ( .A(n18342), .B(n18341), .Z(n18343) );
  NAND U18710 ( .A(b[0]), .B(a[245]), .Z(n18273) );
  XNOR U18711 ( .A(b[1]), .B(n18273), .Z(n18275) );
  NANDN U18712 ( .A(b[0]), .B(a[244]), .Z(n18274) );
  NAND U18713 ( .A(n18275), .B(n18274), .Z(n18344) );
  XNOR U18714 ( .A(n18343), .B(n18344), .Z(n18362) );
  NAND U18715 ( .A(n33), .B(n18276), .Z(n18278) );
  XOR U18716 ( .A(b[5]), .B(a[241]), .Z(n18353) );
  NAND U18717 ( .A(n19342), .B(n18353), .Z(n18277) );
  AND U18718 ( .A(n18278), .B(n18277), .Z(n18386) );
  NAND U18719 ( .A(n34), .B(n18279), .Z(n18281) );
  XOR U18720 ( .A(b[7]), .B(a[239]), .Z(n18356) );
  NAND U18721 ( .A(n19486), .B(n18356), .Z(n18280) );
  AND U18722 ( .A(n18281), .B(n18280), .Z(n18384) );
  NAND U18723 ( .A(n31), .B(n18282), .Z(n18284) );
  XOR U18724 ( .A(b[3]), .B(a[243]), .Z(n18359) );
  NAND U18725 ( .A(n32), .B(n18359), .Z(n18283) );
  NAND U18726 ( .A(n18284), .B(n18283), .Z(n18383) );
  XNOR U18727 ( .A(n18384), .B(n18383), .Z(n18385) );
  XOR U18728 ( .A(n18386), .B(n18385), .Z(n18363) );
  XOR U18729 ( .A(n18362), .B(n18363), .Z(n18365) );
  XOR U18730 ( .A(n18364), .B(n18365), .Z(n18336) );
  NANDN U18731 ( .A(n18286), .B(n18285), .Z(n18290) );
  OR U18732 ( .A(n18288), .B(n18287), .Z(n18289) );
  AND U18733 ( .A(n18290), .B(n18289), .Z(n18335) );
  XNOR U18734 ( .A(n18336), .B(n18335), .Z(n18338) );
  NAND U18735 ( .A(n18291), .B(n19724), .Z(n18293) );
  XOR U18736 ( .A(b[11]), .B(a[235]), .Z(n18368) );
  NAND U18737 ( .A(n19692), .B(n18368), .Z(n18292) );
  AND U18738 ( .A(n18293), .B(n18292), .Z(n18379) );
  NAND U18739 ( .A(n19838), .B(n18294), .Z(n18296) );
  XOR U18740 ( .A(b[15]), .B(a[231]), .Z(n18371) );
  NAND U18741 ( .A(n19805), .B(n18371), .Z(n18295) );
  AND U18742 ( .A(n18296), .B(n18295), .Z(n18378) );
  NAND U18743 ( .A(n35), .B(n18297), .Z(n18299) );
  XOR U18744 ( .A(b[9]), .B(a[237]), .Z(n18374) );
  NAND U18745 ( .A(n19598), .B(n18374), .Z(n18298) );
  NAND U18746 ( .A(n18299), .B(n18298), .Z(n18377) );
  XOR U18747 ( .A(n18378), .B(n18377), .Z(n18380) );
  XOR U18748 ( .A(n18379), .B(n18380), .Z(n18390) );
  NANDN U18749 ( .A(n18301), .B(n18300), .Z(n18305) );
  OR U18750 ( .A(n18303), .B(n18302), .Z(n18304) );
  AND U18751 ( .A(n18305), .B(n18304), .Z(n18389) );
  XNOR U18752 ( .A(n18390), .B(n18389), .Z(n18391) );
  NANDN U18753 ( .A(n18307), .B(n18306), .Z(n18311) );
  NANDN U18754 ( .A(n18309), .B(n18308), .Z(n18310) );
  NAND U18755 ( .A(n18311), .B(n18310), .Z(n18392) );
  XNOR U18756 ( .A(n18391), .B(n18392), .Z(n18337) );
  XOR U18757 ( .A(n18338), .B(n18337), .Z(n18396) );
  NANDN U18758 ( .A(n18313), .B(n18312), .Z(n18317) );
  NANDN U18759 ( .A(n18315), .B(n18314), .Z(n18316) );
  AND U18760 ( .A(n18317), .B(n18316), .Z(n18395) );
  XNOR U18761 ( .A(n18396), .B(n18395), .Z(n18397) );
  XOR U18762 ( .A(n18398), .B(n18397), .Z(n18330) );
  NANDN U18763 ( .A(n18319), .B(n18318), .Z(n18323) );
  NAND U18764 ( .A(n18321), .B(n18320), .Z(n18322) );
  AND U18765 ( .A(n18323), .B(n18322), .Z(n18329) );
  XNOR U18766 ( .A(n18330), .B(n18329), .Z(n18331) );
  XNOR U18767 ( .A(n18332), .B(n18331), .Z(n18401) );
  XNOR U18768 ( .A(sreg[485]), .B(n18401), .Z(n18403) );
  NANDN U18769 ( .A(sreg[484]), .B(n18324), .Z(n18328) );
  NAND U18770 ( .A(n18326), .B(n18325), .Z(n18327) );
  NAND U18771 ( .A(n18328), .B(n18327), .Z(n18402) );
  XNOR U18772 ( .A(n18403), .B(n18402), .Z(c[485]) );
  NANDN U18773 ( .A(n18330), .B(n18329), .Z(n18334) );
  NANDN U18774 ( .A(n18332), .B(n18331), .Z(n18333) );
  AND U18775 ( .A(n18334), .B(n18333), .Z(n18409) );
  NANDN U18776 ( .A(n18336), .B(n18335), .Z(n18340) );
  NAND U18777 ( .A(n18338), .B(n18337), .Z(n18339) );
  AND U18778 ( .A(n18340), .B(n18339), .Z(n18475) );
  NANDN U18779 ( .A(n18342), .B(n18341), .Z(n18346) );
  NANDN U18780 ( .A(n18344), .B(n18343), .Z(n18345) );
  AND U18781 ( .A(n18346), .B(n18345), .Z(n18462) );
  NAND U18782 ( .A(b[0]), .B(a[246]), .Z(n18347) );
  XNOR U18783 ( .A(b[1]), .B(n18347), .Z(n18349) );
  NANDN U18784 ( .A(b[0]), .B(a[245]), .Z(n18348) );
  NAND U18785 ( .A(n18349), .B(n18348), .Z(n18442) );
  NAND U18786 ( .A(n19808), .B(n18350), .Z(n18352) );
  XOR U18787 ( .A(b[13]), .B(a[234]), .Z(n18445) );
  NAND U18788 ( .A(n19768), .B(n18445), .Z(n18351) );
  AND U18789 ( .A(n18352), .B(n18351), .Z(n18440) );
  AND U18790 ( .A(b[15]), .B(a[230]), .Z(n18439) );
  XNOR U18791 ( .A(n18440), .B(n18439), .Z(n18441) );
  XNOR U18792 ( .A(n18442), .B(n18441), .Z(n18460) );
  NAND U18793 ( .A(n33), .B(n18353), .Z(n18355) );
  XOR U18794 ( .A(b[5]), .B(a[242]), .Z(n18451) );
  NAND U18795 ( .A(n19342), .B(n18451), .Z(n18354) );
  AND U18796 ( .A(n18355), .B(n18354), .Z(n18436) );
  NAND U18797 ( .A(n34), .B(n18356), .Z(n18358) );
  XOR U18798 ( .A(b[7]), .B(a[240]), .Z(n18454) );
  NAND U18799 ( .A(n19486), .B(n18454), .Z(n18357) );
  AND U18800 ( .A(n18358), .B(n18357), .Z(n18434) );
  NAND U18801 ( .A(n31), .B(n18359), .Z(n18361) );
  XOR U18802 ( .A(a[244]), .B(b[3]), .Z(n18457) );
  NAND U18803 ( .A(n32), .B(n18457), .Z(n18360) );
  NAND U18804 ( .A(n18361), .B(n18360), .Z(n18433) );
  XNOR U18805 ( .A(n18434), .B(n18433), .Z(n18435) );
  XOR U18806 ( .A(n18436), .B(n18435), .Z(n18461) );
  XOR U18807 ( .A(n18460), .B(n18461), .Z(n18463) );
  XOR U18808 ( .A(n18462), .B(n18463), .Z(n18413) );
  NANDN U18809 ( .A(n18363), .B(n18362), .Z(n18367) );
  OR U18810 ( .A(n18365), .B(n18364), .Z(n18366) );
  AND U18811 ( .A(n18367), .B(n18366), .Z(n18412) );
  XNOR U18812 ( .A(n18413), .B(n18412), .Z(n18415) );
  NAND U18813 ( .A(n18368), .B(n19724), .Z(n18370) );
  XOR U18814 ( .A(b[11]), .B(a[236]), .Z(n18418) );
  NAND U18815 ( .A(n19692), .B(n18418), .Z(n18369) );
  AND U18816 ( .A(n18370), .B(n18369), .Z(n18429) );
  NAND U18817 ( .A(n19838), .B(n18371), .Z(n18373) );
  XOR U18818 ( .A(b[15]), .B(a[232]), .Z(n18421) );
  NAND U18819 ( .A(n19805), .B(n18421), .Z(n18372) );
  AND U18820 ( .A(n18373), .B(n18372), .Z(n18428) );
  NAND U18821 ( .A(n35), .B(n18374), .Z(n18376) );
  XOR U18822 ( .A(b[9]), .B(a[238]), .Z(n18424) );
  NAND U18823 ( .A(n19598), .B(n18424), .Z(n18375) );
  NAND U18824 ( .A(n18376), .B(n18375), .Z(n18427) );
  XOR U18825 ( .A(n18428), .B(n18427), .Z(n18430) );
  XOR U18826 ( .A(n18429), .B(n18430), .Z(n18467) );
  NANDN U18827 ( .A(n18378), .B(n18377), .Z(n18382) );
  OR U18828 ( .A(n18380), .B(n18379), .Z(n18381) );
  AND U18829 ( .A(n18382), .B(n18381), .Z(n18466) );
  XNOR U18830 ( .A(n18467), .B(n18466), .Z(n18468) );
  NANDN U18831 ( .A(n18384), .B(n18383), .Z(n18388) );
  NANDN U18832 ( .A(n18386), .B(n18385), .Z(n18387) );
  NAND U18833 ( .A(n18388), .B(n18387), .Z(n18469) );
  XNOR U18834 ( .A(n18468), .B(n18469), .Z(n18414) );
  XOR U18835 ( .A(n18415), .B(n18414), .Z(n18473) );
  NANDN U18836 ( .A(n18390), .B(n18389), .Z(n18394) );
  NANDN U18837 ( .A(n18392), .B(n18391), .Z(n18393) );
  AND U18838 ( .A(n18394), .B(n18393), .Z(n18472) );
  XNOR U18839 ( .A(n18473), .B(n18472), .Z(n18474) );
  XOR U18840 ( .A(n18475), .B(n18474), .Z(n18407) );
  NANDN U18841 ( .A(n18396), .B(n18395), .Z(n18400) );
  NAND U18842 ( .A(n18398), .B(n18397), .Z(n18399) );
  AND U18843 ( .A(n18400), .B(n18399), .Z(n18406) );
  XNOR U18844 ( .A(n18407), .B(n18406), .Z(n18408) );
  XNOR U18845 ( .A(n18409), .B(n18408), .Z(n18478) );
  XNOR U18846 ( .A(sreg[486]), .B(n18478), .Z(n18480) );
  NANDN U18847 ( .A(sreg[485]), .B(n18401), .Z(n18405) );
  NAND U18848 ( .A(n18403), .B(n18402), .Z(n18404) );
  NAND U18849 ( .A(n18405), .B(n18404), .Z(n18479) );
  XNOR U18850 ( .A(n18480), .B(n18479), .Z(c[486]) );
  NANDN U18851 ( .A(n18407), .B(n18406), .Z(n18411) );
  NANDN U18852 ( .A(n18409), .B(n18408), .Z(n18410) );
  AND U18853 ( .A(n18411), .B(n18410), .Z(n18486) );
  NANDN U18854 ( .A(n18413), .B(n18412), .Z(n18417) );
  NAND U18855 ( .A(n18415), .B(n18414), .Z(n18416) );
  AND U18856 ( .A(n18417), .B(n18416), .Z(n18552) );
  NAND U18857 ( .A(n18418), .B(n19724), .Z(n18420) );
  XOR U18858 ( .A(b[11]), .B(a[237]), .Z(n18522) );
  NAND U18859 ( .A(n19692), .B(n18522), .Z(n18419) );
  AND U18860 ( .A(n18420), .B(n18419), .Z(n18533) );
  NAND U18861 ( .A(n19838), .B(n18421), .Z(n18423) );
  XOR U18862 ( .A(b[15]), .B(a[233]), .Z(n18525) );
  NAND U18863 ( .A(n19805), .B(n18525), .Z(n18422) );
  AND U18864 ( .A(n18423), .B(n18422), .Z(n18532) );
  NAND U18865 ( .A(n35), .B(n18424), .Z(n18426) );
  XOR U18866 ( .A(b[9]), .B(a[239]), .Z(n18528) );
  NAND U18867 ( .A(n19598), .B(n18528), .Z(n18425) );
  NAND U18868 ( .A(n18426), .B(n18425), .Z(n18531) );
  XOR U18869 ( .A(n18532), .B(n18531), .Z(n18534) );
  XOR U18870 ( .A(n18533), .B(n18534), .Z(n18544) );
  NANDN U18871 ( .A(n18428), .B(n18427), .Z(n18432) );
  OR U18872 ( .A(n18430), .B(n18429), .Z(n18431) );
  AND U18873 ( .A(n18432), .B(n18431), .Z(n18543) );
  XNOR U18874 ( .A(n18544), .B(n18543), .Z(n18545) );
  NANDN U18875 ( .A(n18434), .B(n18433), .Z(n18438) );
  NANDN U18876 ( .A(n18436), .B(n18435), .Z(n18437) );
  NAND U18877 ( .A(n18438), .B(n18437), .Z(n18546) );
  XNOR U18878 ( .A(n18545), .B(n18546), .Z(n18492) );
  NANDN U18879 ( .A(n18440), .B(n18439), .Z(n18444) );
  NANDN U18880 ( .A(n18442), .B(n18441), .Z(n18443) );
  AND U18881 ( .A(n18444), .B(n18443), .Z(n18518) );
  NAND U18882 ( .A(n19808), .B(n18445), .Z(n18447) );
  XOR U18883 ( .A(b[13]), .B(a[235]), .Z(n18501) );
  NAND U18884 ( .A(n19768), .B(n18501), .Z(n18446) );
  AND U18885 ( .A(n18447), .B(n18446), .Z(n18496) );
  AND U18886 ( .A(b[15]), .B(a[231]), .Z(n18495) );
  XNOR U18887 ( .A(n18496), .B(n18495), .Z(n18497) );
  NAND U18888 ( .A(b[0]), .B(a[247]), .Z(n18448) );
  XNOR U18889 ( .A(b[1]), .B(n18448), .Z(n18450) );
  NANDN U18890 ( .A(b[0]), .B(a[246]), .Z(n18449) );
  NAND U18891 ( .A(n18450), .B(n18449), .Z(n18498) );
  XNOR U18892 ( .A(n18497), .B(n18498), .Z(n18516) );
  NAND U18893 ( .A(n33), .B(n18451), .Z(n18453) );
  XOR U18894 ( .A(b[5]), .B(a[243]), .Z(n18507) );
  NAND U18895 ( .A(n19342), .B(n18507), .Z(n18452) );
  AND U18896 ( .A(n18453), .B(n18452), .Z(n18540) );
  NAND U18897 ( .A(n34), .B(n18454), .Z(n18456) );
  XOR U18898 ( .A(b[7]), .B(a[241]), .Z(n18510) );
  NAND U18899 ( .A(n19486), .B(n18510), .Z(n18455) );
  AND U18900 ( .A(n18456), .B(n18455), .Z(n18538) );
  NAND U18901 ( .A(n31), .B(n18457), .Z(n18459) );
  XOR U18902 ( .A(b[3]), .B(a[245]), .Z(n18513) );
  NAND U18903 ( .A(n32), .B(n18513), .Z(n18458) );
  NAND U18904 ( .A(n18459), .B(n18458), .Z(n18537) );
  XNOR U18905 ( .A(n18538), .B(n18537), .Z(n18539) );
  XOR U18906 ( .A(n18540), .B(n18539), .Z(n18517) );
  XOR U18907 ( .A(n18516), .B(n18517), .Z(n18519) );
  XOR U18908 ( .A(n18518), .B(n18519), .Z(n18490) );
  NANDN U18909 ( .A(n18461), .B(n18460), .Z(n18465) );
  OR U18910 ( .A(n18463), .B(n18462), .Z(n18464) );
  AND U18911 ( .A(n18465), .B(n18464), .Z(n18489) );
  XNOR U18912 ( .A(n18490), .B(n18489), .Z(n18491) );
  XOR U18913 ( .A(n18492), .B(n18491), .Z(n18550) );
  NANDN U18914 ( .A(n18467), .B(n18466), .Z(n18471) );
  NANDN U18915 ( .A(n18469), .B(n18468), .Z(n18470) );
  AND U18916 ( .A(n18471), .B(n18470), .Z(n18549) );
  XNOR U18917 ( .A(n18550), .B(n18549), .Z(n18551) );
  XOR U18918 ( .A(n18552), .B(n18551), .Z(n18484) );
  NANDN U18919 ( .A(n18473), .B(n18472), .Z(n18477) );
  NAND U18920 ( .A(n18475), .B(n18474), .Z(n18476) );
  AND U18921 ( .A(n18477), .B(n18476), .Z(n18483) );
  XNOR U18922 ( .A(n18484), .B(n18483), .Z(n18485) );
  XNOR U18923 ( .A(n18486), .B(n18485), .Z(n18555) );
  XNOR U18924 ( .A(sreg[487]), .B(n18555), .Z(n18557) );
  NANDN U18925 ( .A(sreg[486]), .B(n18478), .Z(n18482) );
  NAND U18926 ( .A(n18480), .B(n18479), .Z(n18481) );
  NAND U18927 ( .A(n18482), .B(n18481), .Z(n18556) );
  XNOR U18928 ( .A(n18557), .B(n18556), .Z(c[487]) );
  NANDN U18929 ( .A(n18484), .B(n18483), .Z(n18488) );
  NANDN U18930 ( .A(n18486), .B(n18485), .Z(n18487) );
  AND U18931 ( .A(n18488), .B(n18487), .Z(n18563) );
  NANDN U18932 ( .A(n18490), .B(n18489), .Z(n18494) );
  NAND U18933 ( .A(n18492), .B(n18491), .Z(n18493) );
  AND U18934 ( .A(n18494), .B(n18493), .Z(n18629) );
  NANDN U18935 ( .A(n18496), .B(n18495), .Z(n18500) );
  NANDN U18936 ( .A(n18498), .B(n18497), .Z(n18499) );
  AND U18937 ( .A(n18500), .B(n18499), .Z(n18616) );
  NAND U18938 ( .A(n19808), .B(n18501), .Z(n18503) );
  XOR U18939 ( .A(b[13]), .B(a[236]), .Z(n18602) );
  NAND U18940 ( .A(n19768), .B(n18602), .Z(n18502) );
  AND U18941 ( .A(n18503), .B(n18502), .Z(n18594) );
  AND U18942 ( .A(b[15]), .B(a[232]), .Z(n18593) );
  XNOR U18943 ( .A(n18594), .B(n18593), .Z(n18595) );
  NAND U18944 ( .A(b[0]), .B(a[248]), .Z(n18504) );
  XNOR U18945 ( .A(b[1]), .B(n18504), .Z(n18506) );
  NANDN U18946 ( .A(b[0]), .B(a[247]), .Z(n18505) );
  NAND U18947 ( .A(n18506), .B(n18505), .Z(n18596) );
  XNOR U18948 ( .A(n18595), .B(n18596), .Z(n18614) );
  NAND U18949 ( .A(n33), .B(n18507), .Z(n18509) );
  XOR U18950 ( .A(b[5]), .B(a[244]), .Z(n18605) );
  NAND U18951 ( .A(n19342), .B(n18605), .Z(n18508) );
  AND U18952 ( .A(n18509), .B(n18508), .Z(n18590) );
  NAND U18953 ( .A(n34), .B(n18510), .Z(n18512) );
  XOR U18954 ( .A(b[7]), .B(a[242]), .Z(n18608) );
  NAND U18955 ( .A(n19486), .B(n18608), .Z(n18511) );
  AND U18956 ( .A(n18512), .B(n18511), .Z(n18588) );
  NAND U18957 ( .A(n31), .B(n18513), .Z(n18515) );
  XOR U18958 ( .A(a[246]), .B(b[3]), .Z(n18611) );
  NAND U18959 ( .A(n32), .B(n18611), .Z(n18514) );
  NAND U18960 ( .A(n18515), .B(n18514), .Z(n18587) );
  XNOR U18961 ( .A(n18588), .B(n18587), .Z(n18589) );
  XOR U18962 ( .A(n18590), .B(n18589), .Z(n18615) );
  XOR U18963 ( .A(n18614), .B(n18615), .Z(n18617) );
  XOR U18964 ( .A(n18616), .B(n18617), .Z(n18567) );
  NANDN U18965 ( .A(n18517), .B(n18516), .Z(n18521) );
  OR U18966 ( .A(n18519), .B(n18518), .Z(n18520) );
  AND U18967 ( .A(n18521), .B(n18520), .Z(n18566) );
  XNOR U18968 ( .A(n18567), .B(n18566), .Z(n18569) );
  NAND U18969 ( .A(n18522), .B(n19724), .Z(n18524) );
  XOR U18970 ( .A(b[11]), .B(a[238]), .Z(n18572) );
  NAND U18971 ( .A(n19692), .B(n18572), .Z(n18523) );
  AND U18972 ( .A(n18524), .B(n18523), .Z(n18583) );
  NAND U18973 ( .A(n19838), .B(n18525), .Z(n18527) );
  XOR U18974 ( .A(b[15]), .B(a[234]), .Z(n18575) );
  NAND U18975 ( .A(n19805), .B(n18575), .Z(n18526) );
  AND U18976 ( .A(n18527), .B(n18526), .Z(n18582) );
  NAND U18977 ( .A(n35), .B(n18528), .Z(n18530) );
  XOR U18978 ( .A(b[9]), .B(a[240]), .Z(n18578) );
  NAND U18979 ( .A(n19598), .B(n18578), .Z(n18529) );
  NAND U18980 ( .A(n18530), .B(n18529), .Z(n18581) );
  XOR U18981 ( .A(n18582), .B(n18581), .Z(n18584) );
  XOR U18982 ( .A(n18583), .B(n18584), .Z(n18621) );
  NANDN U18983 ( .A(n18532), .B(n18531), .Z(n18536) );
  OR U18984 ( .A(n18534), .B(n18533), .Z(n18535) );
  AND U18985 ( .A(n18536), .B(n18535), .Z(n18620) );
  XNOR U18986 ( .A(n18621), .B(n18620), .Z(n18622) );
  NANDN U18987 ( .A(n18538), .B(n18537), .Z(n18542) );
  NANDN U18988 ( .A(n18540), .B(n18539), .Z(n18541) );
  NAND U18989 ( .A(n18542), .B(n18541), .Z(n18623) );
  XNOR U18990 ( .A(n18622), .B(n18623), .Z(n18568) );
  XOR U18991 ( .A(n18569), .B(n18568), .Z(n18627) );
  NANDN U18992 ( .A(n18544), .B(n18543), .Z(n18548) );
  NANDN U18993 ( .A(n18546), .B(n18545), .Z(n18547) );
  AND U18994 ( .A(n18548), .B(n18547), .Z(n18626) );
  XNOR U18995 ( .A(n18627), .B(n18626), .Z(n18628) );
  XOR U18996 ( .A(n18629), .B(n18628), .Z(n18561) );
  NANDN U18997 ( .A(n18550), .B(n18549), .Z(n18554) );
  NAND U18998 ( .A(n18552), .B(n18551), .Z(n18553) );
  AND U18999 ( .A(n18554), .B(n18553), .Z(n18560) );
  XNOR U19000 ( .A(n18561), .B(n18560), .Z(n18562) );
  XNOR U19001 ( .A(n18563), .B(n18562), .Z(n18632) );
  XNOR U19002 ( .A(sreg[488]), .B(n18632), .Z(n18634) );
  NANDN U19003 ( .A(sreg[487]), .B(n18555), .Z(n18559) );
  NAND U19004 ( .A(n18557), .B(n18556), .Z(n18558) );
  NAND U19005 ( .A(n18559), .B(n18558), .Z(n18633) );
  XNOR U19006 ( .A(n18634), .B(n18633), .Z(c[488]) );
  NANDN U19007 ( .A(n18561), .B(n18560), .Z(n18565) );
  NANDN U19008 ( .A(n18563), .B(n18562), .Z(n18564) );
  AND U19009 ( .A(n18565), .B(n18564), .Z(n18640) );
  NANDN U19010 ( .A(n18567), .B(n18566), .Z(n18571) );
  NAND U19011 ( .A(n18569), .B(n18568), .Z(n18570) );
  AND U19012 ( .A(n18571), .B(n18570), .Z(n18706) );
  NAND U19013 ( .A(n18572), .B(n19724), .Z(n18574) );
  XOR U19014 ( .A(b[11]), .B(a[239]), .Z(n18676) );
  NAND U19015 ( .A(n19692), .B(n18676), .Z(n18573) );
  AND U19016 ( .A(n18574), .B(n18573), .Z(n18687) );
  NAND U19017 ( .A(n19838), .B(n18575), .Z(n18577) );
  XOR U19018 ( .A(b[15]), .B(a[235]), .Z(n18679) );
  NAND U19019 ( .A(n19805), .B(n18679), .Z(n18576) );
  AND U19020 ( .A(n18577), .B(n18576), .Z(n18686) );
  NAND U19021 ( .A(n35), .B(n18578), .Z(n18580) );
  XOR U19022 ( .A(b[9]), .B(a[241]), .Z(n18682) );
  NAND U19023 ( .A(n19598), .B(n18682), .Z(n18579) );
  NAND U19024 ( .A(n18580), .B(n18579), .Z(n18685) );
  XOR U19025 ( .A(n18686), .B(n18685), .Z(n18688) );
  XOR U19026 ( .A(n18687), .B(n18688), .Z(n18698) );
  NANDN U19027 ( .A(n18582), .B(n18581), .Z(n18586) );
  OR U19028 ( .A(n18584), .B(n18583), .Z(n18585) );
  AND U19029 ( .A(n18586), .B(n18585), .Z(n18697) );
  XNOR U19030 ( .A(n18698), .B(n18697), .Z(n18699) );
  NANDN U19031 ( .A(n18588), .B(n18587), .Z(n18592) );
  NANDN U19032 ( .A(n18590), .B(n18589), .Z(n18591) );
  NAND U19033 ( .A(n18592), .B(n18591), .Z(n18700) );
  XNOR U19034 ( .A(n18699), .B(n18700), .Z(n18646) );
  NANDN U19035 ( .A(n18594), .B(n18593), .Z(n18598) );
  NANDN U19036 ( .A(n18596), .B(n18595), .Z(n18597) );
  AND U19037 ( .A(n18598), .B(n18597), .Z(n18672) );
  NAND U19038 ( .A(b[0]), .B(a[249]), .Z(n18599) );
  XNOR U19039 ( .A(b[1]), .B(n18599), .Z(n18601) );
  NANDN U19040 ( .A(b[0]), .B(a[248]), .Z(n18600) );
  NAND U19041 ( .A(n18601), .B(n18600), .Z(n18652) );
  NAND U19042 ( .A(n19808), .B(n18602), .Z(n18604) );
  XOR U19043 ( .A(b[13]), .B(a[237]), .Z(n18655) );
  NAND U19044 ( .A(n19768), .B(n18655), .Z(n18603) );
  AND U19045 ( .A(n18604), .B(n18603), .Z(n18650) );
  AND U19046 ( .A(b[15]), .B(a[233]), .Z(n18649) );
  XNOR U19047 ( .A(n18650), .B(n18649), .Z(n18651) );
  XNOR U19048 ( .A(n18652), .B(n18651), .Z(n18670) );
  NAND U19049 ( .A(n33), .B(n18605), .Z(n18607) );
  XOR U19050 ( .A(b[5]), .B(a[245]), .Z(n18661) );
  NAND U19051 ( .A(n19342), .B(n18661), .Z(n18606) );
  AND U19052 ( .A(n18607), .B(n18606), .Z(n18694) );
  NAND U19053 ( .A(n34), .B(n18608), .Z(n18610) );
  XOR U19054 ( .A(b[7]), .B(a[243]), .Z(n18664) );
  NAND U19055 ( .A(n19486), .B(n18664), .Z(n18609) );
  AND U19056 ( .A(n18610), .B(n18609), .Z(n18692) );
  NAND U19057 ( .A(n31), .B(n18611), .Z(n18613) );
  XOR U19058 ( .A(a[247]), .B(b[3]), .Z(n18667) );
  NAND U19059 ( .A(n32), .B(n18667), .Z(n18612) );
  NAND U19060 ( .A(n18613), .B(n18612), .Z(n18691) );
  XNOR U19061 ( .A(n18692), .B(n18691), .Z(n18693) );
  XOR U19062 ( .A(n18694), .B(n18693), .Z(n18671) );
  XOR U19063 ( .A(n18670), .B(n18671), .Z(n18673) );
  XOR U19064 ( .A(n18672), .B(n18673), .Z(n18644) );
  NANDN U19065 ( .A(n18615), .B(n18614), .Z(n18619) );
  OR U19066 ( .A(n18617), .B(n18616), .Z(n18618) );
  AND U19067 ( .A(n18619), .B(n18618), .Z(n18643) );
  XNOR U19068 ( .A(n18644), .B(n18643), .Z(n18645) );
  XOR U19069 ( .A(n18646), .B(n18645), .Z(n18704) );
  NANDN U19070 ( .A(n18621), .B(n18620), .Z(n18625) );
  NANDN U19071 ( .A(n18623), .B(n18622), .Z(n18624) );
  AND U19072 ( .A(n18625), .B(n18624), .Z(n18703) );
  XNOR U19073 ( .A(n18704), .B(n18703), .Z(n18705) );
  XOR U19074 ( .A(n18706), .B(n18705), .Z(n18638) );
  NANDN U19075 ( .A(n18627), .B(n18626), .Z(n18631) );
  NAND U19076 ( .A(n18629), .B(n18628), .Z(n18630) );
  AND U19077 ( .A(n18631), .B(n18630), .Z(n18637) );
  XNOR U19078 ( .A(n18638), .B(n18637), .Z(n18639) );
  XNOR U19079 ( .A(n18640), .B(n18639), .Z(n18709) );
  XNOR U19080 ( .A(sreg[489]), .B(n18709), .Z(n18711) );
  NANDN U19081 ( .A(sreg[488]), .B(n18632), .Z(n18636) );
  NAND U19082 ( .A(n18634), .B(n18633), .Z(n18635) );
  NAND U19083 ( .A(n18636), .B(n18635), .Z(n18710) );
  XNOR U19084 ( .A(n18711), .B(n18710), .Z(c[489]) );
  NANDN U19085 ( .A(n18638), .B(n18637), .Z(n18642) );
  NANDN U19086 ( .A(n18640), .B(n18639), .Z(n18641) );
  AND U19087 ( .A(n18642), .B(n18641), .Z(n18717) );
  NANDN U19088 ( .A(n18644), .B(n18643), .Z(n18648) );
  NAND U19089 ( .A(n18646), .B(n18645), .Z(n18647) );
  AND U19090 ( .A(n18648), .B(n18647), .Z(n18783) );
  NANDN U19091 ( .A(n18650), .B(n18649), .Z(n18654) );
  NANDN U19092 ( .A(n18652), .B(n18651), .Z(n18653) );
  AND U19093 ( .A(n18654), .B(n18653), .Z(n18749) );
  NAND U19094 ( .A(n19808), .B(n18655), .Z(n18657) );
  XOR U19095 ( .A(b[13]), .B(a[238]), .Z(n18732) );
  NAND U19096 ( .A(n19768), .B(n18732), .Z(n18656) );
  AND U19097 ( .A(n18657), .B(n18656), .Z(n18727) );
  AND U19098 ( .A(b[15]), .B(a[234]), .Z(n18726) );
  XNOR U19099 ( .A(n18727), .B(n18726), .Z(n18728) );
  NAND U19100 ( .A(b[0]), .B(a[250]), .Z(n18658) );
  XNOR U19101 ( .A(b[1]), .B(n18658), .Z(n18660) );
  NANDN U19102 ( .A(b[0]), .B(a[249]), .Z(n18659) );
  NAND U19103 ( .A(n18660), .B(n18659), .Z(n18729) );
  XNOR U19104 ( .A(n18728), .B(n18729), .Z(n18747) );
  NAND U19105 ( .A(n33), .B(n18661), .Z(n18663) );
  XOR U19106 ( .A(b[5]), .B(a[246]), .Z(n18738) );
  NAND U19107 ( .A(n19342), .B(n18738), .Z(n18662) );
  AND U19108 ( .A(n18663), .B(n18662), .Z(n18771) );
  NAND U19109 ( .A(n34), .B(n18664), .Z(n18666) );
  XOR U19110 ( .A(b[7]), .B(a[244]), .Z(n18741) );
  NAND U19111 ( .A(n19486), .B(n18741), .Z(n18665) );
  AND U19112 ( .A(n18666), .B(n18665), .Z(n18769) );
  NAND U19113 ( .A(n31), .B(n18667), .Z(n18669) );
  XOR U19114 ( .A(a[248]), .B(b[3]), .Z(n18744) );
  NAND U19115 ( .A(n32), .B(n18744), .Z(n18668) );
  NAND U19116 ( .A(n18669), .B(n18668), .Z(n18768) );
  XNOR U19117 ( .A(n18769), .B(n18768), .Z(n18770) );
  XOR U19118 ( .A(n18771), .B(n18770), .Z(n18748) );
  XOR U19119 ( .A(n18747), .B(n18748), .Z(n18750) );
  XOR U19120 ( .A(n18749), .B(n18750), .Z(n18721) );
  NANDN U19121 ( .A(n18671), .B(n18670), .Z(n18675) );
  OR U19122 ( .A(n18673), .B(n18672), .Z(n18674) );
  AND U19123 ( .A(n18675), .B(n18674), .Z(n18720) );
  XNOR U19124 ( .A(n18721), .B(n18720), .Z(n18723) );
  NAND U19125 ( .A(n18676), .B(n19724), .Z(n18678) );
  XOR U19126 ( .A(b[11]), .B(a[240]), .Z(n18753) );
  NAND U19127 ( .A(n19692), .B(n18753), .Z(n18677) );
  AND U19128 ( .A(n18678), .B(n18677), .Z(n18764) );
  NAND U19129 ( .A(n19838), .B(n18679), .Z(n18681) );
  XOR U19130 ( .A(b[15]), .B(a[236]), .Z(n18756) );
  NAND U19131 ( .A(n19805), .B(n18756), .Z(n18680) );
  AND U19132 ( .A(n18681), .B(n18680), .Z(n18763) );
  NAND U19133 ( .A(n35), .B(n18682), .Z(n18684) );
  XOR U19134 ( .A(b[9]), .B(a[242]), .Z(n18759) );
  NAND U19135 ( .A(n19598), .B(n18759), .Z(n18683) );
  NAND U19136 ( .A(n18684), .B(n18683), .Z(n18762) );
  XOR U19137 ( .A(n18763), .B(n18762), .Z(n18765) );
  XOR U19138 ( .A(n18764), .B(n18765), .Z(n18775) );
  NANDN U19139 ( .A(n18686), .B(n18685), .Z(n18690) );
  OR U19140 ( .A(n18688), .B(n18687), .Z(n18689) );
  AND U19141 ( .A(n18690), .B(n18689), .Z(n18774) );
  XNOR U19142 ( .A(n18775), .B(n18774), .Z(n18776) );
  NANDN U19143 ( .A(n18692), .B(n18691), .Z(n18696) );
  NANDN U19144 ( .A(n18694), .B(n18693), .Z(n18695) );
  NAND U19145 ( .A(n18696), .B(n18695), .Z(n18777) );
  XNOR U19146 ( .A(n18776), .B(n18777), .Z(n18722) );
  XOR U19147 ( .A(n18723), .B(n18722), .Z(n18781) );
  NANDN U19148 ( .A(n18698), .B(n18697), .Z(n18702) );
  NANDN U19149 ( .A(n18700), .B(n18699), .Z(n18701) );
  AND U19150 ( .A(n18702), .B(n18701), .Z(n18780) );
  XNOR U19151 ( .A(n18781), .B(n18780), .Z(n18782) );
  XOR U19152 ( .A(n18783), .B(n18782), .Z(n18715) );
  NANDN U19153 ( .A(n18704), .B(n18703), .Z(n18708) );
  NAND U19154 ( .A(n18706), .B(n18705), .Z(n18707) );
  AND U19155 ( .A(n18708), .B(n18707), .Z(n18714) );
  XNOR U19156 ( .A(n18715), .B(n18714), .Z(n18716) );
  XNOR U19157 ( .A(n18717), .B(n18716), .Z(n18786) );
  XNOR U19158 ( .A(sreg[490]), .B(n18786), .Z(n18788) );
  NANDN U19159 ( .A(sreg[489]), .B(n18709), .Z(n18713) );
  NAND U19160 ( .A(n18711), .B(n18710), .Z(n18712) );
  NAND U19161 ( .A(n18713), .B(n18712), .Z(n18787) );
  XNOR U19162 ( .A(n18788), .B(n18787), .Z(c[490]) );
  NANDN U19163 ( .A(n18715), .B(n18714), .Z(n18719) );
  NANDN U19164 ( .A(n18717), .B(n18716), .Z(n18718) );
  AND U19165 ( .A(n18719), .B(n18718), .Z(n18794) );
  NANDN U19166 ( .A(n18721), .B(n18720), .Z(n18725) );
  NAND U19167 ( .A(n18723), .B(n18722), .Z(n18724) );
  AND U19168 ( .A(n18725), .B(n18724), .Z(n18860) );
  NANDN U19169 ( .A(n18727), .B(n18726), .Z(n18731) );
  NANDN U19170 ( .A(n18729), .B(n18728), .Z(n18730) );
  AND U19171 ( .A(n18731), .B(n18730), .Z(n18847) );
  NAND U19172 ( .A(n19808), .B(n18732), .Z(n18734) );
  XOR U19173 ( .A(b[13]), .B(a[239]), .Z(n18830) );
  NAND U19174 ( .A(n19768), .B(n18830), .Z(n18733) );
  AND U19175 ( .A(n18734), .B(n18733), .Z(n18825) );
  AND U19176 ( .A(b[15]), .B(a[235]), .Z(n18824) );
  XNOR U19177 ( .A(n18825), .B(n18824), .Z(n18826) );
  NAND U19178 ( .A(b[0]), .B(a[251]), .Z(n18735) );
  XNOR U19179 ( .A(b[1]), .B(n18735), .Z(n18737) );
  NANDN U19180 ( .A(b[0]), .B(a[250]), .Z(n18736) );
  NAND U19181 ( .A(n18737), .B(n18736), .Z(n18827) );
  XNOR U19182 ( .A(n18826), .B(n18827), .Z(n18845) );
  NAND U19183 ( .A(n33), .B(n18738), .Z(n18740) );
  XOR U19184 ( .A(b[5]), .B(a[247]), .Z(n18836) );
  NAND U19185 ( .A(n19342), .B(n18836), .Z(n18739) );
  AND U19186 ( .A(n18740), .B(n18739), .Z(n18821) );
  NAND U19187 ( .A(n34), .B(n18741), .Z(n18743) );
  XOR U19188 ( .A(b[7]), .B(a[245]), .Z(n18839) );
  NAND U19189 ( .A(n19486), .B(n18839), .Z(n18742) );
  AND U19190 ( .A(n18743), .B(n18742), .Z(n18819) );
  NAND U19191 ( .A(n31), .B(n18744), .Z(n18746) );
  XOR U19192 ( .A(a[249]), .B(b[3]), .Z(n18842) );
  NAND U19193 ( .A(n32), .B(n18842), .Z(n18745) );
  NAND U19194 ( .A(n18746), .B(n18745), .Z(n18818) );
  XNOR U19195 ( .A(n18819), .B(n18818), .Z(n18820) );
  XOR U19196 ( .A(n18821), .B(n18820), .Z(n18846) );
  XOR U19197 ( .A(n18845), .B(n18846), .Z(n18848) );
  XOR U19198 ( .A(n18847), .B(n18848), .Z(n18798) );
  NANDN U19199 ( .A(n18748), .B(n18747), .Z(n18752) );
  OR U19200 ( .A(n18750), .B(n18749), .Z(n18751) );
  AND U19201 ( .A(n18752), .B(n18751), .Z(n18797) );
  XNOR U19202 ( .A(n18798), .B(n18797), .Z(n18800) );
  NAND U19203 ( .A(n18753), .B(n19724), .Z(n18755) );
  XOR U19204 ( .A(b[11]), .B(a[241]), .Z(n18803) );
  NAND U19205 ( .A(n19692), .B(n18803), .Z(n18754) );
  AND U19206 ( .A(n18755), .B(n18754), .Z(n18814) );
  NAND U19207 ( .A(n19838), .B(n18756), .Z(n18758) );
  XOR U19208 ( .A(b[15]), .B(a[237]), .Z(n18806) );
  NAND U19209 ( .A(n19805), .B(n18806), .Z(n18757) );
  AND U19210 ( .A(n18758), .B(n18757), .Z(n18813) );
  NAND U19211 ( .A(n35), .B(n18759), .Z(n18761) );
  XOR U19212 ( .A(b[9]), .B(a[243]), .Z(n18809) );
  NAND U19213 ( .A(n19598), .B(n18809), .Z(n18760) );
  NAND U19214 ( .A(n18761), .B(n18760), .Z(n18812) );
  XOR U19215 ( .A(n18813), .B(n18812), .Z(n18815) );
  XOR U19216 ( .A(n18814), .B(n18815), .Z(n18852) );
  NANDN U19217 ( .A(n18763), .B(n18762), .Z(n18767) );
  OR U19218 ( .A(n18765), .B(n18764), .Z(n18766) );
  AND U19219 ( .A(n18767), .B(n18766), .Z(n18851) );
  XNOR U19220 ( .A(n18852), .B(n18851), .Z(n18853) );
  NANDN U19221 ( .A(n18769), .B(n18768), .Z(n18773) );
  NANDN U19222 ( .A(n18771), .B(n18770), .Z(n18772) );
  NAND U19223 ( .A(n18773), .B(n18772), .Z(n18854) );
  XNOR U19224 ( .A(n18853), .B(n18854), .Z(n18799) );
  XOR U19225 ( .A(n18800), .B(n18799), .Z(n18858) );
  NANDN U19226 ( .A(n18775), .B(n18774), .Z(n18779) );
  NANDN U19227 ( .A(n18777), .B(n18776), .Z(n18778) );
  AND U19228 ( .A(n18779), .B(n18778), .Z(n18857) );
  XNOR U19229 ( .A(n18858), .B(n18857), .Z(n18859) );
  XOR U19230 ( .A(n18860), .B(n18859), .Z(n18792) );
  NANDN U19231 ( .A(n18781), .B(n18780), .Z(n18785) );
  NAND U19232 ( .A(n18783), .B(n18782), .Z(n18784) );
  AND U19233 ( .A(n18785), .B(n18784), .Z(n18791) );
  XNOR U19234 ( .A(n18792), .B(n18791), .Z(n18793) );
  XNOR U19235 ( .A(n18794), .B(n18793), .Z(n18863) );
  XNOR U19236 ( .A(sreg[491]), .B(n18863), .Z(n18865) );
  NANDN U19237 ( .A(sreg[490]), .B(n18786), .Z(n18790) );
  NAND U19238 ( .A(n18788), .B(n18787), .Z(n18789) );
  NAND U19239 ( .A(n18790), .B(n18789), .Z(n18864) );
  XNOR U19240 ( .A(n18865), .B(n18864), .Z(c[491]) );
  NANDN U19241 ( .A(n18792), .B(n18791), .Z(n18796) );
  NANDN U19242 ( .A(n18794), .B(n18793), .Z(n18795) );
  AND U19243 ( .A(n18796), .B(n18795), .Z(n18871) );
  NANDN U19244 ( .A(n18798), .B(n18797), .Z(n18802) );
  NAND U19245 ( .A(n18800), .B(n18799), .Z(n18801) );
  AND U19246 ( .A(n18802), .B(n18801), .Z(n18933) );
  NAND U19247 ( .A(n18803), .B(n19724), .Z(n18805) );
  XOR U19248 ( .A(b[11]), .B(a[242]), .Z(n18903) );
  NAND U19249 ( .A(n19692), .B(n18903), .Z(n18804) );
  AND U19250 ( .A(n18805), .B(n18804), .Z(n18915) );
  NAND U19251 ( .A(n19838), .B(n18806), .Z(n18808) );
  XOR U19252 ( .A(b[15]), .B(a[238]), .Z(n18906) );
  NAND U19253 ( .A(n19805), .B(n18906), .Z(n18807) );
  AND U19254 ( .A(n18808), .B(n18807), .Z(n18913) );
  NAND U19255 ( .A(n35), .B(n18809), .Z(n18811) );
  XOR U19256 ( .A(b[9]), .B(a[244]), .Z(n18909) );
  NAND U19257 ( .A(n19598), .B(n18909), .Z(n18810) );
  NAND U19258 ( .A(n18811), .B(n18810), .Z(n18912) );
  XNOR U19259 ( .A(n18913), .B(n18912), .Z(n18914) );
  XOR U19260 ( .A(n18915), .B(n18914), .Z(n18925) );
  NANDN U19261 ( .A(n18813), .B(n18812), .Z(n18817) );
  OR U19262 ( .A(n18815), .B(n18814), .Z(n18816) );
  AND U19263 ( .A(n18817), .B(n18816), .Z(n18924) );
  XOR U19264 ( .A(n18925), .B(n18924), .Z(n18926) );
  NANDN U19265 ( .A(n18819), .B(n18818), .Z(n18823) );
  NANDN U19266 ( .A(n18821), .B(n18820), .Z(n18822) );
  NAND U19267 ( .A(n18823), .B(n18822), .Z(n18927) );
  XNOR U19268 ( .A(n18926), .B(n18927), .Z(n18877) );
  NANDN U19269 ( .A(n18825), .B(n18824), .Z(n18829) );
  NANDN U19270 ( .A(n18827), .B(n18826), .Z(n18828) );
  AND U19271 ( .A(n18829), .B(n18828), .Z(n18902) );
  NAND U19272 ( .A(n19808), .B(n18830), .Z(n18832) );
  XOR U19273 ( .A(b[13]), .B(a[240]), .Z(n18887) );
  NAND U19274 ( .A(n19768), .B(n18887), .Z(n18831) );
  AND U19275 ( .A(n18832), .B(n18831), .Z(n18879) );
  AND U19276 ( .A(b[15]), .B(a[236]), .Z(n18878) );
  XNOR U19277 ( .A(n18879), .B(n18878), .Z(n18880) );
  NAND U19278 ( .A(b[0]), .B(a[252]), .Z(n18833) );
  XNOR U19279 ( .A(b[1]), .B(n18833), .Z(n18835) );
  NANDN U19280 ( .A(b[0]), .B(a[251]), .Z(n18834) );
  NAND U19281 ( .A(n18835), .B(n18834), .Z(n18881) );
  XNOR U19282 ( .A(n18880), .B(n18881), .Z(n18900) );
  NAND U19283 ( .A(n33), .B(n18836), .Z(n18838) );
  XOR U19284 ( .A(a[248]), .B(b[5]), .Z(n18890) );
  NAND U19285 ( .A(n19342), .B(n18890), .Z(n18837) );
  NAND U19286 ( .A(n18838), .B(n18837), .Z(n18921) );
  NAND U19287 ( .A(n34), .B(n18839), .Z(n18841) );
  XOR U19288 ( .A(b[7]), .B(a[246]), .Z(n18893) );
  NAND U19289 ( .A(n19486), .B(n18893), .Z(n18840) );
  NAND U19290 ( .A(n18841), .B(n18840), .Z(n18919) );
  NAND U19291 ( .A(n31), .B(n18842), .Z(n18844) );
  XOR U19292 ( .A(a[250]), .B(b[3]), .Z(n18896) );
  NAND U19293 ( .A(n32), .B(n18896), .Z(n18843) );
  NAND U19294 ( .A(n18844), .B(n18843), .Z(n18918) );
  XNOR U19295 ( .A(n18900), .B(n18899), .Z(n18901) );
  XNOR U19296 ( .A(n18902), .B(n18901), .Z(n18874) );
  NANDN U19297 ( .A(n18846), .B(n18845), .Z(n18850) );
  OR U19298 ( .A(n18848), .B(n18847), .Z(n18849) );
  AND U19299 ( .A(n18850), .B(n18849), .Z(n18875) );
  XNOR U19300 ( .A(n18874), .B(n18875), .Z(n18876) );
  XOR U19301 ( .A(n18877), .B(n18876), .Z(n18931) );
  NANDN U19302 ( .A(n18852), .B(n18851), .Z(n18856) );
  NANDN U19303 ( .A(n18854), .B(n18853), .Z(n18855) );
  AND U19304 ( .A(n18856), .B(n18855), .Z(n18930) );
  XNOR U19305 ( .A(n18931), .B(n18930), .Z(n18932) );
  XOR U19306 ( .A(n18933), .B(n18932), .Z(n18869) );
  NANDN U19307 ( .A(n18858), .B(n18857), .Z(n18862) );
  NAND U19308 ( .A(n18860), .B(n18859), .Z(n18861) );
  AND U19309 ( .A(n18862), .B(n18861), .Z(n18868) );
  XNOR U19310 ( .A(n18869), .B(n18868), .Z(n18870) );
  XNOR U19311 ( .A(n18871), .B(n18870), .Z(n18936) );
  XNOR U19312 ( .A(sreg[492]), .B(n18936), .Z(n18938) );
  NANDN U19313 ( .A(sreg[491]), .B(n18863), .Z(n18867) );
  NAND U19314 ( .A(n18865), .B(n18864), .Z(n18866) );
  NAND U19315 ( .A(n18867), .B(n18866), .Z(n18937) );
  XNOR U19316 ( .A(n18938), .B(n18937), .Z(c[492]) );
  NANDN U19317 ( .A(n18869), .B(n18868), .Z(n18873) );
  NANDN U19318 ( .A(n18871), .B(n18870), .Z(n18872) );
  AND U19319 ( .A(n18873), .B(n18872), .Z(n18944) );
  NANDN U19320 ( .A(n18879), .B(n18878), .Z(n18883) );
  NANDN U19321 ( .A(n18881), .B(n18880), .Z(n18882) );
  NAND U19322 ( .A(n18883), .B(n18882), .Z(n18977) );
  NAND U19323 ( .A(b[0]), .B(a[253]), .Z(n18884) );
  XNOR U19324 ( .A(b[1]), .B(n18884), .Z(n18886) );
  NANDN U19325 ( .A(b[0]), .B(a[252]), .Z(n18885) );
  NAND U19326 ( .A(n18886), .B(n18885), .Z(n18956) );
  NAND U19327 ( .A(n19808), .B(n18887), .Z(n18889) );
  XOR U19328 ( .A(b[13]), .B(a[241]), .Z(n18959) );
  NAND U19329 ( .A(n19768), .B(n18959), .Z(n18888) );
  NAND U19330 ( .A(n18889), .B(n18888), .Z(n18954) );
  AND U19331 ( .A(b[15]), .B(a[237]), .Z(n18953) );
  XNOR U19332 ( .A(n18956), .B(n18955), .Z(n18975) );
  NAND U19333 ( .A(n33), .B(n18890), .Z(n18892) );
  XOR U19334 ( .A(a[249]), .B(b[5]), .Z(n18965) );
  NAND U19335 ( .A(n19342), .B(n18965), .Z(n18891) );
  NAND U19336 ( .A(n18892), .B(n18891), .Z(n18998) );
  NAND U19337 ( .A(n34), .B(n18893), .Z(n18895) );
  XOR U19338 ( .A(b[7]), .B(a[247]), .Z(n18968) );
  NAND U19339 ( .A(n19486), .B(n18968), .Z(n18894) );
  NAND U19340 ( .A(n18895), .B(n18894), .Z(n18996) );
  NAND U19341 ( .A(n31), .B(n18896), .Z(n18898) );
  XOR U19342 ( .A(a[251]), .B(b[3]), .Z(n18971) );
  NAND U19343 ( .A(n32), .B(n18971), .Z(n18897) );
  NAND U19344 ( .A(n18898), .B(n18897), .Z(n18995) );
  XOR U19345 ( .A(n18975), .B(n18974), .Z(n18976) );
  XOR U19346 ( .A(n18947), .B(n18948), .Z(n18950) );
  NAND U19347 ( .A(n18903), .B(n19724), .Z(n18905) );
  XOR U19348 ( .A(b[11]), .B(a[243]), .Z(n18980) );
  NAND U19349 ( .A(n19692), .B(n18980), .Z(n18904) );
  NAND U19350 ( .A(n18905), .B(n18904), .Z(n18992) );
  NAND U19351 ( .A(n19838), .B(n18906), .Z(n18908) );
  XOR U19352 ( .A(b[15]), .B(a[239]), .Z(n18983) );
  NAND U19353 ( .A(n19805), .B(n18983), .Z(n18907) );
  NAND U19354 ( .A(n18908), .B(n18907), .Z(n18990) );
  NAND U19355 ( .A(n35), .B(n18909), .Z(n18911) );
  XOR U19356 ( .A(b[9]), .B(a[245]), .Z(n18986) );
  NAND U19357 ( .A(n19598), .B(n18986), .Z(n18910) );
  NAND U19358 ( .A(n18911), .B(n18910), .Z(n18989) );
  NANDN U19359 ( .A(n18913), .B(n18912), .Z(n18917) );
  NANDN U19360 ( .A(n18915), .B(n18914), .Z(n18916) );
  AND U19361 ( .A(n18917), .B(n18916), .Z(n19002) );
  XOR U19362 ( .A(n19001), .B(n19002), .Z(n19003) );
  NAND U19363 ( .A(n18919), .B(n18918), .Z(n18923) );
  NAND U19364 ( .A(n18921), .B(n18920), .Z(n18922) );
  AND U19365 ( .A(n18923), .B(n18922), .Z(n19004) );
  XOR U19366 ( .A(n18950), .B(n18949), .Z(n19008) );
  NAND U19367 ( .A(n18925), .B(n18924), .Z(n18929) );
  NANDN U19368 ( .A(n18927), .B(n18926), .Z(n18928) );
  AND U19369 ( .A(n18929), .B(n18928), .Z(n19007) );
  XNOR U19370 ( .A(n19008), .B(n19007), .Z(n19009) );
  XOR U19371 ( .A(n19010), .B(n19009), .Z(n18942) );
  NANDN U19372 ( .A(n18931), .B(n18930), .Z(n18935) );
  NAND U19373 ( .A(n18933), .B(n18932), .Z(n18934) );
  AND U19374 ( .A(n18935), .B(n18934), .Z(n18941) );
  XNOR U19375 ( .A(n18942), .B(n18941), .Z(n18943) );
  XNOR U19376 ( .A(n18944), .B(n18943), .Z(n19013) );
  XNOR U19377 ( .A(sreg[493]), .B(n19013), .Z(n19015) );
  NANDN U19378 ( .A(sreg[492]), .B(n18936), .Z(n18940) );
  NAND U19379 ( .A(n18938), .B(n18937), .Z(n18939) );
  NAND U19380 ( .A(n18940), .B(n18939), .Z(n19014) );
  XNOR U19381 ( .A(n19015), .B(n19014), .Z(c[493]) );
  NANDN U19382 ( .A(n18942), .B(n18941), .Z(n18946) );
  NANDN U19383 ( .A(n18944), .B(n18943), .Z(n18945) );
  AND U19384 ( .A(n18946), .B(n18945), .Z(n19021) );
  NAND U19385 ( .A(n18948), .B(n18947), .Z(n18952) );
  NAND U19386 ( .A(n18950), .B(n18949), .Z(n18951) );
  AND U19387 ( .A(n18952), .B(n18951), .Z(n19087) );
  NAND U19388 ( .A(n18954), .B(n18953), .Z(n18958) );
  NANDN U19389 ( .A(n18956), .B(n18955), .Z(n18957) );
  NAND U19390 ( .A(n18958), .B(n18957), .Z(n19054) );
  NAND U19391 ( .A(n19808), .B(n18959), .Z(n18961) );
  XOR U19392 ( .A(b[13]), .B(a[242]), .Z(n19039) );
  NAND U19393 ( .A(n19768), .B(n19039), .Z(n18960) );
  NAND U19394 ( .A(n18961), .B(n18960), .Z(n19031) );
  AND U19395 ( .A(b[15]), .B(a[238]), .Z(n19030) );
  NAND U19396 ( .A(b[0]), .B(a[254]), .Z(n18962) );
  XNOR U19397 ( .A(b[1]), .B(n18962), .Z(n18964) );
  NANDN U19398 ( .A(b[0]), .B(a[253]), .Z(n18963) );
  NAND U19399 ( .A(n18964), .B(n18963), .Z(n19033) );
  XNOR U19400 ( .A(n19032), .B(n19033), .Z(n19052) );
  NAND U19401 ( .A(n33), .B(n18965), .Z(n18967) );
  XOR U19402 ( .A(a[250]), .B(b[5]), .Z(n19042) );
  NAND U19403 ( .A(n19342), .B(n19042), .Z(n18966) );
  NAND U19404 ( .A(n18967), .B(n18966), .Z(n19075) );
  NAND U19405 ( .A(n34), .B(n18968), .Z(n18970) );
  XOR U19406 ( .A(b[7]), .B(a[248]), .Z(n19045) );
  NAND U19407 ( .A(n19486), .B(n19045), .Z(n18969) );
  NAND U19408 ( .A(n18970), .B(n18969), .Z(n19073) );
  NAND U19409 ( .A(n31), .B(n18971), .Z(n18973) );
  XOR U19410 ( .A(a[252]), .B(b[3]), .Z(n19048) );
  NAND U19411 ( .A(n32), .B(n19048), .Z(n18972) );
  NAND U19412 ( .A(n18973), .B(n18972), .Z(n19072) );
  XOR U19413 ( .A(n19052), .B(n19051), .Z(n19053) );
  NAND U19414 ( .A(n18975), .B(n18974), .Z(n18979) );
  NAND U19415 ( .A(n18977), .B(n18976), .Z(n18978) );
  AND U19416 ( .A(n18979), .B(n18978), .Z(n19025) );
  XOR U19417 ( .A(n19024), .B(n19025), .Z(n19027) );
  NAND U19418 ( .A(n18980), .B(n19724), .Z(n18982) );
  XOR U19419 ( .A(b[11]), .B(a[244]), .Z(n19057) );
  NAND U19420 ( .A(n19692), .B(n19057), .Z(n18981) );
  NAND U19421 ( .A(n18982), .B(n18981), .Z(n19069) );
  NAND U19422 ( .A(n19838), .B(n18983), .Z(n18985) );
  XOR U19423 ( .A(b[15]), .B(a[240]), .Z(n19060) );
  NAND U19424 ( .A(n19805), .B(n19060), .Z(n18984) );
  NAND U19425 ( .A(n18985), .B(n18984), .Z(n19067) );
  NAND U19426 ( .A(n35), .B(n18986), .Z(n18988) );
  XOR U19427 ( .A(b[9]), .B(a[246]), .Z(n19063) );
  NAND U19428 ( .A(n19598), .B(n19063), .Z(n18987) );
  NAND U19429 ( .A(n18988), .B(n18987), .Z(n19066) );
  NAND U19430 ( .A(n18990), .B(n18989), .Z(n18994) );
  NAND U19431 ( .A(n18992), .B(n18991), .Z(n18993) );
  AND U19432 ( .A(n18994), .B(n18993), .Z(n19079) );
  XOR U19433 ( .A(n19078), .B(n19079), .Z(n19080) );
  NAND U19434 ( .A(n18996), .B(n18995), .Z(n19000) );
  NAND U19435 ( .A(n18998), .B(n18997), .Z(n18999) );
  AND U19436 ( .A(n19000), .B(n18999), .Z(n19081) );
  XNOR U19437 ( .A(n19027), .B(n19026), .Z(n19085) );
  NAND U19438 ( .A(n19002), .B(n19001), .Z(n19006) );
  NAND U19439 ( .A(n19004), .B(n19003), .Z(n19005) );
  AND U19440 ( .A(n19006), .B(n19005), .Z(n19084) );
  XOR U19441 ( .A(n19087), .B(n19086), .Z(n19019) );
  NANDN U19442 ( .A(n19008), .B(n19007), .Z(n19012) );
  NAND U19443 ( .A(n19010), .B(n19009), .Z(n19011) );
  AND U19444 ( .A(n19012), .B(n19011), .Z(n19018) );
  XNOR U19445 ( .A(n19019), .B(n19018), .Z(n19020) );
  XNOR U19446 ( .A(n19021), .B(n19020), .Z(n19090) );
  XNOR U19447 ( .A(sreg[494]), .B(n19090), .Z(n19092) );
  NANDN U19448 ( .A(sreg[493]), .B(n19013), .Z(n19017) );
  NAND U19449 ( .A(n19015), .B(n19014), .Z(n19016) );
  NAND U19450 ( .A(n19017), .B(n19016), .Z(n19091) );
  XNOR U19451 ( .A(n19092), .B(n19091), .Z(c[494]) );
  NANDN U19452 ( .A(n19019), .B(n19018), .Z(n19023) );
  NANDN U19453 ( .A(n19021), .B(n19020), .Z(n19022) );
  NAND U19454 ( .A(n19023), .B(n19022), .Z(n19103) );
  NAND U19455 ( .A(n19025), .B(n19024), .Z(n19029) );
  NAND U19456 ( .A(n19027), .B(n19026), .Z(n19028) );
  AND U19457 ( .A(n19029), .B(n19028), .Z(n19166) );
  NAND U19458 ( .A(n19031), .B(n19030), .Z(n19035) );
  NANDN U19459 ( .A(n19033), .B(n19032), .Z(n19034) );
  NAND U19460 ( .A(n19035), .B(n19034), .Z(n19133) );
  NAND U19461 ( .A(b[0]), .B(a[255]), .Z(n19036) );
  XNOR U19462 ( .A(b[1]), .B(n19036), .Z(n19038) );
  NANDN U19463 ( .A(b[0]), .B(a[254]), .Z(n19037) );
  NAND U19464 ( .A(n19038), .B(n19037), .Z(n19115) );
  NAND U19465 ( .A(n19808), .B(n19039), .Z(n19041) );
  XOR U19466 ( .A(b[13]), .B(a[243]), .Z(n19118) );
  NAND U19467 ( .A(n19768), .B(n19118), .Z(n19040) );
  NAND U19468 ( .A(n19041), .B(n19040), .Z(n19113) );
  AND U19469 ( .A(b[15]), .B(a[239]), .Z(n19112) );
  XNOR U19470 ( .A(n19115), .B(n19114), .Z(n19131) );
  NAND U19471 ( .A(n33), .B(n19042), .Z(n19044) );
  XOR U19472 ( .A(a[251]), .B(b[5]), .Z(n19121) );
  NAND U19473 ( .A(n19342), .B(n19121), .Z(n19043) );
  NAND U19474 ( .A(n19044), .B(n19043), .Z(n19154) );
  NAND U19475 ( .A(n34), .B(n19045), .Z(n19047) );
  XOR U19476 ( .A(b[7]), .B(a[249]), .Z(n19124) );
  NAND U19477 ( .A(n19486), .B(n19124), .Z(n19046) );
  NAND U19478 ( .A(n19047), .B(n19046), .Z(n19152) );
  NAND U19479 ( .A(n31), .B(n19048), .Z(n19050) );
  XOR U19480 ( .A(a[253]), .B(b[3]), .Z(n19127) );
  NAND U19481 ( .A(n32), .B(n19127), .Z(n19049) );
  NAND U19482 ( .A(n19050), .B(n19049), .Z(n19151) );
  XOR U19483 ( .A(n19131), .B(n19130), .Z(n19132) );
  NAND U19484 ( .A(n19052), .B(n19051), .Z(n19056) );
  NAND U19485 ( .A(n19054), .B(n19053), .Z(n19055) );
  AND U19486 ( .A(n19056), .B(n19055), .Z(n19107) );
  XOR U19487 ( .A(n19106), .B(n19107), .Z(n19109) );
  NAND U19488 ( .A(n19057), .B(n19724), .Z(n19059) );
  XOR U19489 ( .A(b[11]), .B(a[245]), .Z(n19136) );
  NAND U19490 ( .A(n19692), .B(n19136), .Z(n19058) );
  NAND U19491 ( .A(n19059), .B(n19058), .Z(n19148) );
  NAND U19492 ( .A(n19838), .B(n19060), .Z(n19062) );
  XOR U19493 ( .A(b[15]), .B(a[241]), .Z(n19139) );
  NAND U19494 ( .A(n19805), .B(n19139), .Z(n19061) );
  NAND U19495 ( .A(n19062), .B(n19061), .Z(n19146) );
  NAND U19496 ( .A(n35), .B(n19063), .Z(n19065) );
  XOR U19497 ( .A(b[9]), .B(a[247]), .Z(n19142) );
  NAND U19498 ( .A(n19598), .B(n19142), .Z(n19064) );
  NAND U19499 ( .A(n19065), .B(n19064), .Z(n19145) );
  NAND U19500 ( .A(n19067), .B(n19066), .Z(n19071) );
  NAND U19501 ( .A(n19069), .B(n19068), .Z(n19070) );
  AND U19502 ( .A(n19071), .B(n19070), .Z(n19158) );
  XOR U19503 ( .A(n19157), .B(n19158), .Z(n19159) );
  NAND U19504 ( .A(n19073), .B(n19072), .Z(n19077) );
  NAND U19505 ( .A(n19075), .B(n19074), .Z(n19076) );
  AND U19506 ( .A(n19077), .B(n19076), .Z(n19160) );
  XNOR U19507 ( .A(n19109), .B(n19108), .Z(n19164) );
  NAND U19508 ( .A(n19079), .B(n19078), .Z(n19083) );
  NAND U19509 ( .A(n19081), .B(n19080), .Z(n19082) );
  AND U19510 ( .A(n19083), .B(n19082), .Z(n19163) );
  XNOR U19511 ( .A(n19166), .B(n19165), .Z(n19101) );
  NAND U19512 ( .A(n19085), .B(n19084), .Z(n19089) );
  NAND U19513 ( .A(n19087), .B(n19086), .Z(n19088) );
  AND U19514 ( .A(n19089), .B(n19088), .Z(n19100) );
  XNOR U19515 ( .A(sreg[495]), .B(n19095), .Z(n19097) );
  NANDN U19516 ( .A(sreg[494]), .B(n19090), .Z(n19094) );
  NAND U19517 ( .A(n19092), .B(n19091), .Z(n19093) );
  NAND U19518 ( .A(n19094), .B(n19093), .Z(n19096) );
  XNOR U19519 ( .A(n19097), .B(n19096), .Z(c[495]) );
  NANDN U19520 ( .A(sreg[495]), .B(n19095), .Z(n19099) );
  NAND U19521 ( .A(n19097), .B(n19096), .Z(n19098) );
  AND U19522 ( .A(n19099), .B(n19098), .Z(n19170) );
  NAND U19523 ( .A(n19101), .B(n19100), .Z(n19105) );
  NAND U19524 ( .A(n19103), .B(n19102), .Z(n19104) );
  AND U19525 ( .A(n19105), .B(n19104), .Z(n19174) );
  NAND U19526 ( .A(n19107), .B(n19106), .Z(n19111) );
  NAND U19527 ( .A(n19109), .B(n19108), .Z(n19110) );
  AND U19528 ( .A(n19111), .B(n19110), .Z(n19237) );
  NAND U19529 ( .A(n19113), .B(n19112), .Z(n19117) );
  NANDN U19530 ( .A(n19115), .B(n19114), .Z(n19116) );
  NAND U19531 ( .A(n19117), .B(n19116), .Z(n19225) );
  NAND U19532 ( .A(n19808), .B(n19118), .Z(n19120) );
  XOR U19533 ( .A(b[13]), .B(a[244]), .Z(n19213) );
  NAND U19534 ( .A(n19768), .B(n19213), .Z(n19119) );
  NAND U19535 ( .A(n19120), .B(n19119), .Z(n19207) );
  AND U19536 ( .A(b[15]), .B(a[240]), .Z(n19204) );
  NAND U19537 ( .A(n33), .B(n19121), .Z(n19123) );
  XOR U19538 ( .A(a[252]), .B(b[5]), .Z(n19219) );
  NAND U19539 ( .A(n19342), .B(n19219), .Z(n19122) );
  NAND U19540 ( .A(n19123), .B(n19122), .Z(n19201) );
  NAND U19541 ( .A(n34), .B(n19124), .Z(n19126) );
  XOR U19542 ( .A(a[250]), .B(b[7]), .Z(n19189) );
  NAND U19543 ( .A(n19486), .B(n19189), .Z(n19125) );
  NAND U19544 ( .A(n19126), .B(n19125), .Z(n19199) );
  NAND U19545 ( .A(n31), .B(n19127), .Z(n19129) );
  XOR U19546 ( .A(a[254]), .B(b[3]), .Z(n19216) );
  NAND U19547 ( .A(n32), .B(n19216), .Z(n19128) );
  NAND U19548 ( .A(n19129), .B(n19128), .Z(n19198) );
  XOR U19549 ( .A(n19223), .B(n19222), .Z(n19224) );
  NAND U19550 ( .A(n19131), .B(n19130), .Z(n19135) );
  NAND U19551 ( .A(n19133), .B(n19132), .Z(n19134) );
  AND U19552 ( .A(n19135), .B(n19134), .Z(n19178) );
  XOR U19553 ( .A(n19177), .B(n19178), .Z(n19180) );
  NAND U19554 ( .A(n19136), .B(n19724), .Z(n19138) );
  XOR U19555 ( .A(b[11]), .B(a[246]), .Z(n19186) );
  NAND U19556 ( .A(n19692), .B(n19186), .Z(n19137) );
  NAND U19557 ( .A(n19138), .B(n19137), .Z(n19195) );
  NAND U19558 ( .A(n19838), .B(n19139), .Z(n19141) );
  XOR U19559 ( .A(b[15]), .B(a[242]), .Z(n19210) );
  NAND U19560 ( .A(n19805), .B(n19210), .Z(n19140) );
  NAND U19561 ( .A(n19141), .B(n19140), .Z(n19193) );
  NAND U19562 ( .A(n35), .B(n19142), .Z(n19144) );
  XOR U19563 ( .A(b[9]), .B(a[248]), .Z(n19183) );
  NAND U19564 ( .A(n19598), .B(n19183), .Z(n19143) );
  NAND U19565 ( .A(n19144), .B(n19143), .Z(n19192) );
  NAND U19566 ( .A(n19146), .B(n19145), .Z(n19150) );
  NAND U19567 ( .A(n19148), .B(n19147), .Z(n19149) );
  AND U19568 ( .A(n19150), .B(n19149), .Z(n19229) );
  XOR U19569 ( .A(n19228), .B(n19229), .Z(n19230) );
  NAND U19570 ( .A(n19152), .B(n19151), .Z(n19156) );
  NAND U19571 ( .A(n19154), .B(n19153), .Z(n19155) );
  AND U19572 ( .A(n19156), .B(n19155), .Z(n19231) );
  XNOR U19573 ( .A(n19180), .B(n19179), .Z(n19235) );
  NAND U19574 ( .A(n19158), .B(n19157), .Z(n19162) );
  NAND U19575 ( .A(n19160), .B(n19159), .Z(n19161) );
  AND U19576 ( .A(n19162), .B(n19161), .Z(n19234) );
  XNOR U19577 ( .A(n19237), .B(n19236), .Z(n19172) );
  NAND U19578 ( .A(n19164), .B(n19163), .Z(n19168) );
  NAND U19579 ( .A(n19166), .B(n19165), .Z(n19167) );
  AND U19580 ( .A(n19168), .B(n19167), .Z(n19171) );
  XOR U19581 ( .A(n19174), .B(n19173), .Z(n19169) );
  XOR U19582 ( .A(n19170), .B(n19169), .Z(c[496]) );
  AND U19583 ( .A(n19170), .B(n19169), .Z(n19241) );
  NAND U19584 ( .A(n19172), .B(n19171), .Z(n19176) );
  NANDN U19585 ( .A(n19174), .B(n19173), .Z(n19175) );
  AND U19586 ( .A(n19176), .B(n19175), .Z(n19245) );
  NAND U19587 ( .A(n19178), .B(n19177), .Z(n19182) );
  NAND U19588 ( .A(n19180), .B(n19179), .Z(n19181) );
  AND U19589 ( .A(n19182), .B(n19181), .Z(n19306) );
  NAND U19590 ( .A(n35), .B(n19183), .Z(n19185) );
  XOR U19591 ( .A(b[9]), .B(a[249]), .Z(n19272) );
  NAND U19592 ( .A(n19598), .B(n19272), .Z(n19184) );
  NAND U19593 ( .A(n19185), .B(n19184), .Z(n19278) );
  NAND U19594 ( .A(n19186), .B(n19724), .Z(n19188) );
  XOR U19595 ( .A(b[11]), .B(a[247]), .Z(n19260) );
  NAND U19596 ( .A(n19692), .B(n19260), .Z(n19187) );
  NAND U19597 ( .A(n19188), .B(n19187), .Z(n19276) );
  NAND U19598 ( .A(n34), .B(n19189), .Z(n19191) );
  XOR U19599 ( .A(a[251]), .B(b[7]), .Z(n19266) );
  NAND U19600 ( .A(n19486), .B(n19266), .Z(n19190) );
  NAND U19601 ( .A(n19191), .B(n19190), .Z(n19275) );
  NAND U19602 ( .A(n19193), .B(n19192), .Z(n19197) );
  NAND U19603 ( .A(n19195), .B(n19194), .Z(n19196) );
  AND U19604 ( .A(n19197), .B(n19196), .Z(n19298) );
  XOR U19605 ( .A(n19297), .B(n19298), .Z(n19299) );
  NAND U19606 ( .A(n19199), .B(n19198), .Z(n19203) );
  NAND U19607 ( .A(n19201), .B(n19200), .Z(n19202) );
  AND U19608 ( .A(n19203), .B(n19202), .Z(n19300) );
  NAND U19609 ( .A(n19205), .B(n19204), .Z(n19209) );
  NAND U19610 ( .A(n19207), .B(n19206), .Z(n19208) );
  NAND U19611 ( .A(n19209), .B(n19208), .Z(n19294) );
  NAND U19612 ( .A(n19838), .B(n19210), .Z(n19212) );
  XOR U19613 ( .A(b[15]), .B(a[243]), .Z(n19257) );
  NAND U19614 ( .A(n19805), .B(n19257), .Z(n19211) );
  NAND U19615 ( .A(n19212), .B(n19211), .Z(n19288) );
  AND U19616 ( .A(b[15]), .B(a[241]), .Z(n19408) );
  NAND U19617 ( .A(n19808), .B(n19213), .Z(n19215) );
  XOR U19618 ( .A(b[13]), .B(a[245]), .Z(n19263) );
  NAND U19619 ( .A(n19768), .B(n19263), .Z(n19214) );
  NAND U19620 ( .A(n19215), .B(n19214), .Z(n19286) );
  XNOR U19621 ( .A(n19408), .B(n19286), .Z(n19287) );
  NAND U19622 ( .A(n31), .B(n19216), .Z(n19218) );
  XOR U19623 ( .A(a[255]), .B(b[3]), .Z(n19254) );
  NAND U19624 ( .A(n32), .B(n19254), .Z(n19217) );
  NAND U19625 ( .A(n19218), .B(n19217), .Z(n19283) );
  NAND U19626 ( .A(n33), .B(n19219), .Z(n19221) );
  XOR U19627 ( .A(a[253]), .B(b[5]), .Z(n19269) );
  NAND U19628 ( .A(n19342), .B(n19269), .Z(n19220) );
  NAND U19629 ( .A(n19221), .B(n19220), .Z(n19281) );
  XNOR U19630 ( .A(b[1]), .B(n19281), .Z(n19282) );
  XOR U19631 ( .A(n19292), .B(n19291), .Z(n19293) );
  NAND U19632 ( .A(n19223), .B(n19222), .Z(n19227) );
  NAND U19633 ( .A(n19225), .B(n19224), .Z(n19226) );
  AND U19634 ( .A(n19227), .B(n19226), .Z(n19249) );
  XOR U19635 ( .A(n19248), .B(n19249), .Z(n19250) );
  XNOR U19636 ( .A(n19251), .B(n19250), .Z(n19304) );
  NAND U19637 ( .A(n19229), .B(n19228), .Z(n19233) );
  NAND U19638 ( .A(n19231), .B(n19230), .Z(n19232) );
  AND U19639 ( .A(n19233), .B(n19232), .Z(n19303) );
  XNOR U19640 ( .A(n19306), .B(n19305), .Z(n19243) );
  NAND U19641 ( .A(n19235), .B(n19234), .Z(n19239) );
  NAND U19642 ( .A(n19237), .B(n19236), .Z(n19238) );
  AND U19643 ( .A(n19239), .B(n19238), .Z(n19242) );
  XOR U19644 ( .A(n19245), .B(n19244), .Z(n19240) );
  XOR U19645 ( .A(n19241), .B(n19240), .Z(c[497]) );
  AND U19646 ( .A(n19241), .B(n19240), .Z(n19310) );
  NAND U19647 ( .A(n19243), .B(n19242), .Z(n19247) );
  NANDN U19648 ( .A(n19245), .B(n19244), .Z(n19246) );
  AND U19649 ( .A(n19247), .B(n19246), .Z(n19314) );
  NAND U19650 ( .A(n19249), .B(n19248), .Z(n19253) );
  NAND U19651 ( .A(n19251), .B(n19250), .Z(n19252) );
  AND U19652 ( .A(n19253), .B(n19252), .Z(n19376) );
  NAND U19653 ( .A(n32), .B(b[3]), .Z(n19256) );
  NANDN U19654 ( .A(n29), .B(n19254), .Z(n19255) );
  AND U19655 ( .A(n19256), .B(n19255), .Z(n19361) );
  NAND U19656 ( .A(b[15]), .B(a[242]), .Z(n19362) );
  XOR U19657 ( .A(n19361), .B(n19362), .Z(n19363) );
  XNOR U19658 ( .A(n19408), .B(n19363), .Z(n19358) );
  NAND U19659 ( .A(n19838), .B(n19257), .Z(n19259) );
  XOR U19660 ( .A(b[15]), .B(a[244]), .Z(n19329) );
  NAND U19661 ( .A(n19805), .B(n19329), .Z(n19258) );
  NAND U19662 ( .A(n19259), .B(n19258), .Z(n19356) );
  NAND U19663 ( .A(n19260), .B(n19724), .Z(n19262) );
  XOR U19664 ( .A(b[11]), .B(a[248]), .Z(n19345) );
  NAND U19665 ( .A(n19692), .B(n19345), .Z(n19261) );
  NAND U19666 ( .A(n19262), .B(n19261), .Z(n19355) );
  XOR U19667 ( .A(n19358), .B(n19357), .Z(n19326) );
  NAND U19668 ( .A(n19808), .B(n19263), .Z(n19265) );
  XOR U19669 ( .A(b[13]), .B(a[246]), .Z(n19338) );
  NAND U19670 ( .A(n19768), .B(n19338), .Z(n19264) );
  NAND U19671 ( .A(n19265), .B(n19264), .Z(n19324) );
  NAND U19672 ( .A(n34), .B(n19266), .Z(n19268) );
  XOR U19673 ( .A(a[252]), .B(b[7]), .Z(n19335) );
  NAND U19674 ( .A(n19486), .B(n19335), .Z(n19267) );
  NAND U19675 ( .A(n19268), .B(n19267), .Z(n19352) );
  NAND U19676 ( .A(n33), .B(n19269), .Z(n19271) );
  XOR U19677 ( .A(a[254]), .B(b[5]), .Z(n19341) );
  NAND U19678 ( .A(n19342), .B(n19341), .Z(n19270) );
  NAND U19679 ( .A(n19271), .B(n19270), .Z(n19350) );
  NAND U19680 ( .A(n35), .B(n19272), .Z(n19274) );
  XOR U19681 ( .A(b[9]), .B(a[250]), .Z(n19332) );
  NAND U19682 ( .A(n19598), .B(n19332), .Z(n19273) );
  NAND U19683 ( .A(n19274), .B(n19273), .Z(n19349) );
  XOR U19684 ( .A(n19326), .B(n19325), .Z(n19320) );
  NAND U19685 ( .A(n19276), .B(n19275), .Z(n19280) );
  NAND U19686 ( .A(n19278), .B(n19277), .Z(n19279) );
  NAND U19687 ( .A(n19280), .B(n19279), .Z(n19318) );
  NANDN U19688 ( .A(b[1]), .B(n19281), .Z(n19285) );
  NAND U19689 ( .A(n19283), .B(n19282), .Z(n19284) );
  NAND U19690 ( .A(n19285), .B(n19284), .Z(n19317) );
  XNOR U19691 ( .A(n19320), .B(n19319), .Z(n19370) );
  IV U19692 ( .A(n19408), .Z(n19364) );
  NAND U19693 ( .A(n19364), .B(n19286), .Z(n19290) );
  NAND U19694 ( .A(n19288), .B(n19287), .Z(n19289) );
  AND U19695 ( .A(n19290), .B(n19289), .Z(n19367) );
  NAND U19696 ( .A(n19292), .B(n19291), .Z(n19296) );
  NAND U19697 ( .A(n19294), .B(n19293), .Z(n19295) );
  AND U19698 ( .A(n19296), .B(n19295), .Z(n19368) );
  NAND U19699 ( .A(n19298), .B(n19297), .Z(n19302) );
  NAND U19700 ( .A(n19300), .B(n19299), .Z(n19301) );
  AND U19701 ( .A(n19302), .B(n19301), .Z(n19374) );
  XOR U19702 ( .A(n19373), .B(n19374), .Z(n19375) );
  XNOR U19703 ( .A(n19376), .B(n19375), .Z(n19312) );
  NAND U19704 ( .A(n19304), .B(n19303), .Z(n19308) );
  NAND U19705 ( .A(n19306), .B(n19305), .Z(n19307) );
  AND U19706 ( .A(n19308), .B(n19307), .Z(n19311) );
  XOR U19707 ( .A(n19314), .B(n19313), .Z(n19309) );
  XOR U19708 ( .A(n19310), .B(n19309), .Z(c[498]) );
  AND U19709 ( .A(n19310), .B(n19309), .Z(n19380) );
  NAND U19710 ( .A(n19312), .B(n19311), .Z(n19316) );
  NANDN U19711 ( .A(n19314), .B(n19313), .Z(n19315) );
  AND U19712 ( .A(n19316), .B(n19315), .Z(n19384) );
  NAND U19713 ( .A(n19318), .B(n19317), .Z(n19322) );
  NAND U19714 ( .A(n19320), .B(n19319), .Z(n19321) );
  NAND U19715 ( .A(n19322), .B(n19321), .Z(n19388) );
  NAND U19716 ( .A(n19324), .B(n19323), .Z(n19328) );
  NAND U19717 ( .A(n19326), .B(n19325), .Z(n19327) );
  NAND U19718 ( .A(n19328), .B(n19327), .Z(n19394) );
  NAND U19719 ( .A(n19838), .B(n19329), .Z(n19331) );
  XOR U19720 ( .A(b[15]), .B(a[245]), .Z(n19417) );
  NAND U19721 ( .A(n19805), .B(n19417), .Z(n19330) );
  NAND U19722 ( .A(n19331), .B(n19330), .Z(n19436) );
  NAND U19723 ( .A(n35), .B(n19332), .Z(n19334) );
  XOR U19724 ( .A(b[9]), .B(a[251]), .Z(n19424) );
  NAND U19725 ( .A(n19598), .B(n19424), .Z(n19333) );
  NAND U19726 ( .A(n19334), .B(n19333), .Z(n19402) );
  NAND U19727 ( .A(n34), .B(n19335), .Z(n19337) );
  XOR U19728 ( .A(a[253]), .B(b[7]), .Z(n19427) );
  NAND U19729 ( .A(n19486), .B(n19427), .Z(n19336) );
  NAND U19730 ( .A(n19337), .B(n19336), .Z(n19400) );
  NAND U19731 ( .A(n19808), .B(n19338), .Z(n19340) );
  XOR U19732 ( .A(b[13]), .B(a[247]), .Z(n19433) );
  NAND U19733 ( .A(n19768), .B(n19433), .Z(n19339) );
  NAND U19734 ( .A(n19340), .B(n19339), .Z(n19399) );
  NAND U19735 ( .A(n33), .B(n19341), .Z(n19344) );
  XOR U19736 ( .A(a[255]), .B(b[5]), .Z(n19420) );
  NAND U19737 ( .A(n19342), .B(n19420), .Z(n19343) );
  NAND U19738 ( .A(n19344), .B(n19343), .Z(n19412) );
  NAND U19739 ( .A(n19345), .B(n19724), .Z(n19347) );
  XOR U19740 ( .A(b[11]), .B(a[249]), .Z(n19430) );
  NAND U19741 ( .A(n19692), .B(n19430), .Z(n19346) );
  NAND U19742 ( .A(n19347), .B(n19346), .Z(n19411) );
  AND U19743 ( .A(b[15]), .B(a[243]), .Z(n19405) );
  XNOR U19744 ( .A(n19348), .B(n19405), .Z(n19407) );
  XOR U19745 ( .A(n19408), .B(n19407), .Z(n19413) );
  XOR U19746 ( .A(n19414), .B(n19413), .Z(n19437) );
  XOR U19747 ( .A(n19438), .B(n19437), .Z(n19393) );
  NAND U19748 ( .A(n19350), .B(n19349), .Z(n19354) );
  NAND U19749 ( .A(n19352), .B(n19351), .Z(n19353) );
  NAND U19750 ( .A(n19354), .B(n19353), .Z(n19444) );
  NAND U19751 ( .A(n19356), .B(n19355), .Z(n19360) );
  NAND U19752 ( .A(n19358), .B(n19357), .Z(n19359) );
  NAND U19753 ( .A(n19360), .B(n19359), .Z(n19442) );
  OR U19754 ( .A(n19362), .B(n19361), .Z(n19366) );
  NAND U19755 ( .A(n19364), .B(n19363), .Z(n19365) );
  NAND U19756 ( .A(n19366), .B(n19365), .Z(n19441) );
  XOR U19757 ( .A(n19396), .B(n19395), .Z(n19387) );
  NAND U19758 ( .A(n19368), .B(n19367), .Z(n19372) );
  NAND U19759 ( .A(n19370), .B(n19369), .Z(n19371) );
  AND U19760 ( .A(n19372), .B(n19371), .Z(n19389) );
  XNOR U19761 ( .A(n19390), .B(n19389), .Z(n19382) );
  NAND U19762 ( .A(n19374), .B(n19373), .Z(n19378) );
  NAND U19763 ( .A(n19376), .B(n19375), .Z(n19377) );
  AND U19764 ( .A(n19378), .B(n19377), .Z(n19381) );
  XOR U19765 ( .A(n19384), .B(n19383), .Z(n19379) );
  XOR U19766 ( .A(n19380), .B(n19379), .Z(c[499]) );
  AND U19767 ( .A(n19380), .B(n19379), .Z(n19448) );
  NAND U19768 ( .A(n19382), .B(n19381), .Z(n19386) );
  NANDN U19769 ( .A(n19384), .B(n19383), .Z(n19385) );
  AND U19770 ( .A(n19386), .B(n19385), .Z(n19452) );
  NAND U19771 ( .A(n19388), .B(n19387), .Z(n19392) );
  NAND U19772 ( .A(n19390), .B(n19389), .Z(n19391) );
  AND U19773 ( .A(n19392), .B(n19391), .Z(n19450) );
  NAND U19774 ( .A(n19394), .B(n19393), .Z(n19398) );
  NAND U19775 ( .A(n19396), .B(n19395), .Z(n19397) );
  AND U19776 ( .A(n19398), .B(n19397), .Z(n19458) );
  NAND U19777 ( .A(n19400), .B(n19399), .Z(n19404) );
  NAND U19778 ( .A(n19402), .B(n19401), .Z(n19403) );
  AND U19779 ( .A(n19404), .B(n19403), .Z(n19470) );
  NAND U19780 ( .A(n19406), .B(n19405), .Z(n19410) );
  NAND U19781 ( .A(n19408), .B(n19407), .Z(n19409) );
  AND U19782 ( .A(n19410), .B(n19409), .Z(n19467) );
  NAND U19783 ( .A(n19412), .B(n19411), .Z(n19416) );
  NAND U19784 ( .A(n19414), .B(n19413), .Z(n19415) );
  AND U19785 ( .A(n19416), .B(n19415), .Z(n19468) );
  XNOR U19786 ( .A(n19470), .B(n19469), .Z(n19464) );
  NAND U19787 ( .A(n19838), .B(n19417), .Z(n19419) );
  XOR U19788 ( .A(b[15]), .B(a[246]), .Z(n19499) );
  NAND U19789 ( .A(n19805), .B(n19499), .Z(n19418) );
  NAND U19790 ( .A(n19419), .B(n19418), .Z(n19504) );
  AND U19791 ( .A(b[15]), .B(a[244]), .Z(n19554) );
  AND U19792 ( .A(n19420), .B(n33), .Z(n19423) );
  XOR U19793 ( .A(b[4]), .B(b[3]), .Z(n19421) );
  NAND U19794 ( .A(b[5]), .B(n19421), .Z(n19422) );
  NANDN U19795 ( .A(n19423), .B(n19422), .Z(n19502) );
  XNOR U19796 ( .A(n19554), .B(n19502), .Z(n19503) );
  NAND U19797 ( .A(n35), .B(n19424), .Z(n19426) );
  XOR U19798 ( .A(a[252]), .B(b[9]), .Z(n19493) );
  NAND U19799 ( .A(n19598), .B(n19493), .Z(n19425) );
  NAND U19800 ( .A(n19426), .B(n19425), .Z(n19482) );
  NAND U19801 ( .A(n34), .B(n19427), .Z(n19429) );
  XOR U19802 ( .A(a[254]), .B(b[7]), .Z(n19485) );
  NAND U19803 ( .A(n19486), .B(n19485), .Z(n19428) );
  NAND U19804 ( .A(n19429), .B(n19428), .Z(n19480) );
  NAND U19805 ( .A(n19430), .B(n19724), .Z(n19432) );
  XOR U19806 ( .A(b[11]), .B(a[250]), .Z(n19489) );
  NAND U19807 ( .A(n19692), .B(n19489), .Z(n19431) );
  NAND U19808 ( .A(n19432), .B(n19431), .Z(n19479) );
  XOR U19809 ( .A(b[13]), .B(a[248]), .Z(n19496) );
  XOR U19810 ( .A(n19473), .B(n19474), .Z(n19476) );
  XNOR U19811 ( .A(n19475), .B(n19476), .Z(n19462) );
  NAND U19812 ( .A(n19436), .B(n19435), .Z(n19440) );
  NAND U19813 ( .A(n19438), .B(n19437), .Z(n19439) );
  NAND U19814 ( .A(n19440), .B(n19439), .Z(n19461) );
  XOR U19815 ( .A(n19462), .B(n19461), .Z(n19463) );
  NAND U19816 ( .A(n19442), .B(n19441), .Z(n19446) );
  NAND U19817 ( .A(n19444), .B(n19443), .Z(n19445) );
  AND U19818 ( .A(n19446), .B(n19445), .Z(n19456) );
  XOR U19819 ( .A(n19455), .B(n19456), .Z(n19457) );
  XOR U19820 ( .A(n19458), .B(n19457), .Z(n19449) );
  XOR U19821 ( .A(n19450), .B(n19449), .Z(n19451) );
  XOR U19822 ( .A(n19452), .B(n19451), .Z(n19447) );
  XOR U19823 ( .A(n19448), .B(n19447), .Z(c[500]) );
  AND U19824 ( .A(n19448), .B(n19447), .Z(n19506) );
  NAND U19825 ( .A(n19450), .B(n19449), .Z(n19454) );
  NANDN U19826 ( .A(n19452), .B(n19451), .Z(n19453) );
  AND U19827 ( .A(n19454), .B(n19453), .Z(n19510) );
  NAND U19828 ( .A(n19456), .B(n19455), .Z(n19460) );
  NAND U19829 ( .A(n19458), .B(n19457), .Z(n19459) );
  NAND U19830 ( .A(n19460), .B(n19459), .Z(n19508) );
  NAND U19831 ( .A(n19462), .B(n19461), .Z(n19466) );
  NAND U19832 ( .A(n19464), .B(n19463), .Z(n19465) );
  AND U19833 ( .A(n19466), .B(n19465), .Z(n19516) );
  NAND U19834 ( .A(n19468), .B(n19467), .Z(n19472) );
  NAND U19835 ( .A(n19470), .B(n19469), .Z(n19471) );
  NAND U19836 ( .A(n19472), .B(n19471), .Z(n19514) );
  NAND U19837 ( .A(n19474), .B(n19473), .Z(n19478) );
  NAND U19838 ( .A(n19476), .B(n19475), .Z(n19477) );
  NAND U19839 ( .A(n19478), .B(n19477), .Z(n19522) );
  NAND U19840 ( .A(n19480), .B(n19479), .Z(n19484) );
  NAND U19841 ( .A(n19482), .B(n19481), .Z(n19483) );
  NAND U19842 ( .A(n19484), .B(n19483), .Z(n19562) );
  NAND U19843 ( .A(n34), .B(n19485), .Z(n19488) );
  XOR U19844 ( .A(a[255]), .B(b[7]), .Z(n19537) );
  NAND U19845 ( .A(n19486), .B(n19537), .Z(n19487) );
  NAND U19846 ( .A(n19488), .B(n19487), .Z(n19548) );
  NAND U19847 ( .A(n19489), .B(n19724), .Z(n19491) );
  XOR U19848 ( .A(b[11]), .B(a[251]), .Z(n19525) );
  NAND U19849 ( .A(n19692), .B(n19525), .Z(n19490) );
  NAND U19850 ( .A(n19491), .B(n19490), .Z(n19547) );
  XNOR U19851 ( .A(n19554), .B(n19492), .Z(n19556) );
  AND U19852 ( .A(b[15]), .B(a[245]), .Z(n19555) );
  XOR U19853 ( .A(n19556), .B(n19555), .Z(n19549) );
  XOR U19854 ( .A(n19550), .B(n19549), .Z(n19560) );
  NAND U19855 ( .A(n35), .B(n19493), .Z(n19495) );
  XOR U19856 ( .A(a[253]), .B(b[9]), .Z(n19528) );
  NAND U19857 ( .A(n19598), .B(n19528), .Z(n19494) );
  NAND U19858 ( .A(n19495), .B(n19494), .Z(n19544) );
  NAND U19859 ( .A(n19808), .B(n19496), .Z(n19498) );
  XOR U19860 ( .A(b[13]), .B(a[249]), .Z(n19531) );
  NAND U19861 ( .A(n19768), .B(n19531), .Z(n19497) );
  NAND U19862 ( .A(n19498), .B(n19497), .Z(n19542) );
  NAND U19863 ( .A(n19838), .B(n19499), .Z(n19501) );
  XOR U19864 ( .A(b[15]), .B(a[247]), .Z(n19534) );
  NAND U19865 ( .A(n19805), .B(n19534), .Z(n19500) );
  NAND U19866 ( .A(n19501), .B(n19500), .Z(n19541) );
  XOR U19867 ( .A(n19560), .B(n19559), .Z(n19561) );
  XOR U19868 ( .A(n19519), .B(n19520), .Z(n19521) );
  XOR U19869 ( .A(n19516), .B(n19515), .Z(n19507) );
  XOR U19870 ( .A(n19510), .B(n19509), .Z(n19505) );
  XOR U19871 ( .A(n19506), .B(n19505), .Z(c[501]) );
  AND U19872 ( .A(n19506), .B(n19505), .Z(n19566) );
  NAND U19873 ( .A(n19508), .B(n19507), .Z(n19512) );
  NANDN U19874 ( .A(n19510), .B(n19509), .Z(n19511) );
  AND U19875 ( .A(n19512), .B(n19511), .Z(n19570) );
  NAND U19876 ( .A(n19514), .B(n19513), .Z(n19518) );
  NAND U19877 ( .A(n19516), .B(n19515), .Z(n19517) );
  NAND U19878 ( .A(n19518), .B(n19517), .Z(n19568) );
  NAND U19879 ( .A(n19520), .B(n19519), .Z(n19524) );
  NAND U19880 ( .A(n19522), .B(n19521), .Z(n19523) );
  NAND U19881 ( .A(n19524), .B(n19523), .Z(n19576) );
  NAND U19882 ( .A(n19525), .B(n19724), .Z(n19527) );
  XOR U19883 ( .A(b[11]), .B(a[252]), .Z(n19594) );
  NAND U19884 ( .A(n19692), .B(n19594), .Z(n19526) );
  NAND U19885 ( .A(n19527), .B(n19526), .Z(n19585) );
  NAND U19886 ( .A(n35), .B(n19528), .Z(n19530) );
  XOR U19887 ( .A(a[254]), .B(b[9]), .Z(n19597) );
  NAND U19888 ( .A(n19598), .B(n19597), .Z(n19529) );
  NAND U19889 ( .A(n19530), .B(n19529), .Z(n19583) );
  NAND U19890 ( .A(n19808), .B(n19531), .Z(n19533) );
  XOR U19891 ( .A(b[13]), .B(a[250]), .Z(n19601) );
  NAND U19892 ( .A(n19768), .B(n19601), .Z(n19532) );
  NAND U19893 ( .A(n19533), .B(n19532), .Z(n19582) );
  NAND U19894 ( .A(n19838), .B(n19534), .Z(n19536) );
  XOR U19895 ( .A(b[15]), .B(a[248]), .Z(n19591) );
  NAND U19896 ( .A(n19805), .B(n19591), .Z(n19535) );
  AND U19897 ( .A(n19536), .B(n19535), .Z(n19590) );
  AND U19898 ( .A(b[15]), .B(a[246]), .Z(n19644) );
  AND U19899 ( .A(n19537), .B(n34), .Z(n19540) );
  XOR U19900 ( .A(b[6]), .B(b[5]), .Z(n19538) );
  NAND U19901 ( .A(b[7]), .B(n19538), .Z(n19539) );
  NANDN U19902 ( .A(n19540), .B(n19539), .Z(n19588) );
  XNOR U19903 ( .A(n19644), .B(n19588), .Z(n19589) );
  XOR U19904 ( .A(n19590), .B(n19589), .Z(n19604) );
  XOR U19905 ( .A(n19605), .B(n19604), .Z(n19607) );
  NAND U19906 ( .A(n19542), .B(n19541), .Z(n19546) );
  NAND U19907 ( .A(n19544), .B(n19543), .Z(n19545) );
  AND U19908 ( .A(n19546), .B(n19545), .Z(n19606) );
  XNOR U19909 ( .A(n19607), .B(n19606), .Z(n19581) );
  NAND U19910 ( .A(n19548), .B(n19547), .Z(n19552) );
  NAND U19911 ( .A(n19550), .B(n19549), .Z(n19551) );
  NAND U19912 ( .A(n19552), .B(n19551), .Z(n19580) );
  NAND U19913 ( .A(n19554), .B(n19553), .Z(n19558) );
  NAND U19914 ( .A(n19556), .B(n19555), .Z(n19557) );
  AND U19915 ( .A(n19558), .B(n19557), .Z(n19579) );
  NAND U19916 ( .A(n19560), .B(n19559), .Z(n19564) );
  NAND U19917 ( .A(n19562), .B(n19561), .Z(n19563) );
  AND U19918 ( .A(n19564), .B(n19563), .Z(n19574) );
  XOR U19919 ( .A(n19570), .B(n19569), .Z(n19565) );
  XOR U19920 ( .A(n19566), .B(n19565), .Z(c[502]) );
  AND U19921 ( .A(n19566), .B(n19565), .Z(n19611) );
  NAND U19922 ( .A(n19568), .B(n19567), .Z(n19572) );
  NANDN U19923 ( .A(n19570), .B(n19569), .Z(n19571) );
  AND U19924 ( .A(n19572), .B(n19571), .Z(n19615) );
  NAND U19925 ( .A(n19574), .B(n19573), .Z(n19578) );
  NAND U19926 ( .A(n19576), .B(n19575), .Z(n19577) );
  NAND U19927 ( .A(n19578), .B(n19577), .Z(n19613) );
  NAND U19928 ( .A(n19583), .B(n19582), .Z(n19587) );
  NAND U19929 ( .A(n19585), .B(n19584), .Z(n19586) );
  NAND U19930 ( .A(n19587), .B(n19586), .Z(n19627) );
  NAND U19931 ( .A(n19838), .B(n19591), .Z(n19593) );
  XOR U19932 ( .A(b[15]), .B(a[249]), .Z(n19636) );
  NAND U19933 ( .A(n19805), .B(n19636), .Z(n19592) );
  NAND U19934 ( .A(n19593), .B(n19592), .Z(n19659) );
  NAND U19935 ( .A(n19594), .B(n19724), .Z(n19596) );
  XOR U19936 ( .A(b[11]), .B(a[253]), .Z(n19653) );
  NAND U19937 ( .A(n19692), .B(n19653), .Z(n19595) );
  NAND U19938 ( .A(n19596), .B(n19595), .Z(n19657) );
  NAND U19939 ( .A(n35), .B(n19597), .Z(n19600) );
  XOR U19940 ( .A(a[255]), .B(b[9]), .Z(n19639) );
  NAND U19941 ( .A(n19598), .B(n19639), .Z(n19599) );
  NAND U19942 ( .A(n19600), .B(n19599), .Z(n19631) );
  NAND U19943 ( .A(n19808), .B(n19601), .Z(n19603) );
  XOR U19944 ( .A(b[13]), .B(a[251]), .Z(n19650) );
  NAND U19945 ( .A(n19768), .B(n19650), .Z(n19602) );
  NAND U19946 ( .A(n19603), .B(n19602), .Z(n19630) );
  AND U19947 ( .A(b[15]), .B(a[247]), .Z(n19647) );
  XOR U19948 ( .A(n19646), .B(n19647), .Z(n19645) );
  XOR U19949 ( .A(n19644), .B(n19645), .Z(n19632) );
  XOR U19950 ( .A(n19633), .B(n19632), .Z(n19656) );
  NAND U19951 ( .A(n19605), .B(n19604), .Z(n19609) );
  NAND U19952 ( .A(n19607), .B(n19606), .Z(n19608) );
  NAND U19953 ( .A(n19609), .B(n19608), .Z(n19618) );
  XOR U19954 ( .A(n19619), .B(n19618), .Z(n19620) );
  XNOR U19955 ( .A(n19621), .B(n19620), .Z(n19612) );
  XOR U19956 ( .A(n19615), .B(n19614), .Z(n19610) );
  XOR U19957 ( .A(n19611), .B(n19610), .Z(c[503]) );
  AND U19958 ( .A(n19611), .B(n19610), .Z(n19663) );
  NAND U19959 ( .A(n19613), .B(n19612), .Z(n19617) );
  NANDN U19960 ( .A(n19615), .B(n19614), .Z(n19616) );
  AND U19961 ( .A(n19617), .B(n19616), .Z(n19667) );
  NAND U19962 ( .A(n19619), .B(n19618), .Z(n19623) );
  NANDN U19963 ( .A(n19621), .B(n19620), .Z(n19622) );
  NAND U19964 ( .A(n19623), .B(n19622), .Z(n19665) );
  NAND U19965 ( .A(n19625), .B(n19624), .Z(n19629) );
  NAND U19966 ( .A(n19627), .B(n19626), .Z(n19628) );
  AND U19967 ( .A(n19629), .B(n19628), .Z(n19673) );
  NAND U19968 ( .A(n19631), .B(n19630), .Z(n19635) );
  NAND U19969 ( .A(n19633), .B(n19632), .Z(n19634) );
  NAND U19970 ( .A(n19635), .B(n19634), .Z(n19677) );
  NAND U19971 ( .A(n19838), .B(n19636), .Z(n19638) );
  XOR U19972 ( .A(b[15]), .B(a[250]), .Z(n19698) );
  NAND U19973 ( .A(n19805), .B(n19698), .Z(n19637) );
  NAND U19974 ( .A(n19638), .B(n19637), .Z(n19690) );
  IV U19975 ( .A(n19690), .Z(n19643) );
  AND U19976 ( .A(b[15]), .B(a[248]), .Z(n19732) );
  AND U19977 ( .A(n19639), .B(n35), .Z(n19642) );
  XOR U19978 ( .A(b[8]), .B(b[7]), .Z(n19640) );
  NAND U19979 ( .A(b[9]), .B(n19640), .Z(n19641) );
  NANDN U19980 ( .A(n19642), .B(n19641), .Z(n19688) );
  XNOR U19981 ( .A(n19732), .B(n19688), .Z(n19689) );
  XNOR U19982 ( .A(n19643), .B(n19689), .Z(n19676) );
  AND U19983 ( .A(n19645), .B(n19644), .Z(n19649) );
  NAND U19984 ( .A(n19647), .B(n19646), .Z(n19648) );
  NANDN U19985 ( .A(n19649), .B(n19648), .Z(n19685) );
  NAND U19986 ( .A(n19808), .B(n19650), .Z(n19652) );
  XOR U19987 ( .A(b[13]), .B(a[252]), .Z(n19695) );
  NAND U19988 ( .A(n19768), .B(n19695), .Z(n19651) );
  NAND U19989 ( .A(n19652), .B(n19651), .Z(n19683) );
  NAND U19990 ( .A(n19653), .B(n19724), .Z(n19655) );
  XOR U19991 ( .A(b[11]), .B(a[254]), .Z(n19691) );
  NAND U19992 ( .A(n19692), .B(n19691), .Z(n19654) );
  NAND U19993 ( .A(n19655), .B(n19654), .Z(n19682) );
  XNOR U19994 ( .A(n19679), .B(n19678), .Z(n19671) );
  NAND U19995 ( .A(n19657), .B(n19656), .Z(n19661) );
  NAND U19996 ( .A(n19659), .B(n19658), .Z(n19660) );
  AND U19997 ( .A(n19661), .B(n19660), .Z(n19670) );
  XOR U19998 ( .A(n19673), .B(n19672), .Z(n19664) );
  XOR U19999 ( .A(n19667), .B(n19666), .Z(n19662) );
  XOR U20000 ( .A(n19663), .B(n19662), .Z(c[504]) );
  AND U20001 ( .A(n19663), .B(n19662), .Z(n19702) );
  NAND U20002 ( .A(n19665), .B(n19664), .Z(n19669) );
  NANDN U20003 ( .A(n19667), .B(n19666), .Z(n19668) );
  AND U20004 ( .A(n19669), .B(n19668), .Z(n19706) );
  NAND U20005 ( .A(n19671), .B(n19670), .Z(n19675) );
  NAND U20006 ( .A(n19673), .B(n19672), .Z(n19674) );
  NAND U20007 ( .A(n19675), .B(n19674), .Z(n19704) );
  NAND U20008 ( .A(n19677), .B(n19676), .Z(n19681) );
  NAND U20009 ( .A(n19679), .B(n19678), .Z(n19680) );
  AND U20010 ( .A(n19681), .B(n19680), .Z(n19741) );
  NAND U20011 ( .A(n19683), .B(n19682), .Z(n19687) );
  NAND U20012 ( .A(n19685), .B(n19684), .Z(n19686) );
  NAND U20013 ( .A(n19687), .B(n19686), .Z(n19739) );
  NAND U20014 ( .A(n19691), .B(n19724), .Z(n19694) );
  XOR U20015 ( .A(a[255]), .B(b[11]), .Z(n19725) );
  NAND U20016 ( .A(n19692), .B(n19725), .Z(n19693) );
  NAND U20017 ( .A(n19694), .B(n19693), .Z(n19710) );
  NAND U20018 ( .A(n19808), .B(n19695), .Z(n19697) );
  XOR U20019 ( .A(b[13]), .B(a[253]), .Z(n19729) );
  NAND U20020 ( .A(n19768), .B(n19729), .Z(n19696) );
  NAND U20021 ( .A(n19697), .B(n19696), .Z(n19716) );
  NAND U20022 ( .A(n19838), .B(n19698), .Z(n19700) );
  XOR U20023 ( .A(b[15]), .B(a[251]), .Z(n19721) );
  NAND U20024 ( .A(n19805), .B(n19721), .Z(n19699) );
  NAND U20025 ( .A(n19700), .B(n19699), .Z(n19715) );
  AND U20026 ( .A(b[15]), .B(a[249]), .Z(n19735) );
  XOR U20027 ( .A(n19734), .B(n19735), .Z(n19733) );
  XOR U20028 ( .A(n19732), .B(n19733), .Z(n19717) );
  XOR U20029 ( .A(n19718), .B(n19717), .Z(n19709) );
  XOR U20030 ( .A(n19741), .B(n19740), .Z(n19703) );
  XOR U20031 ( .A(n19706), .B(n19705), .Z(n19701) );
  XOR U20032 ( .A(n19702), .B(n19701), .Z(c[505]) );
  AND U20033 ( .A(n19702), .B(n19701), .Z(n19745) );
  NAND U20034 ( .A(n19704), .B(n19703), .Z(n19708) );
  NANDN U20035 ( .A(n19706), .B(n19705), .Z(n19707) );
  AND U20036 ( .A(n19708), .B(n19707), .Z(n19749) );
  NAND U20037 ( .A(n19710), .B(n19709), .Z(n19714) );
  NAND U20038 ( .A(n19712), .B(n19711), .Z(n19713) );
  NAND U20039 ( .A(n19714), .B(n19713), .Z(n19755) );
  NAND U20040 ( .A(n19716), .B(n19715), .Z(n19720) );
  NAND U20041 ( .A(n19718), .B(n19717), .Z(n19719) );
  NAND U20042 ( .A(n19720), .B(n19719), .Z(n19753) );
  NAND U20043 ( .A(n19838), .B(n19721), .Z(n19723) );
  XOR U20044 ( .A(b[15]), .B(a[252]), .Z(n19764) );
  NAND U20045 ( .A(n19805), .B(n19764), .Z(n19722) );
  NAND U20046 ( .A(n19723), .B(n19722), .Z(n19775) );
  AND U20047 ( .A(b[15]), .B(a[250]), .Z(n19798) );
  AND U20048 ( .A(n19725), .B(n19724), .Z(n19728) );
  XOR U20049 ( .A(b[10]), .B(b[9]), .Z(n19726) );
  NAND U20050 ( .A(b[11]), .B(n19726), .Z(n19727) );
  NANDN U20051 ( .A(n19728), .B(n19727), .Z(n19772) );
  XNOR U20052 ( .A(n19798), .B(n19772), .Z(n19774) );
  NAND U20053 ( .A(n19808), .B(n19729), .Z(n19731) );
  XOR U20054 ( .A(b[13]), .B(a[254]), .Z(n19767) );
  NAND U20055 ( .A(n19768), .B(n19767), .Z(n19730) );
  NAND U20056 ( .A(n19731), .B(n19730), .Z(n19759) );
  AND U20057 ( .A(n19733), .B(n19732), .Z(n19737) );
  NAND U20058 ( .A(n19735), .B(n19734), .Z(n19736) );
  NANDN U20059 ( .A(n19737), .B(n19736), .Z(n19758) );
  XOR U20060 ( .A(n19761), .B(n19760), .Z(n19752) );
  NAND U20061 ( .A(n19739), .B(n19738), .Z(n19743) );
  NANDN U20062 ( .A(n19741), .B(n19740), .Z(n19742) );
  AND U20063 ( .A(n19743), .B(n19742), .Z(n19747) );
  XOR U20064 ( .A(n19746), .B(n19747), .Z(n19748) );
  XOR U20065 ( .A(n19749), .B(n19748), .Z(n19744) );
  XOR U20066 ( .A(n19745), .B(n19744), .Z(c[506]) );
  AND U20067 ( .A(n19745), .B(n19744), .Z(n19779) );
  NAND U20068 ( .A(n19747), .B(n19746), .Z(n19751) );
  NANDN U20069 ( .A(n19749), .B(n19748), .Z(n19750) );
  AND U20070 ( .A(n19751), .B(n19750), .Z(n19783) );
  NAND U20071 ( .A(n19753), .B(n19752), .Z(n19757) );
  NAND U20072 ( .A(n19755), .B(n19754), .Z(n19756) );
  AND U20073 ( .A(n19757), .B(n19756), .Z(n19781) );
  NAND U20074 ( .A(n19759), .B(n19758), .Z(n19763) );
  NAND U20075 ( .A(n19761), .B(n19760), .Z(n19762) );
  AND U20076 ( .A(n19763), .B(n19762), .Z(n19789) );
  NAND U20077 ( .A(n19838), .B(n19764), .Z(n19766) );
  XOR U20078 ( .A(b[15]), .B(a[253]), .Z(n19804) );
  NAND U20079 ( .A(n19805), .B(n19804), .Z(n19765) );
  NAND U20080 ( .A(n19766), .B(n19765), .Z(n19793) );
  NAND U20081 ( .A(n19808), .B(n19767), .Z(n19770) );
  XOR U20082 ( .A(a[255]), .B(b[13]), .Z(n19809) );
  NAND U20083 ( .A(n19768), .B(n19809), .Z(n19769) );
  NAND U20084 ( .A(n19770), .B(n19769), .Z(n19792) );
  IV U20085 ( .A(n19798), .Z(n19773) );
  AND U20086 ( .A(b[15]), .B(a[251]), .Z(n19800) );
  XNOR U20087 ( .A(n19771), .B(n19800), .Z(n19799) );
  XNOR U20088 ( .A(n19773), .B(n19799), .Z(n19794) );
  XNOR U20089 ( .A(n19795), .B(n19794), .Z(n19787) );
  NAND U20090 ( .A(n19773), .B(n19772), .Z(n19777) );
  NAND U20091 ( .A(n19775), .B(n19774), .Z(n19776) );
  AND U20092 ( .A(n19777), .B(n19776), .Z(n19786) );
  XOR U20093 ( .A(n19789), .B(n19788), .Z(n19780) );
  XOR U20094 ( .A(n19781), .B(n19780), .Z(n19782) );
  XOR U20095 ( .A(n19783), .B(n19782), .Z(n19778) );
  XOR U20096 ( .A(n19779), .B(n19778), .Z(c[507]) );
  AND U20097 ( .A(n19779), .B(n19778), .Z(n19814) );
  NAND U20098 ( .A(n19781), .B(n19780), .Z(n19785) );
  NANDN U20099 ( .A(n19783), .B(n19782), .Z(n19784) );
  AND U20100 ( .A(n19785), .B(n19784), .Z(n19818) );
  NAND U20101 ( .A(n19787), .B(n19786), .Z(n19791) );
  NAND U20102 ( .A(n19789), .B(n19788), .Z(n19790) );
  NAND U20103 ( .A(n19791), .B(n19790), .Z(n19816) );
  NAND U20104 ( .A(n19793), .B(n19792), .Z(n19797) );
  NAND U20105 ( .A(n19795), .B(n19794), .Z(n19796) );
  AND U20106 ( .A(n19797), .B(n19796), .Z(n19833) );
  AND U20107 ( .A(n19799), .B(n19798), .Z(n19803) );
  NAND U20108 ( .A(n19801), .B(n19800), .Z(n19802) );
  NANDN U20109 ( .A(n19803), .B(n19802), .Z(n19831) );
  NAND U20110 ( .A(n19838), .B(n19804), .Z(n19807) );
  XOR U20111 ( .A(b[15]), .B(a[254]), .Z(n19822) );
  NAND U20112 ( .A(n19805), .B(n19822), .Z(n19806) );
  NAND U20113 ( .A(n19807), .B(n19806), .Z(n19827) );
  AND U20114 ( .A(b[15]), .B(a[252]), .Z(n19844) );
  AND U20115 ( .A(n19809), .B(n19808), .Z(n19812) );
  XOR U20116 ( .A(b[12]), .B(b[11]), .Z(n19810) );
  NAND U20117 ( .A(b[13]), .B(n19810), .Z(n19811) );
  NANDN U20118 ( .A(n19812), .B(n19811), .Z(n19825) );
  XNOR U20119 ( .A(n19844), .B(n19825), .Z(n19826) );
  XOR U20120 ( .A(n19833), .B(n19832), .Z(n19815) );
  XOR U20121 ( .A(n19818), .B(n19817), .Z(n19813) );
  XOR U20122 ( .A(n19814), .B(n19813), .Z(c[508]) );
  AND U20123 ( .A(n19814), .B(n19813), .Z(n19837) );
  NAND U20124 ( .A(n19816), .B(n19815), .Z(n19820) );
  NANDN U20125 ( .A(n19818), .B(n19817), .Z(n19819) );
  AND U20126 ( .A(n19820), .B(n19819), .Z(n19852) );
  AND U20127 ( .A(b[15]), .B(a[253]), .Z(n19845) );
  XOR U20128 ( .A(n19821), .B(n19845), .Z(n19843) );
  XNOR U20129 ( .A(n19844), .B(n19843), .Z(n19855) );
  NAND U20130 ( .A(n19838), .B(n19822), .Z(n19824) );
  XNOR U20131 ( .A(a[255]), .B(b[15]), .Z(n19839) );
  OR U20132 ( .A(n19839), .B(n19840), .Z(n19823) );
  NAND U20133 ( .A(n19824), .B(n19823), .Z(n19856) );
  NANDN U20134 ( .A(n19844), .B(n19825), .Z(n19829) );
  NAND U20135 ( .A(n19827), .B(n19826), .Z(n19828) );
  NAND U20136 ( .A(n19829), .B(n19828), .Z(n19857) );
  XNOR U20137 ( .A(n19858), .B(n19857), .Z(n19850) );
  NAND U20138 ( .A(n19831), .B(n19830), .Z(n19835) );
  NANDN U20139 ( .A(n19833), .B(n19832), .Z(n19834) );
  AND U20140 ( .A(n19835), .B(n19834), .Z(n19849) );
  XOR U20141 ( .A(n19852), .B(n19851), .Z(n19836) );
  XOR U20142 ( .A(n19837), .B(n19836), .Z(c[509]) );
  AND U20143 ( .A(n19837), .B(n19836), .Z(n19862) );
  NANDN U20144 ( .A(n19839), .B(n19838), .Z(n19842) );
  NANDN U20145 ( .A(n19840), .B(b[15]), .Z(n19841) );
  NAND U20146 ( .A(n19842), .B(n19841), .Z(n19874) );
  ANDN U20147 ( .B(n19844), .A(n19843), .Z(n19848) );
  NAND U20148 ( .A(n19846), .B(n19845), .Z(n19847) );
  NANDN U20149 ( .A(n19848), .B(n19847), .Z(n19873) );
  XOR U20150 ( .A(n19874), .B(n19873), .Z(n19872) );
  NAND U20151 ( .A(b[15]), .B(a[254]), .Z(n19871) );
  XOR U20152 ( .A(n19872), .B(n19871), .Z(n19865) );
  NAND U20153 ( .A(n19850), .B(n19849), .Z(n19854) );
  NANDN U20154 ( .A(n19852), .B(n19851), .Z(n19853) );
  NAND U20155 ( .A(n19854), .B(n19853), .Z(n19863) );
  NAND U20156 ( .A(n19856), .B(n19855), .Z(n19860) );
  NAND U20157 ( .A(n19858), .B(n19857), .Z(n19859) );
  AND U20158 ( .A(n19860), .B(n19859), .Z(n19864) );
  XOR U20159 ( .A(n19865), .B(n19866), .Z(n19861) );
  XOR U20160 ( .A(n19862), .B(n19861), .Z(c[510]) );
  NAND U20161 ( .A(n19862), .B(n19861), .Z(n19870) );
  AND U20162 ( .A(n19864), .B(n19863), .Z(n19868) );
  ANDN U20163 ( .B(n19866), .A(n19865), .Z(n19867) );
  OR U20164 ( .A(n19868), .B(n19867), .Z(n19869) );
  AND U20165 ( .A(n19870), .B(n19869), .Z(n19883) );
  NAND U20166 ( .A(n19872), .B(n19871), .Z(n19876) );
  NAND U20167 ( .A(n19874), .B(n19873), .Z(n19875) );
  AND U20168 ( .A(n19876), .B(n19875), .Z(n19881) );
  XNOR U20169 ( .A(a[255]), .B(a[254]), .Z(n19877) );
  XNOR U20170 ( .A(n19878), .B(n19877), .Z(n19879) );
  NAND U20171 ( .A(b[15]), .B(n19879), .Z(n19880) );
  XNOR U20172 ( .A(n19881), .B(n19880), .Z(n19882) );
  XNOR U20173 ( .A(n19883), .B(n19882), .Z(c[511]) );
endmodule

