
module hamming_N1600_CC32 ( clk, rst, x, y, o );
  input [49:0] x;
  input [49:0] y;
  output [10:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302;
  wire   [10:0] oglobal;

  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  OR U53 ( .A(n65), .B(n64), .Z(n1) );
  NANDN U54 ( .A(n67), .B(n66), .Z(n2) );
  NAND U55 ( .A(n1), .B(n2), .Z(n167) );
  XOR U56 ( .A(n171), .B(n170), .Z(n180) );
  NAND U57 ( .A(n39), .B(n40), .Z(n3) );
  XOR U58 ( .A(n40), .B(n39), .Z(n4) );
  NANDN U59 ( .A(n41), .B(n4), .Z(n5) );
  NAND U60 ( .A(n3), .B(n5), .Z(n186) );
  NAND U61 ( .A(n200), .B(n199), .Z(n6) );
  XOR U62 ( .A(n199), .B(n200), .Z(n7) );
  NAND U63 ( .A(n7), .B(n198), .Z(n8) );
  NAND U64 ( .A(n6), .B(n8), .Z(n232) );
  NAND U65 ( .A(n166), .B(n165), .Z(n9) );
  XOR U66 ( .A(n165), .B(n166), .Z(n10) );
  NANDN U67 ( .A(n167), .B(n10), .Z(n11) );
  NAND U68 ( .A(n9), .B(n11), .Z(n239) );
  XNOR U69 ( .A(n33), .B(n34), .Z(n35) );
  XNOR U70 ( .A(n201), .B(n202), .Z(n203) );
  XNOR U71 ( .A(n208), .B(n209), .Z(n210) );
  OR U72 ( .A(n49), .B(n48), .Z(n12) );
  NANDN U73 ( .A(n51), .B(n50), .Z(n13) );
  NAND U74 ( .A(n12), .B(n13), .Z(n215) );
  XNOR U75 ( .A(n168), .B(n169), .Z(n171) );
  OR U76 ( .A(n69), .B(n68), .Z(n14) );
  NANDN U77 ( .A(n71), .B(n70), .Z(n15) );
  AND U78 ( .A(n14), .B(n15), .Z(n166) );
  OR U79 ( .A(n138), .B(n137), .Z(n16) );
  NANDN U80 ( .A(n140), .B(n139), .Z(n17) );
  NAND U81 ( .A(n16), .B(n17), .Z(n162) );
  NANDN U82 ( .A(n74), .B(n73), .Z(n18) );
  NANDN U83 ( .A(n75), .B(n76), .Z(n19) );
  NAND U84 ( .A(n18), .B(n19), .Z(n199) );
  XNOR U85 ( .A(n278), .B(n279), .Z(n269) );
  XNOR U86 ( .A(x[44]), .B(y[44]), .Z(n140) );
  XNOR U87 ( .A(x[48]), .B(y[48]), .Z(n138) );
  XNOR U88 ( .A(x[46]), .B(y[46]), .Z(n137) );
  XOR U89 ( .A(n138), .B(n137), .Z(n139) );
  XOR U90 ( .A(n140), .B(n139), .Z(n41) );
  XNOR U91 ( .A(x[40]), .B(y[40]), .Z(n110) );
  XOR U92 ( .A(x[42]), .B(y[42]), .Z(n108) );
  XNOR U93 ( .A(oglobal[0]), .B(n108), .Z(n109) );
  XOR U94 ( .A(n110), .B(n109), .Z(n40) );
  XNOR U95 ( .A(x[4]), .B(y[4]), .Z(n128) );
  XNOR U96 ( .A(x[6]), .B(y[6]), .Z(n126) );
  XNOR U97 ( .A(x[8]), .B(y[8]), .Z(n125) );
  XNOR U98 ( .A(n126), .B(n125), .Z(n127) );
  XNOR U99 ( .A(n128), .B(n127), .Z(n76) );
  XNOR U100 ( .A(x[10]), .B(y[10]), .Z(n134) );
  XNOR U101 ( .A(x[14]), .B(y[14]), .Z(n132) );
  XNOR U102 ( .A(x[12]), .B(y[12]), .Z(n131) );
  XNOR U103 ( .A(n132), .B(n131), .Z(n133) );
  XNOR U104 ( .A(n134), .B(n133), .Z(n73) );
  XNOR U105 ( .A(x[16]), .B(y[16]), .Z(n105) );
  XNOR U106 ( .A(x[20]), .B(y[20]), .Z(n103) );
  XNOR U107 ( .A(x[18]), .B(y[18]), .Z(n102) );
  XNOR U108 ( .A(n103), .B(n102), .Z(n104) );
  XOR U109 ( .A(n105), .B(n104), .Z(n74) );
  XOR U110 ( .A(n73), .B(n74), .Z(n75) );
  XOR U111 ( .A(n76), .B(n75), .Z(n39) );
  XOR U112 ( .A(n40), .B(n39), .Z(n20) );
  XNOR U113 ( .A(n41), .B(n20), .Z(n23) );
  XNOR U114 ( .A(x[37]), .B(y[37]), .Z(n45) );
  XNOR U115 ( .A(x[45]), .B(y[45]), .Z(n42) );
  XNOR U116 ( .A(x[35]), .B(y[35]), .Z(n43) );
  XOR U117 ( .A(n42), .B(n43), .Z(n44) );
  XOR U118 ( .A(n45), .B(n44), .Z(n33) );
  XNOR U119 ( .A(x[29]), .B(y[29]), .Z(n61) );
  XNOR U120 ( .A(x[27]), .B(y[27]), .Z(n58) );
  XNOR U121 ( .A(x[49]), .B(y[49]), .Z(n59) );
  XOR U122 ( .A(n58), .B(n59), .Z(n60) );
  XNOR U123 ( .A(n61), .B(n60), .Z(n34) );
  XNOR U124 ( .A(x[33]), .B(y[33]), .Z(n55) );
  XNOR U125 ( .A(x[31]), .B(y[31]), .Z(n52) );
  XNOR U126 ( .A(x[47]), .B(y[47]), .Z(n53) );
  XOR U127 ( .A(n52), .B(n53), .Z(n54) );
  XNOR U128 ( .A(n55), .B(n54), .Z(n36) );
  XOR U129 ( .A(n35), .B(n36), .Z(n90) );
  XNOR U130 ( .A(x[1]), .B(y[1]), .Z(n150) );
  XNOR U131 ( .A(x[2]), .B(y[2]), .Z(n148) );
  XNOR U132 ( .A(x[0]), .B(y[0]), .Z(n147) );
  XNOR U133 ( .A(n148), .B(n147), .Z(n149) );
  XNOR U134 ( .A(n150), .B(n149), .Z(n77) );
  XNOR U135 ( .A(x[7]), .B(y[7]), .Z(n144) );
  XNOR U136 ( .A(x[5]), .B(y[5]), .Z(n142) );
  XNOR U137 ( .A(x[3]), .B(y[3]), .Z(n141) );
  XNOR U138 ( .A(n142), .B(n141), .Z(n143) );
  XOR U139 ( .A(n144), .B(n143), .Z(n78) );
  XOR U140 ( .A(n77), .B(n78), .Z(n80) );
  XNOR U141 ( .A(x[11]), .B(y[11]), .Z(n154) );
  XNOR U142 ( .A(x[9]), .B(y[9]), .Z(n153) );
  XNOR U143 ( .A(n154), .B(n153), .Z(n156) );
  XNOR U144 ( .A(x[13]), .B(y[13]), .Z(n155) );
  XOR U145 ( .A(n156), .B(n155), .Z(n79) );
  XOR U146 ( .A(n80), .B(n79), .Z(n91) );
  XNOR U147 ( .A(n90), .B(n91), .Z(n92) );
  XNOR U148 ( .A(x[28]), .B(y[28]), .Z(n116) );
  XNOR U149 ( .A(x[32]), .B(y[32]), .Z(n114) );
  XNOR U150 ( .A(x[30]), .B(y[30]), .Z(n113) );
  XNOR U151 ( .A(n114), .B(n113), .Z(n115) );
  XNOR U152 ( .A(n116), .B(n115), .Z(n83) );
  XNOR U153 ( .A(x[34]), .B(y[34]), .Z(n122) );
  XNOR U154 ( .A(x[38]), .B(y[38]), .Z(n120) );
  XNOR U155 ( .A(x[36]), .B(y[36]), .Z(n119) );
  XNOR U156 ( .A(n120), .B(n119), .Z(n121) );
  XOR U157 ( .A(n122), .B(n121), .Z(n84) );
  XNOR U158 ( .A(n83), .B(n84), .Z(n85) );
  XNOR U159 ( .A(x[22]), .B(y[22]), .Z(n99) );
  XNOR U160 ( .A(x[26]), .B(y[26]), .Z(n97) );
  XNOR U161 ( .A(x[24]), .B(y[24]), .Z(n96) );
  XNOR U162 ( .A(n97), .B(n96), .Z(n98) );
  XOR U163 ( .A(n99), .B(n98), .Z(n86) );
  XOR U164 ( .A(n85), .B(n86), .Z(n93) );
  XNOR U165 ( .A(n92), .B(n93), .Z(n22) );
  XNOR U166 ( .A(x[19]), .B(y[19]), .Z(n67) );
  XNOR U167 ( .A(x[15]), .B(y[15]), .Z(n65) );
  XNOR U168 ( .A(x[17]), .B(y[17]), .Z(n64) );
  XOR U169 ( .A(n65), .B(n64), .Z(n66) );
  XOR U170 ( .A(n67), .B(n66), .Z(n27) );
  XNOR U171 ( .A(x[25]), .B(y[25]), .Z(n71) );
  XNOR U172 ( .A(x[21]), .B(y[21]), .Z(n69) );
  XNOR U173 ( .A(x[23]), .B(y[23]), .Z(n68) );
  XOR U174 ( .A(n69), .B(n68), .Z(n70) );
  XNOR U175 ( .A(n71), .B(n70), .Z(n28) );
  XNOR U176 ( .A(n27), .B(n28), .Z(n29) );
  XNOR U177 ( .A(x[41]), .B(y[41]), .Z(n51) );
  XNOR U178 ( .A(x[43]), .B(y[43]), .Z(n49) );
  XNOR U179 ( .A(x[39]), .B(y[39]), .Z(n48) );
  XOR U180 ( .A(n49), .B(n48), .Z(n50) );
  XNOR U181 ( .A(n51), .B(n50), .Z(n30) );
  XOR U182 ( .A(n29), .B(n30), .Z(n21) );
  XNOR U183 ( .A(n22), .B(n21), .Z(n24) );
  XOR U184 ( .A(n23), .B(n24), .Z(o[0]) );
  NANDN U185 ( .A(n22), .B(n21), .Z(n26) );
  NAND U186 ( .A(n24), .B(n23), .Z(n25) );
  NAND U187 ( .A(n26), .B(n25), .Z(n220) );
  NANDN U188 ( .A(n28), .B(n27), .Z(n32) );
  NANDN U189 ( .A(n30), .B(n29), .Z(n31) );
  NAND U190 ( .A(n32), .B(n31), .Z(n174) );
  NANDN U191 ( .A(n34), .B(n33), .Z(n38) );
  NANDN U192 ( .A(n36), .B(n35), .Z(n37) );
  AND U193 ( .A(n38), .B(n37), .Z(n175) );
  XNOR U194 ( .A(n174), .B(n175), .Z(n176) );
  OR U195 ( .A(n43), .B(n42), .Z(n47) );
  NANDN U196 ( .A(n45), .B(n44), .Z(n46) );
  AND U197 ( .A(n47), .B(n46), .Z(n207) );
  XOR U198 ( .A(oglobal[1]), .B(n207), .Z(n214) );
  XOR U199 ( .A(n214), .B(n215), .Z(n217) );
  OR U200 ( .A(n53), .B(n52), .Z(n57) );
  NANDN U201 ( .A(n55), .B(n54), .Z(n56) );
  NAND U202 ( .A(n57), .B(n56), .Z(n216) );
  XOR U203 ( .A(n217), .B(n216), .Z(n187) );
  XOR U204 ( .A(n186), .B(n187), .Z(n189) );
  OR U205 ( .A(n59), .B(n58), .Z(n63) );
  NANDN U206 ( .A(n61), .B(n60), .Z(n62) );
  AND U207 ( .A(n63), .B(n62), .Z(n165) );
  XOR U208 ( .A(n167), .B(n166), .Z(n72) );
  XOR U209 ( .A(n165), .B(n72), .Z(n188) );
  XNOR U210 ( .A(n189), .B(n188), .Z(n177) );
  XNOR U211 ( .A(n176), .B(n177), .Z(n221) );
  XNOR U212 ( .A(n220), .B(n221), .Z(n222) );
  NANDN U213 ( .A(n78), .B(n77), .Z(n82) );
  OR U214 ( .A(n80), .B(n79), .Z(n81) );
  NAND U215 ( .A(n82), .B(n81), .Z(n200) );
  NANDN U216 ( .A(n84), .B(n83), .Z(n88) );
  NANDN U217 ( .A(n86), .B(n85), .Z(n87) );
  NAND U218 ( .A(n88), .B(n87), .Z(n198) );
  XNOR U219 ( .A(n200), .B(n198), .Z(n89) );
  XOR U220 ( .A(n199), .B(n89), .Z(n194) );
  NANDN U221 ( .A(n91), .B(n90), .Z(n95) );
  NAND U222 ( .A(n93), .B(n92), .Z(n94) );
  NAND U223 ( .A(n95), .B(n94), .Z(n192) );
  OR U224 ( .A(n97), .B(n96), .Z(n101) );
  OR U225 ( .A(n99), .B(n98), .Z(n100) );
  NAND U226 ( .A(n101), .B(n100), .Z(n209) );
  OR U227 ( .A(n103), .B(n102), .Z(n107) );
  OR U228 ( .A(n105), .B(n104), .Z(n106) );
  AND U229 ( .A(n107), .B(n106), .Z(n208) );
  NAND U230 ( .A(n108), .B(oglobal[0]), .Z(n112) );
  OR U231 ( .A(n110), .B(n109), .Z(n111) );
  AND U232 ( .A(n112), .B(n111), .Z(n211) );
  XNOR U233 ( .A(n210), .B(n211), .Z(n183) );
  OR U234 ( .A(n114), .B(n113), .Z(n118) );
  OR U235 ( .A(n116), .B(n115), .Z(n117) );
  NAND U236 ( .A(n118), .B(n117), .Z(n169) );
  OR U237 ( .A(n120), .B(n119), .Z(n124) );
  OR U238 ( .A(n122), .B(n121), .Z(n123) );
  AND U239 ( .A(n124), .B(n123), .Z(n168) );
  OR U240 ( .A(n126), .B(n125), .Z(n130) );
  OR U241 ( .A(n128), .B(n127), .Z(n129) );
  NAND U242 ( .A(n130), .B(n129), .Z(n160) );
  OR U243 ( .A(n132), .B(n131), .Z(n136) );
  OR U244 ( .A(n134), .B(n133), .Z(n135) );
  NAND U245 ( .A(n136), .B(n135), .Z(n159) );
  XNOR U246 ( .A(n160), .B(n159), .Z(n161) );
  XOR U247 ( .A(n161), .B(n162), .Z(n170) );
  OR U248 ( .A(n142), .B(n141), .Z(n146) );
  OR U249 ( .A(n144), .B(n143), .Z(n145) );
  NAND U250 ( .A(n146), .B(n145), .Z(n204) );
  OR U251 ( .A(n148), .B(n147), .Z(n152) );
  OR U252 ( .A(n150), .B(n149), .Z(n151) );
  NAND U253 ( .A(n152), .B(n151), .Z(n202) );
  OR U254 ( .A(n154), .B(n153), .Z(n158) );
  OR U255 ( .A(n156), .B(n155), .Z(n157) );
  AND U256 ( .A(n158), .B(n157), .Z(n201) );
  XNOR U257 ( .A(n204), .B(n203), .Z(n181) );
  XOR U258 ( .A(n180), .B(n181), .Z(n182) );
  XNOR U259 ( .A(n183), .B(n182), .Z(n193) );
  XNOR U260 ( .A(n192), .B(n193), .Z(n195) );
  XOR U261 ( .A(n194), .B(n195), .Z(n223) );
  XOR U262 ( .A(n222), .B(n223), .Z(o[1]) );
  OR U263 ( .A(n160), .B(n159), .Z(n164) );
  OR U264 ( .A(n162), .B(n161), .Z(n163) );
  NAND U265 ( .A(n164), .B(n163), .Z(n242) );
  NANDN U266 ( .A(n169), .B(n168), .Z(n173) );
  NAND U267 ( .A(n171), .B(n170), .Z(n172) );
  AND U268 ( .A(n173), .B(n172), .Z(n240) );
  XNOR U269 ( .A(n239), .B(n240), .Z(n241) );
  XNOR U270 ( .A(n242), .B(n241), .Z(n254) );
  NANDN U271 ( .A(n175), .B(n174), .Z(n179) );
  NANDN U272 ( .A(n177), .B(n176), .Z(n178) );
  NAND U273 ( .A(n179), .B(n178), .Z(n251) );
  NAND U274 ( .A(n181), .B(n180), .Z(n185) );
  NANDN U275 ( .A(n183), .B(n182), .Z(n184) );
  AND U276 ( .A(n185), .B(n184), .Z(n252) );
  XNOR U277 ( .A(n251), .B(n252), .Z(n253) );
  XOR U278 ( .A(n254), .B(n253), .Z(n257) );
  NANDN U279 ( .A(n187), .B(n186), .Z(n191) );
  NANDN U280 ( .A(n189), .B(n188), .Z(n190) );
  NAND U281 ( .A(n191), .B(n190), .Z(n229) );
  NANDN U282 ( .A(n193), .B(n192), .Z(n197) );
  NAND U283 ( .A(n195), .B(n194), .Z(n196) );
  NAND U284 ( .A(n197), .B(n196), .Z(n226) );
  NANDN U285 ( .A(n202), .B(n201), .Z(n206) );
  NANDN U286 ( .A(n204), .B(n203), .Z(n205) );
  AND U287 ( .A(n206), .B(n205), .Z(n233) );
  XOR U288 ( .A(n232), .B(n233), .Z(n235) );
  ANDN U289 ( .B(oglobal[1]), .A(n207), .Z(n238) );
  XOR U290 ( .A(oglobal[2]), .B(n238), .Z(n248) );
  NANDN U291 ( .A(n209), .B(n208), .Z(n213) );
  NAND U292 ( .A(n211), .B(n210), .Z(n212) );
  AND U293 ( .A(n213), .B(n212), .Z(n245) );
  NANDN U294 ( .A(n215), .B(n214), .Z(n219) );
  OR U295 ( .A(n217), .B(n216), .Z(n218) );
  AND U296 ( .A(n219), .B(n218), .Z(n246) );
  XOR U297 ( .A(n245), .B(n246), .Z(n247) );
  XOR U298 ( .A(n248), .B(n247), .Z(n234) );
  XOR U299 ( .A(n235), .B(n234), .Z(n227) );
  XNOR U300 ( .A(n226), .B(n227), .Z(n228) );
  XNOR U301 ( .A(n229), .B(n228), .Z(n258) );
  XNOR U302 ( .A(n257), .B(n258), .Z(n259) );
  NANDN U303 ( .A(n221), .B(n220), .Z(n225) );
  NAND U304 ( .A(n223), .B(n222), .Z(n224) );
  AND U305 ( .A(n225), .B(n224), .Z(n260) );
  XNOR U306 ( .A(n259), .B(n260), .Z(o[2]) );
  NANDN U307 ( .A(n227), .B(n226), .Z(n231) );
  NAND U308 ( .A(n229), .B(n228), .Z(n230) );
  NAND U309 ( .A(n231), .B(n230), .Z(n264) );
  NANDN U310 ( .A(n233), .B(n232), .Z(n237) );
  OR U311 ( .A(n235), .B(n234), .Z(n236) );
  NAND U312 ( .A(n237), .B(n236), .Z(n270) );
  AND U313 ( .A(n238), .B(oglobal[2]), .Z(n275) );
  XOR U314 ( .A(oglobal[3]), .B(n275), .Z(n279) );
  NANDN U315 ( .A(n240), .B(n239), .Z(n244) );
  NAND U316 ( .A(n242), .B(n241), .Z(n243) );
  AND U317 ( .A(n244), .B(n243), .Z(n276) );
  OR U318 ( .A(n246), .B(n245), .Z(n250) );
  NANDN U319 ( .A(n248), .B(n247), .Z(n249) );
  AND U320 ( .A(n250), .B(n249), .Z(n277) );
  XOR U321 ( .A(n276), .B(n277), .Z(n278) );
  XNOR U322 ( .A(n270), .B(n269), .Z(n272) );
  NANDN U323 ( .A(n252), .B(n251), .Z(n256) );
  NANDN U324 ( .A(n254), .B(n253), .Z(n255) );
  NAND U325 ( .A(n256), .B(n255), .Z(n271) );
  XOR U326 ( .A(n272), .B(n271), .Z(n263) );
  XNOR U327 ( .A(n264), .B(n263), .Z(n266) );
  NANDN U328 ( .A(n258), .B(n257), .Z(n262) );
  NANDN U329 ( .A(n260), .B(n259), .Z(n261) );
  AND U330 ( .A(n262), .B(n261), .Z(n265) );
  XOR U331 ( .A(n266), .B(n265), .Z(o[3]) );
  NAND U332 ( .A(n264), .B(n263), .Z(n268) );
  OR U333 ( .A(n266), .B(n265), .Z(n267) );
  NAND U334 ( .A(n268), .B(n267), .Z(n282) );
  OR U335 ( .A(n270), .B(n269), .Z(n274) );
  OR U336 ( .A(n272), .B(n271), .Z(n273) );
  AND U337 ( .A(n274), .B(n273), .Z(n283) );
  XNOR U338 ( .A(n282), .B(n283), .Z(n284) );
  NAND U339 ( .A(n275), .B(oglobal[3]), .Z(n288) );
  XOR U340 ( .A(oglobal[4]), .B(n288), .Z(n290) );
  OR U341 ( .A(n277), .B(n276), .Z(n281) );
  NANDN U342 ( .A(n279), .B(n278), .Z(n280) );
  NAND U343 ( .A(n281), .B(n280), .Z(n289) );
  XNOR U344 ( .A(n290), .B(n289), .Z(n285) );
  XNOR U345 ( .A(n284), .B(n285), .Z(o[4]) );
  NANDN U346 ( .A(n283), .B(n282), .Z(n287) );
  NANDN U347 ( .A(n285), .B(n284), .Z(n286) );
  NAND U348 ( .A(n287), .B(n286), .Z(n293) );
  XNOR U349 ( .A(n293), .B(oglobal[5]), .Z(n295) );
  NANDN U350 ( .A(n288), .B(oglobal[4]), .Z(n292) );
  OR U351 ( .A(n290), .B(n289), .Z(n291) );
  AND U352 ( .A(n292), .B(n291), .Z(n294) );
  XOR U353 ( .A(n295), .B(n294), .Z(o[5]) );
  NAND U354 ( .A(n293), .B(oglobal[5]), .Z(n297) );
  OR U355 ( .A(n295), .B(n294), .Z(n296) );
  AND U356 ( .A(n297), .B(n296), .Z(n298) );
  XNOR U357 ( .A(oglobal[6]), .B(n298), .Z(o[6]) );
  NANDN U358 ( .A(n298), .B(oglobal[6]), .Z(n299) );
  XNOR U359 ( .A(n299), .B(oglobal[7]), .Z(o[7]) );
  NANDN U360 ( .A(n299), .B(oglobal[7]), .Z(n300) );
  XNOR U361 ( .A(n300), .B(oglobal[8]), .Z(o[8]) );
  NANDN U362 ( .A(n300), .B(oglobal[8]), .Z(n301) );
  XNOR U363 ( .A(oglobal[9]), .B(n301), .Z(o[9]) );
  NANDN U364 ( .A(n301), .B(oglobal[9]), .Z(n302) );
  XNOR U365 ( .A(oglobal[10]), .B(n302), .Z(o[10]) );
endmodule

