
module hamming_N16000_CC2_DW01_add_0 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61;

  XNOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U4 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U16 ( .A(B[2]), .B(A[2]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(SUM[1]) );
  XOR U18 ( .A(B[1]), .B(A[1]), .Z(n18) );
  XOR U19 ( .A(A[13]), .B(n19), .Z(SUM[13]) );
  NAND U20 ( .A(n20), .B(n21), .Z(n19) );
  NAND U21 ( .A(B[12]), .B(n22), .Z(n21) );
  NANDN U22 ( .A(A[12]), .B(n23), .Z(n22) );
  NANDN U23 ( .A(n23), .B(A[12]), .Z(n20) );
  XOR U24 ( .A(n23), .B(n24), .Z(SUM[12]) );
  XNOR U25 ( .A(B[12]), .B(A[12]), .Z(n24) );
  AND U26 ( .A(n25), .B(n26), .Z(n23) );
  NAND U27 ( .A(B[11]), .B(n27), .Z(n26) );
  NANDN U28 ( .A(A[11]), .B(n28), .Z(n27) );
  NANDN U29 ( .A(n28), .B(A[11]), .Z(n25) );
  XOR U30 ( .A(n28), .B(n29), .Z(SUM[11]) );
  XNOR U31 ( .A(B[11]), .B(A[11]), .Z(n29) );
  AND U32 ( .A(n30), .B(n31), .Z(n28) );
  NAND U33 ( .A(B[10]), .B(n32), .Z(n31) );
  NANDN U34 ( .A(A[10]), .B(n33), .Z(n32) );
  NANDN U35 ( .A(n33), .B(A[10]), .Z(n30) );
  XOR U36 ( .A(n33), .B(n34), .Z(SUM[10]) );
  XNOR U37 ( .A(B[10]), .B(A[10]), .Z(n34) );
  AND U38 ( .A(n35), .B(n36), .Z(n33) );
  NAND U39 ( .A(B[9]), .B(n37), .Z(n36) );
  OR U40 ( .A(n1), .B(A[9]), .Z(n37) );
  NAND U41 ( .A(A[9]), .B(n1), .Z(n35) );
  NAND U42 ( .A(n38), .B(n39), .Z(n1) );
  NAND U43 ( .A(B[8]), .B(n40), .Z(n39) );
  NANDN U44 ( .A(A[8]), .B(n3), .Z(n40) );
  NANDN U45 ( .A(n3), .B(A[8]), .Z(n38) );
  AND U46 ( .A(n41), .B(n42), .Z(n3) );
  NAND U47 ( .A(B[7]), .B(n43), .Z(n42) );
  NANDN U48 ( .A(A[7]), .B(n5), .Z(n43) );
  NANDN U49 ( .A(n5), .B(A[7]), .Z(n41) );
  AND U50 ( .A(n44), .B(n45), .Z(n5) );
  NAND U51 ( .A(B[6]), .B(n46), .Z(n45) );
  NANDN U52 ( .A(A[6]), .B(n7), .Z(n46) );
  NANDN U53 ( .A(n7), .B(A[6]), .Z(n44) );
  AND U54 ( .A(n47), .B(n48), .Z(n7) );
  NAND U55 ( .A(B[5]), .B(n49), .Z(n48) );
  NANDN U56 ( .A(A[5]), .B(n9), .Z(n49) );
  NANDN U57 ( .A(n9), .B(A[5]), .Z(n47) );
  AND U58 ( .A(n50), .B(n51), .Z(n9) );
  NAND U59 ( .A(B[4]), .B(n52), .Z(n51) );
  NANDN U60 ( .A(A[4]), .B(n11), .Z(n52) );
  NANDN U61 ( .A(n11), .B(A[4]), .Z(n50) );
  AND U62 ( .A(n53), .B(n54), .Z(n11) );
  NAND U63 ( .A(B[3]), .B(n55), .Z(n54) );
  NANDN U64 ( .A(A[3]), .B(n13), .Z(n55) );
  NANDN U65 ( .A(n13), .B(A[3]), .Z(n53) );
  AND U66 ( .A(n56), .B(n57), .Z(n13) );
  NAND U67 ( .A(B[2]), .B(n58), .Z(n57) );
  NANDN U68 ( .A(A[2]), .B(n15), .Z(n58) );
  NANDN U69 ( .A(n15), .B(A[2]), .Z(n56) );
  AND U70 ( .A(n59), .B(n60), .Z(n15) );
  NAND U71 ( .A(B[1]), .B(n61), .Z(n60) );
  OR U72 ( .A(n17), .B(A[1]), .Z(n61) );
  NAND U73 ( .A(A[1]), .B(n17), .Z(n59) );
  AND U74 ( .A(B[0]), .B(A[0]), .Z(n17) );
  XOR U75 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_1 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57;

  IV U1 ( .A(B[12]), .Z(n1) );
  XNOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  XOR U20 ( .A(n20), .B(n1), .Z(SUM[12]) );
  AND U21 ( .A(n21), .B(n22), .Z(n20) );
  NAND U22 ( .A(B[11]), .B(n23), .Z(n22) );
  NANDN U23 ( .A(A[11]), .B(n24), .Z(n23) );
  NANDN U24 ( .A(n24), .B(A[11]), .Z(n21) );
  XOR U25 ( .A(n24), .B(n25), .Z(SUM[11]) );
  XNOR U26 ( .A(B[11]), .B(A[11]), .Z(n25) );
  AND U27 ( .A(n26), .B(n27), .Z(n24) );
  NAND U28 ( .A(B[10]), .B(n28), .Z(n27) );
  NANDN U29 ( .A(A[10]), .B(n29), .Z(n28) );
  NANDN U30 ( .A(n29), .B(A[10]), .Z(n26) );
  XOR U31 ( .A(n29), .B(n30), .Z(SUM[10]) );
  XNOR U32 ( .A(B[10]), .B(A[10]), .Z(n30) );
  AND U33 ( .A(n31), .B(n32), .Z(n29) );
  NAND U34 ( .A(B[9]), .B(n33), .Z(n32) );
  OR U35 ( .A(n2), .B(A[9]), .Z(n33) );
  NAND U36 ( .A(A[9]), .B(n2), .Z(n31) );
  NAND U37 ( .A(n34), .B(n35), .Z(n2) );
  NAND U38 ( .A(B[8]), .B(n36), .Z(n35) );
  NANDN U39 ( .A(A[8]), .B(n4), .Z(n36) );
  NANDN U40 ( .A(n4), .B(A[8]), .Z(n34) );
  AND U41 ( .A(n37), .B(n38), .Z(n4) );
  NAND U42 ( .A(B[7]), .B(n39), .Z(n38) );
  NANDN U43 ( .A(A[7]), .B(n6), .Z(n39) );
  NANDN U44 ( .A(n6), .B(A[7]), .Z(n37) );
  AND U45 ( .A(n40), .B(n41), .Z(n6) );
  NAND U46 ( .A(B[6]), .B(n42), .Z(n41) );
  NANDN U47 ( .A(A[6]), .B(n8), .Z(n42) );
  NANDN U48 ( .A(n8), .B(A[6]), .Z(n40) );
  AND U49 ( .A(n43), .B(n44), .Z(n8) );
  NAND U50 ( .A(B[5]), .B(n45), .Z(n44) );
  NANDN U51 ( .A(A[5]), .B(n10), .Z(n45) );
  NANDN U52 ( .A(n10), .B(A[5]), .Z(n43) );
  AND U53 ( .A(n46), .B(n47), .Z(n10) );
  NAND U54 ( .A(B[4]), .B(n48), .Z(n47) );
  NANDN U55 ( .A(A[4]), .B(n12), .Z(n48) );
  NANDN U56 ( .A(n12), .B(A[4]), .Z(n46) );
  AND U57 ( .A(n49), .B(n50), .Z(n12) );
  NAND U58 ( .A(B[3]), .B(n51), .Z(n50) );
  NANDN U59 ( .A(A[3]), .B(n14), .Z(n51) );
  NANDN U60 ( .A(n14), .B(A[3]), .Z(n49) );
  AND U61 ( .A(n52), .B(n53), .Z(n14) );
  NAND U62 ( .A(B[2]), .B(n54), .Z(n53) );
  NANDN U63 ( .A(A[2]), .B(n16), .Z(n54) );
  NANDN U64 ( .A(n16), .B(A[2]), .Z(n52) );
  AND U65 ( .A(n55), .B(n56), .Z(n16) );
  NAND U66 ( .A(B[1]), .B(n57), .Z(n56) );
  OR U67 ( .A(n18), .B(A[1]), .Z(n57) );
  NAND U68 ( .A(A[1]), .B(n18), .Z(n55) );
  AND U69 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U70 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_2 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56;

  NAND U1 ( .A(n20), .B(n21), .Z(SUM[12]) );
  XNOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  NAND U20 ( .A(B[11]), .B(n22), .Z(n21) );
  NANDN U21 ( .A(A[11]), .B(n23), .Z(n22) );
  NANDN U22 ( .A(n23), .B(A[11]), .Z(n20) );
  XOR U23 ( .A(n23), .B(n24), .Z(SUM[11]) );
  XNOR U24 ( .A(B[11]), .B(A[11]), .Z(n24) );
  AND U25 ( .A(n25), .B(n26), .Z(n23) );
  NAND U26 ( .A(B[10]), .B(n27), .Z(n26) );
  NANDN U27 ( .A(A[10]), .B(n28), .Z(n27) );
  NANDN U28 ( .A(n28), .B(A[10]), .Z(n25) );
  XOR U29 ( .A(n28), .B(n29), .Z(SUM[10]) );
  XNOR U30 ( .A(B[10]), .B(A[10]), .Z(n29) );
  AND U31 ( .A(n30), .B(n31), .Z(n28) );
  NAND U32 ( .A(B[9]), .B(n32), .Z(n31) );
  OR U33 ( .A(n2), .B(A[9]), .Z(n32) );
  NAND U34 ( .A(A[9]), .B(n2), .Z(n30) );
  NAND U35 ( .A(n33), .B(n34), .Z(n2) );
  NAND U36 ( .A(B[8]), .B(n35), .Z(n34) );
  NANDN U37 ( .A(A[8]), .B(n4), .Z(n35) );
  NANDN U38 ( .A(n4), .B(A[8]), .Z(n33) );
  AND U39 ( .A(n36), .B(n37), .Z(n4) );
  NAND U40 ( .A(B[7]), .B(n38), .Z(n37) );
  NANDN U41 ( .A(A[7]), .B(n6), .Z(n38) );
  NANDN U42 ( .A(n6), .B(A[7]), .Z(n36) );
  AND U43 ( .A(n39), .B(n40), .Z(n6) );
  NAND U44 ( .A(B[6]), .B(n41), .Z(n40) );
  NANDN U45 ( .A(A[6]), .B(n8), .Z(n41) );
  NANDN U46 ( .A(n8), .B(A[6]), .Z(n39) );
  AND U47 ( .A(n42), .B(n43), .Z(n8) );
  NAND U48 ( .A(B[5]), .B(n44), .Z(n43) );
  NANDN U49 ( .A(A[5]), .B(n10), .Z(n44) );
  NANDN U50 ( .A(n10), .B(A[5]), .Z(n42) );
  AND U51 ( .A(n45), .B(n46), .Z(n10) );
  NAND U52 ( .A(B[4]), .B(n47), .Z(n46) );
  NANDN U53 ( .A(A[4]), .B(n12), .Z(n47) );
  NANDN U54 ( .A(n12), .B(A[4]), .Z(n45) );
  AND U55 ( .A(n48), .B(n49), .Z(n12) );
  NAND U56 ( .A(B[3]), .B(n50), .Z(n49) );
  NANDN U57 ( .A(A[3]), .B(n14), .Z(n50) );
  NANDN U58 ( .A(n14), .B(A[3]), .Z(n48) );
  AND U59 ( .A(n51), .B(n52), .Z(n14) );
  NAND U60 ( .A(B[2]), .B(n53), .Z(n52) );
  NANDN U61 ( .A(A[2]), .B(n16), .Z(n53) );
  NANDN U62 ( .A(n16), .B(A[2]), .Z(n51) );
  AND U63 ( .A(n54), .B(n55), .Z(n16) );
  NAND U64 ( .A(B[1]), .B(n56), .Z(n55) );
  OR U65 ( .A(n18), .B(A[1]), .Z(n56) );
  NAND U66 ( .A(A[1]), .B(n18), .Z(n54) );
  AND U67 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U68 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_3 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51;

  NAND U1 ( .A(n20), .B(n21), .Z(SUM[11]) );
  XNOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  NAND U20 ( .A(B[10]), .B(n22), .Z(n21) );
  NANDN U21 ( .A(A[10]), .B(n23), .Z(n22) );
  NANDN U22 ( .A(n23), .B(A[10]), .Z(n20) );
  XOR U23 ( .A(n23), .B(n24), .Z(SUM[10]) );
  XNOR U24 ( .A(B[10]), .B(A[10]), .Z(n24) );
  AND U25 ( .A(n25), .B(n26), .Z(n23) );
  NAND U26 ( .A(B[9]), .B(n27), .Z(n26) );
  OR U27 ( .A(n2), .B(A[9]), .Z(n27) );
  NAND U28 ( .A(A[9]), .B(n2), .Z(n25) );
  NAND U29 ( .A(n28), .B(n29), .Z(n2) );
  NAND U30 ( .A(B[8]), .B(n30), .Z(n29) );
  NANDN U31 ( .A(A[8]), .B(n4), .Z(n30) );
  NANDN U32 ( .A(n4), .B(A[8]), .Z(n28) );
  AND U33 ( .A(n31), .B(n32), .Z(n4) );
  NAND U34 ( .A(B[7]), .B(n33), .Z(n32) );
  NANDN U35 ( .A(A[7]), .B(n6), .Z(n33) );
  NANDN U36 ( .A(n6), .B(A[7]), .Z(n31) );
  AND U37 ( .A(n34), .B(n35), .Z(n6) );
  NAND U38 ( .A(B[6]), .B(n36), .Z(n35) );
  NANDN U39 ( .A(A[6]), .B(n8), .Z(n36) );
  NANDN U40 ( .A(n8), .B(A[6]), .Z(n34) );
  AND U41 ( .A(n37), .B(n38), .Z(n8) );
  NAND U42 ( .A(B[5]), .B(n39), .Z(n38) );
  NANDN U43 ( .A(A[5]), .B(n10), .Z(n39) );
  NANDN U44 ( .A(n10), .B(A[5]), .Z(n37) );
  AND U45 ( .A(n40), .B(n41), .Z(n10) );
  NAND U46 ( .A(B[4]), .B(n42), .Z(n41) );
  NANDN U47 ( .A(A[4]), .B(n12), .Z(n42) );
  NANDN U48 ( .A(n12), .B(A[4]), .Z(n40) );
  AND U49 ( .A(n43), .B(n44), .Z(n12) );
  NAND U50 ( .A(B[3]), .B(n45), .Z(n44) );
  NANDN U51 ( .A(A[3]), .B(n14), .Z(n45) );
  NANDN U52 ( .A(n14), .B(A[3]), .Z(n43) );
  AND U53 ( .A(n46), .B(n47), .Z(n14) );
  NAND U54 ( .A(B[2]), .B(n48), .Z(n47) );
  NANDN U55 ( .A(A[2]), .B(n16), .Z(n48) );
  NANDN U56 ( .A(n16), .B(A[2]), .Z(n46) );
  AND U57 ( .A(n49), .B(n50), .Z(n16) );
  NAND U58 ( .A(B[1]), .B(n51), .Z(n50) );
  OR U59 ( .A(n18), .B(A[1]), .Z(n51) );
  NAND U60 ( .A(A[1]), .B(n18), .Z(n49) );
  AND U61 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U62 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_4 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51;

  NAND U1 ( .A(n20), .B(n21), .Z(SUM[11]) );
  XNOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  NAND U20 ( .A(B[10]), .B(n22), .Z(n21) );
  NANDN U21 ( .A(A[10]), .B(n23), .Z(n22) );
  NANDN U22 ( .A(n23), .B(A[10]), .Z(n20) );
  XOR U23 ( .A(n23), .B(n24), .Z(SUM[10]) );
  XNOR U24 ( .A(B[10]), .B(A[10]), .Z(n24) );
  AND U25 ( .A(n25), .B(n26), .Z(n23) );
  NAND U26 ( .A(B[9]), .B(n27), .Z(n26) );
  OR U27 ( .A(n2), .B(A[9]), .Z(n27) );
  NAND U28 ( .A(A[9]), .B(n2), .Z(n25) );
  NAND U29 ( .A(n28), .B(n29), .Z(n2) );
  NAND U30 ( .A(B[8]), .B(n30), .Z(n29) );
  NANDN U31 ( .A(A[8]), .B(n4), .Z(n30) );
  NANDN U32 ( .A(n4), .B(A[8]), .Z(n28) );
  AND U33 ( .A(n31), .B(n32), .Z(n4) );
  NAND U34 ( .A(B[7]), .B(n33), .Z(n32) );
  NANDN U35 ( .A(A[7]), .B(n6), .Z(n33) );
  NANDN U36 ( .A(n6), .B(A[7]), .Z(n31) );
  AND U37 ( .A(n34), .B(n35), .Z(n6) );
  NAND U38 ( .A(B[6]), .B(n36), .Z(n35) );
  NANDN U39 ( .A(A[6]), .B(n8), .Z(n36) );
  NANDN U40 ( .A(n8), .B(A[6]), .Z(n34) );
  AND U41 ( .A(n37), .B(n38), .Z(n8) );
  NAND U42 ( .A(B[5]), .B(n39), .Z(n38) );
  NANDN U43 ( .A(A[5]), .B(n10), .Z(n39) );
  NANDN U44 ( .A(n10), .B(A[5]), .Z(n37) );
  AND U45 ( .A(n40), .B(n41), .Z(n10) );
  NAND U46 ( .A(B[4]), .B(n42), .Z(n41) );
  NANDN U47 ( .A(A[4]), .B(n12), .Z(n42) );
  NANDN U48 ( .A(n12), .B(A[4]), .Z(n40) );
  AND U49 ( .A(n43), .B(n44), .Z(n12) );
  NAND U50 ( .A(B[3]), .B(n45), .Z(n44) );
  NANDN U51 ( .A(A[3]), .B(n14), .Z(n45) );
  NANDN U52 ( .A(n14), .B(A[3]), .Z(n43) );
  AND U53 ( .A(n46), .B(n47), .Z(n14) );
  NAND U54 ( .A(B[2]), .B(n48), .Z(n47) );
  NANDN U55 ( .A(A[2]), .B(n16), .Z(n48) );
  NANDN U56 ( .A(n16), .B(A[2]), .Z(n46) );
  AND U57 ( .A(n49), .B(n50), .Z(n16) );
  NAND U58 ( .A(B[1]), .B(n51), .Z(n50) );
  OR U59 ( .A(n18), .B(A[1]), .Z(n51) );
  NAND U60 ( .A(A[1]), .B(n18), .Z(n49) );
  AND U61 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U62 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_5 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49;

  AND U1 ( .A(B[10]), .B(n2), .Z(SUM[11]) );
  IV U2 ( .A(n22), .Z(n2) );
  IV U3 ( .A(B[10]), .Z(n3) );
  XNOR U4 ( .A(n4), .B(n5), .Z(SUM[9]) );
  XNOR U5 ( .A(B[9]), .B(A[9]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[8]) );
  XNOR U7 ( .A(B[8]), .B(A[8]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[7]) );
  XNOR U9 ( .A(B[7]), .B(A[7]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[6]) );
  XNOR U11 ( .A(B[6]), .B(A[6]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[5]) );
  XNOR U13 ( .A(B[5]), .B(A[5]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[4]) );
  XNOR U15 ( .A(B[4]), .B(A[4]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[3]) );
  XNOR U17 ( .A(B[3]), .B(A[3]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[2]) );
  XNOR U19 ( .A(B[2]), .B(A[2]), .Z(n19) );
  XOR U20 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U21 ( .A(B[1]), .B(A[1]), .Z(n21) );
  XOR U22 ( .A(n22), .B(n3), .Z(SUM[10]) );
  AND U23 ( .A(n23), .B(n24), .Z(n22) );
  NAND U24 ( .A(B[9]), .B(n25), .Z(n24) );
  OR U25 ( .A(n4), .B(A[9]), .Z(n25) );
  NAND U26 ( .A(A[9]), .B(n4), .Z(n23) );
  NAND U27 ( .A(n26), .B(n27), .Z(n4) );
  NAND U28 ( .A(B[8]), .B(n28), .Z(n27) );
  NANDN U29 ( .A(A[8]), .B(n6), .Z(n28) );
  NANDN U30 ( .A(n6), .B(A[8]), .Z(n26) );
  AND U31 ( .A(n29), .B(n30), .Z(n6) );
  NAND U32 ( .A(B[7]), .B(n31), .Z(n30) );
  NANDN U33 ( .A(A[7]), .B(n8), .Z(n31) );
  NANDN U34 ( .A(n8), .B(A[7]), .Z(n29) );
  AND U35 ( .A(n32), .B(n33), .Z(n8) );
  NAND U36 ( .A(B[6]), .B(n34), .Z(n33) );
  NANDN U37 ( .A(A[6]), .B(n10), .Z(n34) );
  NANDN U38 ( .A(n10), .B(A[6]), .Z(n32) );
  AND U39 ( .A(n35), .B(n36), .Z(n10) );
  NAND U40 ( .A(B[5]), .B(n37), .Z(n36) );
  NANDN U41 ( .A(A[5]), .B(n12), .Z(n37) );
  NANDN U42 ( .A(n12), .B(A[5]), .Z(n35) );
  AND U43 ( .A(n38), .B(n39), .Z(n12) );
  NAND U44 ( .A(B[4]), .B(n40), .Z(n39) );
  NANDN U45 ( .A(A[4]), .B(n14), .Z(n40) );
  NANDN U46 ( .A(n14), .B(A[4]), .Z(n38) );
  AND U47 ( .A(n41), .B(n42), .Z(n14) );
  NAND U48 ( .A(B[3]), .B(n43), .Z(n42) );
  NANDN U49 ( .A(A[3]), .B(n16), .Z(n43) );
  NANDN U50 ( .A(n16), .B(A[3]), .Z(n41) );
  AND U51 ( .A(n44), .B(n45), .Z(n16) );
  NAND U52 ( .A(B[2]), .B(n46), .Z(n45) );
  NANDN U53 ( .A(A[2]), .B(n18), .Z(n46) );
  NANDN U54 ( .A(n18), .B(A[2]), .Z(n44) );
  AND U55 ( .A(n47), .B(n48), .Z(n18) );
  NAND U56 ( .A(B[1]), .B(n49), .Z(n48) );
  OR U57 ( .A(n20), .B(A[1]), .Z(n49) );
  NAND U58 ( .A(A[1]), .B(n20), .Z(n47) );
  AND U59 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U60 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_6 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46;

  NAND U1 ( .A(n20), .B(n21), .Z(SUM[10]) );
  XNOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  NAND U20 ( .A(B[9]), .B(n22), .Z(n21) );
  OR U21 ( .A(n2), .B(A[9]), .Z(n22) );
  NAND U22 ( .A(A[9]), .B(n2), .Z(n20) );
  NAND U23 ( .A(n23), .B(n24), .Z(n2) );
  NAND U24 ( .A(B[8]), .B(n25), .Z(n24) );
  NANDN U25 ( .A(A[8]), .B(n4), .Z(n25) );
  NANDN U26 ( .A(n4), .B(A[8]), .Z(n23) );
  AND U27 ( .A(n26), .B(n27), .Z(n4) );
  NAND U28 ( .A(B[7]), .B(n28), .Z(n27) );
  NANDN U29 ( .A(A[7]), .B(n6), .Z(n28) );
  NANDN U30 ( .A(n6), .B(A[7]), .Z(n26) );
  AND U31 ( .A(n29), .B(n30), .Z(n6) );
  NAND U32 ( .A(B[6]), .B(n31), .Z(n30) );
  NANDN U33 ( .A(A[6]), .B(n8), .Z(n31) );
  NANDN U34 ( .A(n8), .B(A[6]), .Z(n29) );
  AND U35 ( .A(n32), .B(n33), .Z(n8) );
  NAND U36 ( .A(B[5]), .B(n34), .Z(n33) );
  NANDN U37 ( .A(A[5]), .B(n10), .Z(n34) );
  NANDN U38 ( .A(n10), .B(A[5]), .Z(n32) );
  AND U39 ( .A(n35), .B(n36), .Z(n10) );
  NAND U40 ( .A(B[4]), .B(n37), .Z(n36) );
  NANDN U41 ( .A(A[4]), .B(n12), .Z(n37) );
  NANDN U42 ( .A(n12), .B(A[4]), .Z(n35) );
  AND U43 ( .A(n38), .B(n39), .Z(n12) );
  NAND U44 ( .A(B[3]), .B(n40), .Z(n39) );
  NANDN U45 ( .A(A[3]), .B(n14), .Z(n40) );
  NANDN U46 ( .A(n14), .B(A[3]), .Z(n38) );
  AND U47 ( .A(n41), .B(n42), .Z(n14) );
  NAND U48 ( .A(B[2]), .B(n43), .Z(n42) );
  NANDN U49 ( .A(A[2]), .B(n16), .Z(n43) );
  NANDN U50 ( .A(n16), .B(A[2]), .Z(n41) );
  AND U51 ( .A(n44), .B(n45), .Z(n16) );
  NAND U52 ( .A(B[1]), .B(n46), .Z(n45) );
  OR U53 ( .A(n18), .B(A[1]), .Z(n46) );
  NAND U54 ( .A(A[1]), .B(n18), .Z(n44) );
  AND U55 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U56 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_7 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46;

  NAND U1 ( .A(n20), .B(n21), .Z(SUM[10]) );
  XNOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  NAND U20 ( .A(B[9]), .B(n22), .Z(n21) );
  OR U21 ( .A(n2), .B(A[9]), .Z(n22) );
  NAND U22 ( .A(A[9]), .B(n2), .Z(n20) );
  NAND U23 ( .A(n23), .B(n24), .Z(n2) );
  NAND U24 ( .A(B[8]), .B(n25), .Z(n24) );
  NANDN U25 ( .A(A[8]), .B(n4), .Z(n25) );
  NANDN U26 ( .A(n4), .B(A[8]), .Z(n23) );
  AND U27 ( .A(n26), .B(n27), .Z(n4) );
  NAND U28 ( .A(B[7]), .B(n28), .Z(n27) );
  NANDN U29 ( .A(A[7]), .B(n6), .Z(n28) );
  NANDN U30 ( .A(n6), .B(A[7]), .Z(n26) );
  AND U31 ( .A(n29), .B(n30), .Z(n6) );
  NAND U32 ( .A(B[6]), .B(n31), .Z(n30) );
  NANDN U33 ( .A(A[6]), .B(n8), .Z(n31) );
  NANDN U34 ( .A(n8), .B(A[6]), .Z(n29) );
  AND U35 ( .A(n32), .B(n33), .Z(n8) );
  NAND U36 ( .A(B[5]), .B(n34), .Z(n33) );
  NANDN U37 ( .A(A[5]), .B(n10), .Z(n34) );
  NANDN U38 ( .A(n10), .B(A[5]), .Z(n32) );
  AND U39 ( .A(n35), .B(n36), .Z(n10) );
  NAND U40 ( .A(B[4]), .B(n37), .Z(n36) );
  NANDN U41 ( .A(A[4]), .B(n12), .Z(n37) );
  NANDN U42 ( .A(n12), .B(A[4]), .Z(n35) );
  AND U43 ( .A(n38), .B(n39), .Z(n12) );
  NAND U44 ( .A(B[3]), .B(n40), .Z(n39) );
  NANDN U45 ( .A(A[3]), .B(n14), .Z(n40) );
  NANDN U46 ( .A(n14), .B(A[3]), .Z(n38) );
  AND U47 ( .A(n41), .B(n42), .Z(n14) );
  NAND U48 ( .A(B[2]), .B(n43), .Z(n42) );
  NANDN U49 ( .A(A[2]), .B(n16), .Z(n43) );
  NANDN U50 ( .A(n16), .B(A[2]), .Z(n41) );
  AND U51 ( .A(n44), .B(n45), .Z(n16) );
  NAND U52 ( .A(B[1]), .B(n46), .Z(n45) );
  OR U53 ( .A(n18), .B(A[1]), .Z(n46) );
  NAND U54 ( .A(A[1]), .B(n18), .Z(n44) );
  AND U55 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U56 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_8 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46;

  NAND U1 ( .A(n20), .B(n21), .Z(SUM[10]) );
  XNOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  NAND U20 ( .A(B[9]), .B(n22), .Z(n21) );
  OR U21 ( .A(n2), .B(A[9]), .Z(n22) );
  NAND U22 ( .A(A[9]), .B(n2), .Z(n20) );
  NAND U23 ( .A(n23), .B(n24), .Z(n2) );
  NAND U24 ( .A(B[8]), .B(n25), .Z(n24) );
  NANDN U25 ( .A(A[8]), .B(n4), .Z(n25) );
  NANDN U26 ( .A(n4), .B(A[8]), .Z(n23) );
  AND U27 ( .A(n26), .B(n27), .Z(n4) );
  NAND U28 ( .A(B[7]), .B(n28), .Z(n27) );
  NANDN U29 ( .A(A[7]), .B(n6), .Z(n28) );
  NANDN U30 ( .A(n6), .B(A[7]), .Z(n26) );
  AND U31 ( .A(n29), .B(n30), .Z(n6) );
  NAND U32 ( .A(B[6]), .B(n31), .Z(n30) );
  NANDN U33 ( .A(A[6]), .B(n8), .Z(n31) );
  NANDN U34 ( .A(n8), .B(A[6]), .Z(n29) );
  AND U35 ( .A(n32), .B(n33), .Z(n8) );
  NAND U36 ( .A(B[5]), .B(n34), .Z(n33) );
  NANDN U37 ( .A(A[5]), .B(n10), .Z(n34) );
  NANDN U38 ( .A(n10), .B(A[5]), .Z(n32) );
  AND U39 ( .A(n35), .B(n36), .Z(n10) );
  NAND U40 ( .A(B[4]), .B(n37), .Z(n36) );
  NANDN U41 ( .A(A[4]), .B(n12), .Z(n37) );
  NANDN U42 ( .A(n12), .B(A[4]), .Z(n35) );
  AND U43 ( .A(n38), .B(n39), .Z(n12) );
  NAND U44 ( .A(B[3]), .B(n40), .Z(n39) );
  NANDN U45 ( .A(A[3]), .B(n14), .Z(n40) );
  NANDN U46 ( .A(n14), .B(A[3]), .Z(n38) );
  AND U47 ( .A(n41), .B(n42), .Z(n14) );
  NAND U48 ( .A(B[2]), .B(n43), .Z(n42) );
  NANDN U49 ( .A(A[2]), .B(n16), .Z(n43) );
  NANDN U50 ( .A(n16), .B(A[2]), .Z(n41) );
  AND U51 ( .A(n44), .B(n45), .Z(n16) );
  NAND U52 ( .A(B[1]), .B(n46), .Z(n45) );
  OR U53 ( .A(n18), .B(A[1]), .Z(n46) );
  NAND U54 ( .A(A[1]), .B(n18), .Z(n44) );
  AND U55 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U56 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_9 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46;

  NAND U1 ( .A(n20), .B(n21), .Z(SUM[10]) );
  XNOR U2 ( .A(n2), .B(n3), .Z(SUM[9]) );
  XNOR U3 ( .A(B[9]), .B(A[9]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n15) );
  XOR U16 ( .A(n16), .B(n17), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n17) );
  XOR U18 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n19) );
  NAND U20 ( .A(B[9]), .B(n22), .Z(n21) );
  OR U21 ( .A(n2), .B(A[9]), .Z(n22) );
  NAND U22 ( .A(A[9]), .B(n2), .Z(n20) );
  NAND U23 ( .A(n23), .B(n24), .Z(n2) );
  NAND U24 ( .A(B[8]), .B(n25), .Z(n24) );
  NANDN U25 ( .A(A[8]), .B(n4), .Z(n25) );
  NANDN U26 ( .A(n4), .B(A[8]), .Z(n23) );
  AND U27 ( .A(n26), .B(n27), .Z(n4) );
  NAND U28 ( .A(B[7]), .B(n28), .Z(n27) );
  NANDN U29 ( .A(A[7]), .B(n6), .Z(n28) );
  NANDN U30 ( .A(n6), .B(A[7]), .Z(n26) );
  AND U31 ( .A(n29), .B(n30), .Z(n6) );
  NAND U32 ( .A(B[6]), .B(n31), .Z(n30) );
  NANDN U33 ( .A(A[6]), .B(n8), .Z(n31) );
  NANDN U34 ( .A(n8), .B(A[6]), .Z(n29) );
  AND U35 ( .A(n32), .B(n33), .Z(n8) );
  NAND U36 ( .A(B[5]), .B(n34), .Z(n33) );
  NANDN U37 ( .A(A[5]), .B(n10), .Z(n34) );
  NANDN U38 ( .A(n10), .B(A[5]), .Z(n32) );
  AND U39 ( .A(n35), .B(n36), .Z(n10) );
  NAND U40 ( .A(B[4]), .B(n37), .Z(n36) );
  NANDN U41 ( .A(A[4]), .B(n12), .Z(n37) );
  NANDN U42 ( .A(n12), .B(A[4]), .Z(n35) );
  AND U43 ( .A(n38), .B(n39), .Z(n12) );
  NAND U44 ( .A(B[3]), .B(n40), .Z(n39) );
  NANDN U45 ( .A(A[3]), .B(n14), .Z(n40) );
  NANDN U46 ( .A(n14), .B(A[3]), .Z(n38) );
  AND U47 ( .A(n41), .B(n42), .Z(n14) );
  NAND U48 ( .A(B[2]), .B(n43), .Z(n42) );
  NANDN U49 ( .A(A[2]), .B(n16), .Z(n43) );
  NANDN U50 ( .A(n16), .B(A[2]), .Z(n41) );
  AND U51 ( .A(n44), .B(n45), .Z(n16) );
  NAND U52 ( .A(B[1]), .B(n46), .Z(n45) );
  OR U53 ( .A(n18), .B(A[1]), .Z(n46) );
  NAND U54 ( .A(A[1]), .B(n18), .Z(n44) );
  AND U55 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U56 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_10 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43;

  AND U1 ( .A(B[9]), .B(n19), .Z(SUM[10]) );
  IV U2 ( .A(B[9]), .Z(n2) );
  XNOR U3 ( .A(n19), .B(n2), .Z(SUM[9]) );
  XOR U4 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U5 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U6 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U7 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U8 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U9 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U10 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U11 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U12 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U13 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U14 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U15 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U16 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U17 ( .A(B[2]), .B(A[2]), .Z(n16) );
  XOR U18 ( .A(n17), .B(n18), .Z(SUM[1]) );
  XOR U19 ( .A(B[1]), .B(A[1]), .Z(n18) );
  NAND U20 ( .A(n20), .B(n21), .Z(n19) );
  NAND U21 ( .A(B[8]), .B(n22), .Z(n21) );
  NANDN U22 ( .A(A[8]), .B(n3), .Z(n22) );
  NANDN U23 ( .A(n3), .B(A[8]), .Z(n20) );
  AND U24 ( .A(n23), .B(n24), .Z(n3) );
  NAND U25 ( .A(B[7]), .B(n25), .Z(n24) );
  NANDN U26 ( .A(A[7]), .B(n5), .Z(n25) );
  NANDN U27 ( .A(n5), .B(A[7]), .Z(n23) );
  AND U28 ( .A(n26), .B(n27), .Z(n5) );
  NAND U29 ( .A(B[6]), .B(n28), .Z(n27) );
  NANDN U30 ( .A(A[6]), .B(n7), .Z(n28) );
  NANDN U31 ( .A(n7), .B(A[6]), .Z(n26) );
  AND U32 ( .A(n29), .B(n30), .Z(n7) );
  NAND U33 ( .A(B[5]), .B(n31), .Z(n30) );
  NANDN U34 ( .A(A[5]), .B(n9), .Z(n31) );
  NANDN U35 ( .A(n9), .B(A[5]), .Z(n29) );
  AND U36 ( .A(n32), .B(n33), .Z(n9) );
  NAND U37 ( .A(B[4]), .B(n34), .Z(n33) );
  NANDN U38 ( .A(A[4]), .B(n11), .Z(n34) );
  NANDN U39 ( .A(n11), .B(A[4]), .Z(n32) );
  AND U40 ( .A(n35), .B(n36), .Z(n11) );
  NAND U41 ( .A(B[3]), .B(n37), .Z(n36) );
  NANDN U42 ( .A(A[3]), .B(n13), .Z(n37) );
  NANDN U43 ( .A(n13), .B(A[3]), .Z(n35) );
  AND U44 ( .A(n38), .B(n39), .Z(n13) );
  NAND U45 ( .A(B[2]), .B(n40), .Z(n39) );
  NANDN U46 ( .A(A[2]), .B(n15), .Z(n40) );
  NANDN U47 ( .A(n15), .B(A[2]), .Z(n38) );
  AND U48 ( .A(n41), .B(n42), .Z(n15) );
  NAND U49 ( .A(B[1]), .B(n43), .Z(n42) );
  OR U50 ( .A(n17), .B(A[1]), .Z(n43) );
  NAND U51 ( .A(A[1]), .B(n17), .Z(n41) );
  AND U52 ( .A(B[0]), .B(A[0]), .Z(n17) );
  XOR U53 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_11 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[8]) );
  XNOR U2 ( .A(B[8]), .B(A[8]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[7]) );
  XNOR U4 ( .A(B[7]), .B(A[7]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[6]) );
  XNOR U6 ( .A(B[6]), .B(A[6]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[5]) );
  XNOR U8 ( .A(B[5]), .B(A[5]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[4]) );
  XNOR U10 ( .A(B[4]), .B(A[4]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[2]) );
  XNOR U14 ( .A(B[2]), .B(A[2]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[1]) );
  XOR U16 ( .A(B[1]), .B(A[1]), .Z(n16) );
  NAND U17 ( .A(n17), .B(n18), .Z(SUM[9]) );
  NAND U18 ( .A(B[8]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[8]), .B(n1), .Z(n19) );
  NANDN U20 ( .A(n1), .B(A[8]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n1) );
  NAND U22 ( .A(B[7]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[7]), .B(n3), .Z(n22) );
  NANDN U24 ( .A(n3), .B(A[7]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n3) );
  NAND U26 ( .A(B[6]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[6]), .B(n5), .Z(n25) );
  NANDN U28 ( .A(n5), .B(A[6]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n5) );
  NAND U30 ( .A(B[5]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[5]), .B(n7), .Z(n28) );
  NANDN U32 ( .A(n7), .B(A[5]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n7) );
  NAND U34 ( .A(B[4]), .B(n31), .Z(n30) );
  NANDN U35 ( .A(A[4]), .B(n9), .Z(n31) );
  NANDN U36 ( .A(n9), .B(A[4]), .Z(n29) );
  AND U37 ( .A(n32), .B(n33), .Z(n9) );
  NAND U38 ( .A(B[3]), .B(n34), .Z(n33) );
  NANDN U39 ( .A(A[3]), .B(n11), .Z(n34) );
  NANDN U40 ( .A(n11), .B(A[3]), .Z(n32) );
  AND U41 ( .A(n35), .B(n36), .Z(n11) );
  NAND U42 ( .A(B[2]), .B(n37), .Z(n36) );
  NANDN U43 ( .A(A[2]), .B(n13), .Z(n37) );
  NANDN U44 ( .A(n13), .B(A[2]), .Z(n35) );
  AND U45 ( .A(n38), .B(n39), .Z(n13) );
  NAND U46 ( .A(B[1]), .B(n40), .Z(n39) );
  OR U47 ( .A(n15), .B(A[1]), .Z(n40) );
  NAND U48 ( .A(A[1]), .B(n15), .Z(n38) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n15) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_12 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[8]) );
  XNOR U2 ( .A(B[8]), .B(A[8]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[7]) );
  XNOR U4 ( .A(B[7]), .B(A[7]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[6]) );
  XNOR U6 ( .A(B[6]), .B(A[6]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[5]) );
  XNOR U8 ( .A(B[5]), .B(A[5]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[4]) );
  XNOR U10 ( .A(B[4]), .B(A[4]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[2]) );
  XNOR U14 ( .A(B[2]), .B(A[2]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[1]) );
  XOR U16 ( .A(B[1]), .B(A[1]), .Z(n16) );
  NAND U17 ( .A(n17), .B(n18), .Z(SUM[9]) );
  NAND U18 ( .A(B[8]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[8]), .B(n1), .Z(n19) );
  NANDN U20 ( .A(n1), .B(A[8]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n1) );
  NAND U22 ( .A(B[7]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[7]), .B(n3), .Z(n22) );
  NANDN U24 ( .A(n3), .B(A[7]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n3) );
  NAND U26 ( .A(B[6]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[6]), .B(n5), .Z(n25) );
  NANDN U28 ( .A(n5), .B(A[6]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n5) );
  NAND U30 ( .A(B[5]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[5]), .B(n7), .Z(n28) );
  NANDN U32 ( .A(n7), .B(A[5]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n7) );
  NAND U34 ( .A(B[4]), .B(n31), .Z(n30) );
  NANDN U35 ( .A(A[4]), .B(n9), .Z(n31) );
  NANDN U36 ( .A(n9), .B(A[4]), .Z(n29) );
  AND U37 ( .A(n32), .B(n33), .Z(n9) );
  NAND U38 ( .A(B[3]), .B(n34), .Z(n33) );
  NANDN U39 ( .A(A[3]), .B(n11), .Z(n34) );
  NANDN U40 ( .A(n11), .B(A[3]), .Z(n32) );
  AND U41 ( .A(n35), .B(n36), .Z(n11) );
  NAND U42 ( .A(B[2]), .B(n37), .Z(n36) );
  NANDN U43 ( .A(A[2]), .B(n13), .Z(n37) );
  NANDN U44 ( .A(n13), .B(A[2]), .Z(n35) );
  AND U45 ( .A(n38), .B(n39), .Z(n13) );
  NAND U46 ( .A(B[1]), .B(n40), .Z(n39) );
  OR U47 ( .A(n15), .B(A[1]), .Z(n40) );
  NAND U48 ( .A(A[1]), .B(n15), .Z(n38) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n15) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_13 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[8]) );
  XNOR U2 ( .A(B[8]), .B(A[8]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[7]) );
  XNOR U4 ( .A(B[7]), .B(A[7]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[6]) );
  XNOR U6 ( .A(B[6]), .B(A[6]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[5]) );
  XNOR U8 ( .A(B[5]), .B(A[5]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[4]) );
  XNOR U10 ( .A(B[4]), .B(A[4]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[2]) );
  XNOR U14 ( .A(B[2]), .B(A[2]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[1]) );
  XOR U16 ( .A(B[1]), .B(A[1]), .Z(n16) );
  NAND U17 ( .A(n17), .B(n18), .Z(SUM[9]) );
  NAND U18 ( .A(B[8]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[8]), .B(n1), .Z(n19) );
  NANDN U20 ( .A(n1), .B(A[8]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n1) );
  NAND U22 ( .A(B[7]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[7]), .B(n3), .Z(n22) );
  NANDN U24 ( .A(n3), .B(A[7]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n3) );
  NAND U26 ( .A(B[6]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[6]), .B(n5), .Z(n25) );
  NANDN U28 ( .A(n5), .B(A[6]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n5) );
  NAND U30 ( .A(B[5]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[5]), .B(n7), .Z(n28) );
  NANDN U32 ( .A(n7), .B(A[5]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n7) );
  NAND U34 ( .A(B[4]), .B(n31), .Z(n30) );
  NANDN U35 ( .A(A[4]), .B(n9), .Z(n31) );
  NANDN U36 ( .A(n9), .B(A[4]), .Z(n29) );
  AND U37 ( .A(n32), .B(n33), .Z(n9) );
  NAND U38 ( .A(B[3]), .B(n34), .Z(n33) );
  NANDN U39 ( .A(A[3]), .B(n11), .Z(n34) );
  NANDN U40 ( .A(n11), .B(A[3]), .Z(n32) );
  AND U41 ( .A(n35), .B(n36), .Z(n11) );
  NAND U42 ( .A(B[2]), .B(n37), .Z(n36) );
  NANDN U43 ( .A(A[2]), .B(n13), .Z(n37) );
  NANDN U44 ( .A(n13), .B(A[2]), .Z(n35) );
  AND U45 ( .A(n38), .B(n39), .Z(n13) );
  NAND U46 ( .A(B[1]), .B(n40), .Z(n39) );
  OR U47 ( .A(n15), .B(A[1]), .Z(n40) );
  NAND U48 ( .A(A[1]), .B(n15), .Z(n38) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n15) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_14 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[8]) );
  XNOR U2 ( .A(B[8]), .B(A[8]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[7]) );
  XNOR U4 ( .A(B[7]), .B(A[7]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[6]) );
  XNOR U6 ( .A(B[6]), .B(A[6]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[5]) );
  XNOR U8 ( .A(B[5]), .B(A[5]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[4]) );
  XNOR U10 ( .A(B[4]), .B(A[4]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[2]) );
  XNOR U14 ( .A(B[2]), .B(A[2]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[1]) );
  XOR U16 ( .A(B[1]), .B(A[1]), .Z(n16) );
  NAND U17 ( .A(n17), .B(n18), .Z(SUM[9]) );
  NAND U18 ( .A(B[8]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[8]), .B(n1), .Z(n19) );
  NANDN U20 ( .A(n1), .B(A[8]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n1) );
  NAND U22 ( .A(B[7]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[7]), .B(n3), .Z(n22) );
  NANDN U24 ( .A(n3), .B(A[7]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n3) );
  NAND U26 ( .A(B[6]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[6]), .B(n5), .Z(n25) );
  NANDN U28 ( .A(n5), .B(A[6]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n5) );
  NAND U30 ( .A(B[5]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[5]), .B(n7), .Z(n28) );
  NANDN U32 ( .A(n7), .B(A[5]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n7) );
  NAND U34 ( .A(B[4]), .B(n31), .Z(n30) );
  NANDN U35 ( .A(A[4]), .B(n9), .Z(n31) );
  NANDN U36 ( .A(n9), .B(A[4]), .Z(n29) );
  AND U37 ( .A(n32), .B(n33), .Z(n9) );
  NAND U38 ( .A(B[3]), .B(n34), .Z(n33) );
  NANDN U39 ( .A(A[3]), .B(n11), .Z(n34) );
  NANDN U40 ( .A(n11), .B(A[3]), .Z(n32) );
  AND U41 ( .A(n35), .B(n36), .Z(n11) );
  NAND U42 ( .A(B[2]), .B(n37), .Z(n36) );
  NANDN U43 ( .A(A[2]), .B(n13), .Z(n37) );
  NANDN U44 ( .A(n13), .B(A[2]), .Z(n35) );
  AND U45 ( .A(n38), .B(n39), .Z(n13) );
  NAND U46 ( .A(B[1]), .B(n40), .Z(n39) );
  OR U47 ( .A(n15), .B(A[1]), .Z(n40) );
  NAND U48 ( .A(A[1]), .B(n15), .Z(n38) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n15) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_15 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[8]) );
  XNOR U2 ( .A(B[8]), .B(A[8]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[7]) );
  XNOR U4 ( .A(B[7]), .B(A[7]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[6]) );
  XNOR U6 ( .A(B[6]), .B(A[6]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[5]) );
  XNOR U8 ( .A(B[5]), .B(A[5]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[4]) );
  XNOR U10 ( .A(B[4]), .B(A[4]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[2]) );
  XNOR U14 ( .A(B[2]), .B(A[2]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[1]) );
  XOR U16 ( .A(B[1]), .B(A[1]), .Z(n16) );
  NAND U17 ( .A(n17), .B(n18), .Z(SUM[9]) );
  NAND U18 ( .A(B[8]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[8]), .B(n1), .Z(n19) );
  NANDN U20 ( .A(n1), .B(A[8]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n1) );
  NAND U22 ( .A(B[7]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[7]), .B(n3), .Z(n22) );
  NANDN U24 ( .A(n3), .B(A[7]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n3) );
  NAND U26 ( .A(B[6]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[6]), .B(n5), .Z(n25) );
  NANDN U28 ( .A(n5), .B(A[6]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n5) );
  NAND U30 ( .A(B[5]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[5]), .B(n7), .Z(n28) );
  NANDN U32 ( .A(n7), .B(A[5]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n7) );
  NAND U34 ( .A(B[4]), .B(n31), .Z(n30) );
  NANDN U35 ( .A(A[4]), .B(n9), .Z(n31) );
  NANDN U36 ( .A(n9), .B(A[4]), .Z(n29) );
  AND U37 ( .A(n32), .B(n33), .Z(n9) );
  NAND U38 ( .A(B[3]), .B(n34), .Z(n33) );
  NANDN U39 ( .A(A[3]), .B(n11), .Z(n34) );
  NANDN U40 ( .A(n11), .B(A[3]), .Z(n32) );
  AND U41 ( .A(n35), .B(n36), .Z(n11) );
  NAND U42 ( .A(B[2]), .B(n37), .Z(n36) );
  NANDN U43 ( .A(A[2]), .B(n13), .Z(n37) );
  NANDN U44 ( .A(n13), .B(A[2]), .Z(n35) );
  AND U45 ( .A(n38), .B(n39), .Z(n13) );
  NAND U46 ( .A(B[1]), .B(n40), .Z(n39) );
  OR U47 ( .A(n15), .B(A[1]), .Z(n40) );
  NAND U48 ( .A(A[1]), .B(n15), .Z(n38) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n15) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_16 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[8]) );
  XNOR U2 ( .A(B[8]), .B(A[8]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[7]) );
  XNOR U4 ( .A(B[7]), .B(A[7]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[6]) );
  XNOR U6 ( .A(B[6]), .B(A[6]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[5]) );
  XNOR U8 ( .A(B[5]), .B(A[5]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[4]) );
  XNOR U10 ( .A(B[4]), .B(A[4]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[2]) );
  XNOR U14 ( .A(B[2]), .B(A[2]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[1]) );
  XOR U16 ( .A(B[1]), .B(A[1]), .Z(n16) );
  NAND U17 ( .A(n17), .B(n18), .Z(SUM[9]) );
  NAND U18 ( .A(B[8]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[8]), .B(n1), .Z(n19) );
  NANDN U20 ( .A(n1), .B(A[8]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n1) );
  NAND U22 ( .A(B[7]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[7]), .B(n3), .Z(n22) );
  NANDN U24 ( .A(n3), .B(A[7]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n3) );
  NAND U26 ( .A(B[6]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[6]), .B(n5), .Z(n25) );
  NANDN U28 ( .A(n5), .B(A[6]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n5) );
  NAND U30 ( .A(B[5]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[5]), .B(n7), .Z(n28) );
  NANDN U32 ( .A(n7), .B(A[5]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n7) );
  NAND U34 ( .A(B[4]), .B(n31), .Z(n30) );
  NANDN U35 ( .A(A[4]), .B(n9), .Z(n31) );
  NANDN U36 ( .A(n9), .B(A[4]), .Z(n29) );
  AND U37 ( .A(n32), .B(n33), .Z(n9) );
  NAND U38 ( .A(B[3]), .B(n34), .Z(n33) );
  NANDN U39 ( .A(A[3]), .B(n11), .Z(n34) );
  NANDN U40 ( .A(n11), .B(A[3]), .Z(n32) );
  AND U41 ( .A(n35), .B(n36), .Z(n11) );
  NAND U42 ( .A(B[2]), .B(n37), .Z(n36) );
  NANDN U43 ( .A(A[2]), .B(n13), .Z(n37) );
  NANDN U44 ( .A(n13), .B(A[2]), .Z(n35) );
  AND U45 ( .A(n38), .B(n39), .Z(n13) );
  NAND U46 ( .A(B[1]), .B(n40), .Z(n39) );
  OR U47 ( .A(n15), .B(A[1]), .Z(n40) );
  NAND U48 ( .A(A[1]), .B(n15), .Z(n38) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n15) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_17 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[8]) );
  XNOR U2 ( .A(B[8]), .B(A[8]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[7]) );
  XNOR U4 ( .A(B[7]), .B(A[7]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[6]) );
  XNOR U6 ( .A(B[6]), .B(A[6]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[5]) );
  XNOR U8 ( .A(B[5]), .B(A[5]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[4]) );
  XNOR U10 ( .A(B[4]), .B(A[4]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[2]) );
  XNOR U14 ( .A(B[2]), .B(A[2]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[1]) );
  XOR U16 ( .A(B[1]), .B(A[1]), .Z(n16) );
  NAND U17 ( .A(n17), .B(n18), .Z(SUM[9]) );
  NAND U18 ( .A(B[8]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[8]), .B(n1), .Z(n19) );
  NANDN U20 ( .A(n1), .B(A[8]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n1) );
  NAND U22 ( .A(B[7]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[7]), .B(n3), .Z(n22) );
  NANDN U24 ( .A(n3), .B(A[7]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n3) );
  NAND U26 ( .A(B[6]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[6]), .B(n5), .Z(n25) );
  NANDN U28 ( .A(n5), .B(A[6]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n5) );
  NAND U30 ( .A(B[5]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[5]), .B(n7), .Z(n28) );
  NANDN U32 ( .A(n7), .B(A[5]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n7) );
  NAND U34 ( .A(B[4]), .B(n31), .Z(n30) );
  NANDN U35 ( .A(A[4]), .B(n9), .Z(n31) );
  NANDN U36 ( .A(n9), .B(A[4]), .Z(n29) );
  AND U37 ( .A(n32), .B(n33), .Z(n9) );
  NAND U38 ( .A(B[3]), .B(n34), .Z(n33) );
  NANDN U39 ( .A(A[3]), .B(n11), .Z(n34) );
  NANDN U40 ( .A(n11), .B(A[3]), .Z(n32) );
  AND U41 ( .A(n35), .B(n36), .Z(n11) );
  NAND U42 ( .A(B[2]), .B(n37), .Z(n36) );
  NANDN U43 ( .A(A[2]), .B(n13), .Z(n37) );
  NANDN U44 ( .A(n13), .B(A[2]), .Z(n35) );
  AND U45 ( .A(n38), .B(n39), .Z(n13) );
  NAND U46 ( .A(B[1]), .B(n40), .Z(n39) );
  OR U47 ( .A(n15), .B(A[1]), .Z(n40) );
  NAND U48 ( .A(A[1]), .B(n15), .Z(n38) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n15) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_18 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[8]) );
  XNOR U2 ( .A(B[8]), .B(A[8]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[7]) );
  XNOR U4 ( .A(B[7]), .B(A[7]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[6]) );
  XNOR U6 ( .A(B[6]), .B(A[6]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[5]) );
  XNOR U8 ( .A(B[5]), .B(A[5]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[4]) );
  XNOR U10 ( .A(B[4]), .B(A[4]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[2]) );
  XNOR U14 ( .A(B[2]), .B(A[2]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[1]) );
  XOR U16 ( .A(B[1]), .B(A[1]), .Z(n16) );
  NAND U17 ( .A(n17), .B(n18), .Z(SUM[9]) );
  NAND U18 ( .A(B[8]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[8]), .B(n1), .Z(n19) );
  NANDN U20 ( .A(n1), .B(A[8]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n1) );
  NAND U22 ( .A(B[7]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[7]), .B(n3), .Z(n22) );
  NANDN U24 ( .A(n3), .B(A[7]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n3) );
  NAND U26 ( .A(B[6]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[6]), .B(n5), .Z(n25) );
  NANDN U28 ( .A(n5), .B(A[6]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n5) );
  NAND U30 ( .A(B[5]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[5]), .B(n7), .Z(n28) );
  NANDN U32 ( .A(n7), .B(A[5]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n7) );
  NAND U34 ( .A(B[4]), .B(n31), .Z(n30) );
  NANDN U35 ( .A(A[4]), .B(n9), .Z(n31) );
  NANDN U36 ( .A(n9), .B(A[4]), .Z(n29) );
  AND U37 ( .A(n32), .B(n33), .Z(n9) );
  NAND U38 ( .A(B[3]), .B(n34), .Z(n33) );
  NANDN U39 ( .A(A[3]), .B(n11), .Z(n34) );
  NANDN U40 ( .A(n11), .B(A[3]), .Z(n32) );
  AND U41 ( .A(n35), .B(n36), .Z(n11) );
  NAND U42 ( .A(B[2]), .B(n37), .Z(n36) );
  NANDN U43 ( .A(A[2]), .B(n13), .Z(n37) );
  NANDN U44 ( .A(n13), .B(A[2]), .Z(n35) );
  AND U45 ( .A(n38), .B(n39), .Z(n13) );
  NAND U46 ( .A(B[1]), .B(n40), .Z(n39) );
  OR U47 ( .A(n15), .B(A[1]), .Z(n40) );
  NAND U48 ( .A(A[1]), .B(n15), .Z(n38) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n15) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_19 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[8]) );
  XNOR U2 ( .A(B[8]), .B(A[8]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[7]) );
  XNOR U4 ( .A(B[7]), .B(A[7]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[6]) );
  XNOR U6 ( .A(B[6]), .B(A[6]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[5]) );
  XNOR U8 ( .A(B[5]), .B(A[5]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[4]) );
  XNOR U10 ( .A(B[4]), .B(A[4]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[2]) );
  XNOR U14 ( .A(B[2]), .B(A[2]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[1]) );
  XOR U16 ( .A(B[1]), .B(A[1]), .Z(n16) );
  NAND U17 ( .A(n17), .B(n18), .Z(SUM[9]) );
  NAND U18 ( .A(B[8]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[8]), .B(n1), .Z(n19) );
  NANDN U20 ( .A(n1), .B(A[8]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n1) );
  NAND U22 ( .A(B[7]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[7]), .B(n3), .Z(n22) );
  NANDN U24 ( .A(n3), .B(A[7]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n3) );
  NAND U26 ( .A(B[6]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[6]), .B(n5), .Z(n25) );
  NANDN U28 ( .A(n5), .B(A[6]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n5) );
  NAND U30 ( .A(B[5]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[5]), .B(n7), .Z(n28) );
  NANDN U32 ( .A(n7), .B(A[5]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n7) );
  NAND U34 ( .A(B[4]), .B(n31), .Z(n30) );
  NANDN U35 ( .A(A[4]), .B(n9), .Z(n31) );
  NANDN U36 ( .A(n9), .B(A[4]), .Z(n29) );
  AND U37 ( .A(n32), .B(n33), .Z(n9) );
  NAND U38 ( .A(B[3]), .B(n34), .Z(n33) );
  NANDN U39 ( .A(A[3]), .B(n11), .Z(n34) );
  NANDN U40 ( .A(n11), .B(A[3]), .Z(n32) );
  AND U41 ( .A(n35), .B(n36), .Z(n11) );
  NAND U42 ( .A(B[2]), .B(n37), .Z(n36) );
  NANDN U43 ( .A(A[2]), .B(n13), .Z(n37) );
  NANDN U44 ( .A(n13), .B(A[2]), .Z(n35) );
  AND U45 ( .A(n38), .B(n39), .Z(n13) );
  NAND U46 ( .A(B[1]), .B(n40), .Z(n39) );
  OR U47 ( .A(n15), .B(A[1]), .Z(n40) );
  NAND U48 ( .A(A[1]), .B(n15), .Z(n38) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n15) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_20 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[8]) );
  XNOR U2 ( .A(B[8]), .B(A[8]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[7]) );
  XNOR U4 ( .A(B[7]), .B(A[7]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[6]) );
  XNOR U6 ( .A(B[6]), .B(A[6]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[5]) );
  XNOR U8 ( .A(B[5]), .B(A[5]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[4]) );
  XNOR U10 ( .A(B[4]), .B(A[4]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[2]) );
  XNOR U14 ( .A(B[2]), .B(A[2]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[1]) );
  XOR U16 ( .A(B[1]), .B(A[1]), .Z(n16) );
  NAND U17 ( .A(n17), .B(n18), .Z(SUM[9]) );
  NAND U18 ( .A(B[8]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[8]), .B(n1), .Z(n19) );
  NANDN U20 ( .A(n1), .B(A[8]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n1) );
  NAND U22 ( .A(B[7]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[7]), .B(n3), .Z(n22) );
  NANDN U24 ( .A(n3), .B(A[7]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n3) );
  NAND U26 ( .A(B[6]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[6]), .B(n5), .Z(n25) );
  NANDN U28 ( .A(n5), .B(A[6]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n5) );
  NAND U30 ( .A(B[5]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[5]), .B(n7), .Z(n28) );
  NANDN U32 ( .A(n7), .B(A[5]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n7) );
  NAND U34 ( .A(B[4]), .B(n31), .Z(n30) );
  NANDN U35 ( .A(A[4]), .B(n9), .Z(n31) );
  NANDN U36 ( .A(n9), .B(A[4]), .Z(n29) );
  AND U37 ( .A(n32), .B(n33), .Z(n9) );
  NAND U38 ( .A(B[3]), .B(n34), .Z(n33) );
  NANDN U39 ( .A(A[3]), .B(n11), .Z(n34) );
  NANDN U40 ( .A(n11), .B(A[3]), .Z(n32) );
  AND U41 ( .A(n35), .B(n36), .Z(n11) );
  NAND U42 ( .A(B[2]), .B(n37), .Z(n36) );
  NANDN U43 ( .A(A[2]), .B(n13), .Z(n37) );
  NANDN U44 ( .A(n13), .B(A[2]), .Z(n35) );
  AND U45 ( .A(n38), .B(n39), .Z(n13) );
  NAND U46 ( .A(B[1]), .B(n40), .Z(n39) );
  OR U47 ( .A(n15), .B(A[1]), .Z(n40) );
  NAND U48 ( .A(A[1]), .B(n15), .Z(n38) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n15) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_21 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_22 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_23 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_24 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_25 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_26 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_27 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_28 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_29 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_30 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_31 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_32 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_33 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_34 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_35 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_36 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_37 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_38 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_39 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_40 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_41 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n16), .B(n17), .Z(SUM[8]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[7]) );
  XNOR U3 ( .A(B[7]), .B(A[7]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[6]) );
  XNOR U5 ( .A(B[6]), .B(A[6]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[5]) );
  XNOR U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U9 ( .A(B[4]), .B(A[4]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U11 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[2]) );
  XNOR U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR U14 ( .A(n14), .B(n15), .Z(SUM[1]) );
  XOR U15 ( .A(B[1]), .B(A[1]), .Z(n15) );
  NAND U16 ( .A(B[7]), .B(n18), .Z(n17) );
  NANDN U17 ( .A(A[7]), .B(n2), .Z(n18) );
  NANDN U18 ( .A(n2), .B(A[7]), .Z(n16) );
  AND U19 ( .A(n19), .B(n20), .Z(n2) );
  NAND U20 ( .A(B[6]), .B(n21), .Z(n20) );
  NANDN U21 ( .A(A[6]), .B(n4), .Z(n21) );
  NANDN U22 ( .A(n4), .B(A[6]), .Z(n19) );
  AND U23 ( .A(n22), .B(n23), .Z(n4) );
  NAND U24 ( .A(B[5]), .B(n24), .Z(n23) );
  NANDN U25 ( .A(A[5]), .B(n6), .Z(n24) );
  NANDN U26 ( .A(n6), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n25), .B(n26), .Z(n6) );
  NAND U28 ( .A(B[4]), .B(n27), .Z(n26) );
  NANDN U29 ( .A(A[4]), .B(n8), .Z(n27) );
  NANDN U30 ( .A(n8), .B(A[4]), .Z(n25) );
  AND U31 ( .A(n28), .B(n29), .Z(n8) );
  NAND U32 ( .A(B[3]), .B(n30), .Z(n29) );
  NANDN U33 ( .A(A[3]), .B(n10), .Z(n30) );
  NANDN U34 ( .A(n10), .B(A[3]), .Z(n28) );
  AND U35 ( .A(n31), .B(n32), .Z(n10) );
  NAND U36 ( .A(B[2]), .B(n33), .Z(n32) );
  NANDN U37 ( .A(A[2]), .B(n12), .Z(n33) );
  NANDN U38 ( .A(n12), .B(A[2]), .Z(n31) );
  AND U39 ( .A(n34), .B(n35), .Z(n12) );
  NAND U40 ( .A(B[1]), .B(n36), .Z(n35) );
  OR U41 ( .A(n14), .B(A[1]), .Z(n36) );
  NAND U42 ( .A(A[1]), .B(n14), .Z(n34) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n14) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_42 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_43 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_44 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_45 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_46 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_47 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_48 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_49 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_50 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_51 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_52 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_53 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_54 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_55 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_56 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_57 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_58 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_59 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_60 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_61 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_62 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_63 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_64 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_65 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_66 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_67 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_68 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_69 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_70 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_71 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_72 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_73 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_74 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_75 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_76 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_77 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_78 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_79 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_80 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_81 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_82 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n14), .B(n15), .Z(SUM[7]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[6]) );
  XNOR U3 ( .A(B[6]), .B(A[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[5]) );
  XNOR U5 ( .A(B[5]), .B(A[5]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  NAND U14 ( .A(B[6]), .B(n16), .Z(n15) );
  NANDN U15 ( .A(A[6]), .B(n2), .Z(n16) );
  NANDN U16 ( .A(n2), .B(A[6]), .Z(n14) );
  AND U17 ( .A(n17), .B(n18), .Z(n2) );
  NAND U18 ( .A(B[5]), .B(n19), .Z(n18) );
  NANDN U19 ( .A(A[5]), .B(n4), .Z(n19) );
  NANDN U20 ( .A(n4), .B(A[5]), .Z(n17) );
  AND U21 ( .A(n20), .B(n21), .Z(n4) );
  NAND U22 ( .A(B[4]), .B(n22), .Z(n21) );
  NANDN U23 ( .A(A[4]), .B(n6), .Z(n22) );
  NANDN U24 ( .A(n6), .B(A[4]), .Z(n20) );
  AND U25 ( .A(n23), .B(n24), .Z(n6) );
  NAND U26 ( .A(B[3]), .B(n25), .Z(n24) );
  NANDN U27 ( .A(A[3]), .B(n8), .Z(n25) );
  NANDN U28 ( .A(n8), .B(A[3]), .Z(n23) );
  AND U29 ( .A(n26), .B(n27), .Z(n8) );
  NAND U30 ( .A(B[2]), .B(n28), .Z(n27) );
  NANDN U31 ( .A(A[2]), .B(n10), .Z(n28) );
  NANDN U32 ( .A(n10), .B(A[2]), .Z(n26) );
  AND U33 ( .A(n29), .B(n30), .Z(n10) );
  NAND U34 ( .A(B[1]), .B(n31), .Z(n30) );
  OR U35 ( .A(n12), .B(A[1]), .Z(n31) );
  NAND U36 ( .A(A[1]), .B(n12), .Z(n29) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_83 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29;

  AND U1 ( .A(B[6]), .B(n2), .Z(SUM[7]) );
  IV U2 ( .A(n4), .Z(n2) );
  IV U3 ( .A(B[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n3), .Z(SUM[6]) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[5]) );
  XNOR U6 ( .A(B[5]), .B(A[5]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[4]) );
  XNOR U8 ( .A(B[4]), .B(A[4]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[3]) );
  XNOR U10 ( .A(B[3]), .B(A[3]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[2]) );
  XNOR U12 ( .A(B[2]), .B(A[2]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[1]) );
  XOR U14 ( .A(B[1]), .B(A[1]), .Z(n14) );
  AND U15 ( .A(n15), .B(n16), .Z(n4) );
  NAND U16 ( .A(B[5]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[5]), .B(n5), .Z(n17) );
  NANDN U18 ( .A(n5), .B(A[5]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n5) );
  NAND U20 ( .A(B[4]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[4]), .B(n7), .Z(n20) );
  NANDN U22 ( .A(n7), .B(A[4]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n7) );
  NAND U24 ( .A(B[3]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[3]), .B(n9), .Z(n23) );
  NANDN U26 ( .A(n9), .B(A[3]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n9) );
  NAND U28 ( .A(B[2]), .B(n26), .Z(n25) );
  NANDN U29 ( .A(A[2]), .B(n11), .Z(n26) );
  NANDN U30 ( .A(n11), .B(A[2]), .Z(n24) );
  AND U31 ( .A(n27), .B(n28), .Z(n11) );
  NAND U32 ( .A(B[1]), .B(n29), .Z(n28) );
  OR U33 ( .A(n13), .B(A[1]), .Z(n29) );
  NAND U34 ( .A(A[1]), .B(n13), .Z(n27) );
  AND U35 ( .A(B[0]), .B(A[0]), .Z(n13) );
  XOR U36 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_84 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_85 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_86 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_87 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_88 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_89 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_90 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_91 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_92 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_93 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_94 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_95 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_96 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_97 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_98 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_99 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_100 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_101 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_102 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_103 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_104 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_105 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_106 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_107 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_108 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_109 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_110 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_111 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_112 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_113 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_114 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_115 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_116 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_117 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_118 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_119 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_120 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_121 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_122 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_123 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_124 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_125 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_126 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_127 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_128 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_129 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_130 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_131 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_132 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_133 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_134 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_135 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_136 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_137 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_138 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_139 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_140 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_141 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_142 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_143 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_144 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_145 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_146 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_147 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_148 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_149 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_150 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_151 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_152 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_153 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_154 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_155 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_156 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_157 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_158 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_159 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_160 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_161 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_162 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_163 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_164 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_165 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_166 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n12), .B(n13), .Z(SUM[6]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[5]) );
  XNOR U3 ( .A(B[5]), .B(A[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[4]) );
  XNOR U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[3]) );
  XNOR U7 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[2]) );
  XNOR U9 ( .A(B[2]), .B(A[2]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[1]) );
  XOR U11 ( .A(B[1]), .B(A[1]), .Z(n11) );
  NAND U12 ( .A(B[5]), .B(n14), .Z(n13) );
  NANDN U13 ( .A(A[5]), .B(n2), .Z(n14) );
  NANDN U14 ( .A(n2), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n15), .B(n16), .Z(n2) );
  NAND U16 ( .A(B[4]), .B(n17), .Z(n16) );
  NANDN U17 ( .A(A[4]), .B(n4), .Z(n17) );
  NANDN U18 ( .A(n4), .B(A[4]), .Z(n15) );
  AND U19 ( .A(n18), .B(n19), .Z(n4) );
  NAND U20 ( .A(B[3]), .B(n20), .Z(n19) );
  NANDN U21 ( .A(A[3]), .B(n6), .Z(n20) );
  NANDN U22 ( .A(n6), .B(A[3]), .Z(n18) );
  AND U23 ( .A(n21), .B(n22), .Z(n6) );
  NAND U24 ( .A(B[2]), .B(n23), .Z(n22) );
  NANDN U25 ( .A(A[2]), .B(n8), .Z(n23) );
  NANDN U26 ( .A(n8), .B(A[2]), .Z(n21) );
  AND U27 ( .A(n24), .B(n25), .Z(n8) );
  NAND U28 ( .A(B[1]), .B(n26), .Z(n25) );
  OR U29 ( .A(n10), .B(A[1]), .Z(n26) );
  NAND U30 ( .A(A[1]), .B(n10), .Z(n24) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n10) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_167 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_168 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_169 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_170 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_171 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_172 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_173 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_174 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_175 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_176 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_177 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_178 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_179 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_180 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_181 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_182 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_183 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_184 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_185 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_186 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_187 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_188 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_189 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_190 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_191 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_192 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_193 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_194 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_195 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_196 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_197 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_198 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_199 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_200 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_201 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_202 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_203 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_204 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_205 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_206 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_207 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_208 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_209 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_210 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_211 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_212 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_213 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_214 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_215 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_216 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_217 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_218 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_219 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_220 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_221 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_222 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_223 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_224 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_225 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_226 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_227 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_228 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_229 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_230 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_231 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_232 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_233 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_234 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_235 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_236 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_237 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_238 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_239 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_240 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_241 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_242 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_243 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_244 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_245 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_246 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_247 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_248 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_249 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_250 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_251 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_252 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_253 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_254 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_255 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_256 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_257 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_258 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_259 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_260 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_261 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_262 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_263 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_264 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_265 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_266 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_267 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_268 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_269 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_270 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_271 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_272 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_273 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_274 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_275 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_276 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_277 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_278 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_279 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_280 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_281 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_282 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_283 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_284 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_285 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_286 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_287 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_288 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_289 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_290 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_291 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_292 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_293 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_294 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_295 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_296 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_297 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_298 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_299 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_300 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_301 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_302 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_303 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_304 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_305 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_306 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_307 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_308 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_309 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_310 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_311 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_312 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_313 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_314 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_315 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_316 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_317 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_318 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_319 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_320 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_321 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_322 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_323 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_324 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_325 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_326 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_327 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_328 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_329 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_330 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_331 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_332 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XOR U2 ( .A(n2), .B(n3), .Z(SUM[4]) );
  XNOR U3 ( .A(B[4]), .B(A[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n5), .Z(SUM[3]) );
  XNOR U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[2]) );
  XNOR U7 ( .A(B[2]), .B(A[2]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[1]) );
  XOR U9 ( .A(B[1]), .B(A[1]), .Z(n9) );
  NAND U10 ( .A(B[4]), .B(n12), .Z(n11) );
  NANDN U11 ( .A(A[4]), .B(n2), .Z(n12) );
  NANDN U12 ( .A(n2), .B(A[4]), .Z(n10) );
  AND U13 ( .A(n13), .B(n14), .Z(n2) );
  NAND U14 ( .A(B[3]), .B(n15), .Z(n14) );
  NANDN U15 ( .A(A[3]), .B(n4), .Z(n15) );
  NANDN U16 ( .A(n4), .B(A[3]), .Z(n13) );
  AND U17 ( .A(n16), .B(n17), .Z(n4) );
  NAND U18 ( .A(B[2]), .B(n18), .Z(n17) );
  NANDN U19 ( .A(A[2]), .B(n6), .Z(n18) );
  NANDN U20 ( .A(n6), .B(A[2]), .Z(n16) );
  AND U21 ( .A(n19), .B(n20), .Z(n6) );
  NAND U22 ( .A(B[1]), .B(n21), .Z(n20) );
  OR U23 ( .A(n8), .B(A[1]), .Z(n21) );
  NAND U24 ( .A(A[1]), .B(n8), .Z(n19) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n8) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2_DW01_add_333 ( A, B, CI, SUM, CO );
  input [12:0] A;
  input [12:0] B;
  output [12:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19;

  AND U1 ( .A(B[4]), .B(n2), .Z(SUM[5]) );
  IV U2 ( .A(n4), .Z(n2) );
  IV U3 ( .A(B[4]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n3), .Z(SUM[4]) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[3]) );
  XNOR U6 ( .A(B[3]), .B(A[3]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[2]) );
  XNOR U8 ( .A(B[2]), .B(A[2]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[1]) );
  XOR U10 ( .A(B[1]), .B(A[1]), .Z(n10) );
  AND U11 ( .A(n11), .B(n12), .Z(n4) );
  NAND U12 ( .A(B[3]), .B(n13), .Z(n12) );
  NANDN U13 ( .A(A[3]), .B(n5), .Z(n13) );
  NANDN U14 ( .A(n5), .B(A[3]), .Z(n11) );
  AND U15 ( .A(n14), .B(n15), .Z(n5) );
  NAND U16 ( .A(B[2]), .B(n16), .Z(n15) );
  NANDN U17 ( .A(A[2]), .B(n7), .Z(n16) );
  NANDN U18 ( .A(n7), .B(A[2]), .Z(n14) );
  AND U19 ( .A(n17), .B(n18), .Z(n7) );
  NAND U20 ( .A(B[1]), .B(n19), .Z(n18) );
  OR U21 ( .A(n9), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(A[1]), .B(n9), .Z(n17) );
  AND U23 ( .A(B[0]), .B(A[0]), .Z(n9) );
  XOR U24 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC2 ( clk, rst, x, y, o );
  input [7999:0] x;
  input [7999:0] y;
  output [13:0] o;
  input clk, rst;
  wire   N60579, N60580, N60581, N60582, N60592, N60593, N60594, N60595,
         N60596, N60605, N60606, N60607, N60608, N60609, N60618, N60619,
         N60620, N60621, N60622, N60631, N60632, N60633, N60634, N60635,
         N60644, N60645, N60646, N60647, N60648, N60657, N60658, N60659,
         N60660, N60661, N60670, N60671, N60672, N60673, N60674, N60683,
         N60684, N60685, N60686, N60687, N60696, N60697, N60698, N60699,
         N60700, N60709, N60710, N60711, N60712, N60713, N60722, N60723,
         N60724, N60725, N60726, N60735, N60736, N60737, N60738, N60739,
         N60748, N60749, N60750, N60751, N60752, N60761, N60762, N60763,
         N60764, N60765, N60774, N60775, N60776, N60777, N60778, N60787,
         N60788, N60789, N60790, N60791, N60800, N60801, N60802, N60803,
         N60804, N60813, N60814, N60815, N60816, N60817, N60826, N60827,
         N60828, N60829, N60830, N60839, N60840, N60841, N60842, N60843,
         N60852, N60853, N60854, N60855, N60856, N60865, N60866, N60867,
         N60868, N60869, N60878, N60879, N60880, N60881, N60882, N60891,
         N60892, N60893, N60894, N60895, N60904, N60905, N60906, N60907,
         N60908, N60917, N60918, N60919, N60920, N60921, N60930, N60931,
         N60932, N60933, N60934, N60943, N60944, N60945, N60946, N60947,
         N60956, N60957, N60958, N60959, N60960, N60969, N60970, N60971,
         N60972, N60973, N60982, N60983, N60984, N60985, N60986, N60995,
         N60996, N60997, N60998, N60999, N61008, N61009, N61010, N61011,
         N61012, N61021, N61022, N61023, N61024, N61025, N61034, N61035,
         N61036, N61037, N61038, N61047, N61048, N61049, N61050, N61051,
         N61060, N61061, N61062, N61063, N61064, N61073, N61074, N61075,
         N61076, N61077, N61086, N61087, N61088, N61089, N61090, N61099,
         N61100, N61101, N61102, N61103, N61112, N61113, N61114, N61115,
         N61116, N61125, N61126, N61127, N61128, N61129, N61138, N61139,
         N61140, N61141, N61142, N61151, N61152, N61153, N61154, N61155,
         N61164, N61165, N61166, N61167, N61168, N61177, N61178, N61179,
         N61180, N61181, N61190, N61191, N61192, N61193, N61194, N61203,
         N61204, N61205, N61206, N61207, N61216, N61217, N61218, N61219,
         N61220, N61229, N61230, N61231, N61232, N61233, N61242, N61243,
         N61244, N61245, N61246, N61255, N61256, N61257, N61258, N61259,
         N61268, N61269, N61270, N61271, N61272, N61281, N61282, N61283,
         N61284, N61285, N61294, N61295, N61296, N61297, N61298, N61307,
         N61308, N61309, N61310, N61311, N61320, N61321, N61322, N61323,
         N61324, N61333, N61334, N61335, N61336, N61337, N61346, N61347,
         N61348, N61349, N61350, N61359, N61360, N61361, N61362, N61363,
         N61372, N61373, N61374, N61375, N61376, N61385, N61386, N61387,
         N61388, N61389, N61398, N61399, N61400, N61401, N61402, N61411,
         N61412, N61413, N61414, N61415, N61424, N61425, N61426, N61427,
         N61428, N61437, N61438, N61439, N61440, N61441, N61450, N61451,
         N61452, N61453, N61454, N61463, N61464, N61465, N61466, N61467,
         N61476, N61477, N61478, N61479, N61480, N61489, N61490, N61491,
         N61492, N61493, N61502, N61503, N61504, N61505, N61506, N61515,
         N61516, N61517, N61518, N61519, N61528, N61529, N61530, N61531,
         N61532, N61541, N61542, N61543, N61544, N61545, N61554, N61555,
         N61556, N61557, N61558, N61567, N61568, N61569, N61570, N61571,
         N61580, N61581, N61582, N61583, N61584, N61593, N61594, N61595,
         N61596, N61597, N61606, N61607, N61608, N61609, N61610, N61619,
         N61620, N61621, N61622, N61623, N61632, N61633, N61634, N61635,
         N61636, N61645, N61646, N61647, N61648, N61649, N61658, N61659,
         N61660, N61661, N61662, N61671, N61672, N61673, N61674, N61675,
         N61684, N61685, N61686, N61687, N61688, N61697, N61698, N61699,
         N61700, N61701, N61710, N61711, N61712, N61713, N61714, N61723,
         N61724, N61725, N61726, N61727, N61736, N61737, N61738, N61739,
         N61740, N61749, N61750, N61751, N61752, N61753, N61762, N61763,
         N61764, N61765, N61766, N61775, N61776, N61777, N61778, N61779,
         N61788, N61789, N61790, N61791, N61792, N61801, N61802, N61803,
         N61804, N61805, N61814, N61815, N61816, N61817, N61818, N61827,
         N61828, N61829, N61830, N61831, N61840, N61841, N61842, N61843,
         N61844, N61853, N61854, N61855, N61856, N61857, N61866, N61867,
         N61868, N61869, N61870, N61879, N61880, N61881, N61882, N61883,
         N61892, N61893, N61894, N61895, N61896, N61905, N61906, N61907,
         N61908, N61909, N61918, N61919, N61920, N61921, N61922, N61931,
         N61932, N61933, N61934, N61935, N61944, N61945, N61946, N61947,
         N61948, N61957, N61958, N61959, N61960, N61961, N61970, N61971,
         N61972, N61973, N61974, N61983, N61984, N61985, N61986, N61987,
         N61996, N61997, N61998, N61999, N62000, N62009, N62010, N62011,
         N62012, N62013, N62022, N62023, N62024, N62025, N62026, N62035,
         N62036, N62037, N62038, N62039, N62048, N62049, N62050, N62051,
         N62052, N62061, N62062, N62063, N62064, N62065, N62074, N62075,
         N62076, N62077, N62078, N62087, N62088, N62089, N62090, N62091,
         N62100, N62101, N62102, N62103, N62104, N62113, N62114, N62115,
         N62116, N62117, N62126, N62127, N62128, N62129, N62130, N62139,
         N62140, N62141, N62142, N62143, N62152, N62153, N62154, N62155,
         N62156, N62165, N62166, N62167, N62168, N62169, N62178, N62179,
         N62180, N62181, N62182, N62191, N62192, N62193, N62194, N62195,
         N62204, N62205, N62206, N62207, N62208, N62217, N62218, N62219,
         N62220, N62221, N62230, N62231, N62232, N62233, N62234, N62243,
         N62244, N62245, N62246, N62247, N62256, N62257, N62258, N62259,
         N62260, N62269, N62270, N62271, N62272, N62273, N62282, N62283,
         N62284, N62285, N62286, N62295, N62296, N62297, N62298, N62299,
         N62308, N62309, N62310, N62311, N62312, N62321, N62322, N62323,
         N62324, N62325, N62334, N62335, N62336, N62337, N62338, N62347,
         N62348, N62349, N62350, N62351, N62360, N62361, N62362, N62363,
         N62364, N62373, N62374, N62375, N62376, N62377, N62386, N62387,
         N62388, N62389, N62390, N62399, N62400, N62401, N62402, N62403,
         N62412, N62413, N62414, N62415, N62416, N62425, N62426, N62427,
         N62428, N62429, N62438, N62439, N62440, N62441, N62442, N62451,
         N62452, N62453, N62454, N62455, N62464, N62465, N62466, N62467,
         N62468, N62477, N62478, N62479, N62480, N62481, N62490, N62491,
         N62492, N62493, N62494, N62503, N62504, N62505, N62506, N62507,
         N62516, N62517, N62518, N62519, N62520, N62529, N62530, N62531,
         N62532, N62533, N62542, N62543, N62544, N62545, N62546, N62555,
         N62556, N62557, N62558, N62559, N62568, N62569, N62570, N62571,
         N62572, N62581, N62582, N62583, N62584, N62585, N62594, N62595,
         N62596, N62597, N62598, N62607, N62608, N62609, N62610, N62611,
         N62620, N62621, N62622, N62623, N62624, N62633, N62634, N62635,
         N62636, N62637, N62646, N62647, N62648, N62649, N62650, N62659,
         N62660, N62661, N62662, N62663, N62672, N62673, N62674, N62675,
         N62676, N62685, N62686, N62687, N62688, N62689, N62698, N62699,
         N62700, N62701, N62702, N62711, N62712, N62713, N62714, N62715,
         N62724, N62725, N62726, N62727, N62728, N62737, N62738, N62739,
         N62740, N62741, N62750, N62751, N62752, N62753, N62754, N62763,
         N62764, N62765, N62766, N62767, N62776, N62777, N62778, N62779,
         N62780, N62789, N62790, N62791, N62792, N62793, N62802, N62803,
         N62804, N62805, N62806, N62815, N62816, N62817, N62818, N62819,
         N62828, N62829, N62830, N62831, N62832, N62841, N62842, N62843,
         N62844, N62845, N62854, N62855, N62856, N62857, N62858, N62867,
         N62868, N62869, N62870, N62871, N62880, N62881, N62882, N62883,
         N62884, N62893, N62894, N62895, N62896, N62897, N62906, N62907,
         N62908, N62909, N62910, N62919, N62920, N62921, N62922, N62923,
         N62932, N62933, N62934, N62935, N62936, N62945, N62946, N62947,
         N62948, N62949, N62958, N62959, N62960, N62961, N62962, N62971,
         N62972, N62973, N62974, N62975, N62984, N62985, N62986, N62987,
         N62988, N62997, N62998, N62999, N63000, N63001, N63010, N63011,
         N63012, N63013, N63014, N63023, N63024, N63025, N63026, N63027,
         N63036, N63037, N63038, N63039, N63040, N63049, N63050, N63051,
         N63052, N63053, N63062, N63063, N63064, N63065, N63066, N63075,
         N63076, N63077, N63078, N63079, N63088, N63089, N63090, N63091,
         N63092, N63101, N63102, N63103, N63104, N63105, N63114, N63115,
         N63116, N63117, N63118, N63127, N63128, N63129, N63130, N63131,
         N63140, N63141, N63142, N63143, N63144, N63153, N63154, N63155,
         N63156, N63157, N63166, N63167, N63168, N63169, N63170, N63179,
         N63180, N63181, N63182, N63183, N63192, N63193, N63194, N63195,
         N63196, N63205, N63206, N63207, N63208, N63209, N63218, N63219,
         N63220, N63221, N63222, N63231, N63232, N63233, N63234, N63235,
         N63244, N63245, N63246, N63247, N63248, N63257, N63258, N63259,
         N63260, N63261, N63270, N63271, N63272, N63273, N63274, N63283,
         N63284, N63285, N63286, N63287, N63296, N63297, N63298, N63299,
         N63300, N63309, N63310, N63311, N63312, N63313, N63322, N63323,
         N63324, N63325, N63326, N63335, N63336, N63337, N63338, N63339,
         N63348, N63349, N63350, N63351, N63352, N63361, N63362, N63363,
         N63364, N63365, N63374, N63375, N63376, N63377, N63378, N63387,
         N63388, N63389, N63390, N63391, N63400, N63401, N63402, N63403,
         N63404, N63413, N63414, N63415, N63416, N63417, N63426, N63427,
         N63428, N63429, N63430, N63439, N63440, N63441, N63442, N63443,
         N63452, N63453, N63454, N63455, N63456, N63465, N63466, N63467,
         N63468, N63469, N63478, N63479, N63480, N63481, N63482, N63491,
         N63492, N63493, N63494, N63495, N63504, N63505, N63506, N63507,
         N63508, N63517, N63518, N63519, N63520, N63521, N63530, N63531,
         N63532, N63533, N63534, N63543, N63544, N63545, N63546, N63547,
         N63556, N63557, N63558, N63559, N63560, N63569, N63570, N63571,
         N63572, N63573, N63582, N63583, N63584, N63585, N63586, N63595,
         N63596, N63597, N63598, N63599, N63608, N63609, N63610, N63611,
         N63612, N63621, N63622, N63623, N63624, N63625, N63634, N63635,
         N63636, N63637, N63638, N63647, N63648, N63649, N63650, N63651,
         N63660, N63661, N63662, N63663, N63664, N63673, N63674, N63675,
         N63676, N63677, N63686, N63687, N63688, N63689, N63690, N63699,
         N63700, N63701, N63702, N63703, N63712, N63713, N63714, N63715,
         N63716, N63725, N63726, N63727, N63728, N63729, N63738, N63739,
         N63740, N63741, N63742, N63751, N63752, N63753, N63754, N63755,
         N63764, N63765, N63766, N63767, N63768, N63777, N63778, N63779,
         N63780, N63781, N63790, N63791, N63792, N63793, N63794, N63803,
         N63804, N63805, N63806, N63807, N63816, N63817, N63818, N63819,
         N63820, N63829, N63830, N63831, N63832, N63833, N63842, N63843,
         N63844, N63845, N63846, N63855, N63856, N63857, N63858, N63859,
         N63868, N63869, N63870, N63871, N63872, N63881, N63882, N63883,
         N63884, N63885, N63894, N63895, N63896, N63897, N63898, N63907,
         N63908, N63909, N63910, N63911, N63920, N63921, N63922, N63923,
         N63924, N63933, N63934, N63935, N63936, N63937, N63946, N63947,
         N63948, N63949, N63950, N63959, N63960, N63961, N63962, N63963,
         N63972, N63973, N63974, N63975, N63976, N63985, N63986, N63987,
         N63988, N63989, N63998, N63999, N64000, N64001, N64002, N64011,
         N64012, N64013, N64014, N64015, N64024, N64025, N64026, N64027,
         N64028, N64037, N64038, N64039, N64040, N64041, N64050, N64051,
         N64052, N64053, N64054, N64063, N64064, N64065, N64066, N64067,
         N64076, N64077, N64078, N64079, N64080, N64089, N64090, N64091,
         N64092, N64093, N64102, N64103, N64104, N64105, N64106, N64115,
         N64116, N64117, N64118, N64119, N64128, N64129, N64130, N64131,
         N64132, N64141, N64142, N64143, N64144, N64145, N64154, N64155,
         N64156, N64157, N64158, N64167, N64168, N64169, N64170, N64171,
         N64180, N64181, N64182, N64183, N64184, N64193, N64194, N64195,
         N64196, N64197, N64206, N64207, N64208, N64209, N64210, N64219,
         N64220, N64221, N64222, N64223, N64232, N64233, N64234, N64235,
         N64236, N64245, N64246, N64247, N64248, N64249, N64258, N64259,
         N64260, N64261, N64262, N64271, N64272, N64273, N64274, N64275,
         N64284, N64285, N64286, N64287, N64288, N64297, N64298, N64299,
         N64300, N64301, N64310, N64311, N64312, N64313, N64314, N64323,
         N64324, N64325, N64326, N64327, N64336, N64337, N64338, N64339,
         N64340, N64349, N64350, N64351, N64352, N64353, N64362, N64363,
         N64364, N64365, N64366, N64375, N64376, N64377, N64378, N64379,
         N64388, N64389, N64390, N64391, N64392, N64401, N64402, N64403,
         N64404, N64405, N64414, N64415, N64416, N64417, N64418, N64427,
         N64428, N64429, N64430, N64431, N64440, N64441, N64442, N64443,
         N64444, N64453, N64454, N64455, N64456, N64457, N64466, N64467,
         N64468, N64469, N64470, N64479, N64480, N64481, N64482, N64483,
         N64492, N64493, N64494, N64495, N64496, N64505, N64506, N64507,
         N64508, N64509, N64518, N64519, N64520, N64521, N64522, N64531,
         N64532, N64533, N64534, N64535, N64544, N64545, N64546, N64547,
         N64548, N64557, N64558, N64559, N64560, N64561, N64570, N64571,
         N64572, N64573, N64574, N64583, N64584, N64585, N64586, N64587,
         N64596, N64597, N64598, N64599, N64600, N64609, N64610, N64611,
         N64612, N64613, N64622, N64623, N64624, N64625, N64626, N64635,
         N64636, N64637, N64638, N64639, N64648, N64649, N64650, N64651,
         N64652, N64661, N64662, N64663, N64664, N64665, N64674, N64675,
         N64676, N64677, N64678, N64687, N64688, N64689, N64690, N64691,
         N64700, N64701, N64702, N64703, N64704, N64713, N64714, N64715,
         N64716, N64717, N64726, N64727, N64728, N64729, N64730, N64739,
         N64740, N64741, N64742, N64743, N64752, N64753, N64754, N64755,
         N64756, N64765, N64766, N64767, N64768, N64769, N64778, N64779,
         N64780, N64781, N64782, N64791, N64792, N64793, N64794, N64795,
         N64804, N64805, N64806, N64807, N64808, N64817, N64818, N64819,
         N64820, N64821, N64830, N64831, N64832, N64833, N64834, N64843,
         N64844, N64845, N64846, N64847, N64856, N64857, N64858, N64859,
         N64860, N64869, N64870, N64871, N64872, N64873, N64882, N64883,
         N64884, N64885, N64886, N64895, N64896, N64897, N64898, N64899,
         N64908, N64909, N64910, N64911, N64912, N64921, N64922, N64923,
         N64924, N64925, N64926, N64934, N64935, N64936, N64937, N64938,
         N64939, N64947, N64948, N64949, N64950, N64951, N64952, N64960,
         N64961, N64962, N64963, N64964, N64965, N64973, N64974, N64975,
         N64976, N64977, N64978, N64986, N64987, N64988, N64989, N64990,
         N64991, N64999, N65000, N65001, N65002, N65003, N65004, N65012,
         N65013, N65014, N65015, N65016, N65017, N65025, N65026, N65027,
         N65028, N65029, N65030, N65038, N65039, N65040, N65041, N65042,
         N65043, N65051, N65052, N65053, N65054, N65055, N65056, N65064,
         N65065, N65066, N65067, N65068, N65069, N65077, N65078, N65079,
         N65080, N65081, N65082, N65090, N65091, N65092, N65093, N65094,
         N65095, N65103, N65104, N65105, N65106, N65107, N65108, N65116,
         N65117, N65118, N65119, N65120, N65121, N65129, N65130, N65131,
         N65132, N65133, N65134, N65142, N65143, N65144, N65145, N65146,
         N65147, N65155, N65156, N65157, N65158, N65159, N65160, N65168,
         N65169, N65170, N65171, N65172, N65173, N65181, N65182, N65183,
         N65184, N65185, N65186, N65194, N65195, N65196, N65197, N65198,
         N65199, N65207, N65208, N65209, N65210, N65211, N65212, N65220,
         N65221, N65222, N65223, N65224, N65225, N65233, N65234, N65235,
         N65236, N65237, N65238, N65246, N65247, N65248, N65249, N65250,
         N65251, N65259, N65260, N65261, N65262, N65263, N65264, N65272,
         N65273, N65274, N65275, N65276, N65277, N65285, N65286, N65287,
         N65288, N65289, N65290, N65298, N65299, N65300, N65301, N65302,
         N65303, N65311, N65312, N65313, N65314, N65315, N65316, N65324,
         N65325, N65326, N65327, N65328, N65329, N65337, N65338, N65339,
         N65340, N65341, N65342, N65350, N65351, N65352, N65353, N65354,
         N65355, N65363, N65364, N65365, N65366, N65367, N65368, N65376,
         N65377, N65378, N65379, N65380, N65381, N65389, N65390, N65391,
         N65392, N65393, N65394, N65402, N65403, N65404, N65405, N65406,
         N65407, N65415, N65416, N65417, N65418, N65419, N65420, N65428,
         N65429, N65430, N65431, N65432, N65433, N65441, N65442, N65443,
         N65444, N65445, N65446, N65454, N65455, N65456, N65457, N65458,
         N65459, N65467, N65468, N65469, N65470, N65471, N65472, N65480,
         N65481, N65482, N65483, N65484, N65485, N65493, N65494, N65495,
         N65496, N65497, N65498, N65506, N65507, N65508, N65509, N65510,
         N65511, N65519, N65520, N65521, N65522, N65523, N65524, N65532,
         N65533, N65534, N65535, N65536, N65537, N65545, N65546, N65547,
         N65548, N65549, N65550, N65558, N65559, N65560, N65561, N65562,
         N65563, N65571, N65572, N65573, N65574, N65575, N65576, N65584,
         N65585, N65586, N65587, N65588, N65589, N65597, N65598, N65599,
         N65600, N65601, N65602, N65610, N65611, N65612, N65613, N65614,
         N65615, N65623, N65624, N65625, N65626, N65627, N65628, N65636,
         N65637, N65638, N65639, N65640, N65641, N65649, N65650, N65651,
         N65652, N65653, N65654, N65662, N65663, N65664, N65665, N65666,
         N65667, N65675, N65676, N65677, N65678, N65679, N65680, N65688,
         N65689, N65690, N65691, N65692, N65693, N65701, N65702, N65703,
         N65704, N65705, N65706, N65714, N65715, N65716, N65717, N65718,
         N65719, N65727, N65728, N65729, N65730, N65731, N65732, N65740,
         N65741, N65742, N65743, N65744, N65745, N65753, N65754, N65755,
         N65756, N65757, N65758, N65766, N65767, N65768, N65769, N65770,
         N65771, N65779, N65780, N65781, N65782, N65783, N65784, N65792,
         N65793, N65794, N65795, N65796, N65797, N65805, N65806, N65807,
         N65808, N65809, N65810, N65818, N65819, N65820, N65821, N65822,
         N65823, N65831, N65832, N65833, N65834, N65835, N65836, N65844,
         N65845, N65846, N65847, N65848, N65849, N65857, N65858, N65859,
         N65860, N65861, N65862, N65870, N65871, N65872, N65873, N65874,
         N65875, N65883, N65884, N65885, N65886, N65887, N65888, N65896,
         N65897, N65898, N65899, N65900, N65901, N65909, N65910, N65911,
         N65912, N65913, N65914, N65922, N65923, N65924, N65925, N65926,
         N65927, N65935, N65936, N65937, N65938, N65939, N65940, N65948,
         N65949, N65950, N65951, N65952, N65953, N65961, N65962, N65963,
         N65964, N65965, N65966, N65974, N65975, N65976, N65977, N65978,
         N65979, N65987, N65988, N65989, N65990, N65991, N65992, N66000,
         N66001, N66002, N66003, N66004, N66005, N66013, N66014, N66015,
         N66016, N66017, N66018, N66026, N66027, N66028, N66029, N66030,
         N66031, N66039, N66040, N66041, N66042, N66043, N66044, N66052,
         N66053, N66054, N66055, N66056, N66057, N66065, N66066, N66067,
         N66068, N66069, N66070, N66078, N66079, N66080, N66081, N66082,
         N66083, N66091, N66092, N66093, N66094, N66095, N66096, N66104,
         N66105, N66106, N66107, N66108, N66109, N66117, N66118, N66119,
         N66120, N66121, N66122, N66130, N66131, N66132, N66133, N66134,
         N66135, N66143, N66144, N66145, N66146, N66147, N66148, N66156,
         N66157, N66158, N66159, N66160, N66161, N66169, N66170, N66171,
         N66172, N66173, N66174, N66182, N66183, N66184, N66185, N66186,
         N66187, N66195, N66196, N66197, N66198, N66199, N66200, N66208,
         N66209, N66210, N66211, N66212, N66213, N66221, N66222, N66223,
         N66224, N66225, N66226, N66234, N66235, N66236, N66237, N66238,
         N66239, N66247, N66248, N66249, N66250, N66251, N66252, N66260,
         N66261, N66262, N66263, N66264, N66265, N66273, N66274, N66275,
         N66276, N66277, N66278, N66286, N66287, N66288, N66289, N66290,
         N66291, N66299, N66300, N66301, N66302, N66303, N66304, N66312,
         N66313, N66314, N66315, N66316, N66317, N66325, N66326, N66327,
         N66328, N66329, N66330, N66338, N66339, N66340, N66341, N66342,
         N66343, N66351, N66352, N66353, N66354, N66355, N66356, N66364,
         N66365, N66366, N66367, N66368, N66369, N66377, N66378, N66379,
         N66380, N66381, N66382, N66390, N66391, N66392, N66393, N66394,
         N66395, N66403, N66404, N66405, N66406, N66407, N66408, N66416,
         N66417, N66418, N66419, N66420, N66421, N66429, N66430, N66431,
         N66432, N66433, N66434, N66442, N66443, N66444, N66445, N66446,
         N66447, N66455, N66456, N66457, N66458, N66459, N66460, N66468,
         N66469, N66470, N66471, N66472, N66473, N66481, N66482, N66483,
         N66484, N66485, N66486, N66494, N66495, N66496, N66497, N66498,
         N66499, N66507, N66508, N66509, N66510, N66511, N66512, N66520,
         N66521, N66522, N66523, N66524, N66525, N66533, N66534, N66535,
         N66536, N66537, N66538, N66546, N66547, N66548, N66549, N66550,
         N66551, N66559, N66560, N66561, N66562, N66563, N66564, N66572,
         N66573, N66574, N66575, N66576, N66577, N66585, N66586, N66587,
         N66588, N66589, N66590, N66598, N66599, N66600, N66601, N66602,
         N66603, N66611, N66612, N66613, N66614, N66615, N66616, N66624,
         N66625, N66626, N66627, N66628, N66629, N66637, N66638, N66639,
         N66640, N66641, N66642, N66650, N66651, N66652, N66653, N66654,
         N66655, N66663, N66664, N66665, N66666, N66667, N66668, N66676,
         N66677, N66678, N66679, N66680, N66681, N66689, N66690, N66691,
         N66692, N66693, N66694, N66702, N66703, N66704, N66705, N66706,
         N66707, N66715, N66716, N66717, N66718, N66719, N66720, N66728,
         N66729, N66730, N66731, N66732, N66733, N66741, N66742, N66743,
         N66744, N66745, N66746, N66754, N66755, N66756, N66757, N66758,
         N66759, N66767, N66768, N66769, N66770, N66771, N66772, N66780,
         N66781, N66782, N66783, N66784, N66785, N66793, N66794, N66795,
         N66796, N66797, N66798, N66806, N66807, N66808, N66809, N66810,
         N66811, N66819, N66820, N66821, N66822, N66823, N66824, N66832,
         N66833, N66834, N66835, N66836, N66837, N66845, N66846, N66847,
         N66848, N66849, N66850, N66858, N66859, N66860, N66861, N66862,
         N66863, N66871, N66872, N66873, N66874, N66875, N66876, N66884,
         N66885, N66886, N66887, N66888, N66889, N66897, N66898, N66899,
         N66900, N66901, N66902, N66910, N66911, N66912, N66913, N66914,
         N66915, N66923, N66924, N66925, N66926, N66927, N66928, N66936,
         N66937, N66938, N66939, N66940, N66941, N66949, N66950, N66951,
         N66952, N66953, N66954, N66962, N66963, N66964, N66965, N66966,
         N66967, N66975, N66976, N66977, N66978, N66979, N66980, N66988,
         N66989, N66990, N66991, N66992, N66993, N67001, N67002, N67003,
         N67004, N67005, N67006, N67014, N67015, N67016, N67017, N67018,
         N67019, N67027, N67028, N67029, N67030, N67031, N67032, N67040,
         N67041, N67042, N67043, N67044, N67045, N67053, N67054, N67055,
         N67056, N67057, N67058, N67066, N67067, N67068, N67069, N67070,
         N67071, N67079, N67080, N67081, N67082, N67083, N67084, N67092,
         N67093, N67094, N67095, N67096, N67097, N67098, N67105, N67106,
         N67107, N67108, N67109, N67110, N67111, N67118, N67119, N67120,
         N67121, N67122, N67123, N67124, N67131, N67132, N67133, N67134,
         N67135, N67136, N67137, N67144, N67145, N67146, N67147, N67148,
         N67149, N67150, N67157, N67158, N67159, N67160, N67161, N67162,
         N67163, N67170, N67171, N67172, N67173, N67174, N67175, N67176,
         N67183, N67184, N67185, N67186, N67187, N67188, N67189, N67196,
         N67197, N67198, N67199, N67200, N67201, N67202, N67209, N67210,
         N67211, N67212, N67213, N67214, N67215, N67222, N67223, N67224,
         N67225, N67226, N67227, N67228, N67235, N67236, N67237, N67238,
         N67239, N67240, N67241, N67248, N67249, N67250, N67251, N67252,
         N67253, N67254, N67261, N67262, N67263, N67264, N67265, N67266,
         N67267, N67274, N67275, N67276, N67277, N67278, N67279, N67280,
         N67287, N67288, N67289, N67290, N67291, N67292, N67293, N67300,
         N67301, N67302, N67303, N67304, N67305, N67306, N67313, N67314,
         N67315, N67316, N67317, N67318, N67319, N67326, N67327, N67328,
         N67329, N67330, N67331, N67332, N67339, N67340, N67341, N67342,
         N67343, N67344, N67345, N67352, N67353, N67354, N67355, N67356,
         N67357, N67358, N67365, N67366, N67367, N67368, N67369, N67370,
         N67371, N67378, N67379, N67380, N67381, N67382, N67383, N67384,
         N67391, N67392, N67393, N67394, N67395, N67396, N67397, N67404,
         N67405, N67406, N67407, N67408, N67409, N67410, N67417, N67418,
         N67419, N67420, N67421, N67422, N67423, N67430, N67431, N67432,
         N67433, N67434, N67435, N67436, N67443, N67444, N67445, N67446,
         N67447, N67448, N67449, N67456, N67457, N67458, N67459, N67460,
         N67461, N67462, N67469, N67470, N67471, N67472, N67473, N67474,
         N67475, N67482, N67483, N67484, N67485, N67486, N67487, N67488,
         N67495, N67496, N67497, N67498, N67499, N67500, N67501, N67508,
         N67509, N67510, N67511, N67512, N67513, N67514, N67521, N67522,
         N67523, N67524, N67525, N67526, N67527, N67534, N67535, N67536,
         N67537, N67538, N67539, N67540, N67547, N67548, N67549, N67550,
         N67551, N67552, N67553, N67560, N67561, N67562, N67563, N67564,
         N67565, N67566, N67573, N67574, N67575, N67576, N67577, N67578,
         N67579, N67586, N67587, N67588, N67589, N67590, N67591, N67592,
         N67599, N67600, N67601, N67602, N67603, N67604, N67605, N67612,
         N67613, N67614, N67615, N67616, N67617, N67618, N67625, N67626,
         N67627, N67628, N67629, N67630, N67631, N67638, N67639, N67640,
         N67641, N67642, N67643, N67644, N67651, N67652, N67653, N67654,
         N67655, N67656, N67657, N67664, N67665, N67666, N67667, N67668,
         N67669, N67670, N67677, N67678, N67679, N67680, N67681, N67682,
         N67683, N67690, N67691, N67692, N67693, N67694, N67695, N67696,
         N67703, N67704, N67705, N67706, N67707, N67708, N67709, N67716,
         N67717, N67718, N67719, N67720, N67721, N67722, N67729, N67730,
         N67731, N67732, N67733, N67734, N67735, N67742, N67743, N67744,
         N67745, N67746, N67747, N67748, N67755, N67756, N67757, N67758,
         N67759, N67760, N67761, N67768, N67769, N67770, N67771, N67772,
         N67773, N67774, N67781, N67782, N67783, N67784, N67785, N67786,
         N67787, N67794, N67795, N67796, N67797, N67798, N67799, N67800,
         N67807, N67808, N67809, N67810, N67811, N67812, N67813, N67820,
         N67821, N67822, N67823, N67824, N67825, N67826, N67833, N67834,
         N67835, N67836, N67837, N67838, N67839, N67846, N67847, N67848,
         N67849, N67850, N67851, N67852, N67859, N67860, N67861, N67862,
         N67863, N67864, N67865, N67872, N67873, N67874, N67875, N67876,
         N67877, N67878, N67885, N67886, N67887, N67888, N67889, N67890,
         N67891, N67898, N67899, N67900, N67901, N67902, N67903, N67904,
         N67911, N67912, N67913, N67914, N67915, N67916, N67917, N67924,
         N67925, N67926, N67927, N67928, N67929, N67930, N67937, N67938,
         N67939, N67940, N67941, N67942, N67943, N67950, N67951, N67952,
         N67953, N67954, N67955, N67956, N67963, N67964, N67965, N67966,
         N67967, N67968, N67969, N67976, N67977, N67978, N67979, N67980,
         N67981, N67982, N67989, N67990, N67991, N67992, N67993, N67994,
         N67995, N68002, N68003, N68004, N68005, N68006, N68007, N68008,
         N68015, N68016, N68017, N68018, N68019, N68020, N68021, N68028,
         N68029, N68030, N68031, N68032, N68033, N68034, N68041, N68042,
         N68043, N68044, N68045, N68046, N68047, N68054, N68055, N68056,
         N68057, N68058, N68059, N68060, N68067, N68068, N68069, N68070,
         N68071, N68072, N68073, N68080, N68081, N68082, N68083, N68084,
         N68085, N68086, N68093, N68094, N68095, N68096, N68097, N68098,
         N68099, N68106, N68107, N68108, N68109, N68110, N68111, N68112,
         N68119, N68120, N68121, N68122, N68123, N68124, N68125, N68132,
         N68133, N68134, N68135, N68136, N68137, N68138, N68145, N68146,
         N68147, N68148, N68149, N68150, N68151, N68158, N68159, N68160,
         N68161, N68162, N68163, N68164, N68171, N68172, N68173, N68174,
         N68175, N68176, N68177, N68178, N68184, N68185, N68186, N68187,
         N68188, N68189, N68190, N68191, N68197, N68198, N68199, N68200,
         N68201, N68202, N68203, N68204, N68210, N68211, N68212, N68213,
         N68214, N68215, N68216, N68217, N68223, N68224, N68225, N68226,
         N68227, N68228, N68229, N68230, N68236, N68237, N68238, N68239,
         N68240, N68241, N68242, N68243, N68249, N68250, N68251, N68252,
         N68253, N68254, N68255, N68256, N68262, N68263, N68264, N68265,
         N68266, N68267, N68268, N68269, N68275, N68276, N68277, N68278,
         N68279, N68280, N68281, N68282, N68288, N68289, N68290, N68291,
         N68292, N68293, N68294, N68295, N68301, N68302, N68303, N68304,
         N68305, N68306, N68307, N68308, N68314, N68315, N68316, N68317,
         N68318, N68319, N68320, N68321, N68327, N68328, N68329, N68330,
         N68331, N68332, N68333, N68334, N68340, N68341, N68342, N68343,
         N68344, N68345, N68346, N68347, N68353, N68354, N68355, N68356,
         N68357, N68358, N68359, N68360, N68366, N68367, N68368, N68369,
         N68370, N68371, N68372, N68373, N68379, N68380, N68381, N68382,
         N68383, N68384, N68385, N68386, N68392, N68393, N68394, N68395,
         N68396, N68397, N68398, N68399, N68405, N68406, N68407, N68408,
         N68409, N68410, N68411, N68412, N68418, N68419, N68420, N68421,
         N68422, N68423, N68424, N68425, N68431, N68432, N68433, N68434,
         N68435, N68436, N68437, N68438, N68444, N68445, N68446, N68447,
         N68448, N68449, N68450, N68451, N68457, N68458, N68459, N68460,
         N68461, N68462, N68463, N68464, N68470, N68471, N68472, N68473,
         N68474, N68475, N68476, N68477, N68483, N68484, N68485, N68486,
         N68487, N68488, N68489, N68490, N68496, N68497, N68498, N68499,
         N68500, N68501, N68502, N68503, N68509, N68510, N68511, N68512,
         N68513, N68514, N68515, N68516, N68522, N68523, N68524, N68525,
         N68526, N68527, N68528, N68529, N68535, N68536, N68537, N68538,
         N68539, N68540, N68541, N68542, N68548, N68549, N68550, N68551,
         N68552, N68553, N68554, N68555, N68561, N68562, N68563, N68564,
         N68565, N68566, N68567, N68568, N68574, N68575, N68576, N68577,
         N68578, N68579, N68580, N68581, N68587, N68588, N68589, N68590,
         N68591, N68592, N68593, N68594, N68600, N68601, N68602, N68603,
         N68604, N68605, N68606, N68607, N68613, N68614, N68615, N68616,
         N68617, N68618, N68619, N68620, N68626, N68627, N68628, N68629,
         N68630, N68631, N68632, N68633, N68639, N68640, N68641, N68642,
         N68643, N68644, N68645, N68646, N68652, N68653, N68654, N68655,
         N68656, N68657, N68658, N68659, N68665, N68666, N68667, N68668,
         N68669, N68670, N68671, N68672, N68678, N68679, N68680, N68681,
         N68682, N68683, N68684, N68685, N68691, N68692, N68693, N68694,
         N68695, N68696, N68697, N68698, N68704, N68705, N68706, N68707,
         N68708, N68709, N68710, N68711, N68717, N68718, N68719, N68720,
         N68721, N68722, N68723, N68724, N68725, N68730, N68731, N68732,
         N68733, N68734, N68735, N68736, N68737, N68738, N68743, N68744,
         N68745, N68746, N68747, N68748, N68749, N68750, N68751, N68756,
         N68757, N68758, N68759, N68760, N68761, N68762, N68763, N68764,
         N68769, N68770, N68771, N68772, N68773, N68774, N68775, N68776,
         N68777, N68782, N68783, N68784, N68785, N68786, N68787, N68788,
         N68789, N68790, N68795, N68796, N68797, N68798, N68799, N68800,
         N68801, N68802, N68803, N68808, N68809, N68810, N68811, N68812,
         N68813, N68814, N68815, N68816, N68821, N68822, N68823, N68824,
         N68825, N68826, N68827, N68828, N68829, N68834, N68835, N68836,
         N68837, N68838, N68839, N68840, N68841, N68842, N68847, N68848,
         N68849, N68850, N68851, N68852, N68853, N68854, N68855, N68860,
         N68861, N68862, N68863, N68864, N68865, N68866, N68867, N68868,
         N68873, N68874, N68875, N68876, N68877, N68878, N68879, N68880,
         N68881, N68886, N68887, N68888, N68889, N68890, N68891, N68892,
         N68893, N68894, N68899, N68900, N68901, N68902, N68903, N68904,
         N68905, N68906, N68907, N68912, N68913, N68914, N68915, N68916,
         N68917, N68918, N68919, N68920, N68925, N68926, N68927, N68928,
         N68929, N68930, N68931, N68932, N68933, N68938, N68939, N68940,
         N68941, N68942, N68943, N68944, N68945, N68946, N68951, N68952,
         N68953, N68954, N68955, N68956, N68957, N68958, N68959, N68964,
         N68965, N68966, N68967, N68968, N68969, N68970, N68971, N68972,
         N68977, N68978, N68979, N68980, N68981, N68982, N68983, N68984,
         N68985, N68990, N68991, N68992, N68993, N68994, N68995, N68996,
         N68997, N68998, N68999, N69003, N69004, N69005, N69006, N69007,
         N69008, N69009, N69010, N69011, N69012, N69016, N69017, N69018,
         N69019, N69020, N69021, N69022, N69023, N69024, N69025, N69029,
         N69030, N69031, N69032, N69033, N69034, N69035, N69036, N69037,
         N69038, N69042, N69043, N69044, N69045, N69046, N69047, N69048,
         N69049, N69050, N69051, N69055, N69056, N69057, N69058, N69059,
         N69060, N69061, N69062, N69063, N69064, N69068, N69069, N69070,
         N69071, N69072, N69073, N69074, N69075, N69076, N69077, N69081,
         N69082, N69083, N69084, N69085, N69086, N69087, N69088, N69089,
         N69090, N69094, N69095, N69096, N69097, N69098, N69099, N69100,
         N69101, N69102, N69103, N69107, N69108, N69109, N69110, N69111,
         N69112, N69113, N69114, N69115, N69116, N69120, N69121, N69122,
         N69123, N69124, N69125, N69126, N69127, N69128, N69129, N69130,
         N69133, N69134, N69135, N69136, N69137, N69138, N69139, N69140,
         N69141, N69142, N69143, N69146, N69147, N69148, N69149, N69150,
         N69151, N69152, N69153, N69154, N69155, N69156, N69159, N69160,
         N69161, N69162, N69163, N69164, N69165, N69166, N69167, N69168,
         N69169, N69172, N69173, N69174, N69175, N69176, N69177, N69178,
         N69179, N69180, N69181, N69182, N69185, N69186, N69187, N69188,
         N69189, N69190, N69191, N69192, N69193, N69194, N69195, N69196,
         N69198, N69199, N69200, N69201, N69202, N69203, N69204, N69205,
         N69206, N69207, N69208, N69209, N69211, N69212, N69213, N69214,
         N69215, N69216, N69217, N69218, N69219, N69220, N69221, N69222,
         N69224, N69225, N69226, N69227, N69228, N69229, N69230, N69231,
         N69232, N69233, N69234, N69235, N69236, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
         n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
         n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
         n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
         n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
         n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
         n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
         n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
         n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
         n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
         n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
         n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603,
         n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
         n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
         n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
         n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731,
         n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
         n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
         n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
         n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
         n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
         n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
         n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
         n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
         n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
         n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
         n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
         n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
         n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
         n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123,
         n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
         n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
         n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
         n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
         n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
         n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
         n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
         n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411,
         n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
         n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
         n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
         n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
         n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
         n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
         n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
         n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
         n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683,
         n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
         n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699,
         n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
         n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875,
         n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
         n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
         n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
         n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
         n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
         n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
         n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
         n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
         n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
         n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
         n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
         n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
         n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
         n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
         n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
         n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
         n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
         n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
         n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
         n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
         n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
         n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
         n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
         n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
         n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547,
         n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
         n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
         n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643,
         n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
         n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
         n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667,
         n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
         n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
         n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691,
         n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
         n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707,
         n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715,
         n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723,
         n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
         n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739,
         n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747,
         n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
         n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763,
         n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
         n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779,
         n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
         n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
         n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
         n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811,
         n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819,
         n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
         n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835,
         n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
         n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851,
         n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
         n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
         n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
         n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883,
         n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891,
         n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
         n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907,
         n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915,
         n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923,
         n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931,
         n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
         n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
         n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955,
         n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963,
         n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971,
         n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979,
         n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
         n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995,
         n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003,
         n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
         n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
         n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027,
         n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035,
         n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043,
         n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
         n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
         n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
         n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
         n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
         n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
         n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099,
         n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107,
         n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
         n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
         n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131,
         n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
         n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147,
         n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155,
         n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
         n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171,
         n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
         n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187,
         n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195,
         n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
         n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211,
         n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219,
         n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227,
         n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235,
         n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243,
         n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251,
         n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259,
         n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267,
         n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275,
         n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283,
         n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291,
         n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299,
         n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307,
         n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315,
         n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323,
         n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331,
         n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339,
         n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347,
         n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355,
         n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363,
         n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371,
         n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379,
         n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387,
         n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395,
         n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403,
         n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411,
         n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419,
         n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427,
         n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435,
         n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443,
         n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451,
         n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459,
         n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467,
         n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475,
         n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483,
         n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491,
         n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499,
         n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507,
         n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515,
         n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523,
         n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531,
         n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539,
         n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547,
         n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555,
         n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563,
         n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571,
         n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579,
         n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587,
         n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595,
         n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603,
         n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611,
         n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619,
         n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627,
         n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635,
         n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643,
         n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651,
         n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659,
         n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667,
         n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675,
         n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683,
         n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691,
         n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699,
         n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707,
         n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715,
         n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723,
         n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731,
         n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739,
         n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747,
         n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755,
         n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763,
         n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771,
         n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779,
         n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787,
         n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795,
         n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803,
         n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811,
         n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819,
         n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827,
         n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835,
         n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843,
         n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851,
         n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859,
         n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867,
         n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875,
         n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883,
         n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891,
         n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899,
         n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907,
         n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915,
         n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923,
         n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931,
         n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939,
         n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947,
         n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955,
         n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963,
         n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971,
         n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979,
         n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987,
         n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995,
         n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003,
         n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011,
         n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019,
         n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027,
         n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035,
         n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043,
         n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051,
         n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059,
         n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067,
         n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075,
         n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083,
         n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091,
         n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099,
         n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107,
         n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115,
         n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123,
         n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131,
         n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139,
         n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147,
         n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155,
         n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163,
         n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171,
         n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179,
         n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187,
         n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195,
         n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203,
         n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211,
         n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219,
         n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227,
         n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235,
         n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243,
         n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251,
         n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259,
         n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267,
         n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275,
         n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283,
         n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291,
         n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299,
         n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307,
         n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315,
         n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323,
         n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331,
         n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339,
         n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347,
         n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355,
         n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363,
         n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371,
         n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379,
         n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387,
         n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395,
         n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403,
         n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411,
         n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419,
         n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427,
         n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435,
         n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443,
         n22444, n22445, n22446, n22447, n22448, n22449, n22450, n22451,
         n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459,
         n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467,
         n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475,
         n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483,
         n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491,
         n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499,
         n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507,
         n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515,
         n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523,
         n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531,
         n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539,
         n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547,
         n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555,
         n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563,
         n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571,
         n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579,
         n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587,
         n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595,
         n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603,
         n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611,
         n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619,
         n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627,
         n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635,
         n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643,
         n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651,
         n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659,
         n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667,
         n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675,
         n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683,
         n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691,
         n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699,
         n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707,
         n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715,
         n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723,
         n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731,
         n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739,
         n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747,
         n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755,
         n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763,
         n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771,
         n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779,
         n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787,
         n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795,
         n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803,
         n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811,
         n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819,
         n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827,
         n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835,
         n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843,
         n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851,
         n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859,
         n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867,
         n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875,
         n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883,
         n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891,
         n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899,
         n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907,
         n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915,
         n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923,
         n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931,
         n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939,
         n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947,
         n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955,
         n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963,
         n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971,
         n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979,
         n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987,
         n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995,
         n22996, n22997, n22998, n22999, n23000, n23001, n23002, n23003,
         n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011,
         n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019,
         n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027,
         n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035,
         n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043,
         n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051,
         n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059,
         n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067,
         n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075,
         n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083,
         n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091,
         n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099,
         n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107,
         n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115,
         n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123,
         n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131,
         n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139,
         n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147,
         n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155,
         n23156, n23157, n23158, n23159, n23160, n23161, n23162, n23163,
         n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171,
         n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179,
         n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187,
         n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195,
         n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23203,
         n23204, n23205, n23206, n23207, n23208, n23209, n23210, n23211,
         n23212, n23213, n23214, n23215, n23216, n23217, n23218, n23219,
         n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227,
         n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235,
         n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243,
         n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251,
         n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259,
         n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267,
         n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275,
         n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283,
         n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291,
         n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299,
         n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307,
         n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315,
         n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323,
         n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331,
         n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339,
         n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347,
         n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23355,
         n23356, n23357, n23358, n23359, n23360, n23361, n23362, n23363,
         n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371,
         n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379,
         n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387,
         n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395,
         n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403,
         n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411,
         n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419,
         n23420, n23421, n23422, n23423, n23424, n23425, n23426, n23427,
         n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435,
         n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443,
         n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451,
         n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459,
         n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467,
         n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475,
         n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483,
         n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491,
         n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499,
         n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507,
         n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515,
         n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523,
         n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531,
         n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539,
         n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547,
         n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555,
         n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563,
         n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571,
         n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579,
         n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587,
         n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595,
         n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603,
         n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611,
         n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619,
         n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627,
         n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635,
         n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643,
         n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651,
         n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659,
         n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667,
         n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675,
         n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683,
         n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691,
         n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699,
         n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707,
         n23708, n23709, n23710, n23711, n23712, n23713, n23714, n23715,
         n23716, n23717, n23718, n23719, n23720, n23721, n23722, n23723,
         n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731,
         n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739,
         n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747,
         n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755,
         n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763,
         n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771,
         n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779,
         n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787,
         n23788, n23789, n23790, n23791, n23792, n23793, n23794, n23795,
         n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803,
         n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811,
         n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819,
         n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827,
         n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835,
         n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843,
         n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23851,
         n23852, n23853, n23854, n23855, n23856, n23857, n23858, n23859,
         n23860, n23861, n23862, n23863, n23864, n23865, n23866, n23867,
         n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875,
         n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883,
         n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891,
         n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899,
         n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907,
         n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915,
         n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923,
         n23924, n23925, n23926, n23927, n23928, n23929, n23930, n23931,
         n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939,
         n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947,
         n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955,
         n23956, n23957, n23958, n23959, n23960, n23961, n23962, n23963,
         n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971,
         n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979,
         n23980, n23981, n23982, n23983, n23984, n23985, n23986, n23987,
         n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995,
         n23996, n23997, n23998, n23999, n24000, n24001, n24002, n24003,
         n24004, n24005, n24006, n24007, n24008, n24009, n24010, n24011,
         n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019,
         n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027,
         n24028, n24029, n24030, n24031, n24032, n24033, n24034, n24035,
         n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043,
         n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051,
         n24052, n24053, n24054, n24055, n24056, n24057, n24058, n24059,
         n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067,
         n24068, n24069, n24070, n24071, n24072, n24073, n24074, n24075,
         n24076, n24077, n24078, n24079, n24080, n24081, n24082, n24083,
         n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091,
         n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099,
         n24100, n24101, n24102, n24103, n24104, n24105, n24106, n24107,
         n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115,
         n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123,
         n24124, n24125, n24126, n24127, n24128, n24129, n24130, n24131,
         n24132, n24133, n24134, n24135, n24136, n24137, n24138, n24139,
         n24140, n24141, n24142, n24143, n24144, n24145, n24146, n24147,
         n24148, n24149, n24150, n24151, n24152, n24153, n24154, n24155,
         n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163,
         n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171,
         n24172, n24173, n24174, n24175, n24176, n24177, n24178, n24179,
         n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187,
         n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195,
         n24196, n24197, n24198, n24199, n24200, n24201, n24202, n24203,
         n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211,
         n24212, n24213, n24214, n24215, n24216, n24217, n24218, n24219,
         n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227,
         n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235,
         n24236, n24237, n24238, n24239, n24240, n24241, n24242, n24243,
         n24244, n24245, n24246, n24247, n24248, n24249, n24250, n24251,
         n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259,
         n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267,
         n24268, n24269, n24270, n24271, n24272, n24273, n24274, n24275,
         n24276, n24277, n24278, n24279, n24280, n24281, n24282, n24283,
         n24284, n24285, n24286, n24287, n24288, n24289, n24290, n24291,
         n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299,
         n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307,
         n24308, n24309, n24310, n24311, n24312, n24313, n24314, n24315,
         n24316, n24317, n24318, n24319, n24320, n24321, n24322, n24323,
         n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331,
         n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339,
         n24340, n24341, n24342, n24343, n24344, n24345, n24346, n24347,
         n24348, n24349, n24350, n24351, n24352, n24353, n24354, n24355,
         n24356, n24357, n24358, n24359, n24360, n24361, n24362, n24363,
         n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371,
         n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379,
         n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387,
         n24388, n24389, n24390, n24391, n24392, n24393, n24394, n24395,
         n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403,
         n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411,
         n24412, n24413, n24414, n24415, n24416, n24417, n24418, n24419,
         n24420, n24421, n24422, n24423, n24424, n24425, n24426, n24427,
         n24428, n24429, n24430, n24431, n24432, n24433, n24434, n24435,
         n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443,
         n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451,
         n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459,
         n24460, n24461, n24462, n24463, n24464, n24465, n24466, n24467,
         n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475,
         n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483,
         n24484, n24485, n24486, n24487, n24488, n24489, n24490, n24491,
         n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499,
         n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507,
         n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515,
         n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523,
         n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531,
         n24532, n24533, n24534, n24535, n24536, n24537, n24538, n24539,
         n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547,
         n24548, n24549, n24550, n24551, n24552, n24553, n24554, n24555,
         n24556, n24557, n24558, n24559, n24560, n24561, n24562, n24563,
         n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571,
         n24572, n24573, n24574, n24575, n24576, n24577, n24578, n24579,
         n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587,
         n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595,
         n24596, n24597, n24598, n24599, n24600, n24601, n24602, n24603,
         n24604, n24605, n24606, n24607, n24608, n24609, n24610, n24611,
         n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619,
         n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627,
         n24628, n24629, n24630, n24631, n24632, n24633, n24634, n24635,
         n24636, n24637, n24638, n24639, n24640, n24641, n24642, n24643,
         n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651,
         n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659,
         n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667,
         n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675,
         n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683,
         n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691,
         n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699,
         n24700, n24701, n24702, n24703, n24704, n24705, n24706, n24707,
         n24708, n24709, n24710, n24711, n24712, n24713, n24714, n24715,
         n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723,
         n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731,
         n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739,
         n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747,
         n24748, n24749, n24750, n24751, n24752, n24753, n24754, n24755,
         n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763,
         n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771,
         n24772, n24773, n24774, n24775, n24776, n24777, n24778, n24779,
         n24780, n24781, n24782, n24783, n24784, n24785, n24786, n24787,
         n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795,
         n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803,
         n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811,
         n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819,
         n24820, n24821, n24822, n24823, n24824, n24825, n24826, n24827,
         n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835,
         n24836, n24837, n24838, n24839, n24840, n24841, n24842, n24843,
         n24844, n24845, n24846, n24847, n24848, n24849, n24850, n24851,
         n24852, n24853, n24854, n24855, n24856, n24857, n24858, n24859,
         n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867,
         n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875,
         n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883,
         n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891,
         n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899,
         n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907,
         n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915,
         n24916, n24917, n24918, n24919, n24920, n24921, n24922, n24923,
         n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931,
         n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939,
         n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947,
         n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955,
         n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963,
         n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24971,
         n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979,
         n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987,
         n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995,
         n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003,
         n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011,
         n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019,
         n25020, n25021, n25022, n25023, n25024, n25025, n25026, n25027,
         n25028, n25029, n25030, n25031, n25032, n25033, n25034, n25035,
         n25036, n25037, n25038, n25039, n25040, n25041, n25042, n25043,
         n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25051,
         n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059,
         n25060, n25061, n25062, n25063, n25064, n25065, n25066, n25067,
         n25068, n25069, n25070, n25071, n25072, n25073, n25074, n25075,
         n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083,
         n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091,
         n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099,
         n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107,
         n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115,
         n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123,
         n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131,
         n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139,
         n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147,
         n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155,
         n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163,
         n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171,
         n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179,
         n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187,
         n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195,
         n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203,
         n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211,
         n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219,
         n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227,
         n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235,
         n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243,
         n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251,
         n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259,
         n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267,
         n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275,
         n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283,
         n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291,
         n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299,
         n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307,
         n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315,
         n25316, n25317, n25318, n25319, n25320, n25321, n25322, n25323,
         n25324, n25325, n25326, n25327, n25328, n25329, n25330, n25331,
         n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339,
         n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347,
         n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355,
         n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363,
         n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371,
         n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379,
         n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387,
         n25388, n25389, n25390, n25391, n25392, n25393, n25394, n25395,
         n25396, n25397, n25398, n25399, n25400, n25401, n25402, n25403,
         n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411,
         n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419,
         n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427,
         n25428, n25429, n25430, n25431, n25432, n25433, n25434, n25435,
         n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443,
         n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451,
         n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459,
         n25460, n25461, n25462, n25463, n25464, n25465, n25466, n25467,
         n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475,
         n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483,
         n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491,
         n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499,
         n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507,
         n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515,
         n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523,
         n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531,
         n25532, n25533, n25534, n25535, n25536, n25537, n25538, n25539,
         n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547,
         n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555,
         n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563,
         n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571,
         n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579,
         n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587,
         n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595,
         n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603,
         n25604, n25605, n25606, n25607, n25608, n25609, n25610, n25611,
         n25612, n25613, n25614, n25615, n25616, n25617, n25618, n25619,
         n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627,
         n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635,
         n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643,
         n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651,
         n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659,
         n25660, n25661, n25662, n25663, n25664, n25665, n25666, n25667,
         n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675,
         n25676, n25677, n25678, n25679, n25680, n25681, n25682, n25683,
         n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691,
         n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699,
         n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707,
         n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715,
         n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723,
         n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731,
         n25732, n25733, n25734, n25735, n25736, n25737, n25738, n25739,
         n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747,
         n25748, n25749, n25750, n25751, n25752, n25753, n25754, n25755,
         n25756, n25757, n25758, n25759, n25760, n25761, n25762, n25763,
         n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771,
         n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779,
         n25780, n25781, n25782, n25783, n25784, n25785, n25786, n25787,
         n25788, n25789, n25790, n25791, n25792, n25793, n25794, n25795,
         n25796, n25797, n25798, n25799, n25800, n25801, n25802, n25803,
         n25804, n25805, n25806, n25807, n25808, n25809, n25810, n25811,
         n25812, n25813, n25814, n25815, n25816, n25817, n25818, n25819,
         n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827,
         n25828, n25829, n25830, n25831, n25832, n25833, n25834, n25835,
         n25836, n25837, n25838, n25839, n25840, n25841, n25842, n25843,
         n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851,
         n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859,
         n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867,
         n25868, n25869, n25870, n25871, n25872, n25873, n25874, n25875,
         n25876, n25877, n25878, n25879, n25880, n25881, n25882, n25883,
         n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891,
         n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899,
         n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907,
         n25908, n25909, n25910, n25911, n25912, n25913, n25914, n25915,
         n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923,
         n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931,
         n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939,
         n25940, n25941, n25942, n25943, n25944, n25945, n25946, n25947,
         n25948, n25949, n25950, n25951, n25952, n25953, n25954, n25955,
         n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963,
         n25964, n25965, n25966, n25967, n25968, n25969, n25970, n25971,
         n25972, n25973, n25974, n25975, n25976, n25977, n25978, n25979,
         n25980, n25981, n25982, n25983, n25984, n25985, n25986, n25987,
         n25988, n25989, n25990, n25991, n25992, n25993, n25994, n25995,
         n25996, n25997, n25998, n25999, n26000, n26001, n26002, n26003,
         n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011,
         n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26019,
         n26020, n26021, n26022, n26023, n26024, n26025, n26026, n26027,
         n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035,
         n26036, n26037, n26038, n26039, n26040, n26041, n26042, n26043,
         n26044, n26045, n26046, n26047, n26048, n26049, n26050, n26051,
         n26052, n26053, n26054, n26055, n26056, n26057, n26058, n26059,
         n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067,
         n26068, n26069, n26070, n26071, n26072, n26073, n26074, n26075,
         n26076, n26077, n26078, n26079, n26080, n26081, n26082, n26083,
         n26084, n26085, n26086, n26087, n26088, n26089, n26090, n26091,
         n26092, n26093, n26094, n26095, n26096, n26097, n26098, n26099,
         n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26107,
         n26108, n26109, n26110, n26111, n26112, n26113, n26114, n26115,
         n26116, n26117, n26118, n26119, n26120, n26121, n26122, n26123,
         n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131,
         n26132, n26133, n26134, n26135, n26136, n26137, n26138, n26139,
         n26140, n26141, n26142, n26143, n26144, n26145, n26146, n26147,
         n26148, n26149, n26150, n26151, n26152, n26153, n26154, n26155,
         n26156, n26157, n26158, n26159, n26160, n26161, n26162, n26163,
         n26164, n26165, n26166, n26167, n26168, n26169, n26170, n26171,
         n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26179,
         n26180, n26181, n26182, n26183, n26184, n26185, n26186, n26187,
         n26188, n26189, n26190, n26191, n26192, n26193, n26194, n26195,
         n26196, n26197, n26198, n26199, n26200, n26201, n26202, n26203,
         n26204, n26205, n26206, n26207, n26208, n26209, n26210, n26211,
         n26212, n26213, n26214, n26215, n26216, n26217, n26218, n26219,
         n26220, n26221, n26222, n26223, n26224, n26225, n26226, n26227,
         n26228, n26229, n26230, n26231, n26232, n26233, n26234, n26235,
         n26236, n26237, n26238, n26239, n26240, n26241, n26242, n26243,
         n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251,
         n26252, n26253, n26254, n26255, n26256, n26257, n26258, n26259,
         n26260, n26261, n26262, n26263, n26264, n26265, n26266, n26267,
         n26268, n26269, n26270, n26271, n26272, n26273, n26274, n26275,
         n26276, n26277, n26278, n26279, n26280, n26281, n26282, n26283,
         n26284, n26285, n26286, n26287, n26288, n26289, n26290, n26291,
         n26292, n26293, n26294, n26295, n26296, n26297, n26298, n26299,
         n26300, n26301, n26302, n26303, n26304, n26305, n26306, n26307,
         n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315,
         n26316, n26317, n26318, n26319, n26320, n26321, n26322, n26323,
         n26324, n26325, n26326, n26327, n26328, n26329, n26330, n26331,
         n26332, n26333, n26334, n26335, n26336, n26337, n26338, n26339,
         n26340, n26341, n26342, n26343, n26344, n26345, n26346, n26347,
         n26348, n26349, n26350, n26351, n26352, n26353, n26354, n26355,
         n26356, n26357, n26358, n26359, n26360, n26361, n26362, n26363,
         n26364, n26365, n26366, n26367, n26368, n26369, n26370, n26371,
         n26372, n26373, n26374, n26375, n26376, n26377, n26378, n26379,
         n26380, n26381, n26382, n26383, n26384, n26385, n26386, n26387,
         n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395,
         n26396, n26397, n26398, n26399, n26400, n26401, n26402, n26403,
         n26404, n26405, n26406, n26407, n26408, n26409, n26410, n26411,
         n26412, n26413, n26414, n26415, n26416, n26417, n26418, n26419,
         n26420, n26421, n26422, n26423, n26424, n26425, n26426, n26427,
         n26428, n26429, n26430, n26431, n26432, n26433, n26434, n26435,
         n26436, n26437, n26438, n26439, n26440, n26441, n26442, n26443,
         n26444, n26445, n26446, n26447, n26448, n26449, n26450, n26451,
         n26452, n26453, n26454, n26455, n26456, n26457, n26458, n26459,
         n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467,
         n26468, n26469, n26470, n26471, n26472, n26473, n26474, n26475,
         n26476, n26477, n26478, n26479, n26480, n26481, n26482, n26483,
         n26484, n26485, n26486, n26487, n26488, n26489, n26490, n26491,
         n26492, n26493, n26494, n26495, n26496, n26497, n26498, n26499,
         n26500, n26501, n26502, n26503, n26504, n26505, n26506, n26507,
         n26508, n26509, n26510, n26511, n26512, n26513, n26514, n26515,
         n26516, n26517, n26518, n26519, n26520, n26521, n26522, n26523,
         n26524, n26525, n26526, n26527, n26528, n26529, n26530, n26531,
         n26532, n26533, n26534, n26535, n26536, n26537, n26538, n26539,
         n26540, n26541, n26542, n26543, n26544, n26545, n26546, n26547,
         n26548, n26549, n26550, n26551, n26552, n26553, n26554, n26555,
         n26556, n26557, n26558, n26559, n26560, n26561, n26562, n26563,
         n26564, n26565, n26566, n26567, n26568, n26569, n26570, n26571,
         n26572, n26573, n26574, n26575, n26576, n26577, n26578, n26579,
         n26580, n26581, n26582, n26583, n26584, n26585, n26586, n26587,
         n26588, n26589, n26590, n26591, n26592, n26593, n26594, n26595,
         n26596, n26597, n26598, n26599, n26600, n26601, n26602, n26603,
         n26604, n26605, n26606, n26607, n26608, n26609, n26610, n26611,
         n26612, n26613, n26614, n26615, n26616, n26617, n26618, n26619,
         n26620, n26621, n26622, n26623, n26624, n26625, n26626, n26627,
         n26628, n26629, n26630, n26631, n26632, n26633, n26634, n26635,
         n26636, n26637, n26638, n26639, n26640, n26641, n26642, n26643,
         n26644, n26645, n26646, n26647, n26648, n26649, n26650, n26651,
         n26652, n26653, n26654, n26655, n26656, n26657, n26658, n26659,
         n26660, n26661, n26662, n26663, n26664, n26665, n26666, n26667,
         n26668, n26669, n26670, n26671, n26672, n26673, n26674, n26675,
         n26676, n26677, n26678, n26679, n26680, n26681, n26682, n26683,
         n26684, n26685, n26686, n26687, n26688, n26689, n26690, n26691,
         n26692, n26693, n26694, n26695, n26696, n26697, n26698, n26699,
         n26700, n26701, n26702, n26703, n26704, n26705, n26706, n26707,
         n26708, n26709, n26710, n26711, n26712, n26713, n26714, n26715,
         n26716, n26717, n26718, n26719, n26720, n26721, n26722, n26723,
         n26724, n26725, n26726, n26727, n26728, n26729, n26730, n26731,
         n26732, n26733, n26734, n26735, n26736, n26737, n26738, n26739,
         n26740, n26741, n26742, n26743, n26744, n26745, n26746, n26747,
         n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755,
         n26756, n26757, n26758, n26759, n26760, n26761, n26762, n26763,
         n26764, n26765, n26766, n26767, n26768, n26769, n26770, n26771,
         n26772, n26773, n26774, n26775, n26776, n26777, n26778, n26779,
         n26780, n26781, n26782, n26783, n26784, n26785, n26786, n26787,
         n26788, n26789, n26790, n26791, n26792, n26793, n26794, n26795,
         n26796, n26797, n26798, n26799, n26800, n26801, n26802, n26803,
         n26804, n26805, n26806, n26807, n26808, n26809, n26810, n26811,
         n26812, n26813, n26814, n26815, n26816, n26817, n26818, n26819,
         n26820, n26821, n26822, n26823, n26824, n26825, n26826, n26827,
         n26828, n26829, n26830, n26831, n26832, n26833, n26834, n26835,
         n26836, n26837, n26838, n26839, n26840, n26841, n26842, n26843,
         n26844, n26845, n26846, n26847, n26848, n26849, n26850, n26851,
         n26852, n26853, n26854, n26855, n26856, n26857, n26858, n26859,
         n26860, n26861, n26862, n26863, n26864, n26865, n26866, n26867,
         n26868, n26869, n26870, n26871, n26872, n26873, n26874, n26875,
         n26876, n26877, n26878, n26879, n26880, n26881, n26882, n26883,
         n26884, n26885, n26886, n26887, n26888, n26889, n26890, n26891,
         n26892, n26893, n26894, n26895, n26896, n26897, n26898, n26899,
         n26900, n26901, n26902, n26903, n26904, n26905, n26906, n26907,
         n26908, n26909, n26910, n26911, n26912, n26913, n26914, n26915,
         n26916, n26917, n26918, n26919, n26920, n26921, n26922, n26923,
         n26924, n26925, n26926, n26927, n26928, n26929, n26930, n26931,
         n26932, n26933, n26934, n26935, n26936, n26937, n26938, n26939,
         n26940, n26941, n26942, n26943, n26944, n26945, n26946, n26947,
         n26948, n26949, n26950, n26951, n26952, n26953, n26954, n26955,
         n26956, n26957, n26958, n26959, n26960, n26961, n26962, n26963,
         n26964, n26965, n26966, n26967, n26968, n26969, n26970, n26971,
         n26972, n26973, n26974, n26975, n26976, n26977, n26978, n26979,
         n26980, n26981, n26982, n26983, n26984, n26985, n26986, n26987,
         n26988, n26989, n26990, n26991, n26992, n26993, n26994, n26995,
         n26996, n26997, n26998, n26999, n27000, n27001, n27002, n27003,
         n27004, n27005, n27006, n27007, n27008, n27009, n27010, n27011,
         n27012, n27013, n27014, n27015, n27016, n27017, n27018, n27019,
         n27020, n27021, n27022, n27023, n27024, n27025, n27026, n27027,
         n27028, n27029, n27030, n27031, n27032, n27033, n27034, n27035,
         n27036, n27037, n27038, n27039, n27040, n27041, n27042, n27043,
         n27044, n27045, n27046, n27047, n27048, n27049, n27050, n27051,
         n27052, n27053, n27054, n27055, n27056, n27057, n27058, n27059,
         n27060, n27061, n27062, n27063, n27064, n27065, n27066, n27067,
         n27068, n27069, n27070, n27071, n27072, n27073, n27074, n27075,
         n27076, n27077, n27078, n27079, n27080, n27081, n27082, n27083,
         n27084, n27085, n27086, n27087, n27088, n27089, n27090, n27091,
         n27092, n27093, n27094, n27095, n27096, n27097, n27098, n27099,
         n27100, n27101, n27102, n27103, n27104, n27105, n27106, n27107,
         n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115,
         n27116, n27117, n27118, n27119, n27120, n27121, n27122, n27123,
         n27124, n27125, n27126, n27127, n27128, n27129, n27130, n27131,
         n27132, n27133, n27134, n27135, n27136, n27137, n27138, n27139,
         n27140, n27141, n27142, n27143, n27144, n27145, n27146, n27147,
         n27148, n27149, n27150, n27151, n27152, n27153, n27154, n27155,
         n27156, n27157, n27158, n27159, n27160, n27161, n27162, n27163,
         n27164, n27165, n27166, n27167, n27168, n27169, n27170, n27171,
         n27172, n27173, n27174, n27175, n27176, n27177, n27178, n27179,
         n27180, n27181, n27182, n27183, n27184, n27185, n27186, n27187,
         n27188, n27189, n27190, n27191, n27192, n27193, n27194, n27195,
         n27196, n27197, n27198, n27199, n27200, n27201, n27202, n27203,
         n27204, n27205, n27206, n27207, n27208, n27209, n27210, n27211,
         n27212, n27213, n27214, n27215, n27216, n27217, n27218, n27219,
         n27220, n27221, n27222, n27223, n27224, n27225, n27226, n27227,
         n27228, n27229, n27230, n27231, n27232, n27233, n27234, n27235,
         n27236, n27237, n27238, n27239, n27240, n27241, n27242, n27243,
         n27244, n27245, n27246, n27247, n27248, n27249, n27250, n27251,
         n27252, n27253, n27254, n27255, n27256, n27257, n27258, n27259,
         n27260, n27261, n27262, n27263, n27264, n27265, n27266, n27267,
         n27268, n27269, n27270, n27271, n27272, n27273, n27274, n27275,
         n27276, n27277, n27278, n27279, n27280, n27281, n27282, n27283,
         n27284, n27285, n27286, n27287, n27288, n27289, n27290, n27291,
         n27292, n27293, n27294, n27295, n27296, n27297, n27298, n27299,
         n27300, n27301, n27302, n27303, n27304, n27305, n27306, n27307,
         n27308, n27309, n27310, n27311, n27312, n27313, n27314, n27315,
         n27316, n27317, n27318, n27319, n27320, n27321, n27322, n27323,
         n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331,
         n27332, n27333, n27334, n27335, n27336, n27337, n27338, n27339,
         n27340, n27341, n27342, n27343, n27344, n27345, n27346, n27347,
         n27348, n27349, n27350, n27351, n27352, n27353, n27354, n27355,
         n27356, n27357, n27358, n27359, n27360, n27361, n27362, n27363,
         n27364, n27365, n27366, n27367, n27368, n27369, n27370, n27371,
         n27372, n27373, n27374, n27375, n27376, n27377, n27378, n27379,
         n27380, n27381, n27382, n27383, n27384, n27385, n27386, n27387,
         n27388, n27389, n27390, n27391, n27392, n27393, n27394, n27395,
         n27396, n27397, n27398, n27399, n27400, n27401, n27402, n27403,
         n27404, n27405, n27406, n27407, n27408, n27409, n27410, n27411,
         n27412, n27413, n27414, n27415, n27416, n27417, n27418, n27419,
         n27420, n27421, n27422, n27423, n27424, n27425, n27426, n27427,
         n27428, n27429, n27430, n27431, n27432, n27433, n27434, n27435,
         n27436, n27437, n27438, n27439, n27440, n27441, n27442, n27443,
         n27444, n27445, n27446, n27447, n27448, n27449, n27450, n27451,
         n27452, n27453, n27454, n27455, n27456, n27457, n27458, n27459,
         n27460, n27461, n27462, n27463, n27464, n27465, n27466, n27467,
         n27468, n27469, n27470, n27471, n27472, n27473, n27474, n27475,
         n27476, n27477, n27478, n27479, n27480, n27481, n27482, n27483,
         n27484, n27485, n27486, n27487, n27488, n27489, n27490, n27491,
         n27492, n27493, n27494, n27495, n27496, n27497, n27498, n27499,
         n27500, n27501, n27502, n27503, n27504, n27505, n27506, n27507,
         n27508, n27509, n27510, n27511, n27512, n27513, n27514, n27515,
         n27516, n27517, n27518, n27519, n27520, n27521, n27522, n27523,
         n27524, n27525, n27526, n27527, n27528, n27529, n27530, n27531,
         n27532, n27533, n27534, n27535, n27536, n27537, n27538, n27539,
         n27540, n27541, n27542, n27543, n27544, n27545, n27546, n27547,
         n27548, n27549, n27550, n27551, n27552, n27553, n27554, n27555,
         n27556, n27557, n27558, n27559, n27560, n27561, n27562, n27563,
         n27564, n27565, n27566, n27567, n27568, n27569, n27570, n27571,
         n27572, n27573, n27574, n27575, n27576, n27577, n27578, n27579,
         n27580, n27581, n27582, n27583, n27584, n27585, n27586, n27587,
         n27588, n27589, n27590, n27591, n27592, n27593, n27594, n27595,
         n27596, n27597, n27598, n27599, n27600, n27601, n27602, n27603,
         n27604, n27605, n27606, n27607, n27608, n27609, n27610, n27611,
         n27612, n27613, n27614, n27615, n27616, n27617, n27618, n27619,
         n27620, n27621, n27622, n27623, n27624, n27625, n27626, n27627,
         n27628, n27629, n27630, n27631, n27632, n27633, n27634, n27635,
         n27636, n27637, n27638, n27639, n27640, n27641, n27642, n27643,
         n27644, n27645, n27646, n27647, n27648, n27649, n27650, n27651,
         n27652, n27653, n27654, n27655, n27656, n27657, n27658, n27659,
         n27660, n27661, n27662, n27663, n27664, n27665, n27666, n27667,
         n27668, n27669, n27670, n27671, n27672, n27673, n27674, n27675,
         n27676, n27677, n27678, n27679, n27680, n27681, n27682, n27683,
         n27684, n27685, n27686, n27687, n27688, n27689, n27690, n27691,
         n27692, n27693, n27694, n27695, n27696, n27697, n27698, n27699,
         n27700, n27701, n27702, n27703, n27704, n27705, n27706, n27707,
         n27708, n27709, n27710, n27711, n27712, n27713, n27714, n27715,
         n27716, n27717, n27718, n27719, n27720, n27721, n27722, n27723,
         n27724, n27725, n27726, n27727, n27728, n27729, n27730, n27731,
         n27732, n27733, n27734, n27735, n27736, n27737, n27738, n27739,
         n27740, n27741, n27742, n27743, n27744, n27745, n27746, n27747,
         n27748, n27749, n27750, n27751, n27752, n27753, n27754, n27755,
         n27756, n27757, n27758, n27759, n27760, n27761, n27762, n27763,
         n27764, n27765, n27766, n27767, n27768, n27769, n27770, n27771,
         n27772, n27773, n27774, n27775, n27776, n27777, n27778, n27779,
         n27780, n27781, n27782, n27783, n27784, n27785, n27786, n27787,
         n27788, n27789, n27790, n27791, n27792, n27793, n27794, n27795,
         n27796, n27797, n27798, n27799, n27800, n27801, n27802, n27803,
         n27804, n27805, n27806, n27807, n27808, n27809, n27810, n27811,
         n27812, n27813, n27814, n27815, n27816, n27817, n27818, n27819,
         n27820, n27821, n27822, n27823, n27824, n27825, n27826, n27827,
         n27828, n27829, n27830, n27831, n27832, n27833, n27834, n27835,
         n27836, n27837, n27838, n27839, n27840, n27841, n27842, n27843,
         n27844, n27845, n27846, n27847, n27848, n27849, n27850, n27851,
         n27852, n27853, n27854, n27855, n27856, n27857, n27858, n27859,
         n27860, n27861, n27862, n27863, n27864, n27865, n27866, n27867,
         n27868, n27869, n27870, n27871, n27872, n27873, n27874, n27875,
         n27876, n27877, n27878, n27879, n27880, n27881, n27882, n27883,
         n27884, n27885, n27886, n27887, n27888, n27889, n27890, n27891,
         n27892, n27893, n27894, n27895, n27896, n27897, n27898, n27899,
         n27900, n27901, n27902, n27903, n27904, n27905, n27906, n27907,
         n27908, n27909, n27910, n27911, n27912, n27913, n27914, n27915,
         n27916, n27917, n27918, n27919, n27920, n27921, n27922, n27923,
         n27924, n27925, n27926, n27927, n27928, n27929, n27930, n27931,
         n27932, n27933, n27934, n27935, n27936, n27937, n27938, n27939,
         n27940, n27941, n27942, n27943, n27944, n27945, n27946, n27947,
         n27948, n27949, n27950, n27951, n27952, n27953, n27954, n27955,
         n27956, n27957, n27958, n27959, n27960, n27961, n27962, n27963,
         n27964, n27965, n27966, n27967, n27968, n27969, n27970, n27971,
         n27972, n27973, n27974, n27975, n27976, n27977, n27978, n27979,
         n27980, n27981, n27982, n27983, n27984, n27985, n27986, n27987,
         n27988, n27989, n27990, n27991, n27992, n27993, n27994, n27995,
         n27996, n27997, n27998, n27999, n28000, n28001, n28002, n28003,
         n28004, n28005, n28006, n28007, n28008, n28009, n28010, n28011,
         n28012, n28013, n28014, n28015, n28016, n28017, n28018, n28019,
         n28020, n28021, n28022, n28023, n28024, n28025, n28026, n28027,
         n28028, n28029, n28030, n28031, n28032, n28033, n28034, n28035,
         n28036, n28037, n28038, n28039, n28040, n28041, n28042, n28043,
         n28044, n28045, n28046, n28047, n28048, n28049, n28050, n28051,
         n28052, n28053, n28054, n28055, n28056, n28057, n28058, n28059,
         n28060, n28061, n28062, n28063, n28064, n28065, n28066, n28067,
         n28068, n28069, n28070, n28071, n28072, n28073, n28074, n28075,
         n28076, n28077, n28078, n28079, n28080, n28081, n28082, n28083,
         n28084, n28085, n28086, n28087, n28088, n28089, n28090, n28091,
         n28092, n28093, n28094, n28095, n28096, n28097, n28098, n28099,
         n28100, n28101, n28102, n28103, n28104, n28105, n28106, n28107,
         n28108, n28109, n28110, n28111, n28112, n28113, n28114, n28115,
         n28116, n28117, n28118, n28119, n28120, n28121, n28122, n28123,
         n28124, n28125, n28126, n28127, n28128, n28129, n28130, n28131,
         n28132, n28133, n28134, n28135, n28136, n28137, n28138, n28139,
         n28140, n28141, n28142, n28143, n28144, n28145, n28146, n28147,
         n28148, n28149, n28150, n28151, n28152, n28153, n28154, n28155,
         n28156, n28157, n28158, n28159, n28160, n28161, n28162, n28163,
         n28164, n28165, n28166, n28167, n28168, n28169, n28170, n28171,
         n28172, n28173, n28174, n28175, n28176, n28177, n28178, n28179,
         n28180, n28181, n28182, n28183, n28184, n28185, n28186, n28187,
         n28188, n28189, n28190, n28191, n28192, n28193, n28194, n28195,
         n28196, n28197, n28198, n28199, n28200, n28201, n28202, n28203,
         n28204, n28205, n28206, n28207, n28208, n28209, n28210, n28211,
         n28212, n28213, n28214, n28215, n28216, n28217, n28218, n28219,
         n28220, n28221, n28222, n28223, n28224, n28225, n28226, n28227,
         n28228, n28229, n28230, n28231, n28232, n28233, n28234, n28235,
         n28236, n28237, n28238, n28239, n28240, n28241, n28242, n28243,
         n28244, n28245, n28246, n28247, n28248, n28249, n28250, n28251,
         n28252, n28253, n28254, n28255, n28256, n28257, n28258, n28259,
         n28260, n28261, n28262, n28263, n28264, n28265, n28266, n28267,
         n28268, n28269, n28270, n28271, n28272, n28273, n28274, n28275,
         n28276, n28277, n28278, n28279, n28280, n28281, n28282, n28283,
         n28284, n28285, n28286, n28287, n28288, n28289, n28290, n28291,
         n28292, n28293, n28294, n28295, n28296, n28297, n28298, n28299,
         n28300, n28301, n28302, n28303, n28304, n28305, n28306, n28307,
         n28308, n28309, n28310, n28311, n28312, n28313, n28314, n28315,
         n28316, n28317, n28318, n28319, n28320, n28321, n28322, n28323,
         n28324, n28325, n28326, n28327, n28328, n28329, n28330, n28331,
         n28332, n28333, n28334, n28335, n28336, n28337, n28338, n28339,
         n28340, n28341, n28342, n28343, n28344, n28345, n28346, n28347,
         n28348, n28349, n28350, n28351, n28352, n28353, n28354, n28355,
         n28356, n28357, n28358, n28359, n28360, n28361, n28362, n28363,
         n28364, n28365, n28366, n28367, n28368, n28369, n28370, n28371,
         n28372, n28373, n28374, n28375, n28376, n28377, n28378, n28379,
         n28380, n28381, n28382, n28383, n28384, n28385, n28386, n28387,
         n28388, n28389, n28390, n28391, n28392, n28393, n28394, n28395,
         n28396, n28397, n28398, n28399, n28400, n28401, n28402, n28403,
         n28404, n28405, n28406, n28407, n28408, n28409, n28410, n28411,
         n28412, n28413, n28414, n28415, n28416, n28417, n28418, n28419,
         n28420, n28421, n28422, n28423, n28424, n28425, n28426, n28427,
         n28428, n28429, n28430, n28431, n28432, n28433, n28434, n28435,
         n28436, n28437, n28438, n28439, n28440, n28441, n28442, n28443,
         n28444, n28445, n28446, n28447, n28448, n28449, n28450, n28451,
         n28452, n28453, n28454, n28455, n28456, n28457, n28458, n28459,
         n28460, n28461, n28462, n28463, n28464, n28465, n28466, n28467,
         n28468, n28469, n28470, n28471, n28472, n28473, n28474, n28475,
         n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483,
         n28484, n28485, n28486, n28487, n28488, n28489, n28490, n28491,
         n28492, n28493, n28494, n28495, n28496, n28497, n28498, n28499,
         n28500, n28501, n28502, n28503, n28504, n28505, n28506, n28507,
         n28508, n28509, n28510, n28511, n28512, n28513, n28514, n28515,
         n28516, n28517, n28518, n28519, n28520, n28521, n28522, n28523,
         n28524, n28525, n28526, n28527, n28528, n28529, n28530, n28531,
         n28532, n28533, n28534, n28535, n28536, n28537, n28538, n28539,
         n28540, n28541, n28542, n28543, n28544, n28545, n28546, n28547,
         n28548, n28549, n28550, n28551, n28552, n28553, n28554, n28555,
         n28556, n28557, n28558, n28559, n28560, n28561, n28562, n28563,
         n28564, n28565, n28566, n28567, n28568, n28569, n28570, n28571,
         n28572, n28573, n28574, n28575, n28576, n28577, n28578, n28579,
         n28580, n28581, n28582, n28583, n28584, n28585, n28586, n28587,
         n28588, n28589, n28590, n28591, n28592, n28593, n28594, n28595,
         n28596, n28597, n28598, n28599, n28600, n28601, n28602, n28603,
         n28604, n28605, n28606, n28607, n28608, n28609, n28610, n28611,
         n28612, n28613, n28614, n28615, n28616, n28617, n28618, n28619,
         n28620, n28621, n28622, n28623, n28624, n28625, n28626, n28627,
         n28628, n28629, n28630, n28631, n28632, n28633, n28634, n28635,
         n28636, n28637, n28638, n28639, n28640, n28641, n28642, n28643,
         n28644, n28645, n28646, n28647, n28648, n28649, n28650, n28651,
         n28652, n28653, n28654, n28655, n28656, n28657, n28658, n28659,
         n28660, n28661, n28662, n28663, n28664, n28665, n28666, n28667,
         n28668, n28669, n28670, n28671, n28672, n28673, n28674, n28675,
         n28676, n28677, n28678, n28679, n28680, n28681, n28682, n28683,
         n28684, n28685, n28686, n28687, n28688, n28689, n28690, n28691,
         n28692, n28693, n28694, n28695, n28696, n28697, n28698, n28699,
         n28700, n28701, n28702, n28703, n28704, n28705, n28706, n28707,
         n28708, n28709, n28710, n28711, n28712, n28713, n28714, n28715,
         n28716, n28717, n28718, n28719, n28720, n28721, n28722, n28723,
         n28724, n28725, n28726, n28727, n28728, n28729, n28730, n28731,
         n28732, n28733, n28734, n28735, n28736, n28737, n28738, n28739,
         n28740, n28741, n28742, n28743, n28744, n28745, n28746, n28747,
         n28748, n28749, n28750, n28751, n28752, n28753, n28754, n28755,
         n28756, n28757, n28758, n28759, n28760, n28761, n28762, n28763,
         n28764, n28765, n28766, n28767, n28768, n28769, n28770, n28771,
         n28772, n28773, n28774, n28775, n28776, n28777, n28778, n28779,
         n28780, n28781, n28782, n28783, n28784, n28785, n28786, n28787,
         n28788, n28789, n28790, n28791, n28792, n28793, n28794, n28795,
         n28796, n28797, n28798, n28799, n28800, n28801, n28802, n28803,
         n28804, n28805, n28806, n28807, n28808, n28809, n28810, n28811,
         n28812, n28813, n28814, n28815, n28816, n28817, n28818, n28819,
         n28820, n28821, n28822, n28823, n28824, n28825, n28826, n28827,
         n28828, n28829, n28830, n28831, n28832, n28833, n28834, n28835,
         n28836, n28837, n28838, n28839, n28840, n28841, n28842, n28843,
         n28844, n28845, n28846, n28847, n28848, n28849, n28850, n28851,
         n28852, n28853, n28854, n28855, n28856, n28857, n28858, n28859,
         n28860, n28861, n28862, n28863, n28864, n28865, n28866, n28867,
         n28868, n28869, n28870, n28871, n28872, n28873, n28874, n28875,
         n28876, n28877, n28878, n28879, n28880, n28881, n28882, n28883,
         n28884, n28885, n28886, n28887, n28888, n28889, n28890, n28891,
         n28892, n28893, n28894, n28895, n28896, n28897, n28898, n28899,
         n28900, n28901, n28902, n28903, n28904, n28905, n28906, n28907,
         n28908, n28909, n28910, n28911, n28912, n28913, n28914, n28915,
         n28916, n28917, n28918, n28919, n28920, n28921, n28922, n28923,
         n28924, n28925, n28926, n28927, n28928, n28929, n28930, n28931,
         n28932, n28933, n28934, n28935, n28936, n28937, n28938, n28939,
         n28940, n28941, n28942, n28943, n28944, n28945, n28946, n28947,
         n28948, n28949, n28950, n28951, n28952, n28953, n28954, n28955,
         n28956, n28957, n28958, n28959, n28960, n28961, n28962, n28963,
         n28964, n28965, n28966, n28967, n28968, n28969, n28970, n28971,
         n28972, n28973, n28974, n28975, n28976, n28977, n28978, n28979,
         n28980, n28981, n28982, n28983, n28984, n28985, n28986, n28987,
         n28988, n28989, n28990, n28991, n28992, n28993, n28994, n28995,
         n28996, n28997, n28998, n28999, n29000, n29001, n29002, n29003,
         n29004, n29005, n29006, n29007, n29008, n29009, n29010, n29011,
         n29012, n29013, n29014, n29015, n29016, n29017, n29018, n29019,
         n29020, n29021, n29022, n29023, n29024, n29025, n29026, n29027,
         n29028, n29029, n29030, n29031, n29032, n29033, n29034, n29035,
         n29036, n29037, n29038, n29039, n29040, n29041, n29042, n29043,
         n29044, n29045, n29046, n29047, n29048, n29049, n29050, n29051,
         n29052, n29053, n29054, n29055, n29056, n29057, n29058, n29059,
         n29060, n29061, n29062, n29063, n29064, n29065, n29066, n29067,
         n29068, n29069, n29070, n29071, n29072, n29073, n29074, n29075,
         n29076, n29077, n29078, n29079, n29080, n29081, n29082, n29083,
         n29084, n29085, n29086, n29087, n29088, n29089, n29090, n29091,
         n29092, n29093, n29094, n29095, n29096, n29097, n29098, n29099,
         n29100, n29101, n29102, n29103, n29104, n29105, n29106, n29107,
         n29108, n29109, n29110, n29111, n29112, n29113, n29114, n29115,
         n29116, n29117, n29118, n29119, n29120, n29121, n29122, n29123,
         n29124, n29125, n29126, n29127, n29128, n29129, n29130, n29131,
         n29132, n29133, n29134, n29135, n29136, n29137, n29138, n29139,
         n29140, n29141, n29142, n29143, n29144, n29145, n29146, n29147,
         n29148, n29149, n29150, n29151, n29152, n29153, n29154, n29155,
         n29156, n29157, n29158, n29159, n29160, n29161, n29162, n29163,
         n29164, n29165, n29166, n29167, n29168, n29169, n29170, n29171,
         n29172, n29173, n29174, n29175, n29176, n29177, n29178, n29179,
         n29180, n29181, n29182, n29183, n29184, n29185, n29186, n29187,
         n29188, n29189, n29190, n29191, n29192, n29193, n29194, n29195,
         n29196, n29197, n29198, n29199, n29200, n29201, n29202, n29203,
         n29204, n29205, n29206, n29207, n29208, n29209, n29210, n29211,
         n29212, n29213, n29214, n29215, n29216, n29217, n29218, n29219,
         n29220, n29221, n29222, n29223, n29224, n29225, n29226, n29227,
         n29228, n29229, n29230, n29231, n29232, n29233, n29234, n29235,
         n29236, n29237, n29238, n29239, n29240, n29241, n29242, n29243,
         n29244, n29245, n29246, n29247, n29248, n29249, n29250, n29251,
         n29252, n29253, n29254, n29255, n29256, n29257, n29258, n29259,
         n29260, n29261, n29262, n29263, n29264, n29265, n29266, n29267,
         n29268, n29269, n29270, n29271, n29272, n29273, n29274, n29275,
         n29276, n29277, n29278, n29279, n29280, n29281, n29282, n29283,
         n29284, n29285, n29286, n29287, n29288, n29289, n29290, n29291,
         n29292, n29293, n29294, n29295, n29296, n29297, n29298, n29299,
         n29300, n29301, n29302, n29303, n29304, n29305, n29306, n29307,
         n29308, n29309, n29310, n29311, n29312, n29313, n29314, n29315,
         n29316, n29317, n29318, n29319, n29320, n29321, n29322, n29323,
         n29324, n29325, n29326, n29327, n29328, n29329, n29330, n29331,
         n29332, n29333, n29334, n29335, n29336, n29337, n29338, n29339,
         n29340, n29341, n29342, n29343, n29344, n29345, n29346, n29347,
         n29348, n29349, n29350, n29351, n29352, n29353, n29354, n29355,
         n29356, n29357, n29358, n29359, n29360, n29361, n29362, n29363,
         n29364, n29365, n29366, n29367, n29368, n29369, n29370, n29371,
         n29372, n29373, n29374, n29375, n29376, n29377, n29378, n29379,
         n29380, n29381, n29382, n29383, n29384, n29385, n29386, n29387,
         n29388, n29389, n29390, n29391, n29392, n29393, n29394, n29395,
         n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403,
         n29404, n29405, n29406, n29407, n29408, n29409, n29410, n29411,
         n29412, n29413, n29414, n29415, n29416, n29417, n29418, n29419,
         n29420, n29421, n29422, n29423, n29424, n29425, n29426, n29427,
         n29428, n29429, n29430, n29431, n29432, n29433, n29434, n29435,
         n29436, n29437, n29438, n29439, n29440, n29441, n29442, n29443,
         n29444, n29445, n29446, n29447, n29448, n29449, n29450, n29451,
         n29452, n29453, n29454, n29455, n29456, n29457, n29458, n29459,
         n29460, n29461, n29462, n29463, n29464, n29465, n29466, n29467,
         n29468, n29469, n29470, n29471, n29472, n29473, n29474, n29475,
         n29476, n29477, n29478, n29479, n29480, n29481, n29482, n29483,
         n29484, n29485, n29486, n29487, n29488, n29489, n29490, n29491,
         n29492, n29493, n29494, n29495, n29496, n29497, n29498, n29499,
         n29500, n29501, n29502, n29503, n29504, n29505, n29506, n29507,
         n29508, n29509, n29510, n29511, n29512, n29513, n29514, n29515,
         n29516, n29517, n29518, n29519, n29520, n29521, n29522, n29523,
         n29524, n29525, n29526, n29527, n29528, n29529, n29530, n29531,
         n29532, n29533, n29534, n29535, n29536, n29537, n29538, n29539,
         n29540, n29541, n29542, n29543, n29544, n29545, n29546, n29547,
         n29548, n29549, n29550, n29551, n29552, n29553, n29554, n29555,
         n29556, n29557, n29558, n29559, n29560, n29561, n29562, n29563,
         n29564, n29565, n29566, n29567, n29568, n29569, n29570, n29571,
         n29572, n29573, n29574, n29575, n29576, n29577, n29578, n29579,
         n29580, n29581, n29582, n29583, n29584, n29585, n29586, n29587,
         n29588, n29589, n29590, n29591, n29592, n29593, n29594, n29595,
         n29596, n29597, n29598, n29599, n29600, n29601, n29602, n29603,
         n29604, n29605, n29606, n29607, n29608, n29609, n29610, n29611,
         n29612, n29613, n29614, n29615, n29616, n29617, n29618, n29619,
         n29620, n29621, n29622, n29623, n29624, n29625, n29626, n29627,
         n29628, n29629, n29630, n29631, n29632, n29633, n29634, n29635,
         n29636, n29637, n29638, n29639, n29640, n29641, n29642, n29643,
         n29644, n29645, n29646, n29647, n29648, n29649, n29650, n29651,
         n29652, n29653, n29654, n29655, n29656, n29657, n29658, n29659,
         n29660, n29661, n29662, n29663, n29664, n29665, n29666, n29667,
         n29668, n29669, n29670, n29671, n29672, n29673, n29674, n29675,
         n29676, n29677, n29678, n29679, n29680, n29681, n29682, n29683,
         n29684, n29685, n29686, n29687, n29688, n29689, n29690, n29691,
         n29692, n29693, n29694, n29695, n29696, n29697, n29698, n29699,
         n29700, n29701, n29702, n29703, n29704, n29705, n29706, n29707,
         n29708, n29709, n29710, n29711, n29712, n29713, n29714, n29715,
         n29716, n29717, n29718, n29719, n29720, n29721, n29722, n29723,
         n29724, n29725, n29726, n29727, n29728, n29729, n29730, n29731,
         n29732, n29733, n29734, n29735, n29736, n29737, n29738, n29739,
         n29740, n29741, n29742, n29743, n29744, n29745, n29746, n29747,
         n29748, n29749, n29750, n29751, n29752, n29753, n29754, n29755,
         n29756, n29757, n29758, n29759, n29760, n29761, n29762, n29763,
         n29764, n29765, n29766, n29767, n29768, n29769, n29770, n29771,
         n29772, n29773, n29774, n29775, n29776, n29777, n29778, n29779,
         n29780, n29781, n29782, n29783, n29784, n29785, n29786, n29787,
         n29788, n29789, n29790, n29791, n29792, n29793, n29794, n29795,
         n29796, n29797, n29798, n29799, n29800, n29801, n29802, n29803,
         n29804, n29805, n29806, n29807, n29808, n29809, n29810, n29811,
         n29812, n29813, n29814, n29815, n29816, n29817, n29818, n29819,
         n29820, n29821, n29822, n29823, n29824, n29825, n29826, n29827,
         n29828, n29829, n29830, n29831, n29832, n29833, n29834, n29835,
         n29836, n29837, n29838, n29839, n29840, n29841, n29842, n29843,
         n29844, n29845, n29846, n29847, n29848, n29849, n29850, n29851,
         n29852, n29853, n29854, n29855, n29856, n29857, n29858, n29859,
         n29860, n29861, n29862, n29863, n29864, n29865, n29866, n29867,
         n29868, n29869, n29870, n29871, n29872, n29873, n29874, n29875,
         n29876, n29877, n29878, n29879, n29880, n29881, n29882, n29883,
         n29884, n29885, n29886, n29887, n29888, n29889, n29890, n29891,
         n29892, n29893, n29894, n29895, n29896, n29897, n29898, n29899,
         n29900, n29901, n29902, n29903, n29904, n29905, n29906, n29907,
         n29908, n29909, n29910, n29911, n29912, n29913, n29914, n29915,
         n29916, n29917, n29918, n29919, n29920, n29921, n29922, n29923,
         n29924, n29925, n29926, n29927, n29928, n29929, n29930, n29931,
         n29932, n29933, n29934, n29935, n29936, n29937, n29938, n29939,
         n29940, n29941, n29942, n29943, n29944, n29945, n29946, n29947,
         n29948, n29949, n29950, n29951, n29952, n29953, n29954, n29955,
         n29956, n29957, n29958, n29959, n29960, n29961, n29962, n29963,
         n29964, n29965, n29966, n29967, n29968, n29969, n29970, n29971,
         n29972, n29973, n29974, n29975, n29976, n29977, n29978, n29979,
         n29980, n29981, n29982, n29983, n29984, n29985, n29986, n29987,
         n29988, n29989, n29990, n29991, n29992, n29993, n29994, n29995,
         n29996, n29997, n29998, n29999, n30000, n30001, n30002, n30003,
         n30004, n30005, n30006, n30007, n30008, n30009, n30010, n30011,
         n30012, n30013, n30014, n30015, n30016, n30017, n30018, n30019,
         n30020, n30021, n30022, n30023, n30024, n30025, n30026, n30027,
         n30028, n30029, n30030, n30031, n30032, n30033, n30034, n30035,
         n30036, n30037, n30038, n30039, n30040, n30041, n30042, n30043,
         n30044, n30045, n30046, n30047, n30048, n30049, n30050, n30051,
         n30052, n30053, n30054, n30055, n30056, n30057, n30058, n30059,
         n30060, n30061, n30062, n30063, n30064, n30065, n30066, n30067,
         n30068, n30069, n30070, n30071, n30072, n30073, n30074, n30075,
         n30076, n30077, n30078, n30079, n30080, n30081, n30082, n30083,
         n30084, n30085, n30086, n30087, n30088, n30089, n30090, n30091,
         n30092, n30093, n30094, n30095, n30096, n30097, n30098, n30099,
         n30100, n30101, n30102, n30103, n30104, n30105, n30106, n30107,
         n30108, n30109, n30110, n30111, n30112, n30113, n30114, n30115,
         n30116, n30117, n30118, n30119, n30120, n30121, n30122, n30123,
         n30124, n30125, n30126, n30127, n30128, n30129, n30130, n30131,
         n30132, n30133, n30134, n30135, n30136, n30137, n30138, n30139,
         n30140, n30141, n30142, n30143, n30144, n30145, n30146, n30147,
         n30148, n30149, n30150, n30151, n30152, n30153, n30154, n30155,
         n30156, n30157, n30158, n30159, n30160, n30161, n30162, n30163,
         n30164, n30165, n30166, n30167, n30168, n30169, n30170, n30171,
         n30172, n30173, n30174, n30175, n30176, n30177, n30178, n30179,
         n30180, n30181, n30182, n30183, n30184, n30185, n30186, n30187,
         n30188, n30189, n30190, n30191, n30192, n30193, n30194, n30195,
         n30196, n30197, n30198, n30199, n30200, n30201, n30202, n30203,
         n30204, n30205, n30206, n30207, n30208, n30209, n30210, n30211,
         n30212, n30213, n30214, n30215, n30216, n30217, n30218, n30219,
         n30220, n30221, n30222, n30223, n30224, n30225, n30226, n30227,
         n30228, n30229, n30230, n30231, n30232, n30233, n30234, n30235,
         n30236, n30237, n30238, n30239, n30240, n30241, n30242, n30243,
         n30244, n30245, n30246, n30247, n30248, n30249, n30250, n30251,
         n30252, n30253, n30254, n30255, n30256, n30257, n30258, n30259,
         n30260, n30261, n30262, n30263, n30264, n30265, n30266, n30267,
         n30268, n30269, n30270, n30271, n30272, n30273, n30274, n30275,
         n30276, n30277, n30278, n30279, n30280, n30281, n30282, n30283,
         n30284, n30285, n30286, n30287, n30288, n30289, n30290, n30291,
         n30292, n30293, n30294, n30295, n30296, n30297, n30298, n30299,
         n30300, n30301, n30302, n30303, n30304, n30305, n30306, n30307,
         n30308, n30309, n30310, n30311, n30312, n30313, n30314, n30315,
         n30316, n30317, n30318, n30319, n30320, n30321, n30322, n30323,
         n30324, n30325, n30326, n30327, n30328, n30329, n30330, n30331,
         n30332, n30333, n30334, n30335, n30336, n30337, n30338, n30339,
         n30340, n30341, n30342, n30343, n30344, n30345, n30346, n30347,
         n30348, n30349, n30350, n30351, n30352, n30353, n30354, n30355,
         n30356, n30357, n30358, n30359, n30360, n30361, n30362, n30363,
         n30364, n30365, n30366, n30367, n30368, n30369, n30370, n30371,
         n30372, n30373, n30374, n30375, n30376, n30377, n30378, n30379,
         n30380, n30381, n30382, n30383, n30384, n30385, n30386, n30387,
         n30388, n30389, n30390, n30391, n30392, n30393, n30394, n30395,
         n30396, n30397, n30398, n30399, n30400, n30401, n30402, n30403,
         n30404, n30405, n30406, n30407, n30408, n30409, n30410, n30411,
         n30412, n30413, n30414, n30415, n30416, n30417, n30418, n30419,
         n30420, n30421, n30422, n30423, n30424, n30425, n30426, n30427,
         n30428, n30429, n30430, n30431, n30432, n30433, n30434, n30435,
         n30436, n30437, n30438, n30439, n30440, n30441, n30442, n30443,
         n30444, n30445, n30446, n30447, n30448, n30449, n30450, n30451,
         n30452, n30453, n30454, n30455, n30456, n30457, n30458, n30459,
         n30460, n30461, n30462, n30463, n30464, n30465, n30466, n30467,
         n30468, n30469, n30470, n30471, n30472, n30473, n30474, n30475,
         n30476, n30477, n30478, n30479, n30480, n30481, n30482, n30483,
         n30484, n30485, n30486, n30487, n30488, n30489, n30490, n30491,
         n30492, n30493, n30494, n30495, n30496, n30497, n30498, n30499,
         n30500, n30501, n30502, n30503, n30504, n30505, n30506, n30507,
         n30508, n30509, n30510, n30511, n30512, n30513, n30514, n30515,
         n30516, n30517, n30518, n30519, n30520, n30521, n30522, n30523,
         n30524, n30525, n30526, n30527, n30528, n30529, n30530, n30531,
         n30532, n30533, n30534, n30535, n30536, n30537, n30538, n30539,
         n30540, n30541, n30542, n30543, n30544, n30545, n30546, n30547,
         n30548, n30549, n30550, n30551, n30552, n30553, n30554, n30555,
         n30556, n30557, n30558, n30559, n30560, n30561, n30562, n30563,
         n30564, n30565, n30566, n30567, n30568, n30569, n30570, n30571,
         n30572, n30573, n30574, n30575, n30576, n30577, n30578, n30579,
         n30580, n30581, n30582, n30583, n30584, n30585, n30586, n30587,
         n30588, n30589, n30590, n30591, n30592, n30593, n30594, n30595,
         n30596, n30597, n30598, n30599, n30600, n30601, n30602, n30603,
         n30604, n30605, n30606, n30607, n30608, n30609, n30610, n30611,
         n30612, n30613, n30614, n30615, n30616, n30617, n30618, n30619,
         n30620, n30621, n30622, n30623, n30624, n30625, n30626, n30627,
         n30628, n30629, n30630, n30631, n30632, n30633, n30634, n30635,
         n30636, n30637, n30638, n30639, n30640, n30641, n30642, n30643,
         n30644, n30645, n30646, n30647, n30648, n30649, n30650, n30651,
         n30652, n30653, n30654, n30655, n30656, n30657, n30658, n30659,
         n30660, n30661, n30662, n30663, n30664, n30665, n30666, n30667,
         n30668, n30669, n30670, n30671, n30672, n30673, n30674, n30675,
         n30676, n30677, n30678, n30679, n30680, n30681, n30682, n30683,
         n30684, n30685, n30686, n30687, n30688, n30689, n30690, n30691,
         n30692, n30693, n30694, n30695, n30696, n30697, n30698, n30699,
         n30700, n30701, n30702, n30703, n30704, n30705, n30706, n30707,
         n30708, n30709, n30710, n30711, n30712, n30713, n30714, n30715,
         n30716, n30717, n30718, n30719, n30720, n30721, n30722, n30723,
         n30724, n30725, n30726, n30727, n30728, n30729, n30730, n30731,
         n30732, n30733, n30734, n30735, n30736, n30737, n30738, n30739,
         n30740, n30741, n30742, n30743, n30744, n30745, n30746, n30747,
         n30748, n30749, n30750, n30751, n30752, n30753, n30754, n30755,
         n30756, n30757, n30758, n30759, n30760, n30761, n30762, n30763,
         n30764, n30765, n30766, n30767, n30768, n30769, n30770, n30771,
         n30772, n30773, n30774, n30775, n30776, n30777, n30778, n30779,
         n30780, n30781, n30782, n30783, n30784, n30785, n30786, n30787,
         n30788, n30789, n30790, n30791, n30792, n30793, n30794, n30795,
         n30796, n30797, n30798, n30799, n30800, n30801, n30802, n30803,
         n30804, n30805, n30806, n30807, n30808, n30809, n30810, n30811,
         n30812, n30813, n30814, n30815, n30816, n30817, n30818, n30819,
         n30820, n30821, n30822, n30823, n30824, n30825, n30826, n30827,
         n30828, n30829, n30830, n30831, n30832, n30833, n30834, n30835,
         n30836, n30837, n30838, n30839, n30840, n30841, n30842, n30843,
         n30844, n30845, n30846, n30847, n30848, n30849, n30850, n30851,
         n30852, n30853, n30854, n30855, n30856, n30857, n30858, n30859,
         n30860, n30861, n30862, n30863, n30864, n30865, n30866, n30867,
         n30868, n30869, n30870, n30871, n30872, n30873, n30874, n30875,
         n30876, n30877, n30878, n30879, n30880, n30881, n30882, n30883,
         n30884, n30885, n30886, n30887, n30888, n30889, n30890, n30891,
         n30892, n30893, n30894, n30895, n30896, n30897, n30898, n30899,
         n30900, n30901, n30902, n30903, n30904, n30905, n30906, n30907,
         n30908, n30909, n30910, n30911, n30912, n30913, n30914, n30915,
         n30916, n30917, n30918, n30919, n30920, n30921, n30922, n30923,
         n30924, n30925, n30926, n30927, n30928, n30929, n30930, n30931,
         n30932, n30933, n30934, n30935, n30936, n30937, n30938, n30939,
         n30940, n30941, n30942, n30943, n30944, n30945, n30946, n30947,
         n30948, n30949, n30950, n30951, n30952, n30953, n30954, n30955,
         n30956, n30957, n30958, n30959, n30960, n30961, n30962, n30963,
         n30964, n30965, n30966, n30967, n30968, n30969, n30970, n30971,
         n30972, n30973, n30974, n30975, n30976, n30977, n30978, n30979,
         n30980, n30981, n30982, n30983, n30984, n30985, n30986, n30987,
         n30988, n30989, n30990, n30991, n30992, n30993, n30994, n30995,
         n30996, n30997, n30998, n30999, n31000, n31001, n31002, n31003,
         n31004, n31005, n31006, n31007, n31008, n31009, n31010, n31011,
         n31012, n31013, n31014, n31015, n31016, n31017, n31018, n31019,
         n31020, n31021, n31022, n31023, n31024, n31025, n31026, n31027,
         n31028, n31029, n31030, n31031, n31032, n31033, n31034, n31035,
         n31036, n31037, n31038, n31039, n31040, n31041, n31042, n31043,
         n31044, n31045, n31046, n31047, n31048, n31049, n31050, n31051,
         n31052, n31053, n31054, n31055, n31056, n31057, n31058, n31059,
         n31060, n31061, n31062, n31063, n31064, n31065, n31066, n31067,
         n31068, n31069, n31070, n31071, n31072, n31073, n31074, n31075,
         n31076, n31077, n31078, n31079, n31080, n31081, n31082, n31083,
         n31084, n31085, n31086, n31087, n31088, n31089, n31090, n31091,
         n31092, n31093, n31094, n31095, n31096, n31097, n31098, n31099,
         n31100, n31101, n31102, n31103, n31104, n31105, n31106, n31107,
         n31108, n31109, n31110, n31111, n31112, n31113, n31114, n31115,
         n31116, n31117, n31118, n31119, n31120, n31121, n31122, n31123,
         n31124, n31125, n31126, n31127, n31128, n31129, n31130, n31131,
         n31132, n31133, n31134, n31135, n31136, n31137, n31138, n31139,
         n31140, n31141, n31142, n31143, n31144, n31145, n31146, n31147,
         n31148, n31149, n31150, n31151, n31152, n31153, n31154, n31155,
         n31156, n31157, n31158, n31159, n31160, n31161, n31162, n31163,
         n31164, n31165, n31166, n31167, n31168, n31169, n31170, n31171,
         n31172, n31173, n31174, n31175, n31176, n31177, n31178, n31179,
         n31180, n31181, n31182, n31183, n31184, n31185, n31186, n31187,
         n31188, n31189, n31190, n31191, n31192, n31193, n31194, n31195,
         n31196, n31197, n31198, n31199, n31200, n31201, n31202, n31203,
         n31204, n31205, n31206, n31207, n31208, n31209, n31210, n31211,
         n31212, n31213, n31214, n31215, n31216, n31217, n31218, n31219,
         n31220, n31221, n31222, n31223, n31224, n31225, n31226, n31227,
         n31228, n31229, n31230, n31231, n31232, n31233, n31234, n31235,
         n31236, n31237, n31238, n31239, n31240, n31241, n31242, n31243,
         n31244, n31245, n31246, n31247, n31248, n31249, n31250, n31251,
         n31252, n31253, n31254, n31255, n31256, n31257, n31258, n31259,
         n31260, n31261, n31262, n31263, n31264, n31265, n31266, n31267,
         n31268, n31269, n31270, n31271, n31272, n31273, n31274, n31275,
         n31276, n31277, n31278, n31279, n31280, n31281, n31282, n31283,
         n31284, n31285, n31286, n31287, n31288, n31289, n31290, n31291,
         n31292, n31293, n31294, n31295, n31296, n31297, n31298, n31299,
         n31300, n31301, n31302, n31303, n31304, n31305, n31306, n31307,
         n31308, n31309, n31310, n31311, n31312, n31313, n31314, n31315,
         n31316, n31317, n31318, n31319, n31320, n31321, n31322, n31323,
         n31324, n31325, n31326, n31327, n31328, n31329, n31330, n31331,
         n31332, n31333, n31334, n31335, n31336, n31337, n31338, n31339,
         n31340, n31341, n31342, n31343, n31344, n31345, n31346, n31347,
         n31348, n31349, n31350, n31351, n31352, n31353, n31354, n31355,
         n31356, n31357, n31358, n31359, n31360, n31361, n31362, n31363,
         n31364, n31365, n31366, n31367, n31368, n31369, n31370, n31371,
         n31372, n31373, n31374, n31375, n31376, n31377, n31378, n31379,
         n31380, n31381, n31382, n31383, n31384, n31385, n31386, n31387,
         n31388, n31389, n31390, n31391, n31392, n31393, n31394, n31395,
         n31396, n31397, n31398, n31399, n31400, n31401, n31402, n31403,
         n31404, n31405, n31406, n31407, n31408, n31409, n31410, n31411,
         n31412, n31413, n31414, n31415, n31416, n31417, n31418, n31419,
         n31420, n31421, n31422, n31423, n31424, n31425, n31426, n31427,
         n31428, n31429, n31430, n31431, n31432, n31433, n31434, n31435,
         n31436, n31437, n31438, n31439, n31440, n31441, n31442, n31443,
         n31444, n31445, n31446, n31447, n31448, n31449, n31450, n31451,
         n31452, n31453, n31454, n31455, n31456, n31457, n31458, n31459,
         n31460, n31461, n31462, n31463, n31464, n31465, n31466, n31467,
         n31468, n31469, n31470, n31471, n31472, n31473, n31474, n31475,
         n31476, n31477, n31478, n31479, n31480, n31481, n31482, n31483,
         n31484, n31485, n31486, n31487, n31488, n31489, n31490, n31491,
         n31492, n31493, n31494, n31495, n31496, n31497, n31498, n31499,
         n31500, n31501, n31502, n31503, n31504, n31505, n31506, n31507,
         n31508, n31509, n31510, n31511, n31512, n31513, n31514, n31515,
         n31516, n31517, n31518, n31519, n31520, n31521, n31522, n31523,
         n31524, n31525, n31526, n31527, n31528, n31529, n31530, n31531,
         n31532, n31533, n31534, n31535, n31536, n31537, n31538, n31539,
         n31540, n31541, n31542, n31543, n31544, n31545, n31546, n31547,
         n31548, n31549, n31550, n31551, n31552, n31553, n31554, n31555,
         n31556, n31557, n31558, n31559, n31560, n31561, n31562, n31563,
         n31564, n31565, n31566, n31567, n31568, n31569, n31570, n31571,
         n31572, n31573, n31574, n31575, n31576, n31577, n31578, n31579,
         n31580, n31581, n31582, n31583, n31584, n31585, n31586, n31587,
         n31588, n31589, n31590, n31591, n31592, n31593, n31594, n31595,
         n31596, n31597, n31598, n31599, n31600, n31601, n31602, n31603,
         n31604, n31605, n31606, n31607, n31608, n31609, n31610, n31611,
         n31612, n31613, n31614, n31615, n31616, n31617, n31618, n31619,
         n31620, n31621, n31622, n31623, n31624, n31625, n31626, n31627,
         n31628, n31629, n31630, n31631, n31632, n31633, n31634, n31635,
         n31636, n31637, n31638, n31639, n31640, n31641, n31642, n31643,
         n31644, n31645, n31646, n31647, n31648, n31649, n31650, n31651,
         n31652, n31653, n31654, n31655, n31656, n31657, n31658, n31659,
         n31660, n31661, n31662, n31663, n31664, n31665, n31666, n31667,
         n31668, n31669, n31670, n31671, n31672, n31673, n31674, n31675,
         n31676, n31677, n31678, n31679, n31680, n31681, n31682, n31683,
         n31684, n31685, n31686, n31687, n31688, n31689, n31690, n31691,
         n31692, n31693, n31694, n31695, n31696, n31697, n31698, n31699,
         n31700, n31701, n31702, n31703, n31704, n31705, n31706, n31707,
         n31708, n31709, n31710, n31711, n31712, n31713, n31714, n31715,
         n31716, n31717, n31718, n31719, n31720, n31721, n31722, n31723,
         n31724, n31725, n31726, n31727, n31728, n31729, n31730, n31731,
         n31732, n31733, n31734, n31735, n31736, n31737, n31738, n31739,
         n31740, n31741, n31742, n31743, n31744, n31745, n31746, n31747,
         n31748, n31749, n31750, n31751, n31752, n31753, n31754, n31755,
         n31756, n31757, n31758, n31759, n31760, n31761, n31762, n31763,
         n31764, n31765, n31766, n31767, n31768, n31769, n31770, n31771,
         n31772, n31773, n31774, n31775, n31776, n31777, n31778, n31779,
         n31780, n31781, n31782, n31783, n31784, n31785, n31786, n31787,
         n31788, n31789, n31790, n31791, n31792, n31793, n31794, n31795,
         n31796, n31797, n31798, n31799, n31800, n31801, n31802, n31803,
         n31804, n31805, n31806, n31807, n31808, n31809, n31810, n31811,
         n31812, n31813, n31814, n31815, n31816, n31817, n31818, n31819,
         n31820, n31821, n31822, n31823, n31824, n31825, n31826, n31827,
         n31828, n31829, n31830, n31831, n31832, n31833, n31834, n31835,
         n31836, n31837, n31838, n31839, n31840, n31841, n31842, n31843,
         n31844, n31845, n31846, n31847, n31848, n31849, n31850, n31851,
         n31852, n31853, n31854, n31855, n31856, n31857, n31858, n31859,
         n31860, n31861, n31862, n31863, n31864, n31865, n31866, n31867,
         n31868, n31869, n31870, n31871, n31872, n31873, n31874, n31875,
         n31876, n31877, n31878, n31879, n31880, n31881, n31882, n31883,
         n31884, n31885, n31886, n31887, n31888, n31889, n31890, n31891,
         n31892, n31893, n31894, n31895, n31896, n31897, n31898, n31899,
         n31900, n31901, n31902, n31903, n31904, n31905, n31906, n31907,
         n31908, n31909, n31910, n31911, n31912, n31913, n31914, n31915,
         n31916, n31917, n31918, n31919, n31920, n31921, n31922, n31923,
         n31924, n31925, n31926, n31927, n31928, n31929, n31930, n31931,
         n31932, n31933, n31934, n31935, n31936, n31937, n31938, n31939,
         n31940, n31941, n31942, n31943, n31944, n31945, n31946, n31947,
         n31948, n31949, n31950, n31951, n31952, n31953, n31954, n31955,
         n31956, n31957, n31958, n31959, n31960, n31961, n31962, n31963,
         n31964, n31965, n31966, n31967, n31968, n31969, n31970, n31971,
         n31972, n31973, n31974, n31975, n31976, n31977, n31978, n31979,
         n31980, n31981, n31982, n31983, n31984, n31985, n31986, n31987,
         n31988, n31989, n31990, n31991, n31992, n31993, n31994, n31995,
         n31996, n31997, n31998, n31999, n32000, n32001, n32002, n32003,
         n32004, n32005, n32006, n32007, n32008, n32009, n32010, n32011,
         n32012, n32013, n32014, n32015, n32016, n32017, n32018, n32019,
         n32020, n32021, n32022, n32023, n32024, n32025, n32026, n32027,
         n32028, n32029, n32030, n32031, n32032, n32033, n32034, n32035,
         n32036, n32037, n32038, n32039, n32040, n32041, n32042, n32043,
         n32044, n32045, n32046, n32047, n32048, n32049, n32050, n32051,
         n32052, n32053, n32054, n32055, n32056, n32057, n32058, n32059,
         n32060, n32061, n32062, n32063, n32064, n32065, n32066, n32067,
         n32068, n32069, n32070, n32071, n32072, n32073, n32074, n32075,
         n32076, n32077, n32078, n32079, n32080, n32081, n32082, n32083,
         n32084, n32085, n32086, n32087, n32088, n32089, n32090, n32091,
         n32092, n32093, n32094, n32095, n32096, n32097, n32098, n32099,
         n32100, n32101, n32102, n32103, n32104, n32105, n32106, n32107,
         n32108, n32109, n32110, n32111, n32112, n32113, n32114, n32115,
         n32116, n32117, n32118, n32119, n32120, n32121, n32122, n32123,
         n32124, n32125, n32126, n32127, n32128, n32129, n32130, n32131,
         n32132, n32133, n32134, n32135, n32136, n32137, n32138, n32139,
         n32140, n32141, n32142, n32143, n32144, n32145, n32146, n32147,
         n32148, n32149, n32150, n32151, n32152, n32153, n32154, n32155,
         n32156, n32157, n32158, n32159, n32160, n32161, n32162, n32163,
         n32164, n32165, n32166, n32167, n32168, n32169, n32170, n32171,
         n32172, n32173, n32174, n32175, n32176, n32177, n32178, n32179,
         n32180, n32181, n32182, n32183, n32184, n32185, n32186, n32187,
         n32188, n32189, n32190, n32191, n32192, n32193, n32194, n32195,
         n32196, n32197, n32198, n32199, n32200, n32201, n32202, n32203,
         n32204, n32205, n32206, n32207, n32208, n32209, n32210, n32211,
         n32212, n32213, n32214, n32215, n32216, n32217, n32218, n32219,
         n32220, n32221, n32222, n32223, n32224, n32225, n32226, n32227,
         n32228, n32229, n32230, n32231, n32232, n32233, n32234, n32235,
         n32236, n32237, n32238, n32239, n32240, n32241, n32242, n32243,
         n32244, n32245, n32246, n32247, n32248, n32249, n32250, n32251,
         n32252, n32253, n32254, n32255, n32256, n32257, n32258, n32259,
         n32260, n32261, n32262, n32263, n32264, n32265, n32266, n32267,
         n32268, n32269, n32270, n32271, n32272, n32273, n32274, n32275,
         n32276, n32277, n32278, n32279, n32280, n32281, n32282, n32283,
         n32284, n32285, n32286, n32287, n32288, n32289, n32290, n32291,
         n32292, n32293, n32294, n32295, n32296, n32297, n32298, n32299,
         n32300, n32301, n32302, n32303, n32304, n32305, n32306, n32307,
         n32308, n32309, n32310, n32311, n32312, n32313, n32314, n32315,
         n32316, n32317, n32318, n32319, n32320, n32321, n32322, n32323,
         n32324, n32325, n32326, n32327, n32328, n32329, n32330, n32331,
         n32332, n32333, n32334, n32335, n32336, n32337, n32338, n32339,
         n32340, n32341, n32342, n32343, n32344, n32345, n32346, n32347,
         n32348, n32349, n32350, n32351, n32352, n32353, n32354, n32355,
         n32356, n32357, n32358, n32359, n32360, n32361, n32362, n32363,
         n32364, n32365, n32366, n32367, n32368, n32369, n32370, n32371,
         n32372, n32373, n32374, n32375, n32376, n32377, n32378, n32379,
         n32380, n32381, n32382, n32383, n32384, n32385, n32386, n32387,
         n32388, n32389, n32390, n32391, n32392, n32393, n32394, n32395,
         n32396, n32397, n32398, n32399, n32400, n32401, n32402, n32403,
         n32404, n32405, n32406, n32407, n32408, n32409, n32410, n32411,
         n32412, n32413, n32414, n32415, n32416, n32417, n32418, n32419,
         n32420, n32421, n32422, n32423, n32424, n32425, n32426, n32427,
         n32428, n32429, n32430, n32431, n32432, n32433, n32434, n32435,
         n32436, n32437, n32438, n32439, n32440, n32441, n32442, n32443,
         n32444, n32445, n32446, n32447, n32448, n32449, n32450, n32451,
         n32452, n32453, n32454, n32455, n32456, n32457, n32458, n32459,
         n32460, n32461, n32462, n32463, n32464, n32465, n32466, n32467,
         n32468, n32469, n32470, n32471, n32472, n32473, n32474, n32475,
         n32476, n32477, n32478, n32479, n32480, n32481, n32482, n32483,
         n32484, n32485, n32486, n32487, n32488, n32489, n32490, n32491,
         n32492, n32493, n32494, n32495, n32496, n32497, n32498, n32499,
         n32500, n32501, n32502, n32503, n32504, n32505, n32506, n32507,
         n32508, n32509, n32510, n32511, n32512, n32513, n32514, n32515,
         n32516, n32517, n32518, n32519, n32520, n32521, n32522, n32523,
         n32524, n32525, n32526, n32527, n32528, n32529, n32530, n32531,
         n32532, n32533, n32534, n32535, n32536, n32537, n32538, n32539,
         n32540, n32541, n32542, n32543, n32544, n32545, n32546, n32547,
         n32548, n32549, n32550, n32551, n32552, n32553, n32554, n32555,
         n32556, n32557, n32558, n32559, n32560, n32561, n32562, n32563,
         n32564, n32565, n32566, n32567, n32568, n32569, n32570, n32571,
         n32572, n32573, n32574, n32575, n32576, n32577, n32578, n32579,
         n32580, n32581, n32582, n32583, n32584, n32585, n32586, n32587,
         n32588, n32589, n32590, n32591, n32592, n32593, n32594, n32595,
         n32596, n32597, n32598, n32599, n32600, n32601, n32602, n32603,
         n32604, n32605, n32606, n32607, n32608, n32609, n32610, n32611,
         n32612, n32613, n32614, n32615, n32616, n32617, n32618, n32619,
         n32620, n32621, n32622, n32623, n32624, n32625, n32626, n32627,
         n32628, n32629, n32630, n32631, n32632, n32633, n32634, n32635,
         n32636, n32637, n32638, n32639, n32640, n32641, n32642, n32643,
         n32644, n32645, n32646, n32647, n32648, n32649, n32650, n32651,
         n32652, n32653, n32654, n32655, n32656, n32657, n32658, n32659,
         n32660, n32661, n32662, n32663, n32664, n32665, n32666, n32667,
         n32668, n32669, n32670, n32671, n32672, n32673, n32674, n32675,
         n32676, n32677, n32678, n32679, n32680, n32681, n32682, n32683,
         n32684, n32685, n32686, n32687, n32688, n32689, n32690, n32691,
         n32692, n32693, n32694, n32695, n32696, n32697, n32698, n32699,
         n32700, n32701, n32702, n32703, n32704, n32705, n32706, n32707,
         n32708, n32709, n32710, n32711, n32712, n32713, n32714, n32715,
         n32716, n32717, n32718, n32719, n32720, n32721, n32722, n32723,
         n32724, n32725, n32726, n32727, n32728, n32729, n32730, n32731,
         n32732, n32733, n32734, n32735, n32736, n32737, n32738, n32739,
         n32740, n32741, n32742, n32743, n32744, n32745, n32746, n32747,
         n32748, n32749, n32750, n32751, n32752, n32753, n32754, n32755,
         n32756, n32757, n32758, n32759, n32760, n32761, n32762, n32763,
         n32764, n32765, n32766, n32767, n32768, n32769, n32770, n32771,
         n32772, n32773, n32774, n32775, n32776, n32777, n32778, n32779,
         n32780, n32781, n32782, n32783, n32784, n32785, n32786, n32787,
         n32788, n32789, n32790, n32791, n32792, n32793, n32794, n32795,
         n32796, n32797, n32798, n32799, n32800, n32801, n32802, n32803,
         n32804, n32805, n32806, n32807, n32808, n32809, n32810, n32811,
         n32812, n32813, n32814, n32815, n32816, n32817, n32818, n32819,
         n32820, n32821, n32822, n32823, n32824, n32825, n32826, n32827,
         n32828, n32829, n32830, n32831, n32832, n32833, n32834, n32835,
         n32836, n32837, n32838, n32839, n32840, n32841, n32842, n32843,
         n32844, n32845, n32846, n32847, n32848, n32849, n32850, n32851,
         n32852, n32853, n32854, n32855, n32856, n32857, n32858, n32859,
         n32860, n32861, n32862, n32863, n32864, n32865, n32866, n32867,
         n32868, n32869, n32870, n32871, n32872, n32873, n32874, n32875,
         n32876, n32877, n32878, n32879, n32880, n32881, n32882, n32883,
         n32884, n32885, n32886, n32887, n32888, n32889, n32890, n32891,
         n32892, n32893, n32894, n32895, n32896, n32897, n32898, n32899,
         n32900, n32901, n32902, n32903, n32904, n32905, n32906, n32907,
         n32908, n32909, n32910, n32911, n32912, n32913, n32914, n32915,
         n32916, n32917, n32918, n32919, n32920, n32921, n32922, n32923,
         n32924, n32925, n32926, n32927, n32928, n32929, n32930, n32931,
         n32932, n32933, n32934, n32935, n32936, n32937, n32938, n32939,
         n32940, n32941, n32942, n32943, n32944, n32945, n32946, n32947,
         n32948, n32949, n32950, n32951, n32952, n32953, n32954, n32955,
         n32956, n32957, n32958, n32959, n32960, n32961, n32962, n32963,
         n32964, n32965, n32966, n32967, n32968, n32969, n32970, n32971,
         n32972, n32973, n32974, n32975, n32976, n32977, n32978, n32979,
         n32980, n32981, n32982, n32983, n32984, n32985, n32986, n32987,
         n32988, n32989, n32990, n32991, n32992, n32993, n32994, n32995,
         n32996, n32997, n32998, n32999, n33000, n33001, n33002, n33003,
         n33004, n33005, n33006, n33007, n33008, n33009, n33010, n33011,
         n33012, n33013, n33014, n33015, n33016, n33017, n33018, n33019,
         n33020, n33021, n33022, n33023, n33024, n33025, n33026, n33027,
         n33028, n33029, n33030, n33031, n33032, n33033, n33034, n33035,
         n33036, n33037, n33038, n33039, n33040, n33041, n33042, n33043,
         n33044, n33045, n33046, n33047, n33048, n33049, n33050, n33051,
         n33052, n33053, n33054, n33055, n33056, n33057, n33058, n33059,
         n33060, n33061, n33062, n33063, n33064, n33065, n33066, n33067,
         n33068, n33069, n33070, n33071, n33072, n33073, n33074, n33075,
         n33076, n33077, n33078, n33079, n33080, n33081, n33082, n33083,
         n33084, n33085, n33086, n33087, n33088, n33089, n33090, n33091,
         n33092, n33093, n33094, n33095, n33096, n33097, n33098, n33099,
         n33100, n33101, n33102, n33103, n33104, n33105, n33106, n33107,
         n33108, n33109, n33110, n33111, n33112, n33113, n33114, n33115,
         n33116, n33117, n33118, n33119, n33120, n33121, n33122, n33123,
         n33124, n33125, n33126, n33127, n33128, n33129, n33130, n33131,
         n33132, n33133, n33134, n33135, n33136, n33137, n33138, n33139,
         n33140, n33141, n33142, n33143, n33144, n33145, n33146, n33147,
         n33148, n33149, n33150, n33151, n33152, n33153, n33154, n33155,
         n33156, n33157, n33158, n33159, n33160, n33161, n33162, n33163,
         n33164, n33165, n33166, n33167, n33168, n33169, n33170, n33171,
         n33172, n33173, n33174, n33175, n33176, n33177, n33178, n33179,
         n33180, n33181, n33182, n33183, n33184, n33185, n33186, n33187,
         n33188, n33189, n33190, n33191, n33192, n33193, n33194, n33195,
         n33196, n33197, n33198, n33199, n33200, n33201, n33202, n33203,
         n33204, n33205, n33206, n33207, n33208, n33209, n33210, n33211,
         n33212, n33213, n33214, n33215, n33216, n33217, n33218, n33219,
         n33220, n33221, n33222, n33223, n33224, n33225, n33226, n33227,
         n33228, n33229, n33230, n33231, n33232, n33233, n33234, n33235,
         n33236, n33237, n33238, n33239, n33240, n33241, n33242, n33243,
         n33244, n33245, n33246, n33247, n33248, n33249, n33250, n33251,
         n33252, n33253, n33254, n33255, n33256, n33257, n33258, n33259,
         n33260, n33261, n33262, n33263, n33264, n33265, n33266, n33267,
         n33268, n33269, n33270, n33271, n33272, n33273, n33274, n33275,
         n33276, n33277, n33278, n33279, n33280, n33281, n33282, n33283,
         n33284, n33285, n33286, n33287, n33288, n33289, n33290, n33291,
         n33292, n33293, n33294, n33295, n33296, n33297, n33298, n33299,
         n33300, n33301, n33302, n33303, n33304, n33305, n33306, n33307,
         n33308, n33309, n33310, n33311, n33312, n33313, n33314, n33315,
         n33316, n33317, n33318, n33319, n33320, n33321, n33322, n33323,
         n33324, n33325, n33326, n33327, n33328, n33329, n33330, n33331,
         n33332, n33333, n33334, n33335, n33336, n33337, n33338, n33339,
         n33340, n33341, n33342, n33343, n33344, n33345, n33346, n33347,
         n33348, n33349, n33350, n33351, n33352, n33353, n33354, n33355,
         n33356, n33357, n33358, n33359, n33360, n33361, n33362, n33363,
         n33364, n33365, n33366, n33367, n33368, n33369, n33370, n33371,
         n33372, n33373, n33374, n33375, n33376, n33377, n33378, n33379,
         n33380, n33381, n33382, n33383, n33384, n33385, n33386, n33387,
         n33388, n33389, n33390, n33391, n33392, n33393, n33394, n33395,
         n33396, n33397, n33398, n33399, n33400, n33401, n33402, n33403,
         n33404, n33405, n33406, n33407, n33408, n33409, n33410, n33411,
         n33412, n33413, n33414, n33415, n33416, n33417, n33418, n33419,
         n33420, n33421, n33422, n33423, n33424, n33425, n33426, n33427,
         n33428, n33429, n33430, n33431, n33432, n33433, n33434, n33435,
         n33436, n33437, n33438, n33439, n33440, n33441, n33442, n33443,
         n33444, n33445, n33446, n33447, n33448, n33449, n33450, n33451,
         n33452, n33453, n33454, n33455, n33456, n33457, n33458, n33459,
         n33460, n33461, n33462, n33463, n33464, n33465, n33466, n33467,
         n33468, n33469, n33470, n33471, n33472, n33473, n33474, n33475,
         n33476, n33477, n33478, n33479, n33480, n33481, n33482, n33483,
         n33484, n33485, n33486, n33487, n33488, n33489, n33490, n33491,
         n33492, n33493, n33494, n33495, n33496, n33497, n33498, n33499,
         n33500, n33501, n33502, n33503, n33504, n33505, n33506, n33507,
         n33508, n33509, n33510, n33511, n33512, n33513, n33514, n33515,
         n33516, n33517, n33518, n33519, n33520, n33521, n33522, n33523,
         n33524, n33525, n33526, n33527, n33528, n33529, n33530, n33531,
         n33532, n33533, n33534, n33535, n33536, n33537, n33538, n33539,
         n33540, n33541, n33542, n33543, n33544, n33545, n33546, n33547,
         n33548, n33549, n33550, n33551, n33552, n33553, n33554, n33555,
         n33556, n33557, n33558, n33559, n33560, n33561, n33562, n33563,
         n33564, n33565, n33566, n33567, n33568, n33569, n33570, n33571,
         n33572, n33573, n33574, n33575, n33576, n33577, n33578, n33579,
         n33580, n33581, n33582, n33583, n33584, n33585, n33586, n33587,
         n33588, n33589, n33590, n33591, n33592, n33593, n33594, n33595,
         n33596, n33597, n33598, n33599, n33600, n33601, n33602, n33603,
         n33604, n33605, n33606, n33607, n33608, n33609, n33610, n33611,
         n33612, n33613, n33614, n33615, n33616, n33617, n33618, n33619,
         n33620, n33621, n33622, n33623, n33624, n33625, n33626, n33627,
         n33628, n33629, n33630, n33631, n33632, n33633, n33634, n33635,
         n33636, n33637, n33638, n33639, n33640, n33641, n33642, n33643,
         n33644, n33645, n33646, n33647, n33648, n33649, n33650, n33651,
         n33652, n33653, n33654, n33655, n33656, n33657, n33658, n33659,
         n33660, n33661, n33662, n33663, n33664, n33665, n33666, n33667,
         n33668, n33669, n33670, n33671, n33672, n33673, n33674, n33675,
         n33676, n33677, n33678, n33679, n33680, n33681, n33682, n33683,
         n33684, n33685, n33686, n33687, n33688, n33689, n33690, n33691,
         n33692, n33693, n33694, n33695, n33696, n33697, n33698, n33699,
         n33700, n33701, n33702, n33703, n33704, n33705, n33706, n33707,
         n33708, n33709, n33710, n33711, n33712, n33713, n33714, n33715,
         n33716, n33717, n33718, n33719, n33720, n33721, n33722, n33723,
         n33724, n33725, n33726, n33727, n33728, n33729, n33730, n33731,
         n33732, n33733, n33734, n33735, n33736, n33737, n33738, n33739,
         n33740, n33741, n33742, n33743, n33744, n33745, n33746, n33747,
         n33748, n33749, n33750, n33751, n33752, n33753, n33754, n33755,
         n33756, n33757, n33758, n33759, n33760, n33761, n33762, n33763,
         n33764, n33765, n33766, n33767, n33768, n33769, n33770, n33771,
         n33772, n33773, n33774, n33775, n33776, n33777, n33778, n33779,
         n33780, n33781, n33782, n33783, n33784, n33785, n33786, n33787,
         n33788, n33789, n33790, n33791, n33792, n33793, n33794, n33795,
         n33796, n33797, n33798, n33799, n33800, n33801, n33802, n33803,
         n33804, n33805, n33806, n33807, n33808, n33809, n33810, n33811,
         n33812, n33813, n33814, n33815, n33816, n33817, n33818, n33819,
         n33820, n33821, n33822, n33823, n33824, n33825, n33826, n33827,
         n33828, n33829, n33830, n33831, n33832, n33833, n33834, n33835,
         n33836, n33837, n33838, n33839, n33840, n33841, n33842, n33843,
         n33844, n33845, n33846, n33847, n33848, n33849, n33850, n33851,
         n33852, n33853, n33854, n33855, n33856, n33857, n33858, n33859,
         n33860, n33861, n33862, n33863, n33864, n33865, n33866, n33867,
         n33868, n33869, n33870, n33871, n33872, n33873, n33874, n33875,
         n33876, n33877, n33878, n33879, n33880, n33881, n33882, n33883,
         n33884, n33885, n33886, n33887, n33888, n33889, n33890, n33891,
         n33892, n33893, n33894, n33895, n33896, n33897, n33898, n33899,
         n33900, n33901, n33902, n33903, n33904, n33905, n33906, n33907,
         n33908, n33909, n33910, n33911, n33912, n33913, n33914, n33915,
         n33916, n33917, n33918, n33919, n33920, n33921, n33922, n33923,
         n33924, n33925, n33926, n33927, n33928, n33929, n33930, n33931,
         n33932, n33933, n33934, n33935, n33936, n33937, n33938, n33939,
         n33940, n33941, n33942, n33943, n33944, n33945, n33946, n33947,
         n33948, n33949, n33950, n33951, n33952, n33953, n33954, n33955,
         n33956, n33957, n33958, n33959, n33960, n33961, n33962, n33963,
         n33964, n33965, n33966, n33967, n33968, n33969, n33970, n33971,
         n33972, n33973, n33974, n33975, n33976, n33977, n33978, n33979,
         n33980, n33981, n33982, n33983, n33984, n33985, n33986, n33987,
         n33988, n33989, n33990, n33991, n33992, n33993, n33994, n33995,
         n33996, n33997, n33998, n33999, n34000, n34001, n34002, n34003,
         n34004, n34005, n34006, n34007, n34008, n34009, n34010, n34011,
         n34012, n34013, n34014, n34015, n34016, n34017, n34018, n34019,
         n34020, n34021, n34022, n34023, n34024, n34025, n34026, n34027,
         n34028, n34029, n34030, n34031, n34032, n34033, n34034, n34035,
         n34036, n34037, n34038, n34039, n34040, n34041, n34042, n34043,
         n34044, n34045, n34046, n34047, n34048, n34049, n34050, n34051,
         n34052, n34053, n34054, n34055, n34056, n34057, n34058, n34059,
         n34060, n34061, n34062, n34063, n34064, n34065, n34066, n34067,
         n34068, n34069, n34070, n34071, n34072, n34073, n34074, n34075,
         n34076, n34077, n34078, n34079, n34080, n34081, n34082, n34083,
         n34084, n34085, n34086, n34087, n34088, n34089, n34090, n34091,
         n34092, n34093, n34094, n34095, n34096, n34097, n34098, n34099,
         n34100, n34101, n34102, n34103, n34104, n34105, n34106, n34107,
         n34108, n34109, n34110, n34111, n34112, n34113, n34114, n34115,
         n34116, n34117, n34118, n34119, n34120, n34121, n34122, n34123,
         n34124, n34125, n34126, n34127, n34128, n34129, n34130, n34131,
         n34132, n34133, n34134, n34135, n34136, n34137, n34138, n34139,
         n34140, n34141, n34142, n34143, n34144, n34145, n34146, n34147,
         n34148, n34149, n34150, n34151, n34152, n34153, n34154, n34155,
         n34156, n34157, n34158, n34159, n34160, n34161, n34162, n34163,
         n34164, n34165, n34166, n34167, n34168, n34169, n34170, n34171,
         n34172, n34173, n34174, n34175, n34176, n34177, n34178, n34179,
         n34180, n34181, n34182, n34183, n34184, n34185, n34186, n34187,
         n34188, n34189, n34190, n34191, n34192, n34193, n34194, n34195,
         n34196, n34197, n34198, n34199, n34200, n34201, n34202, n34203,
         n34204, n34205, n34206, n34207, n34208, n34209, n34210, n34211,
         n34212, n34213, n34214, n34215, n34216, n34217, n34218, n34219,
         n34220, n34221, n34222, n34223, n34224, n34225, n34226, n34227,
         n34228, n34229, n34230, n34231, n34232, n34233, n34234, n34235,
         n34236, n34237, n34238, n34239, n34240, n34241, n34242, n34243,
         n34244, n34245, n34246, n34247, n34248, n34249, n34250, n34251,
         n34252, n34253, n34254, n34255, n34256, n34257, n34258, n34259,
         n34260, n34261, n34262, n34263, n34264, n34265, n34266, n34267,
         n34268, n34269, n34270, n34271, n34272, n34273, n34274, n34275,
         n34276, n34277, n34278, n34279, n34280, n34281, n34282, n34283,
         n34284, n34285, n34286, n34287, n34288, n34289, n34290, n34291,
         n34292, n34293, n34294, n34295, n34296, n34297, n34298, n34299,
         n34300, n34301, n34302, n34303, n34304, n34305, n34306, n34307,
         n34308, n34309, n34310, n34311, n34312, n34313, n34314, n34315,
         n34316, n34317, n34318, n34319, n34320, n34321, n34322, n34323,
         n34324, n34325, n34326, n34327, n34328, n34329, n34330, n34331,
         n34332, n34333, n34334, n34335, n34336, n34337, n34338, n34339,
         n34340, n34341, n34342, n34343, n34344, n34345, n34346, n34347,
         n34348, n34349, n34350, n34351, n34352, n34353, n34354, n34355,
         n34356, n34357, n34358, n34359, n34360, n34361, n34362, n34363,
         n34364, n34365, n34366, n34367, n34368, n34369, n34370, n34371,
         n34372, n34373, n34374, n34375, n34376, n34377, n34378, n34379,
         n34380, n34381, n34382, n34383, n34384, n34385, n34386, n34387,
         n34388, n34389, n34390, n34391, n34392, n34393, n34394, n34395,
         n34396, n34397, n34398, n34399, n34400, n34401, n34402, n34403,
         n34404, n34405, n34406, n34407, n34408, n34409, n34410, n34411,
         n34412, n34413, n34414, n34415, n34416, n34417, n34418, n34419,
         n34420, n34421, n34422, n34423, n34424, n34425, n34426, n34427,
         n34428, n34429, n34430, n34431, n34432, n34433, n34434, n34435,
         n34436, n34437, n34438, n34439, n34440, n34441, n34442, n34443,
         n34444, n34445, n34446, n34447, n34448, n34449, n34450, n34451,
         n34452, n34453, n34454, n34455, n34456, n34457, n34458, n34459,
         n34460, n34461, n34462, n34463, n34464, n34465, n34466, n34467,
         n34468, n34469, n34470, n34471, n34472, n34473, n34474, n34475,
         n34476, n34477, n34478, n34479, n34480, n34481, n34482, n34483,
         n34484, n34485, n34486, n34487, n34488, n34489, n34490, n34491,
         n34492, n34493, n34494, n34495, n34496, n34497, n34498, n34499,
         n34500, n34501, n34502, n34503, n34504, n34505, n34506, n34507,
         n34508, n34509, n34510, n34511, n34512, n34513, n34514, n34515,
         n34516, n34517, n34518, n34519, n34520, n34521, n34522, n34523,
         n34524, n34525, n34526, n34527, n34528, n34529, n34530, n34531,
         n34532, n34533, n34534, n34535, n34536, n34537, n34538, n34539,
         n34540, n34541, n34542, n34543, n34544, n34545, n34546, n34547,
         n34548, n34549, n34550, n34551, n34552, n34553, n34554, n34555,
         n34556, n34557, n34558, n34559, n34560, n34561, n34562, n34563,
         n34564, n34565, n34566, n34567, n34568, n34569, n34570, n34571,
         n34572, n34573, n34574, n34575, n34576, n34577, n34578, n34579,
         n34580, n34581, n34582, n34583, n34584, n34585, n34586, n34587,
         n34588, n34589, n34590, n34591, n34592, n34593, n34594, n34595,
         n34596, n34597, n34598, n34599, n34600, n34601, n34602, n34603,
         n34604, n34605, n34606, n34607, n34608, n34609, n34610, n34611,
         n34612, n34613, n34614, n34615, n34616, n34617, n34618, n34619,
         n34620, n34621, n34622, n34623, n34624, n34625, n34626, n34627,
         n34628, n34629, n34630, n34631, n34632, n34633, n34634, n34635,
         n34636, n34637, n34638, n34639, n34640, n34641, n34642, n34643,
         n34644, n34645, n34646, n34647, n34648, n34649, n34650, n34651,
         n34652, n34653, n34654, n34655, n34656, n34657, n34658, n34659,
         n34660, n34661, n34662, n34663, n34664, n34665, n34666, n34667,
         n34668, n34669, n34670, n34671, n34672, n34673, n34674, n34675,
         n34676, n34677, n34678, n34679, n34680, n34681, n34682, n34683,
         n34684, n34685, n34686, n34687, n34688, n34689, n34690, n34691,
         n34692, n34693, n34694, n34695, n34696, n34697, n34698, n34699,
         n34700, n34701, n34702, n34703, n34704, n34705, n34706, n34707,
         n34708, n34709, n34710, n34711, n34712, n34713, n34714, n34715,
         n34716, n34717, n34718, n34719, n34720, n34721, n34722, n34723,
         n34724, n34725, n34726, n34727, n34728, n34729, n34730, n34731,
         n34732, n34733, n34734, n34735, n34736, n34737, n34738, n34739,
         n34740, n34741, n34742, n34743, n34744, n34745, n34746, n34747,
         n34748, n34749, n34750, n34751, n34752, n34753, n34754, n34755,
         n34756, n34757, n34758, n34759, n34760, n34761, n34762, n34763,
         n34764, n34765, n34766, n34767, n34768, n34769, n34770, n34771,
         n34772, n34773, n34774, n34775, n34776, n34777, n34778, n34779,
         n34780, n34781, n34782, n34783, n34784, n34785, n34786, n34787,
         n34788, n34789, n34790, n34791, n34792, n34793, n34794, n34795,
         n34796, n34797, n34798, n34799, n34800, n34801, n34802, n34803,
         n34804, n34805, n34806, n34807, n34808, n34809, n34810, n34811,
         n34812, n34813, n34814, n34815, n34816, n34817, n34818, n34819,
         n34820, n34821, n34822, n34823, n34824, n34825, n34826, n34827,
         n34828, n34829, n34830, n34831, n34832, n34833, n34834, n34835,
         n34836, n34837, n34838, n34839, n34840, n34841, n34842, n34843,
         n34844, n34845, n34846, n34847, n34848, n34849, n34850, n34851,
         n34852, n34853, n34854, n34855, n34856, n34857, n34858, n34859,
         n34860, n34861, n34862, n34863, n34864, n34865, n34866, n34867,
         n34868, n34869, n34870, n34871, n34872, n34873, n34874, n34875,
         n34876, n34877, n34878, n34879, n34880, n34881, n34882, n34883,
         n34884, n34885, n34886, n34887, n34888, n34889, n34890, n34891,
         n34892, n34893, n34894, n34895, n34896, n34897, n34898, n34899,
         n34900, n34901, n34902, n34903, n34904, n34905, n34906, n34907,
         n34908, n34909, n34910, n34911, n34912, n34913, n34914, n34915,
         n34916, n34917, n34918, n34919, n34920, n34921, n34922, n34923,
         n34924, n34925, n34926, n34927, n34928, n34929, n34930, n34931,
         n34932, n34933, n34934, n34935, n34936, n34937, n34938, n34939,
         n34940, n34941, n34942, n34943, n34944, n34945, n34946, n34947,
         n34948, n34949, n34950, n34951, n34952, n34953, n34954, n34955,
         n34956, n34957, n34958, n34959, n34960, n34961, n34962, n34963,
         n34964, n34965, n34966, n34967, n34968, n34969, n34970, n34971,
         n34972, n34973, n34974, n34975, n34976, n34977, n34978, n34979,
         n34980, n34981, n34982, n34983, n34984, n34985, n34986, n34987,
         n34988, n34989, n34990, n34991, n34992, n34993, n34994, n34995,
         n34996, n34997, n34998, n34999, n35000, n35001, n35002, n35003,
         n35004, n35005, n35006, n35007, n35008, n35009, n35010, n35011,
         n35012, n35013, n35014, n35015, n35016, n35017, n35018, n35019,
         n35020, n35021, n35022, n35023, n35024, n35025, n35026, n35027,
         n35028, n35029, n35030, n35031, n35032, n35033, n35034, n35035,
         n35036, n35037, n35038, n35039, n35040, n35041, n35042, n35043,
         n35044, n35045, n35046, n35047, n35048, n35049, n35050, n35051,
         n35052, n35053, n35054, n35055, n35056, n35057, n35058, n35059,
         n35060, n35061, n35062, n35063, n35064, n35065, n35066, n35067,
         n35068, n35069, n35070, n35071, n35072, n35073, n35074, n35075,
         n35076, n35077, n35078, n35079, n35080, n35081, n35082, n35083,
         n35084, n35085, n35086, n35087, n35088, n35089, n35090, n35091,
         n35092, n35093, n35094, n35095, n35096, n35097, n35098, n35099,
         n35100, n35101, n35102, n35103, n35104, n35105, n35106, n35107,
         n35108, n35109, n35110, n35111, n35112, n35113, n35114, n35115,
         n35116, n35117, n35118, n35119, n35120, n35121, n35122, n35123,
         n35124, n35125, n35126, n35127, n35128, n35129, n35130, n35131,
         n35132, n35133, n35134, n35135, n35136, n35137, n35138, n35139,
         n35140, n35141, n35142, n35143, n35144, n35145, n35146, n35147,
         n35148, n35149, n35150, n35151, n35152, n35153, n35154, n35155,
         n35156, n35157, n35158, n35159, n35160, n35161, n35162, n35163,
         n35164, n35165, n35166, n35167, n35168, n35169, n35170, n35171,
         n35172, n35173, n35174, n35175, n35176, n35177, n35178, n35179,
         n35180, n35181, n35182, n35183, n35184, n35185, n35186, n35187,
         n35188, n35189, n35190, n35191, n35192, n35193, n35194, n35195,
         n35196, n35197, n35198, n35199, n35200, n35201, n35202, n35203,
         n35204, n35205, n35206, n35207, n35208, n35209, n35210, n35211,
         n35212, n35213, n35214, n35215, n35216, n35217, n35218, n35219,
         n35220, n35221, n35222, n35223, n35224, n35225, n35226, n35227,
         n35228, n35229, n35230, n35231, n35232, n35233, n35234, n35235,
         n35236, n35237, n35238, n35239, n35240, n35241, n35242, n35243,
         n35244, n35245, n35246, n35247, n35248, n35249, n35250, n35251,
         n35252, n35253, n35254, n35255, n35256, n35257, n35258, n35259,
         n35260, n35261, n35262, n35263, n35264, n35265, n35266, n35267,
         n35268, n35269, n35270, n35271, n35272, n35273, n35274, n35275,
         n35276, n35277, n35278, n35279, n35280, n35281, n35282, n35283,
         n35284, n35285, n35286, n35287, n35288, n35289, n35290, n35291,
         n35292, n35293, n35294, n35295, n35296, n35297, n35298, n35299,
         n35300, n35301, n35302, n35303, n35304, n35305, n35306, n35307,
         n35308, n35309, n35310, n35311, n35312, n35313, n35314, n35315,
         n35316, n35317, n35318, n35319, n35320, n35321, n35322, n35323,
         n35324, n35325, n35326, n35327, n35328, n35329, n35330, n35331,
         n35332, n35333, n35334, n35335, n35336, n35337, n35338, n35339,
         n35340, n35341, n35342, n35343, n35344, n35345, n35346, n35347,
         n35348, n35349, n35350, n35351, n35352, n35353, n35354, n35355,
         n35356, n35357, n35358, n35359, n35360, n35361, n35362, n35363,
         n35364, n35365, n35366, n35367, n35368, n35369, n35370, n35371,
         n35372, n35373, n35374, n35375, n35376, n35377, n35378, n35379,
         n35380, n35381, n35382, n35383, n35384, n35385, n35386, n35387,
         n35388, n35389, n35390, n35391, n35392, n35393, n35394, n35395,
         n35396, n35397, n35398, n35399, n35400, n35401, n35402, n35403,
         n35404, n35405, n35406, n35407, n35408, n35409, n35410, n35411,
         n35412, n35413, n35414, n35415, n35416, n35417, n35418, n35419,
         n35420, n35421, n35422, n35423, n35424, n35425, n35426, n35427,
         n35428, n35429, n35430, n35431, n35432, n35433, n35434, n35435,
         n35436, n35437, n35438, n35439, n35440, n35441, n35442, n35443,
         n35444, n35445, n35446, n35447, n35448, n35449, n35450, n35451,
         n35452, n35453, n35454, n35455, n35456, n35457, n35458, n35459,
         n35460, n35461, n35462, n35463, n35464, n35465, n35466, n35467,
         n35468, n35469, n35470, n35471, n35472, n35473, n35474, n35475,
         n35476, n35477, n35478, n35479, n35480, n35481, n35482, n35483,
         n35484, n35485, n35486, n35487, n35488, n35489, n35490, n35491,
         n35492, n35493, n35494, n35495, n35496, n35497, n35498, n35499,
         n35500, n35501, n35502, n35503, n35504, n35505, n35506, n35507,
         n35508, n35509, n35510, n35511, n35512, n35513, n35514, n35515,
         n35516, n35517, n35518, n35519, n35520, n35521, n35522, n35523,
         n35524, n35525, n35526, n35527, n35528, n35529, n35530, n35531,
         n35532, n35533, n35534, n35535, n35536, n35537, n35538, n35539,
         n35540, n35541, n35542, n35543, n35544, n35545, n35546, n35547,
         n35548, n35549, n35550, n35551, n35552, n35553, n35554, n35555,
         n35556, n35557, n35558, n35559, n35560, n35561, n35562, n35563,
         n35564, n35565, n35566, n35567, n35568, n35569, n35570, n35571,
         n35572, n35573, n35574, n35575, n35576, n35577, n35578, n35579,
         n35580, n35581, n35582, n35583, n35584, n35585, n35586, n35587,
         n35588, n35589, n35590, n35591, n35592, n35593, n35594, n35595,
         n35596, n35597, n35598, n35599, n35600, n35601, n35602, n35603,
         n35604, n35605, n35606, n35607, n35608, n35609, n35610, n35611,
         n35612, n35613, n35614, n35615, n35616, n35617, n35618, n35619,
         n35620, n35621, n35622, n35623, n35624, n35625, n35626, n35627,
         n35628, n35629, n35630, n35631, n35632, n35633, n35634, n35635,
         n35636, n35637, n35638, n35639, n35640, n35641, n35642, n35643,
         n35644, n35645, n35646, n35647, n35648, n35649, n35650, n35651,
         n35652, n35653, n35654, n35655, n35656, n35657, n35658, n35659,
         n35660, n35661, n35662, n35663, n35664, n35665, n35666, n35667,
         n35668, n35669, n35670, n35671, n35672, n35673, n35674, n35675,
         n35676, n35677, n35678, n35679, n35680, n35681, n35682, n35683,
         n35684, n35685, n35686, n35687, n35688, n35689, n35690, n35691,
         n35692, n35693, n35694, n35695, n35696, n35697, n35698, n35699,
         n35700, n35701, n35702, n35703, n35704, n35705, n35706, n35707,
         n35708, n35709, n35710, n35711, n35712, n35713, n35714, n35715,
         n35716, n35717, n35718, n35719, n35720, n35721, n35722, n35723,
         n35724, n35725, n35726, n35727, n35728, n35729, n35730, n35731,
         n35732, n35733, n35734, n35735, n35736, n35737, n35738, n35739,
         n35740, n35741, n35742, n35743, n35744, n35745, n35746, n35747,
         n35748, n35749, n35750, n35751, n35752, n35753, n35754, n35755,
         n35756, n35757, n35758, n35759, n35760, n35761, n35762, n35763,
         n35764, n35765, n35766, n35767, n35768, n35769, n35770, n35771,
         n35772, n35773, n35774, n35775, n35776, n35777, n35778, n35779,
         n35780, n35781, n35782, n35783, n35784, n35785, n35786, n35787,
         n35788, n35789, n35790, n35791, n35792, n35793, n35794, n35795,
         n35796, n35797, n35798, n35799, n35800, n35801, n35802, n35803,
         n35804, n35805, n35806, n35807, n35808, n35809, n35810, n35811,
         n35812, n35813, n35814, n35815, n35816, n35817, n35818, n35819,
         n35820, n35821, n35822, n35823, n35824, n35825, n35826, n35827,
         n35828, n35829, n35830, n35831, n35832, n35833, n35834, n35835,
         n35836, n35837, n35838, n35839, n35840, n35841, n35842, n35843,
         n35844, n35845, n35846, n35847, n35848, n35849, n35850, n35851,
         n35852, n35853, n35854, n35855, n35856, n35857, n35858, n35859,
         n35860, n35861, n35862, n35863, n35864, n35865, n35866, n35867,
         n35868, n35869, n35870, n35871, n35872, n35873, n35874, n35875,
         n35876, n35877, n35878, n35879, n35880, n35881, n35882, n35883,
         n35884, n35885, n35886, n35887, n35888, n35889, n35890, n35891,
         n35892, n35893, n35894, n35895, n35896, n35897, n35898, n35899,
         n35900, n35901, n35902, n35903, n35904, n35905, n35906, n35907,
         n35908, n35909, n35910, n35911, n35912, n35913, n35914, n35915,
         n35916, n35917, n35918, n35919, n35920, n35921, n35922, n35923,
         n35924, n35925, n35926, n35927, n35928, n35929, n35930, n35931,
         n35932, n35933, n35934, n35935, n35936, n35937, n35938, n35939,
         n35940, n35941, n35942, n35943, n35944, n35945, n35946, n35947,
         n35948, n35949, n35950, n35951, n35952, n35953, n35954, n35955,
         n35956, n35957, n35958, n35959, n35960, n35961, n35962, n35963,
         n35964, n35965, n35966, n35967, n35968, n35969, n35970, n35971,
         n35972, n35973, n35974, n35975, n35976, n35977, n35978, n35979,
         n35980, n35981, n35982, n35983, n35984, n35985, n35986, n35987,
         n35988, n35989, n35990, n35991, n35992, n35993, n35994, n35995,
         n35996, n35997, n35998, n35999, n36000, n36001, n36002, n36003,
         n36004, n36005, n36006, n36007, n36008, n36009, n36010, n36011,
         n36012, n36013, n36014, n36015, n36016, n36017, n36018, n36019,
         n36020, n36021, n36022, n36023, n36024, n36025, n36026, n36027,
         n36028, n36029, n36030, n36031, n36032, n36033, n36034, n36035,
         n36036, n36037, n36038, n36039, n36040, n36041, n36042, n36043,
         n36044, n36045, n36046, n36047, n36048, n36049, n36050, n36051,
         n36052, n36053, n36054, n36055, n36056, n36057, n36058, n36059,
         n36060, n36061, n36062, n36063, n36064, n36065, n36066, n36067,
         n36068, n36069, n36070, n36071, n36072, n36073, n36074, n36075,
         n36076, n36077, n36078, n36079, n36080, n36081, n36082, n36083,
         n36084, n36085, n36086, n36087, n36088, n36089, n36090, n36091,
         n36092, n36093, n36094, n36095, n36096, n36097, n36098, n36099,
         n36100, n36101, n36102, n36103, n36104, n36105, n36106, n36107,
         n36108, n36109, n36110, n36111, n36112, n36113, n36114, n36115,
         n36116, n36117, n36118, n36119, n36120, n36121, n36122, n36123,
         n36124, n36125, n36126, n36127, n36128, n36129, n36130, n36131,
         n36132, n36133, n36134, n36135, n36136, n36137, n36138, n36139,
         n36140, n36141, n36142, n36143, n36144, n36145, n36146, n36147,
         n36148, n36149, n36150, n36151, n36152, n36153, n36154, n36155,
         n36156, n36157, n36158, n36159, n36160, n36161, n36162, n36163,
         n36164, n36165, n36166, n36167, n36168, n36169, n36170, n36171,
         n36172, n36173, n36174, n36175, n36176, n36177, n36178, n36179,
         n36180, n36181, n36182, n36183, n36184, n36185, n36186, n36187,
         n36188, n36189, n36190, n36191, n36192, n36193, n36194, n36195,
         n36196, n36197, n36198, n36199, n36200, n36201, n36202, n36203,
         n36204, n36205, n36206, n36207, n36208, n36209, n36210, n36211,
         n36212, n36213, n36214, n36215, n36216, n36217, n36218, n36219,
         n36220, n36221, n36222, n36223, n36224, n36225, n36226, n36227,
         n36228, n36229, n36230, n36231, n36232, n36233, n36234, n36235,
         n36236, n36237, n36238, n36239, n36240, n36241, n36242, n36243,
         n36244, n36245, n36246, n36247, n36248, n36249, n36250, n36251,
         n36252, n36253, n36254, n36255, n36256, n36257, n36258, n36259,
         n36260, n36261, n36262, n36263, n36264, n36265, n36266, n36267,
         n36268, n36269, n36270, n36271, n36272, n36273, n36274, n36275,
         n36276, n36277, n36278, n36279, n36280, n36281, n36282, n36283,
         n36284, n36285, n36286, n36287, n36288, n36289, n36290, n36291,
         n36292, n36293, n36294, n36295, n36296, n36297, n36298, n36299,
         n36300, n36301, n36302, n36303, n36304, n36305, n36306, n36307,
         n36308, n36309, n36310, n36311, n36312, n36313, n36314, n36315,
         n36316, n36317, n36318, n36319, n36320, n36321, n36322, n36323,
         n36324, n36325, n36326, n36327, n36328, n36329, n36330, n36331,
         n36332, n36333, n36334, n36335, n36336, n36337, n36338, n36339,
         n36340, n36341, n36342, n36343, n36344, n36345, n36346, n36347,
         n36348, n36349, n36350, n36351, n36352, n36353, n36354, n36355,
         n36356, n36357, n36358, n36359, n36360, n36361, n36362, n36363,
         n36364, n36365, n36366, n36367, n36368, n36369, n36370, n36371,
         n36372, n36373, n36374, n36375, n36376, n36377, n36378, n36379,
         n36380, n36381, n36382, n36383, n36384, n36385, n36386, n36387,
         n36388, n36389, n36390, n36391, n36392, n36393, n36394, n36395,
         n36396, n36397, n36398, n36399, n36400, n36401, n36402, n36403,
         n36404, n36405, n36406, n36407, n36408, n36409, n36410, n36411,
         n36412, n36413, n36414, n36415, n36416, n36417, n36418, n36419,
         n36420, n36421, n36422, n36423, n36424, n36425, n36426, n36427,
         n36428, n36429, n36430, n36431, n36432, n36433, n36434, n36435,
         n36436, n36437, n36438, n36439, n36440, n36441, n36442, n36443,
         n36444, n36445, n36446, n36447, n36448, n36449, n36450, n36451,
         n36452, n36453, n36454, n36455, n36456, n36457, n36458, n36459,
         n36460, n36461, n36462, n36463, n36464, n36465, n36466, n36467,
         n36468, n36469, n36470, n36471, n36472, n36473, n36474, n36475,
         n36476, n36477, n36478, n36479, n36480, n36481, n36482, n36483,
         n36484, n36485, n36486, n36487, n36488, n36489, n36490, n36491,
         n36492, n36493, n36494, n36495, n36496, n36497, n36498, n36499,
         n36500, n36501, n36502, n36503, n36504, n36505, n36506, n36507,
         n36508, n36509, n36510, n36511, n36512, n36513, n36514, n36515,
         n36516, n36517, n36518, n36519, n36520, n36521, n36522, n36523,
         n36524, n36525, n36526, n36527, n36528, n36529, n36530, n36531,
         n36532, n36533, n36534, n36535, n36536, n36537, n36538, n36539,
         n36540, n36541, n36542, n36543, n36544, n36545, n36546, n36547,
         n36548, n36549, n36550, n36551, n36552, n36553, n36554, n36555,
         n36556, n36557, n36558, n36559, n36560, n36561, n36562, n36563,
         n36564, n36565, n36566, n36567, n36568, n36569, n36570, n36571,
         n36572, n36573, n36574, n36575, n36576, n36577, n36578, n36579,
         n36580, n36581, n36582, n36583, n36584, n36585, n36586, n36587,
         n36588, n36589, n36590, n36591, n36592, n36593, n36594, n36595,
         n36596, n36597, n36598, n36599, n36600, n36601, n36602, n36603,
         n36604, n36605, n36606, n36607, n36608, n36609, n36610, n36611,
         n36612, n36613, n36614, n36615, n36616, n36617, n36618, n36619,
         n36620, n36621, n36622, n36623, n36624, n36625, n36626, n36627,
         n36628, n36629, n36630, n36631, n36632, n36633, n36634, n36635,
         n36636, n36637, n36638, n36639, n36640, n36641, n36642, n36643,
         n36644, n36645, n36646, n36647, n36648, n36649, n36650, n36651,
         n36652, n36653, n36654, n36655, n36656, n36657, n36658, n36659,
         n36660, n36661, n36662, n36663, n36664, n36665, n36666, n36667,
         n36668, n36669, n36670, n36671, n36672, n36673, n36674, n36675,
         n36676, n36677, n36678, n36679, n36680, n36681, n36682, n36683,
         n36684, n36685, n36686, n36687, n36688, n36689, n36690, n36691,
         n36692, n36693, n36694, n36695, n36696, n36697, n36698, n36699,
         n36700, n36701, n36702, n36703, n36704, n36705, n36706, n36707,
         n36708, n36709, n36710, n36711, n36712, n36713, n36714, n36715,
         n36716, n36717, n36718, n36719, n36720, n36721, n36722, n36723,
         n36724, n36725, n36726, n36727, n36728, n36729, n36730, n36731,
         n36732, n36733, n36734, n36735, n36736, n36737, n36738, n36739,
         n36740, n36741, n36742, n36743, n36744, n36745, n36746, n36747,
         n36748, n36749, n36750, n36751, n36752, n36753, n36754, n36755,
         n36756, n36757, n36758, n36759, n36760, n36761, n36762, n36763,
         n36764, n36765, n36766, n36767, n36768, n36769, n36770, n36771,
         n36772, n36773, n36774, n36775, n36776, n36777, n36778, n36779,
         n36780, n36781, n36782, n36783, n36784, n36785, n36786, n36787,
         n36788, n36789, n36790, n36791, n36792, n36793, n36794, n36795,
         n36796, n36797, n36798, n36799, n36800, n36801, n36802, n36803,
         n36804, n36805, n36806, n36807, n36808, n36809, n36810, n36811,
         n36812, n36813, n36814, n36815, n36816, n36817, n36818, n36819,
         n36820, n36821, n36822, n36823, n36824, n36825, n36826, n36827,
         n36828, n36829, n36830, n36831, n36832, n36833, n36834, n36835,
         n36836, n36837, n36838, n36839, n36840, n36841, n36842, n36843,
         n36844, n36845, n36846, n36847, n36848, n36849, n36850, n36851,
         n36852, n36853, n36854, n36855, n36856, n36857, n36858, n36859,
         n36860, n36861, n36862, n36863, n36864, n36865, n36866, n36867,
         n36868, n36869, n36870, n36871, n36872, n36873, n36874, n36875,
         n36876, n36877, n36878, n36879, n36880, n36881, n36882, n36883,
         n36884, n36885, n36886, n36887, n36888, n36889, n36890, n36891,
         n36892, n36893, n36894, n36895, n36896, n36897, n36898, n36899,
         n36900, n36901, n36902, n36903, n36904, n36905, n36906, n36907,
         n36908, n36909, n36910, n36911, n36912, n36913, n36914, n36915,
         n36916, n36917, n36918, n36919, n36920, n36921, n36922, n36923,
         n36924, n36925, n36926, n36927, n36928, n36929, n36930, n36931,
         n36932, n36933, n36934, n36935, n36936, n36937, n36938, n36939,
         n36940, n36941, n36942, n36943, n36944, n36945, n36946, n36947,
         n36948, n36949, n36950, n36951, n36952, n36953, n36954, n36955,
         n36956, n36957, n36958, n36959, n36960, n36961, n36962, n36963,
         n36964, n36965, n36966, n36967, n36968, n36969, n36970, n36971,
         n36972, n36973, n36974, n36975, n36976, n36977, n36978, n36979,
         n36980, n36981, n36982, n36983, n36984, n36985, n36986, n36987,
         n36988, n36989, n36990, n36991, n36992, n36993, n36994, n36995,
         n36996, n36997, n36998, n36999, n37000, n37001, n37002, n37003,
         n37004, n37005, n37006, n37007, n37008, n37009, n37010, n37011,
         n37012, n37013, n37014, n37015, n37016, n37017, n37018, n37019,
         n37020, n37021, n37022, n37023, n37024, n37025, n37026, n37027,
         n37028, n37029, n37030, n37031, n37032, n37033, n37034, n37035,
         n37036, n37037, n37038, n37039, n37040, n37041, n37042, n37043,
         n37044, n37045, n37046, n37047, n37048, n37049, n37050, n37051,
         n37052, n37053, n37054, n37055, n37056, n37057, n37058, n37059,
         n37060, n37061, n37062, n37063, n37064, n37065, n37066, n37067,
         n37068, n37069, n37070, n37071, n37072, n37073, n37074, n37075,
         n37076, n37077, n37078, n37079, n37080, n37081, n37082, n37083,
         n37084, n37085, n37086, n37087, n37088, n37089, n37090, n37091,
         n37092, n37093, n37094, n37095, n37096, n37097, n37098, n37099,
         n37100, n37101, n37102, n37103, n37104, n37105, n37106, n37107,
         n37108, n37109, n37110, n37111, n37112, n37113, n37114, n37115,
         n37116, n37117, n37118, n37119, n37120, n37121, n37122, n37123,
         n37124, n37125, n37126, n37127, n37128, n37129, n37130, n37131,
         n37132, n37133, n37134, n37135, n37136, n37137, n37138, n37139,
         n37140, n37141, n37142, n37143, n37144, n37145, n37146, n37147,
         n37148, n37149, n37150, n37151, n37152, n37153, n37154, n37155,
         n37156, n37157, n37158, n37159, n37160, n37161, n37162, n37163,
         n37164, n37165, n37166, n37167, n37168, n37169, n37170, n37171,
         n37172, n37173, n37174, n37175, n37176, n37177, n37178, n37179,
         n37180, n37181, n37182, n37183, n37184, n37185, n37186, n37187,
         n37188, n37189, n37190, n37191, n37192, n37193, n37194, n37195,
         n37196, n37197, n37198, n37199, n37200, n37201, n37202, n37203,
         n37204, n37205, n37206, n37207, n37208, n37209, n37210, n37211,
         n37212, n37213, n37214, n37215, n37216, n37217, n37218, n37219,
         n37220, n37221, n37222, n37223, n37224, n37225, n37226, n37227,
         n37228, n37229, n37230, n37231, n37232, n37233, n37234, n37235,
         n37236, n37237, n37238, n37239, n37240, n37241, n37242, n37243,
         n37244, n37245, n37246, n37247, n37248, n37249, n37250, n37251,
         n37252, n37253, n37254, n37255, n37256, n37257, n37258, n37259,
         n37260, n37261, n37262, n37263, n37264, n37265, n37266, n37267,
         n37268, n37269, n37270, n37271, n37272, n37273, n37274, n37275,
         n37276, n37277, n37278, n37279, n37280, n37281, n37282, n37283,
         n37284, n37285, n37286, n37287, n37288, n37289, n37290, n37291,
         n37292, n37293, n37294, n37295, n37296, n37297, n37298, n37299,
         n37300, n37301, n37302, n37303, n37304, n37305, n37306, n37307,
         n37308, n37309, n37310, n37311, n37312, n37313, n37314, n37315,
         n37316, n37317, n37318, n37319, n37320, n37321, n37322, n37323,
         n37324, n37325, n37326, n37327, n37328, n37329, n37330, n37331,
         n37332, n37333, n37334, n37335, n37336, n37337, n37338, n37339,
         n37340, n37341, n37342, n37343, n37344, n37345, n37346, n37347,
         n37348, n37349, n37350, n37351, n37352, n37353, n37354, n37355,
         n37356, n37357, n37358, n37359, n37360, n37361, n37362, n37363,
         n37364, n37365, n37366, n37367, n37368, n37369, n37370, n37371,
         n37372, n37373, n37374, n37375, n37376, n37377, n37378, n37379,
         n37380, n37381, n37382, n37383, n37384, n37385, n37386, n37387,
         n37388, n37389, n37390, n37391, n37392, n37393, n37394, n37395,
         n37396, n37397, n37398, n37399, n37400, n37401, n37402, n37403,
         n37404, n37405, n37406, n37407, n37408, n37409, n37410, n37411,
         n37412, n37413, n37414, n37415, n37416, n37417, n37418, n37419,
         n37420, n37421, n37422, n37423, n37424, n37425, n37426, n37427,
         n37428, n37429, n37430, n37431, n37432, n37433, n37434, n37435,
         n37436, n37437, n37438, n37439, n37440, n37441, n37442, n37443,
         n37444, n37445, n37446, n37447, n37448, n37449, n37450, n37451,
         n37452, n37453, n37454, n37455, n37456, n37457, n37458, n37459,
         n37460, n37461, n37462, n37463, n37464, n37465, n37466, n37467,
         n37468, n37469, n37470, n37471, n37472, n37473, n37474, n37475,
         n37476, n37477, n37478, n37479, n37480, n37481, n37482, n37483,
         n37484, n37485, n37486, n37487, n37488, n37489, n37490, n37491,
         n37492, n37493, n37494, n37495, n37496, n37497, n37498, n37499,
         n37500, n37501, n37502, n37503, n37504, n37505, n37506, n37507,
         n37508, n37509, n37510, n37511, n37512, n37513, n37514, n37515,
         n37516, n37517, n37518, n37519, n37520, n37521, n37522, n37523,
         n37524, n37525, n37526, n37527, n37528, n37529, n37530, n37531,
         n37532, n37533, n37534, n37535, n37536, n37537, n37538, n37539,
         n37540, n37541, n37542, n37543, n37544, n37545, n37546, n37547,
         n37548, n37549, n37550, n37551, n37552, n37553, n37554, n37555,
         n37556, n37557, n37558, n37559, n37560, n37561, n37562, n37563,
         n37564, n37565, n37566, n37567, n37568, n37569, n37570, n37571,
         n37572, n37573, n37574, n37575, n37576, n37577, n37578, n37579,
         n37580, n37581, n37582, n37583, n37584, n37585, n37586, n37587,
         n37588, n37589, n37590, n37591, n37592, n37593, n37594, n37595,
         n37596, n37597, n37598, n37599, n37600, n37601, n37602, n37603,
         n37604, n37605, n37606, n37607, n37608, n37609, n37610, n37611,
         n37612, n37613, n37614, n37615, n37616, n37617, n37618, n37619,
         n37620, n37621, n37622, n37623, n37624, n37625, n37626, n37627,
         n37628, n37629, n37630, n37631, n37632, n37633, n37634, n37635,
         n37636, n37637, n37638, n37639, n37640, n37641, n37642, n37643,
         n37644, n37645, n37646, n37647, n37648, n37649, n37650, n37651,
         n37652, n37653, n37654, n37655, n37656, n37657, n37658, n37659,
         n37660, n37661, n37662, n37663, n37664, n37665, n37666, n37667,
         n37668, n37669, n37670, n37671, n37672, n37673, n37674, n37675,
         n37676, n37677, n37678, n37679, n37680, n37681, n37682, n37683,
         n37684, n37685, n37686, n37687, n37688, n37689, n37690, n37691,
         n37692, n37693, n37694, n37695, n37696, n37697, n37698, n37699,
         n37700, n37701, n37702, n37703, n37704, n37705, n37706, n37707,
         n37708, n37709, n37710, n37711, n37712, n37713, n37714, n37715,
         n37716, n37717, n37718, n37719, n37720, n37721, n37722, n37723,
         n37724, n37725, n37726, n37727, n37728, n37729, n37730, n37731,
         n37732, n37733, n37734, n37735, n37736, n37737, n37738, n37739,
         n37740, n37741, n37742, n37743, n37744, n37745, n37746, n37747,
         n37748, n37749, n37750, n37751, n37752, n37753, n37754, n37755,
         n37756, n37757, n37758, n37759, n37760, n37761, n37762, n37763,
         n37764, n37765, n37766, n37767, n37768, n37769, n37770, n37771,
         n37772, n37773, n37774, n37775, n37776, n37777, n37778, n37779,
         n37780, n37781, n37782, n37783, n37784, n37785, n37786, n37787,
         n37788, n37789, n37790, n37791, n37792, n37793, n37794, n37795,
         n37796, n37797, n37798, n37799, n37800, n37801, n37802, n37803,
         n37804, n37805, n37806, n37807, n37808, n37809, n37810, n37811,
         n37812, n37813, n37814, n37815, n37816, n37817, n37818, n37819,
         n37820, n37821, n37822, n37823, n37824, n37825, n37826, n37827,
         n37828, n37829, n37830, n37831, n37832, n37833, n37834, n37835,
         n37836, n37837, n37838, n37839, n37840, n37841, n37842, n37843,
         n37844, n37845, n37846, n37847, n37848, n37849, n37850, n37851,
         n37852, n37853, n37854, n37855, n37856, n37857, n37858, n37859,
         n37860, n37861, n37862, n37863, n37864, n37865, n37866, n37867,
         n37868, n37869, n37870, n37871, n37872, n37873, n37874, n37875,
         n37876, n37877, n37878, n37879, n37880, n37881, n37882, n37883,
         n37884, n37885, n37886, n37887, n37888, n37889, n37890, n37891,
         n37892, n37893, n37894, n37895, n37896, n37897, n37898, n37899,
         n37900, n37901, n37902, n37903, n37904, n37905, n37906, n37907,
         n37908, n37909, n37910, n37911, n37912, n37913, n37914, n37915,
         n37916, n37917, n37918, n37919, n37920, n37921, n37922, n37923,
         n37924, n37925, n37926, n37927, n37928, n37929, n37930, n37931,
         n37932, n37933, n37934, n37935, n37936, n37937, n37938, n37939,
         n37940, n37941, n37942, n37943, n37944, n37945, n37946, n37947,
         n37948, n37949, n37950, n37951, n37952, n37953, n37954, n37955,
         n37956, n37957, n37958, n37959, n37960, n37961, n37962, n37963,
         n37964, n37965, n37966, n37967, n37968, n37969, n37970, n37971,
         n37972, n37973, n37974, n37975, n37976, n37977, n37978, n37979,
         n37980, n37981, n37982, n37983, n37984, n37985, n37986, n37987,
         n37988, n37989, n37990, n37991, n37992, n37993, n37994, n37995,
         n37996, n37997, n37998, n37999, n38000, n38001, n38002, n38003,
         n38004, n38005, n38006, n38007, n38008, n38009, n38010, n38011,
         n38012, n38013, n38014, n38015, n38016, n38017, n38018, n38019,
         n38020, n38021, n38022, n38023, n38024, n38025, n38026, n38027,
         n38028, n38029, n38030, n38031, n38032, n38033, n38034, n38035,
         n38036, n38037, n38038, n38039, n38040, n38041, n38042, n38043,
         n38044, n38045, n38046, n38047, n38048, n38049, n38050, n38051,
         n38052, n38053, n38054, n38055, n38056, n38057, n38058, n38059,
         n38060, n38061, n38062, n38063, n38064, n38065, n38066, n38067,
         n38068, n38069, n38070, n38071, n38072, n38073, n38074, n38075,
         n38076, n38077, n38078, n38079, n38080, n38081, n38082, n38083,
         n38084, n38085, n38086, n38087, n38088, n38089, n38090, n38091,
         n38092, n38093, n38094, n38095, n38096, n38097, n38098, n38099,
         n38100, n38101, n38102, n38103, n38104, n38105, n38106, n38107,
         n38108, n38109, n38110, n38111, n38112, n38113, n38114, n38115,
         n38116, n38117, n38118, n38119, n38120, n38121, n38122, n38123,
         n38124, n38125, n38126, n38127, n38128, n38129, n38130, n38131,
         n38132, n38133, n38134, n38135, n38136, n38137, n38138, n38139,
         n38140, n38141, n38142, n38143, n38144, n38145, n38146, n38147,
         n38148, n38149, n38150, n38151, n38152, n38153, n38154, n38155,
         n38156, n38157, n38158, n38159, n38160, n38161, n38162, n38163,
         n38164, n38165, n38166, n38167, n38168, n38169, n38170, n38171,
         n38172, n38173, n38174, n38175, n38176, n38177, n38178, n38179,
         n38180, n38181, n38182, n38183, n38184, n38185, n38186, n38187,
         n38188, n38189, n38190, n38191, n38192, n38193, n38194, n38195,
         n38196, n38197, n38198, n38199, n38200, n38201, n38202, n38203,
         n38204, n38205, n38206, n38207, n38208, n38209, n38210, n38211,
         n38212, n38213, n38214, n38215, n38216, n38217, n38218, n38219,
         n38220, n38221, n38222, n38223, n38224, n38225, n38226, n38227,
         n38228, n38229, n38230, n38231, n38232, n38233, n38234, n38235,
         n38236, n38237, n38238, n38239, n38240, n38241, n38242, n38243,
         n38244, n38245, n38246, n38247, n38248, n38249, n38250, n38251,
         n38252, n38253, n38254, n38255, n38256, n38257, n38258, n38259,
         n38260, n38261, n38262, n38263, n38264, n38265, n38266, n38267,
         n38268, n38269, n38270, n38271, n38272, n38273, n38274, n38275,
         n38276, n38277, n38278, n38279, n38280, n38281, n38282, n38283,
         n38284, n38285, n38286, n38287, n38288, n38289, n38290, n38291,
         n38292, n38293, n38294, n38295, n38296, n38297, n38298, n38299,
         n38300, n38301, n38302, n38303, n38304, n38305, n38306, n38307,
         n38308, n38309, n38310, n38311, n38312, n38313, n38314, n38315,
         n38316, n38317, n38318, n38319, n38320, n38321, n38322, n38323,
         n38324, n38325, n38326, n38327, n38328, n38329, n38330, n38331,
         n38332, n38333, n38334, n38335, n38336, n38337, n38338, n38339,
         n38340, n38341, n38342, n38343, n38344, n38345, n38346, n38347,
         n38348, n38349, n38350, n38351, n38352, n38353, n38354, n38355,
         n38356, n38357, n38358, n38359, n38360, n38361, n38362, n38363,
         n38364, n38365, n38366, n38367, n38368, n38369, n38370, n38371,
         n38372, n38373, n38374, n38375, n38376, n38377, n38378, n38379,
         n38380, n38381, n38382, n38383, n38384, n38385, n38386, n38387,
         n38388, n38389, n38390, n38391, n38392, n38393, n38394, n38395,
         n38396, n38397, n38398, n38399, n38400, n38401, n38402, n38403,
         n38404, n38405, n38406, n38407, n38408, n38409, n38410, n38411,
         n38412, n38413, n38414, n38415, n38416, n38417, n38418, n38419,
         n38420, n38421, n38422, n38423, n38424, n38425, n38426, n38427,
         n38428, n38429, n38430, n38431, n38432, n38433, n38434, n38435,
         n38436, n38437, n38438, n38439, n38440, n38441, n38442, n38443,
         n38444, n38445, n38446, n38447, n38448, n38449, n38450, n38451,
         n38452, n38453, n38454, n38455, n38456, n38457, n38458, n38459,
         n38460, n38461, n38462, n38463, n38464, n38465, n38466, n38467,
         n38468, n38469, n38470, n38471, n38472, n38473, n38474, n38475,
         n38476, n38477, n38478, n38479, n38480, n38481, n38482, n38483,
         n38484, n38485, n38486, n38487, n38488, n38489, n38490, n38491,
         n38492, n38493, n38494, n38495, n38496, n38497, n38498, n38499,
         n38500, n38501, n38502, n38503, n38504, n38505, n38506, n38507,
         n38508, n38509, n38510, n38511, n38512, n38513, n38514, n38515,
         n38516, n38517, n38518, n38519, n38520, n38521, n38522, n38523,
         n38524, n38525, n38526, n38527, n38528, n38529, n38530, n38531,
         n38532, n38533, n38534, n38535, n38536, n38537, n38538, n38539,
         n38540, n38541, n38542, n38543, n38544, n38545, n38546, n38547,
         n38548, n38549, n38550, n38551, n38552, n38553, n38554, n38555,
         n38556, n38557, n38558, n38559, n38560, n38561, n38562, n38563,
         n38564, n38565, n38566, n38567, n38568, n38569, n38570, n38571,
         n38572, n38573, n38574, n38575, n38576, n38577, n38578, n38579,
         n38580, n38581, n38582, n38583, n38584, n38585, n38586, n38587,
         n38588, n38589, n38590, n38591, n38592, n38593, n38594, n38595,
         n38596, n38597, n38598, n38599, n38600, n38601, n38602, n38603,
         n38604, n38605, n38606, n38607, n38608, n38609, n38610, n38611,
         n38612, n38613, n38614, n38615, n38616, n38617, n38618, n38619,
         n38620, n38621, n38622, n38623, n38624, n38625, n38626, n38627,
         n38628, n38629, n38630, n38631, n38632, n38633, n38634, n38635,
         n38636, n38637, n38638, n38639, n38640, n38641, n38642, n38643,
         n38644, n38645, n38646, n38647, n38648, n38649, n38650, n38651,
         n38652, n38653, n38654, n38655, n38656, n38657, n38658, n38659,
         n38660, n38661, n38662, n38663, n38664, n38665, n38666, n38667,
         n38668, n38669, n38670, n38671, n38672, n38673, n38674, n38675,
         n38676, n38677, n38678, n38679, n38680, n38681, n38682, n38683,
         n38684, n38685, n38686, n38687, n38688, n38689, n38690, n38691,
         n38692, n38693, n38694, n38695, n38696, n38697, n38698, n38699,
         n38700, n38701, n38702, n38703, n38704, n38705, n38706, n38707,
         n38708, n38709, n38710, n38711, n38712, n38713, n38714, n38715,
         n38716, n38717, n38718, n38719, n38720, n38721, n38722, n38723,
         n38724, n38725, n38726, n38727, n38728, n38729, n38730, n38731,
         n38732, n38733, n38734, n38735, n38736, n38737, n38738, n38739,
         n38740, n38741, n38742, n38743, n38744, n38745, n38746, n38747,
         n38748, n38749, n38750, n38751, n38752, n38753, n38754, n38755,
         n38756, n38757, n38758, n38759, n38760, n38761, n38762, n38763,
         n38764, n38765, n38766, n38767, n38768, n38769, n38770, n38771,
         n38772, n38773, n38774, n38775, n38776, n38777, n38778, n38779,
         n38780, n38781, n38782, n38783, n38784, n38785, n38786, n38787,
         n38788, n38789, n38790, n38791, n38792, n38793, n38794, n38795,
         n38796, n38797, n38798, n38799, n38800, n38801, n38802, n38803,
         n38804, n38805, n38806, n38807, n38808, n38809, n38810, n38811,
         n38812, n38813, n38814, n38815, n38816, n38817, n38818, n38819,
         n38820, n38821, n38822, n38823, n38824, n38825, n38826, n38827,
         n38828, n38829, n38830, n38831, n38832, n38833, n38834, n38835,
         n38836, n38837, n38838, n38839, n38840, n38841, n38842, n38843,
         n38844, n38845, n38846, n38847, n38848, n38849, n38850, n38851,
         n38852, n38853, n38854, n38855, n38856, n38857, n38858, n38859,
         n38860, n38861, n38862, n38863, n38864, n38865, n38866, n38867,
         n38868, n38869, n38870, n38871, n38872, n38873, n38874, n38875,
         n38876, n38877, n38878, n38879, n38880, n38881, n38882, n38883,
         n38884, n38885, n38886, n38887, n38888, n38889, n38890, n38891,
         n38892, n38893, n38894, n38895, n38896, n38897, n38898, n38899,
         n38900, n38901, n38902, n38903, n38904, n38905, n38906, n38907,
         n38908, n38909, n38910, n38911, n38912, n38913, n38914, n38915,
         n38916, n38917, n38918, n38919, n38920, n38921, n38922, n38923,
         n38924, n38925, n38926, n38927, n38928, n38929, n38930, n38931,
         n38932, n38933, n38934, n38935, n38936, n38937, n38938, n38939,
         n38940, n38941, n38942, n38943, n38944, n38945, n38946, n38947,
         n38948, n38949, n38950, n38951, n38952, n38953, n38954, n38955,
         n38956, n38957, n38958, n38959, n38960, n38961, n38962, n38963,
         n38964, n38965, n38966, n38967, n38968, n38969, n38970, n38971,
         n38972, n38973, n38974, n38975, n38976, n38977, n38978, n38979,
         n38980, n38981, n38982, n38983, n38984, n38985, n38986, n38987,
         n38988, n38989, n38990, n38991, n38992, n38993, n38994, n38995,
         n38996, n38997, n38998, n38999, n39000, n39001, n39002, n39003,
         n39004, n39005, n39006, n39007, n39008, n39009, n39010, n39011,
         n39012, n39013, n39014, n39015, n39016, n39017, n39018, n39019,
         n39020, n39021, n39022, n39023, n39024, n39025, n39026, n39027,
         n39028, n39029, n39030, n39031, n39032, n39033, n39034, n39035,
         n39036, n39037, n39038, n39039, n39040, n39041, n39042, n39043,
         n39044, n39045, n39046, n39047, n39048, n39049, n39050, n39051,
         n39052, n39053, n39054, n39055, n39056, n39057, n39058, n39059,
         n39060, n39061, n39062, n39063, n39064, n39065, n39066, n39067,
         n39068, n39069, n39070, n39071, n39072, n39073, n39074, n39075,
         n39076, n39077, n39078, n39079, n39080, n39081, n39082, n39083,
         n39084, n39085, n39086, n39087, n39088, n39089, n39090, n39091,
         n39092, n39093, n39094, n39095, n39096, n39097, n39098, n39099,
         n39100, n39101, n39102, n39103, n39104, n39105, n39106, n39107,
         n39108, n39109, n39110, n39111, n39112, n39113, n39114, n39115,
         n39116, n39117, n39118, n39119, n39120, n39121, n39122, n39123,
         n39124, n39125, n39126, n39127, n39128, n39129, n39130, n39131,
         n39132, n39133, n39134, n39135, n39136, n39137, n39138, n39139,
         n39140, n39141, n39142, n39143, n39144, n39145, n39146, n39147,
         n39148, n39149, n39150, n39151, n39152, n39153, n39154, n39155,
         n39156, n39157, n39158, n39159, n39160, n39161, n39162, n39163,
         n39164, n39165, n39166, n39167, n39168, n39169, n39170, n39171,
         n39172, n39173, n39174, n39175, n39176, n39177, n39178, n39179,
         n39180, n39181, n39182, n39183, n39184, n39185, n39186, n39187,
         n39188, n39189, n39190, n39191, n39192, n39193, n39194, n39195,
         n39196, n39197, n39198, n39199, n39200, n39201, n39202, n39203,
         n39204, n39205, n39206, n39207, n39208, n39209, n39210, n39211,
         n39212, n39213, n39214, n39215, n39216, n39217, n39218, n39219,
         n39220, n39221, n39222, n39223, n39224, n39225, n39226, n39227,
         n39228, n39229, n39230, n39231, n39232, n39233, n39234, n39235,
         n39236, n39237, n39238, n39239, n39240, n39241, n39242, n39243,
         n39244, n39245, n39246, n39247, n39248, n39249, n39250, n39251,
         n39252, n39253, n39254, n39255, n39256, n39257, n39258, n39259,
         n39260, n39261, n39262, n39263, n39264, n39265, n39266, n39267,
         n39268, n39269, n39270, n39271, n39272, n39273, n39274, n39275,
         n39276, n39277, n39278, n39279, n39280, n39281, n39282, n39283,
         n39284, n39285, n39286, n39287, n39288, n39289, n39290, n39291,
         n39292, n39293, n39294, n39295, n39296, n39297, n39298, n39299,
         n39300, n39301, n39302, n39303, n39304, n39305, n39306, n39307,
         n39308, n39309, n39310, n39311, n39312, n39313, n39314, n39315,
         n39316, n39317, n39318, n39319, n39320, n39321, n39322, n39323,
         n39324, n39325, n39326, n39327, n39328, n39329, n39330, n39331,
         n39332, n39333, n39334, n39335, n39336, n39337, n39338, n39339,
         n39340, n39341, n39342, n39343, n39344, n39345, n39346, n39347,
         n39348, n39349, n39350, n39351, n39352, n39353, n39354, n39355,
         n39356, n39357, n39358, n39359, n39360, n39361, n39362, n39363,
         n39364, n39365, n39366, n39367, n39368, n39369, n39370, n39371,
         n39372, n39373, n39374, n39375, n39376, n39377, n39378, n39379,
         n39380, n39381, n39382, n39383, n39384, n39385, n39386, n39387,
         n39388, n39389, n39390, n39391, n39392, n39393, n39394, n39395,
         n39396, n39397, n39398, n39399, n39400, n39401, n39402, n39403,
         n39404, n39405, n39406, n39407, n39408, n39409, n39410, n39411,
         n39412, n39413, n39414, n39415, n39416, n39417, n39418, n39419,
         n39420, n39421, n39422, n39423, n39424, n39425, n39426, n39427,
         n39428, n39429, n39430, n39431, n39432, n39433, n39434, n39435,
         n39436, n39437, n39438, n39439, n39440, n39441, n39442, n39443,
         n39444, n39445, n39446, n39447, n39448, n39449, n39450, n39451,
         n39452, n39453, n39454, n39455, n39456, n39457, n39458, n39459,
         n39460, n39461, n39462, n39463, n39464, n39465, n39466, n39467,
         n39468, n39469, n39470, n39471, n39472, n39473, n39474, n39475,
         n39476, n39477, n39478, n39479, n39480, n39481, n39482, n39483,
         n39484, n39485, n39486, n39487, n39488, n39489, n39490, n39491,
         n39492, n39493, n39494, n39495, n39496, n39497, n39498, n39499,
         n39500, n39501, n39502, n39503, n39504, n39505, n39506, n39507,
         n39508, n39509, n39510, n39511, n39512, n39513, n39514, n39515,
         n39516, n39517, n39518, n39519, n39520, n39521, n39522, n39523,
         n39524, n39525, n39526, n39527, n39528, n39529, n39530, n39531,
         n39532, n39533, n39534, n39535, n39536, n39537, n39538, n39539,
         n39540, n39541, n39542, n39543, n39544, n39545, n39546, n39547,
         n39548, n39549, n39550, n39551, n39552, n39553, n39554, n39555,
         n39556, n39557, n39558, n39559, n39560, n39561, n39562, n39563,
         n39564, n39565, n39566, n39567, n39568, n39569, n39570, n39571,
         n39572, n39573, n39574, n39575, n39576, n39577, n39578, n39579,
         n39580, n39581, n39582, n39583, n39584, n39585, n39586, n39587,
         n39588, n39589, n39590, n39591, n39592, n39593, n39594, n39595,
         n39596, n39597, n39598, n39599, n39600, n39601, n39602, n39603,
         n39604, n39605, n39606, n39607, n39608, n39609, n39610, n39611,
         n39612, n39613, n39614, n39615, n39616, n39617, n39618, n39619,
         n39620, n39621, n39622, n39623, n39624, n39625, n39626, n39627,
         n39628, n39629, n39630, n39631, n39632, n39633, n39634, n39635,
         n39636, n39637, n39638, n39639, n39640, n39641, n39642, n39643,
         n39644, n39645, n39646, n39647, n39648, n39649, n39650, n39651,
         n39652, n39653, n39654, n39655, n39656, n39657, n39658, n39659,
         n39660, n39661, n39662, n39663, n39664, n39665, n39666, n39667,
         n39668, n39669, n39670, n39671, n39672, n39673, n39674, n39675,
         n39676, n39677, n39678, n39679, n39680, n39681, n39682, n39683,
         n39684, n39685, n39686, n39687, n39688, n39689, n39690, n39691,
         n39692, n39693, n39694, n39695, n39696, n39697, n39698, n39699,
         n39700, n39701, n39702, n39703, n39704, n39705, n39706, n39707,
         n39708, n39709, n39710, n39711, n39712, n39713, n39714, n39715,
         n39716, n39717, n39718, n39719, n39720, n39721, n39722, n39723,
         n39724, n39725, n39726, n39727, n39728, n39729, n39730, n39731,
         n39732, n39733, n39734, n39735, n39736, n39737, n39738, n39739,
         n39740, n39741, n39742, n39743, n39744, n39745, n39746, n39747,
         n39748, n39749, n39750, n39751, n39752, n39753, n39754, n39755,
         n39756, n39757, n39758, n39759, n39760, n39761, n39762, n39763,
         n39764, n39765, n39766, n39767, n39768, n39769, n39770, n39771,
         n39772, n39773, n39774, n39775, n39776, n39777, n39778, n39779,
         n39780, n39781, n39782, n39783, n39784, n39785, n39786, n39787,
         n39788, n39789, n39790, n39791, n39792, n39793, n39794, n39795,
         n39796, n39797, n39798, n39799, n39800, n39801, n39802, n39803,
         n39804, n39805, n39806, n39807, n39808, n39809, n39810, n39811,
         n39812, n39813, n39814, n39815, n39816, n39817, n39818, n39819,
         n39820, n39821, n39822, n39823, n39824, n39825, n39826, n39827,
         n39828, n39829, n39830, n39831, n39832, n39833, n39834, n39835,
         n39836, n39837, n39838, n39839, n39840, n39841, n39842, n39843,
         n39844, n39845, n39846, n39847, n39848, n39849, n39850, n39851,
         n39852, n39853, n39854, n39855, n39856, n39857, n39858, n39859,
         n39860, n39861, n39862, n39863, n39864, n39865, n39866, n39867,
         n39868, n39869, n39870, n39871, n39872, n39873, n39874, n39875,
         n39876, n39877, n39878, n39879, n39880, n39881, n39882, n39883,
         n39884, n39885, n39886, n39887, n39888, n39889, n39890, n39891,
         n39892, n39893, n39894, n39895, n39896, n39897, n39898, n39899,
         n39900, n39901, n39902, n39903, n39904, n39905, n39906, n39907,
         n39908, n39909, n39910, n39911, n39912, n39913, n39914, n39915,
         n39916, n39917, n39918, n39919, n39920, n39921, n39922, n39923,
         n39924, n39925, n39926, n39927, n39928, n39929, n39930, n39931,
         n39932, n39933, n39934, n39935, n39936, n39937, n39938, n39939,
         n39940, n39941, n39942, n39943, n39944, n39945, n39946, n39947,
         n39948, n39949, n39950, n39951, n39952, n39953, n39954, n39955,
         n39956, n39957, n39958, n39959, n39960, n39961, n39962, n39963,
         n39964, n39965, n39966, n39967, n39968, n39969, n39970, n39971,
         n39972, n39973, n39974, n39975, n39976, n39977, n39978, n39979,
         n39980, n39981, n39982, n39983, n39984, n39985, n39986, n39987,
         n39988, n39989, n39990, n39991, n39992, n39993, n39994, n39995,
         n39996, n39997, n39998, n39999, n40000, n40001, n40002, n40003,
         n40004, n40005, n40006, n40007, n40008, n40009, n40010, n40011,
         n40012, n40013, n40014, n40015, n40016, n40017, n40018, n40019,
         n40020, n40021, n40022, n40023, n40024, n40025, n40026, n40027,
         n40028, n40029, n40030, n40031, n40032, n40033, n40034, n40035,
         n40036, n40037, n40038, n40039, n40040, n40041, n40042, n40043,
         n40044, n40045, n40046, n40047, n40048, n40049, n40050, n40051,
         n40052, n40053, n40054, n40055, n40056, n40057, n40058, n40059,
         n40060, n40061, n40062, n40063, n40064, n40065, n40066, n40067,
         n40068, n40069, n40070, n40071, n40072, n40073, n40074, n40075,
         n40076, n40077, n40078, n40079, n40080, n40081, n40082, n40083,
         n40084, n40085, n40086, n40087, n40088, n40089, n40090, n40091,
         n40092, n40093, n40094, n40095, n40096, n40097, n40098, n40099,
         n40100, n40101, n40102, n40103, n40104, n40105, n40106, n40107,
         n40108, n40109, n40110, n40111, n40112, n40113, n40114, n40115,
         n40116, n40117, n40118, n40119, n40120, n40121, n40122, n40123,
         n40124, n40125, n40126, n40127, n40128, n40129, n40130, n40131,
         n40132, n40133, n40134, n40135, n40136, n40137, n40138, n40139,
         n40140, n40141, n40142, n40143, n40144, n40145, n40146, n40147,
         n40148, n40149, n40150, n40151, n40152, n40153, n40154, n40155,
         n40156, n40157, n40158, n40159, n40160, n40161, n40162, n40163,
         n40164, n40165, n40166, n40167, n40168, n40169, n40170, n40171,
         n40172, n40173, n40174, n40175, n40176, n40177, n40178, n40179,
         n40180, n40181, n40182, n40183, n40184, n40185, n40186, n40187,
         n40188, n40189, n40190, n40191, n40192, n40193, n40194, n40195,
         n40196, n40197, n40198, n40199, n40200, n40201, n40202, n40203,
         n40204, n40205, n40206, n40207, n40208, n40209, n40210, n40211,
         n40212, n40213, n40214, n40215, n40216, n40217, n40218, n40219,
         n40220, n40221, n40222, n40223, n40224, n40225, n40226, n40227,
         n40228, n40229, n40230, n40231, n40232, n40233, n40234, n40235,
         n40236, n40237, n40238, n40239, n40240, n40241, n40242, n40243,
         n40244, n40245, n40246, n40247, n40248, n40249, n40250, n40251,
         n40252, n40253, n40254, n40255, n40256, n40257, n40258, n40259,
         n40260, n40261, n40262, n40263, n40264, n40265, n40266, n40267,
         n40268, n40269, n40270, n40271, n40272, n40273, n40274, n40275,
         n40276, n40277, n40278, n40279, n40280, n40281, n40282, n40283,
         n40284, n40285, n40286, n40287, n40288, n40289, n40290, n40291,
         n40292, n40293, n40294, n40295, n40296, n40297, n40298, n40299,
         n40300, n40301, n40302, n40303, n40304, n40305, n40306, n40307,
         n40308, n40309, n40310, n40311, n40312, n40313, n40314, n40315,
         n40316, n40317, n40318, n40319, n40320, n40321, n40322, n40323,
         n40324, n40325, n40326, n40327, n40328, n40329, n40330, n40331,
         n40332, n40333, n40334, n40335, n40336, n40337, n40338, n40339,
         n40340, n40341, n40342, n40343, n40344, n40345, n40346, n40347,
         n40348, n40349, n40350, n40351, n40352, n40353, n40354, n40355,
         n40356, n40357, n40358, n40359, n40360, n40361, n40362, n40363,
         n40364, n40365, n40366, n40367, n40368, n40369, n40370, n40371,
         n40372, n40373, n40374, n40375, n40376, n40377, n40378, n40379,
         n40380, n40381, n40382, n40383, n40384, n40385, n40386, n40387,
         n40388, n40389, n40390, n40391, n40392, n40393, n40394, n40395,
         n40396, n40397, n40398, n40399, n40400, n40401, n40402, n40403,
         n40404, n40405, n40406, n40407, n40408, n40409, n40410, n40411,
         n40412, n40413, n40414, n40415, n40416, n40417, n40418, n40419,
         n40420, n40421, n40422, n40423, n40424, n40425, n40426, n40427,
         n40428, n40429, n40430, n40431, n40432, n40433, n40434, n40435,
         n40436, n40437, n40438, n40439, n40440, n40441, n40442, n40443,
         n40444, n40445, n40446, n40447, n40448, n40449, n40450, n40451,
         n40452, n40453, n40454, n40455, n40456, n40457, n40458, n40459,
         n40460, n40461, n40462, n40463, n40464, n40465, n40466, n40467,
         n40468, n40469, n40470, n40471, n40472, n40473, n40474, n40475,
         n40476, n40477, n40478, n40479, n40480, n40481, n40482, n40483,
         n40484, n40485, n40486, n40487, n40488, n40489, n40490, n40491,
         n40492, n40493, n40494, n40495, n40496, n40497, n40498, n40499,
         n40500, n40501, n40502, n40503, n40504, n40505, n40506, n40507,
         n40508, n40509, n40510, n40511, n40512, n40513, n40514, n40515,
         n40516, n40517, n40518, n40519, n40520, n40521, n40522, n40523,
         n40524, n40525, n40526, n40527, n40528, n40529, n40530, n40531,
         n40532, n40533, n40534, n40535, n40536, n40537, n40538, n40539,
         n40540, n40541, n40542, n40543, n40544, n40545, n40546, n40547,
         n40548, n40549, n40550, n40551, n40552, n40553, n40554, n40555,
         n40556, n40557, n40558, n40559, n40560, n40561, n40562, n40563,
         n40564, n40565, n40566, n40567, n40568, n40569, n40570, n40571,
         n40572, n40573, n40574, n40575, n40576, n40577, n40578, n40579,
         n40580, n40581, n40582, n40583, n40584, n40585, n40586, n40587,
         n40588, n40589, n40590, n40591, n40592, n40593, n40594, n40595,
         n40596, n40597, n40598, n40599, n40600, n40601, n40602, n40603,
         n40604, n40605, n40606, n40607, n40608, n40609, n40610, n40611,
         n40612, n40613, n40614, n40615, n40616, n40617, n40618, n40619,
         n40620, n40621, n40622, n40623, n40624, n40625, n40626, n40627,
         n40628, n40629, n40630, n40631, n40632, n40633, n40634, n40635,
         n40636, n40637, n40638, n40639, n40640, n40641, n40642, n40643,
         n40644, n40645, n40646, n40647, n40648, n40649, n40650, n40651,
         n40652, n40653, n40654, n40655, n40656, n40657, n40658, n40659,
         n40660, n40661, n40662, n40663, n40664, n40665, n40666, n40667,
         n40668, n40669, n40670, n40671, n40672, n40673, n40674, n40675,
         n40676, n40677, n40678, n40679, n40680, n40681, n40682, n40683,
         n40684, n40685, n40686, n40687, n40688, n40689, n40690, n40691,
         n40692, n40693, n40694, n40695, n40696, n40697, n40698, n40699,
         n40700, n40701, n40702, n40703, n40704, n40705, n40706, n40707,
         n40708, n40709, n40710, n40711, n40712, n40713, n40714, n40715,
         n40716, n40717, n40718, n40719, n40720, n40721, n40722, n40723,
         n40724, n40725, n40726, n40727, n40728, n40729, n40730, n40731,
         n40732, n40733, n40734, n40735, n40736, n40737, n40738, n40739,
         n40740, n40741, n40742, n40743, n40744, n40745, n40746, n40747,
         n40748, n40749, n40750, n40751, n40752, n40753, n40754, n40755,
         n40756, n40757, n40758, n40759, n40760, n40761, n40762, n40763,
         n40764, n40765, n40766, n40767, n40768, n40769, n40770, n40771,
         n40772, n40773, n40774, n40775, n40776, n40777, n40778, n40779,
         n40780, n40781, n40782, n40783, n40784, n40785, n40786, n40787,
         n40788, n40789, n40790, n40791, n40792, n40793, n40794, n40795,
         n40796, n40797, n40798, n40799, n40800, n40801, n40802, n40803,
         n40804, n40805, n40806, n40807, n40808, n40809, n40810, n40811,
         n40812, n40813, n40814, n40815, n40816, n40817, n40818, n40819,
         n40820, n40821, n40822, n40823, n40824, n40825, n40826, n40827,
         n40828, n40829, n40830, n40831, n40832, n40833, n40834, n40835,
         n40836, n40837, n40838, n40839, n40840, n40841, n40842, n40843,
         n40844, n40845, n40846, n40847, n40848, n40849, n40850, n40851,
         n40852, n40853, n40854, n40855, n40856, n40857, n40858, n40859,
         n40860, n40861, n40862, n40863, n40864, n40865, n40866, n40867,
         n40868, n40869, n40870, n40871, n40872, n40873, n40874, n40875,
         n40876, n40877, n40878, n40879, n40880, n40881, n40882, n40883,
         n40884, n40885, n40886, n40887, n40888, n40889, n40890, n40891,
         n40892, n40893, n40894, n40895, n40896, n40897, n40898, n40899,
         n40900, n40901, n40902, n40903, n40904, n40905, n40906, n40907,
         n40908, n40909, n40910, n40911, n40912, n40913, n40914, n40915,
         n40916, n40917, n40918, n40919, n40920, n40921, n40922, n40923,
         n40924, n40925, n40926, n40927, n40928, n40929, n40930, n40931,
         n40932, n40933, n40934, n40935, n40936, n40937, n40938, n40939,
         n40940, n40941, n40942, n40943, n40944, n40945, n40946, n40947,
         n40948, n40949, n40950, n40951, n40952, n40953, n40954, n40955,
         n40956, n40957, n40958, n40959, n40960, n40961, n40962, n40963,
         n40964, n40965, n40966, n40967, n40968, n40969, n40970, n40971,
         n40972, n40973, n40974, n40975, n40976, n40977, n40978, n40979,
         n40980, n40981, n40982, n40983, n40984, n40985, n40986, n40987,
         n40988, n40989, n40990, n40991, n40992, n40993, n40994, n40995,
         n40996, n40997, n40998, n40999, n41000, n41001, n41002, n41003,
         n41004, n41005, n41006, n41007, n41008, n41009, n41010, n41011,
         n41012, n41013, n41014, n41015, n41016, n41017, n41018, n41019,
         n41020, n41021, n41022, n41023, n41024, n41025, n41026, n41027,
         n41028, n41029, n41030, n41031, n41032, n41033, n41034, n41035,
         n41036, n41037, n41038, n41039, n41040, n41041, n41042, n41043,
         n41044, n41045, n41046, n41047, n41048, n41049, n41050, n41051,
         n41052, n41053, n41054, n41055, n41056, n41057, n41058, n41059,
         n41060, n41061, n41062, n41063, n41064, n41065, n41066, n41067,
         n41068, n41069, n41070, n41071, n41072, n41073, n41074, n41075,
         n41076, n41077, n41078, n41079, n41080, n41081, n41082, n41083,
         n41084, n41085, n41086, n41087, n41088, n41089, n41090, n41091,
         n41092, n41093, n41094, n41095, n41096, n41097, n41098, n41099,
         n41100, n41101, n41102, n41103, n41104, n41105, n41106, n41107,
         n41108, n41109, n41110, n41111, n41112, n41113, n41114, n41115,
         n41116, n41117, n41118, n41119, n41120, n41121, n41122, n41123,
         n41124, n41125, n41126, n41127, n41128, n41129, n41130, n41131,
         n41132, n41133, n41134, n41135, n41136, n41137, n41138, n41139,
         n41140, n41141, n41142, n41143, n41144, n41145, n41146, n41147,
         n41148, n41149, n41150, n41151, n41152, n41153, n41154, n41155,
         n41156, n41157, n41158, n41159, n41160, n41161, n41162, n41163,
         n41164, n41165, n41166, n41167, n41168, n41169, n41170, n41171,
         n41172, n41173, n41174, n41175, n41176, n41177, n41178, n41179,
         n41180, n41181, n41182, n41183, n41184, n41185, n41186, n41187,
         n41188, n41189, n41190, n41191, n41192, n41193, n41194, n41195,
         n41196, n41197, n41198, n41199, n41200, n41201, n41202, n41203,
         n41204, n41205, n41206, n41207, n41208, n41209, n41210, n41211,
         n41212, n41213, n41214, n41215, n41216, n41217, n41218, n41219,
         n41220, n41221, n41222, n41223, n41224, n41225, n41226, n41227,
         n41228, n41229, n41230, n41231, n41232, n41233, n41234, n41235,
         n41236, n41237, n41238, n41239, n41240, n41241, n41242, n41243,
         n41244, n41245, n41246, n41247, n41248, n41249, n41250, n41251,
         n41252, n41253, n41254, n41255, n41256, n41257, n41258, n41259,
         n41260, n41261, n41262, n41263, n41264, n41265, n41266, n41267,
         n41268, n41269, n41270, n41271, n41272, n41273, n41274, n41275,
         n41276, n41277, n41278, n41279, n41280, n41281, n41282, n41283,
         n41284, n41285, n41286, n41287, n41288, n41289, n41290, n41291,
         n41292, n41293, n41294, n41295, n41296, n41297, n41298, n41299,
         n41300, n41301, n41302, n41303, n41304, n41305, n41306, n41307,
         n41308, n41309, n41310, n41311, n41312, n41313, n41314, n41315,
         n41316, n41317, n41318, n41319, n41320, n41321, n41322, n41323,
         n41324, n41325, n41326, n41327, n41328, n41329, n41330, n41331,
         n41332, n41333, n41334, n41335, n41336, n41337, n41338, n41339,
         n41340, n41341, n41342, n41343, n41344, n41345, n41346, n41347,
         n41348, n41349, n41350, n41351, n41352, n41353, n41354, n41355,
         n41356, n41357, n41358, n41359, n41360, n41361, n41362, n41363,
         n41364, n41365, n41366, n41367, n41368, n41369, n41370, n41371,
         n41372, n41373, n41374, n41375, n41376, n41377, n41378, n41379,
         n41380, n41381, n41382, n41383, n41384, n41385, n41386, n41387,
         n41388, n41389, n41390, n41391, n41392, n41393, n41394, n41395,
         n41396, n41397, n41398, n41399, n41400, n41401, n41402, n41403,
         n41404, n41405, n41406, n41407, n41408, n41409, n41410, n41411,
         n41412, n41413, n41414, n41415, n41416, n41417, n41418, n41419,
         n41420, n41421, n41422, n41423, n41424, n41425, n41426, n41427,
         n41428, n41429, n41430, n41431, n41432, n41433, n41434, n41435,
         n41436, n41437, n41438, n41439, n41440, n41441, n41442, n41443,
         n41444, n41445, n41446, n41447, n41448, n41449, n41450, n41451,
         n41452, n41453, n41454, n41455, n41456, n41457, n41458, n41459,
         n41460, n41461, n41462, n41463, n41464, n41465, n41466, n41467,
         n41468, n41469, n41470, n41471, n41472, n41473, n41474, n41475,
         n41476, n41477, n41478, n41479, n41480, n41481, n41482, n41483,
         n41484, n41485, n41486, n41487, n41488, n41489, n41490, n41491,
         n41492, n41493, n41494, n41495, n41496, n41497, n41498, n41499,
         n41500, n41501, n41502, n41503, n41504, n41505, n41506, n41507,
         n41508, n41509, n41510, n41511, n41512, n41513, n41514, n41515,
         n41516, n41517, n41518, n41519, n41520, n41521, n41522, n41523,
         n41524, n41525, n41526, n41527, n41528, n41529, n41530, n41531,
         n41532, n41533, n41534, n41535, n41536, n41537, n41538, n41539,
         n41540, n41541, n41542, n41543, n41544, n41545, n41546, n41547,
         n41548, n41549, n41550, n41551, n41552, n41553, n41554, n41555,
         n41556, n41557, n41558, n41559, n41560, n41561, n41562, n41563,
         n41564, n41565, n41566, n41567, n41568, n41569, n41570, n41571,
         n41572, n41573, n41574, n41575, n41576, n41577, n41578, n41579,
         n41580, n41581, n41582, n41583, n41584, n41585, n41586, n41587,
         n41588, n41589, n41590, n41591, n41592, n41593, n41594, n41595,
         n41596, n41597, n41598, n41599, n41600, n41601, n41602, n41603,
         n41604, n41605, n41606, n41607, n41608, n41609, n41610, n41611,
         n41612, n41613, n41614, n41615, n41616, n41617, n41618, n41619,
         n41620, n41621, n41622, n41623, n41624, n41625, n41626, n41627,
         n41628, n41629, n41630, n41631, n41632, n41633, n41634, n41635,
         n41636, n41637, n41638, n41639, n41640, n41641, n41642, n41643,
         n41644, n41645, n41646, n41647, n41648, n41649, n41650, n41651,
         n41652, n41653, n41654, n41655, n41656, n41657, n41658, n41659,
         n41660, n41661, n41662, n41663, n41664, n41665, n41666, n41667,
         n41668, n41669, n41670, n41671, n41672, n41673, n41674, n41675,
         n41676, n41677, n41678, n41679, n41680, n41681, n41682, n41683,
         n41684, n41685, n41686, n41687, n41688, n41689, n41690, n41691,
         n41692, n41693, n41694, n41695, n41696, n41697, n41698, n41699,
         n41700, n41701, n41702, n41703, n41704, n41705, n41706, n41707,
         n41708, n41709, n41710, n41711, n41712, n41713, n41714, n41715,
         n41716, n41717, n41718, n41719, n41720, n41721, n41722, n41723,
         n41724, n41725, n41726, n41727, n41728, n41729, n41730, n41731,
         n41732, n41733, n41734, n41735, n41736, n41737, n41738, n41739,
         n41740, n41741, n41742, n41743, n41744, n41745, n41746, n41747,
         n41748, n41749, n41750, n41751, n41752, n41753, n41754, n41755,
         n41756, n41757, n41758, n41759, n41760, n41761, n41762, n41763,
         n41764, n41765, n41766, n41767, n41768, n41769, n41770, n41771,
         n41772, n41773, n41774, n41775, n41776, n41777, n41778, n41779,
         n41780, n41781, n41782, n41783, n41784, n41785, n41786, n41787,
         n41788, n41789, n41790, n41791, n41792, n41793, n41794, n41795,
         n41796, n41797, n41798, n41799, n41800, n41801, n41802, n41803,
         n41804, n41805, n41806, n41807, n41808, n41809, n41810, n41811,
         n41812, n41813, n41814, n41815, n41816, n41817, n41818, n41819,
         n41820, n41821, n41822, n41823, n41824, n41825, n41826, n41827,
         n41828, n41829, n41830, n41831, n41832, n41833, n41834, n41835,
         n41836, n41837, n41838, n41839, n41840, n41841, n41842, n41843,
         n41844, n41845, n41846, n41847, n41848, n41849, n41850, n41851,
         n41852, n41853, n41854, n41855, n41856, n41857, n41858, n41859,
         n41860, n41861, n41862, n41863, n41864, n41865, n41866, n41867,
         n41868, n41869, n41870, n41871, n41872, n41873, n41874, n41875,
         n41876, n41877, n41878, n41879, n41880, n41881, n41882, n41883,
         n41884, n41885, n41886, n41887, n41888, n41889, n41890, n41891,
         n41892, n41893, n41894, n41895, n41896, n41897, n41898, n41899,
         n41900, n41901, n41902, n41903, n41904, n41905, n41906, n41907,
         n41908, n41909, n41910, n41911, n41912, n41913, n41914, n41915,
         n41916, n41917, n41918, n41919, n41920, n41921, n41922, n41923,
         n41924, n41925, n41926, n41927, n41928, n41929, n41930, n41931,
         n41932, n41933, n41934, n41935, n41936, n41937, n41938, n41939,
         n41940, n41941, n41942, n41943, n41944, n41945, n41946, n41947,
         n41948, n41949, n41950, n41951, n41952, n41953, n41954, n41955,
         n41956, n41957, n41958, n41959, n41960, n41961, n41962, n41963,
         n41964, n41965, n41966, n41967, n41968, n41969, n41970, n41971,
         n41972, n41973, n41974, n41975, n41976, n41977, n41978, n41979,
         n41980, n41981, n41982, n41983, n41984, n41985, n41986, n41987,
         n41988, n41989, n41990, n41991, n41992, n41993, n41994, n41995,
         n41996, n41997, n41998, n41999, n42000, n42001, n42002, n42003,
         n42004, n42005, n42006, n42007, n42008, n42009, n42010, n42011,
         n42012, n42013, n42014, n42015, n42016, n42017, n42018, n42019,
         n42020, n42021, n42022, n42023, n42024, n42025, n42026, n42027,
         n42028, n42029, n42030, n42031, n42032, n42033, n42034, n42035,
         n42036, n42037, n42038, n42039, n42040, n42041, n42042, n42043,
         n42044, n42045, n42046, n42047, n42048, n42049, n42050, n42051,
         n42052, n42053, n42054, n42055, n42056, n42057, n42058, n42059,
         n42060, n42061, n42062, n42063, n42064, n42065, n42066, n42067,
         n42068, n42069, n42070, n42071, n42072, n42073, n42074, n42075,
         n42076, n42077, n42078, n42079, n42080, n42081, n42082, n42083,
         n42084, n42085, n42086, n42087, n42088, n42089, n42090, n42091,
         n42092, n42093, n42094, n42095, n42096, n42097, n42098, n42099,
         n42100, n42101, n42102, n42103, n42104, n42105, n42106, n42107,
         n42108, n42109, n42110, n42111, n42112, n42113, n42114, n42115,
         n42116, n42117, n42118, n42119, n42120, n42121, n42122, n42123,
         n42124, n42125, n42126, n42127, n42128, n42129, n42130, n42131,
         n42132, n42133, n42134, n42135, n42136, n42137, n42138, n42139,
         n42140, n42141, n42142, n42143, n42144, n42145, n42146, n42147,
         n42148, n42149, n42150, n42151, n42152, n42153, n42154, n42155,
         n42156, n42157, n42158, n42159, n42160, n42161, n42162, n42163,
         n42164, n42165, n42166, n42167, n42168, n42169, n42170, n42171,
         n42172, n42173, n42174, n42175, n42176, n42177, n42178, n42179,
         n42180, n42181, n42182, n42183, n42184, n42185, n42186, n42187,
         n42188, n42189, n42190, n42191, n42192, n42193, n42194, n42195,
         n42196, n42197, n42198, n42199, n42200, n42201, n42202, n42203,
         n42204, n42205, n42206, n42207, n42208, n42209, n42210, n42211,
         n42212, n42213, n42214, n42215, n42216, n42217, n42218, n42219,
         n42220, n42221, n42222, n42223, n42224, n42225, n42226, n42227,
         n42228, n42229, n42230, n42231, n42232, n42233, n42234, n42235,
         n42236, n42237, n42238, n42239, n42240, n42241, n42242, n42243,
         n42244, n42245, n42246, n42247, n42248, n42249, n42250, n42251,
         n42252, n42253, n42254, n42255, n42256, n42257, n42258, n42259,
         n42260, n42261, n42262, n42263, n42264, n42265, n42266, n42267,
         n42268, n42269, n42270, n42271, n42272, n42273, n42274, n42275,
         n42276, n42277, n42278, n42279, n42280, n42281, n42282, n42283,
         n42284, n42285, n42286, n42287, n42288, n42289, n42290, n42291,
         n42292, n42293, n42294, n42295, n42296, n42297, n42298, n42299,
         n42300, n42301, n42302, n42303, n42304, n42305, n42306, n42307,
         n42308, n42309, n42310, n42311, n42312, n42313, n42314, n42315,
         n42316, n42317, n42318, n42319, n42320, n42321, n42322, n42323,
         n42324, n42325, n42326, n42327, n42328, n42329, n42330, n42331,
         n42332, n42333, n42334, n42335, n42336, n42337, n42338, n42339,
         n42340, n42341, n42342, n42343, n42344, n42345, n42346, n42347,
         n42348, n42349, n42350, n42351, n42352, n42353, n42354, n42355,
         n42356, n42357, n42358, n42359, n42360, n42361, n42362, n42363,
         n42364, n42365, n42366, n42367, n42368, n42369, n42370, n42371,
         n42372, n42373, n42374, n42375, n42376, n42377, n42378, n42379,
         n42380, n42381, n42382, n42383, n42384, n42385, n42386, n42387,
         n42388, n42389, n42390, n42391, n42392, n42393, n42394, n42395,
         n42396, n42397, n42398, n42399, n42400, n42401, n42402, n42403,
         n42404, n42405, n42406, n42407, n42408, n42409, n42410, n42411,
         n42412, n42413, n42414, n42415, n42416, n42417, n42418, n42419,
         n42420, n42421, n42422, n42423, n42424, n42425, n42426, n42427,
         n42428, n42429, n42430, n42431, n42432, n42433, n42434, n42435,
         n42436, n42437, n42438, n42439, n42440, n42441, n42442, n42443,
         n42444, n42445, n42446, n42447, n42448, n42449, n42450, n42451,
         n42452, n42453, n42454, n42455, n42456, n42457, n42458, n42459,
         n42460, n42461, n42462, n42463, n42464, n42465, n42466, n42467,
         n42468, n42469, n42470, n42471, n42472, n42473, n42474, n42475,
         n42476, n42477, n42478, n42479, n42480, n42481, n42482, n42483,
         n42484, n42485, n42486, n42487, n42488, n42489, n42490, n42491,
         n42492, n42493, n42494, n42495, n42496, n42497, n42498, n42499,
         n42500, n42501, n42502, n42503, n42504, n42505, n42506, n42507,
         n42508, n42509, n42510, n42511, n42512, n42513, n42514, n42515,
         n42516, n42517, n42518, n42519, n42520, n42521, n42522, n42523,
         n42524, n42525, n42526, n42527, n42528, n42529, n42530, n42531,
         n42532, n42533, n42534, n42535, n42536, n42537, n42538, n42539,
         n42540, n42541, n42542, n42543, n42544, n42545, n42546, n42547,
         n42548, n42549, n42550, n42551, n42552, n42553, n42554, n42555,
         n42556, n42557, n42558, n42559, n42560, n42561, n42562, n42563,
         n42564, n42565, n42566, n42567, n42568, n42569, n42570, n42571,
         n42572, n42573, n42574, n42575, n42576, n42577, n42578, n42579,
         n42580, n42581, n42582, n42583, n42584, n42585, n42586, n42587,
         n42588, n42589, n42590, n42591, n42592, n42593, n42594, n42595,
         n42596, n42597, n42598, n42599, n42600, n42601, n42602, n42603,
         n42604, n42605, n42606, n42607, n42608, n42609, n42610, n42611,
         n42612, n42613, n42614, n42615, n42616, n42617, n42618, n42619,
         n42620, n42621, n42622, n42623, n42624, n42625, n42626, n42627,
         n42628, n42629, n42630, n42631, n42632, n42633, n42634, n42635,
         n42636, n42637, n42638, n42639, n42640, n42641, n42642, n42643,
         n42644, n42645, n42646, n42647, n42648, n42649, n42650, n42651,
         n42652, n42653, n42654, n42655, n42656, n42657, n42658, n42659,
         n42660, n42661, n42662, n42663, n42664, n42665, n42666, n42667,
         n42668, n42669, n42670, n42671, n42672, n42673, n42674, n42675,
         n42676, n42677, n42678, n42679, n42680, n42681, n42682, n42683,
         n42684, n42685, n42686, n42687, n42688, n42689, n42690, n42691,
         n42692, n42693, n42694, n42695, n42696, n42697, n42698, n42699,
         n42700, n42701, n42702, n42703, n42704, n42705, n42706, n42707,
         n42708, n42709, n42710, n42711, n42712, n42713, n42714, n42715,
         n42716, n42717, n42718, n42719, n42720, n42721, n42722, n42723,
         n42724, n42725, n42726, n42727, n42728, n42729, n42730, n42731,
         n42732, n42733, n42734, n42735, n42736, n42737, n42738, n42739,
         n42740, n42741, n42742, n42743, n42744, n42745, n42746, n42747,
         n42748, n42749, n42750, n42751, n42752, n42753, n42754, n42755,
         n42756, n42757, n42758, n42759, n42760, n42761, n42762, n42763,
         n42764, n42765, n42766, n42767, n42768, n42769, n42770, n42771,
         n42772, n42773, n42774, n42775, n42776, n42777, n42778, n42779,
         n42780, n42781, n42782, n42783, n42784, n42785, n42786, n42787,
         n42788, n42789, n42790, n42791, n42792, n42793, n42794, n42795,
         n42796, n42797, n42798, n42799, n42800, n42801, n42802, n42803,
         n42804, n42805, n42806, n42807, n42808, n42809, n42810, n42811,
         n42812, n42813, n42814, n42815, n42816, n42817, n42818, n42819,
         n42820, n42821, n42822, n42823, n42824, n42825, n42826, n42827,
         n42828, n42829, n42830, n42831, n42832, n42833, n42834, n42835,
         n42836, n42837, n42838, n42839, n42840, n42841, n42842, n42843,
         n42844, n42845, n42846, n42847, n42848, n42849, n42850, n42851,
         n42852, n42853, n42854, n42855, n42856, n42857, n42858, n42859,
         n42860, n42861, n42862, n42863, n42864, n42865, n42866, n42867,
         n42868, n42869, n42870, n42871, n42872, n42873, n42874, n42875,
         n42876, n42877, n42878, n42879, n42880, n42881, n42882, n42883,
         n42884, n42885, n42886, n42887, n42888, n42889, n42890, n42891,
         n42892, n42893, n42894, n42895, n42896, n42897, n42898, n42899,
         n42900, n42901, n42902, n42903, n42904, n42905, n42906, n42907,
         n42908, n42909, n42910, n42911, n42912, n42913, n42914, n42915,
         n42916, n42917, n42918, n42919, n42920, n42921, n42922, n42923,
         n42924, n42925, n42926, n42927, n42928, n42929, n42930, n42931,
         n42932, n42933, n42934, n42935, n42936, n42937, n42938, n42939,
         n42940, n42941, n42942, n42943, n42944, n42945, n42946, n42947,
         n42948, n42949, n42950, n42951, n42952, n42953, n42954, n42955,
         n42956, n42957, n42958, n42959, n42960, n42961, n42962, n42963,
         n42964, n42965, n42966, n42967, n42968, n42969, n42970, n42971,
         n42972, n42973, n42974, n42975, n42976, n42977, n42978, n42979,
         n42980, n42981, n42982, n42983, n42984, n42985, n42986, n42987,
         n42988, n42989, n42990, n42991, n42992, n42993, n42994, n42995,
         n42996, n42997, n42998, n42999, n43000, n43001, n43002, n43003,
         n43004, n43005, n43006, n43007, n43008, n43009, n43010, n43011,
         n43012, n43013, n43014, n43015, n43016, n43017, n43018, n43019,
         n43020, n43021, n43022, n43023, n43024, n43025, n43026, n43027,
         n43028, n43029, n43030, n43031, n43032, n43033, n43034, n43035,
         n43036, n43037, n43038, n43039, n43040, n43041, n43042, n43043,
         n43044, n43045, n43046, n43047, n43048, n43049, n43050, n43051,
         n43052, n43053, n43054, n43055, n43056, n43057, n43058, n43059,
         n43060, n43061, n43062, n43063, n43064, n43065, n43066, n43067,
         n43068, n43069, n43070, n43071, n43072, n43073, n43074, n43075,
         n43076, n43077, n43078, n43079, n43080, n43081, n43082, n43083,
         n43084, n43085, n43086, n43087, n43088, n43089, n43090, n43091,
         n43092, n43093, n43094, n43095, n43096, n43097, n43098, n43099,
         n43100, n43101, n43102, n43103, n43104, n43105, n43106, n43107,
         n43108, n43109, n43110, n43111, n43112, n43113, n43114, n43115,
         n43116, n43117, n43118, n43119, n43120, n43121, n43122, n43123,
         n43124, n43125, n43126, n43127, n43128, n43129, n43130, n43131,
         n43132, n43133, n43134, n43135, n43136, n43137, n43138, n43139,
         n43140, n43141, n43142, n43143, n43144, n43145, n43146, n43147,
         n43148, n43149, n43150, n43151, n43152, n43153, n43154, n43155,
         n43156, n43157, n43158, n43159, n43160, n43161, n43162, n43163,
         n43164, n43165, n43166, n43167, n43168, n43169, n43170, n43171,
         n43172, n43173, n43174, n43175, n43176, n43177, n43178, n43179,
         n43180, n43181, n43182, n43183, n43184, n43185, n43186, n43187,
         n43188, n43189, n43190, n43191, n43192, n43193, n43194, n43195,
         n43196, n43197, n43198, n43199, n43200, n43201, n43202, n43203,
         n43204, n43205, n43206, n43207, n43208, n43209, n43210, n43211,
         n43212, n43213, n43214, n43215, n43216, n43217, n43218, n43219,
         n43220, n43221, n43222, n43223, n43224, n43225, n43226, n43227,
         n43228, n43229, n43230, n43231, n43232, n43233, n43234, n43235,
         n43236, n43237, n43238, n43239, n43240, n43241, n43242, n43243,
         n43244, n43245, n43246, n43247, n43248, n43249, n43250, n43251,
         n43252, n43253, n43254, n43255, n43256, n43257, n43258, n43259,
         n43260, n43261, n43262, n43263, n43264, n43265, n43266, n43267,
         n43268, n43269, n43270, n43271, n43272, n43273, n43274, n43275,
         n43276, n43277, n43278, n43279, n43280, n43281, n43282, n43283,
         n43284, n43285, n43286, n43287, n43288, n43289, n43290, n43291,
         n43292, n43293, n43294, n43295, n43296, n43297, n43298, n43299,
         n43300, n43301, n43302, n43303, n43304, n43305, n43306, n43307,
         n43308, n43309, n43310, n43311, n43312, n43313, n43314, n43315,
         n43316, n43317, n43318, n43319, n43320, n43321, n43322, n43323,
         n43324, n43325, n43326, n43327, n43328, n43329, n43330, n43331,
         n43332, n43333, n43334, n43335, n43336, n43337, n43338, n43339,
         n43340, n43341, n43342, n43343, n43344, n43345, n43346, n43347,
         n43348, n43349, n43350, n43351, n43352, n43353, n43354, n43355,
         n43356, n43357, n43358, n43359, n43360, n43361, n43362, n43363,
         n43364, n43365, n43366, n43367, n43368, n43369, n43370, n43371,
         n43372, n43373, n43374, n43375, n43376, n43377, n43378, n43379,
         n43380, n43381, n43382, n43383, n43384, n43385, n43386, n43387,
         n43388, n43389, n43390, n43391, n43392, n43393, n43394, n43395,
         n43396, n43397, n43398, n43399, n43400, n43401, n43402, n43403,
         n43404, n43405, n43406, n43407, n43408, n43409, n43410, n43411,
         n43412, n43413, n43414, n43415, n43416, n43417, n43418, n43419,
         n43420, n43421, n43422, n43423, n43424, n43425, n43426, n43427,
         n43428, n43429, n43430, n43431, n43432, n43433, n43434, n43435,
         n43436, n43437, n43438, n43439, n43440, n43441, n43442, n43443,
         n43444, n43445, n43446, n43447, n43448, n43449, n43450, n43451,
         n43452, n43453, n43454, n43455, n43456, n43457, n43458, n43459,
         n43460, n43461, n43462, n43463, n43464, n43465, n43466, n43467,
         n43468, n43469, n43470, n43471, n43472, n43473, n43474, n43475,
         n43476, n43477, n43478, n43479, n43480, n43481, n43482, n43483,
         n43484, n43485, n43486, n43487, n43488, n43489, n43490, n43491,
         n43492, n43493, n43494, n43495, n43496, n43497, n43498, n43499,
         n43500, n43501, n43502, n43503, n43504, n43505, n43506, n43507,
         n43508, n43509, n43510, n43511, n43512, n43513, n43514, n43515,
         n43516, n43517, n43518, n43519, n43520, n43521, n43522, n43523,
         n43524, n43525, n43526, n43527, n43528, n43529, n43530, n43531,
         n43532, n43533, n43534, n43535, n43536, n43537, n43538, n43539,
         n43540, n43541, n43542, n43543, n43544, n43545, n43546, n43547,
         n43548, n43549, n43550, n43551, n43552, n43553, n43554, n43555,
         n43556, n43557, n43558, n43559, n43560, n43561, n43562, n43563,
         n43564, n43565, n43566, n43567, n43568, n43569, n43570, n43571,
         n43572, n43573, n43574, n43575, n43576, n43577, n43578, n43579,
         n43580, n43581, n43582, n43583, n43584, n43585, n43586, n43587,
         n43588, n43589, n43590, n43591, n43592, n43593, n43594, n43595,
         n43596, n43597, n43598, n43599, n43600, n43601, n43602, n43603,
         n43604, n43605, n43606, n43607, n43608, n43609, n43610, n43611,
         n43612, n43613, n43614, n43615, n43616, n43617, n43618, n43619,
         n43620, n43621, n43622, n43623, n43624, n43625, n43626, n43627,
         n43628, n43629, n43630, n43631, n43632, n43633, n43634, n43635,
         n43636, n43637, n43638, n43639, n43640, n43641, n43642, n43643,
         n43644, n43645, n43646, n43647, n43648, n43649, n43650, n43651,
         n43652, n43653, n43654, n43655, n43656, n43657, n43658, n43659,
         n43660, n43661, n43662, n43663, n43664, n43665, n43666, n43667,
         n43668, n43669, n43670, n43671, n43672, n43673, n43674, n43675,
         n43676, n43677, n43678, n43679, n43680, n43681, n43682, n43683,
         n43684, n43685, n43686, n43687, n43688, n43689, n43690, n43691,
         n43692, n43693, n43694, n43695, n43696, n43697, n43698, n43699,
         n43700, n43701, n43702, n43703, n43704, n43705, n43706, n43707,
         n43708, n43709, n43710, n43711, n43712, n43713, n43714, n43715,
         n43716, n43717, n43718, n43719, n43720, n43721, n43722, n43723,
         n43724, n43725, n43726, n43727, n43728, n43729, n43730, n43731,
         n43732, n43733, n43734, n43735, n43736, n43737, n43738, n43739,
         n43740, n43741, n43742, n43743, n43744, n43745, n43746, n43747,
         n43748, n43749, n43750, n43751, n43752, n43753, n43754, n43755,
         n43756, n43757, n43758, n43759, n43760, n43761, n43762, n43763,
         n43764, n43765, n43766, n43767, n43768, n43769, n43770, n43771,
         n43772, n43773, n43774, n43775, n43776, n43777, n43778, n43779,
         n43780, n43781, n43782, n43783, n43784, n43785, n43786, n43787,
         n43788, n43789, n43790, n43791, n43792, n43793, n43794, n43795,
         n43796, n43797, n43798, n43799, n43800, n43801, n43802, n43803,
         n43804, n43805, n43806, n43807, n43808, n43809, n43810, n43811,
         n43812, n43813, n43814, n43815, n43816, n43817, n43818, n43819,
         n43820, n43821, n43822, n43823, n43824, n43825, n43826, n43827,
         n43828, n43829, n43830, n43831, n43832, n43833, n43834, n43835,
         n43836, n43837, n43838, n43839, n43840, n43841, n43842, n43843,
         n43844, n43845, n43846, n43847, n43848, n43849, n43850, n43851,
         n43852, n43853, n43854, n43855, n43856, n43857, n43858, n43859,
         n43860, n43861, n43862, n43863, n43864, n43865, n43866, n43867,
         n43868, n43869, n43870, n43871, n43872, n43873, n43874, n43875,
         n43876, n43877, n43878, n43879, n43880, n43881, n43882, n43883,
         n43884, n43885, n43886, n43887, n43888, n43889, n43890, n43891,
         n43892, n43893, n43894, n43895, n43896, n43897, n43898, n43899,
         n43900, n43901, n43902, n43903, n43904, n43905, n43906, n43907,
         n43908, n43909, n43910, n43911, n43912, n43913, n43914, n43915,
         n43916, n43917, n43918, n43919, n43920, n43921, n43922, n43923,
         n43924, n43925, n43926, n43927, n43928, n43929, n43930, n43931,
         n43932, n43933, n43934, n43935, n43936, n43937, n43938, n43939,
         n43940, n43941, n43942, n43943, n43944, n43945, n43946, n43947,
         n43948, n43949, n43950, n43951, n43952, n43953, n43954, n43955,
         n43956, n43957, n43958, n43959, n43960, n43961, n43962, n43963,
         n43964, n43965, n43966, n43967, n43968, n43969, n43970, n43971,
         n43972, n43973, n43974, n43975, n43976, n43977, n43978, n43979,
         n43980, n43981, n43982, n43983, n43984, n43985, n43986, n43987,
         n43988, n43989, n43990, n43991, n43992, n43993, n43994, n43995,
         n43996, n43997, n43998, n43999, n44000, n44001, n44002, n44003,
         n44004, n44005, n44006, n44007, n44008, n44009, n44010, n44011,
         n44012, n44013, n44014, n44015, n44016, n44017, n44018, n44019,
         n44020, n44021, n44022, n44023, n44024, n44025, n44026, n44027,
         n44028, n44029, n44030, n44031, n44032, n44033, n44034, n44035,
         n44036, n44037, n44038, n44039, n44040, n44041, n44042, n44043,
         n44044, n44045, n44046, n44047, n44048, n44049, n44050, n44051,
         n44052, n44053, n44054, n44055, n44056, n44057, n44058, n44059,
         n44060, n44061, n44062, n44063, n44064, n44065, n44066, n44067,
         n44068, n44069, n44070, n44071, n44072, n44073, n44074, n44075,
         n44076, n44077, n44078, n44079, n44080, n44081, n44082, n44083,
         n44084, n44085, n44086, n44087, n44088, n44089, n44090, n44091,
         n44092, n44093, n44094, n44095, n44096, n44097, n44098, n44099,
         n44100, n44101, n44102, n44103, n44104, n44105, n44106, n44107,
         n44108, n44109, n44110, n44111, n44112, n44113, n44114, n44115,
         n44116, n44117, n44118, n44119, n44120, n44121, n44122, n44123,
         n44124, n44125, n44126, n44127, n44128, n44129, n44130, n44131,
         n44132, n44133, n44134, n44135, n44136, n44137, n44138, n44139,
         n44140, n44141, n44142, n44143, n44144, n44145, n44146, n44147,
         n44148, n44149, n44150, n44151, n44152, n44153, n44154, n44155,
         n44156, n44157, n44158, n44159, n44160, n44161, n44162, n44163,
         n44164, n44165, n44166, n44167, n44168, n44169, n44170, n44171,
         n44172, n44173, n44174, n44175, n44176, n44177, n44178, n44179,
         n44180, n44181, n44182, n44183, n44184, n44185, n44186, n44187,
         n44188, n44189, n44190, n44191, n44192, n44193, n44194, n44195,
         n44196, n44197, n44198, n44199, n44200, n44201, n44202, n44203,
         n44204, n44205, n44206, n44207, n44208, n44209, n44210, n44211,
         n44212, n44213, n44214, n44215, n44216, n44217, n44218, n44219,
         n44220, n44221, n44222, n44223, n44224, n44225, n44226, n44227,
         n44228, n44229, n44230, n44231, n44232, n44233, n44234, n44235,
         n44236, n44237, n44238, n44239, n44240, n44241, n44242, n44243,
         n44244, n44245, n44246, n44247, n44248, n44249, n44250, n44251,
         n44252, n44253, n44254, n44255, n44256, n44257, n44258, n44259,
         n44260, n44261, n44262, n44263, n44264, n44265, n44266, n44267,
         n44268, n44269, n44270, n44271, n44272, n44273, n44274, n44275,
         n44276, n44277, n44278, n44279, n44280, n44281, n44282, n44283,
         n44284, n44285, n44286, n44287, n44288, n44289, n44290, n44291,
         n44292, n44293, n44294, n44295, n44296, n44297, n44298, n44299,
         n44300, n44301, n44302, n44303, n44304, n44305, n44306, n44307,
         n44308, n44309, n44310, n44311, n44312, n44313, n44314, n44315,
         n44316, n44317, n44318, n44319, n44320, n44321, n44322, n44323,
         n44324, n44325, n44326, n44327, n44328, n44329, n44330, n44331,
         n44332, n44333, n44334, n44335, n44336, n44337, n44338, n44339,
         n44340, n44341, n44342, n44343, n44344, n44345, n44346, n44347,
         n44348, n44349, n44350, n44351, n44352, n44353, n44354, n44355,
         n44356, n44357, n44358, n44359, n44360, n44361, n44362, n44363,
         n44364, n44365, n44366, n44367, n44368, n44369, n44370, n44371,
         n44372, n44373, n44374, n44375, n44376, n44377, n44378, n44379,
         n44380, n44381, n44382, n44383, n44384, n44385, n44386, n44387,
         n44388, n44389, n44390, n44391, n44392, n44393, n44394, n44395,
         n44396, n44397, n44398, n44399, n44400, n44401, n44402, n44403,
         n44404, n44405, n44406, n44407, n44408, n44409, n44410, n44411,
         n44412, n44413, n44414, n44415, n44416, n44417, n44418, n44419,
         n44420, n44421, n44422, n44423, n44424, n44425, n44426, n44427,
         n44428, n44429, n44430, n44431, n44432, n44433, n44434, n44435,
         n44436, n44437, n44438, n44439, n44440, n44441, n44442, n44443,
         n44444, n44445, n44446, n44447, n44448, n44449, n44450, n44451,
         n44452, n44453, n44454, n44455, n44456, n44457, n44458, n44459,
         n44460, n44461, n44462, n44463, n44464, n44465, n44466, n44467,
         n44468, n44469, n44470, n44471, n44472, n44473, n44474, n44475,
         n44476, n44477, n44478, n44479, n44480, n44481, n44482, n44483,
         n44484, n44485, n44486, n44487, n44488, n44489, n44490, n44491,
         n44492, n44493, n44494, n44495, n44496, n44497, n44498, n44499,
         n44500, n44501, n44502, n44503, n44504, n44505, n44506, n44507,
         n44508, n44509, n44510, n44511, n44512, n44513, n44514, n44515,
         n44516, n44517, n44518, n44519, n44520, n44521, n44522, n44523,
         n44524, n44525, n44526, n44527, n44528, n44529, n44530, n44531,
         n44532, n44533, n44534, n44535, n44536, n44537, n44538, n44539,
         n44540, n44541, n44542, n44543, n44544, n44545, n44546, n44547,
         n44548, n44549, n44550, n44551, n44552, n44553, n44554, n44555,
         n44556, n44557, n44558, n44559, n44560, n44561, n44562, n44563,
         n44564, n44565, n44566, n44567, n44568, n44569, n44570, n44571,
         n44572, n44573, n44574, n44575, n44576, n44577, n44578, n44579,
         n44580, n44581, n44582, n44583, n44584, n44585, n44586, n44587,
         n44588, n44589, n44590, n44591, n44592, n44593, n44594, n44595,
         n44596, n44597, n44598, n44599, n44600, n44601, n44602, n44603,
         n44604, n44605, n44606, n44607, n44608, n44609, n44610, n44611,
         n44612, n44613, n44614, n44615, n44616, n44617, n44618, n44619,
         n44620, n44621, n44622, n44623, n44624, n44625, n44626, n44627,
         n44628, n44629, n44630, n44631, n44632, n44633, n44634, n44635,
         n44636, n44637, n44638, n44639, n44640, n44641, n44642, n44643,
         n44644, n44645, n44646, n44647, n44648, n44649, n44650, n44651,
         n44652, n44653, n44654, n44655, n44656, n44657, n44658, n44659,
         n44660, n44661, n44662, n44663, n44664, n44665, n44666, n44667,
         n44668, n44669, n44670, n44671, n44672, n44673, n44674, n44675,
         n44676, n44677, n44678, n44679, n44680, n44681, n44682, n44683,
         n44684, n44685, n44686, n44687, n44688, n44689, n44690, n44691,
         n44692, n44693, n44694, n44695, n44696, n44697, n44698, n44699,
         n44700, n44701, n44702, n44703, n44704, n44705, n44706, n44707,
         n44708, n44709, n44710, n44711, n44712, n44713, n44714, n44715,
         n44716, n44717, n44718, n44719, n44720, n44721, n44722, n44723,
         n44724, n44725, n44726, n44727, n44728, n44729, n44730, n44731,
         n44732, n44733, n44734, n44735, n44736, n44737, n44738, n44739,
         n44740, n44741, n44742, n44743, n44744, n44745, n44746, n44747,
         n44748, n44749, n44750, n44751, n44752, n44753, n44754, n44755,
         n44756, n44757, n44758, n44759, n44760, n44761, n44762, n44763,
         n44764, n44765, n44766, n44767, n44768, n44769, n44770, n44771,
         n44772, n44773, n44774, n44775, n44776, n44777, n44778, n44779,
         n44780, n44781, n44782, n44783, n44784, n44785, n44786, n44787,
         n44788, n44789, n44790, n44791, n44792, n44793, n44794, n44795,
         n44796, n44797, n44798, n44799, n44800, n44801, n44802, n44803,
         n44804, n44805, n44806, n44807, n44808, n44809, n44810, n44811,
         n44812, n44813, n44814, n44815, n44816, n44817, n44818, n44819,
         n44820, n44821, n44822, n44823, n44824, n44825, n44826, n44827,
         n44828, n44829, n44830, n44831, n44832, n44833, n44834, n44835,
         n44836, n44837, n44838, n44839, n44840, n44841, n44842, n44843,
         n44844, n44845, n44846, n44847, n44848, n44849, n44850, n44851,
         n44852, n44853, n44854, n44855, n44856, n44857, n44858, n44859,
         n44860, n44861, n44862, n44863, n44864, n44865, n44866, n44867,
         n44868, n44869, n44870, n44871, n44872, n44873, n44874, n44875,
         n44876, n44877, n44878, n44879, n44880, n44881, n44882, n44883,
         n44884, n44885, n44886, n44887, n44888, n44889, n44890, n44891,
         n44892, n44893, n44894, n44895, n44896, n44897, n44898, n44899,
         n44900, n44901, n44902, n44903, n44904, n44905, n44906, n44907,
         n44908, n44909, n44910, n44911, n44912, n44913, n44914, n44915,
         n44916, n44917, n44918, n44919, n44920, n44921, n44922, n44923,
         n44924, n44925, n44926, n44927, n44928, n44929, n44930, n44931,
         n44932, n44933, n44934, n44935, n44936, n44937, n44938, n44939,
         n44940, n44941, n44942, n44943, n44944, n44945, n44946, n44947,
         n44948, n44949, n44950, n44951, n44952, n44953, n44954, n44955,
         n44956, n44957, n44958, n44959, n44960, n44961, n44962, n44963,
         n44964, n44965, n44966, n44967, n44968, n44969, n44970, n44971,
         n44972, n44973, n44974, n44975, n44976, n44977, n44978, n44979,
         n44980, n44981, n44982, n44983, n44984, n44985, n44986, n44987,
         n44988, n44989, n44990, n44991, n44992, n44993, n44994, n44995,
         n44996, n44997, n44998, n44999, n45000, n45001, n45002, n45003,
         n45004, n45005, n45006, n45007, n45008, n45009, n45010, n45011,
         n45012, n45013, n45014, n45015, n45016, n45017, n45018, n45019,
         n45020, n45021, n45022, n45023, n45024, n45025, n45026, n45027,
         n45028, n45029, n45030, n45031, n45032, n45033, n45034, n45035,
         n45036, n45037, n45038, n45039, n45040, n45041, n45042, n45043,
         n45044, n45045, n45046, n45047, n45048, n45049, n45050, n45051,
         n45052, n45053, n45054, n45055, n45056, n45057, n45058, n45059,
         n45060, n45061, n45062, n45063, n45064, n45065, n45066, n45067,
         n45068, n45069, n45070, n45071, n45072, n45073, n45074, n45075,
         n45076, n45077, n45078, n45079, n45080, n45081, n45082, n45083,
         n45084, n45085, n45086, n45087, n45088, n45089, n45090, n45091,
         n45092, n45093, n45094, n45095, n45096, n45097, n45098, n45099,
         n45100, n45101, n45102, n45103, n45104, n45105, n45106, n45107,
         n45108, n45109, n45110, n45111, n45112, n45113, n45114, n45115,
         n45116, n45117, n45118, n45119, n45120, n45121, n45122, n45123,
         n45124, n45125, n45126, n45127, n45128, n45129, n45130, n45131,
         n45132, n45133, n45134, n45135, n45136, n45137, n45138, n45139,
         n45140, n45141, n45142, n45143, n45144, n45145, n45146, n45147,
         n45148, n45149, n45150, n45151, n45152, n45153, n45154, n45155,
         n45156, n45157, n45158, n45159, n45160, n45161, n45162, n45163,
         n45164, n45165, n45166, n45167, n45168, n45169, n45170, n45171,
         n45172, n45173, n45174, n45175, n45176, n45177, n45178, n45179,
         n45180, n45181, n45182, n45183, n45184, n45185, n45186, n45187,
         n45188, n45189, n45190, n45191, n45192, n45193, n45194, n45195,
         n45196, n45197, n45198, n45199, n45200, n45201, n45202, n45203,
         n45204, n45205, n45206, n45207, n45208, n45209, n45210, n45211,
         n45212, n45213, n45214, n45215, n45216, n45217, n45218, n45219,
         n45220, n45221, n45222, n45223, n45224, n45225, n45226, n45227,
         n45228, n45229, n45230, n45231, n45232, n45233, n45234, n45235,
         n45236, n45237, n45238, n45239, n45240, n45241, n45242, n45243,
         n45244, n45245, n45246, n45247, n45248, n45249, n45250, n45251,
         n45252, n45253, n45254, n45255, n45256, n45257, n45258, n45259,
         n45260, n45261, n45262, n45263, n45264, n45265, n45266, n45267,
         n45268, n45269, n45270, n45271, n45272, n45273, n45274, n45275,
         n45276, n45277, n45278, n45279, n45280, n45281, n45282, n45283,
         n45284, n45285, n45286, n45287, n45288, n45289, n45290, n45291,
         n45292, n45293, n45294, n45295, n45296, n45297, n45298, n45299,
         n45300, n45301, n45302, n45303, n45304, n45305, n45306, n45307,
         n45308, n45309, n45310, n45311, n45312, n45313, n45314, n45315,
         n45316, n45317, n45318, n45319, n45320, n45321, n45322, n45323,
         n45324, n45325, n45326, n45327, n45328, n45329, n45330, n45331,
         n45332, n45333, n45334, n45335, n45336, n45337, n45338, n45339,
         n45340, n45341, n45342, n45343, n45344, n45345, n45346, n45347,
         n45348, n45349, n45350, n45351, n45352, n45353, n45354, n45355,
         n45356, n45357, n45358, n45359, n45360, n45361, n45362, n45363,
         n45364, n45365, n45366, n45367, n45368, n45369, n45370, n45371,
         n45372, n45373, n45374, n45375, n45376, n45377, n45378, n45379,
         n45380, n45381, n45382, n45383, n45384, n45385, n45386, n45387,
         n45388, n45389, n45390, n45391, n45392, n45393, n45394, n45395,
         n45396, n45397, n45398, n45399, n45400, n45401, n45402, n45403,
         n45404, n45405, n45406, n45407, n45408, n45409, n45410, n45411,
         n45412, n45413, n45414, n45415, n45416, n45417, n45418, n45419,
         n45420, n45421, n45422, n45423, n45424, n45425, n45426, n45427,
         n45428, n45429, n45430, n45431, n45432, n45433, n45434, n45435,
         n45436, n45437, n45438, n45439, n45440, n45441, n45442, n45443,
         n45444, n45445, n45446, n45447, n45448, n45449, n45450, n45451,
         n45452, n45453, n45454, n45455, n45456, n45457, n45458, n45459,
         n45460, n45461, n45462, n45463, n45464, n45465, n45466, n45467,
         n45468, n45469, n45470, n45471, n45472, n45473, n45474, n45475,
         n45476, n45477, n45478, n45479, n45480, n45481, n45482, n45483,
         n45484, n45485, n45486, n45487, n45488, n45489, n45490, n45491,
         n45492, n45493, n45494, n45495, n45496, n45497, n45498, n45499,
         n45500, n45501, n45502, n45503, n45504, n45505, n45506, n45507,
         n45508, n45509, n45510, n45511, n45512, n45513, n45514, n45515,
         n45516, n45517, n45518, n45519, n45520, n45521, n45522, n45523,
         n45524, n45525, n45526, n45527, n45528, n45529, n45530, n45531,
         n45532, n45533, n45534, n45535, n45536, n45537, n45538, n45539,
         n45540, n45541, n45542, n45543, n45544, n45545, n45546, n45547,
         n45548, n45549, n45550, n45551, n45552, n45553, n45554, n45555,
         n45556, n45557, n45558, n45559, n45560, n45561, n45562, n45563,
         n45564, n45565, n45566, n45567, n45568, n45569, n45570, n45571,
         n45572, n45573, n45574, n45575, n45576, n45577, n45578, n45579,
         n45580, n45581, n45582, n45583, n45584, n45585, n45586, n45587,
         n45588, n45589, n45590, n45591, n45592, n45593, n45594, n45595,
         n45596, n45597, n45598, n45599, n45600, n45601, n45602, n45603,
         n45604, n45605, n45606, n45607, n45608, n45609, n45610, n45611,
         n45612, n45613, n45614, n45615, n45616, n45617, n45618, n45619,
         n45620, n45621, n45622, n45623, n45624, n45625, n45626, n45627,
         n45628, n45629, n45630, n45631, n45632, n45633, n45634, n45635,
         n45636, n45637, n45638, n45639, n45640, n45641, n45642, n45643,
         n45644, n45645, n45646, n45647, n45648, n45649, n45650, n45651,
         n45652, n45653, n45654, n45655, n45656, n45657, n45658, n45659,
         n45660, n45661, n45662, n45663, n45664, n45665, n45666, n45667,
         n45668, n45669, n45670, n45671, n45672, n45673, n45674, n45675,
         n45676, n45677, n45678, n45679, n45680, n45681, n45682, n45683,
         n45684, n45685, n45686, n45687, n45688, n45689, n45690, n45691,
         n45692, n45693, n45694, n45695, n45696, n45697, n45698, n45699,
         n45700, n45701, n45702, n45703, n45704, n45705, n45706, n45707,
         n45708, n45709, n45710, n45711, n45712, n45713, n45714, n45715,
         n45716, n45717, n45718, n45719, n45720, n45721, n45722, n45723,
         n45724, n45725, n45726, n45727, n45728, n45729, n45730, n45731,
         n45732, n45733, n45734, n45735, n45736, n45737, n45738, n45739,
         n45740, n45741, n45742, n45743, n45744, n45745, n45746, n45747,
         n45748, n45749, n45750, n45751, n45752, n45753, n45754, n45755,
         n45756, n45757, n45758, n45759, n45760, n45761, n45762, n45763,
         n45764, n45765, n45766, n45767, n45768, n45769, n45770, n45771,
         n45772, n45773, n45774, n45775, n45776, n45777, n45778, n45779,
         n45780, n45781, n45782, n45783, n45784, n45785, n45786, n45787,
         n45788, n45789, n45790, n45791, n45792, n45793, n45794, n45795,
         n45796, n45797, n45798, n45799, n45800, n45801, n45802, n45803,
         n45804, n45805, n45806, n45807, n45808, n45809, n45810, n45811,
         n45812, n45813, n45814, n45815, n45816, n45817, n45818, n45819,
         n45820, n45821, n45822, n45823, n45824, n45825, n45826, n45827,
         n45828, n45829, n45830, n45831, n45832, n45833, n45834, n45835,
         n45836, n45837, n45838, n45839, n45840, n45841, n45842, n45843,
         n45844, n45845, n45846, n45847, n45848, n45849, n45850, n45851,
         n45852, n45853, n45854, n45855, n45856, n45857, n45858, n45859,
         n45860, n45861, n45862, n45863, n45864, n45865, n45866, n45867,
         n45868, n45869, n45870, n45871, n45872, n45873, n45874, n45875,
         n45876, n45877, n45878, n45879, n45880, n45881, n45882, n45883,
         n45884, n45885, n45886, n45887, n45888, n45889, n45890, n45891,
         n45892, n45893, n45894, n45895, n45896, n45897, n45898, n45899,
         n45900, n45901, n45902, n45903, n45904, n45905, n45906, n45907,
         n45908, n45909, n45910, n45911, n45912, n45913, n45914, n45915,
         n45916, n45917, n45918, n45919, n45920, n45921, n45922, n45923,
         n45924, n45925, n45926, n45927, n45928, n45929, n45930, n45931,
         n45932, n45933, n45934, n45935, n45936, n45937, n45938, n45939,
         n45940, n45941, n45942, n45943, n45944, n45945, n45946, n45947,
         n45948, n45949, n45950, n45951, n45952, n45953, n45954, n45955,
         n45956, n45957, n45958, n45959, n45960, n45961, n45962, n45963,
         n45964, n45965, n45966, n45967, n45968, n45969, n45970, n45971,
         n45972, n45973, n45974, n45975, n45976, n45977, n45978, n45979,
         n45980, n45981, n45982, n45983, n45984, n45985, n45986, n45987,
         n45988, n45989, n45990, n45991, n45992, n45993, n45994, n45995,
         n45996, n45997, n45998, n45999, n46000, n46001, n46002, n46003,
         n46004, n46005, n46006, n46007, n46008, n46009, n46010, n46011,
         n46012, n46013, n46014, n46015, n46016, n46017, n46018, n46019,
         n46020, n46021, n46022, n46023, n46024, n46025, n46026, n46027,
         n46028, n46029, n46030, n46031, n46032, n46033, n46034, n46035,
         n46036, n46037, n46038, n46039, n46040, n46041, n46042, n46043,
         n46044, n46045, n46046, n46047, n46048, n46049, n46050, n46051,
         n46052, n46053, n46054, n46055, n46056, n46057, n46058, n46059,
         n46060, n46061, n46062, n46063, n46064, n46065, n46066, n46067,
         n46068, n46069, n46070, n46071, n46072, n46073, n46074, n46075,
         n46076, n46077, n46078, n46079, n46080, n46081, n46082, n46083,
         n46084, n46085, n46086, n46087, n46088, n46089, n46090, n46091,
         n46092, n46093, n46094, n46095, n46096, n46097, n46098, n46099,
         n46100, n46101, n46102, n46103, n46104, n46105, n46106, n46107,
         n46108, n46109, n46110, n46111, n46112, n46113, n46114, n46115,
         n46116, n46117, n46118, n46119, n46120, n46121, n46122, n46123,
         n46124, n46125, n46126, n46127, n46128, n46129, n46130, n46131,
         n46132, n46133, n46134, n46135, n46136, n46137, n46138, n46139,
         n46140, n46141, n46142, n46143, n46144, n46145, n46146, n46147,
         n46148, n46149, n46150, n46151, n46152, n46153, n46154, n46155,
         n46156, n46157, n46158, n46159, n46160, n46161, n46162, n46163,
         n46164, n46165, n46166, n46167, n46168, n46169, n46170, n46171,
         n46172, n46173, n46174, n46175, n46176, n46177, n46178, n46179,
         n46180, n46181, n46182, n46183, n46184, n46185, n46186, n46187,
         n46188, n46189, n46190, n46191, n46192, n46193, n46194, n46195,
         n46196, n46197, n46198, n46199, n46200, n46201, n46202, n46203,
         n46204, n46205, n46206, n46207, n46208, n46209, n46210, n46211,
         n46212, n46213, n46214, n46215, n46216, n46217, n46218, n46219,
         n46220, n46221, n46222, n46223, n46224, n46225, n46226, n46227,
         n46228, n46229, n46230, n46231, n46232, n46233, n46234, n46235,
         n46236, n46237, n46238, n46239, n46240, n46241, n46242, n46243,
         n46244, n46245, n46246, n46247, n46248, n46249, n46250, n46251,
         n46252, n46253, n46254, n46255, n46256, n46257, n46258, n46259,
         n46260, n46261, n46262, n46263, n46264, n46265, n46266, n46267,
         n46268, n46269, n46270, n46271, n46272, n46273, n46274, n46275,
         n46276, n46277, n46278, n46279, n46280, n46281, n46282, n46283,
         n46284, n46285, n46286, n46287, n46288, n46289, n46290, n46291,
         n46292, n46293, n46294, n46295, n46296, n46297, n46298, n46299,
         n46300, n46301, n46302, n46303, n46304, n46305, n46306, n46307,
         n46308, n46309, n46310, n46311, n46312, n46313, n46314, n46315,
         n46316, n46317, n46318, n46319, n46320, n46321, n46322, n46323,
         n46324, n46325, n46326, n46327, n46328, n46329, n46330, n46331,
         n46332, n46333, n46334, n46335, n46336, n46337, n46338, n46339,
         n46340, n46341, n46342, n46343, n46344, n46345, n46346, n46347,
         n46348, n46349, n46350, n46351, n46352, n46353, n46354, n46355,
         n46356, n46357, n46358, n46359, n46360, n46361, n46362, n46363,
         n46364, n46365, n46366, n46367, n46368, n46369, n46370, n46371,
         n46372, n46373, n46374, n46375, n46376, n46377, n46378, n46379,
         n46380, n46381, n46382, n46383, n46384, n46385, n46386, n46387,
         n46388, n46389, n46390, n46391, n46392, n46393, n46394, n46395,
         n46396, n46397, n46398, n46399, n46400, n46401, n46402, n46403,
         n46404, n46405, n46406, n46407, n46408, n46409, n46410, n46411,
         n46412, n46413, n46414, n46415, n46416, n46417, n46418, n46419,
         n46420, n46421, n46422, n46423, n46424, n46425, n46426, n46427,
         n46428, n46429, n46430, n46431, n46432, n46433, n46434, n46435,
         n46436, n46437, n46438, n46439, n46440, n46441, n46442, n46443,
         n46444, n46445, n46446, n46447, n46448, n46449, n46450, n46451,
         n46452, n46453, n46454, n46455, n46456, n46457, n46458, n46459,
         n46460, n46461, n46462, n46463, n46464, n46465, n46466, n46467,
         n46468, n46469, n46470, n46471, n46472, n46473, n46474, n46475,
         n46476, n46477, n46478, n46479, n46480, n46481, n46482, n46483,
         n46484, n46485, n46486, n46487, n46488, n46489, n46490, n46491,
         n46492, n46493, n46494, n46495, n46496, n46497, n46498, n46499,
         n46500, n46501, n46502, n46503, n46504, n46505, n46506, n46507,
         n46508, n46509, n46510, n46511, n46512, n46513, n46514, n46515,
         n46516, n46517, n46518, n46519, n46520, n46521, n46522, n46523,
         n46524, n46525, n46526, n46527, n46528, n46529, n46530, n46531,
         n46532, n46533, n46534, n46535, n46536, n46537, n46538, n46539,
         n46540, n46541, n46542, n46543, n46544, n46545, n46546, n46547,
         n46548, n46549, n46550, n46551, n46552, n46553, n46554, n46555,
         n46556, n46557, n46558, n46559, n46560, n46561, n46562, n46563,
         n46564, n46565, n46566, n46567, n46568, n46569, n46570, n46571,
         n46572, n46573, n46574, n46575, n46576, n46577, n46578, n46579,
         n46580, n46581, n46582, n46583, n46584, n46585, n46586, n46587,
         n46588, n46589, n46590, n46591, n46592, n46593, n46594, n46595,
         n46596, n46597, n46598, n46599, n46600, n46601, n46602, n46603,
         n46604, n46605, n46606, n46607, n46608, n46609, n46610, n46611,
         n46612, n46613, n46614, n46615, n46616, n46617, n46618, n46619,
         n46620, n46621, n46622, n46623, n46624, n46625, n46626, n46627,
         n46628, n46629, n46630, n46631, n46632, n46633, n46634, n46635,
         n46636, n46637, n46638, n46639, n46640, n46641, n46642, n46643,
         n46644, n46645, n46646, n46647, n46648, n46649, n46650, n46651,
         n46652, n46653, n46654, n46655, n46656, n46657, n46658, n46659,
         n46660, n46661, n46662, n46663, n46664, n46665, n46666, n46667,
         n46668, n46669, n46670, n46671, n46672, n46673, n46674, n46675,
         n46676, n46677, n46678, n46679, n46680, n46681, n46682, n46683,
         n46684, n46685, n46686, n46687, n46688, n46689, n46690, n46691,
         n46692, n46693, n46694, n46695, n46696, n46697, n46698, n46699,
         n46700, n46701, n46702, n46703, n46704, n46705, n46706, n46707,
         n46708, n46709, n46710, n46711, n46712, n46713, n46714, n46715,
         n46716, n46717, n46718, n46719, n46720, n46721, n46722, n46723,
         n46724, n46725, n46726, n46727, n46728, n46729, n46730, n46731,
         n46732, n46733, n46734, n46735, n46736, n46737, n46738, n46739,
         n46740, n46741, n46742, n46743, n46744, n46745, n46746, n46747,
         n46748, n46749, n46750, n46751, n46752, n46753, n46754, n46755,
         n46756, n46757, n46758, n46759, n46760, n46761, n46762, n46763,
         n46764, n46765, n46766, n46767, n46768, n46769, n46770, n46771,
         n46772, n46773, n46774, n46775, n46776, n46777, n46778, n46779,
         n46780, n46781, n46782, n46783, n46784, n46785, n46786, n46787,
         n46788, n46789, n46790, n46791, n46792, n46793, n46794, n46795,
         n46796, n46797, n46798, n46799, n46800, n46801, n46802, n46803,
         n46804, n46805, n46806, n46807, n46808, n46809, n46810, n46811,
         n46812, n46813, n46814, n46815, n46816, n46817, n46818, n46819,
         n46820, n46821, n46822, n46823, n46824, n46825, n46826, n46827,
         n46828, n46829, n46830, n46831, n46832, n46833, n46834, n46835,
         n46836, n46837, n46838, n46839, n46840, n46841, n46842, n46843,
         n46844, n46845, n46846, n46847, n46848, n46849, n46850, n46851,
         n46852, n46853, n46854, n46855, n46856, n46857, n46858, n46859,
         n46860, n46861, n46862, n46863, n46864, n46865, n46866, n46867,
         n46868, n46869, n46870, n46871, n46872, n46873, n46874, n46875,
         n46876, n46877, n46878, n46879, n46880, n46881, n46882, n46883,
         n46884, n46885, n46886, n46887, n46888, n46889, n46890, n46891,
         n46892, n46893, n46894, n46895, n46896, n46897, n46898, n46899,
         n46900, n46901, n46902, n46903, n46904, n46905, n46906, n46907,
         n46908, n46909, n46910, n46911, n46912, n46913, n46914, n46915,
         n46916, n46917, n46918, n46919, n46920, n46921, n46922, n46923,
         n46924, n46925, n46926, n46927, n46928, n46929, n46930, n46931,
         n46932, n46933, n46934, n46935, n46936, n46937, n46938, n46939,
         n46940, n46941, n46942, n46943, n46944, n46945, n46946, n46947,
         n46948, n46949, n46950, n46951, n46952, n46953, n46954, n46955,
         n46956, n46957, n46958, n46959, n46960, n46961, n46962, n46963,
         n46964, n46965, n46966, n46967, n46968, n46969, n46970, n46971,
         n46972, n46973, n46974, n46975, n46976, n46977, n46978, n46979,
         n46980, n46981, n46982, n46983, n46984, n46985, n46986, n46987,
         n46988, n46989, n46990, n46991, n46992, n46993, n46994, n46995,
         n46996, n46997, n46998, n46999, n47000, n47001, n47002, n47003,
         n47004, n47005, n47006, n47007, n47008, n47009, n47010, n47011,
         n47012, n47013, n47014, n47015, n47016, n47017, n47018, n47019,
         n47020, n47021, n47022, n47023, n47024, n47025, n47026, n47027,
         n47028, n47029, n47030, n47031, n47032, n47033, n47034, n47035,
         n47036, n47037, n47038, n47039, n47040, n47041, n47042, n47043,
         n47044, n47045, n47046, n47047, n47048, n47049, n47050, n47051,
         n47052, n47053, n47054, n47055, n47056, n47057, n47058, n47059,
         n47060, n47061, n47062, n47063, n47064, n47065, n47066, n47067,
         n47068, n47069, n47070, n47071, n47072, n47073, n47074, n47075,
         n47076, n47077, n47078, n47079, n47080, n47081, n47082, n47083,
         n47084, n47085, n47086, n47087, n47088, n47089, n47090, n47091,
         n47092, n47093, n47094, n47095, n47096, n47097, n47098, n47099,
         n47100, n47101, n47102, n47103, n47104, n47105, n47106, n47107,
         n47108, n47109, n47110, n47111, n47112, n47113, n47114, n47115,
         n47116, n47117, n47118, n47119, n47120, n47121, n47122, n47123,
         n47124, n47125, n47126, n47127, n47128, n47129, n47130, n47131,
         n47132, n47133, n47134, n47135, n47136, n47137, n47138, n47139,
         n47140, n47141, n47142, n47143, n47144, n47145, n47146, n47147,
         n47148, n47149, n47150, n47151, n47152, n47153, n47154, n47155,
         n47156, n47157, n47158, n47159, n47160, n47161, n47162, n47163,
         n47164, n47165, n47166, n47167, n47168, n47169, n47170, n47171,
         n47172, n47173, n47174, n47175, n47176, n47177, n47178, n47179,
         n47180, n47181, n47182, n47183, n47184, n47185, n47186, n47187,
         n47188, n47189, n47190, n47191, n47192, n47193, n47194, n47195,
         n47196, n47197, n47198, n47199, n47200, n47201, n47202, n47203,
         n47204, n47205, n47206, n47207, n47208, n47209, n47210, n47211,
         n47212, n47213, n47214, n47215, n47216, n47217, n47218, n47219,
         n47220, n47221, n47222, n47223, n47224, n47225, n47226, n47227,
         n47228, n47229, n47230, n47231, n47232, n47233, n47234, n47235,
         n47236, n47237, n47238, n47239, n47240, n47241, n47242, n47243,
         n47244, n47245, n47246, n47247, n47248, n47249, n47250, n47251,
         n47252, n47253, n47254, n47255, n47256, n47257, n47258, n47259,
         n47260, n47261, n47262, n47263, n47264, n47265, n47266, n47267,
         n47268, n47269, n47270, n47271, n47272, n47273, n47274, n47275,
         n47276, n47277, n47278, n47279, n47280, n47281, n47282, n47283,
         n47284, n47285, n47286, n47287, n47288, n47289, n47290, n47291,
         n47292, n47293, n47294, n47295, n47296, n47297, n47298, n47299,
         n47300, n47301, n47302, n47303, n47304, n47305, n47306, n47307,
         n47308, n47309, n47310, n47311, n47312, n47313, n47314, n47315,
         n47316, n47317, n47318, n47319, n47320, n47321, n47322, n47323,
         n47324, n47325, n47326, n47327, n47328, n47329, n47330, n47331,
         n47332, n47333, n47334, n47335, n47336, n47337, n47338, n47339,
         n47340, n47341, n47342, n47343, n47344, n47345, n47346, n47347,
         n47348, n47349, n47350, n47351, n47352, n47353, n47354, n47355,
         n47356, n47357, n47358, n47359, n47360, n47361, n47362, n47363,
         n47364, n47365, n47366, n47367, n47368, n47369, n47370, n47371,
         n47372, n47373, n47374, n47375, n47376, n47377, n47378, n47379,
         n47380, n47381, n47382, n47383, n47384, n47385, n47386, n47387,
         n47388, n47389, n47390, n47391, n47392, n47393, n47394, n47395,
         n47396, n47397, n47398, n47399, n47400, n47401, n47402, n47403,
         n47404, n47405, n47406, n47407, n47408, n47409, n47410, n47411,
         n47412, n47413, n47414, n47415, n47416, n47417, n47418, n47419,
         n47420, n47421, n47422, n47423, n47424, n47425, n47426, n47427,
         n47428, n47429, n47430, n47431, n47432, n47433, n47434, n47435,
         n47436, n47437, n47438, n47439, n47440, n47441, n47442, n47443,
         n47444, n47445, n47446, n47447, n47448, n47449, n47450, n47451,
         n47452, n47453, n47454, n47455, n47456, n47457, n47458, n47459,
         n47460, n47461, n47462, n47463, n47464, n47465, n47466, n47467,
         n47468, n47469, n47470, n47471, n47472, n47473, n47474, n47475,
         n47476, n47477, n47478, n47479, n47480, n47481, n47482, n47483,
         n47484, n47485, n47486, n47487, n47488, n47489, n47490, n47491,
         n47492, n47493, n47494, n47495, n47496, n47497, n47498, n47499,
         n47500, n47501, n47502, n47503, n47504, n47505, n47506, n47507,
         n47508, n47509, n47510, n47511, n47512, n47513, n47514, n47515,
         n47516, n47517, n47518, n47519, n47520, n47521, n47522, n47523,
         n47524, n47525, n47526, n47527, n47528, n47529, n47530, n47531,
         n47532, n47533, n47534, n47535, n47536, n47537, n47538, n47539,
         n47540, n47541, n47542, n47543, n47544, n47545, n47546, n47547,
         n47548, n47549, n47550, n47551, n47552, n47553, n47554, n47555,
         n47556, n47557, n47558, n47559, n47560, n47561, n47562, n47563,
         n47564, n47565, n47566, n47567, n47568, n47569, n47570, n47571,
         n47572, n47573, n47574, n47575, n47576, n47577, n47578, n47579,
         n47580, n47581, n47582, n47583, n47584, n47585, n47586, n47587,
         n47588, n47589, n47590, n47591, n47592, n47593, n47594, n47595,
         n47596, n47597, n47598, n47599, n47600, n47601, n47602, n47603,
         n47604, n47605, n47606, n47607, n47608, n47609, n47610, n47611,
         n47612, n47613, n47614, n47615, n47616, n47617, n47618, n47619,
         n47620, n47621, n47622, n47623, n47624, n47625, n47626, n47627,
         n47628, n47629, n47630, n47631, n47632, n47633, n47634, n47635,
         n47636, n47637, n47638, n47639, n47640, n47641, n47642, n47643,
         n47644, n47645, n47646, n47647, n47648, n47649, n47650, n47651,
         n47652, n47653, n47654, n47655, n47656, n47657, n47658, n47659,
         n47660, n47661, n47662, n47663, n47664, n47665, n47666, n47667,
         n47668, n47669, n47670, n47671, n47672, n47673, n47674, n47675,
         n47676, n47677, n47678, n47679, n47680, n47681, n47682, n47683,
         n47684, n47685, n47686, n47687, n47688, n47689, n47690, n47691,
         n47692, n47693, n47694, n47695, n47696, n47697, n47698, n47699,
         n47700, n47701, n47702, n47703, n47704, n47705, n47706, n47707,
         n47708, n47709, n47710, n47711, n47712, n47713, n47714, n47715,
         n47716, n47717, n47718, n47719, n47720, n47721, n47722, n47723,
         n47724, n47725, n47726, n47727, n47728, n47729, n47730, n47731,
         n47732, n47733, n47734, n47735, n47736, n47737, n47738, n47739,
         n47740, n47741, n47742, n47743, n47744, n47745, n47746, n47747,
         n47748, n47749, n47750, n47751, n47752, n47753, n47754, n47755,
         n47756, n47757, n47758, n47759, n47760, n47761, n47762, n47763,
         n47764, n47765, n47766, n47767, n47768, n47769, n47770, n47771,
         n47772, n47773, n47774, n47775, n47776, n47777, n47778, n47779,
         n47780, n47781, n47782, n47783, n47784, n47785, n47786, n47787,
         n47788, n47789, n47790, n47791, n47792, n47793, n47794, n47795,
         n47796, n47797, n47798, n47799, n47800, n47801, n47802, n47803,
         n47804, n47805, n47806, n47807, n47808, n47809, n47810, n47811,
         n47812, n47813, n47814, n47815, n47816, n47817, n47818, n47819,
         n47820, n47821, n47822, n47823, n47824, n47825, n47826, n47827,
         n47828, n47829, n47830, n47831, n47832, n47833, n47834, n47835,
         n47836, n47837, n47838, n47839, n47840, n47841, n47842, n47843,
         n47844, n47845, n47846, n47847, n47848, n47849, n47850, n47851,
         n47852, n47853, n47854, n47855, n47856, n47857, n47858, n47859,
         n47860, n47861, n47862, n47863, n47864, n47865, n47866, n47867,
         n47868, n47869, n47870, n47871, n47872, n47873, n47874, n47875,
         n47876, n47877, n47878, n47879, n47880, n47881, n47882, n47883,
         n47884, n47885, n47886, n47887, n47888, n47889, n47890, n47891,
         n47892, n47893, n47894, n47895, n47896, n47897, n47898, n47899,
         n47900, n47901, n47902, n47903, n47904, n47905, n47906, n47907,
         n47908, n47909, n47910, n47911, n47912, n47913, n47914, n47915,
         n47916, n47917, n47918, n47919, n47920, n47921, n47922, n47923,
         n47924, n47925, n47926, n47927, n47928, n47929, n47930, n47931,
         n47932, n47933, n47934, n47935, n47936, n47937, n47938, n47939,
         n47940, n47941, n47942, n47943, n47944, n47945, n47946, n47947,
         n47948, n47949, n47950, n47951, n47952, n47953, n47954, n47955,
         n47956, n47957, n47958, n47959, n47960, n47961, n47962, n47963,
         n47964, n47965, n47966, n47967, n47968, n47969, n47970, n47971,
         n47972, n47973, n47974, n47975, n47976, n47977, n47978, n47979,
         n47980, n47981, n47982, n47983, n47984, n47985, n47986, n47987,
         n47988, n47989, n47990, n47991, n47992, n47993, n47994, n47995,
         n47996, n47997, n47998, n47999, n48000, n48001, n48002, n48003,
         n48004, n48005, n48006, n48007, n48008, n48009, n48010, n48011,
         n48012, n48013, n48014, n48015, n48016, n48017, n48018, n48019,
         n48020, n48021, n48022, n48023, n48024, n48025, n48026, n48027,
         n48028, n48029, n48030, n48031, n48032, n48033, n48034, n48035,
         n48036, n48037, n48038, n48039, n48040, n48041, n48042, n48043,
         n48044, n48045, n48046, n48047, n48048, n48049, n48050, n48051,
         n48052, n48053, n48054, n48055, n48056, n48057, n48058, n48059,
         n48060, n48061, n48062, n48063, n48064, n48065, n48066, n48067,
         n48068, n48069, n48070, n48071, n48072, n48073, n48074, n48075,
         n48076, n48077, n48078, n48079, n48080, n48081, n48082, n48083,
         n48084, n48085, n48086, n48087, n48088, n48089, n48090, n48091,
         n48092, n48093, n48094, n48095, n48096, n48097, n48098, n48099,
         n48100, n48101, n48102, n48103, n48104, n48105, n48106, n48107,
         n48108, n48109, n48110, n48111, n48112, n48113, n48114, n48115,
         n48116, n48117, n48118, n48119, n48120, n48121, n48122, n48123,
         n48124, n48125, n48126, n48127, n48128, n48129, n48130, n48131,
         n48132, n48133, n48134, n48135, n48136, n48137, n48138, n48139,
         n48140, n48141, n48142, n48143, n48144, n48145, n48146, n48147,
         n48148, n48149, n48150, n48151, n48152, n48153, n48154, n48155,
         n48156, n48157, n48158, n48159, n48160, n48161, n48162, n48163,
         n48164, n48165, n48166, n48167, n48168, n48169, n48170, n48171,
         n48172, n48173, n48174, n48175, n48176, n48177, n48178, n48179,
         n48180, n48181, n48182, n48183, n48184, n48185, n48186, n48187,
         n48188, n48189, n48190, n48191, n48192, n48193, n48194, n48195,
         n48196, n48197, n48198, n48199, n48200, n48201, n48202, n48203,
         n48204, n48205, n48206, n48207, n48208, n48209, n48210, n48211,
         n48212, n48213, n48214, n48215, n48216, n48217, n48218, n48219,
         n48220, n48221, n48222, n48223, n48224, n48225, n48226, n48227,
         n48228, n48229, n48230, n48231, n48232, n48233, n48234, n48235,
         n48236, n48237, n48238, n48239, n48240, n48241, n48242, n48243,
         n48244, n48245, n48246, n48247, n48248, n48249, n48250, n48251,
         n48252, n48253, n48254, n48255, n48256, n48257, n48258, n48259,
         n48260, n48261, n48262, n48263, n48264, n48265, n48266, n48267,
         n48268, n48269, n48270, n48271, n48272, n48273, n48274, n48275,
         n48276, n48277, n48278, n48279, n48280, n48281, n48282, n48283,
         n48284, n48285, n48286, n48287, n48288, n48289, n48290, n48291,
         n48292, n48293, n48294, n48295, n48296, n48297, n48298, n48299,
         n48300, n48301, n48302, n48303, n48304, n48305, n48306, n48307,
         n48308, n48309, n48310, n48311, n48312, n48313, n48314, n48315,
         n48316, n48317, n48318, n48319, n48320, n48321, n48322, n48323,
         n48324, n48325, n48326, n48327, n48328, n48329, n48330, n48331,
         n48332, n48333, n48334, n48335, n48336, n48337, n48338, n48339,
         n48340, n48341, n48342, n48343, n48344, n48345, n48346, n48347,
         n48348, n48349, n48350, n48351, n48352, n48353, n48354, n48355,
         n48356, n48357, n48358, n48359, n48360, n48361, n48362, n48363,
         n48364, n48365, n48366, n48367, n48368, n48369, n48370, n48371,
         n48372, n48373, n48374, n48375, n48376, n48377, n48378, n48379,
         n48380, n48381, n48382, n48383, n48384, n48385, n48386, n48387,
         n48388, n48389, n48390, n48391, n48392, n48393, n48394, n48395,
         n48396, n48397, n48398, n48399, n48400, n48401, n48402, n48403,
         n48404, n48405, n48406, n48407, n48408, n48409, n48410, n48411,
         n48412, n48413, n48414, n48415, n48416, n48417, n48418, n48419,
         n48420, n48421, n48422, n48423, n48424, n48425, n48426, n48427,
         n48428, n48429, n48430, n48431, n48432, n48433, n48434, n48435,
         n48436, n48437, n48438, n48439, n48440, n48441, n48442, n48443,
         n48444, n48445, n48446, n48447, n48448, n48449, n48450, n48451,
         n48452, n48453, n48454, n48455, n48456, n48457, n48458, n48459,
         n48460, n48461, n48462, n48463, n48464, n48465, n48466, n48467,
         n48468, n48469, n48470, n48471, n48472, n48473, n48474, n48475,
         n48476, n48477, n48478, n48479, n48480, n48481, n48482, n48483,
         n48484, n48485, n48486, n48487, n48488, n48489, n48490, n48491,
         n48492, n48493, n48494, n48495, n48496, n48497, n48498, n48499,
         n48500, n48501, n48502, n48503, n48504, n48505, n48506, n48507,
         n48508, n48509, n48510, n48511, n48512, n48513, n48514, n48515,
         n48516, n48517, n48518, n48519, n48520, n48521, n48522, n48523,
         n48524, n48525, n48526, n48527, n48528, n48529, n48530, n48531,
         n48532, n48533, n48534, n48535, n48536, n48537, n48538, n48539,
         n48540, n48541, n48542, n48543, n48544, n48545, n48546, n48547,
         n48548, n48549, n48550, n48551, n48552, n48553, n48554, n48555,
         n48556, n48557, n48558, n48559, n48560, n48561, n48562, n48563,
         n48564, n48565, n48566, n48567, n48568, n48569, n48570, n48571,
         n48572, n48573, n48574, n48575, n48576, n48577, n48578, n48579,
         n48580, n48581, n48582, n48583, n48584, n48585, n48586, n48587,
         n48588, n48589, n48590, n48591, n48592, n48593, n48594, n48595,
         n48596, n48597, n48598, n48599, n48600, n48601, n48602, n48603,
         n48604, n48605, n48606, n48607, n48608, n48609, n48610, n48611,
         n48612, n48613, n48614, n48615, n48616, n48617, n48618, n48619,
         n48620, n48621, n48622, n48623, n48624, n48625, n48626, n48627,
         n48628, n48629, n48630, n48631, n48632, n48633, n48634, n48635,
         n48636, n48637, n48638, n48639, n48640, n48641, n48642, n48643,
         n48644, n48645, n48646, n48647, n48648, n48649, n48650, n48651,
         n48652, n48653, n48654, n48655, n48656, n48657, n48658, n48659,
         n48660, n48661, n48662, n48663, n48664, n48665, n48666, n48667,
         n48668, n48669, n48670, n48671, n48672, n48673, n48674, n48675,
         n48676, n48677, n48678, n48679, n48680, n48681, n48682, n48683,
         n48684, n48685, n48686, n48687, n48688, n48689, n48690, n48691,
         n48692, n48693, n48694, n48695, n48696, n48697, n48698, n48699,
         n48700, n48701, n48702, n48703, n48704, n48705, n48706, n48707,
         n48708, n48709, n48710, n48711, n48712, n48713, n48714, n48715,
         n48716, n48717, n48718, n48719, n48720, n48721, n48722, n48723,
         n48724, n48725, n48726, n48727, n48728, n48729, n48730, n48731,
         n48732, n48733, n48734, n48735, n48736, n48737, n48738, n48739,
         n48740, n48741, n48742, n48743, n48744, n48745, n48746, n48747,
         n48748, n48749, n48750, n48751, n48752, n48753, n48754, n48755,
         n48756, n48757, n48758, n48759, n48760, n48761, n48762, n48763,
         n48764, n48765, n48766, n48767, n48768, n48769, n48770, n48771,
         n48772, n48773, n48774, n48775, n48776, n48777, n48778, n48779,
         n48780, n48781, n48782, n48783, n48784, n48785, n48786, n48787,
         n48788, n48789, n48790, n48791, n48792, n48793, n48794, n48795,
         n48796, n48797, n48798, n48799, n48800, n48801, n48802, n48803,
         n48804, n48805, n48806, n48807, n48808, n48809, n48810, n48811,
         n48812, n48813, n48814, n48815, n48816, n48817, n48818, n48819,
         n48820, n48821, n48822, n48823, n48824, n48825, n48826, n48827,
         n48828, n48829, n48830, n48831, n48832, n48833, n48834, n48835,
         n48836, n48837, n48838, n48839, n48840, n48841, n48842, n48843,
         n48844, n48845, n48846, n48847, n48848, n48849, n48850, n48851,
         n48852, n48853, n48854, n48855, n48856, n48857, n48858, n48859,
         n48860, n48861, n48862, n48863, n48864, n48865, n48866, n48867,
         n48868, n48869, n48870, n48871, n48872, n48873, n48874, n48875,
         n48876, n48877, n48878, n48879, n48880, n48881, n48882, n48883,
         n48884, n48885, n48886, n48887, n48888, n48889, n48890, n48891,
         n48892, n48893, n48894, n48895, n48896, n48897, n48898, n48899,
         n48900, n48901, n48902, n48903, n48904, n48905, n48906, n48907,
         n48908, n48909, n48910, n48911, n48912, n48913, n48914, n48915,
         n48916, n48917, n48918, n48919, n48920, n48921, n48922, n48923,
         n48924, n48925, n48926, n48927, n48928, n48929, n48930, n48931,
         n48932, n48933, n48934, n48935, n48936, n48937, n48938, n48939,
         n48940, n48941, n48942, n48943, n48944, n48945, n48946, n48947,
         n48948, n48949, n48950, n48951, n48952, n48953, n48954, n48955,
         n48956, n48957, n48958, n48959, n48960, n48961, n48962, n48963,
         n48964, n48965, n48966, n48967, n48968, n48969, n48970, n48971,
         n48972, n48973, n48974, n48975, n48976, n48977, n48978, n48979,
         n48980, n48981, n48982, n48983, n48984, n48985, n48986, n48987,
         n48988, n48989, n48990, n48991, n48992, n48993, n48994, n48995,
         n48996, n48997, n48998, n48999, n49000, n49001, n49002, n49003,
         n49004, n49005, n49006, n49007, n49008, n49009, n49010, n49011,
         n49012, n49013, n49014, n49015, n49016, n49017, n49018, n49019,
         n49020, n49021, n49022, n49023, n49024, n49025, n49026, n49027,
         n49028, n49029, n49030, n49031, n49032, n49033, n49034, n49035,
         n49036, n49037, n49038, n49039, n49040, n49041, n49042, n49043,
         n49044, n49045, n49046, n49047, n49048, n49049, n49050, n49051,
         n49052, n49053, n49054, n49055, n49056, n49057, n49058, n49059,
         n49060, n49061, n49062, n49063, n49064, n49065, n49066, n49067,
         n49068, n49069, n49070, n49071, n49072, n49073, n49074, n49075,
         n49076, n49077, n49078, n49079, n49080, n49081, n49082, n49083,
         n49084, n49085, n49086, n49087, n49088, n49089, n49090, n49091,
         n49092, n49093, n49094, n49095, n49096, n49097, n49098, n49099,
         n49100, n49101, n49102, n49103, n49104, n49105, n49106, n49107,
         n49108, n49109, n49110, n49111, n49112, n49113, n49114, n49115,
         n49116, n49117, n49118, n49119, n49120, n49121, n49122, n49123,
         n49124, n49125, n49126, n49127, n49128, n49129, n49130, n49131,
         n49132, n49133, n49134, n49135, n49136, n49137, n49138, n49139,
         n49140, n49141, n49142, n49143, n49144, n49145, n49146, n49147,
         n49148, n49149, n49150, n49151, n49152, n49153, n49154, n49155,
         n49156, n49157, n49158, n49159, n49160, n49161, n49162, n49163,
         n49164, n49165, n49166, n49167, n49168, n49169, n49170, n49171,
         n49172, n49173, n49174, n49175, n49176, n49177, n49178, n49179,
         n49180, n49181, n49182, n49183, n49184, n49185, n49186, n49187,
         n49188, n49189, n49190, n49191, n49192, n49193, n49194, n49195,
         n49196, n49197, n49198, n49199, n49200, n49201, n49202, n49203,
         n49204, n49205, n49206, n49207, n49208, n49209, n49210, n49211,
         n49212, n49213, n49214, n49215, n49216, n49217, n49218, n49219,
         n49220, n49221, n49222, n49223, n49224, n49225, n49226, n49227,
         n49228, n49229, n49230, n49231, n49232, n49233, n49234, n49235,
         n49236, n49237, n49238, n49239, n49240, n49241, n49242, n49243,
         n49244, n49245, n49246, n49247, n49248, n49249, n49250, n49251,
         n49252, n49253, n49254, n49255, n49256, n49257, n49258, n49259,
         n49260, n49261, n49262, n49263, n49264, n49265, n49266, n49267,
         n49268, n49269, n49270, n49271, n49272, n49273, n49274, n49275,
         n49276, n49277, n49278, n49279, n49280, n49281, n49282, n49283,
         n49284, n49285, n49286, n49287, n49288, n49289, n49290, n49291,
         n49292, n49293, n49294, n49295, n49296, n49297, n49298, n49299,
         n49300, n49301, n49302, n49303, n49304, n49305, n49306, n49307,
         n49308, n49309, n49310, n49311, n49312, n49313, n49314, n49315,
         n49316, n49317, n49318, n49319, n49320, n49321, n49322, n49323,
         n49324, n49325, n49326, n49327, n49328, n49329, n49330, n49331,
         n49332, n49333, n49334, n49335, n49336, n49337, n49338, n49339,
         n49340, n49341, n49342, n49343, n49344, n49345, n49346, n49347,
         n49348, n49349, n49350, n49351, n49352, n49353, n49354, n49355,
         n49356, n49357, n49358, n49359, n49360, n49361, n49362, n49363,
         n49364, n49365, n49366, n49367, n49368, n49369, n49370, n49371,
         n49372, n49373, n49374, n49375, n49376, n49377, n49378, n49379,
         n49380, n49381, n49382, n49383, n49384, n49385, n49386, n49387,
         n49388, n49389, n49390, n49391, n49392, n49393, n49394, n49395,
         n49396, n49397, n49398, n49399, n49400, n49401, n49402, n49403,
         n49404, n49405, n49406, n49407, n49408, n49409, n49410, n49411,
         n49412, n49413, n49414, n49415, n49416, n49417, n49418, n49419,
         n49420, n49421, n49422, n49423, n49424, n49425, n49426, n49427,
         n49428, n49429, n49430, n49431, n49432, n49433, n49434, n49435,
         n49436, n49437, n49438, n49439, n49440, n49441, n49442, n49443,
         n49444, n49445, n49446, n49447, n49448, n49449, n49450, n49451,
         n49452, n49453, n49454, n49455, n49456, n49457, n49458, n49459,
         n49460, n49461, n49462, n49463, n49464, n49465, n49466, n49467,
         n49468, n49469, n49470, n49471, n49472, n49473, n49474, n49475,
         n49476, n49477, n49478, n49479, n49480, n49481, n49482, n49483,
         n49484, n49485, n49486, n49487, n49488, n49489, n49490, n49491,
         n49492, n49493, n49494, n49495, n49496, n49497, n49498, n49499,
         n49500, n49501, n49502, n49503, n49504, n49505, n49506, n49507,
         n49508, n49509, n49510, n49511, n49512, n49513, n49514, n49515,
         n49516, n49517, n49518, n49519, n49520, n49521, n49522, n49523,
         n49524, n49525, n49526, n49527, n49528, n49529, n49530, n49531,
         n49532, n49533, n49534, n49535, n49536, n49537, n49538, n49539,
         n49540, n49541, n49542, n49543, n49544, n49545, n49546, n49547,
         n49548, n49549, n49550, n49551, n49552, n49553, n49554, n49555,
         n49556, n49557, n49558, n49559, n49560, n49561, n49562, n49563,
         n49564, n49565, n49566, n49567, n49568, n49569, n49570, n49571,
         n49572, n49573, n49574, n49575, n49576, n49577, n49578, n49579,
         n49580, n49581, n49582, n49583, n49584, n49585, n49586, n49587,
         n49588, n49589, n49590, n49591, n49592, n49593, n49594, n49595,
         n49596, n49597, n49598, n49599, n49600, n49601, n49602, n49603,
         n49604, n49605, n49606, n49607, n49608, n49609, n49610, n49611,
         n49612, n49613, n49614, n49615, n49616, n49617, n49618, n49619,
         n49620, n49621, n49622, n49623, n49624, n49625, n49626, n49627,
         n49628, n49629, n49630, n49631, n49632, n49633, n49634, n49635,
         n49636, n49637, n49638, n49639, n49640, n49641, n49642, n49643,
         n49644, n49645, n49646, n49647, n49648, n49649, n49650, n49651,
         n49652, n49653, n49654, n49655, n49656, n49657, n49658, n49659,
         n49660, n49661, n49662, n49663, n49664, n49665, n49666, n49667,
         n49668, n49669, n49670, n49671, n49672, n49673, n49674, n49675,
         n49676, n49677, n49678, n49679, n49680, n49681, n49682, n49683,
         n49684, n49685, n49686, n49687, n49688, n49689, n49690, n49691,
         n49692, n49693, n49694, n49695, n49696, n49697, n49698, n49699,
         n49700, n49701, n49702, n49703, n49704, n49705, n49706, n49707,
         n49708, n49709, n49710, n49711, n49712, n49713, n49714, n49715,
         n49716, n49717, n49718, n49719, n49720, n49721, n49722, n49723,
         n49724, n49725, n49726, n49727, n49728, n49729, n49730, n49731,
         n49732, n49733, n49734, n49735, n49736, n49737, n49738, n49739,
         n49740, n49741, n49742, n49743, n49744, n49745, n49746, n49747,
         n49748, n49749, n49750, n49751, n49752, n49753, n49754, n49755,
         n49756, n49757, n49758, n49759, n49760, n49761, n49762, n49763,
         n49764, n49765, n49766, n49767, n49768, n49769, n49770, n49771,
         n49772, n49773, n49774, n49775, n49776, n49777, n49778, n49779,
         n49780, n49781, n49782, n49783, n49784, n49785, n49786, n49787,
         n49788, n49789, n49790, n49791, n49792, n49793, n49794, n49795,
         n49796, n49797, n49798, n49799, n49800, n49801, n49802, n49803,
         n49804, n49805, n49806, n49807, n49808, n49809, n49810, n49811,
         n49812, n49813, n49814, n49815, n49816, n49817, n49818, n49819,
         n49820, n49821, n49822, n49823, n49824, n49825, n49826, n49827,
         n49828, n49829, n49830, n49831, n49832, n49833, n49834, n49835,
         n49836, n49837, n49838, n49839, n49840, n49841, n49842, n49843,
         n49844, n49845, n49846, n49847, n49848, n49849, n49850, n49851,
         n49852, n49853, n49854, n49855, n49856, n49857, n49858, n49859,
         n49860, n49861, n49862, n49863, n49864, n49865, n49866, n49867,
         n49868, n49869, n49870, n49871, n49872, n49873, n49874, n49875,
         n49876, n49877, n49878, n49879, n49880, n49881, n49882, n49883,
         n49884, n49885, n49886, n49887, n49888, n49889, n49890, n49891,
         n49892, n49893, n49894, n49895, n49896, n49897, n49898, n49899,
         n49900, n49901, n49902, n49903, n49904, n49905, n49906, n49907,
         n49908, n49909, n49910, n49911, n49912, n49913, n49914, n49915,
         n49916, n49917, n49918, n49919, n49920, n49921, n49922, n49923,
         n49924, n49925, n49926, n49927, n49928, n49929, n49930, n49931,
         n49932, n49933, n49934, n49935, n49936, n49937, n49938, n49939,
         n49940, n49941, n49942, n49943, n49944, n49945, n49946, n49947,
         n49948, n49949, n49950, n49951, n49952, n49953, n49954, n49955,
         n49956, n49957, n49958, n49959, n49960, n49961, n49962, n49963,
         n49964, n49965, n49966, n49967, n49968, n49969, n49970, n49971,
         n49972, n49973, n49974, n49975, n49976, n49977, n49978, n49979,
         n49980, n49981, n49982, n49983, n49984, n49985, n49986, n49987,
         n49988, n49989, n49990, n49991, n49992, n49993, n49994, n49995,
         n49996, n49997, n49998, n49999, n50000, n50001, n50002, n50003,
         n50004, n50005, n50006, n50007, n50008, n50009, n50010, n50011,
         n50012, n50013, n50014, n50015, n50016, n50017, n50018, n50019,
         n50020, n50021, n50022, n50023, n50024, n50025, n50026, n50027,
         n50028, n50029, n50030, n50031, n50032, n50033, n50034, n50035,
         n50036, n50037, n50038, n50039, n50040, n50041, n50042, n50043,
         n50044, n50045, n50046, n50047, n50048, n50049, n50050, n50051,
         n50052, n50053, n50054, n50055, n50056, n50057, n50058, n50059,
         n50060, n50061, n50062, n50063, n50064, n50065, n50066, n50067,
         n50068, n50069, n50070, n50071, n50072, n50073, n50074, n50075,
         n50076, n50077, n50078, n50079, n50080, n50081, n50082, n50083,
         n50084, n50085, n50086, n50087, n50088, n50089, n50090, n50091,
         n50092, n50093, n50094, n50095, n50096, n50097, n50098, n50099,
         n50100, n50101, n50102, n50103, n50104, n50105, n50106, n50107,
         n50108, n50109, n50110, n50111, n50112, n50113, n50114, n50115,
         n50116, n50117, n50118, n50119, n50120, n50121, n50122, n50123,
         n50124, n50125, n50126, n50127, n50128, n50129, n50130, n50131,
         n50132, n50133, n50134, n50135, n50136, n50137, n50138, n50139,
         n50140, n50141, n50142, n50143, n50144, n50145, n50146, n50147,
         n50148, n50149, n50150, n50151, n50152, n50153, n50154, n50155,
         n50156, n50157, n50158, n50159, n50160, n50161, n50162, n50163,
         n50164, n50165, n50166, n50167, n50168, n50169, n50170, n50171,
         n50172, n50173, n50174, n50175, n50176, n50177, n50178, n50179,
         n50180, n50181, n50182, n50183, n50184, n50185, n50186, n50187,
         n50188, n50189, n50190, n50191, n50192, n50193, n50194, n50195,
         n50196, n50197, n50198, n50199, n50200, n50201, n50202, n50203,
         n50204, n50205, n50206, n50207, n50208, n50209, n50210, n50211,
         n50212, n50213, n50214, n50215, n50216, n50217, n50218, n50219,
         n50220, n50221, n50222, n50223, n50224, n50225, n50226, n50227,
         n50228, n50229, n50230, n50231, n50232, n50233, n50234, n50235,
         n50236, n50237, n50238, n50239, n50240, n50241, n50242, n50243,
         n50244, n50245, n50246, n50247, n50248, n50249, n50250, n50251,
         n50252, n50253, n50254, n50255, n50256, n50257, n50258, n50259,
         n50260, n50261, n50262, n50263, n50264, n50265, n50266, n50267,
         n50268, n50269, n50270, n50271, n50272, n50273, n50274, n50275,
         n50276, n50277, n50278, n50279, n50280, n50281, n50282, n50283,
         n50284, n50285, n50286, n50287, n50288, n50289, n50290, n50291,
         n50292, n50293, n50294, n50295, n50296, n50297, n50298, n50299,
         n50300, n50301, n50302, n50303, n50304, n50305, n50306, n50307,
         n50308, n50309, n50310, n50311, n50312, n50313, n50314, n50315,
         n50316, n50317, n50318, n50319, n50320, n50321, n50322, n50323,
         n50324, n50325, n50326, n50327, n50328, n50329, n50330, n50331,
         n50332, n50333, n50334, n50335, n50336, n50337, n50338, n50339,
         n50340, n50341, n50342, n50343, n50344, n50345, n50346, n50347,
         n50348, n50349, n50350, n50351, n50352, n50353, n50354, n50355,
         n50356, n50357, n50358, n50359, n50360, n50361, n50362, n50363,
         n50364, n50365, n50366, n50367, n50368, n50369, n50370, n50371,
         n50372, n50373, n50374, n50375, n50376, n50377, n50378, n50379,
         n50380, n50381, n50382, n50383, n50384, n50385, n50386, n50387,
         n50388, n50389, n50390, n50391, n50392, n50393, n50394, n50395,
         n50396, n50397, n50398, n50399, n50400, n50401, n50402, n50403,
         n50404, n50405, n50406, n50407, n50408, n50409, n50410, n50411,
         n50412, n50413, n50414, n50415, n50416, n50417, n50418, n50419,
         n50420, n50421, n50422, n50423, n50424, n50425, n50426, n50427,
         n50428, n50429, n50430, n50431, n50432, n50433, n50434, n50435,
         n50436, n50437, n50438, n50439, n50440, n50441, n50442, n50443,
         n50444, n50445, n50446, n50447, n50448, n50449, n50450, n50451,
         n50452, n50453, n50454, n50455, n50456, n50457, n50458, n50459,
         n50460, n50461, n50462, n50463, n50464, n50465, n50466, n50467,
         n50468, n50469, n50470, n50471, n50472, n50473, n50474, n50475,
         n50476, n50477, n50478, n50479, n50480, n50481, n50482, n50483,
         n50484, n50485, n50486, n50487, n50488, n50489, n50490, n50491,
         n50492, n50493, n50494, n50495, n50496, n50497, n50498, n50499,
         n50500, n50501, n50502, n50503, n50504, n50505, n50506, n50507,
         n50508, n50509, n50510, n50511, n50512, n50513, n50514, n50515,
         n50516, n50517, n50518, n50519, n50520, n50521, n50522, n50523,
         n50524, n50525, n50526, n50527, n50528, n50529, n50530, n50531,
         n50532, n50533, n50534, n50535, n50536, n50537, n50538, n50539,
         n50540, n50541, n50542, n50543, n50544, n50545, n50546, n50547,
         n50548, n50549, n50550, n50551, n50552, n50553, n50554, n50555,
         n50556, n50557, n50558, n50559, n50560, n50561, n50562, n50563,
         n50564, n50565, n50566, n50567, n50568, n50569, n50570, n50571,
         n50572, n50573, n50574, n50575, n50576, n50577, n50578, n50579,
         n50580, n50581, n50582, n50583, n50584, n50585, n50586, n50587,
         n50588, n50589, n50590, n50591, n50592, n50593, n50594, n50595,
         n50596, n50597, n50598, n50599, n50600, n50601, n50602, n50603,
         n50604, n50605, n50606, n50607, n50608, n50609, n50610, n50611,
         n50612, n50613, n50614, n50615, n50616, n50617, n50618, n50619,
         n50620, n50621, n50622, n50623, n50624, n50625, n50626, n50627,
         n50628, n50629, n50630, n50631, n50632, n50633, n50634, n50635,
         n50636, n50637, n50638, n50639, n50640, n50641, n50642, n50643,
         n50644, n50645, n50646, n50647, n50648, n50649, n50650, n50651,
         n50652, n50653, n50654, n50655, n50656, n50657, n50658, n50659,
         n50660, n50661, n50662, n50663, n50664, n50665, n50666, n50667,
         n50668, n50669, n50670, n50671, n50672, n50673, n50674, n50675,
         n50676, n50677, n50678, n50679, n50680, n50681, n50682, n50683,
         n50684, n50685, n50686, n50687, n50688, n50689, n50690, n50691,
         n50692, n50693, n50694, n50695, n50696, n50697, n50698, n50699,
         n50700, n50701, n50702, n50703, n50704, n50705, n50706, n50707,
         n50708, n50709, n50710, n50711, n50712, n50713, n50714, n50715,
         n50716, n50717, n50718, n50719, n50720, n50721, n50722, n50723,
         n50724, n50725, n50726, n50727, n50728, n50729, n50730, n50731,
         n50732, n50733, n50734, n50735, n50736, n50737, n50738, n50739,
         n50740, n50741, n50742, n50743, n50744, n50745, n50746, n50747,
         n50748, n50749, n50750, n50751, n50752, n50753, n50754, n50755,
         n50756, n50757, n50758, n50759, n50760, n50761, n50762, n50763,
         n50764, n50765, n50766, n50767, n50768, n50769, n50770, n50771,
         n50772, n50773, n50774, n50775, n50776, n50777, n50778, n50779,
         n50780, n50781, n50782, n50783, n50784, n50785, n50786, n50787,
         n50788, n50789, n50790, n50791, n50792, n50793, n50794, n50795,
         n50796, n50797, n50798, n50799, n50800, n50801, n50802, n50803,
         n50804, n50805, n50806, n50807, n50808, n50809, n50810, n50811,
         n50812, n50813, n50814, n50815, n50816, n50817, n50818, n50819,
         n50820, n50821, n50822, n50823, n50824, n50825, n50826, n50827,
         n50828, n50829, n50830, n50831, n50832, n50833, n50834, n50835,
         n50836, n50837, n50838, n50839, n50840, n50841, n50842, n50843,
         n50844, n50845, n50846, n50847, n50848, n50849, n50850, n50851,
         n50852, n50853, n50854, n50855, n50856, n50857, n50858, n50859,
         n50860, n50861, n50862, n50863, n50864, n50865, n50866, n50867,
         n50868, n50869, n50870, n50871, n50872, n50873, n50874, n50875,
         n50876, n50877, n50878, n50879, n50880, n50881, n50882, n50883,
         n50884, n50885, n50886, n50887, n50888, n50889, n50890, n50891,
         n50892, n50893, n50894, n50895, n50896, n50897, n50898, n50899,
         n50900, n50901, n50902, n50903, n50904, n50905, n50906, n50907,
         n50908, n50909, n50910, n50911, n50912, n50913, n50914, n50915,
         n50916, n50917, n50918, n50919, n50920, n50921, n50922, n50923,
         n50924, n50925, n50926, n50927, n50928, n50929, n50930, n50931,
         n50932, n50933, n50934, n50935, n50936, n50937, n50938, n50939,
         n50940, n50941, n50942, n50943, n50944, n50945, n50946, n50947,
         n50948, n50949, n50950, n50951, n50952, n50953, n50954, n50955,
         n50956, n50957, n50958, n50959, n50960, n50961, n50962, n50963,
         n50964, n50965, n50966, n50967, n50968, n50969, n50970, n50971,
         n50972, n50973, n50974, n50975, n50976, n50977, n50978, n50979,
         n50980, n50981, n50982, n50983, n50984, n50985, n50986, n50987,
         n50988, n50989, n50990, n50991, n50992, n50993, n50994, n50995,
         n50996, n50997, n50998, n50999, n51000, n51001, n51002, n51003,
         n51004, n51005, n51006, n51007, n51008, n51009, n51010, n51011,
         n51012, n51013, n51014, n51015, n51016, n51017, n51018, n51019,
         n51020, n51021, n51022, n51023, n51024, n51025, n51026, n51027,
         n51028, n51029, n51030, n51031, n51032, n51033, n51034, n51035,
         n51036, n51037, n51038, n51039, n51040, n51041, n51042, n51043,
         n51044, n51045, n51046, n51047, n51048, n51049, n51050, n51051,
         n51052, n51053, n51054, n51055, n51056, n51057, n51058, n51059,
         n51060, n51061, n51062, n51063, n51064, n51065, n51066, n51067,
         n51068, n51069, n51070, n51071, n51072, n51073, n51074, n51075,
         n51076, n51077, n51078, n51079, n51080, n51081, n51082, n51083,
         n51084, n51085, n51086, n51087, n51088, n51089, n51090, n51091,
         n51092, n51093, n51094, n51095, n51096, n51097, n51098, n51099,
         n51100, n51101, n51102, n51103, n51104, n51105, n51106, n51107,
         n51108, n51109, n51110, n51111, n51112, n51113, n51114, n51115,
         n51116, n51117, n51118, n51119, n51120, n51121, n51122, n51123,
         n51124, n51125, n51126, n51127, n51128, n51129, n51130, n51131,
         n51132, n51133, n51134, n51135, n51136, n51137, n51138, n51139,
         n51140, n51141, n51142, n51143, n51144, n51145, n51146, n51147,
         n51148, n51149, n51150, n51151, n51152, n51153, n51154, n51155,
         n51156, n51157, n51158, n51159, n51160, n51161, n51162, n51163,
         n51164, n51165, n51166, n51167, n51168, n51169, n51170, n51171,
         n51172, n51173, n51174, n51175, n51176, n51177, n51178, n51179,
         n51180, n51181, n51182, n51183, n51184, n51185, n51186, n51187,
         n51188, n51189, n51190, n51191, n51192, n51193, n51194, n51195,
         n51196, n51197, n51198, n51199, n51200, n51201, n51202, n51203,
         n51204, n51205, n51206, n51207, n51208, n51209, n51210, n51211,
         n51212, n51213, n51214, n51215, n51216, n51217, n51218, n51219,
         n51220, n51221, n51222, n51223, n51224, n51225, n51226, n51227,
         n51228, n51229, n51230, n51231, n51232, n51233, n51234, n51235,
         n51236, n51237, n51238, n51239, n51240, n51241, n51242, n51243,
         n51244, n51245, n51246, n51247, n51248, n51249, n51250, n51251,
         n51252, n51253, n51254, n51255, n51256, n51257, n51258, n51259,
         n51260, n51261, n51262, n51263, n51264, n51265, n51266, n51267,
         n51268, n51269, n51270, n51271, n51272, n51273, n51274, n51275,
         n51276, n51277, n51278, n51279, n51280, n51281, n51282, n51283,
         n51284, n51285, n51286, n51287, n51288, n51289, n51290, n51291,
         n51292, n51293, n51294, n51295, n51296, n51297, n51298, n51299,
         n51300, n51301, n51302, n51303, n51304, n51305, n51306, n51307,
         n51308, n51309, n51310, n51311, n51312, n51313, n51314, n51315,
         n51316, n51317, n51318, n51319, n51320, n51321, n51322, n51323,
         n51324, n51325, n51326, n51327, n51328, n51329, n51330, n51331,
         n51332, n51333, n51334, n51335, n51336, n51337, n51338, n51339,
         n51340, n51341, n51342, n51343, n51344, n51345, n51346, n51347,
         n51348, n51349, n51350, n51351, n51352, n51353, n51354, n51355,
         n51356, n51357, n51358, n51359, n51360, n51361, n51362, n51363,
         n51364, n51365, n51366, n51367, n51368, n51369, n51370, n51371,
         n51372, n51373, n51374, n51375, n51376, n51377, n51378, n51379,
         n51380, n51381, n51382, n51383, n51384, n51385, n51386, n51387,
         n51388, n51389, n51390, n51391, n51392, n51393, n51394, n51395,
         n51396, n51397, n51398, n51399, n51400, n51401, n51402, n51403,
         n51404, n51405, n51406, n51407, n51408, n51409, n51410, n51411,
         n51412, n51413, n51414, n51415, n51416, n51417, n51418, n51419,
         n51420, n51421, n51422, n51423, n51424, n51425, n51426, n51427,
         n51428, n51429, n51430, n51431, n51432, n51433, n51434, n51435,
         n51436, n51437, n51438, n51439, n51440, n51441, n51442, n51443,
         n51444, n51445, n51446, n51447, n51448, n51449, n51450, n51451,
         n51452, n51453, n51454, n51455, n51456, n51457, n51458, n51459,
         n51460, n51461, n51462, n51463, n51464, n51465, n51466, n51467,
         n51468, n51469, n51470, n51471, n51472, n51473, n51474, n51475,
         n51476, n51477, n51478, n51479, n51480, n51481, n51482, n51483,
         n51484, n51485, n51486, n51487, n51488, n51489, n51490, n51491,
         n51492, n51493, n51494, n51495, n51496, n51497, n51498, n51499,
         n51500, n51501, n51502, n51503, n51504, n51505, n51506, n51507,
         n51508, n51509, n51510, n51511, n51512, n51513, n51514, n51515,
         n51516, n51517, n51518, n51519, n51520, n51521, n51522, n51523,
         n51524, n51525, n51526, n51527, n51528, n51529, n51530, n51531,
         n51532, n51533, n51534, n51535, n51536, n51537, n51538, n51539,
         n51540, n51541, n51542, n51543, n51544, n51545, n51546, n51547,
         n51548, n51549, n51550, n51551, n51552, n51553, n51554, n51555,
         n51556, n51557, n51558, n51559, n51560, n51561, n51562, n51563,
         n51564, n51565, n51566, n51567, n51568, n51569, n51570, n51571,
         n51572, n51573, n51574, n51575, n51576, n51577, n51578, n51579,
         n51580, n51581, n51582, n51583, n51584, n51585, n51586, n51587,
         n51588, n51589, n51590, n51591, n51592, n51593, n51594, n51595,
         n51596, n51597, n51598, n51599, n51600, n51601, n51602, n51603,
         n51604, n51605, n51606, n51607, n51608, n51609, n51610, n51611,
         n51612, n51613, n51614, n51615, n51616, n51617, n51618, n51619,
         n51620, n51621, n51622, n51623, n51624, n51625, n51626, n51627,
         n51628, n51629, n51630, n51631, n51632, n51633, n51634, n51635,
         n51636, n51637, n51638, n51639, n51640, n51641, n51642, n51643,
         n51644, n51645, n51646, n51647, n51648, n51649, n51650, n51651,
         n51652, n51653, n51654, n51655, n51656, n51657, n51658, n51659,
         n51660, n51661, n51662, n51663, n51664, n51665, n51666, n51667,
         n51668, n51669, n51670, n51671, n51672, n51673, n51674, n51675,
         n51676, n51677, n51678, n51679, n51680, n51681, n51682, n51683,
         n51684, n51685, n51686, n51687, n51688, n51689, n51690, n51691,
         n51692, n51693, n51694, n51695, n51696, n51697, n51698, n51699,
         n51700, n51701, n51702, n51703, n51704, n51705, n51706, n51707,
         n51708, n51709, n51710, n51711, n51712, n51713, n51714, n51715,
         n51716, n51717, n51718, n51719, n51720, n51721, n51722, n51723,
         n51724, n51725, n51726, n51727, n51728, n51729, n51730, n51731,
         n51732, n51733, n51734, n51735, n51736, n51737, n51738, n51739,
         n51740, n51741, n51742, n51743, n51744, n51745, n51746, n51747,
         n51748, n51749, n51750, n51751, n51752, n51753, n51754, n51755,
         n51756, n51757, n51758, n51759, n51760, n51761, n51762, n51763,
         n51764, n51765, n51766, n51767, n51768, n51769, n51770, n51771,
         n51772, n51773, n51774, n51775, n51776, n51777, n51778, n51779,
         n51780, n51781, n51782, n51783, n51784, n51785, n51786, n51787,
         n51788, n51789, n51790, n51791, n51792, n51793, n51794, n51795,
         n51796, n51797, n51798, n51799, n51800, n51801, n51802, n51803,
         n51804, n51805, n51806, n51807, n51808, n51809, n51810, n51811,
         n51812, n51813, n51814, n51815, n51816, n51817, n51818, n51819,
         n51820, n51821, n51822, n51823, n51824, n51825, n51826, n51827,
         n51828, n51829, n51830, n51831, n51832, n51833, n51834, n51835,
         n51836, n51837, n51838, n51839, n51840, n51841, n51842, n51843,
         n51844, n51845, n51846, n51847, n51848, n51849, n51850, n51851,
         n51852, n51853, n51854, n51855, n51856, n51857, n51858, n51859,
         n51860, n51861, n51862, n51863, n51864, n51865, n51866, n51867,
         n51868, n51869, n51870, n51871, n51872, n51873, n51874, n51875,
         n51876, n51877, n51878, n51879, n51880, n51881, n51882, n51883,
         n51884, n51885, n51886, n51887, n51888, n51889, n51890, n51891,
         n51892, n51893, n51894, n51895, n51896, n51897, n51898, n51899,
         n51900, n51901, n51902, n51903, n51904, n51905, n51906, n51907,
         n51908, n51909, n51910, n51911, n51912, n51913, n51914, n51915,
         n51916, n51917, n51918, n51919, n51920, n51921, n51922, n51923,
         n51924, n51925, n51926, n51927, n51928, n51929, n51930, n51931,
         n51932, n51933, n51934, n51935, n51936, n51937, n51938, n51939,
         n51940, n51941, n51942, n51943, n51944, n51945, n51946, n51947,
         n51948, n51949, n51950, n51951, n51952, n51953, n51954, n51955,
         n51956, n51957, n51958, n51959, n51960, n51961, n51962, n51963,
         n51964, n51965, n51966, n51967, n51968, n51969, n51970, n51971,
         n51972, n51973, n51974, n51975, n51976, n51977, n51978, n51979,
         n51980, n51981, n51982, n51983, n51984, n51985, n51986, n51987,
         n51988, n51989, n51990, n51991, n51992, n51993, n51994, n51995,
         n51996, n51997, n51998, n51999, n52000, n52001, n52002, n52003,
         n52004, n52005, n52006, n52007, n52008, n52009, n52010, n52011,
         n52012, n52013, n52014, n52015, n52016, n52017, n52018, n52019,
         n52020, n52021, n52022, n52023, n52024, n52025, n52026, n52027,
         n52028, n52029, n52030, n52031, n52032, n52033, n52034, n52035,
         n52036, n52037, n52038, n52039, n52040, n52041, n52042, n52043,
         n52044, n52045, n52046, n52047, n52048, n52049, n52050, n52051,
         n52052, n52053, n52054, n52055, n52056, n52057, n52058, n52059,
         n52060, n52061, n52062, n52063, n52064, n52065, n52066, n52067,
         n52068, n52069, n52070, n52071, n52072, n52073, n52074, n52075,
         n52076, n52077, n52078, n52079, n52080, n52081, n52082, n52083,
         n52084, n52085, n52086, n52087, n52088, n52089, n52090, n52091,
         n52092, n52093, n52094, n52095, n52096, n52097, n52098, n52099,
         n52100, n52101, n52102, n52103, n52104, n52105, n52106, n52107,
         n52108, n52109, n52110, n52111, n52112, n52113, n52114, n52115,
         n52116, n52117, n52118, n52119, n52120, n52121, n52122, n52123,
         n52124, n52125, n52126, n52127, n52128, n52129, n52130, n52131,
         n52132, n52133, n52134, n52135, n52136, n52137, n52138, n52139,
         n52140, n52141, n52142, n52143, n52144, n52145, n52146, n52147,
         n52148, n52149, n52150, n52151, n52152, n52153, n52154, n52155,
         n52156, n52157, n52158, n52159, n52160, n52161, n52162, n52163,
         n52164, n52165, n52166, n52167, n52168, n52169, n52170, n52171,
         n52172, n52173, n52174, n52175, n52176, n52177, n52178, n52179,
         n52180, n52181, n52182, n52183, n52184, n52185, n52186, n52187,
         n52188, n52189, n52190, n52191, n52192, n52193, n52194, n52195,
         n52196, n52197, n52198, n52199, n52200, n52201, n52202, n52203,
         n52204, n52205, n52206, n52207, n52208, n52209, n52210, n52211,
         n52212, n52213, n52214, n52215, n52216, n52217, n52218, n52219,
         n52220, n52221, n52222, n52223, n52224, n52225, n52226, n52227,
         n52228, n52229, n52230, n52231, n52232, n52233, n52234, n52235,
         n52236, n52237, n52238, n52239, n52240, n52241, n52242, n52243,
         n52244, n52245, n52246, n52247, n52248, n52249, n52250, n52251,
         n52252, n52253, n52254, n52255, n52256, n52257, n52258, n52259,
         n52260, n52261, n52262, n52263, n52264, n52265, n52266, n52267,
         n52268, n52269, n52270, n52271, n52272, n52273, n52274, n52275,
         n52276, n52277, n52278, n52279, n52280, n52281, n52282, n52283,
         n52284, n52285, n52286, n52287, n52288, n52289, n52290, n52291,
         n52292, n52293, n52294, n52295, n52296, n52297, n52298, n52299,
         n52300, n52301, n52302, n52303, n52304, n52305, n52306, n52307,
         n52308, n52309, n52310, n52311, n52312, n52313, n52314, n52315,
         n52316, n52317, n52318, n52319, n52320, n52321, n52322, n52323,
         n52324, n52325, n52326, n52327, n52328, n52329, n52330, n52331,
         n52332, n52333, n52334, n52335, n52336, n52337, n52338, n52339,
         n52340, n52341, n52342, n52343, n52344, n52345, n52346, n52347,
         n52348, n52349, n52350, n52351, n52352, n52353, n52354, n52355,
         n52356, n52357, n52358, n52359, n52360, n52361, n52362, n52363,
         n52364, n52365, n52366, n52367, n52368, n52369, n52370, n52371,
         n52372, n52373, n52374, n52375, n52376, n52377, n52378, n52379,
         n52380, n52381, n52382, n52383, n52384, n52385, n52386, n52387,
         n52388, n52389, n52390, n52391, n52392, n52393, n52394, n52395,
         n52396, n52397, n52398, n52399, n52400, n52401, n52402, n52403,
         n52404, n52405, n52406, n52407, n52408, n52409, n52410, n52411,
         n52412, n52413, n52414, n52415, n52416, n52417, n52418, n52419,
         n52420, n52421, n52422, n52423, n52424, n52425, n52426, n52427,
         n52428, n52429, n52430, n52431, n52432, n52433, n52434, n52435,
         n52436, n52437, n52438, n52439, n52440, n52441, n52442, n52443,
         n52444, n52445, n52446, n52447, n52448, n52449, n52450, n52451,
         n52452, n52453, n52454, n52455, n52456, n52457, n52458, n52459,
         n52460, n52461, n52462, n52463, n52464, n52465, n52466, n52467,
         n52468, n52469, n52470, n52471, n52472, n52473, n52474, n52475,
         n52476, n52477, n52478, n52479, n52480, n52481, n52482, n52483,
         n52484, n52485, n52486, n52487, n52488, n52489, n52490, n52491,
         n52492, n52493, n52494, n52495, n52496, n52497, n52498, n52499,
         n52500, n52501, n52502, n52503, n52504, n52505, n52506, n52507,
         n52508, n52509, n52510, n52511, n52512, n52513, n52514, n52515,
         n52516, n52517, n52518, n52519, n52520, n52521, n52522, n52523,
         n52524, n52525, n52526, n52527, n52528, n52529, n52530, n52531,
         n52532, n52533, n52534, n52535, n52536, n52537, n52538, n52539,
         n52540, n52541, n52542, n52543, n52544, n52545, n52546, n52547,
         n52548, n52549, n52550, n52551, n52552, n52553, n52554, n52555,
         n52556, n52557, n52558, n52559, n52560, n52561, n52562, n52563,
         n52564, n52565, n52566, n52567, n52568, n52569, n52570, n52571,
         n52572, n52573, n52574, n52575, n52576, n52577, n52578, n52579,
         n52580, n52581, n52582, n52583, n52584, n52585, n52586, n52587,
         n52588, n52589, n52590, n52591, n52592, n52593, n52594, n52595,
         n52596, n52597, n52598, n52599, n52600, n52601, n52602, n52603,
         n52604, n52605, n52606, n52607, n52608, n52609, n52610, n52611,
         n52612, n52613, n52614, n52615, n52616, n52617, n52618, n52619,
         n52620, n52621, n52622, n52623, n52624, n52625, n52626, n52627,
         n52628, n52629, n52630, n52631, n52632, n52633, n52634, n52635,
         n52636, n52637, n52638, n52639, n52640, n52641, n52642, n52643,
         n52644, n52645, n52646, n52647, n52648, n52649, n52650, n52651,
         n52652, n52653, n52654, n52655, n52656, n52657, n52658, n52659,
         n52660, n52661, n52662, n52663, n52664, n52665, n52666, n52667,
         n52668, n52669, n52670, n52671, n52672, n52673, n52674, n52675,
         n52676, n52677, n52678, n52679, n52680, n52681, n52682, n52683,
         n52684, n52685, n52686, n52687, n52688, n52689, n52690, n52691,
         n52692, n52693, n52694, n52695, n52696, n52697, n52698, n52699,
         n52700, n52701, n52702, n52703, n52704, n52705, n52706, n52707,
         n52708, n52709, n52710, n52711, n52712, n52713, n52714, n52715,
         n52716, n52717, n52718, n52719, n52720, n52721, n52722, n52723,
         n52724, n52725, n52726, n52727, n52728, n52729, n52730, n52731,
         n52732, n52733, n52734, n52735, n52736, n52737, n52738, n52739,
         n52740, n52741, n52742, n52743, n52744, n52745, n52746, n52747,
         n52748, n52749, n52750, n52751, n52752, n52753, n52754, n52755,
         n52756, n52757, n52758, n52759, n52760, n52761, n52762, n52763,
         n52764, n52765, n52766, n52767, n52768, n52769, n52770, n52771,
         n52772, n52773, n52774, n52775, n52776, n52777, n52778, n52779,
         n52780, n52781, n52782, n52783, n52784, n52785, n52786, n52787,
         n52788, n52789, n52790, n52791, n52792, n52793, n52794, n52795,
         n52796, n52797, n52798, n52799, n52800, n52801, n52802, n52803,
         n52804, n52805, n52806, n52807, n52808, n52809, n52810, n52811,
         n52812, n52813, n52814, n52815, n52816, n52817, n52818, n52819,
         n52820, n52821, n52822, n52823, n52824, n52825, n52826, n52827,
         n52828, n52829, n52830, n52831, n52832, n52833, n52834, n52835,
         n52836, n52837, n52838, n52839, n52840, n52841, n52842, n52843,
         n52844, n52845, n52846, n52847, n52848, n52849, n52850, n52851,
         n52852, n52853, n52854, n52855, n52856, n52857, n52858, n52859,
         n52860, n52861, n52862, n52863, n52864, n52865, n52866, n52867,
         n52868, n52869, n52870, n52871, n52872, n52873, n52874, n52875,
         n52876, n52877, n52878, n52879, n52880, n52881, n52882, n52883,
         n52884, n52885, n52886, n52887, n52888, n52889, n52890, n52891,
         n52892, n52893, n52894, n52895, n52896, n52897, n52898, n52899,
         n52900, n52901, n52902, n52903, n52904, n52905, n52906, n52907,
         n52908, n52909, n52910, n52911, n52912, n52913, n52914, n52915,
         n52916, n52917, n52918, n52919, n52920, n52921, n52922, n52923,
         n52924, n52925, n52926, n52927, n52928, n52929, n52930, n52931,
         n52932, n52933, n52934, n52935, n52936, n52937, n52938, n52939,
         n52940, n52941, n52942, n52943, n52944, n52945, n52946, n52947,
         n52948, n52949, n52950, n52951, n52952, n52953, n52954, n52955,
         n52956, n52957, n52958, n52959, n52960, n52961, n52962, n52963,
         n52964, n52965, n52966, n52967, n52968, n52969, n52970, n52971,
         n52972, n52973, n52974, n52975, n52976, n52977, n52978, n52979,
         n52980, n52981, n52982, n52983, n52984, n52985, n52986, n52987,
         n52988, n52989, n52990, n52991, n52992, n52993, n52994, n52995,
         n52996, n52997, n52998, n52999, n53000, n53001, n53002, n53003,
         n53004, n53005, n53006, n53007, n53008, n53009, n53010, n53011,
         n53012, n53013, n53014, n53015, n53016, n53017, n53018, n53019,
         n53020, n53021, n53022, n53023, n53024, n53025, n53026, n53027,
         n53028, n53029, n53030, n53031, n53032, n53033, n53034, n53035,
         n53036, n53037, n53038, n53039, n53040, n53041, n53042, n53043,
         n53044, n53045, n53046, n53047, n53048, n53049, n53050, n53051,
         n53052, n53053, n53054, n53055, n53056, n53057, n53058, n53059,
         n53060, n53061, n53062, n53063, n53064, n53065, n53066, n53067,
         n53068, n53069, n53070, n53071, n53072, n53073, n53074, n53075,
         n53076, n53077, n53078, n53079, n53080, n53081, n53082, n53083,
         n53084, n53085, n53086, n53087, n53088, n53089, n53090, n53091,
         n53092, n53093, n53094, n53095, n53096, n53097, n53098, n53099,
         n53100, n53101, n53102, n53103, n53104, n53105, n53106, n53107,
         n53108, n53109, n53110, n53111, n53112, n53113, n53114, n53115,
         n53116, n53117, n53118, n53119, n53120, n53121, n53122, n53123,
         n53124, n53125, n53126, n53127, n53128, n53129, n53130, n53131,
         n53132, n53133, n53134, n53135, n53136, n53137, n53138, n53139,
         n53140, n53141, n53142, n53143, n53144, n53145, n53146, n53147,
         n53148, n53149, n53150, n53151, n53152, n53153, n53154, n53155,
         n53156, n53157, n53158, n53159, n53160, n53161, n53162, n53163,
         n53164, n53165, n53166, n53167, n53168, n53169, n53170, n53171,
         n53172, n53173, n53174, n53175, n53176, n53177, n53178, n53179,
         n53180, n53181, n53182, n53183, n53184, n53185, n53186, n53187,
         n53188, n53189, n53190, n53191, n53192, n53193, n53194, n53195,
         n53196, n53197, n53198, n53199, n53200, n53201, n53202, n53203,
         n53204, n53205, n53206, n53207, n53208, n53209, n53210, n53211,
         n53212, n53213, n53214, n53215, n53216, n53217, n53218, n53219,
         n53220, n53221, n53222, n53223, n53224, n53225, n53226, n53227,
         n53228, n53229, n53230, n53231, n53232, n53233, n53234, n53235,
         n53236, n53237, n53238, n53239, n53240, n53241, n53242, n53243,
         n53244, n53245, n53246, n53247, n53248, n53249, n53250, n53251,
         n53252, n53253, n53254, n53255, n53256, n53257, n53258, n53259,
         n53260, n53261, n53262, n53263, n53264, n53265, n53266, n53267,
         n53268, n53269, n53270, n53271, n53272, n53273, n53274, n53275,
         n53276, n53277, n53278, n53279, n53280, n53281, n53282, n53283,
         n53284, n53285, n53286, n53287, n53288, n53289, n53290, n53291,
         n53292, n53293, n53294, n53295, n53296, n53297, n53298, n53299,
         n53300, n53301, n53302, n53303, n53304, n53305, n53306, n53307,
         n53308, n53309, n53310, n53311, n53312, n53313, n53314, n53315,
         n53316, n53317, n53318, n53319, n53320, n53321, n53322, n53323,
         n53324, n53325, n53326, n53327, n53328, n53329, n53330, n53331,
         n53332, n53333, n53334, n53335, n53336, n53337, n53338, n53339,
         n53340, n53341, n53342, n53343, n53344, n53345, n53346, n53347,
         n53348, n53349, n53350, n53351, n53352, n53353, n53354, n53355,
         n53356, n53357, n53358, n53359, n53360, n53361, n53362, n53363,
         n53364, n53365, n53366, n53367, n53368, n53369, n53370, n53371,
         n53372, n53373, n53374, n53375, n53376, n53377, n53378, n53379,
         n53380, n53381, n53382, n53383, n53384, n53385, n53386, n53387,
         n53388, n53389, n53390, n53391, n53392, n53393, n53394, n53395,
         n53396, n53397, n53398, n53399, n53400, n53401, n53402, n53403,
         n53404, n53405, n53406, n53407, n53408, n53409, n53410, n53411,
         n53412, n53413, n53414, n53415, n53416, n53417, n53418, n53419,
         n53420, n53421, n53422, n53423, n53424, n53425, n53426, n53427,
         n53428, n53429, n53430, n53431, n53432, n53433, n53434, n53435,
         n53436, n53437, n53438, n53439, n53440, n53441, n53442, n53443,
         n53444, n53445, n53446, n53447, n53448, n53449, n53450, n53451,
         n53452, n53453, n53454, n53455, n53456, n53457, n53458, n53459,
         n53460, n53461, n53462, n53463, n53464, n53465, n53466, n53467,
         n53468, n53469, n53470, n53471, n53472, n53473, n53474, n53475,
         n53476, n53477, n53478, n53479, n53480, n53481, n53482, n53483,
         n53484, n53485, n53486, n53487, n53488, n53489, n53490, n53491,
         n53492, n53493, n53494, n53495, n53496, n53497, n53498, n53499,
         n53500, n53501, n53502, n53503, n53504, n53505, n53506, n53507,
         n53508, n53509, n53510, n53511, n53512, n53513, n53514, n53515,
         n53516, n53517, n53518, n53519, n53520, n53521, n53522, n53523,
         n53524, n53525, n53526, n53527, n53528, n53529, n53530, n53531,
         n53532, n53533, n53534, n53535, n53536, n53537, n53538, n53539,
         n53540, n53541, n53542, n53543, n53544, n53545, n53546, n53547,
         n53548, n53549, n53550, n53551, n53552, n53553, n53554, n53555,
         n53556, n53557, n53558, n53559, n53560, n53561, n53562, n53563,
         n53564, n53565, n53566, n53567, n53568, n53569, n53570, n53571,
         n53572, n53573, n53574, n53575, n53576, n53577, n53578, n53579,
         n53580, n53581, n53582, n53583, n53584, n53585, n53586, n53587,
         n53588, n53589, n53590, n53591, n53592, n53593, n53594, n53595,
         n53596, n53597, n53598, n53599, n53600, n53601, n53602, n53603,
         n53604, n53605, n53606, n53607, n53608, n53609, n53610, n53611,
         n53612, n53613, n53614, n53615, n53616, n53617, n53618, n53619,
         n53620, n53621, n53622, n53623, n53624, n53625, n53626, n53627,
         n53628, n53629, n53630, n53631, n53632, n53633, n53634, n53635,
         n53636, n53637, n53638, n53639, n53640, n53641, n53642, n53643,
         n53644, n53645, n53646, n53647, n53648, n53649, n53650, n53651,
         n53652, n53653, n53654, n53655, n53656, n53657, n53658, n53659,
         n53660, n53661, n53662, n53663, n53664, n53665, n53666, n53667,
         n53668, n53669, n53670, n53671, n53672, n53673, n53674, n53675,
         n53676, n53677, n53678, n53679, n53680, n53681, n53682, n53683,
         n53684, n53685, n53686, n53687, n53688, n53689, n53690, n53691,
         n53692, n53693, n53694, n53695, n53696, n53697, n53698, n53699,
         n53700, n53701, n53702, n53703, n53704, n53705, n53706, n53707,
         n53708, n53709, n53710, n53711, n53712, n53713, n53714, n53715,
         n53716, n53717, n53718, n53719, n53720, n53721, n53722, n53723,
         n53724, n53725, n53726, n53727, n53728, n53729, n53730, n53731,
         n53732, n53733, n53734, n53735, n53736, n53737, n53738, n53739,
         n53740, n53741, n53742, n53743, n53744, n53745, n53746, n53747,
         n53748, n53749, n53750, n53751, n53752, n53753, n53754, n53755,
         n53756, n53757, n53758, n53759, n53760, n53761, n53762, n53763,
         n53764, n53765, n53766, n53767, n53768, n53769, n53770, n53771,
         n53772, n53773, n53774, n53775, n53776, n53777, n53778, n53779,
         n53780, n53781, n53782, n53783, n53784, n53785, n53786, n53787,
         n53788, n53789, n53790, n53791, n53792, n53793, n53794, n53795,
         n53796, n53797, n53798, n53799, n53800, n53801, n53802, n53803,
         n53804, n53805, n53806, n53807, n53808, n53809, n53810, n53811,
         n53812, n53813, n53814, n53815, n53816, n53817, n53818, n53819,
         n53820, n53821, n53822, n53823, n53824, n53825, n53826, n53827,
         n53828, n53829, n53830, n53831, n53832, n53833, n53834, n53835,
         n53836, n53837, n53838, n53839, n53840, n53841, n53842, n53843,
         n53844, n53845, n53846, n53847, n53848, n53849, n53850, n53851,
         n53852, n53853, n53854, n53855, n53856, n53857, n53858, n53859,
         n53860, n53861, n53862, n53863, n53864, n53865, n53866, n53867,
         n53868, n53869, n53870, n53871, n53872, n53873, n53874, n53875,
         n53876, n53877, n53878, n53879, n53880, n53881, n53882, n53883,
         n53884, n53885, n53886, n53887, n53888, n53889, n53890, n53891,
         n53892, n53893, n53894, n53895, n53896, n53897, n53898, n53899,
         n53900, n53901, n53902, n53903, n53904, n53905, n53906, n53907,
         n53908, n53909, n53910, n53911, n53912, n53913, n53914, n53915,
         n53916, n53917, n53918, n53919, n53920, n53921, n53922, n53923,
         n53924, n53925, n53926, n53927, n53928, n53929, n53930, n53931,
         n53932, n53933, n53934, n53935, n53936, n53937, n53938, n53939,
         n53940, n53941, n53942, n53943, n53944, n53945, n53946, n53947,
         n53948, n53949, n53950, n53951, n53952, n53953, n53954, n53955,
         n53956, n53957, n53958, n53959, n53960, n53961, n53962, n53963,
         n53964, n53965, n53966, n53967, n53968, n53969, n53970, n53971,
         n53972, n53973, n53974, n53975, n53976, n53977, n53978, n53979,
         n53980, n53981, n53982, n53983, n53984, n53985, n53986, n53987,
         n53988, n53989, n53990, n53991, n53992, n53993, n53994, n53995,
         n53996, n53997, n53998;
  wire   [12:0] olocal;
  wire   [13:0] oglobal;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131, 
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, SYNOPSYS_UNCONNECTED__137, 
        SYNOPSYS_UNCONNECTED__138, SYNOPSYS_UNCONNECTED__139, 
        SYNOPSYS_UNCONNECTED__140, SYNOPSYS_UNCONNECTED__141, 
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, SYNOPSYS_UNCONNECTED__147, 
        SYNOPSYS_UNCONNECTED__148, SYNOPSYS_UNCONNECTED__149, 
        SYNOPSYS_UNCONNECTED__150, SYNOPSYS_UNCONNECTED__151, 
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, SYNOPSYS_UNCONNECTED__157, 
        SYNOPSYS_UNCONNECTED__158, SYNOPSYS_UNCONNECTED__159, 
        SYNOPSYS_UNCONNECTED__160, SYNOPSYS_UNCONNECTED__161, 
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, SYNOPSYS_UNCONNECTED__167, 
        SYNOPSYS_UNCONNECTED__168, SYNOPSYS_UNCONNECTED__169, 
        SYNOPSYS_UNCONNECTED__170, SYNOPSYS_UNCONNECTED__171, 
        SYNOPSYS_UNCONNECTED__172, SYNOPSYS_UNCONNECTED__173, 
        SYNOPSYS_UNCONNECTED__174, SYNOPSYS_UNCONNECTED__175, 
        SYNOPSYS_UNCONNECTED__176, SYNOPSYS_UNCONNECTED__177, 
        SYNOPSYS_UNCONNECTED__178, SYNOPSYS_UNCONNECTED__179, 
        SYNOPSYS_UNCONNECTED__180, SYNOPSYS_UNCONNECTED__181, 
        SYNOPSYS_UNCONNECTED__182, SYNOPSYS_UNCONNECTED__183, 
        SYNOPSYS_UNCONNECTED__184, SYNOPSYS_UNCONNECTED__185, 
        SYNOPSYS_UNCONNECTED__186, SYNOPSYS_UNCONNECTED__187, 
        SYNOPSYS_UNCONNECTED__188, SYNOPSYS_UNCONNECTED__189, 
        SYNOPSYS_UNCONNECTED__190, SYNOPSYS_UNCONNECTED__191, 
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, SYNOPSYS_UNCONNECTED__197, 
        SYNOPSYS_UNCONNECTED__198, SYNOPSYS_UNCONNECTED__199, 
        SYNOPSYS_UNCONNECTED__200, SYNOPSYS_UNCONNECTED__201, 
        SYNOPSYS_UNCONNECTED__202, SYNOPSYS_UNCONNECTED__203, 
        SYNOPSYS_UNCONNECTED__204, SYNOPSYS_UNCONNECTED__205, 
        SYNOPSYS_UNCONNECTED__206, SYNOPSYS_UNCONNECTED__207, 
        SYNOPSYS_UNCONNECTED__208, SYNOPSYS_UNCONNECTED__209, 
        SYNOPSYS_UNCONNECTED__210, SYNOPSYS_UNCONNECTED__211, 
        SYNOPSYS_UNCONNECTED__212, SYNOPSYS_UNCONNECTED__213, 
        SYNOPSYS_UNCONNECTED__214, SYNOPSYS_UNCONNECTED__215, 
        SYNOPSYS_UNCONNECTED__216, SYNOPSYS_UNCONNECTED__217, 
        SYNOPSYS_UNCONNECTED__218, SYNOPSYS_UNCONNECTED__219, 
        SYNOPSYS_UNCONNECTED__220, SYNOPSYS_UNCONNECTED__221, 
        SYNOPSYS_UNCONNECTED__222, SYNOPSYS_UNCONNECTED__223, 
        SYNOPSYS_UNCONNECTED__224, SYNOPSYS_UNCONNECTED__225, 
        SYNOPSYS_UNCONNECTED__226, SYNOPSYS_UNCONNECTED__227, 
        SYNOPSYS_UNCONNECTED__228, SYNOPSYS_UNCONNECTED__229, 
        SYNOPSYS_UNCONNECTED__230, SYNOPSYS_UNCONNECTED__231, 
        SYNOPSYS_UNCONNECTED__232, SYNOPSYS_UNCONNECTED__233, 
        SYNOPSYS_UNCONNECTED__234, SYNOPSYS_UNCONNECTED__235, 
        SYNOPSYS_UNCONNECTED__236, SYNOPSYS_UNCONNECTED__237, 
        SYNOPSYS_UNCONNECTED__238, SYNOPSYS_UNCONNECTED__239, 
        SYNOPSYS_UNCONNECTED__240, SYNOPSYS_UNCONNECTED__241, 
        SYNOPSYS_UNCONNECTED__242, SYNOPSYS_UNCONNECTED__243, 
        SYNOPSYS_UNCONNECTED__244, SYNOPSYS_UNCONNECTED__245, 
        SYNOPSYS_UNCONNECTED__246, SYNOPSYS_UNCONNECTED__247, 
        SYNOPSYS_UNCONNECTED__248, SYNOPSYS_UNCONNECTED__249, 
        SYNOPSYS_UNCONNECTED__250, SYNOPSYS_UNCONNECTED__251, 
        SYNOPSYS_UNCONNECTED__252, SYNOPSYS_UNCONNECTED__253, 
        SYNOPSYS_UNCONNECTED__254, SYNOPSYS_UNCONNECTED__255, 
        SYNOPSYS_UNCONNECTED__256, SYNOPSYS_UNCONNECTED__257, 
        SYNOPSYS_UNCONNECTED__258, SYNOPSYS_UNCONNECTED__259, 
        SYNOPSYS_UNCONNECTED__260, SYNOPSYS_UNCONNECTED__261, 
        SYNOPSYS_UNCONNECTED__262, SYNOPSYS_UNCONNECTED__263, 
        SYNOPSYS_UNCONNECTED__264, SYNOPSYS_UNCONNECTED__265, 
        SYNOPSYS_UNCONNECTED__266, SYNOPSYS_UNCONNECTED__267, 
        SYNOPSYS_UNCONNECTED__268, SYNOPSYS_UNCONNECTED__269, 
        SYNOPSYS_UNCONNECTED__270, SYNOPSYS_UNCONNECTED__271, 
        SYNOPSYS_UNCONNECTED__272, SYNOPSYS_UNCONNECTED__273, 
        SYNOPSYS_UNCONNECTED__274, SYNOPSYS_UNCONNECTED__275, 
        SYNOPSYS_UNCONNECTED__276, SYNOPSYS_UNCONNECTED__277, 
        SYNOPSYS_UNCONNECTED__278, SYNOPSYS_UNCONNECTED__279, 
        SYNOPSYS_UNCONNECTED__280, SYNOPSYS_UNCONNECTED__281, 
        SYNOPSYS_UNCONNECTED__282, SYNOPSYS_UNCONNECTED__283, 
        SYNOPSYS_UNCONNECTED__284, SYNOPSYS_UNCONNECTED__285, 
        SYNOPSYS_UNCONNECTED__286, SYNOPSYS_UNCONNECTED__287, 
        SYNOPSYS_UNCONNECTED__288, SYNOPSYS_UNCONNECTED__289, 
        SYNOPSYS_UNCONNECTED__290, SYNOPSYS_UNCONNECTED__291, 
        SYNOPSYS_UNCONNECTED__292, SYNOPSYS_UNCONNECTED__293, 
        SYNOPSYS_UNCONNECTED__294, SYNOPSYS_UNCONNECTED__295, 
        SYNOPSYS_UNCONNECTED__296, SYNOPSYS_UNCONNECTED__297, 
        SYNOPSYS_UNCONNECTED__298, SYNOPSYS_UNCONNECTED__299, 
        SYNOPSYS_UNCONNECTED__300, SYNOPSYS_UNCONNECTED__301, 
        SYNOPSYS_UNCONNECTED__302, SYNOPSYS_UNCONNECTED__303, 
        SYNOPSYS_UNCONNECTED__304, SYNOPSYS_UNCONNECTED__305, 
        SYNOPSYS_UNCONNECTED__306, SYNOPSYS_UNCONNECTED__307, 
        SYNOPSYS_UNCONNECTED__308, SYNOPSYS_UNCONNECTED__309, 
        SYNOPSYS_UNCONNECTED__310, SYNOPSYS_UNCONNECTED__311, 
        SYNOPSYS_UNCONNECTED__312, SYNOPSYS_UNCONNECTED__313, 
        SYNOPSYS_UNCONNECTED__314, SYNOPSYS_UNCONNECTED__315, 
        SYNOPSYS_UNCONNECTED__316, SYNOPSYS_UNCONNECTED__317, 
        SYNOPSYS_UNCONNECTED__318, SYNOPSYS_UNCONNECTED__319, 
        SYNOPSYS_UNCONNECTED__320, SYNOPSYS_UNCONNECTED__321, 
        SYNOPSYS_UNCONNECTED__322, SYNOPSYS_UNCONNECTED__323, 
        SYNOPSYS_UNCONNECTED__324, SYNOPSYS_UNCONNECTED__325, 
        SYNOPSYS_UNCONNECTED__326, SYNOPSYS_UNCONNECTED__327, 
        SYNOPSYS_UNCONNECTED__328, SYNOPSYS_UNCONNECTED__329, 
        SYNOPSYS_UNCONNECTED__330, SYNOPSYS_UNCONNECTED__331, 
        SYNOPSYS_UNCONNECTED__332, SYNOPSYS_UNCONNECTED__333, 
        SYNOPSYS_UNCONNECTED__334, SYNOPSYS_UNCONNECTED__335, 
        SYNOPSYS_UNCONNECTED__336, SYNOPSYS_UNCONNECTED__337, 
        SYNOPSYS_UNCONNECTED__338, SYNOPSYS_UNCONNECTED__339, 
        SYNOPSYS_UNCONNECTED__340, SYNOPSYS_UNCONNECTED__341, 
        SYNOPSYS_UNCONNECTED__342, SYNOPSYS_UNCONNECTED__343, 
        SYNOPSYS_UNCONNECTED__344, SYNOPSYS_UNCONNECTED__345, 
        SYNOPSYS_UNCONNECTED__346, SYNOPSYS_UNCONNECTED__347, 
        SYNOPSYS_UNCONNECTED__348, SYNOPSYS_UNCONNECTED__349, 
        SYNOPSYS_UNCONNECTED__350, SYNOPSYS_UNCONNECTED__351, 
        SYNOPSYS_UNCONNECTED__352, SYNOPSYS_UNCONNECTED__353, 
        SYNOPSYS_UNCONNECTED__354, SYNOPSYS_UNCONNECTED__355, 
        SYNOPSYS_UNCONNECTED__356, SYNOPSYS_UNCONNECTED__357, 
        SYNOPSYS_UNCONNECTED__358, SYNOPSYS_UNCONNECTED__359, 
        SYNOPSYS_UNCONNECTED__360, SYNOPSYS_UNCONNECTED__361, 
        SYNOPSYS_UNCONNECTED__362, SYNOPSYS_UNCONNECTED__363, 
        SYNOPSYS_UNCONNECTED__364, SYNOPSYS_UNCONNECTED__365, 
        SYNOPSYS_UNCONNECTED__366, SYNOPSYS_UNCONNECTED__367, 
        SYNOPSYS_UNCONNECTED__368, SYNOPSYS_UNCONNECTED__369, 
        SYNOPSYS_UNCONNECTED__370, SYNOPSYS_UNCONNECTED__371, 
        SYNOPSYS_UNCONNECTED__372, SYNOPSYS_UNCONNECTED__373, 
        SYNOPSYS_UNCONNECTED__374, SYNOPSYS_UNCONNECTED__375, 
        SYNOPSYS_UNCONNECTED__376, SYNOPSYS_UNCONNECTED__377, 
        SYNOPSYS_UNCONNECTED__378, SYNOPSYS_UNCONNECTED__379, 
        SYNOPSYS_UNCONNECTED__380, SYNOPSYS_UNCONNECTED__381, 
        SYNOPSYS_UNCONNECTED__382, SYNOPSYS_UNCONNECTED__383, 
        SYNOPSYS_UNCONNECTED__384, SYNOPSYS_UNCONNECTED__385, 
        SYNOPSYS_UNCONNECTED__386, SYNOPSYS_UNCONNECTED__387, 
        SYNOPSYS_UNCONNECTED__388, SYNOPSYS_UNCONNECTED__389, 
        SYNOPSYS_UNCONNECTED__390, SYNOPSYS_UNCONNECTED__391, 
        SYNOPSYS_UNCONNECTED__392, SYNOPSYS_UNCONNECTED__393, 
        SYNOPSYS_UNCONNECTED__394, SYNOPSYS_UNCONNECTED__395, 
        SYNOPSYS_UNCONNECTED__396, SYNOPSYS_UNCONNECTED__397, 
        SYNOPSYS_UNCONNECTED__398, SYNOPSYS_UNCONNECTED__399, 
        SYNOPSYS_UNCONNECTED__400, SYNOPSYS_UNCONNECTED__401, 
        SYNOPSYS_UNCONNECTED__402, SYNOPSYS_UNCONNECTED__403, 
        SYNOPSYS_UNCONNECTED__404, SYNOPSYS_UNCONNECTED__405, 
        SYNOPSYS_UNCONNECTED__406, SYNOPSYS_UNCONNECTED__407, 
        SYNOPSYS_UNCONNECTED__408, SYNOPSYS_UNCONNECTED__409, 
        SYNOPSYS_UNCONNECTED__410, SYNOPSYS_UNCONNECTED__411, 
        SYNOPSYS_UNCONNECTED__412, SYNOPSYS_UNCONNECTED__413, 
        SYNOPSYS_UNCONNECTED__414, SYNOPSYS_UNCONNECTED__415, 
        SYNOPSYS_UNCONNECTED__416, SYNOPSYS_UNCONNECTED__417, 
        SYNOPSYS_UNCONNECTED__418, SYNOPSYS_UNCONNECTED__419, 
        SYNOPSYS_UNCONNECTED__420, SYNOPSYS_UNCONNECTED__421, 
        SYNOPSYS_UNCONNECTED__422, SYNOPSYS_UNCONNECTED__423, 
        SYNOPSYS_UNCONNECTED__424, SYNOPSYS_UNCONNECTED__425, 
        SYNOPSYS_UNCONNECTED__426, SYNOPSYS_UNCONNECTED__427, 
        SYNOPSYS_UNCONNECTED__428, SYNOPSYS_UNCONNECTED__429, 
        SYNOPSYS_UNCONNECTED__430, SYNOPSYS_UNCONNECTED__431, 
        SYNOPSYS_UNCONNECTED__432, SYNOPSYS_UNCONNECTED__433, 
        SYNOPSYS_UNCONNECTED__434, SYNOPSYS_UNCONNECTED__435, 
        SYNOPSYS_UNCONNECTED__436, SYNOPSYS_UNCONNECTED__437, 
        SYNOPSYS_UNCONNECTED__438, SYNOPSYS_UNCONNECTED__439, 
        SYNOPSYS_UNCONNECTED__440, SYNOPSYS_UNCONNECTED__441, 
        SYNOPSYS_UNCONNECTED__442, SYNOPSYS_UNCONNECTED__443, 
        SYNOPSYS_UNCONNECTED__444, SYNOPSYS_UNCONNECTED__445, 
        SYNOPSYS_UNCONNECTED__446, SYNOPSYS_UNCONNECTED__447, 
        SYNOPSYS_UNCONNECTED__448, SYNOPSYS_UNCONNECTED__449, 
        SYNOPSYS_UNCONNECTED__450, SYNOPSYS_UNCONNECTED__451, 
        SYNOPSYS_UNCONNECTED__452, SYNOPSYS_UNCONNECTED__453, 
        SYNOPSYS_UNCONNECTED__454, SYNOPSYS_UNCONNECTED__455, 
        SYNOPSYS_UNCONNECTED__456, SYNOPSYS_UNCONNECTED__457, 
        SYNOPSYS_UNCONNECTED__458, SYNOPSYS_UNCONNECTED__459, 
        SYNOPSYS_UNCONNECTED__460, SYNOPSYS_UNCONNECTED__461, 
        SYNOPSYS_UNCONNECTED__462, SYNOPSYS_UNCONNECTED__463, 
        SYNOPSYS_UNCONNECTED__464, SYNOPSYS_UNCONNECTED__465, 
        SYNOPSYS_UNCONNECTED__466, SYNOPSYS_UNCONNECTED__467, 
        SYNOPSYS_UNCONNECTED__468, SYNOPSYS_UNCONNECTED__469, 
        SYNOPSYS_UNCONNECTED__470, SYNOPSYS_UNCONNECTED__471, 
        SYNOPSYS_UNCONNECTED__472, SYNOPSYS_UNCONNECTED__473, 
        SYNOPSYS_UNCONNECTED__474, SYNOPSYS_UNCONNECTED__475, 
        SYNOPSYS_UNCONNECTED__476, SYNOPSYS_UNCONNECTED__477, 
        SYNOPSYS_UNCONNECTED__478, SYNOPSYS_UNCONNECTED__479, 
        SYNOPSYS_UNCONNECTED__480, SYNOPSYS_UNCONNECTED__481, 
        SYNOPSYS_UNCONNECTED__482, SYNOPSYS_UNCONNECTED__483, 
        SYNOPSYS_UNCONNECTED__484, SYNOPSYS_UNCONNECTED__485, 
        SYNOPSYS_UNCONNECTED__486, SYNOPSYS_UNCONNECTED__487, 
        SYNOPSYS_UNCONNECTED__488, SYNOPSYS_UNCONNECTED__489, 
        SYNOPSYS_UNCONNECTED__490, SYNOPSYS_UNCONNECTED__491, 
        SYNOPSYS_UNCONNECTED__492, SYNOPSYS_UNCONNECTED__493, 
        SYNOPSYS_UNCONNECTED__494, SYNOPSYS_UNCONNECTED__495, 
        SYNOPSYS_UNCONNECTED__496, SYNOPSYS_UNCONNECTED__497, 
        SYNOPSYS_UNCONNECTED__498, SYNOPSYS_UNCONNECTED__499, 
        SYNOPSYS_UNCONNECTED__500, SYNOPSYS_UNCONNECTED__501, 
        SYNOPSYS_UNCONNECTED__502, SYNOPSYS_UNCONNECTED__503, 
        SYNOPSYS_UNCONNECTED__504, SYNOPSYS_UNCONNECTED__505, 
        SYNOPSYS_UNCONNECTED__506, SYNOPSYS_UNCONNECTED__507, 
        SYNOPSYS_UNCONNECTED__508, SYNOPSYS_UNCONNECTED__509, 
        SYNOPSYS_UNCONNECTED__510, SYNOPSYS_UNCONNECTED__511, 
        SYNOPSYS_UNCONNECTED__512, SYNOPSYS_UNCONNECTED__513, 
        SYNOPSYS_UNCONNECTED__514, SYNOPSYS_UNCONNECTED__515, 
        SYNOPSYS_UNCONNECTED__516, SYNOPSYS_UNCONNECTED__517, 
        SYNOPSYS_UNCONNECTED__518, SYNOPSYS_UNCONNECTED__519, 
        SYNOPSYS_UNCONNECTED__520, SYNOPSYS_UNCONNECTED__521, 
        SYNOPSYS_UNCONNECTED__522, SYNOPSYS_UNCONNECTED__523, 
        SYNOPSYS_UNCONNECTED__524, SYNOPSYS_UNCONNECTED__525, 
        SYNOPSYS_UNCONNECTED__526, SYNOPSYS_UNCONNECTED__527, 
        SYNOPSYS_UNCONNECTED__528, SYNOPSYS_UNCONNECTED__529, 
        SYNOPSYS_UNCONNECTED__530, SYNOPSYS_UNCONNECTED__531, 
        SYNOPSYS_UNCONNECTED__532, SYNOPSYS_UNCONNECTED__533, 
        SYNOPSYS_UNCONNECTED__534, SYNOPSYS_UNCONNECTED__535, 
        SYNOPSYS_UNCONNECTED__536, SYNOPSYS_UNCONNECTED__537, 
        SYNOPSYS_UNCONNECTED__538, SYNOPSYS_UNCONNECTED__539, 
        SYNOPSYS_UNCONNECTED__540, SYNOPSYS_UNCONNECTED__541, 
        SYNOPSYS_UNCONNECTED__542, SYNOPSYS_UNCONNECTED__543, 
        SYNOPSYS_UNCONNECTED__544, SYNOPSYS_UNCONNECTED__545, 
        SYNOPSYS_UNCONNECTED__546, SYNOPSYS_UNCONNECTED__547, 
        SYNOPSYS_UNCONNECTED__548, SYNOPSYS_UNCONNECTED__549, 
        SYNOPSYS_UNCONNECTED__550, SYNOPSYS_UNCONNECTED__551, 
        SYNOPSYS_UNCONNECTED__552, SYNOPSYS_UNCONNECTED__553, 
        SYNOPSYS_UNCONNECTED__554, SYNOPSYS_UNCONNECTED__555, 
        SYNOPSYS_UNCONNECTED__556, SYNOPSYS_UNCONNECTED__557, 
        SYNOPSYS_UNCONNECTED__558, SYNOPSYS_UNCONNECTED__559, 
        SYNOPSYS_UNCONNECTED__560, SYNOPSYS_UNCONNECTED__561, 
        SYNOPSYS_UNCONNECTED__562, SYNOPSYS_UNCONNECTED__563, 
        SYNOPSYS_UNCONNECTED__564, SYNOPSYS_UNCONNECTED__565, 
        SYNOPSYS_UNCONNECTED__566, SYNOPSYS_UNCONNECTED__567, 
        SYNOPSYS_UNCONNECTED__568, SYNOPSYS_UNCONNECTED__569, 
        SYNOPSYS_UNCONNECTED__570, SYNOPSYS_UNCONNECTED__571, 
        SYNOPSYS_UNCONNECTED__572, SYNOPSYS_UNCONNECTED__573, 
        SYNOPSYS_UNCONNECTED__574, SYNOPSYS_UNCONNECTED__575, 
        SYNOPSYS_UNCONNECTED__576, SYNOPSYS_UNCONNECTED__577, 
        SYNOPSYS_UNCONNECTED__578, SYNOPSYS_UNCONNECTED__579, 
        SYNOPSYS_UNCONNECTED__580, SYNOPSYS_UNCONNECTED__581, 
        SYNOPSYS_UNCONNECTED__582, SYNOPSYS_UNCONNECTED__583, 
        SYNOPSYS_UNCONNECTED__584, SYNOPSYS_UNCONNECTED__585, 
        SYNOPSYS_UNCONNECTED__586, SYNOPSYS_UNCONNECTED__587, 
        SYNOPSYS_UNCONNECTED__588, SYNOPSYS_UNCONNECTED__589, 
        SYNOPSYS_UNCONNECTED__590, SYNOPSYS_UNCONNECTED__591, 
        SYNOPSYS_UNCONNECTED__592, SYNOPSYS_UNCONNECTED__593, 
        SYNOPSYS_UNCONNECTED__594, SYNOPSYS_UNCONNECTED__595, 
        SYNOPSYS_UNCONNECTED__596, SYNOPSYS_UNCONNECTED__597, 
        SYNOPSYS_UNCONNECTED__598, SYNOPSYS_UNCONNECTED__599, 
        SYNOPSYS_UNCONNECTED__600, SYNOPSYS_UNCONNECTED__601, 
        SYNOPSYS_UNCONNECTED__602, SYNOPSYS_UNCONNECTED__603, 
        SYNOPSYS_UNCONNECTED__604, SYNOPSYS_UNCONNECTED__605, 
        SYNOPSYS_UNCONNECTED__606, SYNOPSYS_UNCONNECTED__607, 
        SYNOPSYS_UNCONNECTED__608, SYNOPSYS_UNCONNECTED__609, 
        SYNOPSYS_UNCONNECTED__610, SYNOPSYS_UNCONNECTED__611, 
        SYNOPSYS_UNCONNECTED__612, SYNOPSYS_UNCONNECTED__613, 
        SYNOPSYS_UNCONNECTED__614, SYNOPSYS_UNCONNECTED__615, 
        SYNOPSYS_UNCONNECTED__616, SYNOPSYS_UNCONNECTED__617, 
        SYNOPSYS_UNCONNECTED__618, SYNOPSYS_UNCONNECTED__619, 
        SYNOPSYS_UNCONNECTED__620, SYNOPSYS_UNCONNECTED__621, 
        SYNOPSYS_UNCONNECTED__622, SYNOPSYS_UNCONNECTED__623, 
        SYNOPSYS_UNCONNECTED__624, SYNOPSYS_UNCONNECTED__625, 
        SYNOPSYS_UNCONNECTED__626, SYNOPSYS_UNCONNECTED__627, 
        SYNOPSYS_UNCONNECTED__628, SYNOPSYS_UNCONNECTED__629, 
        SYNOPSYS_UNCONNECTED__630, SYNOPSYS_UNCONNECTED__631, 
        SYNOPSYS_UNCONNECTED__632, SYNOPSYS_UNCONNECTED__633, 
        SYNOPSYS_UNCONNECTED__634, SYNOPSYS_UNCONNECTED__635, 
        SYNOPSYS_UNCONNECTED__636, SYNOPSYS_UNCONNECTED__637, 
        SYNOPSYS_UNCONNECTED__638, SYNOPSYS_UNCONNECTED__639, 
        SYNOPSYS_UNCONNECTED__640, SYNOPSYS_UNCONNECTED__641, 
        SYNOPSYS_UNCONNECTED__642, SYNOPSYS_UNCONNECTED__643, 
        SYNOPSYS_UNCONNECTED__644, SYNOPSYS_UNCONNECTED__645, 
        SYNOPSYS_UNCONNECTED__646, SYNOPSYS_UNCONNECTED__647, 
        SYNOPSYS_UNCONNECTED__648, SYNOPSYS_UNCONNECTED__649, 
        SYNOPSYS_UNCONNECTED__650, SYNOPSYS_UNCONNECTED__651, 
        SYNOPSYS_UNCONNECTED__652, SYNOPSYS_UNCONNECTED__653, 
        SYNOPSYS_UNCONNECTED__654, SYNOPSYS_UNCONNECTED__655, 
        SYNOPSYS_UNCONNECTED__656, SYNOPSYS_UNCONNECTED__657, 
        SYNOPSYS_UNCONNECTED__658, SYNOPSYS_UNCONNECTED__659, 
        SYNOPSYS_UNCONNECTED__660, SYNOPSYS_UNCONNECTED__661, 
        SYNOPSYS_UNCONNECTED__662, SYNOPSYS_UNCONNECTED__663, 
        SYNOPSYS_UNCONNECTED__664, SYNOPSYS_UNCONNECTED__665, 
        SYNOPSYS_UNCONNECTED__666, SYNOPSYS_UNCONNECTED__667, 
        SYNOPSYS_UNCONNECTED__668, SYNOPSYS_UNCONNECTED__669, 
        SYNOPSYS_UNCONNECTED__670, SYNOPSYS_UNCONNECTED__671, 
        SYNOPSYS_UNCONNECTED__672, SYNOPSYS_UNCONNECTED__673, 
        SYNOPSYS_UNCONNECTED__674, SYNOPSYS_UNCONNECTED__675, 
        SYNOPSYS_UNCONNECTED__676, SYNOPSYS_UNCONNECTED__677, 
        SYNOPSYS_UNCONNECTED__678, SYNOPSYS_UNCONNECTED__679, 
        SYNOPSYS_UNCONNECTED__680, SYNOPSYS_UNCONNECTED__681, 
        SYNOPSYS_UNCONNECTED__682, SYNOPSYS_UNCONNECTED__683, 
        SYNOPSYS_UNCONNECTED__684, SYNOPSYS_UNCONNECTED__685, 
        SYNOPSYS_UNCONNECTED__686, SYNOPSYS_UNCONNECTED__687, 
        SYNOPSYS_UNCONNECTED__688, SYNOPSYS_UNCONNECTED__689, 
        SYNOPSYS_UNCONNECTED__690, SYNOPSYS_UNCONNECTED__691, 
        SYNOPSYS_UNCONNECTED__692, SYNOPSYS_UNCONNECTED__693, 
        SYNOPSYS_UNCONNECTED__694, SYNOPSYS_UNCONNECTED__695, 
        SYNOPSYS_UNCONNECTED__696, SYNOPSYS_UNCONNECTED__697, 
        SYNOPSYS_UNCONNECTED__698, SYNOPSYS_UNCONNECTED__699, 
        SYNOPSYS_UNCONNECTED__700, SYNOPSYS_UNCONNECTED__701, 
        SYNOPSYS_UNCONNECTED__702, SYNOPSYS_UNCONNECTED__703, 
        SYNOPSYS_UNCONNECTED__704, SYNOPSYS_UNCONNECTED__705, 
        SYNOPSYS_UNCONNECTED__706, SYNOPSYS_UNCONNECTED__707, 
        SYNOPSYS_UNCONNECTED__708, SYNOPSYS_UNCONNECTED__709, 
        SYNOPSYS_UNCONNECTED__710, SYNOPSYS_UNCONNECTED__711, 
        SYNOPSYS_UNCONNECTED__712, SYNOPSYS_UNCONNECTED__713, 
        SYNOPSYS_UNCONNECTED__714, SYNOPSYS_UNCONNECTED__715, 
        SYNOPSYS_UNCONNECTED__716, SYNOPSYS_UNCONNECTED__717, 
        SYNOPSYS_UNCONNECTED__718, SYNOPSYS_UNCONNECTED__719, 
        SYNOPSYS_UNCONNECTED__720, SYNOPSYS_UNCONNECTED__721, 
        SYNOPSYS_UNCONNECTED__722, SYNOPSYS_UNCONNECTED__723, 
        SYNOPSYS_UNCONNECTED__724, SYNOPSYS_UNCONNECTED__725, 
        SYNOPSYS_UNCONNECTED__726, SYNOPSYS_UNCONNECTED__727, 
        SYNOPSYS_UNCONNECTED__728, SYNOPSYS_UNCONNECTED__729, 
        SYNOPSYS_UNCONNECTED__730, SYNOPSYS_UNCONNECTED__731, 
        SYNOPSYS_UNCONNECTED__732, SYNOPSYS_UNCONNECTED__733, 
        SYNOPSYS_UNCONNECTED__734, SYNOPSYS_UNCONNECTED__735, 
        SYNOPSYS_UNCONNECTED__736, SYNOPSYS_UNCONNECTED__737, 
        SYNOPSYS_UNCONNECTED__738, SYNOPSYS_UNCONNECTED__739, 
        SYNOPSYS_UNCONNECTED__740, SYNOPSYS_UNCONNECTED__741, 
        SYNOPSYS_UNCONNECTED__742, SYNOPSYS_UNCONNECTED__743, 
        SYNOPSYS_UNCONNECTED__744, SYNOPSYS_UNCONNECTED__745, 
        SYNOPSYS_UNCONNECTED__746, SYNOPSYS_UNCONNECTED__747, 
        SYNOPSYS_UNCONNECTED__748, SYNOPSYS_UNCONNECTED__749, 
        SYNOPSYS_UNCONNECTED__750, SYNOPSYS_UNCONNECTED__751, 
        SYNOPSYS_UNCONNECTED__752, SYNOPSYS_UNCONNECTED__753, 
        SYNOPSYS_UNCONNECTED__754, SYNOPSYS_UNCONNECTED__755, 
        SYNOPSYS_UNCONNECTED__756, SYNOPSYS_UNCONNECTED__757, 
        SYNOPSYS_UNCONNECTED__758, SYNOPSYS_UNCONNECTED__759, 
        SYNOPSYS_UNCONNECTED__760, SYNOPSYS_UNCONNECTED__761, 
        SYNOPSYS_UNCONNECTED__762, SYNOPSYS_UNCONNECTED__763, 
        SYNOPSYS_UNCONNECTED__764, SYNOPSYS_UNCONNECTED__765, 
        SYNOPSYS_UNCONNECTED__766, SYNOPSYS_UNCONNECTED__767, 
        SYNOPSYS_UNCONNECTED__768, SYNOPSYS_UNCONNECTED__769, 
        SYNOPSYS_UNCONNECTED__770, SYNOPSYS_UNCONNECTED__771, 
        SYNOPSYS_UNCONNECTED__772, SYNOPSYS_UNCONNECTED__773, 
        SYNOPSYS_UNCONNECTED__774, SYNOPSYS_UNCONNECTED__775, 
        SYNOPSYS_UNCONNECTED__776, SYNOPSYS_UNCONNECTED__777, 
        SYNOPSYS_UNCONNECTED__778, SYNOPSYS_UNCONNECTED__779, 
        SYNOPSYS_UNCONNECTED__780, SYNOPSYS_UNCONNECTED__781, 
        SYNOPSYS_UNCONNECTED__782, SYNOPSYS_UNCONNECTED__783, 
        SYNOPSYS_UNCONNECTED__784, SYNOPSYS_UNCONNECTED__785, 
        SYNOPSYS_UNCONNECTED__786, SYNOPSYS_UNCONNECTED__787, 
        SYNOPSYS_UNCONNECTED__788, SYNOPSYS_UNCONNECTED__789, 
        SYNOPSYS_UNCONNECTED__790, SYNOPSYS_UNCONNECTED__791, 
        SYNOPSYS_UNCONNECTED__792, SYNOPSYS_UNCONNECTED__793, 
        SYNOPSYS_UNCONNECTED__794, SYNOPSYS_UNCONNECTED__795, 
        SYNOPSYS_UNCONNECTED__796, SYNOPSYS_UNCONNECTED__797, 
        SYNOPSYS_UNCONNECTED__798, SYNOPSYS_UNCONNECTED__799, 
        SYNOPSYS_UNCONNECTED__800, SYNOPSYS_UNCONNECTED__801, 
        SYNOPSYS_UNCONNECTED__802, SYNOPSYS_UNCONNECTED__803, 
        SYNOPSYS_UNCONNECTED__804, SYNOPSYS_UNCONNECTED__805, 
        SYNOPSYS_UNCONNECTED__806, SYNOPSYS_UNCONNECTED__807, 
        SYNOPSYS_UNCONNECTED__808, SYNOPSYS_UNCONNECTED__809, 
        SYNOPSYS_UNCONNECTED__810, SYNOPSYS_UNCONNECTED__811, 
        SYNOPSYS_UNCONNECTED__812, SYNOPSYS_UNCONNECTED__813, 
        SYNOPSYS_UNCONNECTED__814, SYNOPSYS_UNCONNECTED__815, 
        SYNOPSYS_UNCONNECTED__816, SYNOPSYS_UNCONNECTED__817, 
        SYNOPSYS_UNCONNECTED__818, SYNOPSYS_UNCONNECTED__819, 
        SYNOPSYS_UNCONNECTED__820, SYNOPSYS_UNCONNECTED__821, 
        SYNOPSYS_UNCONNECTED__822, SYNOPSYS_UNCONNECTED__823, 
        SYNOPSYS_UNCONNECTED__824, SYNOPSYS_UNCONNECTED__825, 
        SYNOPSYS_UNCONNECTED__826, SYNOPSYS_UNCONNECTED__827, 
        SYNOPSYS_UNCONNECTED__828, SYNOPSYS_UNCONNECTED__829, 
        SYNOPSYS_UNCONNECTED__830, SYNOPSYS_UNCONNECTED__831, 
        SYNOPSYS_UNCONNECTED__832, SYNOPSYS_UNCONNECTED__833, 
        SYNOPSYS_UNCONNECTED__834, SYNOPSYS_UNCONNECTED__835, 
        SYNOPSYS_UNCONNECTED__836, SYNOPSYS_UNCONNECTED__837, 
        SYNOPSYS_UNCONNECTED__838, SYNOPSYS_UNCONNECTED__839, 
        SYNOPSYS_UNCONNECTED__840, SYNOPSYS_UNCONNECTED__841, 
        SYNOPSYS_UNCONNECTED__842, SYNOPSYS_UNCONNECTED__843, 
        SYNOPSYS_UNCONNECTED__844, SYNOPSYS_UNCONNECTED__845, 
        SYNOPSYS_UNCONNECTED__846, SYNOPSYS_UNCONNECTED__847, 
        SYNOPSYS_UNCONNECTED__848, SYNOPSYS_UNCONNECTED__849, 
        SYNOPSYS_UNCONNECTED__850, SYNOPSYS_UNCONNECTED__851, 
        SYNOPSYS_UNCONNECTED__852, SYNOPSYS_UNCONNECTED__853, 
        SYNOPSYS_UNCONNECTED__854, SYNOPSYS_UNCONNECTED__855, 
        SYNOPSYS_UNCONNECTED__856, SYNOPSYS_UNCONNECTED__857, 
        SYNOPSYS_UNCONNECTED__858, SYNOPSYS_UNCONNECTED__859, 
        SYNOPSYS_UNCONNECTED__860, SYNOPSYS_UNCONNECTED__861, 
        SYNOPSYS_UNCONNECTED__862, SYNOPSYS_UNCONNECTED__863, 
        SYNOPSYS_UNCONNECTED__864, SYNOPSYS_UNCONNECTED__865, 
        SYNOPSYS_UNCONNECTED__866, SYNOPSYS_UNCONNECTED__867, 
        SYNOPSYS_UNCONNECTED__868, SYNOPSYS_UNCONNECTED__869, 
        SYNOPSYS_UNCONNECTED__870, SYNOPSYS_UNCONNECTED__871, 
        SYNOPSYS_UNCONNECTED__872, SYNOPSYS_UNCONNECTED__873, 
        SYNOPSYS_UNCONNECTED__874, SYNOPSYS_UNCONNECTED__875, 
        SYNOPSYS_UNCONNECTED__876, SYNOPSYS_UNCONNECTED__877, 
        SYNOPSYS_UNCONNECTED__878, SYNOPSYS_UNCONNECTED__879, 
        SYNOPSYS_UNCONNECTED__880, SYNOPSYS_UNCONNECTED__881, 
        SYNOPSYS_UNCONNECTED__882, SYNOPSYS_UNCONNECTED__883, 
        SYNOPSYS_UNCONNECTED__884, SYNOPSYS_UNCONNECTED__885, 
        SYNOPSYS_UNCONNECTED__886, SYNOPSYS_UNCONNECTED__887, 
        SYNOPSYS_UNCONNECTED__888, SYNOPSYS_UNCONNECTED__889, 
        SYNOPSYS_UNCONNECTED__890, SYNOPSYS_UNCONNECTED__891, 
        SYNOPSYS_UNCONNECTED__892, SYNOPSYS_UNCONNECTED__893, 
        SYNOPSYS_UNCONNECTED__894, SYNOPSYS_UNCONNECTED__895, 
        SYNOPSYS_UNCONNECTED__896, SYNOPSYS_UNCONNECTED__897, 
        SYNOPSYS_UNCONNECTED__898, SYNOPSYS_UNCONNECTED__899, 
        SYNOPSYS_UNCONNECTED__900, SYNOPSYS_UNCONNECTED__901, 
        SYNOPSYS_UNCONNECTED__902, SYNOPSYS_UNCONNECTED__903, 
        SYNOPSYS_UNCONNECTED__904, SYNOPSYS_UNCONNECTED__905, 
        SYNOPSYS_UNCONNECTED__906, SYNOPSYS_UNCONNECTED__907, 
        SYNOPSYS_UNCONNECTED__908, SYNOPSYS_UNCONNECTED__909, 
        SYNOPSYS_UNCONNECTED__910, SYNOPSYS_UNCONNECTED__911, 
        SYNOPSYS_UNCONNECTED__912, SYNOPSYS_UNCONNECTED__913, 
        SYNOPSYS_UNCONNECTED__914, SYNOPSYS_UNCONNECTED__915, 
        SYNOPSYS_UNCONNECTED__916, SYNOPSYS_UNCONNECTED__917, 
        SYNOPSYS_UNCONNECTED__918, SYNOPSYS_UNCONNECTED__919, 
        SYNOPSYS_UNCONNECTED__920, SYNOPSYS_UNCONNECTED__921, 
        SYNOPSYS_UNCONNECTED__922, SYNOPSYS_UNCONNECTED__923, 
        SYNOPSYS_UNCONNECTED__924, SYNOPSYS_UNCONNECTED__925, 
        SYNOPSYS_UNCONNECTED__926, SYNOPSYS_UNCONNECTED__927, 
        SYNOPSYS_UNCONNECTED__928, SYNOPSYS_UNCONNECTED__929, 
        SYNOPSYS_UNCONNECTED__930, SYNOPSYS_UNCONNECTED__931, 
        SYNOPSYS_UNCONNECTED__932, SYNOPSYS_UNCONNECTED__933, 
        SYNOPSYS_UNCONNECTED__934, SYNOPSYS_UNCONNECTED__935, 
        SYNOPSYS_UNCONNECTED__936, SYNOPSYS_UNCONNECTED__937, 
        SYNOPSYS_UNCONNECTED__938, SYNOPSYS_UNCONNECTED__939, 
        SYNOPSYS_UNCONNECTED__940, SYNOPSYS_UNCONNECTED__941, 
        SYNOPSYS_UNCONNECTED__942, SYNOPSYS_UNCONNECTED__943, 
        SYNOPSYS_UNCONNECTED__944, SYNOPSYS_UNCONNECTED__945, 
        SYNOPSYS_UNCONNECTED__946, SYNOPSYS_UNCONNECTED__947, 
        SYNOPSYS_UNCONNECTED__948, SYNOPSYS_UNCONNECTED__949, 
        SYNOPSYS_UNCONNECTED__950, SYNOPSYS_UNCONNECTED__951, 
        SYNOPSYS_UNCONNECTED__952, SYNOPSYS_UNCONNECTED__953, 
        SYNOPSYS_UNCONNECTED__954, SYNOPSYS_UNCONNECTED__955, 
        SYNOPSYS_UNCONNECTED__956, SYNOPSYS_UNCONNECTED__957, 
        SYNOPSYS_UNCONNECTED__958, SYNOPSYS_UNCONNECTED__959, 
        SYNOPSYS_UNCONNECTED__960, SYNOPSYS_UNCONNECTED__961, 
        SYNOPSYS_UNCONNECTED__962, SYNOPSYS_UNCONNECTED__963, 
        SYNOPSYS_UNCONNECTED__964, SYNOPSYS_UNCONNECTED__965, 
        SYNOPSYS_UNCONNECTED__966, SYNOPSYS_UNCONNECTED__967, 
        SYNOPSYS_UNCONNECTED__968, SYNOPSYS_UNCONNECTED__969, 
        SYNOPSYS_UNCONNECTED__970, SYNOPSYS_UNCONNECTED__971, 
        SYNOPSYS_UNCONNECTED__972, SYNOPSYS_UNCONNECTED__973, 
        SYNOPSYS_UNCONNECTED__974, SYNOPSYS_UNCONNECTED__975, 
        SYNOPSYS_UNCONNECTED__976, SYNOPSYS_UNCONNECTED__977, 
        SYNOPSYS_UNCONNECTED__978, SYNOPSYS_UNCONNECTED__979, 
        SYNOPSYS_UNCONNECTED__980, SYNOPSYS_UNCONNECTED__981, 
        SYNOPSYS_UNCONNECTED__982, SYNOPSYS_UNCONNECTED__983, 
        SYNOPSYS_UNCONNECTED__984, SYNOPSYS_UNCONNECTED__985, 
        SYNOPSYS_UNCONNECTED__986, SYNOPSYS_UNCONNECTED__987, 
        SYNOPSYS_UNCONNECTED__988, SYNOPSYS_UNCONNECTED__989, 
        SYNOPSYS_UNCONNECTED__990, SYNOPSYS_UNCONNECTED__991, 
        SYNOPSYS_UNCONNECTED__992, SYNOPSYS_UNCONNECTED__993, 
        SYNOPSYS_UNCONNECTED__994, SYNOPSYS_UNCONNECTED__995, 
        SYNOPSYS_UNCONNECTED__996, SYNOPSYS_UNCONNECTED__997, 
        SYNOPSYS_UNCONNECTED__998, SYNOPSYS_UNCONNECTED__999, 
        SYNOPSYS_UNCONNECTED__1000, SYNOPSYS_UNCONNECTED__1001, 
        SYNOPSYS_UNCONNECTED__1002, SYNOPSYS_UNCONNECTED__1003, 
        SYNOPSYS_UNCONNECTED__1004, SYNOPSYS_UNCONNECTED__1005, 
        SYNOPSYS_UNCONNECTED__1006, SYNOPSYS_UNCONNECTED__1007, 
        SYNOPSYS_UNCONNECTED__1008, SYNOPSYS_UNCONNECTED__1009, 
        SYNOPSYS_UNCONNECTED__1010, SYNOPSYS_UNCONNECTED__1011, 
        SYNOPSYS_UNCONNECTED__1012, SYNOPSYS_UNCONNECTED__1013, 
        SYNOPSYS_UNCONNECTED__1014, SYNOPSYS_UNCONNECTED__1015, 
        SYNOPSYS_UNCONNECTED__1016, SYNOPSYS_UNCONNECTED__1017, 
        SYNOPSYS_UNCONNECTED__1018, SYNOPSYS_UNCONNECTED__1019, 
        SYNOPSYS_UNCONNECTED__1020, SYNOPSYS_UNCONNECTED__1021, 
        SYNOPSYS_UNCONNECTED__1022, SYNOPSYS_UNCONNECTED__1023, 
        SYNOPSYS_UNCONNECTED__1024, SYNOPSYS_UNCONNECTED__1025, 
        SYNOPSYS_UNCONNECTED__1026, SYNOPSYS_UNCONNECTED__1027, 
        SYNOPSYS_UNCONNECTED__1028, SYNOPSYS_UNCONNECTED__1029, 
        SYNOPSYS_UNCONNECTED__1030, SYNOPSYS_UNCONNECTED__1031, 
        SYNOPSYS_UNCONNECTED__1032, SYNOPSYS_UNCONNECTED__1033, 
        SYNOPSYS_UNCONNECTED__1034, SYNOPSYS_UNCONNECTED__1035, 
        SYNOPSYS_UNCONNECTED__1036, SYNOPSYS_UNCONNECTED__1037, 
        SYNOPSYS_UNCONNECTED__1038, SYNOPSYS_UNCONNECTED__1039, 
        SYNOPSYS_UNCONNECTED__1040, SYNOPSYS_UNCONNECTED__1041, 
        SYNOPSYS_UNCONNECTED__1042, SYNOPSYS_UNCONNECTED__1043, 
        SYNOPSYS_UNCONNECTED__1044, SYNOPSYS_UNCONNECTED__1045, 
        SYNOPSYS_UNCONNECTED__1046, SYNOPSYS_UNCONNECTED__1047, 
        SYNOPSYS_UNCONNECTED__1048, SYNOPSYS_UNCONNECTED__1049, 
        SYNOPSYS_UNCONNECTED__1050, SYNOPSYS_UNCONNECTED__1051, 
        SYNOPSYS_UNCONNECTED__1052, SYNOPSYS_UNCONNECTED__1053, 
        SYNOPSYS_UNCONNECTED__1054, SYNOPSYS_UNCONNECTED__1055, 
        SYNOPSYS_UNCONNECTED__1056, SYNOPSYS_UNCONNECTED__1057, 
        SYNOPSYS_UNCONNECTED__1058, SYNOPSYS_UNCONNECTED__1059, 
        SYNOPSYS_UNCONNECTED__1060, SYNOPSYS_UNCONNECTED__1061, 
        SYNOPSYS_UNCONNECTED__1062, SYNOPSYS_UNCONNECTED__1063, 
        SYNOPSYS_UNCONNECTED__1064, SYNOPSYS_UNCONNECTED__1065, 
        SYNOPSYS_UNCONNECTED__1066, SYNOPSYS_UNCONNECTED__1067, 
        SYNOPSYS_UNCONNECTED__1068, SYNOPSYS_UNCONNECTED__1069, 
        SYNOPSYS_UNCONNECTED__1070, SYNOPSYS_UNCONNECTED__1071, 
        SYNOPSYS_UNCONNECTED__1072, SYNOPSYS_UNCONNECTED__1073, 
        SYNOPSYS_UNCONNECTED__1074, SYNOPSYS_UNCONNECTED__1075, 
        SYNOPSYS_UNCONNECTED__1076, SYNOPSYS_UNCONNECTED__1077, 
        SYNOPSYS_UNCONNECTED__1078, SYNOPSYS_UNCONNECTED__1079, 
        SYNOPSYS_UNCONNECTED__1080, SYNOPSYS_UNCONNECTED__1081, 
        SYNOPSYS_UNCONNECTED__1082, SYNOPSYS_UNCONNECTED__1083, 
        SYNOPSYS_UNCONNECTED__1084, SYNOPSYS_UNCONNECTED__1085, 
        SYNOPSYS_UNCONNECTED__1086, SYNOPSYS_UNCONNECTED__1087, 
        SYNOPSYS_UNCONNECTED__1088, SYNOPSYS_UNCONNECTED__1089, 
        SYNOPSYS_UNCONNECTED__1090, SYNOPSYS_UNCONNECTED__1091, 
        SYNOPSYS_UNCONNECTED__1092, SYNOPSYS_UNCONNECTED__1093, 
        SYNOPSYS_UNCONNECTED__1094, SYNOPSYS_UNCONNECTED__1095, 
        SYNOPSYS_UNCONNECTED__1096, SYNOPSYS_UNCONNECTED__1097, 
        SYNOPSYS_UNCONNECTED__1098, SYNOPSYS_UNCONNECTED__1099, 
        SYNOPSYS_UNCONNECTED__1100, SYNOPSYS_UNCONNECTED__1101, 
        SYNOPSYS_UNCONNECTED__1102, SYNOPSYS_UNCONNECTED__1103, 
        SYNOPSYS_UNCONNECTED__1104, SYNOPSYS_UNCONNECTED__1105, 
        SYNOPSYS_UNCONNECTED__1106, SYNOPSYS_UNCONNECTED__1107, 
        SYNOPSYS_UNCONNECTED__1108, SYNOPSYS_UNCONNECTED__1109, 
        SYNOPSYS_UNCONNECTED__1110, SYNOPSYS_UNCONNECTED__1111, 
        SYNOPSYS_UNCONNECTED__1112, SYNOPSYS_UNCONNECTED__1113, 
        SYNOPSYS_UNCONNECTED__1114, SYNOPSYS_UNCONNECTED__1115, 
        SYNOPSYS_UNCONNECTED__1116, SYNOPSYS_UNCONNECTED__1117, 
        SYNOPSYS_UNCONNECTED__1118, SYNOPSYS_UNCONNECTED__1119, 
        SYNOPSYS_UNCONNECTED__1120, SYNOPSYS_UNCONNECTED__1121, 
        SYNOPSYS_UNCONNECTED__1122, SYNOPSYS_UNCONNECTED__1123, 
        SYNOPSYS_UNCONNECTED__1124, SYNOPSYS_UNCONNECTED__1125, 
        SYNOPSYS_UNCONNECTED__1126, SYNOPSYS_UNCONNECTED__1127, 
        SYNOPSYS_UNCONNECTED__1128, SYNOPSYS_UNCONNECTED__1129, 
        SYNOPSYS_UNCONNECTED__1130, SYNOPSYS_UNCONNECTED__1131, 
        SYNOPSYS_UNCONNECTED__1132, SYNOPSYS_UNCONNECTED__1133, 
        SYNOPSYS_UNCONNECTED__1134, SYNOPSYS_UNCONNECTED__1135, 
        SYNOPSYS_UNCONNECTED__1136, SYNOPSYS_UNCONNECTED__1137, 
        SYNOPSYS_UNCONNECTED__1138, SYNOPSYS_UNCONNECTED__1139, 
        SYNOPSYS_UNCONNECTED__1140, SYNOPSYS_UNCONNECTED__1141, 
        SYNOPSYS_UNCONNECTED__1142, SYNOPSYS_UNCONNECTED__1143, 
        SYNOPSYS_UNCONNECTED__1144, SYNOPSYS_UNCONNECTED__1145, 
        SYNOPSYS_UNCONNECTED__1146, SYNOPSYS_UNCONNECTED__1147, 
        SYNOPSYS_UNCONNECTED__1148, SYNOPSYS_UNCONNECTED__1149, 
        SYNOPSYS_UNCONNECTED__1150, SYNOPSYS_UNCONNECTED__1151, 
        SYNOPSYS_UNCONNECTED__1152, SYNOPSYS_UNCONNECTED__1153, 
        SYNOPSYS_UNCONNECTED__1154, SYNOPSYS_UNCONNECTED__1155, 
        SYNOPSYS_UNCONNECTED__1156, SYNOPSYS_UNCONNECTED__1157, 
        SYNOPSYS_UNCONNECTED__1158, SYNOPSYS_UNCONNECTED__1159, 
        SYNOPSYS_UNCONNECTED__1160, SYNOPSYS_UNCONNECTED__1161, 
        SYNOPSYS_UNCONNECTED__1162, SYNOPSYS_UNCONNECTED__1163, 
        SYNOPSYS_UNCONNECTED__1164, SYNOPSYS_UNCONNECTED__1165, 
        SYNOPSYS_UNCONNECTED__1166, SYNOPSYS_UNCONNECTED__1167, 
        SYNOPSYS_UNCONNECTED__1168, SYNOPSYS_UNCONNECTED__1169, 
        SYNOPSYS_UNCONNECTED__1170, SYNOPSYS_UNCONNECTED__1171, 
        SYNOPSYS_UNCONNECTED__1172, SYNOPSYS_UNCONNECTED__1173, 
        SYNOPSYS_UNCONNECTED__1174, SYNOPSYS_UNCONNECTED__1175, 
        SYNOPSYS_UNCONNECTED__1176, SYNOPSYS_UNCONNECTED__1177, 
        SYNOPSYS_UNCONNECTED__1178, SYNOPSYS_UNCONNECTED__1179, 
        SYNOPSYS_UNCONNECTED__1180, SYNOPSYS_UNCONNECTED__1181, 
        SYNOPSYS_UNCONNECTED__1182, SYNOPSYS_UNCONNECTED__1183, 
        SYNOPSYS_UNCONNECTED__1184, SYNOPSYS_UNCONNECTED__1185, 
        SYNOPSYS_UNCONNECTED__1186, SYNOPSYS_UNCONNECTED__1187, 
        SYNOPSYS_UNCONNECTED__1188, SYNOPSYS_UNCONNECTED__1189, 
        SYNOPSYS_UNCONNECTED__1190, SYNOPSYS_UNCONNECTED__1191, 
        SYNOPSYS_UNCONNECTED__1192, SYNOPSYS_UNCONNECTED__1193, 
        SYNOPSYS_UNCONNECTED__1194, SYNOPSYS_UNCONNECTED__1195, 
        SYNOPSYS_UNCONNECTED__1196, SYNOPSYS_UNCONNECTED__1197, 
        SYNOPSYS_UNCONNECTED__1198, SYNOPSYS_UNCONNECTED__1199, 
        SYNOPSYS_UNCONNECTED__1200, SYNOPSYS_UNCONNECTED__1201, 
        SYNOPSYS_UNCONNECTED__1202, SYNOPSYS_UNCONNECTED__1203, 
        SYNOPSYS_UNCONNECTED__1204, SYNOPSYS_UNCONNECTED__1205, 
        SYNOPSYS_UNCONNECTED__1206, SYNOPSYS_UNCONNECTED__1207, 
        SYNOPSYS_UNCONNECTED__1208, SYNOPSYS_UNCONNECTED__1209, 
        SYNOPSYS_UNCONNECTED__1210, SYNOPSYS_UNCONNECTED__1211, 
        SYNOPSYS_UNCONNECTED__1212, SYNOPSYS_UNCONNECTED__1213, 
        SYNOPSYS_UNCONNECTED__1214, SYNOPSYS_UNCONNECTED__1215, 
        SYNOPSYS_UNCONNECTED__1216, SYNOPSYS_UNCONNECTED__1217, 
        SYNOPSYS_UNCONNECTED__1218, SYNOPSYS_UNCONNECTED__1219, 
        SYNOPSYS_UNCONNECTED__1220, SYNOPSYS_UNCONNECTED__1221, 
        SYNOPSYS_UNCONNECTED__1222, SYNOPSYS_UNCONNECTED__1223, 
        SYNOPSYS_UNCONNECTED__1224, SYNOPSYS_UNCONNECTED__1225, 
        SYNOPSYS_UNCONNECTED__1226, SYNOPSYS_UNCONNECTED__1227, 
        SYNOPSYS_UNCONNECTED__1228, SYNOPSYS_UNCONNECTED__1229, 
        SYNOPSYS_UNCONNECTED__1230, SYNOPSYS_UNCONNECTED__1231, 
        SYNOPSYS_UNCONNECTED__1232, SYNOPSYS_UNCONNECTED__1233, 
        SYNOPSYS_UNCONNECTED__1234, SYNOPSYS_UNCONNECTED__1235, 
        SYNOPSYS_UNCONNECTED__1236, SYNOPSYS_UNCONNECTED__1237, 
        SYNOPSYS_UNCONNECTED__1238, SYNOPSYS_UNCONNECTED__1239, 
        SYNOPSYS_UNCONNECTED__1240, SYNOPSYS_UNCONNECTED__1241, 
        SYNOPSYS_UNCONNECTED__1242, SYNOPSYS_UNCONNECTED__1243, 
        SYNOPSYS_UNCONNECTED__1244, SYNOPSYS_UNCONNECTED__1245, 
        SYNOPSYS_UNCONNECTED__1246, SYNOPSYS_UNCONNECTED__1247, 
        SYNOPSYS_UNCONNECTED__1248, SYNOPSYS_UNCONNECTED__1249, 
        SYNOPSYS_UNCONNECTED__1250, SYNOPSYS_UNCONNECTED__1251, 
        SYNOPSYS_UNCONNECTED__1252, SYNOPSYS_UNCONNECTED__1253, 
        SYNOPSYS_UNCONNECTED__1254, SYNOPSYS_UNCONNECTED__1255, 
        SYNOPSYS_UNCONNECTED__1256, SYNOPSYS_UNCONNECTED__1257, 
        SYNOPSYS_UNCONNECTED__1258, SYNOPSYS_UNCONNECTED__1259, 
        SYNOPSYS_UNCONNECTED__1260, SYNOPSYS_UNCONNECTED__1261, 
        SYNOPSYS_UNCONNECTED__1262, SYNOPSYS_UNCONNECTED__1263, 
        SYNOPSYS_UNCONNECTED__1264, SYNOPSYS_UNCONNECTED__1265, 
        SYNOPSYS_UNCONNECTED__1266, SYNOPSYS_UNCONNECTED__1267, 
        SYNOPSYS_UNCONNECTED__1268, SYNOPSYS_UNCONNECTED__1269, 
        SYNOPSYS_UNCONNECTED__1270, SYNOPSYS_UNCONNECTED__1271, 
        SYNOPSYS_UNCONNECTED__1272, SYNOPSYS_UNCONNECTED__1273, 
        SYNOPSYS_UNCONNECTED__1274, SYNOPSYS_UNCONNECTED__1275, 
        SYNOPSYS_UNCONNECTED__1276, SYNOPSYS_UNCONNECTED__1277, 
        SYNOPSYS_UNCONNECTED__1278, SYNOPSYS_UNCONNECTED__1279, 
        SYNOPSYS_UNCONNECTED__1280, SYNOPSYS_UNCONNECTED__1281, 
        SYNOPSYS_UNCONNECTED__1282, SYNOPSYS_UNCONNECTED__1283, 
        SYNOPSYS_UNCONNECTED__1284, SYNOPSYS_UNCONNECTED__1285, 
        SYNOPSYS_UNCONNECTED__1286, SYNOPSYS_UNCONNECTED__1287, 
        SYNOPSYS_UNCONNECTED__1288, SYNOPSYS_UNCONNECTED__1289, 
        SYNOPSYS_UNCONNECTED__1290, SYNOPSYS_UNCONNECTED__1291, 
        SYNOPSYS_UNCONNECTED__1292, SYNOPSYS_UNCONNECTED__1293, 
        SYNOPSYS_UNCONNECTED__1294, SYNOPSYS_UNCONNECTED__1295, 
        SYNOPSYS_UNCONNECTED__1296, SYNOPSYS_UNCONNECTED__1297, 
        SYNOPSYS_UNCONNECTED__1298, SYNOPSYS_UNCONNECTED__1299, 
        SYNOPSYS_UNCONNECTED__1300, SYNOPSYS_UNCONNECTED__1301, 
        SYNOPSYS_UNCONNECTED__1302, SYNOPSYS_UNCONNECTED__1303, 
        SYNOPSYS_UNCONNECTED__1304, SYNOPSYS_UNCONNECTED__1305, 
        SYNOPSYS_UNCONNECTED__1306, SYNOPSYS_UNCONNECTED__1307, 
        SYNOPSYS_UNCONNECTED__1308, SYNOPSYS_UNCONNECTED__1309, 
        SYNOPSYS_UNCONNECTED__1310, SYNOPSYS_UNCONNECTED__1311, 
        SYNOPSYS_UNCONNECTED__1312, SYNOPSYS_UNCONNECTED__1313, 
        SYNOPSYS_UNCONNECTED__1314, SYNOPSYS_UNCONNECTED__1315, 
        SYNOPSYS_UNCONNECTED__1316, SYNOPSYS_UNCONNECTED__1317, 
        SYNOPSYS_UNCONNECTED__1318, SYNOPSYS_UNCONNECTED__1319, 
        SYNOPSYS_UNCONNECTED__1320, SYNOPSYS_UNCONNECTED__1321, 
        SYNOPSYS_UNCONNECTED__1322, SYNOPSYS_UNCONNECTED__1323, 
        SYNOPSYS_UNCONNECTED__1324, SYNOPSYS_UNCONNECTED__1325, 
        SYNOPSYS_UNCONNECTED__1326, SYNOPSYS_UNCONNECTED__1327, 
        SYNOPSYS_UNCONNECTED__1328, SYNOPSYS_UNCONNECTED__1329, 
        SYNOPSYS_UNCONNECTED__1330, SYNOPSYS_UNCONNECTED__1331, 
        SYNOPSYS_UNCONNECTED__1332, SYNOPSYS_UNCONNECTED__1333, 
        SYNOPSYS_UNCONNECTED__1334, SYNOPSYS_UNCONNECTED__1335, 
        SYNOPSYS_UNCONNECTED__1336, SYNOPSYS_UNCONNECTED__1337, 
        SYNOPSYS_UNCONNECTED__1338, SYNOPSYS_UNCONNECTED__1339, 
        SYNOPSYS_UNCONNECTED__1340, SYNOPSYS_UNCONNECTED__1341, 
        SYNOPSYS_UNCONNECTED__1342, SYNOPSYS_UNCONNECTED__1343, 
        SYNOPSYS_UNCONNECTED__1344, SYNOPSYS_UNCONNECTED__1345, 
        SYNOPSYS_UNCONNECTED__1346, SYNOPSYS_UNCONNECTED__1347, 
        SYNOPSYS_UNCONNECTED__1348, SYNOPSYS_UNCONNECTED__1349, 
        SYNOPSYS_UNCONNECTED__1350, SYNOPSYS_UNCONNECTED__1351, 
        SYNOPSYS_UNCONNECTED__1352, SYNOPSYS_UNCONNECTED__1353, 
        SYNOPSYS_UNCONNECTED__1354, SYNOPSYS_UNCONNECTED__1355, 
        SYNOPSYS_UNCONNECTED__1356, SYNOPSYS_UNCONNECTED__1357, 
        SYNOPSYS_UNCONNECTED__1358, SYNOPSYS_UNCONNECTED__1359, 
        SYNOPSYS_UNCONNECTED__1360, SYNOPSYS_UNCONNECTED__1361, 
        SYNOPSYS_UNCONNECTED__1362, SYNOPSYS_UNCONNECTED__1363, 
        SYNOPSYS_UNCONNECTED__1364, SYNOPSYS_UNCONNECTED__1365, 
        SYNOPSYS_UNCONNECTED__1366, SYNOPSYS_UNCONNECTED__1367, 
        SYNOPSYS_UNCONNECTED__1368, SYNOPSYS_UNCONNECTED__1369, 
        SYNOPSYS_UNCONNECTED__1370, SYNOPSYS_UNCONNECTED__1371, 
        SYNOPSYS_UNCONNECTED__1372, SYNOPSYS_UNCONNECTED__1373, 
        SYNOPSYS_UNCONNECTED__1374, SYNOPSYS_UNCONNECTED__1375, 
        SYNOPSYS_UNCONNECTED__1376, SYNOPSYS_UNCONNECTED__1377, 
        SYNOPSYS_UNCONNECTED__1378, SYNOPSYS_UNCONNECTED__1379, 
        SYNOPSYS_UNCONNECTED__1380, SYNOPSYS_UNCONNECTED__1381, 
        SYNOPSYS_UNCONNECTED__1382, SYNOPSYS_UNCONNECTED__1383, 
        SYNOPSYS_UNCONNECTED__1384, SYNOPSYS_UNCONNECTED__1385, 
        SYNOPSYS_UNCONNECTED__1386, SYNOPSYS_UNCONNECTED__1387, 
        SYNOPSYS_UNCONNECTED__1388, SYNOPSYS_UNCONNECTED__1389, 
        SYNOPSYS_UNCONNECTED__1390, SYNOPSYS_UNCONNECTED__1391, 
        SYNOPSYS_UNCONNECTED__1392, SYNOPSYS_UNCONNECTED__1393, 
        SYNOPSYS_UNCONNECTED__1394, SYNOPSYS_UNCONNECTED__1395, 
        SYNOPSYS_UNCONNECTED__1396, SYNOPSYS_UNCONNECTED__1397, 
        SYNOPSYS_UNCONNECTED__1398, SYNOPSYS_UNCONNECTED__1399, 
        SYNOPSYS_UNCONNECTED__1400, SYNOPSYS_UNCONNECTED__1401, 
        SYNOPSYS_UNCONNECTED__1402, SYNOPSYS_UNCONNECTED__1403, 
        SYNOPSYS_UNCONNECTED__1404, SYNOPSYS_UNCONNECTED__1405, 
        SYNOPSYS_UNCONNECTED__1406, SYNOPSYS_UNCONNECTED__1407, 
        SYNOPSYS_UNCONNECTED__1408, SYNOPSYS_UNCONNECTED__1409, 
        SYNOPSYS_UNCONNECTED__1410, SYNOPSYS_UNCONNECTED__1411, 
        SYNOPSYS_UNCONNECTED__1412, SYNOPSYS_UNCONNECTED__1413, 
        SYNOPSYS_UNCONNECTED__1414, SYNOPSYS_UNCONNECTED__1415, 
        SYNOPSYS_UNCONNECTED__1416, SYNOPSYS_UNCONNECTED__1417, 
        SYNOPSYS_UNCONNECTED__1418, SYNOPSYS_UNCONNECTED__1419, 
        SYNOPSYS_UNCONNECTED__1420, SYNOPSYS_UNCONNECTED__1421, 
        SYNOPSYS_UNCONNECTED__1422, SYNOPSYS_UNCONNECTED__1423, 
        SYNOPSYS_UNCONNECTED__1424, SYNOPSYS_UNCONNECTED__1425, 
        SYNOPSYS_UNCONNECTED__1426, SYNOPSYS_UNCONNECTED__1427, 
        SYNOPSYS_UNCONNECTED__1428, SYNOPSYS_UNCONNECTED__1429, 
        SYNOPSYS_UNCONNECTED__1430, SYNOPSYS_UNCONNECTED__1431, 
        SYNOPSYS_UNCONNECTED__1432, SYNOPSYS_UNCONNECTED__1433, 
        SYNOPSYS_UNCONNECTED__1434, SYNOPSYS_UNCONNECTED__1435, 
        SYNOPSYS_UNCONNECTED__1436, SYNOPSYS_UNCONNECTED__1437, 
        SYNOPSYS_UNCONNECTED__1438, SYNOPSYS_UNCONNECTED__1439, 
        SYNOPSYS_UNCONNECTED__1440, SYNOPSYS_UNCONNECTED__1441, 
        SYNOPSYS_UNCONNECTED__1442, SYNOPSYS_UNCONNECTED__1443, 
        SYNOPSYS_UNCONNECTED__1444, SYNOPSYS_UNCONNECTED__1445, 
        SYNOPSYS_UNCONNECTED__1446, SYNOPSYS_UNCONNECTED__1447, 
        SYNOPSYS_UNCONNECTED__1448, SYNOPSYS_UNCONNECTED__1449, 
        SYNOPSYS_UNCONNECTED__1450, SYNOPSYS_UNCONNECTED__1451, 
        SYNOPSYS_UNCONNECTED__1452, SYNOPSYS_UNCONNECTED__1453, 
        SYNOPSYS_UNCONNECTED__1454, SYNOPSYS_UNCONNECTED__1455, 
        SYNOPSYS_UNCONNECTED__1456, SYNOPSYS_UNCONNECTED__1457, 
        SYNOPSYS_UNCONNECTED__1458, SYNOPSYS_UNCONNECTED__1459, 
        SYNOPSYS_UNCONNECTED__1460, SYNOPSYS_UNCONNECTED__1461, 
        SYNOPSYS_UNCONNECTED__1462, SYNOPSYS_UNCONNECTED__1463, 
        SYNOPSYS_UNCONNECTED__1464, SYNOPSYS_UNCONNECTED__1465, 
        SYNOPSYS_UNCONNECTED__1466, SYNOPSYS_UNCONNECTED__1467, 
        SYNOPSYS_UNCONNECTED__1468, SYNOPSYS_UNCONNECTED__1469, 
        SYNOPSYS_UNCONNECTED__1470, SYNOPSYS_UNCONNECTED__1471, 
        SYNOPSYS_UNCONNECTED__1472, SYNOPSYS_UNCONNECTED__1473, 
        SYNOPSYS_UNCONNECTED__1474, SYNOPSYS_UNCONNECTED__1475, 
        SYNOPSYS_UNCONNECTED__1476, SYNOPSYS_UNCONNECTED__1477, 
        SYNOPSYS_UNCONNECTED__1478, SYNOPSYS_UNCONNECTED__1479, 
        SYNOPSYS_UNCONNECTED__1480, SYNOPSYS_UNCONNECTED__1481, 
        SYNOPSYS_UNCONNECTED__1482, SYNOPSYS_UNCONNECTED__1483, 
        SYNOPSYS_UNCONNECTED__1484, SYNOPSYS_UNCONNECTED__1485, 
        SYNOPSYS_UNCONNECTED__1486, SYNOPSYS_UNCONNECTED__1487, 
        SYNOPSYS_UNCONNECTED__1488, SYNOPSYS_UNCONNECTED__1489, 
        SYNOPSYS_UNCONNECTED__1490, SYNOPSYS_UNCONNECTED__1491, 
        SYNOPSYS_UNCONNECTED__1492, SYNOPSYS_UNCONNECTED__1493, 
        SYNOPSYS_UNCONNECTED__1494, SYNOPSYS_UNCONNECTED__1495, 
        SYNOPSYS_UNCONNECTED__1496, SYNOPSYS_UNCONNECTED__1497, 
        SYNOPSYS_UNCONNECTED__1498, SYNOPSYS_UNCONNECTED__1499, 
        SYNOPSYS_UNCONNECTED__1500, SYNOPSYS_UNCONNECTED__1501, 
        SYNOPSYS_UNCONNECTED__1502, SYNOPSYS_UNCONNECTED__1503, 
        SYNOPSYS_UNCONNECTED__1504, SYNOPSYS_UNCONNECTED__1505, 
        SYNOPSYS_UNCONNECTED__1506, SYNOPSYS_UNCONNECTED__1507, 
        SYNOPSYS_UNCONNECTED__1508, SYNOPSYS_UNCONNECTED__1509, 
        SYNOPSYS_UNCONNECTED__1510, SYNOPSYS_UNCONNECTED__1511, 
        SYNOPSYS_UNCONNECTED__1512, SYNOPSYS_UNCONNECTED__1513, 
        SYNOPSYS_UNCONNECTED__1514, SYNOPSYS_UNCONNECTED__1515, 
        SYNOPSYS_UNCONNECTED__1516, SYNOPSYS_UNCONNECTED__1517, 
        SYNOPSYS_UNCONNECTED__1518, SYNOPSYS_UNCONNECTED__1519, 
        SYNOPSYS_UNCONNECTED__1520, SYNOPSYS_UNCONNECTED__1521, 
        SYNOPSYS_UNCONNECTED__1522, SYNOPSYS_UNCONNECTED__1523, 
        SYNOPSYS_UNCONNECTED__1524, SYNOPSYS_UNCONNECTED__1525, 
        SYNOPSYS_UNCONNECTED__1526, SYNOPSYS_UNCONNECTED__1527, 
        SYNOPSYS_UNCONNECTED__1528, SYNOPSYS_UNCONNECTED__1529, 
        SYNOPSYS_UNCONNECTED__1530, SYNOPSYS_UNCONNECTED__1531, 
        SYNOPSYS_UNCONNECTED__1532, SYNOPSYS_UNCONNECTED__1533, 
        SYNOPSYS_UNCONNECTED__1534, SYNOPSYS_UNCONNECTED__1535, 
        SYNOPSYS_UNCONNECTED__1536, SYNOPSYS_UNCONNECTED__1537, 
        SYNOPSYS_UNCONNECTED__1538, SYNOPSYS_UNCONNECTED__1539, 
        SYNOPSYS_UNCONNECTED__1540, SYNOPSYS_UNCONNECTED__1541, 
        SYNOPSYS_UNCONNECTED__1542, SYNOPSYS_UNCONNECTED__1543, 
        SYNOPSYS_UNCONNECTED__1544, SYNOPSYS_UNCONNECTED__1545, 
        SYNOPSYS_UNCONNECTED__1546, SYNOPSYS_UNCONNECTED__1547, 
        SYNOPSYS_UNCONNECTED__1548, SYNOPSYS_UNCONNECTED__1549, 
        SYNOPSYS_UNCONNECTED__1550, SYNOPSYS_UNCONNECTED__1551, 
        SYNOPSYS_UNCONNECTED__1552, SYNOPSYS_UNCONNECTED__1553, 
        SYNOPSYS_UNCONNECTED__1554, SYNOPSYS_UNCONNECTED__1555, 
        SYNOPSYS_UNCONNECTED__1556, SYNOPSYS_UNCONNECTED__1557, 
        SYNOPSYS_UNCONNECTED__1558, SYNOPSYS_UNCONNECTED__1559, 
        SYNOPSYS_UNCONNECTED__1560, SYNOPSYS_UNCONNECTED__1561, 
        SYNOPSYS_UNCONNECTED__1562, SYNOPSYS_UNCONNECTED__1563, 
        SYNOPSYS_UNCONNECTED__1564, SYNOPSYS_UNCONNECTED__1565, 
        SYNOPSYS_UNCONNECTED__1566, SYNOPSYS_UNCONNECTED__1567, 
        SYNOPSYS_UNCONNECTED__1568, SYNOPSYS_UNCONNECTED__1569, 
        SYNOPSYS_UNCONNECTED__1570, SYNOPSYS_UNCONNECTED__1571, 
        SYNOPSYS_UNCONNECTED__1572, SYNOPSYS_UNCONNECTED__1573, 
        SYNOPSYS_UNCONNECTED__1574, SYNOPSYS_UNCONNECTED__1575, 
        SYNOPSYS_UNCONNECTED__1576, SYNOPSYS_UNCONNECTED__1577, 
        SYNOPSYS_UNCONNECTED__1578, SYNOPSYS_UNCONNECTED__1579, 
        SYNOPSYS_UNCONNECTED__1580, SYNOPSYS_UNCONNECTED__1581, 
        SYNOPSYS_UNCONNECTED__1582, SYNOPSYS_UNCONNECTED__1583, 
        SYNOPSYS_UNCONNECTED__1584, SYNOPSYS_UNCONNECTED__1585, 
        SYNOPSYS_UNCONNECTED__1586, SYNOPSYS_UNCONNECTED__1587, 
        SYNOPSYS_UNCONNECTED__1588, SYNOPSYS_UNCONNECTED__1589, 
        SYNOPSYS_UNCONNECTED__1590, SYNOPSYS_UNCONNECTED__1591, 
        SYNOPSYS_UNCONNECTED__1592, SYNOPSYS_UNCONNECTED__1593, 
        SYNOPSYS_UNCONNECTED__1594, SYNOPSYS_UNCONNECTED__1595, 
        SYNOPSYS_UNCONNECTED__1596, SYNOPSYS_UNCONNECTED__1597, 
        SYNOPSYS_UNCONNECTED__1598, SYNOPSYS_UNCONNECTED__1599, 
        SYNOPSYS_UNCONNECTED__1600, SYNOPSYS_UNCONNECTED__1601, 
        SYNOPSYS_UNCONNECTED__1602, SYNOPSYS_UNCONNECTED__1603, 
        SYNOPSYS_UNCONNECTED__1604, SYNOPSYS_UNCONNECTED__1605, 
        SYNOPSYS_UNCONNECTED__1606, SYNOPSYS_UNCONNECTED__1607, 
        SYNOPSYS_UNCONNECTED__1608, SYNOPSYS_UNCONNECTED__1609, 
        SYNOPSYS_UNCONNECTED__1610, SYNOPSYS_UNCONNECTED__1611, 
        SYNOPSYS_UNCONNECTED__1612, SYNOPSYS_UNCONNECTED__1613, 
        SYNOPSYS_UNCONNECTED__1614, SYNOPSYS_UNCONNECTED__1615, 
        SYNOPSYS_UNCONNECTED__1616, SYNOPSYS_UNCONNECTED__1617, 
        SYNOPSYS_UNCONNECTED__1618, SYNOPSYS_UNCONNECTED__1619, 
        SYNOPSYS_UNCONNECTED__1620, SYNOPSYS_UNCONNECTED__1621, 
        SYNOPSYS_UNCONNECTED__1622, SYNOPSYS_UNCONNECTED__1623, 
        SYNOPSYS_UNCONNECTED__1624, SYNOPSYS_UNCONNECTED__1625, 
        SYNOPSYS_UNCONNECTED__1626, SYNOPSYS_UNCONNECTED__1627, 
        SYNOPSYS_UNCONNECTED__1628, SYNOPSYS_UNCONNECTED__1629, 
        SYNOPSYS_UNCONNECTED__1630, SYNOPSYS_UNCONNECTED__1631, 
        SYNOPSYS_UNCONNECTED__1632, SYNOPSYS_UNCONNECTED__1633, 
        SYNOPSYS_UNCONNECTED__1634, SYNOPSYS_UNCONNECTED__1635, 
        SYNOPSYS_UNCONNECTED__1636, SYNOPSYS_UNCONNECTED__1637, 
        SYNOPSYS_UNCONNECTED__1638, SYNOPSYS_UNCONNECTED__1639, 
        SYNOPSYS_UNCONNECTED__1640, SYNOPSYS_UNCONNECTED__1641, 
        SYNOPSYS_UNCONNECTED__1642, SYNOPSYS_UNCONNECTED__1643, 
        SYNOPSYS_UNCONNECTED__1644, SYNOPSYS_UNCONNECTED__1645, 
        SYNOPSYS_UNCONNECTED__1646, SYNOPSYS_UNCONNECTED__1647, 
        SYNOPSYS_UNCONNECTED__1648, SYNOPSYS_UNCONNECTED__1649, 
        SYNOPSYS_UNCONNECTED__1650, SYNOPSYS_UNCONNECTED__1651, 
        SYNOPSYS_UNCONNECTED__1652, SYNOPSYS_UNCONNECTED__1653, 
        SYNOPSYS_UNCONNECTED__1654, SYNOPSYS_UNCONNECTED__1655, 
        SYNOPSYS_UNCONNECTED__1656, SYNOPSYS_UNCONNECTED__1657, 
        SYNOPSYS_UNCONNECTED__1658, SYNOPSYS_UNCONNECTED__1659, 
        SYNOPSYS_UNCONNECTED__1660, SYNOPSYS_UNCONNECTED__1661, 
        SYNOPSYS_UNCONNECTED__1662, SYNOPSYS_UNCONNECTED__1663, 
        SYNOPSYS_UNCONNECTED__1664, SYNOPSYS_UNCONNECTED__1665, 
        SYNOPSYS_UNCONNECTED__1666, SYNOPSYS_UNCONNECTED__1667, 
        SYNOPSYS_UNCONNECTED__1668, SYNOPSYS_UNCONNECTED__1669, 
        SYNOPSYS_UNCONNECTED__1670, SYNOPSYS_UNCONNECTED__1671, 
        SYNOPSYS_UNCONNECTED__1672, SYNOPSYS_UNCONNECTED__1673, 
        SYNOPSYS_UNCONNECTED__1674, SYNOPSYS_UNCONNECTED__1675, 
        SYNOPSYS_UNCONNECTED__1676, SYNOPSYS_UNCONNECTED__1677, 
        SYNOPSYS_UNCONNECTED__1678, SYNOPSYS_UNCONNECTED__1679, 
        SYNOPSYS_UNCONNECTED__1680, SYNOPSYS_UNCONNECTED__1681, 
        SYNOPSYS_UNCONNECTED__1682, SYNOPSYS_UNCONNECTED__1683, 
        SYNOPSYS_UNCONNECTED__1684, SYNOPSYS_UNCONNECTED__1685, 
        SYNOPSYS_UNCONNECTED__1686, SYNOPSYS_UNCONNECTED__1687, 
        SYNOPSYS_UNCONNECTED__1688, SYNOPSYS_UNCONNECTED__1689, 
        SYNOPSYS_UNCONNECTED__1690, SYNOPSYS_UNCONNECTED__1691, 
        SYNOPSYS_UNCONNECTED__1692, SYNOPSYS_UNCONNECTED__1693, 
        SYNOPSYS_UNCONNECTED__1694, SYNOPSYS_UNCONNECTED__1695, 
        SYNOPSYS_UNCONNECTED__1696, SYNOPSYS_UNCONNECTED__1697, 
        SYNOPSYS_UNCONNECTED__1698, SYNOPSYS_UNCONNECTED__1699, 
        SYNOPSYS_UNCONNECTED__1700, SYNOPSYS_UNCONNECTED__1701, 
        SYNOPSYS_UNCONNECTED__1702, SYNOPSYS_UNCONNECTED__1703, 
        SYNOPSYS_UNCONNECTED__1704, SYNOPSYS_UNCONNECTED__1705, 
        SYNOPSYS_UNCONNECTED__1706, SYNOPSYS_UNCONNECTED__1707, 
        SYNOPSYS_UNCONNECTED__1708, SYNOPSYS_UNCONNECTED__1709, 
        SYNOPSYS_UNCONNECTED__1710, SYNOPSYS_UNCONNECTED__1711, 
        SYNOPSYS_UNCONNECTED__1712, SYNOPSYS_UNCONNECTED__1713, 
        SYNOPSYS_UNCONNECTED__1714, SYNOPSYS_UNCONNECTED__1715, 
        SYNOPSYS_UNCONNECTED__1716, SYNOPSYS_UNCONNECTED__1717, 
        SYNOPSYS_UNCONNECTED__1718, SYNOPSYS_UNCONNECTED__1719, 
        SYNOPSYS_UNCONNECTED__1720, SYNOPSYS_UNCONNECTED__1721, 
        SYNOPSYS_UNCONNECTED__1722, SYNOPSYS_UNCONNECTED__1723, 
        SYNOPSYS_UNCONNECTED__1724, SYNOPSYS_UNCONNECTED__1725, 
        SYNOPSYS_UNCONNECTED__1726, SYNOPSYS_UNCONNECTED__1727, 
        SYNOPSYS_UNCONNECTED__1728, SYNOPSYS_UNCONNECTED__1729, 
        SYNOPSYS_UNCONNECTED__1730, SYNOPSYS_UNCONNECTED__1731, 
        SYNOPSYS_UNCONNECTED__1732, SYNOPSYS_UNCONNECTED__1733, 
        SYNOPSYS_UNCONNECTED__1734, SYNOPSYS_UNCONNECTED__1735, 
        SYNOPSYS_UNCONNECTED__1736, SYNOPSYS_UNCONNECTED__1737, 
        SYNOPSYS_UNCONNECTED__1738, SYNOPSYS_UNCONNECTED__1739, 
        SYNOPSYS_UNCONNECTED__1740, SYNOPSYS_UNCONNECTED__1741, 
        SYNOPSYS_UNCONNECTED__1742, SYNOPSYS_UNCONNECTED__1743, 
        SYNOPSYS_UNCONNECTED__1744, SYNOPSYS_UNCONNECTED__1745, 
        SYNOPSYS_UNCONNECTED__1746, SYNOPSYS_UNCONNECTED__1747, 
        SYNOPSYS_UNCONNECTED__1748, SYNOPSYS_UNCONNECTED__1749, 
        SYNOPSYS_UNCONNECTED__1750, SYNOPSYS_UNCONNECTED__1751, 
        SYNOPSYS_UNCONNECTED__1752, SYNOPSYS_UNCONNECTED__1753, 
        SYNOPSYS_UNCONNECTED__1754, SYNOPSYS_UNCONNECTED__1755, 
        SYNOPSYS_UNCONNECTED__1756, SYNOPSYS_UNCONNECTED__1757, 
        SYNOPSYS_UNCONNECTED__1758, SYNOPSYS_UNCONNECTED__1759, 
        SYNOPSYS_UNCONNECTED__1760, SYNOPSYS_UNCONNECTED__1761, 
        SYNOPSYS_UNCONNECTED__1762, SYNOPSYS_UNCONNECTED__1763, 
        SYNOPSYS_UNCONNECTED__1764, SYNOPSYS_UNCONNECTED__1765, 
        SYNOPSYS_UNCONNECTED__1766, SYNOPSYS_UNCONNECTED__1767, 
        SYNOPSYS_UNCONNECTED__1768, SYNOPSYS_UNCONNECTED__1769, 
        SYNOPSYS_UNCONNECTED__1770, SYNOPSYS_UNCONNECTED__1771, 
        SYNOPSYS_UNCONNECTED__1772, SYNOPSYS_UNCONNECTED__1773, 
        SYNOPSYS_UNCONNECTED__1774, SYNOPSYS_UNCONNECTED__1775, 
        SYNOPSYS_UNCONNECTED__1776, SYNOPSYS_UNCONNECTED__1777, 
        SYNOPSYS_UNCONNECTED__1778, SYNOPSYS_UNCONNECTED__1779, 
        SYNOPSYS_UNCONNECTED__1780, SYNOPSYS_UNCONNECTED__1781, 
        SYNOPSYS_UNCONNECTED__1782, SYNOPSYS_UNCONNECTED__1783, 
        SYNOPSYS_UNCONNECTED__1784, SYNOPSYS_UNCONNECTED__1785, 
        SYNOPSYS_UNCONNECTED__1786, SYNOPSYS_UNCONNECTED__1787, 
        SYNOPSYS_UNCONNECTED__1788, SYNOPSYS_UNCONNECTED__1789, 
        SYNOPSYS_UNCONNECTED__1790, SYNOPSYS_UNCONNECTED__1791, 
        SYNOPSYS_UNCONNECTED__1792, SYNOPSYS_UNCONNECTED__1793, 
        SYNOPSYS_UNCONNECTED__1794, SYNOPSYS_UNCONNECTED__1795, 
        SYNOPSYS_UNCONNECTED__1796, SYNOPSYS_UNCONNECTED__1797, 
        SYNOPSYS_UNCONNECTED__1798, SYNOPSYS_UNCONNECTED__1799, 
        SYNOPSYS_UNCONNECTED__1800, SYNOPSYS_UNCONNECTED__1801, 
        SYNOPSYS_UNCONNECTED__1802, SYNOPSYS_UNCONNECTED__1803, 
        SYNOPSYS_UNCONNECTED__1804, SYNOPSYS_UNCONNECTED__1805, 
        SYNOPSYS_UNCONNECTED__1806, SYNOPSYS_UNCONNECTED__1807, 
        SYNOPSYS_UNCONNECTED__1808, SYNOPSYS_UNCONNECTED__1809, 
        SYNOPSYS_UNCONNECTED__1810, SYNOPSYS_UNCONNECTED__1811, 
        SYNOPSYS_UNCONNECTED__1812, SYNOPSYS_UNCONNECTED__1813, 
        SYNOPSYS_UNCONNECTED__1814, SYNOPSYS_UNCONNECTED__1815, 
        SYNOPSYS_UNCONNECTED__1816, SYNOPSYS_UNCONNECTED__1817, 
        SYNOPSYS_UNCONNECTED__1818, SYNOPSYS_UNCONNECTED__1819, 
        SYNOPSYS_UNCONNECTED__1820, SYNOPSYS_UNCONNECTED__1821, 
        SYNOPSYS_UNCONNECTED__1822, SYNOPSYS_UNCONNECTED__1823, 
        SYNOPSYS_UNCONNECTED__1824, SYNOPSYS_UNCONNECTED__1825, 
        SYNOPSYS_UNCONNECTED__1826, SYNOPSYS_UNCONNECTED__1827, 
        SYNOPSYS_UNCONNECTED__1828, SYNOPSYS_UNCONNECTED__1829, 
        SYNOPSYS_UNCONNECTED__1830, SYNOPSYS_UNCONNECTED__1831, 
        SYNOPSYS_UNCONNECTED__1832, SYNOPSYS_UNCONNECTED__1833, 
        SYNOPSYS_UNCONNECTED__1834, SYNOPSYS_UNCONNECTED__1835, 
        SYNOPSYS_UNCONNECTED__1836, SYNOPSYS_UNCONNECTED__1837, 
        SYNOPSYS_UNCONNECTED__1838, SYNOPSYS_UNCONNECTED__1839, 
        SYNOPSYS_UNCONNECTED__1840, SYNOPSYS_UNCONNECTED__1841, 
        SYNOPSYS_UNCONNECTED__1842, SYNOPSYS_UNCONNECTED__1843, 
        SYNOPSYS_UNCONNECTED__1844, SYNOPSYS_UNCONNECTED__1845, 
        SYNOPSYS_UNCONNECTED__1846, SYNOPSYS_UNCONNECTED__1847, 
        SYNOPSYS_UNCONNECTED__1848, SYNOPSYS_UNCONNECTED__1849, 
        SYNOPSYS_UNCONNECTED__1850, SYNOPSYS_UNCONNECTED__1851, 
        SYNOPSYS_UNCONNECTED__1852, SYNOPSYS_UNCONNECTED__1853, 
        SYNOPSYS_UNCONNECTED__1854, SYNOPSYS_UNCONNECTED__1855, 
        SYNOPSYS_UNCONNECTED__1856, SYNOPSYS_UNCONNECTED__1857, 
        SYNOPSYS_UNCONNECTED__1858, SYNOPSYS_UNCONNECTED__1859, 
        SYNOPSYS_UNCONNECTED__1860, SYNOPSYS_UNCONNECTED__1861, 
        SYNOPSYS_UNCONNECTED__1862, SYNOPSYS_UNCONNECTED__1863, 
        SYNOPSYS_UNCONNECTED__1864, SYNOPSYS_UNCONNECTED__1865, 
        SYNOPSYS_UNCONNECTED__1866, SYNOPSYS_UNCONNECTED__1867, 
        SYNOPSYS_UNCONNECTED__1868, SYNOPSYS_UNCONNECTED__1869, 
        SYNOPSYS_UNCONNECTED__1870, SYNOPSYS_UNCONNECTED__1871, 
        SYNOPSYS_UNCONNECTED__1872, SYNOPSYS_UNCONNECTED__1873, 
        SYNOPSYS_UNCONNECTED__1874, SYNOPSYS_UNCONNECTED__1875, 
        SYNOPSYS_UNCONNECTED__1876, SYNOPSYS_UNCONNECTED__1877, 
        SYNOPSYS_UNCONNECTED__1878, SYNOPSYS_UNCONNECTED__1879, 
        SYNOPSYS_UNCONNECTED__1880, SYNOPSYS_UNCONNECTED__1881, 
        SYNOPSYS_UNCONNECTED__1882, SYNOPSYS_UNCONNECTED__1883, 
        SYNOPSYS_UNCONNECTED__1884, SYNOPSYS_UNCONNECTED__1885, 
        SYNOPSYS_UNCONNECTED__1886, SYNOPSYS_UNCONNECTED__1887, 
        SYNOPSYS_UNCONNECTED__1888, SYNOPSYS_UNCONNECTED__1889, 
        SYNOPSYS_UNCONNECTED__1890, SYNOPSYS_UNCONNECTED__1891, 
        SYNOPSYS_UNCONNECTED__1892, SYNOPSYS_UNCONNECTED__1893, 
        SYNOPSYS_UNCONNECTED__1894, SYNOPSYS_UNCONNECTED__1895, 
        SYNOPSYS_UNCONNECTED__1896, SYNOPSYS_UNCONNECTED__1897, 
        SYNOPSYS_UNCONNECTED__1898, SYNOPSYS_UNCONNECTED__1899, 
        SYNOPSYS_UNCONNECTED__1900, SYNOPSYS_UNCONNECTED__1901, 
        SYNOPSYS_UNCONNECTED__1902, SYNOPSYS_UNCONNECTED__1903, 
        SYNOPSYS_UNCONNECTED__1904, SYNOPSYS_UNCONNECTED__1905, 
        SYNOPSYS_UNCONNECTED__1906, SYNOPSYS_UNCONNECTED__1907, 
        SYNOPSYS_UNCONNECTED__1908, SYNOPSYS_UNCONNECTED__1909, 
        SYNOPSYS_UNCONNECTED__1910, SYNOPSYS_UNCONNECTED__1911, 
        SYNOPSYS_UNCONNECTED__1912, SYNOPSYS_UNCONNECTED__1913, 
        SYNOPSYS_UNCONNECTED__1914, SYNOPSYS_UNCONNECTED__1915, 
        SYNOPSYS_UNCONNECTED__1916, SYNOPSYS_UNCONNECTED__1917, 
        SYNOPSYS_UNCONNECTED__1918, SYNOPSYS_UNCONNECTED__1919, 
        SYNOPSYS_UNCONNECTED__1920, SYNOPSYS_UNCONNECTED__1921, 
        SYNOPSYS_UNCONNECTED__1922, SYNOPSYS_UNCONNECTED__1923, 
        SYNOPSYS_UNCONNECTED__1924, SYNOPSYS_UNCONNECTED__1925, 
        SYNOPSYS_UNCONNECTED__1926, SYNOPSYS_UNCONNECTED__1927, 
        SYNOPSYS_UNCONNECTED__1928, SYNOPSYS_UNCONNECTED__1929, 
        SYNOPSYS_UNCONNECTED__1930, SYNOPSYS_UNCONNECTED__1931, 
        SYNOPSYS_UNCONNECTED__1932, SYNOPSYS_UNCONNECTED__1933, 
        SYNOPSYS_UNCONNECTED__1934, SYNOPSYS_UNCONNECTED__1935, 
        SYNOPSYS_UNCONNECTED__1936, SYNOPSYS_UNCONNECTED__1937, 
        SYNOPSYS_UNCONNECTED__1938, SYNOPSYS_UNCONNECTED__1939, 
        SYNOPSYS_UNCONNECTED__1940, SYNOPSYS_UNCONNECTED__1941, 
        SYNOPSYS_UNCONNECTED__1942, SYNOPSYS_UNCONNECTED__1943, 
        SYNOPSYS_UNCONNECTED__1944, SYNOPSYS_UNCONNECTED__1945, 
        SYNOPSYS_UNCONNECTED__1946, SYNOPSYS_UNCONNECTED__1947, 
        SYNOPSYS_UNCONNECTED__1948, SYNOPSYS_UNCONNECTED__1949, 
        SYNOPSYS_UNCONNECTED__1950, SYNOPSYS_UNCONNECTED__1951, 
        SYNOPSYS_UNCONNECTED__1952, SYNOPSYS_UNCONNECTED__1953, 
        SYNOPSYS_UNCONNECTED__1954, SYNOPSYS_UNCONNECTED__1955, 
        SYNOPSYS_UNCONNECTED__1956, SYNOPSYS_UNCONNECTED__1957, 
        SYNOPSYS_UNCONNECTED__1958, SYNOPSYS_UNCONNECTED__1959, 
        SYNOPSYS_UNCONNECTED__1960, SYNOPSYS_UNCONNECTED__1961, 
        SYNOPSYS_UNCONNECTED__1962, SYNOPSYS_UNCONNECTED__1963, 
        SYNOPSYS_UNCONNECTED__1964, SYNOPSYS_UNCONNECTED__1965, 
        SYNOPSYS_UNCONNECTED__1966, SYNOPSYS_UNCONNECTED__1967, 
        SYNOPSYS_UNCONNECTED__1968, SYNOPSYS_UNCONNECTED__1969, 
        SYNOPSYS_UNCONNECTED__1970, SYNOPSYS_UNCONNECTED__1971, 
        SYNOPSYS_UNCONNECTED__1972, SYNOPSYS_UNCONNECTED__1973, 
        SYNOPSYS_UNCONNECTED__1974, SYNOPSYS_UNCONNECTED__1975, 
        SYNOPSYS_UNCONNECTED__1976, SYNOPSYS_UNCONNECTED__1977, 
        SYNOPSYS_UNCONNECTED__1978, SYNOPSYS_UNCONNECTED__1979, 
        SYNOPSYS_UNCONNECTED__1980, SYNOPSYS_UNCONNECTED__1981, 
        SYNOPSYS_UNCONNECTED__1982, SYNOPSYS_UNCONNECTED__1983, 
        SYNOPSYS_UNCONNECTED__1984, SYNOPSYS_UNCONNECTED__1985, 
        SYNOPSYS_UNCONNECTED__1986, SYNOPSYS_UNCONNECTED__1987, 
        SYNOPSYS_UNCONNECTED__1988, SYNOPSYS_UNCONNECTED__1989, 
        SYNOPSYS_UNCONNECTED__1990, SYNOPSYS_UNCONNECTED__1991, 
        SYNOPSYS_UNCONNECTED__1992, SYNOPSYS_UNCONNECTED__1993, 
        SYNOPSYS_UNCONNECTED__1994, SYNOPSYS_UNCONNECTED__1995, 
        SYNOPSYS_UNCONNECTED__1996, SYNOPSYS_UNCONNECTED__1997, 
        SYNOPSYS_UNCONNECTED__1998, SYNOPSYS_UNCONNECTED__1999, 
        SYNOPSYS_UNCONNECTED__2000, SYNOPSYS_UNCONNECTED__2001, 
        SYNOPSYS_UNCONNECTED__2002, SYNOPSYS_UNCONNECTED__2003;

  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .Q(oglobal[11]) );
  DFF \oglobal_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .Q(oglobal[12]) );
  DFF \oglobal_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .Q(oglobal[13]) );
  hamming_N16000_CC2_DW01_add_0 add_97 ( .A(oglobal), .B({1'b0, olocal}), .CI(
        1'b0), .SUM(o) );
  hamming_N16000_CC2_DW01_add_1 add_2667_root_add_71_I832 ( .A({1'b0, N69222, 
        N69221, N69220, N69219, N69218, N69217, N69216, N69215, N69214, N69213, 
        N69212, N69211}), .B({N69236, N69235, N69234, N69233, N69232, N69231, 
        N69230, N69229, N69228, N69227, N69226, N69225, N69224}), .CI(1'b0), 
        .SUM(olocal) );
  hamming_N16000_CC2_DW01_add_2 add_2668_root_add_71_I832 ( .A({1'b0, N69196, 
        N69195, N69194, N69193, N69192, N69191, N69190, N69189, N69188, N69187, 
        N69186, N69185}), .B({1'b0, N69209, N69208, N69207, N69206, N69205, 
        N69204, N69203, N69202, N69201, N69200, N69199, N69198}), .CI(1'b0), 
        .SUM({N69236, N69235, N69234, N69233, N69232, N69231, N69230, N69229, 
        N69228, N69227, N69226, N69225, N69224}) );
  hamming_N16000_CC2_DW01_add_3 add_2669_root_add_71_I832 ( .A({1'b0, 1'b0, 
        N69169, N69168, N69167, N69166, N69165, N69164, N69163, N69162, N69161, 
        N69160, N69159}), .B({1'b0, 1'b0, N69182, N69181, N69180, N69179, 
        N69178, N69177, N69176, N69175, N69174, N69173, N69172}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__0, N69222, N69221, N69220, N69219, N69218, 
        N69217, N69216, N69215, N69214, N69213, N69212, N69211}) );
  hamming_N16000_CC2_DW01_add_4 add_2670_root_add_71_I832 ( .A({1'b0, 1'b0, 
        N69143, N69142, N69141, N69140, N69139, N69138, N69137, N69136, N69135, 
        N69134, N69133}), .B({1'b0, 1'b0, N69156, N69155, N69154, N69153, 
        N69152, N69151, N69150, N69149, N69148, N69147, N69146}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__1, N69209, N69208, N69207, N69206, N69205, 
        N69204, N69203, N69202, N69201, N69200, N69199, N69198}) );
  hamming_N16000_CC2_DW01_add_5 add_2671_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, N69116, N69115, N69114, N69113, N69112, N69111, N69110, N69109, 
        N69108, N69107}), .B({1'b0, 1'b0, N69130, N69129, N69128, N69127, 
        N69126, N69125, N69124, N69123, N69122, N69121, N69120}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__2, N69196, N69195, N69194, N69193, N69192, 
        N69191, N69190, N69189, N69188, N69187, N69186, N69185}) );
  hamming_N16000_CC2_DW01_add_6 add_2672_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, N69090, N69089, N69088, N69087, N69086, N69085, N69084, N69083, 
        N69082, N69081}), .B({1'b0, 1'b0, 1'b0, N69103, N69102, N69101, N69100, 
        N69099, N69098, N69097, N69096, N69095, N69094}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, N69182, N69181, 
        N69180, N69179, N69178, N69177, N69176, N69175, N69174, N69173, N69172}) );
  hamming_N16000_CC2_DW01_add_7 add_2673_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, N69064, N69063, N69062, N69061, N69060, N69059, N69058, N69057, 
        N69056, N69055}), .B({1'b0, 1'b0, 1'b0, N69077, N69076, N69075, N69074, 
        N69073, N69072, N69071, N69070, N69069, N69068}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, N69169, N69168, 
        N69167, N69166, N69165, N69164, N69163, N69162, N69161, N69160, N69159}) );
  hamming_N16000_CC2_DW01_add_8 add_2674_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, N69038, N69037, N69036, N69035, N69034, N69033, N69032, N69031, 
        N69030, N69029}), .B({1'b0, 1'b0, 1'b0, N69051, N69050, N69049, N69048, 
        N69047, N69046, N69045, N69044, N69043, N69042}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, N69156, N69155, 
        N69154, N69153, N69152, N69151, N69150, N69149, N69148, N69147, N69146}) );
  hamming_N16000_CC2_DW01_add_9 add_2675_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, N69012, N69011, N69010, N69009, N69008, N69007, N69006, N69005, 
        N69004, N69003}), .B({1'b0, 1'b0, 1'b0, N69025, N69024, N69023, N69022, 
        N69021, N69020, N69019, N69018, N69017, N69016}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, N69143, N69142, 
        N69141, N69140, N69139, N69138, N69137, N69136, N69135, N69134, N69133}) );
  hamming_N16000_CC2_DW01_add_10 add_2676_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N68985, N68984, N68983, N68982, N68981, N68980, N68979, 
        N68978, N68977}), .B({1'b0, 1'b0, 1'b0, N68999, N68998, N68997, N68996, 
        N68995, N68994, N68993, N68992, N68991, N68990}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, N69130, N69129, 
        N69128, N69127, N69126, N69125, N69124, N69123, N69122, N69121, N69120}) );
  hamming_N16000_CC2_DW01_add_11 add_2677_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N68959, N68958, N68957, N68956, N68955, N68954, N68953, 
        N68952, N68951}), .B({1'b0, 1'b0, 1'b0, 1'b0, N68972, N68971, N68970, 
        N68969, N68968, N68967, N68966, N68965, N68964}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N69116, N69115, N69114, N69113, N69112, 
        N69111, N69110, N69109, N69108, N69107}) );
  hamming_N16000_CC2_DW01_add_12 add_2678_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N68933, N68932, N68931, N68930, N68929, N68928, N68927, 
        N68926, N68925}), .B({1'b0, 1'b0, 1'b0, 1'b0, N68946, N68945, N68944, 
        N68943, N68942, N68941, N68940, N68939, N68938}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, N69103, N69102, N69101, N69100, N69099, 
        N69098, N69097, N69096, N69095, N69094}) );
  hamming_N16000_CC2_DW01_add_13 add_2679_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N68907, N68906, N68905, N68904, N68903, N68902, N68901, 
        N68900, N68899}), .B({1'b0, 1'b0, 1'b0, 1'b0, N68920, N68919, N68918, 
        N68917, N68916, N68915, N68914, N68913, N68912}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, N69090, N69089, N69088, N69087, N69086, 
        N69085, N69084, N69083, N69082, N69081}) );
  hamming_N16000_CC2_DW01_add_14 add_2680_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N68881, N68880, N68879, N68878, N68877, N68876, N68875, 
        N68874, N68873}), .B({1'b0, 1'b0, 1'b0, 1'b0, N68894, N68893, N68892, 
        N68891, N68890, N68889, N68888, N68887, N68886}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, N69077, N69076, N69075, N69074, N69073, 
        N69072, N69071, N69070, N69069, N69068}) );
  hamming_N16000_CC2_DW01_add_15 add_2681_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N68855, N68854, N68853, N68852, N68851, N68850, N68849, 
        N68848, N68847}), .B({1'b0, 1'b0, 1'b0, 1'b0, N68868, N68867, N68866, 
        N68865, N68864, N68863, N68862, N68861, N68860}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, N69064, N69063, N69062, N69061, N69060, 
        N69059, N69058, N69057, N69056, N69055}) );
  hamming_N16000_CC2_DW01_add_16 add_2682_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N68829, N68828, N68827, N68826, N68825, N68824, N68823, 
        N68822, N68821}), .B({1'b0, 1'b0, 1'b0, 1'b0, N68842, N68841, N68840, 
        N68839, N68838, N68837, N68836, N68835, N68834}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, N69051, N69050, N69049, N69048, N69047, 
        N69046, N69045, N69044, N69043, N69042}) );
  hamming_N16000_CC2_DW01_add_17 add_2683_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N68803, N68802, N68801, N68800, N68799, N68798, N68797, 
        N68796, N68795}), .B({1'b0, 1'b0, 1'b0, 1'b0, N68816, N68815, N68814, 
        N68813, N68812, N68811, N68810, N68809, N68808}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, N69038, N69037, N69036, N69035, N69034, 
        N69033, N69032, N69031, N69030, N69029}) );
  hamming_N16000_CC2_DW01_add_18 add_2684_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N68777, N68776, N68775, N68774, N68773, N68772, N68771, 
        N68770, N68769}), .B({1'b0, 1'b0, 1'b0, 1'b0, N68790, N68789, N68788, 
        N68787, N68786, N68785, N68784, N68783, N68782}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, N69025, N69024, N69023, N69022, N69021, 
        N69020, N69019, N69018, N69017, N69016}) );
  hamming_N16000_CC2_DW01_add_19 add_2685_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N68751, N68750, N68749, N68748, N68747, N68746, N68745, 
        N68744, N68743}), .B({1'b0, 1'b0, 1'b0, 1'b0, N68764, N68763, N68762, 
        N68761, N68760, N68759, N68758, N68757, N68756}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, N69012, N69011, N69010, N69009, N69008, 
        N69007, N69006, N69005, N69004, N69003}) );
  hamming_N16000_CC2_DW01_add_20 add_2686_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N68725, N68724, N68723, N68722, N68721, N68720, N68719, 
        N68718, N68717}), .B({1'b0, 1'b0, 1'b0, 1'b0, N68738, N68737, N68736, 
        N68735, N68734, N68733, N68732, N68731, N68730}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, N68999, N68998, N68997, N68996, N68995, 
        N68994, N68993, N68992, N68991, N68990}) );
  hamming_N16000_CC2_DW01_add_21 add_2687_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68698, N68697, N68696, N68695, N68694, N68693, 
        N68692, N68691}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68711, N68710, 
        N68709, N68708, N68707, N68706, N68705, N68704}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, N68985, N68984, 
        N68983, N68982, N68981, N68980, N68979, N68978, N68977}) );
  hamming_N16000_CC2_DW01_add_22 add_2688_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68672, N68671, N68670, N68669, N68668, N68667, 
        N68666, N68665}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68685, N68684, 
        N68683, N68682, N68681, N68680, N68679, N68678}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, N68972, N68971, 
        N68970, N68969, N68968, N68967, N68966, N68965, N68964}) );
  hamming_N16000_CC2_DW01_add_23 add_2689_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68646, N68645, N68644, N68643, N68642, N68641, 
        N68640, N68639}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68659, N68658, 
        N68657, N68656, N68655, N68654, N68653, N68652}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, N68959, N68958, 
        N68957, N68956, N68955, N68954, N68953, N68952, N68951}) );
  hamming_N16000_CC2_DW01_add_24 add_2690_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68620, N68619, N68618, N68617, N68616, N68615, 
        N68614, N68613}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68633, N68632, 
        N68631, N68630, N68629, N68628, N68627, N68626}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58, N68946, N68945, 
        N68944, N68943, N68942, N68941, N68940, N68939, N68938}) );
  hamming_N16000_CC2_DW01_add_25 add_2691_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68594, N68593, N68592, N68591, N68590, N68589, 
        N68588, N68587}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68607, N68606, 
        N68605, N68604, N68603, N68602, N68601, N68600}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, 
        SYNOPSYS_UNCONNECTED__61, SYNOPSYS_UNCONNECTED__62, N68933, N68932, 
        N68931, N68930, N68929, N68928, N68927, N68926, N68925}) );
  hamming_N16000_CC2_DW01_add_26 add_2692_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68568, N68567, N68566, N68565, N68564, N68563, 
        N68562, N68561}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68581, N68580, 
        N68579, N68578, N68577, N68576, N68575, N68574}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__63, SYNOPSYS_UNCONNECTED__64, 
        SYNOPSYS_UNCONNECTED__65, SYNOPSYS_UNCONNECTED__66, N68920, N68919, 
        N68918, N68917, N68916, N68915, N68914, N68913, N68912}) );
  hamming_N16000_CC2_DW01_add_27 add_2693_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68542, N68541, N68540, N68539, N68538, N68537, 
        N68536, N68535}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68555, N68554, 
        N68553, N68552, N68551, N68550, N68549, N68548}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__67, SYNOPSYS_UNCONNECTED__68, 
        SYNOPSYS_UNCONNECTED__69, SYNOPSYS_UNCONNECTED__70, N68907, N68906, 
        N68905, N68904, N68903, N68902, N68901, N68900, N68899}) );
  hamming_N16000_CC2_DW01_add_28 add_2694_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68516, N68515, N68514, N68513, N68512, N68511, 
        N68510, N68509}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68529, N68528, 
        N68527, N68526, N68525, N68524, N68523, N68522}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__71, SYNOPSYS_UNCONNECTED__72, 
        SYNOPSYS_UNCONNECTED__73, SYNOPSYS_UNCONNECTED__74, N68894, N68893, 
        N68892, N68891, N68890, N68889, N68888, N68887, N68886}) );
  hamming_N16000_CC2_DW01_add_29 add_2695_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68490, N68489, N68488, N68487, N68486, N68485, 
        N68484, N68483}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68503, N68502, 
        N68501, N68500, N68499, N68498, N68497, N68496}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__75, SYNOPSYS_UNCONNECTED__76, 
        SYNOPSYS_UNCONNECTED__77, SYNOPSYS_UNCONNECTED__78, N68881, N68880, 
        N68879, N68878, N68877, N68876, N68875, N68874, N68873}) );
  hamming_N16000_CC2_DW01_add_30 add_2696_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68464, N68463, N68462, N68461, N68460, N68459, 
        N68458, N68457}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68477, N68476, 
        N68475, N68474, N68473, N68472, N68471, N68470}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__79, SYNOPSYS_UNCONNECTED__80, 
        SYNOPSYS_UNCONNECTED__81, SYNOPSYS_UNCONNECTED__82, N68868, N68867, 
        N68866, N68865, N68864, N68863, N68862, N68861, N68860}) );
  hamming_N16000_CC2_DW01_add_31 add_2697_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68438, N68437, N68436, N68435, N68434, N68433, 
        N68432, N68431}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68451, N68450, 
        N68449, N68448, N68447, N68446, N68445, N68444}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__83, SYNOPSYS_UNCONNECTED__84, 
        SYNOPSYS_UNCONNECTED__85, SYNOPSYS_UNCONNECTED__86, N68855, N68854, 
        N68853, N68852, N68851, N68850, N68849, N68848, N68847}) );
  hamming_N16000_CC2_DW01_add_32 add_2698_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68412, N68411, N68410, N68409, N68408, N68407, 
        N68406, N68405}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68425, N68424, 
        N68423, N68422, N68421, N68420, N68419, N68418}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__87, SYNOPSYS_UNCONNECTED__88, 
        SYNOPSYS_UNCONNECTED__89, SYNOPSYS_UNCONNECTED__90, N68842, N68841, 
        N68840, N68839, N68838, N68837, N68836, N68835, N68834}) );
  hamming_N16000_CC2_DW01_add_33 add_2699_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68386, N68385, N68384, N68383, N68382, N68381, 
        N68380, N68379}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68399, N68398, 
        N68397, N68396, N68395, N68394, N68393, N68392}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__91, SYNOPSYS_UNCONNECTED__92, 
        SYNOPSYS_UNCONNECTED__93, SYNOPSYS_UNCONNECTED__94, N68829, N68828, 
        N68827, N68826, N68825, N68824, N68823, N68822, N68821}) );
  hamming_N16000_CC2_DW01_add_34 add_2700_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68360, N68359, N68358, N68357, N68356, N68355, 
        N68354, N68353}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68373, N68372, 
        N68371, N68370, N68369, N68368, N68367, N68366}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__95, SYNOPSYS_UNCONNECTED__96, 
        SYNOPSYS_UNCONNECTED__97, SYNOPSYS_UNCONNECTED__98, N68816, N68815, 
        N68814, N68813, N68812, N68811, N68810, N68809, N68808}) );
  hamming_N16000_CC2_DW01_add_35 add_2701_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68334, N68333, N68332, N68331, N68330, N68329, 
        N68328, N68327}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68347, N68346, 
        N68345, N68344, N68343, N68342, N68341, N68340}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__99, SYNOPSYS_UNCONNECTED__100, 
        SYNOPSYS_UNCONNECTED__101, SYNOPSYS_UNCONNECTED__102, N68803, N68802, 
        N68801, N68800, N68799, N68798, N68797, N68796, N68795}) );
  hamming_N16000_CC2_DW01_add_36 add_2702_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68308, N68307, N68306, N68305, N68304, N68303, 
        N68302, N68301}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68321, N68320, 
        N68319, N68318, N68317, N68316, N68315, N68314}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__103, SYNOPSYS_UNCONNECTED__104, 
        SYNOPSYS_UNCONNECTED__105, SYNOPSYS_UNCONNECTED__106, N68790, N68789, 
        N68788, N68787, N68786, N68785, N68784, N68783, N68782}) );
  hamming_N16000_CC2_DW01_add_37 add_2703_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68282, N68281, N68280, N68279, N68278, N68277, 
        N68276, N68275}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68295, N68294, 
        N68293, N68292, N68291, N68290, N68289, N68288}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__107, SYNOPSYS_UNCONNECTED__108, 
        SYNOPSYS_UNCONNECTED__109, SYNOPSYS_UNCONNECTED__110, N68777, N68776, 
        N68775, N68774, N68773, N68772, N68771, N68770, N68769}) );
  hamming_N16000_CC2_DW01_add_38 add_2704_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68256, N68255, N68254, N68253, N68252, N68251, 
        N68250, N68249}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68269, N68268, 
        N68267, N68266, N68265, N68264, N68263, N68262}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__111, SYNOPSYS_UNCONNECTED__112, 
        SYNOPSYS_UNCONNECTED__113, SYNOPSYS_UNCONNECTED__114, N68764, N68763, 
        N68762, N68761, N68760, N68759, N68758, N68757, N68756}) );
  hamming_N16000_CC2_DW01_add_39 add_2705_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68230, N68229, N68228, N68227, N68226, N68225, 
        N68224, N68223}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68243, N68242, 
        N68241, N68240, N68239, N68238, N68237, N68236}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__115, SYNOPSYS_UNCONNECTED__116, 
        SYNOPSYS_UNCONNECTED__117, SYNOPSYS_UNCONNECTED__118, N68751, N68750, 
        N68749, N68748, N68747, N68746, N68745, N68744, N68743}) );
  hamming_N16000_CC2_DW01_add_40 add_2706_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68204, N68203, N68202, N68201, N68200, N68199, 
        N68198, N68197}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68217, N68216, 
        N68215, N68214, N68213, N68212, N68211, N68210}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__119, SYNOPSYS_UNCONNECTED__120, 
        SYNOPSYS_UNCONNECTED__121, SYNOPSYS_UNCONNECTED__122, N68738, N68737, 
        N68736, N68735, N68734, N68733, N68732, N68731, N68730}) );
  hamming_N16000_CC2_DW01_add_41 add_2707_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N68178, N68177, N68176, N68175, N68174, N68173, 
        N68172, N68171}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68191, N68190, 
        N68189, N68188, N68187, N68186, N68185, N68184}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__123, SYNOPSYS_UNCONNECTED__124, 
        SYNOPSYS_UNCONNECTED__125, SYNOPSYS_UNCONNECTED__126, N68725, N68724, 
        N68723, N68722, N68721, N68720, N68719, N68718, N68717}) );
  hamming_N16000_CC2_DW01_add_42 add_2708_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N68151, N68150, N68149, N68148, N68147, N68146, 
        N68145}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68164, N68163, 
        N68162, N68161, N68160, N68159, N68158}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__127, SYNOPSYS_UNCONNECTED__128, 
        SYNOPSYS_UNCONNECTED__129, SYNOPSYS_UNCONNECTED__130, 
        SYNOPSYS_UNCONNECTED__131, N68711, N68710, N68709, N68708, N68707, 
        N68706, N68705, N68704}) );
  hamming_N16000_CC2_DW01_add_43 add_2709_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N68125, N68124, N68123, N68122, N68121, N68120, 
        N68119}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68138, N68137, 
        N68136, N68135, N68134, N68133, N68132}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__132, SYNOPSYS_UNCONNECTED__133, 
        SYNOPSYS_UNCONNECTED__134, SYNOPSYS_UNCONNECTED__135, 
        SYNOPSYS_UNCONNECTED__136, N68698, N68697, N68696, N68695, N68694, 
        N68693, N68692, N68691}) );
  hamming_N16000_CC2_DW01_add_44 add_2710_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N68099, N68098, N68097, N68096, N68095, N68094, 
        N68093}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68112, N68111, 
        N68110, N68109, N68108, N68107, N68106}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__137, SYNOPSYS_UNCONNECTED__138, 
        SYNOPSYS_UNCONNECTED__139, SYNOPSYS_UNCONNECTED__140, 
        SYNOPSYS_UNCONNECTED__141, N68685, N68684, N68683, N68682, N68681, 
        N68680, N68679, N68678}) );
  hamming_N16000_CC2_DW01_add_45 add_2711_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N68073, N68072, N68071, N68070, N68069, N68068, 
        N68067}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68086, N68085, 
        N68084, N68083, N68082, N68081, N68080}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__142, SYNOPSYS_UNCONNECTED__143, 
        SYNOPSYS_UNCONNECTED__144, SYNOPSYS_UNCONNECTED__145, 
        SYNOPSYS_UNCONNECTED__146, N68672, N68671, N68670, N68669, N68668, 
        N68667, N68666, N68665}) );
  hamming_N16000_CC2_DW01_add_46 add_2712_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N68047, N68046, N68045, N68044, N68043, N68042, 
        N68041}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68060, N68059, 
        N68058, N68057, N68056, N68055, N68054}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__147, SYNOPSYS_UNCONNECTED__148, 
        SYNOPSYS_UNCONNECTED__149, SYNOPSYS_UNCONNECTED__150, 
        SYNOPSYS_UNCONNECTED__151, N68659, N68658, N68657, N68656, N68655, 
        N68654, N68653, N68652}) );
  hamming_N16000_CC2_DW01_add_47 add_2713_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N68021, N68020, N68019, N68018, N68017, N68016, 
        N68015}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68034, N68033, 
        N68032, N68031, N68030, N68029, N68028}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__152, SYNOPSYS_UNCONNECTED__153, 
        SYNOPSYS_UNCONNECTED__154, SYNOPSYS_UNCONNECTED__155, 
        SYNOPSYS_UNCONNECTED__156, N68646, N68645, N68644, N68643, N68642, 
        N68641, N68640, N68639}) );
  hamming_N16000_CC2_DW01_add_48 add_2714_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67995, N67994, N67993, N67992, N67991, N67990, 
        N67989}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N68008, N68007, 
        N68006, N68005, N68004, N68003, N68002}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__157, SYNOPSYS_UNCONNECTED__158, 
        SYNOPSYS_UNCONNECTED__159, SYNOPSYS_UNCONNECTED__160, 
        SYNOPSYS_UNCONNECTED__161, N68633, N68632, N68631, N68630, N68629, 
        N68628, N68627, N68626}) );
  hamming_N16000_CC2_DW01_add_49 add_2715_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67969, N67968, N67967, N67966, N67965, N67964, 
        N67963}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67982, N67981, 
        N67980, N67979, N67978, N67977, N67976}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__162, SYNOPSYS_UNCONNECTED__163, 
        SYNOPSYS_UNCONNECTED__164, SYNOPSYS_UNCONNECTED__165, 
        SYNOPSYS_UNCONNECTED__166, N68620, N68619, N68618, N68617, N68616, 
        N68615, N68614, N68613}) );
  hamming_N16000_CC2_DW01_add_50 add_2716_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67943, N67942, N67941, N67940, N67939, N67938, 
        N67937}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67956, N67955, 
        N67954, N67953, N67952, N67951, N67950}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__167, SYNOPSYS_UNCONNECTED__168, 
        SYNOPSYS_UNCONNECTED__169, SYNOPSYS_UNCONNECTED__170, 
        SYNOPSYS_UNCONNECTED__171, N68607, N68606, N68605, N68604, N68603, 
        N68602, N68601, N68600}) );
  hamming_N16000_CC2_DW01_add_51 add_2717_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67917, N67916, N67915, N67914, N67913, N67912, 
        N67911}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67930, N67929, 
        N67928, N67927, N67926, N67925, N67924}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__172, SYNOPSYS_UNCONNECTED__173, 
        SYNOPSYS_UNCONNECTED__174, SYNOPSYS_UNCONNECTED__175, 
        SYNOPSYS_UNCONNECTED__176, N68594, N68593, N68592, N68591, N68590, 
        N68589, N68588, N68587}) );
  hamming_N16000_CC2_DW01_add_52 add_2718_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67891, N67890, N67889, N67888, N67887, N67886, 
        N67885}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67904, N67903, 
        N67902, N67901, N67900, N67899, N67898}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__177, SYNOPSYS_UNCONNECTED__178, 
        SYNOPSYS_UNCONNECTED__179, SYNOPSYS_UNCONNECTED__180, 
        SYNOPSYS_UNCONNECTED__181, N68581, N68580, N68579, N68578, N68577, 
        N68576, N68575, N68574}) );
  hamming_N16000_CC2_DW01_add_53 add_2719_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67865, N67864, N67863, N67862, N67861, N67860, 
        N67859}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67878, N67877, 
        N67876, N67875, N67874, N67873, N67872}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__182, SYNOPSYS_UNCONNECTED__183, 
        SYNOPSYS_UNCONNECTED__184, SYNOPSYS_UNCONNECTED__185, 
        SYNOPSYS_UNCONNECTED__186, N68568, N68567, N68566, N68565, N68564, 
        N68563, N68562, N68561}) );
  hamming_N16000_CC2_DW01_add_54 add_2720_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67839, N67838, N67837, N67836, N67835, N67834, 
        N67833}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67852, N67851, 
        N67850, N67849, N67848, N67847, N67846}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__187, SYNOPSYS_UNCONNECTED__188, 
        SYNOPSYS_UNCONNECTED__189, SYNOPSYS_UNCONNECTED__190, 
        SYNOPSYS_UNCONNECTED__191, N68555, N68554, N68553, N68552, N68551, 
        N68550, N68549, N68548}) );
  hamming_N16000_CC2_DW01_add_55 add_2721_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67813, N67812, N67811, N67810, N67809, N67808, 
        N67807}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67826, N67825, 
        N67824, N67823, N67822, N67821, N67820}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__192, SYNOPSYS_UNCONNECTED__193, 
        SYNOPSYS_UNCONNECTED__194, SYNOPSYS_UNCONNECTED__195, 
        SYNOPSYS_UNCONNECTED__196, N68542, N68541, N68540, N68539, N68538, 
        N68537, N68536, N68535}) );
  hamming_N16000_CC2_DW01_add_56 add_2722_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67787, N67786, N67785, N67784, N67783, N67782, 
        N67781}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67800, N67799, 
        N67798, N67797, N67796, N67795, N67794}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__197, SYNOPSYS_UNCONNECTED__198, 
        SYNOPSYS_UNCONNECTED__199, SYNOPSYS_UNCONNECTED__200, 
        SYNOPSYS_UNCONNECTED__201, N68529, N68528, N68527, N68526, N68525, 
        N68524, N68523, N68522}) );
  hamming_N16000_CC2_DW01_add_57 add_2723_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67761, N67760, N67759, N67758, N67757, N67756, 
        N67755}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67774, N67773, 
        N67772, N67771, N67770, N67769, N67768}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__202, SYNOPSYS_UNCONNECTED__203, 
        SYNOPSYS_UNCONNECTED__204, SYNOPSYS_UNCONNECTED__205, 
        SYNOPSYS_UNCONNECTED__206, N68516, N68515, N68514, N68513, N68512, 
        N68511, N68510, N68509}) );
  hamming_N16000_CC2_DW01_add_58 add_2724_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67735, N67734, N67733, N67732, N67731, N67730, 
        N67729}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67748, N67747, 
        N67746, N67745, N67744, N67743, N67742}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__207, SYNOPSYS_UNCONNECTED__208, 
        SYNOPSYS_UNCONNECTED__209, SYNOPSYS_UNCONNECTED__210, 
        SYNOPSYS_UNCONNECTED__211, N68503, N68502, N68501, N68500, N68499, 
        N68498, N68497, N68496}) );
  hamming_N16000_CC2_DW01_add_59 add_2725_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67709, N67708, N67707, N67706, N67705, N67704, 
        N67703}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67722, N67721, 
        N67720, N67719, N67718, N67717, N67716}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__212, SYNOPSYS_UNCONNECTED__213, 
        SYNOPSYS_UNCONNECTED__214, SYNOPSYS_UNCONNECTED__215, 
        SYNOPSYS_UNCONNECTED__216, N68490, N68489, N68488, N68487, N68486, 
        N68485, N68484, N68483}) );
  hamming_N16000_CC2_DW01_add_60 add_2726_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67683, N67682, N67681, N67680, N67679, N67678, 
        N67677}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67696, N67695, 
        N67694, N67693, N67692, N67691, N67690}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__217, SYNOPSYS_UNCONNECTED__218, 
        SYNOPSYS_UNCONNECTED__219, SYNOPSYS_UNCONNECTED__220, 
        SYNOPSYS_UNCONNECTED__221, N68477, N68476, N68475, N68474, N68473, 
        N68472, N68471, N68470}) );
  hamming_N16000_CC2_DW01_add_61 add_2727_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67657, N67656, N67655, N67654, N67653, N67652, 
        N67651}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67670, N67669, 
        N67668, N67667, N67666, N67665, N67664}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__222, SYNOPSYS_UNCONNECTED__223, 
        SYNOPSYS_UNCONNECTED__224, SYNOPSYS_UNCONNECTED__225, 
        SYNOPSYS_UNCONNECTED__226, N68464, N68463, N68462, N68461, N68460, 
        N68459, N68458, N68457}) );
  hamming_N16000_CC2_DW01_add_62 add_2728_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67631, N67630, N67629, N67628, N67627, N67626, 
        N67625}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67644, N67643, 
        N67642, N67641, N67640, N67639, N67638}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__227, SYNOPSYS_UNCONNECTED__228, 
        SYNOPSYS_UNCONNECTED__229, SYNOPSYS_UNCONNECTED__230, 
        SYNOPSYS_UNCONNECTED__231, N68451, N68450, N68449, N68448, N68447, 
        N68446, N68445, N68444}) );
  hamming_N16000_CC2_DW01_add_63 add_2729_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67605, N67604, N67603, N67602, N67601, N67600, 
        N67599}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67618, N67617, 
        N67616, N67615, N67614, N67613, N67612}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__232, SYNOPSYS_UNCONNECTED__233, 
        SYNOPSYS_UNCONNECTED__234, SYNOPSYS_UNCONNECTED__235, 
        SYNOPSYS_UNCONNECTED__236, N68438, N68437, N68436, N68435, N68434, 
        N68433, N68432, N68431}) );
  hamming_N16000_CC2_DW01_add_64 add_2730_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67579, N67578, N67577, N67576, N67575, N67574, 
        N67573}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67592, N67591, 
        N67590, N67589, N67588, N67587, N67586}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__237, SYNOPSYS_UNCONNECTED__238, 
        SYNOPSYS_UNCONNECTED__239, SYNOPSYS_UNCONNECTED__240, 
        SYNOPSYS_UNCONNECTED__241, N68425, N68424, N68423, N68422, N68421, 
        N68420, N68419, N68418}) );
  hamming_N16000_CC2_DW01_add_65 add_2731_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67553, N67552, N67551, N67550, N67549, N67548, 
        N67547}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67566, N67565, 
        N67564, N67563, N67562, N67561, N67560}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__242, SYNOPSYS_UNCONNECTED__243, 
        SYNOPSYS_UNCONNECTED__244, SYNOPSYS_UNCONNECTED__245, 
        SYNOPSYS_UNCONNECTED__246, N68412, N68411, N68410, N68409, N68408, 
        N68407, N68406, N68405}) );
  hamming_N16000_CC2_DW01_add_66 add_2732_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67527, N67526, N67525, N67524, N67523, N67522, 
        N67521}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67540, N67539, 
        N67538, N67537, N67536, N67535, N67534}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__247, SYNOPSYS_UNCONNECTED__248, 
        SYNOPSYS_UNCONNECTED__249, SYNOPSYS_UNCONNECTED__250, 
        SYNOPSYS_UNCONNECTED__251, N68399, N68398, N68397, N68396, N68395, 
        N68394, N68393, N68392}) );
  hamming_N16000_CC2_DW01_add_67 add_2733_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67501, N67500, N67499, N67498, N67497, N67496, 
        N67495}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67514, N67513, 
        N67512, N67511, N67510, N67509, N67508}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__252, SYNOPSYS_UNCONNECTED__253, 
        SYNOPSYS_UNCONNECTED__254, SYNOPSYS_UNCONNECTED__255, 
        SYNOPSYS_UNCONNECTED__256, N68386, N68385, N68384, N68383, N68382, 
        N68381, N68380, N68379}) );
  hamming_N16000_CC2_DW01_add_68 add_2734_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67475, N67474, N67473, N67472, N67471, N67470, 
        N67469}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67488, N67487, 
        N67486, N67485, N67484, N67483, N67482}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__257, SYNOPSYS_UNCONNECTED__258, 
        SYNOPSYS_UNCONNECTED__259, SYNOPSYS_UNCONNECTED__260, 
        SYNOPSYS_UNCONNECTED__261, N68373, N68372, N68371, N68370, N68369, 
        N68368, N68367, N68366}) );
  hamming_N16000_CC2_DW01_add_69 add_2735_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67449, N67448, N67447, N67446, N67445, N67444, 
        N67443}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67462, N67461, 
        N67460, N67459, N67458, N67457, N67456}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__262, SYNOPSYS_UNCONNECTED__263, 
        SYNOPSYS_UNCONNECTED__264, SYNOPSYS_UNCONNECTED__265, 
        SYNOPSYS_UNCONNECTED__266, N68360, N68359, N68358, N68357, N68356, 
        N68355, N68354, N68353}) );
  hamming_N16000_CC2_DW01_add_70 add_2736_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67423, N67422, N67421, N67420, N67419, N67418, 
        N67417}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67436, N67435, 
        N67434, N67433, N67432, N67431, N67430}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__267, SYNOPSYS_UNCONNECTED__268, 
        SYNOPSYS_UNCONNECTED__269, SYNOPSYS_UNCONNECTED__270, 
        SYNOPSYS_UNCONNECTED__271, N68347, N68346, N68345, N68344, N68343, 
        N68342, N68341, N68340}) );
  hamming_N16000_CC2_DW01_add_71 add_2737_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67397, N67396, N67395, N67394, N67393, N67392, 
        N67391}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67410, N67409, 
        N67408, N67407, N67406, N67405, N67404}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__272, SYNOPSYS_UNCONNECTED__273, 
        SYNOPSYS_UNCONNECTED__274, SYNOPSYS_UNCONNECTED__275, 
        SYNOPSYS_UNCONNECTED__276, N68334, N68333, N68332, N68331, N68330, 
        N68329, N68328, N68327}) );
  hamming_N16000_CC2_DW01_add_72 add_2738_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67371, N67370, N67369, N67368, N67367, N67366, 
        N67365}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67384, N67383, 
        N67382, N67381, N67380, N67379, N67378}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__277, SYNOPSYS_UNCONNECTED__278, 
        SYNOPSYS_UNCONNECTED__279, SYNOPSYS_UNCONNECTED__280, 
        SYNOPSYS_UNCONNECTED__281, N68321, N68320, N68319, N68318, N68317, 
        N68316, N68315, N68314}) );
  hamming_N16000_CC2_DW01_add_73 add_2739_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67345, N67344, N67343, N67342, N67341, N67340, 
        N67339}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67358, N67357, 
        N67356, N67355, N67354, N67353, N67352}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__282, SYNOPSYS_UNCONNECTED__283, 
        SYNOPSYS_UNCONNECTED__284, SYNOPSYS_UNCONNECTED__285, 
        SYNOPSYS_UNCONNECTED__286, N68308, N68307, N68306, N68305, N68304, 
        N68303, N68302, N68301}) );
  hamming_N16000_CC2_DW01_add_74 add_2740_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67319, N67318, N67317, N67316, N67315, N67314, 
        N67313}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67332, N67331, 
        N67330, N67329, N67328, N67327, N67326}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__287, SYNOPSYS_UNCONNECTED__288, 
        SYNOPSYS_UNCONNECTED__289, SYNOPSYS_UNCONNECTED__290, 
        SYNOPSYS_UNCONNECTED__291, N68295, N68294, N68293, N68292, N68291, 
        N68290, N68289, N68288}) );
  hamming_N16000_CC2_DW01_add_75 add_2741_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67293, N67292, N67291, N67290, N67289, N67288, 
        N67287}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67306, N67305, 
        N67304, N67303, N67302, N67301, N67300}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__292, SYNOPSYS_UNCONNECTED__293, 
        SYNOPSYS_UNCONNECTED__294, SYNOPSYS_UNCONNECTED__295, 
        SYNOPSYS_UNCONNECTED__296, N68282, N68281, N68280, N68279, N68278, 
        N68277, N68276, N68275}) );
  hamming_N16000_CC2_DW01_add_76 add_2742_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67267, N67266, N67265, N67264, N67263, N67262, 
        N67261}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67280, N67279, 
        N67278, N67277, N67276, N67275, N67274}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__297, SYNOPSYS_UNCONNECTED__298, 
        SYNOPSYS_UNCONNECTED__299, SYNOPSYS_UNCONNECTED__300, 
        SYNOPSYS_UNCONNECTED__301, N68269, N68268, N68267, N68266, N68265, 
        N68264, N68263, N68262}) );
  hamming_N16000_CC2_DW01_add_77 add_2743_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67241, N67240, N67239, N67238, N67237, N67236, 
        N67235}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67254, N67253, 
        N67252, N67251, N67250, N67249, N67248}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__302, SYNOPSYS_UNCONNECTED__303, 
        SYNOPSYS_UNCONNECTED__304, SYNOPSYS_UNCONNECTED__305, 
        SYNOPSYS_UNCONNECTED__306, N68256, N68255, N68254, N68253, N68252, 
        N68251, N68250, N68249}) );
  hamming_N16000_CC2_DW01_add_78 add_2744_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67215, N67214, N67213, N67212, N67211, N67210, 
        N67209}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67228, N67227, 
        N67226, N67225, N67224, N67223, N67222}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__307, SYNOPSYS_UNCONNECTED__308, 
        SYNOPSYS_UNCONNECTED__309, SYNOPSYS_UNCONNECTED__310, 
        SYNOPSYS_UNCONNECTED__311, N68243, N68242, N68241, N68240, N68239, 
        N68238, N68237, N68236}) );
  hamming_N16000_CC2_DW01_add_79 add_2745_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67189, N67188, N67187, N67186, N67185, N67184, 
        N67183}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67202, N67201, 
        N67200, N67199, N67198, N67197, N67196}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__312, SYNOPSYS_UNCONNECTED__313, 
        SYNOPSYS_UNCONNECTED__314, SYNOPSYS_UNCONNECTED__315, 
        SYNOPSYS_UNCONNECTED__316, N68230, N68229, N68228, N68227, N68226, 
        N68225, N68224, N68223}) );
  hamming_N16000_CC2_DW01_add_80 add_2746_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67163, N67162, N67161, N67160, N67159, N67158, 
        N67157}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67176, N67175, 
        N67174, N67173, N67172, N67171, N67170}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__317, SYNOPSYS_UNCONNECTED__318, 
        SYNOPSYS_UNCONNECTED__319, SYNOPSYS_UNCONNECTED__320, 
        SYNOPSYS_UNCONNECTED__321, N68217, N68216, N68215, N68214, N68213, 
        N68212, N68211, N68210}) );
  hamming_N16000_CC2_DW01_add_81 add_2747_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67137, N67136, N67135, N67134, N67133, N67132, 
        N67131}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67150, N67149, 
        N67148, N67147, N67146, N67145, N67144}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__322, SYNOPSYS_UNCONNECTED__323, 
        SYNOPSYS_UNCONNECTED__324, SYNOPSYS_UNCONNECTED__325, 
        SYNOPSYS_UNCONNECTED__326, N68204, N68203, N68202, N68201, N68200, 
        N68199, N68198, N68197}) );
  hamming_N16000_CC2_DW01_add_82 add_2748_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, N67111, N67110, N67109, N67108, N67107, N67106, 
        N67105}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67124, N67123, 
        N67122, N67121, N67120, N67119, N67118}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__327, SYNOPSYS_UNCONNECTED__328, 
        SYNOPSYS_UNCONNECTED__329, SYNOPSYS_UNCONNECTED__330, 
        SYNOPSYS_UNCONNECTED__331, N68191, N68190, N68189, N68188, N68187, 
        N68186, N68185, N68184}) );
  hamming_N16000_CC2_DW01_add_83 add_2749_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67084, N67083, N67082, N67081, N67080, 
        N67079}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67098, N67097, 
        N67096, N67095, N67094, N67093, N67092}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__332, SYNOPSYS_UNCONNECTED__333, 
        SYNOPSYS_UNCONNECTED__334, SYNOPSYS_UNCONNECTED__335, 
        SYNOPSYS_UNCONNECTED__336, N68178, N68177, N68176, N68175, N68174, 
        N68173, N68172, N68171}) );
  hamming_N16000_CC2_DW01_add_84 add_2750_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67058, N67057, N67056, N67055, N67054, 
        N67053}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67071, N67070, 
        N67069, N67068, N67067, N67066}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__337, SYNOPSYS_UNCONNECTED__338, 
        SYNOPSYS_UNCONNECTED__339, SYNOPSYS_UNCONNECTED__340, 
        SYNOPSYS_UNCONNECTED__341, SYNOPSYS_UNCONNECTED__342, N68164, N68163, 
        N68162, N68161, N68160, N68159, N68158}) );
  hamming_N16000_CC2_DW01_add_85 add_2751_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67032, N67031, N67030, N67029, N67028, 
        N67027}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67045, N67044, 
        N67043, N67042, N67041, N67040}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__343, SYNOPSYS_UNCONNECTED__344, 
        SYNOPSYS_UNCONNECTED__345, SYNOPSYS_UNCONNECTED__346, 
        SYNOPSYS_UNCONNECTED__347, SYNOPSYS_UNCONNECTED__348, N68151, N68150, 
        N68149, N68148, N68147, N68146, N68145}) );
  hamming_N16000_CC2_DW01_add_86 add_2752_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67006, N67005, N67004, N67003, N67002, 
        N67001}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N67019, N67018, 
        N67017, N67016, N67015, N67014}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__349, SYNOPSYS_UNCONNECTED__350, 
        SYNOPSYS_UNCONNECTED__351, SYNOPSYS_UNCONNECTED__352, 
        SYNOPSYS_UNCONNECTED__353, SYNOPSYS_UNCONNECTED__354, N68138, N68137, 
        N68136, N68135, N68134, N68133, N68132}) );
  hamming_N16000_CC2_DW01_add_87 add_2753_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66980, N66979, N66978, N66977, N66976, 
        N66975}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66993, N66992, 
        N66991, N66990, N66989, N66988}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__355, SYNOPSYS_UNCONNECTED__356, 
        SYNOPSYS_UNCONNECTED__357, SYNOPSYS_UNCONNECTED__358, 
        SYNOPSYS_UNCONNECTED__359, SYNOPSYS_UNCONNECTED__360, N68125, N68124, 
        N68123, N68122, N68121, N68120, N68119}) );
  hamming_N16000_CC2_DW01_add_88 add_2754_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66954, N66953, N66952, N66951, N66950, 
        N66949}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66967, N66966, 
        N66965, N66964, N66963, N66962}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__361, SYNOPSYS_UNCONNECTED__362, 
        SYNOPSYS_UNCONNECTED__363, SYNOPSYS_UNCONNECTED__364, 
        SYNOPSYS_UNCONNECTED__365, SYNOPSYS_UNCONNECTED__366, N68112, N68111, 
        N68110, N68109, N68108, N68107, N68106}) );
  hamming_N16000_CC2_DW01_add_89 add_2755_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66928, N66927, N66926, N66925, N66924, 
        N66923}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66941, N66940, 
        N66939, N66938, N66937, N66936}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__367, SYNOPSYS_UNCONNECTED__368, 
        SYNOPSYS_UNCONNECTED__369, SYNOPSYS_UNCONNECTED__370, 
        SYNOPSYS_UNCONNECTED__371, SYNOPSYS_UNCONNECTED__372, N68099, N68098, 
        N68097, N68096, N68095, N68094, N68093}) );
  hamming_N16000_CC2_DW01_add_90 add_2756_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66902, N66901, N66900, N66899, N66898, 
        N66897}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66915, N66914, 
        N66913, N66912, N66911, N66910}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__373, SYNOPSYS_UNCONNECTED__374, 
        SYNOPSYS_UNCONNECTED__375, SYNOPSYS_UNCONNECTED__376, 
        SYNOPSYS_UNCONNECTED__377, SYNOPSYS_UNCONNECTED__378, N68086, N68085, 
        N68084, N68083, N68082, N68081, N68080}) );
  hamming_N16000_CC2_DW01_add_91 add_2757_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66876, N66875, N66874, N66873, N66872, 
        N66871}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66889, N66888, 
        N66887, N66886, N66885, N66884}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__379, SYNOPSYS_UNCONNECTED__380, 
        SYNOPSYS_UNCONNECTED__381, SYNOPSYS_UNCONNECTED__382, 
        SYNOPSYS_UNCONNECTED__383, SYNOPSYS_UNCONNECTED__384, N68073, N68072, 
        N68071, N68070, N68069, N68068, N68067}) );
  hamming_N16000_CC2_DW01_add_92 add_2758_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66850, N66849, N66848, N66847, N66846, 
        N66845}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66863, N66862, 
        N66861, N66860, N66859, N66858}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__385, SYNOPSYS_UNCONNECTED__386, 
        SYNOPSYS_UNCONNECTED__387, SYNOPSYS_UNCONNECTED__388, 
        SYNOPSYS_UNCONNECTED__389, SYNOPSYS_UNCONNECTED__390, N68060, N68059, 
        N68058, N68057, N68056, N68055, N68054}) );
  hamming_N16000_CC2_DW01_add_93 add_2759_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66824, N66823, N66822, N66821, N66820, 
        N66819}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66837, N66836, 
        N66835, N66834, N66833, N66832}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__391, SYNOPSYS_UNCONNECTED__392, 
        SYNOPSYS_UNCONNECTED__393, SYNOPSYS_UNCONNECTED__394, 
        SYNOPSYS_UNCONNECTED__395, SYNOPSYS_UNCONNECTED__396, N68047, N68046, 
        N68045, N68044, N68043, N68042, N68041}) );
  hamming_N16000_CC2_DW01_add_94 add_2760_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66798, N66797, N66796, N66795, N66794, 
        N66793}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66811, N66810, 
        N66809, N66808, N66807, N66806}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__397, SYNOPSYS_UNCONNECTED__398, 
        SYNOPSYS_UNCONNECTED__399, SYNOPSYS_UNCONNECTED__400, 
        SYNOPSYS_UNCONNECTED__401, SYNOPSYS_UNCONNECTED__402, N68034, N68033, 
        N68032, N68031, N68030, N68029, N68028}) );
  hamming_N16000_CC2_DW01_add_95 add_2761_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66772, N66771, N66770, N66769, N66768, 
        N66767}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66785, N66784, 
        N66783, N66782, N66781, N66780}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__403, SYNOPSYS_UNCONNECTED__404, 
        SYNOPSYS_UNCONNECTED__405, SYNOPSYS_UNCONNECTED__406, 
        SYNOPSYS_UNCONNECTED__407, SYNOPSYS_UNCONNECTED__408, N68021, N68020, 
        N68019, N68018, N68017, N68016, N68015}) );
  hamming_N16000_CC2_DW01_add_96 add_2762_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66746, N66745, N66744, N66743, N66742, 
        N66741}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66759, N66758, 
        N66757, N66756, N66755, N66754}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__409, SYNOPSYS_UNCONNECTED__410, 
        SYNOPSYS_UNCONNECTED__411, SYNOPSYS_UNCONNECTED__412, 
        SYNOPSYS_UNCONNECTED__413, SYNOPSYS_UNCONNECTED__414, N68008, N68007, 
        N68006, N68005, N68004, N68003, N68002}) );
  hamming_N16000_CC2_DW01_add_97 add_2763_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66720, N66719, N66718, N66717, N66716, 
        N66715}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66733, N66732, 
        N66731, N66730, N66729, N66728}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__415, SYNOPSYS_UNCONNECTED__416, 
        SYNOPSYS_UNCONNECTED__417, SYNOPSYS_UNCONNECTED__418, 
        SYNOPSYS_UNCONNECTED__419, SYNOPSYS_UNCONNECTED__420, N67995, N67994, 
        N67993, N67992, N67991, N67990, N67989}) );
  hamming_N16000_CC2_DW01_add_98 add_2764_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66694, N66693, N66692, N66691, N66690, 
        N66689}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66707, N66706, 
        N66705, N66704, N66703, N66702}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__421, SYNOPSYS_UNCONNECTED__422, 
        SYNOPSYS_UNCONNECTED__423, SYNOPSYS_UNCONNECTED__424, 
        SYNOPSYS_UNCONNECTED__425, SYNOPSYS_UNCONNECTED__426, N67982, N67981, 
        N67980, N67979, N67978, N67977, N67976}) );
  hamming_N16000_CC2_DW01_add_99 add_2765_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66668, N66667, N66666, N66665, N66664, 
        N66663}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66681, N66680, 
        N66679, N66678, N66677, N66676}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__427, SYNOPSYS_UNCONNECTED__428, 
        SYNOPSYS_UNCONNECTED__429, SYNOPSYS_UNCONNECTED__430, 
        SYNOPSYS_UNCONNECTED__431, SYNOPSYS_UNCONNECTED__432, N67969, N67968, 
        N67967, N67966, N67965, N67964, N67963}) );
  hamming_N16000_CC2_DW01_add_100 add_2766_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66642, N66641, N66640, N66639, N66638, 
        N66637}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66655, N66654, 
        N66653, N66652, N66651, N66650}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__433, SYNOPSYS_UNCONNECTED__434, 
        SYNOPSYS_UNCONNECTED__435, SYNOPSYS_UNCONNECTED__436, 
        SYNOPSYS_UNCONNECTED__437, SYNOPSYS_UNCONNECTED__438, N67956, N67955, 
        N67954, N67953, N67952, N67951, N67950}) );
  hamming_N16000_CC2_DW01_add_101 add_2767_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66616, N66615, N66614, N66613, N66612, 
        N66611}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66629, N66628, 
        N66627, N66626, N66625, N66624}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__439, SYNOPSYS_UNCONNECTED__440, 
        SYNOPSYS_UNCONNECTED__441, SYNOPSYS_UNCONNECTED__442, 
        SYNOPSYS_UNCONNECTED__443, SYNOPSYS_UNCONNECTED__444, N67943, N67942, 
        N67941, N67940, N67939, N67938, N67937}) );
  hamming_N16000_CC2_DW01_add_102 add_2768_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66590, N66589, N66588, N66587, N66586, 
        N66585}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66603, N66602, 
        N66601, N66600, N66599, N66598}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__445, SYNOPSYS_UNCONNECTED__446, 
        SYNOPSYS_UNCONNECTED__447, SYNOPSYS_UNCONNECTED__448, 
        SYNOPSYS_UNCONNECTED__449, SYNOPSYS_UNCONNECTED__450, N67930, N67929, 
        N67928, N67927, N67926, N67925, N67924}) );
  hamming_N16000_CC2_DW01_add_103 add_2769_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66564, N66563, N66562, N66561, N66560, 
        N66559}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66577, N66576, 
        N66575, N66574, N66573, N66572}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__451, SYNOPSYS_UNCONNECTED__452, 
        SYNOPSYS_UNCONNECTED__453, SYNOPSYS_UNCONNECTED__454, 
        SYNOPSYS_UNCONNECTED__455, SYNOPSYS_UNCONNECTED__456, N67917, N67916, 
        N67915, N67914, N67913, N67912, N67911}) );
  hamming_N16000_CC2_DW01_add_104 add_2770_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66538, N66537, N66536, N66535, N66534, 
        N66533}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66551, N66550, 
        N66549, N66548, N66547, N66546}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__457, SYNOPSYS_UNCONNECTED__458, 
        SYNOPSYS_UNCONNECTED__459, SYNOPSYS_UNCONNECTED__460, 
        SYNOPSYS_UNCONNECTED__461, SYNOPSYS_UNCONNECTED__462, N67904, N67903, 
        N67902, N67901, N67900, N67899, N67898}) );
  hamming_N16000_CC2_DW01_add_105 add_2771_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66512, N66511, N66510, N66509, N66508, 
        N66507}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66525, N66524, 
        N66523, N66522, N66521, N66520}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__463, SYNOPSYS_UNCONNECTED__464, 
        SYNOPSYS_UNCONNECTED__465, SYNOPSYS_UNCONNECTED__466, 
        SYNOPSYS_UNCONNECTED__467, SYNOPSYS_UNCONNECTED__468, N67891, N67890, 
        N67889, N67888, N67887, N67886, N67885}) );
  hamming_N16000_CC2_DW01_add_106 add_2772_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66486, N66485, N66484, N66483, N66482, 
        N66481}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66499, N66498, 
        N66497, N66496, N66495, N66494}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__469, SYNOPSYS_UNCONNECTED__470, 
        SYNOPSYS_UNCONNECTED__471, SYNOPSYS_UNCONNECTED__472, 
        SYNOPSYS_UNCONNECTED__473, SYNOPSYS_UNCONNECTED__474, N67878, N67877, 
        N67876, N67875, N67874, N67873, N67872}) );
  hamming_N16000_CC2_DW01_add_107 add_2773_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66460, N66459, N66458, N66457, N66456, 
        N66455}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66473, N66472, 
        N66471, N66470, N66469, N66468}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__475, SYNOPSYS_UNCONNECTED__476, 
        SYNOPSYS_UNCONNECTED__477, SYNOPSYS_UNCONNECTED__478, 
        SYNOPSYS_UNCONNECTED__479, SYNOPSYS_UNCONNECTED__480, N67865, N67864, 
        N67863, N67862, N67861, N67860, N67859}) );
  hamming_N16000_CC2_DW01_add_108 add_2774_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66434, N66433, N66432, N66431, N66430, 
        N66429}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66447, N66446, 
        N66445, N66444, N66443, N66442}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__481, SYNOPSYS_UNCONNECTED__482, 
        SYNOPSYS_UNCONNECTED__483, SYNOPSYS_UNCONNECTED__484, 
        SYNOPSYS_UNCONNECTED__485, SYNOPSYS_UNCONNECTED__486, N67852, N67851, 
        N67850, N67849, N67848, N67847, N67846}) );
  hamming_N16000_CC2_DW01_add_109 add_2775_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66408, N66407, N66406, N66405, N66404, 
        N66403}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66421, N66420, 
        N66419, N66418, N66417, N66416}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__487, SYNOPSYS_UNCONNECTED__488, 
        SYNOPSYS_UNCONNECTED__489, SYNOPSYS_UNCONNECTED__490, 
        SYNOPSYS_UNCONNECTED__491, SYNOPSYS_UNCONNECTED__492, N67839, N67838, 
        N67837, N67836, N67835, N67834, N67833}) );
  hamming_N16000_CC2_DW01_add_110 add_2776_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66382, N66381, N66380, N66379, N66378, 
        N66377}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66395, N66394, 
        N66393, N66392, N66391, N66390}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__493, SYNOPSYS_UNCONNECTED__494, 
        SYNOPSYS_UNCONNECTED__495, SYNOPSYS_UNCONNECTED__496, 
        SYNOPSYS_UNCONNECTED__497, SYNOPSYS_UNCONNECTED__498, N67826, N67825, 
        N67824, N67823, N67822, N67821, N67820}) );
  hamming_N16000_CC2_DW01_add_111 add_2777_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66356, N66355, N66354, N66353, N66352, 
        N66351}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66369, N66368, 
        N66367, N66366, N66365, N66364}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__499, SYNOPSYS_UNCONNECTED__500, 
        SYNOPSYS_UNCONNECTED__501, SYNOPSYS_UNCONNECTED__502, 
        SYNOPSYS_UNCONNECTED__503, SYNOPSYS_UNCONNECTED__504, N67813, N67812, 
        N67811, N67810, N67809, N67808, N67807}) );
  hamming_N16000_CC2_DW01_add_112 add_2778_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66330, N66329, N66328, N66327, N66326, 
        N66325}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66343, N66342, 
        N66341, N66340, N66339, N66338}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__505, SYNOPSYS_UNCONNECTED__506, 
        SYNOPSYS_UNCONNECTED__507, SYNOPSYS_UNCONNECTED__508, 
        SYNOPSYS_UNCONNECTED__509, SYNOPSYS_UNCONNECTED__510, N67800, N67799, 
        N67798, N67797, N67796, N67795, N67794}) );
  hamming_N16000_CC2_DW01_add_113 add_2779_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66304, N66303, N66302, N66301, N66300, 
        N66299}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66317, N66316, 
        N66315, N66314, N66313, N66312}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__511, SYNOPSYS_UNCONNECTED__512, 
        SYNOPSYS_UNCONNECTED__513, SYNOPSYS_UNCONNECTED__514, 
        SYNOPSYS_UNCONNECTED__515, SYNOPSYS_UNCONNECTED__516, N67787, N67786, 
        N67785, N67784, N67783, N67782, N67781}) );
  hamming_N16000_CC2_DW01_add_114 add_2780_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66278, N66277, N66276, N66275, N66274, 
        N66273}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66291, N66290, 
        N66289, N66288, N66287, N66286}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__517, SYNOPSYS_UNCONNECTED__518, 
        SYNOPSYS_UNCONNECTED__519, SYNOPSYS_UNCONNECTED__520, 
        SYNOPSYS_UNCONNECTED__521, SYNOPSYS_UNCONNECTED__522, N67774, N67773, 
        N67772, N67771, N67770, N67769, N67768}) );
  hamming_N16000_CC2_DW01_add_115 add_2781_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66252, N66251, N66250, N66249, N66248, 
        N66247}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66265, N66264, 
        N66263, N66262, N66261, N66260}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__523, SYNOPSYS_UNCONNECTED__524, 
        SYNOPSYS_UNCONNECTED__525, SYNOPSYS_UNCONNECTED__526, 
        SYNOPSYS_UNCONNECTED__527, SYNOPSYS_UNCONNECTED__528, N67761, N67760, 
        N67759, N67758, N67757, N67756, N67755}) );
  hamming_N16000_CC2_DW01_add_116 add_2782_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66226, N66225, N66224, N66223, N66222, 
        N66221}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66239, N66238, 
        N66237, N66236, N66235, N66234}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__529, SYNOPSYS_UNCONNECTED__530, 
        SYNOPSYS_UNCONNECTED__531, SYNOPSYS_UNCONNECTED__532, 
        SYNOPSYS_UNCONNECTED__533, SYNOPSYS_UNCONNECTED__534, N67748, N67747, 
        N67746, N67745, N67744, N67743, N67742}) );
  hamming_N16000_CC2_DW01_add_117 add_2783_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66200, N66199, N66198, N66197, N66196, 
        N66195}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66213, N66212, 
        N66211, N66210, N66209, N66208}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__535, SYNOPSYS_UNCONNECTED__536, 
        SYNOPSYS_UNCONNECTED__537, SYNOPSYS_UNCONNECTED__538, 
        SYNOPSYS_UNCONNECTED__539, SYNOPSYS_UNCONNECTED__540, N67735, N67734, 
        N67733, N67732, N67731, N67730, N67729}) );
  hamming_N16000_CC2_DW01_add_118 add_2784_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66174, N66173, N66172, N66171, N66170, 
        N66169}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66187, N66186, 
        N66185, N66184, N66183, N66182}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__541, SYNOPSYS_UNCONNECTED__542, 
        SYNOPSYS_UNCONNECTED__543, SYNOPSYS_UNCONNECTED__544, 
        SYNOPSYS_UNCONNECTED__545, SYNOPSYS_UNCONNECTED__546, N67722, N67721, 
        N67720, N67719, N67718, N67717, N67716}) );
  hamming_N16000_CC2_DW01_add_119 add_2785_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66148, N66147, N66146, N66145, N66144, 
        N66143}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66161, N66160, 
        N66159, N66158, N66157, N66156}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__547, SYNOPSYS_UNCONNECTED__548, 
        SYNOPSYS_UNCONNECTED__549, SYNOPSYS_UNCONNECTED__550, 
        SYNOPSYS_UNCONNECTED__551, SYNOPSYS_UNCONNECTED__552, N67709, N67708, 
        N67707, N67706, N67705, N67704, N67703}) );
  hamming_N16000_CC2_DW01_add_120 add_2786_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66122, N66121, N66120, N66119, N66118, 
        N66117}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66135, N66134, 
        N66133, N66132, N66131, N66130}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__553, SYNOPSYS_UNCONNECTED__554, 
        SYNOPSYS_UNCONNECTED__555, SYNOPSYS_UNCONNECTED__556, 
        SYNOPSYS_UNCONNECTED__557, SYNOPSYS_UNCONNECTED__558, N67696, N67695, 
        N67694, N67693, N67692, N67691, N67690}) );
  hamming_N16000_CC2_DW01_add_121 add_2787_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66096, N66095, N66094, N66093, N66092, 
        N66091}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66109, N66108, 
        N66107, N66106, N66105, N66104}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__559, SYNOPSYS_UNCONNECTED__560, 
        SYNOPSYS_UNCONNECTED__561, SYNOPSYS_UNCONNECTED__562, 
        SYNOPSYS_UNCONNECTED__563, SYNOPSYS_UNCONNECTED__564, N67683, N67682, 
        N67681, N67680, N67679, N67678, N67677}) );
  hamming_N16000_CC2_DW01_add_122 add_2788_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66070, N66069, N66068, N66067, N66066, 
        N66065}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66083, N66082, 
        N66081, N66080, N66079, N66078}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__565, SYNOPSYS_UNCONNECTED__566, 
        SYNOPSYS_UNCONNECTED__567, SYNOPSYS_UNCONNECTED__568, 
        SYNOPSYS_UNCONNECTED__569, SYNOPSYS_UNCONNECTED__570, N67670, N67669, 
        N67668, N67667, N67666, N67665, N67664}) );
  hamming_N16000_CC2_DW01_add_123 add_2789_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66044, N66043, N66042, N66041, N66040, 
        N66039}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66057, N66056, 
        N66055, N66054, N66053, N66052}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__571, SYNOPSYS_UNCONNECTED__572, 
        SYNOPSYS_UNCONNECTED__573, SYNOPSYS_UNCONNECTED__574, 
        SYNOPSYS_UNCONNECTED__575, SYNOPSYS_UNCONNECTED__576, N67657, N67656, 
        N67655, N67654, N67653, N67652, N67651}) );
  hamming_N16000_CC2_DW01_add_124 add_2790_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66018, N66017, N66016, N66015, N66014, 
        N66013}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66031, N66030, 
        N66029, N66028, N66027, N66026}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__577, SYNOPSYS_UNCONNECTED__578, 
        SYNOPSYS_UNCONNECTED__579, SYNOPSYS_UNCONNECTED__580, 
        SYNOPSYS_UNCONNECTED__581, SYNOPSYS_UNCONNECTED__582, N67644, N67643, 
        N67642, N67641, N67640, N67639, N67638}) );
  hamming_N16000_CC2_DW01_add_125 add_2791_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65992, N65991, N65990, N65989, N65988, 
        N65987}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N66005, N66004, 
        N66003, N66002, N66001, N66000}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__583, SYNOPSYS_UNCONNECTED__584, 
        SYNOPSYS_UNCONNECTED__585, SYNOPSYS_UNCONNECTED__586, 
        SYNOPSYS_UNCONNECTED__587, SYNOPSYS_UNCONNECTED__588, N67631, N67630, 
        N67629, N67628, N67627, N67626, N67625}) );
  hamming_N16000_CC2_DW01_add_126 add_2792_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65966, N65965, N65964, N65963, N65962, 
        N65961}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65979, N65978, 
        N65977, N65976, N65975, N65974}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__589, SYNOPSYS_UNCONNECTED__590, 
        SYNOPSYS_UNCONNECTED__591, SYNOPSYS_UNCONNECTED__592, 
        SYNOPSYS_UNCONNECTED__593, SYNOPSYS_UNCONNECTED__594, N67618, N67617, 
        N67616, N67615, N67614, N67613, N67612}) );
  hamming_N16000_CC2_DW01_add_127 add_2793_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65940, N65939, N65938, N65937, N65936, 
        N65935}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65953, N65952, 
        N65951, N65950, N65949, N65948}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__595, SYNOPSYS_UNCONNECTED__596, 
        SYNOPSYS_UNCONNECTED__597, SYNOPSYS_UNCONNECTED__598, 
        SYNOPSYS_UNCONNECTED__599, SYNOPSYS_UNCONNECTED__600, N67605, N67604, 
        N67603, N67602, N67601, N67600, N67599}) );
  hamming_N16000_CC2_DW01_add_128 add_2794_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65914, N65913, N65912, N65911, N65910, 
        N65909}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65927, N65926, 
        N65925, N65924, N65923, N65922}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__601, SYNOPSYS_UNCONNECTED__602, 
        SYNOPSYS_UNCONNECTED__603, SYNOPSYS_UNCONNECTED__604, 
        SYNOPSYS_UNCONNECTED__605, SYNOPSYS_UNCONNECTED__606, N67592, N67591, 
        N67590, N67589, N67588, N67587, N67586}) );
  hamming_N16000_CC2_DW01_add_129 add_2795_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65888, N65887, N65886, N65885, N65884, 
        N65883}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65901, N65900, 
        N65899, N65898, N65897, N65896}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__607, SYNOPSYS_UNCONNECTED__608, 
        SYNOPSYS_UNCONNECTED__609, SYNOPSYS_UNCONNECTED__610, 
        SYNOPSYS_UNCONNECTED__611, SYNOPSYS_UNCONNECTED__612, N67579, N67578, 
        N67577, N67576, N67575, N67574, N67573}) );
  hamming_N16000_CC2_DW01_add_130 add_2796_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65862, N65861, N65860, N65859, N65858, 
        N65857}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65875, N65874, 
        N65873, N65872, N65871, N65870}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__613, SYNOPSYS_UNCONNECTED__614, 
        SYNOPSYS_UNCONNECTED__615, SYNOPSYS_UNCONNECTED__616, 
        SYNOPSYS_UNCONNECTED__617, SYNOPSYS_UNCONNECTED__618, N67566, N67565, 
        N67564, N67563, N67562, N67561, N67560}) );
  hamming_N16000_CC2_DW01_add_131 add_2797_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65836, N65835, N65834, N65833, N65832, 
        N65831}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65849, N65848, 
        N65847, N65846, N65845, N65844}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__619, SYNOPSYS_UNCONNECTED__620, 
        SYNOPSYS_UNCONNECTED__621, SYNOPSYS_UNCONNECTED__622, 
        SYNOPSYS_UNCONNECTED__623, SYNOPSYS_UNCONNECTED__624, N67553, N67552, 
        N67551, N67550, N67549, N67548, N67547}) );
  hamming_N16000_CC2_DW01_add_132 add_2798_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65810, N65809, N65808, N65807, N65806, 
        N65805}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65823, N65822, 
        N65821, N65820, N65819, N65818}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__625, SYNOPSYS_UNCONNECTED__626, 
        SYNOPSYS_UNCONNECTED__627, SYNOPSYS_UNCONNECTED__628, 
        SYNOPSYS_UNCONNECTED__629, SYNOPSYS_UNCONNECTED__630, N67540, N67539, 
        N67538, N67537, N67536, N67535, N67534}) );
  hamming_N16000_CC2_DW01_add_133 add_2799_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65784, N65783, N65782, N65781, N65780, 
        N65779}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65797, N65796, 
        N65795, N65794, N65793, N65792}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__631, SYNOPSYS_UNCONNECTED__632, 
        SYNOPSYS_UNCONNECTED__633, SYNOPSYS_UNCONNECTED__634, 
        SYNOPSYS_UNCONNECTED__635, SYNOPSYS_UNCONNECTED__636, N67527, N67526, 
        N67525, N67524, N67523, N67522, N67521}) );
  hamming_N16000_CC2_DW01_add_134 add_2800_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65758, N65757, N65756, N65755, N65754, 
        N65753}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65771, N65770, 
        N65769, N65768, N65767, N65766}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__637, SYNOPSYS_UNCONNECTED__638, 
        SYNOPSYS_UNCONNECTED__639, SYNOPSYS_UNCONNECTED__640, 
        SYNOPSYS_UNCONNECTED__641, SYNOPSYS_UNCONNECTED__642, N67514, N67513, 
        N67512, N67511, N67510, N67509, N67508}) );
  hamming_N16000_CC2_DW01_add_135 add_2801_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65732, N65731, N65730, N65729, N65728, 
        N65727}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65745, N65744, 
        N65743, N65742, N65741, N65740}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__643, SYNOPSYS_UNCONNECTED__644, 
        SYNOPSYS_UNCONNECTED__645, SYNOPSYS_UNCONNECTED__646, 
        SYNOPSYS_UNCONNECTED__647, SYNOPSYS_UNCONNECTED__648, N67501, N67500, 
        N67499, N67498, N67497, N67496, N67495}) );
  hamming_N16000_CC2_DW01_add_136 add_2802_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65706, N65705, N65704, N65703, N65702, 
        N65701}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65719, N65718, 
        N65717, N65716, N65715, N65714}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__649, SYNOPSYS_UNCONNECTED__650, 
        SYNOPSYS_UNCONNECTED__651, SYNOPSYS_UNCONNECTED__652, 
        SYNOPSYS_UNCONNECTED__653, SYNOPSYS_UNCONNECTED__654, N67488, N67487, 
        N67486, N67485, N67484, N67483, N67482}) );
  hamming_N16000_CC2_DW01_add_137 add_2803_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65680, N65679, N65678, N65677, N65676, 
        N65675}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65693, N65692, 
        N65691, N65690, N65689, N65688}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__655, SYNOPSYS_UNCONNECTED__656, 
        SYNOPSYS_UNCONNECTED__657, SYNOPSYS_UNCONNECTED__658, 
        SYNOPSYS_UNCONNECTED__659, SYNOPSYS_UNCONNECTED__660, N67475, N67474, 
        N67473, N67472, N67471, N67470, N67469}) );
  hamming_N16000_CC2_DW01_add_138 add_2804_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65654, N65653, N65652, N65651, N65650, 
        N65649}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65667, N65666, 
        N65665, N65664, N65663, N65662}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__661, SYNOPSYS_UNCONNECTED__662, 
        SYNOPSYS_UNCONNECTED__663, SYNOPSYS_UNCONNECTED__664, 
        SYNOPSYS_UNCONNECTED__665, SYNOPSYS_UNCONNECTED__666, N67462, N67461, 
        N67460, N67459, N67458, N67457, N67456}) );
  hamming_N16000_CC2_DW01_add_139 add_2805_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65628, N65627, N65626, N65625, N65624, 
        N65623}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65641, N65640, 
        N65639, N65638, N65637, N65636}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__667, SYNOPSYS_UNCONNECTED__668, 
        SYNOPSYS_UNCONNECTED__669, SYNOPSYS_UNCONNECTED__670, 
        SYNOPSYS_UNCONNECTED__671, SYNOPSYS_UNCONNECTED__672, N67449, N67448, 
        N67447, N67446, N67445, N67444, N67443}) );
  hamming_N16000_CC2_DW01_add_140 add_2806_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65602, N65601, N65600, N65599, N65598, 
        N65597}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65615, N65614, 
        N65613, N65612, N65611, N65610}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__673, SYNOPSYS_UNCONNECTED__674, 
        SYNOPSYS_UNCONNECTED__675, SYNOPSYS_UNCONNECTED__676, 
        SYNOPSYS_UNCONNECTED__677, SYNOPSYS_UNCONNECTED__678, N67436, N67435, 
        N67434, N67433, N67432, N67431, N67430}) );
  hamming_N16000_CC2_DW01_add_141 add_2807_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65576, N65575, N65574, N65573, N65572, 
        N65571}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65589, N65588, 
        N65587, N65586, N65585, N65584}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__679, SYNOPSYS_UNCONNECTED__680, 
        SYNOPSYS_UNCONNECTED__681, SYNOPSYS_UNCONNECTED__682, 
        SYNOPSYS_UNCONNECTED__683, SYNOPSYS_UNCONNECTED__684, N67423, N67422, 
        N67421, N67420, N67419, N67418, N67417}) );
  hamming_N16000_CC2_DW01_add_142 add_2808_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65550, N65549, N65548, N65547, N65546, 
        N65545}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65563, N65562, 
        N65561, N65560, N65559, N65558}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__685, SYNOPSYS_UNCONNECTED__686, 
        SYNOPSYS_UNCONNECTED__687, SYNOPSYS_UNCONNECTED__688, 
        SYNOPSYS_UNCONNECTED__689, SYNOPSYS_UNCONNECTED__690, N67410, N67409, 
        N67408, N67407, N67406, N67405, N67404}) );
  hamming_N16000_CC2_DW01_add_143 add_2809_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65524, N65523, N65522, N65521, N65520, 
        N65519}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65537, N65536, 
        N65535, N65534, N65533, N65532}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__691, SYNOPSYS_UNCONNECTED__692, 
        SYNOPSYS_UNCONNECTED__693, SYNOPSYS_UNCONNECTED__694, 
        SYNOPSYS_UNCONNECTED__695, SYNOPSYS_UNCONNECTED__696, N67397, N67396, 
        N67395, N67394, N67393, N67392, N67391}) );
  hamming_N16000_CC2_DW01_add_144 add_2810_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65498, N65497, N65496, N65495, N65494, 
        N65493}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65511, N65510, 
        N65509, N65508, N65507, N65506}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__697, SYNOPSYS_UNCONNECTED__698, 
        SYNOPSYS_UNCONNECTED__699, SYNOPSYS_UNCONNECTED__700, 
        SYNOPSYS_UNCONNECTED__701, SYNOPSYS_UNCONNECTED__702, N67384, N67383, 
        N67382, N67381, N67380, N67379, N67378}) );
  hamming_N16000_CC2_DW01_add_145 add_2811_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65472, N65471, N65470, N65469, N65468, 
        N65467}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65485, N65484, 
        N65483, N65482, N65481, N65480}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__703, SYNOPSYS_UNCONNECTED__704, 
        SYNOPSYS_UNCONNECTED__705, SYNOPSYS_UNCONNECTED__706, 
        SYNOPSYS_UNCONNECTED__707, SYNOPSYS_UNCONNECTED__708, N67371, N67370, 
        N67369, N67368, N67367, N67366, N67365}) );
  hamming_N16000_CC2_DW01_add_146 add_2812_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65446, N65445, N65444, N65443, N65442, 
        N65441}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65459, N65458, 
        N65457, N65456, N65455, N65454}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__709, SYNOPSYS_UNCONNECTED__710, 
        SYNOPSYS_UNCONNECTED__711, SYNOPSYS_UNCONNECTED__712, 
        SYNOPSYS_UNCONNECTED__713, SYNOPSYS_UNCONNECTED__714, N67358, N67357, 
        N67356, N67355, N67354, N67353, N67352}) );
  hamming_N16000_CC2_DW01_add_147 add_2813_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65420, N65419, N65418, N65417, N65416, 
        N65415}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65433, N65432, 
        N65431, N65430, N65429, N65428}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__715, SYNOPSYS_UNCONNECTED__716, 
        SYNOPSYS_UNCONNECTED__717, SYNOPSYS_UNCONNECTED__718, 
        SYNOPSYS_UNCONNECTED__719, SYNOPSYS_UNCONNECTED__720, N67345, N67344, 
        N67343, N67342, N67341, N67340, N67339}) );
  hamming_N16000_CC2_DW01_add_148 add_2814_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65394, N65393, N65392, N65391, N65390, 
        N65389}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65407, N65406, 
        N65405, N65404, N65403, N65402}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__721, SYNOPSYS_UNCONNECTED__722, 
        SYNOPSYS_UNCONNECTED__723, SYNOPSYS_UNCONNECTED__724, 
        SYNOPSYS_UNCONNECTED__725, SYNOPSYS_UNCONNECTED__726, N67332, N67331, 
        N67330, N67329, N67328, N67327, N67326}) );
  hamming_N16000_CC2_DW01_add_149 add_2815_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65368, N65367, N65366, N65365, N65364, 
        N65363}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65381, N65380, 
        N65379, N65378, N65377, N65376}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__727, SYNOPSYS_UNCONNECTED__728, 
        SYNOPSYS_UNCONNECTED__729, SYNOPSYS_UNCONNECTED__730, 
        SYNOPSYS_UNCONNECTED__731, SYNOPSYS_UNCONNECTED__732, N67319, N67318, 
        N67317, N67316, N67315, N67314, N67313}) );
  hamming_N16000_CC2_DW01_add_150 add_2816_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65342, N65341, N65340, N65339, N65338, 
        N65337}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65355, N65354, 
        N65353, N65352, N65351, N65350}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__733, SYNOPSYS_UNCONNECTED__734, 
        SYNOPSYS_UNCONNECTED__735, SYNOPSYS_UNCONNECTED__736, 
        SYNOPSYS_UNCONNECTED__737, SYNOPSYS_UNCONNECTED__738, N67306, N67305, 
        N67304, N67303, N67302, N67301, N67300}) );
  hamming_N16000_CC2_DW01_add_151 add_2817_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65316, N65315, N65314, N65313, N65312, 
        N65311}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65329, N65328, 
        N65327, N65326, N65325, N65324}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__739, SYNOPSYS_UNCONNECTED__740, 
        SYNOPSYS_UNCONNECTED__741, SYNOPSYS_UNCONNECTED__742, 
        SYNOPSYS_UNCONNECTED__743, SYNOPSYS_UNCONNECTED__744, N67293, N67292, 
        N67291, N67290, N67289, N67288, N67287}) );
  hamming_N16000_CC2_DW01_add_152 add_2818_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65290, N65289, N65288, N65287, N65286, 
        N65285}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65303, N65302, 
        N65301, N65300, N65299, N65298}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__745, SYNOPSYS_UNCONNECTED__746, 
        SYNOPSYS_UNCONNECTED__747, SYNOPSYS_UNCONNECTED__748, 
        SYNOPSYS_UNCONNECTED__749, SYNOPSYS_UNCONNECTED__750, N67280, N67279, 
        N67278, N67277, N67276, N67275, N67274}) );
  hamming_N16000_CC2_DW01_add_153 add_2819_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65264, N65263, N65262, N65261, N65260, 
        N65259}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65277, N65276, 
        N65275, N65274, N65273, N65272}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__751, SYNOPSYS_UNCONNECTED__752, 
        SYNOPSYS_UNCONNECTED__753, SYNOPSYS_UNCONNECTED__754, 
        SYNOPSYS_UNCONNECTED__755, SYNOPSYS_UNCONNECTED__756, N67267, N67266, 
        N67265, N67264, N67263, N67262, N67261}) );
  hamming_N16000_CC2_DW01_add_154 add_2820_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65238, N65237, N65236, N65235, N65234, 
        N65233}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65251, N65250, 
        N65249, N65248, N65247, N65246}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__757, SYNOPSYS_UNCONNECTED__758, 
        SYNOPSYS_UNCONNECTED__759, SYNOPSYS_UNCONNECTED__760, 
        SYNOPSYS_UNCONNECTED__761, SYNOPSYS_UNCONNECTED__762, N67254, N67253, 
        N67252, N67251, N67250, N67249, N67248}) );
  hamming_N16000_CC2_DW01_add_155 add_2821_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65212, N65211, N65210, N65209, N65208, 
        N65207}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65225, N65224, 
        N65223, N65222, N65221, N65220}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__763, SYNOPSYS_UNCONNECTED__764, 
        SYNOPSYS_UNCONNECTED__765, SYNOPSYS_UNCONNECTED__766, 
        SYNOPSYS_UNCONNECTED__767, SYNOPSYS_UNCONNECTED__768, N67241, N67240, 
        N67239, N67238, N67237, N67236, N67235}) );
  hamming_N16000_CC2_DW01_add_156 add_2822_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65186, N65185, N65184, N65183, N65182, 
        N65181}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65199, N65198, 
        N65197, N65196, N65195, N65194}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__769, SYNOPSYS_UNCONNECTED__770, 
        SYNOPSYS_UNCONNECTED__771, SYNOPSYS_UNCONNECTED__772, 
        SYNOPSYS_UNCONNECTED__773, SYNOPSYS_UNCONNECTED__774, N67228, N67227, 
        N67226, N67225, N67224, N67223, N67222}) );
  hamming_N16000_CC2_DW01_add_157 add_2823_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65160, N65159, N65158, N65157, N65156, 
        N65155}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65173, N65172, 
        N65171, N65170, N65169, N65168}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__775, SYNOPSYS_UNCONNECTED__776, 
        SYNOPSYS_UNCONNECTED__777, SYNOPSYS_UNCONNECTED__778, 
        SYNOPSYS_UNCONNECTED__779, SYNOPSYS_UNCONNECTED__780, N67215, N67214, 
        N67213, N67212, N67211, N67210, N67209}) );
  hamming_N16000_CC2_DW01_add_158 add_2824_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65134, N65133, N65132, N65131, N65130, 
        N65129}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65147, N65146, 
        N65145, N65144, N65143, N65142}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__781, SYNOPSYS_UNCONNECTED__782, 
        SYNOPSYS_UNCONNECTED__783, SYNOPSYS_UNCONNECTED__784, 
        SYNOPSYS_UNCONNECTED__785, SYNOPSYS_UNCONNECTED__786, N67202, N67201, 
        N67200, N67199, N67198, N67197, N67196}) );
  hamming_N16000_CC2_DW01_add_159 add_2825_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65108, N65107, N65106, N65105, N65104, 
        N65103}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65121, N65120, 
        N65119, N65118, N65117, N65116}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__787, SYNOPSYS_UNCONNECTED__788, 
        SYNOPSYS_UNCONNECTED__789, SYNOPSYS_UNCONNECTED__790, 
        SYNOPSYS_UNCONNECTED__791, SYNOPSYS_UNCONNECTED__792, N67189, N67188, 
        N67187, N67186, N67185, N67184, N67183}) );
  hamming_N16000_CC2_DW01_add_160 add_2826_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65082, N65081, N65080, N65079, N65078, 
        N65077}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65095, N65094, 
        N65093, N65092, N65091, N65090}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__793, SYNOPSYS_UNCONNECTED__794, 
        SYNOPSYS_UNCONNECTED__795, SYNOPSYS_UNCONNECTED__796, 
        SYNOPSYS_UNCONNECTED__797, SYNOPSYS_UNCONNECTED__798, N67176, N67175, 
        N67174, N67173, N67172, N67171, N67170}) );
  hamming_N16000_CC2_DW01_add_161 add_2827_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65056, N65055, N65054, N65053, N65052, 
        N65051}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65069, N65068, 
        N65067, N65066, N65065, N65064}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__799, SYNOPSYS_UNCONNECTED__800, 
        SYNOPSYS_UNCONNECTED__801, SYNOPSYS_UNCONNECTED__802, 
        SYNOPSYS_UNCONNECTED__803, SYNOPSYS_UNCONNECTED__804, N67163, N67162, 
        N67161, N67160, N67159, N67158, N67157}) );
  hamming_N16000_CC2_DW01_add_162 add_2828_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65030, N65029, N65028, N65027, N65026, 
        N65025}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65043, N65042, 
        N65041, N65040, N65039, N65038}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__805, SYNOPSYS_UNCONNECTED__806, 
        SYNOPSYS_UNCONNECTED__807, SYNOPSYS_UNCONNECTED__808, 
        SYNOPSYS_UNCONNECTED__809, SYNOPSYS_UNCONNECTED__810, N67150, N67149, 
        N67148, N67147, N67146, N67145, N67144}) );
  hamming_N16000_CC2_DW01_add_163 add_2829_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65004, N65003, N65002, N65001, N65000, 
        N64999}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N65017, N65016, 
        N65015, N65014, N65013, N65012}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__811, SYNOPSYS_UNCONNECTED__812, 
        SYNOPSYS_UNCONNECTED__813, SYNOPSYS_UNCONNECTED__814, 
        SYNOPSYS_UNCONNECTED__815, SYNOPSYS_UNCONNECTED__816, N67137, N67136, 
        N67135, N67134, N67133, N67132, N67131}) );
  hamming_N16000_CC2_DW01_add_164 add_2830_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64978, N64977, N64976, N64975, N64974, 
        N64973}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64991, N64990, 
        N64989, N64988, N64987, N64986}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__817, SYNOPSYS_UNCONNECTED__818, 
        SYNOPSYS_UNCONNECTED__819, SYNOPSYS_UNCONNECTED__820, 
        SYNOPSYS_UNCONNECTED__821, SYNOPSYS_UNCONNECTED__822, N67124, N67123, 
        N67122, N67121, N67120, N67119, N67118}) );
  hamming_N16000_CC2_DW01_add_165 add_2831_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64952, N64951, N64950, N64949, N64948, 
        N64947}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64965, N64964, 
        N64963, N64962, N64961, N64960}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__823, SYNOPSYS_UNCONNECTED__824, 
        SYNOPSYS_UNCONNECTED__825, SYNOPSYS_UNCONNECTED__826, 
        SYNOPSYS_UNCONNECTED__827, SYNOPSYS_UNCONNECTED__828, N67111, N67110, 
        N67109, N67108, N67107, N67106, N67105}) );
  hamming_N16000_CC2_DW01_add_166 add_2832_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64926, N64925, N64924, N64923, N64922, 
        N64921}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64939, N64938, 
        N64937, N64936, N64935, N64934}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__829, SYNOPSYS_UNCONNECTED__830, 
        SYNOPSYS_UNCONNECTED__831, SYNOPSYS_UNCONNECTED__832, 
        SYNOPSYS_UNCONNECTED__833, SYNOPSYS_UNCONNECTED__834, N67098, N67097, 
        N67096, N67095, N67094, N67093, N67092}) );
  hamming_N16000_CC2_DW01_add_167 add_2833_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64899, N64898, N64897, N64896, 
        N64895}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64912, 
        N64911, N64910, N64909, N64908}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__835, SYNOPSYS_UNCONNECTED__836, 
        SYNOPSYS_UNCONNECTED__837, SYNOPSYS_UNCONNECTED__838, 
        SYNOPSYS_UNCONNECTED__839, SYNOPSYS_UNCONNECTED__840, 
        SYNOPSYS_UNCONNECTED__841, N67084, N67083, N67082, N67081, N67080, 
        N67079}) );
  hamming_N16000_CC2_DW01_add_168 add_2834_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64873, N64872, N64871, N64870, 
        N64869}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64886, 
        N64885, N64884, N64883, N64882}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__842, SYNOPSYS_UNCONNECTED__843, 
        SYNOPSYS_UNCONNECTED__844, SYNOPSYS_UNCONNECTED__845, 
        SYNOPSYS_UNCONNECTED__846, SYNOPSYS_UNCONNECTED__847, 
        SYNOPSYS_UNCONNECTED__848, N67071, N67070, N67069, N67068, N67067, 
        N67066}) );
  hamming_N16000_CC2_DW01_add_169 add_2835_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64847, N64846, N64845, N64844, 
        N64843}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64860, 
        N64859, N64858, N64857, N64856}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__849, SYNOPSYS_UNCONNECTED__850, 
        SYNOPSYS_UNCONNECTED__851, SYNOPSYS_UNCONNECTED__852, 
        SYNOPSYS_UNCONNECTED__853, SYNOPSYS_UNCONNECTED__854, 
        SYNOPSYS_UNCONNECTED__855, N67058, N67057, N67056, N67055, N67054, 
        N67053}) );
  hamming_N16000_CC2_DW01_add_170 add_2836_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64821, N64820, N64819, N64818, 
        N64817}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64834, 
        N64833, N64832, N64831, N64830}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__856, SYNOPSYS_UNCONNECTED__857, 
        SYNOPSYS_UNCONNECTED__858, SYNOPSYS_UNCONNECTED__859, 
        SYNOPSYS_UNCONNECTED__860, SYNOPSYS_UNCONNECTED__861, 
        SYNOPSYS_UNCONNECTED__862, N67045, N67044, N67043, N67042, N67041, 
        N67040}) );
  hamming_N16000_CC2_DW01_add_171 add_2837_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64795, N64794, N64793, N64792, 
        N64791}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64808, 
        N64807, N64806, N64805, N64804}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__863, SYNOPSYS_UNCONNECTED__864, 
        SYNOPSYS_UNCONNECTED__865, SYNOPSYS_UNCONNECTED__866, 
        SYNOPSYS_UNCONNECTED__867, SYNOPSYS_UNCONNECTED__868, 
        SYNOPSYS_UNCONNECTED__869, N67032, N67031, N67030, N67029, N67028, 
        N67027}) );
  hamming_N16000_CC2_DW01_add_172 add_2838_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64769, N64768, N64767, N64766, 
        N64765}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64782, 
        N64781, N64780, N64779, N64778}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__870, SYNOPSYS_UNCONNECTED__871, 
        SYNOPSYS_UNCONNECTED__872, SYNOPSYS_UNCONNECTED__873, 
        SYNOPSYS_UNCONNECTED__874, SYNOPSYS_UNCONNECTED__875, 
        SYNOPSYS_UNCONNECTED__876, N67019, N67018, N67017, N67016, N67015, 
        N67014}) );
  hamming_N16000_CC2_DW01_add_173 add_2839_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64743, N64742, N64741, N64740, 
        N64739}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64756, 
        N64755, N64754, N64753, N64752}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__877, SYNOPSYS_UNCONNECTED__878, 
        SYNOPSYS_UNCONNECTED__879, SYNOPSYS_UNCONNECTED__880, 
        SYNOPSYS_UNCONNECTED__881, SYNOPSYS_UNCONNECTED__882, 
        SYNOPSYS_UNCONNECTED__883, N67006, N67005, N67004, N67003, N67002, 
        N67001}) );
  hamming_N16000_CC2_DW01_add_174 add_2840_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64717, N64716, N64715, N64714, 
        N64713}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64730, 
        N64729, N64728, N64727, N64726}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__884, SYNOPSYS_UNCONNECTED__885, 
        SYNOPSYS_UNCONNECTED__886, SYNOPSYS_UNCONNECTED__887, 
        SYNOPSYS_UNCONNECTED__888, SYNOPSYS_UNCONNECTED__889, 
        SYNOPSYS_UNCONNECTED__890, N66993, N66992, N66991, N66990, N66989, 
        N66988}) );
  hamming_N16000_CC2_DW01_add_175 add_2841_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64691, N64690, N64689, N64688, 
        N64687}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64704, 
        N64703, N64702, N64701, N64700}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__891, SYNOPSYS_UNCONNECTED__892, 
        SYNOPSYS_UNCONNECTED__893, SYNOPSYS_UNCONNECTED__894, 
        SYNOPSYS_UNCONNECTED__895, SYNOPSYS_UNCONNECTED__896, 
        SYNOPSYS_UNCONNECTED__897, N66980, N66979, N66978, N66977, N66976, 
        N66975}) );
  hamming_N16000_CC2_DW01_add_176 add_2842_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64665, N64664, N64663, N64662, 
        N64661}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64678, 
        N64677, N64676, N64675, N64674}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__898, SYNOPSYS_UNCONNECTED__899, 
        SYNOPSYS_UNCONNECTED__900, SYNOPSYS_UNCONNECTED__901, 
        SYNOPSYS_UNCONNECTED__902, SYNOPSYS_UNCONNECTED__903, 
        SYNOPSYS_UNCONNECTED__904, N66967, N66966, N66965, N66964, N66963, 
        N66962}) );
  hamming_N16000_CC2_DW01_add_177 add_2843_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64639, N64638, N64637, N64636, 
        N64635}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64652, 
        N64651, N64650, N64649, N64648}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__905, SYNOPSYS_UNCONNECTED__906, 
        SYNOPSYS_UNCONNECTED__907, SYNOPSYS_UNCONNECTED__908, 
        SYNOPSYS_UNCONNECTED__909, SYNOPSYS_UNCONNECTED__910, 
        SYNOPSYS_UNCONNECTED__911, N66954, N66953, N66952, N66951, N66950, 
        N66949}) );
  hamming_N16000_CC2_DW01_add_178 add_2844_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64613, N64612, N64611, N64610, 
        N64609}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64626, 
        N64625, N64624, N64623, N64622}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__912, SYNOPSYS_UNCONNECTED__913, 
        SYNOPSYS_UNCONNECTED__914, SYNOPSYS_UNCONNECTED__915, 
        SYNOPSYS_UNCONNECTED__916, SYNOPSYS_UNCONNECTED__917, 
        SYNOPSYS_UNCONNECTED__918, N66941, N66940, N66939, N66938, N66937, 
        N66936}) );
  hamming_N16000_CC2_DW01_add_179 add_2845_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64587, N64586, N64585, N64584, 
        N64583}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64600, 
        N64599, N64598, N64597, N64596}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__919, SYNOPSYS_UNCONNECTED__920, 
        SYNOPSYS_UNCONNECTED__921, SYNOPSYS_UNCONNECTED__922, 
        SYNOPSYS_UNCONNECTED__923, SYNOPSYS_UNCONNECTED__924, 
        SYNOPSYS_UNCONNECTED__925, N66928, N66927, N66926, N66925, N66924, 
        N66923}) );
  hamming_N16000_CC2_DW01_add_180 add_2846_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64561, N64560, N64559, N64558, 
        N64557}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64574, 
        N64573, N64572, N64571, N64570}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__926, SYNOPSYS_UNCONNECTED__927, 
        SYNOPSYS_UNCONNECTED__928, SYNOPSYS_UNCONNECTED__929, 
        SYNOPSYS_UNCONNECTED__930, SYNOPSYS_UNCONNECTED__931, 
        SYNOPSYS_UNCONNECTED__932, N66915, N66914, N66913, N66912, N66911, 
        N66910}) );
  hamming_N16000_CC2_DW01_add_181 add_2847_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64535, N64534, N64533, N64532, 
        N64531}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64548, 
        N64547, N64546, N64545, N64544}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__933, SYNOPSYS_UNCONNECTED__934, 
        SYNOPSYS_UNCONNECTED__935, SYNOPSYS_UNCONNECTED__936, 
        SYNOPSYS_UNCONNECTED__937, SYNOPSYS_UNCONNECTED__938, 
        SYNOPSYS_UNCONNECTED__939, N66902, N66901, N66900, N66899, N66898, 
        N66897}) );
  hamming_N16000_CC2_DW01_add_182 add_2848_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64509, N64508, N64507, N64506, 
        N64505}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64522, 
        N64521, N64520, N64519, N64518}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__940, SYNOPSYS_UNCONNECTED__941, 
        SYNOPSYS_UNCONNECTED__942, SYNOPSYS_UNCONNECTED__943, 
        SYNOPSYS_UNCONNECTED__944, SYNOPSYS_UNCONNECTED__945, 
        SYNOPSYS_UNCONNECTED__946, N66889, N66888, N66887, N66886, N66885, 
        N66884}) );
  hamming_N16000_CC2_DW01_add_183 add_2849_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64483, N64482, N64481, N64480, 
        N64479}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64496, 
        N64495, N64494, N64493, N64492}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__947, SYNOPSYS_UNCONNECTED__948, 
        SYNOPSYS_UNCONNECTED__949, SYNOPSYS_UNCONNECTED__950, 
        SYNOPSYS_UNCONNECTED__951, SYNOPSYS_UNCONNECTED__952, 
        SYNOPSYS_UNCONNECTED__953, N66876, N66875, N66874, N66873, N66872, 
        N66871}) );
  hamming_N16000_CC2_DW01_add_184 add_2850_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64457, N64456, N64455, N64454, 
        N64453}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64470, 
        N64469, N64468, N64467, N64466}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__954, SYNOPSYS_UNCONNECTED__955, 
        SYNOPSYS_UNCONNECTED__956, SYNOPSYS_UNCONNECTED__957, 
        SYNOPSYS_UNCONNECTED__958, SYNOPSYS_UNCONNECTED__959, 
        SYNOPSYS_UNCONNECTED__960, N66863, N66862, N66861, N66860, N66859, 
        N66858}) );
  hamming_N16000_CC2_DW01_add_185 add_2851_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64431, N64430, N64429, N64428, 
        N64427}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64444, 
        N64443, N64442, N64441, N64440}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__961, SYNOPSYS_UNCONNECTED__962, 
        SYNOPSYS_UNCONNECTED__963, SYNOPSYS_UNCONNECTED__964, 
        SYNOPSYS_UNCONNECTED__965, SYNOPSYS_UNCONNECTED__966, 
        SYNOPSYS_UNCONNECTED__967, N66850, N66849, N66848, N66847, N66846, 
        N66845}) );
  hamming_N16000_CC2_DW01_add_186 add_2852_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64405, N64404, N64403, N64402, 
        N64401}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64418, 
        N64417, N64416, N64415, N64414}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__968, SYNOPSYS_UNCONNECTED__969, 
        SYNOPSYS_UNCONNECTED__970, SYNOPSYS_UNCONNECTED__971, 
        SYNOPSYS_UNCONNECTED__972, SYNOPSYS_UNCONNECTED__973, 
        SYNOPSYS_UNCONNECTED__974, N66837, N66836, N66835, N66834, N66833, 
        N66832}) );
  hamming_N16000_CC2_DW01_add_187 add_2853_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64379, N64378, N64377, N64376, 
        N64375}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64392, 
        N64391, N64390, N64389, N64388}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__975, SYNOPSYS_UNCONNECTED__976, 
        SYNOPSYS_UNCONNECTED__977, SYNOPSYS_UNCONNECTED__978, 
        SYNOPSYS_UNCONNECTED__979, SYNOPSYS_UNCONNECTED__980, 
        SYNOPSYS_UNCONNECTED__981, N66824, N66823, N66822, N66821, N66820, 
        N66819}) );
  hamming_N16000_CC2_DW01_add_188 add_2854_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64353, N64352, N64351, N64350, 
        N64349}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64366, 
        N64365, N64364, N64363, N64362}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__982, SYNOPSYS_UNCONNECTED__983, 
        SYNOPSYS_UNCONNECTED__984, SYNOPSYS_UNCONNECTED__985, 
        SYNOPSYS_UNCONNECTED__986, SYNOPSYS_UNCONNECTED__987, 
        SYNOPSYS_UNCONNECTED__988, N66811, N66810, N66809, N66808, N66807, 
        N66806}) );
  hamming_N16000_CC2_DW01_add_189 add_2855_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64327, N64326, N64325, N64324, 
        N64323}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64340, 
        N64339, N64338, N64337, N64336}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__989, SYNOPSYS_UNCONNECTED__990, 
        SYNOPSYS_UNCONNECTED__991, SYNOPSYS_UNCONNECTED__992, 
        SYNOPSYS_UNCONNECTED__993, SYNOPSYS_UNCONNECTED__994, 
        SYNOPSYS_UNCONNECTED__995, N66798, N66797, N66796, N66795, N66794, 
        N66793}) );
  hamming_N16000_CC2_DW01_add_190 add_2856_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64301, N64300, N64299, N64298, 
        N64297}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64314, 
        N64313, N64312, N64311, N64310}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__996, SYNOPSYS_UNCONNECTED__997, 
        SYNOPSYS_UNCONNECTED__998, SYNOPSYS_UNCONNECTED__999, 
        SYNOPSYS_UNCONNECTED__1000, SYNOPSYS_UNCONNECTED__1001, 
        SYNOPSYS_UNCONNECTED__1002, N66785, N66784, N66783, N66782, N66781, 
        N66780}) );
  hamming_N16000_CC2_DW01_add_191 add_2857_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64275, N64274, N64273, N64272, 
        N64271}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64288, 
        N64287, N64286, N64285, N64284}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1003, SYNOPSYS_UNCONNECTED__1004, 
        SYNOPSYS_UNCONNECTED__1005, SYNOPSYS_UNCONNECTED__1006, 
        SYNOPSYS_UNCONNECTED__1007, SYNOPSYS_UNCONNECTED__1008, 
        SYNOPSYS_UNCONNECTED__1009, N66772, N66771, N66770, N66769, N66768, 
        N66767}) );
  hamming_N16000_CC2_DW01_add_192 add_2858_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64249, N64248, N64247, N64246, 
        N64245}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64262, 
        N64261, N64260, N64259, N64258}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1010, SYNOPSYS_UNCONNECTED__1011, 
        SYNOPSYS_UNCONNECTED__1012, SYNOPSYS_UNCONNECTED__1013, 
        SYNOPSYS_UNCONNECTED__1014, SYNOPSYS_UNCONNECTED__1015, 
        SYNOPSYS_UNCONNECTED__1016, N66759, N66758, N66757, N66756, N66755, 
        N66754}) );
  hamming_N16000_CC2_DW01_add_193 add_2859_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64223, N64222, N64221, N64220, 
        N64219}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64236, 
        N64235, N64234, N64233, N64232}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1017, SYNOPSYS_UNCONNECTED__1018, 
        SYNOPSYS_UNCONNECTED__1019, SYNOPSYS_UNCONNECTED__1020, 
        SYNOPSYS_UNCONNECTED__1021, SYNOPSYS_UNCONNECTED__1022, 
        SYNOPSYS_UNCONNECTED__1023, N66746, N66745, N66744, N66743, N66742, 
        N66741}) );
  hamming_N16000_CC2_DW01_add_194 add_2860_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64197, N64196, N64195, N64194, 
        N64193}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64210, 
        N64209, N64208, N64207, N64206}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1024, SYNOPSYS_UNCONNECTED__1025, 
        SYNOPSYS_UNCONNECTED__1026, SYNOPSYS_UNCONNECTED__1027, 
        SYNOPSYS_UNCONNECTED__1028, SYNOPSYS_UNCONNECTED__1029, 
        SYNOPSYS_UNCONNECTED__1030, N66733, N66732, N66731, N66730, N66729, 
        N66728}) );
  hamming_N16000_CC2_DW01_add_195 add_2861_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64171, N64170, N64169, N64168, 
        N64167}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64184, 
        N64183, N64182, N64181, N64180}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1031, SYNOPSYS_UNCONNECTED__1032, 
        SYNOPSYS_UNCONNECTED__1033, SYNOPSYS_UNCONNECTED__1034, 
        SYNOPSYS_UNCONNECTED__1035, SYNOPSYS_UNCONNECTED__1036, 
        SYNOPSYS_UNCONNECTED__1037, N66720, N66719, N66718, N66717, N66716, 
        N66715}) );
  hamming_N16000_CC2_DW01_add_196 add_2862_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64145, N64144, N64143, N64142, 
        N64141}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64158, 
        N64157, N64156, N64155, N64154}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1038, SYNOPSYS_UNCONNECTED__1039, 
        SYNOPSYS_UNCONNECTED__1040, SYNOPSYS_UNCONNECTED__1041, 
        SYNOPSYS_UNCONNECTED__1042, SYNOPSYS_UNCONNECTED__1043, 
        SYNOPSYS_UNCONNECTED__1044, N66707, N66706, N66705, N66704, N66703, 
        N66702}) );
  hamming_N16000_CC2_DW01_add_197 add_2863_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64119, N64118, N64117, N64116, 
        N64115}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64132, 
        N64131, N64130, N64129, N64128}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1045, SYNOPSYS_UNCONNECTED__1046, 
        SYNOPSYS_UNCONNECTED__1047, SYNOPSYS_UNCONNECTED__1048, 
        SYNOPSYS_UNCONNECTED__1049, SYNOPSYS_UNCONNECTED__1050, 
        SYNOPSYS_UNCONNECTED__1051, N66694, N66693, N66692, N66691, N66690, 
        N66689}) );
  hamming_N16000_CC2_DW01_add_198 add_2864_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64093, N64092, N64091, N64090, 
        N64089}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64106, 
        N64105, N64104, N64103, N64102}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1052, SYNOPSYS_UNCONNECTED__1053, 
        SYNOPSYS_UNCONNECTED__1054, SYNOPSYS_UNCONNECTED__1055, 
        SYNOPSYS_UNCONNECTED__1056, SYNOPSYS_UNCONNECTED__1057, 
        SYNOPSYS_UNCONNECTED__1058, N66681, N66680, N66679, N66678, N66677, 
        N66676}) );
  hamming_N16000_CC2_DW01_add_199 add_2865_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64067, N64066, N64065, N64064, 
        N64063}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64080, 
        N64079, N64078, N64077, N64076}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1059, SYNOPSYS_UNCONNECTED__1060, 
        SYNOPSYS_UNCONNECTED__1061, SYNOPSYS_UNCONNECTED__1062, 
        SYNOPSYS_UNCONNECTED__1063, SYNOPSYS_UNCONNECTED__1064, 
        SYNOPSYS_UNCONNECTED__1065, N66668, N66667, N66666, N66665, N66664, 
        N66663}) );
  hamming_N16000_CC2_DW01_add_200 add_2866_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64041, N64040, N64039, N64038, 
        N64037}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64054, 
        N64053, N64052, N64051, N64050}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1066, SYNOPSYS_UNCONNECTED__1067, 
        SYNOPSYS_UNCONNECTED__1068, SYNOPSYS_UNCONNECTED__1069, 
        SYNOPSYS_UNCONNECTED__1070, SYNOPSYS_UNCONNECTED__1071, 
        SYNOPSYS_UNCONNECTED__1072, N66655, N66654, N66653, N66652, N66651, 
        N66650}) );
  hamming_N16000_CC2_DW01_add_201 add_2867_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64015, N64014, N64013, N64012, 
        N64011}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64028, 
        N64027, N64026, N64025, N64024}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1073, SYNOPSYS_UNCONNECTED__1074, 
        SYNOPSYS_UNCONNECTED__1075, SYNOPSYS_UNCONNECTED__1076, 
        SYNOPSYS_UNCONNECTED__1077, SYNOPSYS_UNCONNECTED__1078, 
        SYNOPSYS_UNCONNECTED__1079, N66642, N66641, N66640, N66639, N66638, 
        N66637}) );
  hamming_N16000_CC2_DW01_add_202 add_2868_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63989, N63988, N63987, N63986, 
        N63985}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N64002, 
        N64001, N64000, N63999, N63998}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1080, SYNOPSYS_UNCONNECTED__1081, 
        SYNOPSYS_UNCONNECTED__1082, SYNOPSYS_UNCONNECTED__1083, 
        SYNOPSYS_UNCONNECTED__1084, SYNOPSYS_UNCONNECTED__1085, 
        SYNOPSYS_UNCONNECTED__1086, N66629, N66628, N66627, N66626, N66625, 
        N66624}) );
  hamming_N16000_CC2_DW01_add_203 add_2869_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63963, N63962, N63961, N63960, 
        N63959}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63976, 
        N63975, N63974, N63973, N63972}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1087, SYNOPSYS_UNCONNECTED__1088, 
        SYNOPSYS_UNCONNECTED__1089, SYNOPSYS_UNCONNECTED__1090, 
        SYNOPSYS_UNCONNECTED__1091, SYNOPSYS_UNCONNECTED__1092, 
        SYNOPSYS_UNCONNECTED__1093, N66616, N66615, N66614, N66613, N66612, 
        N66611}) );
  hamming_N16000_CC2_DW01_add_204 add_2870_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63937, N63936, N63935, N63934, 
        N63933}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63950, 
        N63949, N63948, N63947, N63946}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1094, SYNOPSYS_UNCONNECTED__1095, 
        SYNOPSYS_UNCONNECTED__1096, SYNOPSYS_UNCONNECTED__1097, 
        SYNOPSYS_UNCONNECTED__1098, SYNOPSYS_UNCONNECTED__1099, 
        SYNOPSYS_UNCONNECTED__1100, N66603, N66602, N66601, N66600, N66599, 
        N66598}) );
  hamming_N16000_CC2_DW01_add_205 add_2871_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63911, N63910, N63909, N63908, 
        N63907}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63924, 
        N63923, N63922, N63921, N63920}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1101, SYNOPSYS_UNCONNECTED__1102, 
        SYNOPSYS_UNCONNECTED__1103, SYNOPSYS_UNCONNECTED__1104, 
        SYNOPSYS_UNCONNECTED__1105, SYNOPSYS_UNCONNECTED__1106, 
        SYNOPSYS_UNCONNECTED__1107, N66590, N66589, N66588, N66587, N66586, 
        N66585}) );
  hamming_N16000_CC2_DW01_add_206 add_2872_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63885, N63884, N63883, N63882, 
        N63881}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63898, 
        N63897, N63896, N63895, N63894}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1108, SYNOPSYS_UNCONNECTED__1109, 
        SYNOPSYS_UNCONNECTED__1110, SYNOPSYS_UNCONNECTED__1111, 
        SYNOPSYS_UNCONNECTED__1112, SYNOPSYS_UNCONNECTED__1113, 
        SYNOPSYS_UNCONNECTED__1114, N66577, N66576, N66575, N66574, N66573, 
        N66572}) );
  hamming_N16000_CC2_DW01_add_207 add_2873_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63859, N63858, N63857, N63856, 
        N63855}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63872, 
        N63871, N63870, N63869, N63868}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1115, SYNOPSYS_UNCONNECTED__1116, 
        SYNOPSYS_UNCONNECTED__1117, SYNOPSYS_UNCONNECTED__1118, 
        SYNOPSYS_UNCONNECTED__1119, SYNOPSYS_UNCONNECTED__1120, 
        SYNOPSYS_UNCONNECTED__1121, N66564, N66563, N66562, N66561, N66560, 
        N66559}) );
  hamming_N16000_CC2_DW01_add_208 add_2874_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63833, N63832, N63831, N63830, 
        N63829}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63846, 
        N63845, N63844, N63843, N63842}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1122, SYNOPSYS_UNCONNECTED__1123, 
        SYNOPSYS_UNCONNECTED__1124, SYNOPSYS_UNCONNECTED__1125, 
        SYNOPSYS_UNCONNECTED__1126, SYNOPSYS_UNCONNECTED__1127, 
        SYNOPSYS_UNCONNECTED__1128, N66551, N66550, N66549, N66548, N66547, 
        N66546}) );
  hamming_N16000_CC2_DW01_add_209 add_2875_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63807, N63806, N63805, N63804, 
        N63803}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63820, 
        N63819, N63818, N63817, N63816}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1129, SYNOPSYS_UNCONNECTED__1130, 
        SYNOPSYS_UNCONNECTED__1131, SYNOPSYS_UNCONNECTED__1132, 
        SYNOPSYS_UNCONNECTED__1133, SYNOPSYS_UNCONNECTED__1134, 
        SYNOPSYS_UNCONNECTED__1135, N66538, N66537, N66536, N66535, N66534, 
        N66533}) );
  hamming_N16000_CC2_DW01_add_210 add_2876_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63781, N63780, N63779, N63778, 
        N63777}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63794, 
        N63793, N63792, N63791, N63790}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1136, SYNOPSYS_UNCONNECTED__1137, 
        SYNOPSYS_UNCONNECTED__1138, SYNOPSYS_UNCONNECTED__1139, 
        SYNOPSYS_UNCONNECTED__1140, SYNOPSYS_UNCONNECTED__1141, 
        SYNOPSYS_UNCONNECTED__1142, N66525, N66524, N66523, N66522, N66521, 
        N66520}) );
  hamming_N16000_CC2_DW01_add_211 add_2877_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63755, N63754, N63753, N63752, 
        N63751}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63768, 
        N63767, N63766, N63765, N63764}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1143, SYNOPSYS_UNCONNECTED__1144, 
        SYNOPSYS_UNCONNECTED__1145, SYNOPSYS_UNCONNECTED__1146, 
        SYNOPSYS_UNCONNECTED__1147, SYNOPSYS_UNCONNECTED__1148, 
        SYNOPSYS_UNCONNECTED__1149, N66512, N66511, N66510, N66509, N66508, 
        N66507}) );
  hamming_N16000_CC2_DW01_add_212 add_2878_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63729, N63728, N63727, N63726, 
        N63725}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63742, 
        N63741, N63740, N63739, N63738}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1150, SYNOPSYS_UNCONNECTED__1151, 
        SYNOPSYS_UNCONNECTED__1152, SYNOPSYS_UNCONNECTED__1153, 
        SYNOPSYS_UNCONNECTED__1154, SYNOPSYS_UNCONNECTED__1155, 
        SYNOPSYS_UNCONNECTED__1156, N66499, N66498, N66497, N66496, N66495, 
        N66494}) );
  hamming_N16000_CC2_DW01_add_213 add_2879_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63703, N63702, N63701, N63700, 
        N63699}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63716, 
        N63715, N63714, N63713, N63712}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1157, SYNOPSYS_UNCONNECTED__1158, 
        SYNOPSYS_UNCONNECTED__1159, SYNOPSYS_UNCONNECTED__1160, 
        SYNOPSYS_UNCONNECTED__1161, SYNOPSYS_UNCONNECTED__1162, 
        SYNOPSYS_UNCONNECTED__1163, N66486, N66485, N66484, N66483, N66482, 
        N66481}) );
  hamming_N16000_CC2_DW01_add_214 add_2880_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63677, N63676, N63675, N63674, 
        N63673}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63690, 
        N63689, N63688, N63687, N63686}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1164, SYNOPSYS_UNCONNECTED__1165, 
        SYNOPSYS_UNCONNECTED__1166, SYNOPSYS_UNCONNECTED__1167, 
        SYNOPSYS_UNCONNECTED__1168, SYNOPSYS_UNCONNECTED__1169, 
        SYNOPSYS_UNCONNECTED__1170, N66473, N66472, N66471, N66470, N66469, 
        N66468}) );
  hamming_N16000_CC2_DW01_add_215 add_2881_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63651, N63650, N63649, N63648, 
        N63647}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63664, 
        N63663, N63662, N63661, N63660}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1171, SYNOPSYS_UNCONNECTED__1172, 
        SYNOPSYS_UNCONNECTED__1173, SYNOPSYS_UNCONNECTED__1174, 
        SYNOPSYS_UNCONNECTED__1175, SYNOPSYS_UNCONNECTED__1176, 
        SYNOPSYS_UNCONNECTED__1177, N66460, N66459, N66458, N66457, N66456, 
        N66455}) );
  hamming_N16000_CC2_DW01_add_216 add_2882_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63625, N63624, N63623, N63622, 
        N63621}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63638, 
        N63637, N63636, N63635, N63634}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1178, SYNOPSYS_UNCONNECTED__1179, 
        SYNOPSYS_UNCONNECTED__1180, SYNOPSYS_UNCONNECTED__1181, 
        SYNOPSYS_UNCONNECTED__1182, SYNOPSYS_UNCONNECTED__1183, 
        SYNOPSYS_UNCONNECTED__1184, N66447, N66446, N66445, N66444, N66443, 
        N66442}) );
  hamming_N16000_CC2_DW01_add_217 add_2883_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63599, N63598, N63597, N63596, 
        N63595}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63612, 
        N63611, N63610, N63609, N63608}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1185, SYNOPSYS_UNCONNECTED__1186, 
        SYNOPSYS_UNCONNECTED__1187, SYNOPSYS_UNCONNECTED__1188, 
        SYNOPSYS_UNCONNECTED__1189, SYNOPSYS_UNCONNECTED__1190, 
        SYNOPSYS_UNCONNECTED__1191, N66434, N66433, N66432, N66431, N66430, 
        N66429}) );
  hamming_N16000_CC2_DW01_add_218 add_2884_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63573, N63572, N63571, N63570, 
        N63569}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63586, 
        N63585, N63584, N63583, N63582}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1192, SYNOPSYS_UNCONNECTED__1193, 
        SYNOPSYS_UNCONNECTED__1194, SYNOPSYS_UNCONNECTED__1195, 
        SYNOPSYS_UNCONNECTED__1196, SYNOPSYS_UNCONNECTED__1197, 
        SYNOPSYS_UNCONNECTED__1198, N66421, N66420, N66419, N66418, N66417, 
        N66416}) );
  hamming_N16000_CC2_DW01_add_219 add_2885_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63547, N63546, N63545, N63544, 
        N63543}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63560, 
        N63559, N63558, N63557, N63556}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1199, SYNOPSYS_UNCONNECTED__1200, 
        SYNOPSYS_UNCONNECTED__1201, SYNOPSYS_UNCONNECTED__1202, 
        SYNOPSYS_UNCONNECTED__1203, SYNOPSYS_UNCONNECTED__1204, 
        SYNOPSYS_UNCONNECTED__1205, N66408, N66407, N66406, N66405, N66404, 
        N66403}) );
  hamming_N16000_CC2_DW01_add_220 add_2886_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63521, N63520, N63519, N63518, 
        N63517}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63534, 
        N63533, N63532, N63531, N63530}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1206, SYNOPSYS_UNCONNECTED__1207, 
        SYNOPSYS_UNCONNECTED__1208, SYNOPSYS_UNCONNECTED__1209, 
        SYNOPSYS_UNCONNECTED__1210, SYNOPSYS_UNCONNECTED__1211, 
        SYNOPSYS_UNCONNECTED__1212, N66395, N66394, N66393, N66392, N66391, 
        N66390}) );
  hamming_N16000_CC2_DW01_add_221 add_2887_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63495, N63494, N63493, N63492, 
        N63491}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63508, 
        N63507, N63506, N63505, N63504}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1213, SYNOPSYS_UNCONNECTED__1214, 
        SYNOPSYS_UNCONNECTED__1215, SYNOPSYS_UNCONNECTED__1216, 
        SYNOPSYS_UNCONNECTED__1217, SYNOPSYS_UNCONNECTED__1218, 
        SYNOPSYS_UNCONNECTED__1219, N66382, N66381, N66380, N66379, N66378, 
        N66377}) );
  hamming_N16000_CC2_DW01_add_222 add_2888_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63469, N63468, N63467, N63466, 
        N63465}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63482, 
        N63481, N63480, N63479, N63478}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1220, SYNOPSYS_UNCONNECTED__1221, 
        SYNOPSYS_UNCONNECTED__1222, SYNOPSYS_UNCONNECTED__1223, 
        SYNOPSYS_UNCONNECTED__1224, SYNOPSYS_UNCONNECTED__1225, 
        SYNOPSYS_UNCONNECTED__1226, N66369, N66368, N66367, N66366, N66365, 
        N66364}) );
  hamming_N16000_CC2_DW01_add_223 add_2889_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63443, N63442, N63441, N63440, 
        N63439}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63456, 
        N63455, N63454, N63453, N63452}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1227, SYNOPSYS_UNCONNECTED__1228, 
        SYNOPSYS_UNCONNECTED__1229, SYNOPSYS_UNCONNECTED__1230, 
        SYNOPSYS_UNCONNECTED__1231, SYNOPSYS_UNCONNECTED__1232, 
        SYNOPSYS_UNCONNECTED__1233, N66356, N66355, N66354, N66353, N66352, 
        N66351}) );
  hamming_N16000_CC2_DW01_add_224 add_2890_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63417, N63416, N63415, N63414, 
        N63413}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63430, 
        N63429, N63428, N63427, N63426}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1234, SYNOPSYS_UNCONNECTED__1235, 
        SYNOPSYS_UNCONNECTED__1236, SYNOPSYS_UNCONNECTED__1237, 
        SYNOPSYS_UNCONNECTED__1238, SYNOPSYS_UNCONNECTED__1239, 
        SYNOPSYS_UNCONNECTED__1240, N66343, N66342, N66341, N66340, N66339, 
        N66338}) );
  hamming_N16000_CC2_DW01_add_225 add_2891_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63391, N63390, N63389, N63388, 
        N63387}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63404, 
        N63403, N63402, N63401, N63400}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1241, SYNOPSYS_UNCONNECTED__1242, 
        SYNOPSYS_UNCONNECTED__1243, SYNOPSYS_UNCONNECTED__1244, 
        SYNOPSYS_UNCONNECTED__1245, SYNOPSYS_UNCONNECTED__1246, 
        SYNOPSYS_UNCONNECTED__1247, N66330, N66329, N66328, N66327, N66326, 
        N66325}) );
  hamming_N16000_CC2_DW01_add_226 add_2892_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63365, N63364, N63363, N63362, 
        N63361}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63378, 
        N63377, N63376, N63375, N63374}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1248, SYNOPSYS_UNCONNECTED__1249, 
        SYNOPSYS_UNCONNECTED__1250, SYNOPSYS_UNCONNECTED__1251, 
        SYNOPSYS_UNCONNECTED__1252, SYNOPSYS_UNCONNECTED__1253, 
        SYNOPSYS_UNCONNECTED__1254, N66317, N66316, N66315, N66314, N66313, 
        N66312}) );
  hamming_N16000_CC2_DW01_add_227 add_2893_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63339, N63338, N63337, N63336, 
        N63335}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63352, 
        N63351, N63350, N63349, N63348}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1255, SYNOPSYS_UNCONNECTED__1256, 
        SYNOPSYS_UNCONNECTED__1257, SYNOPSYS_UNCONNECTED__1258, 
        SYNOPSYS_UNCONNECTED__1259, SYNOPSYS_UNCONNECTED__1260, 
        SYNOPSYS_UNCONNECTED__1261, N66304, N66303, N66302, N66301, N66300, 
        N66299}) );
  hamming_N16000_CC2_DW01_add_228 add_2894_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63313, N63312, N63311, N63310, 
        N63309}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63326, 
        N63325, N63324, N63323, N63322}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1262, SYNOPSYS_UNCONNECTED__1263, 
        SYNOPSYS_UNCONNECTED__1264, SYNOPSYS_UNCONNECTED__1265, 
        SYNOPSYS_UNCONNECTED__1266, SYNOPSYS_UNCONNECTED__1267, 
        SYNOPSYS_UNCONNECTED__1268, N66291, N66290, N66289, N66288, N66287, 
        N66286}) );
  hamming_N16000_CC2_DW01_add_229 add_2895_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63287, N63286, N63285, N63284, 
        N63283}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63300, 
        N63299, N63298, N63297, N63296}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1269, SYNOPSYS_UNCONNECTED__1270, 
        SYNOPSYS_UNCONNECTED__1271, SYNOPSYS_UNCONNECTED__1272, 
        SYNOPSYS_UNCONNECTED__1273, SYNOPSYS_UNCONNECTED__1274, 
        SYNOPSYS_UNCONNECTED__1275, N66278, N66277, N66276, N66275, N66274, 
        N66273}) );
  hamming_N16000_CC2_DW01_add_230 add_2896_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63261, N63260, N63259, N63258, 
        N63257}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63274, 
        N63273, N63272, N63271, N63270}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1276, SYNOPSYS_UNCONNECTED__1277, 
        SYNOPSYS_UNCONNECTED__1278, SYNOPSYS_UNCONNECTED__1279, 
        SYNOPSYS_UNCONNECTED__1280, SYNOPSYS_UNCONNECTED__1281, 
        SYNOPSYS_UNCONNECTED__1282, N66265, N66264, N66263, N66262, N66261, 
        N66260}) );
  hamming_N16000_CC2_DW01_add_231 add_2897_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63235, N63234, N63233, N63232, 
        N63231}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63248, 
        N63247, N63246, N63245, N63244}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1283, SYNOPSYS_UNCONNECTED__1284, 
        SYNOPSYS_UNCONNECTED__1285, SYNOPSYS_UNCONNECTED__1286, 
        SYNOPSYS_UNCONNECTED__1287, SYNOPSYS_UNCONNECTED__1288, 
        SYNOPSYS_UNCONNECTED__1289, N66252, N66251, N66250, N66249, N66248, 
        N66247}) );
  hamming_N16000_CC2_DW01_add_232 add_2898_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63209, N63208, N63207, N63206, 
        N63205}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63222, 
        N63221, N63220, N63219, N63218}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1290, SYNOPSYS_UNCONNECTED__1291, 
        SYNOPSYS_UNCONNECTED__1292, SYNOPSYS_UNCONNECTED__1293, 
        SYNOPSYS_UNCONNECTED__1294, SYNOPSYS_UNCONNECTED__1295, 
        SYNOPSYS_UNCONNECTED__1296, N66239, N66238, N66237, N66236, N66235, 
        N66234}) );
  hamming_N16000_CC2_DW01_add_233 add_2899_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63183, N63182, N63181, N63180, 
        N63179}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63196, 
        N63195, N63194, N63193, N63192}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1297, SYNOPSYS_UNCONNECTED__1298, 
        SYNOPSYS_UNCONNECTED__1299, SYNOPSYS_UNCONNECTED__1300, 
        SYNOPSYS_UNCONNECTED__1301, SYNOPSYS_UNCONNECTED__1302, 
        SYNOPSYS_UNCONNECTED__1303, N66226, N66225, N66224, N66223, N66222, 
        N66221}) );
  hamming_N16000_CC2_DW01_add_234 add_2900_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63157, N63156, N63155, N63154, 
        N63153}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63170, 
        N63169, N63168, N63167, N63166}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1304, SYNOPSYS_UNCONNECTED__1305, 
        SYNOPSYS_UNCONNECTED__1306, SYNOPSYS_UNCONNECTED__1307, 
        SYNOPSYS_UNCONNECTED__1308, SYNOPSYS_UNCONNECTED__1309, 
        SYNOPSYS_UNCONNECTED__1310, N66213, N66212, N66211, N66210, N66209, 
        N66208}) );
  hamming_N16000_CC2_DW01_add_235 add_2901_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63131, N63130, N63129, N63128, 
        N63127}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63144, 
        N63143, N63142, N63141, N63140}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1311, SYNOPSYS_UNCONNECTED__1312, 
        SYNOPSYS_UNCONNECTED__1313, SYNOPSYS_UNCONNECTED__1314, 
        SYNOPSYS_UNCONNECTED__1315, SYNOPSYS_UNCONNECTED__1316, 
        SYNOPSYS_UNCONNECTED__1317, N66200, N66199, N66198, N66197, N66196, 
        N66195}) );
  hamming_N16000_CC2_DW01_add_236 add_2902_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63105, N63104, N63103, N63102, 
        N63101}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63118, 
        N63117, N63116, N63115, N63114}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1318, SYNOPSYS_UNCONNECTED__1319, 
        SYNOPSYS_UNCONNECTED__1320, SYNOPSYS_UNCONNECTED__1321, 
        SYNOPSYS_UNCONNECTED__1322, SYNOPSYS_UNCONNECTED__1323, 
        SYNOPSYS_UNCONNECTED__1324, N66187, N66186, N66185, N66184, N66183, 
        N66182}) );
  hamming_N16000_CC2_DW01_add_237 add_2903_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63079, N63078, N63077, N63076, 
        N63075}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63092, 
        N63091, N63090, N63089, N63088}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1325, SYNOPSYS_UNCONNECTED__1326, 
        SYNOPSYS_UNCONNECTED__1327, SYNOPSYS_UNCONNECTED__1328, 
        SYNOPSYS_UNCONNECTED__1329, SYNOPSYS_UNCONNECTED__1330, 
        SYNOPSYS_UNCONNECTED__1331, N66174, N66173, N66172, N66171, N66170, 
        N66169}) );
  hamming_N16000_CC2_DW01_add_238 add_2904_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63053, N63052, N63051, N63050, 
        N63049}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63066, 
        N63065, N63064, N63063, N63062}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1332, SYNOPSYS_UNCONNECTED__1333, 
        SYNOPSYS_UNCONNECTED__1334, SYNOPSYS_UNCONNECTED__1335, 
        SYNOPSYS_UNCONNECTED__1336, SYNOPSYS_UNCONNECTED__1337, 
        SYNOPSYS_UNCONNECTED__1338, N66161, N66160, N66159, N66158, N66157, 
        N66156}) );
  hamming_N16000_CC2_DW01_add_239 add_2905_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63027, N63026, N63025, N63024, 
        N63023}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63040, 
        N63039, N63038, N63037, N63036}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1339, SYNOPSYS_UNCONNECTED__1340, 
        SYNOPSYS_UNCONNECTED__1341, SYNOPSYS_UNCONNECTED__1342, 
        SYNOPSYS_UNCONNECTED__1343, SYNOPSYS_UNCONNECTED__1344, 
        SYNOPSYS_UNCONNECTED__1345, N66148, N66147, N66146, N66145, N66144, 
        N66143}) );
  hamming_N16000_CC2_DW01_add_240 add_2906_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63001, N63000, N62999, N62998, 
        N62997}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N63014, 
        N63013, N63012, N63011, N63010}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1346, SYNOPSYS_UNCONNECTED__1347, 
        SYNOPSYS_UNCONNECTED__1348, SYNOPSYS_UNCONNECTED__1349, 
        SYNOPSYS_UNCONNECTED__1350, SYNOPSYS_UNCONNECTED__1351, 
        SYNOPSYS_UNCONNECTED__1352, N66135, N66134, N66133, N66132, N66131, 
        N66130}) );
  hamming_N16000_CC2_DW01_add_241 add_2907_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62975, N62974, N62973, N62972, 
        N62971}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62988, 
        N62987, N62986, N62985, N62984}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1353, SYNOPSYS_UNCONNECTED__1354, 
        SYNOPSYS_UNCONNECTED__1355, SYNOPSYS_UNCONNECTED__1356, 
        SYNOPSYS_UNCONNECTED__1357, SYNOPSYS_UNCONNECTED__1358, 
        SYNOPSYS_UNCONNECTED__1359, N66122, N66121, N66120, N66119, N66118, 
        N66117}) );
  hamming_N16000_CC2_DW01_add_242 add_2908_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62949, N62948, N62947, N62946, 
        N62945}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62962, 
        N62961, N62960, N62959, N62958}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1360, SYNOPSYS_UNCONNECTED__1361, 
        SYNOPSYS_UNCONNECTED__1362, SYNOPSYS_UNCONNECTED__1363, 
        SYNOPSYS_UNCONNECTED__1364, SYNOPSYS_UNCONNECTED__1365, 
        SYNOPSYS_UNCONNECTED__1366, N66109, N66108, N66107, N66106, N66105, 
        N66104}) );
  hamming_N16000_CC2_DW01_add_243 add_2909_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62923, N62922, N62921, N62920, 
        N62919}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62936, 
        N62935, N62934, N62933, N62932}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1367, SYNOPSYS_UNCONNECTED__1368, 
        SYNOPSYS_UNCONNECTED__1369, SYNOPSYS_UNCONNECTED__1370, 
        SYNOPSYS_UNCONNECTED__1371, SYNOPSYS_UNCONNECTED__1372, 
        SYNOPSYS_UNCONNECTED__1373, N66096, N66095, N66094, N66093, N66092, 
        N66091}) );
  hamming_N16000_CC2_DW01_add_244 add_2910_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62897, N62896, N62895, N62894, 
        N62893}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62910, 
        N62909, N62908, N62907, N62906}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1374, SYNOPSYS_UNCONNECTED__1375, 
        SYNOPSYS_UNCONNECTED__1376, SYNOPSYS_UNCONNECTED__1377, 
        SYNOPSYS_UNCONNECTED__1378, SYNOPSYS_UNCONNECTED__1379, 
        SYNOPSYS_UNCONNECTED__1380, N66083, N66082, N66081, N66080, N66079, 
        N66078}) );
  hamming_N16000_CC2_DW01_add_245 add_2911_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62871, N62870, N62869, N62868, 
        N62867}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62884, 
        N62883, N62882, N62881, N62880}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1381, SYNOPSYS_UNCONNECTED__1382, 
        SYNOPSYS_UNCONNECTED__1383, SYNOPSYS_UNCONNECTED__1384, 
        SYNOPSYS_UNCONNECTED__1385, SYNOPSYS_UNCONNECTED__1386, 
        SYNOPSYS_UNCONNECTED__1387, N66070, N66069, N66068, N66067, N66066, 
        N66065}) );
  hamming_N16000_CC2_DW01_add_246 add_2912_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62845, N62844, N62843, N62842, 
        N62841}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62858, 
        N62857, N62856, N62855, N62854}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1388, SYNOPSYS_UNCONNECTED__1389, 
        SYNOPSYS_UNCONNECTED__1390, SYNOPSYS_UNCONNECTED__1391, 
        SYNOPSYS_UNCONNECTED__1392, SYNOPSYS_UNCONNECTED__1393, 
        SYNOPSYS_UNCONNECTED__1394, N66057, N66056, N66055, N66054, N66053, 
        N66052}) );
  hamming_N16000_CC2_DW01_add_247 add_2913_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62819, N62818, N62817, N62816, 
        N62815}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62832, 
        N62831, N62830, N62829, N62828}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1395, SYNOPSYS_UNCONNECTED__1396, 
        SYNOPSYS_UNCONNECTED__1397, SYNOPSYS_UNCONNECTED__1398, 
        SYNOPSYS_UNCONNECTED__1399, SYNOPSYS_UNCONNECTED__1400, 
        SYNOPSYS_UNCONNECTED__1401, N66044, N66043, N66042, N66041, N66040, 
        N66039}) );
  hamming_N16000_CC2_DW01_add_248 add_2914_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62793, N62792, N62791, N62790, 
        N62789}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62806, 
        N62805, N62804, N62803, N62802}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1402, SYNOPSYS_UNCONNECTED__1403, 
        SYNOPSYS_UNCONNECTED__1404, SYNOPSYS_UNCONNECTED__1405, 
        SYNOPSYS_UNCONNECTED__1406, SYNOPSYS_UNCONNECTED__1407, 
        SYNOPSYS_UNCONNECTED__1408, N66031, N66030, N66029, N66028, N66027, 
        N66026}) );
  hamming_N16000_CC2_DW01_add_249 add_2915_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62767, N62766, N62765, N62764, 
        N62763}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62780, 
        N62779, N62778, N62777, N62776}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1409, SYNOPSYS_UNCONNECTED__1410, 
        SYNOPSYS_UNCONNECTED__1411, SYNOPSYS_UNCONNECTED__1412, 
        SYNOPSYS_UNCONNECTED__1413, SYNOPSYS_UNCONNECTED__1414, 
        SYNOPSYS_UNCONNECTED__1415, N66018, N66017, N66016, N66015, N66014, 
        N66013}) );
  hamming_N16000_CC2_DW01_add_250 add_2916_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62741, N62740, N62739, N62738, 
        N62737}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62754, 
        N62753, N62752, N62751, N62750}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1416, SYNOPSYS_UNCONNECTED__1417, 
        SYNOPSYS_UNCONNECTED__1418, SYNOPSYS_UNCONNECTED__1419, 
        SYNOPSYS_UNCONNECTED__1420, SYNOPSYS_UNCONNECTED__1421, 
        SYNOPSYS_UNCONNECTED__1422, N66005, N66004, N66003, N66002, N66001, 
        N66000}) );
  hamming_N16000_CC2_DW01_add_251 add_2917_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62715, N62714, N62713, N62712, 
        N62711}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62728, 
        N62727, N62726, N62725, N62724}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1423, SYNOPSYS_UNCONNECTED__1424, 
        SYNOPSYS_UNCONNECTED__1425, SYNOPSYS_UNCONNECTED__1426, 
        SYNOPSYS_UNCONNECTED__1427, SYNOPSYS_UNCONNECTED__1428, 
        SYNOPSYS_UNCONNECTED__1429, N65992, N65991, N65990, N65989, N65988, 
        N65987}) );
  hamming_N16000_CC2_DW01_add_252 add_2918_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62689, N62688, N62687, N62686, 
        N62685}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62702, 
        N62701, N62700, N62699, N62698}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1430, SYNOPSYS_UNCONNECTED__1431, 
        SYNOPSYS_UNCONNECTED__1432, SYNOPSYS_UNCONNECTED__1433, 
        SYNOPSYS_UNCONNECTED__1434, SYNOPSYS_UNCONNECTED__1435, 
        SYNOPSYS_UNCONNECTED__1436, N65979, N65978, N65977, N65976, N65975, 
        N65974}) );
  hamming_N16000_CC2_DW01_add_253 add_2919_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62663, N62662, N62661, N62660, 
        N62659}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62676, 
        N62675, N62674, N62673, N62672}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1437, SYNOPSYS_UNCONNECTED__1438, 
        SYNOPSYS_UNCONNECTED__1439, SYNOPSYS_UNCONNECTED__1440, 
        SYNOPSYS_UNCONNECTED__1441, SYNOPSYS_UNCONNECTED__1442, 
        SYNOPSYS_UNCONNECTED__1443, N65966, N65965, N65964, N65963, N65962, 
        N65961}) );
  hamming_N16000_CC2_DW01_add_254 add_2920_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62637, N62636, N62635, N62634, 
        N62633}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62650, 
        N62649, N62648, N62647, N62646}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1444, SYNOPSYS_UNCONNECTED__1445, 
        SYNOPSYS_UNCONNECTED__1446, SYNOPSYS_UNCONNECTED__1447, 
        SYNOPSYS_UNCONNECTED__1448, SYNOPSYS_UNCONNECTED__1449, 
        SYNOPSYS_UNCONNECTED__1450, N65953, N65952, N65951, N65950, N65949, 
        N65948}) );
  hamming_N16000_CC2_DW01_add_255 add_2921_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62611, N62610, N62609, N62608, 
        N62607}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62624, 
        N62623, N62622, N62621, N62620}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1451, SYNOPSYS_UNCONNECTED__1452, 
        SYNOPSYS_UNCONNECTED__1453, SYNOPSYS_UNCONNECTED__1454, 
        SYNOPSYS_UNCONNECTED__1455, SYNOPSYS_UNCONNECTED__1456, 
        SYNOPSYS_UNCONNECTED__1457, N65940, N65939, N65938, N65937, N65936, 
        N65935}) );
  hamming_N16000_CC2_DW01_add_256 add_2922_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62585, N62584, N62583, N62582, 
        N62581}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62598, 
        N62597, N62596, N62595, N62594}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1458, SYNOPSYS_UNCONNECTED__1459, 
        SYNOPSYS_UNCONNECTED__1460, SYNOPSYS_UNCONNECTED__1461, 
        SYNOPSYS_UNCONNECTED__1462, SYNOPSYS_UNCONNECTED__1463, 
        SYNOPSYS_UNCONNECTED__1464, N65927, N65926, N65925, N65924, N65923, 
        N65922}) );
  hamming_N16000_CC2_DW01_add_257 add_2923_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62559, N62558, N62557, N62556, 
        N62555}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62572, 
        N62571, N62570, N62569, N62568}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1465, SYNOPSYS_UNCONNECTED__1466, 
        SYNOPSYS_UNCONNECTED__1467, SYNOPSYS_UNCONNECTED__1468, 
        SYNOPSYS_UNCONNECTED__1469, SYNOPSYS_UNCONNECTED__1470, 
        SYNOPSYS_UNCONNECTED__1471, N65914, N65913, N65912, N65911, N65910, 
        N65909}) );
  hamming_N16000_CC2_DW01_add_258 add_2924_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62533, N62532, N62531, N62530, 
        N62529}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62546, 
        N62545, N62544, N62543, N62542}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1472, SYNOPSYS_UNCONNECTED__1473, 
        SYNOPSYS_UNCONNECTED__1474, SYNOPSYS_UNCONNECTED__1475, 
        SYNOPSYS_UNCONNECTED__1476, SYNOPSYS_UNCONNECTED__1477, 
        SYNOPSYS_UNCONNECTED__1478, N65901, N65900, N65899, N65898, N65897, 
        N65896}) );
  hamming_N16000_CC2_DW01_add_259 add_2925_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62507, N62506, N62505, N62504, 
        N62503}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62520, 
        N62519, N62518, N62517, N62516}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1479, SYNOPSYS_UNCONNECTED__1480, 
        SYNOPSYS_UNCONNECTED__1481, SYNOPSYS_UNCONNECTED__1482, 
        SYNOPSYS_UNCONNECTED__1483, SYNOPSYS_UNCONNECTED__1484, 
        SYNOPSYS_UNCONNECTED__1485, N65888, N65887, N65886, N65885, N65884, 
        N65883}) );
  hamming_N16000_CC2_DW01_add_260 add_2926_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62481, N62480, N62479, N62478, 
        N62477}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62494, 
        N62493, N62492, N62491, N62490}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1486, SYNOPSYS_UNCONNECTED__1487, 
        SYNOPSYS_UNCONNECTED__1488, SYNOPSYS_UNCONNECTED__1489, 
        SYNOPSYS_UNCONNECTED__1490, SYNOPSYS_UNCONNECTED__1491, 
        SYNOPSYS_UNCONNECTED__1492, N65875, N65874, N65873, N65872, N65871, 
        N65870}) );
  hamming_N16000_CC2_DW01_add_261 add_2927_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62455, N62454, N62453, N62452, 
        N62451}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62468, 
        N62467, N62466, N62465, N62464}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1493, SYNOPSYS_UNCONNECTED__1494, 
        SYNOPSYS_UNCONNECTED__1495, SYNOPSYS_UNCONNECTED__1496, 
        SYNOPSYS_UNCONNECTED__1497, SYNOPSYS_UNCONNECTED__1498, 
        SYNOPSYS_UNCONNECTED__1499, N65862, N65861, N65860, N65859, N65858, 
        N65857}) );
  hamming_N16000_CC2_DW01_add_262 add_2928_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62429, N62428, N62427, N62426, 
        N62425}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62442, 
        N62441, N62440, N62439, N62438}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1500, SYNOPSYS_UNCONNECTED__1501, 
        SYNOPSYS_UNCONNECTED__1502, SYNOPSYS_UNCONNECTED__1503, 
        SYNOPSYS_UNCONNECTED__1504, SYNOPSYS_UNCONNECTED__1505, 
        SYNOPSYS_UNCONNECTED__1506, N65849, N65848, N65847, N65846, N65845, 
        N65844}) );
  hamming_N16000_CC2_DW01_add_263 add_2929_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62403, N62402, N62401, N62400, 
        N62399}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62416, 
        N62415, N62414, N62413, N62412}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1507, SYNOPSYS_UNCONNECTED__1508, 
        SYNOPSYS_UNCONNECTED__1509, SYNOPSYS_UNCONNECTED__1510, 
        SYNOPSYS_UNCONNECTED__1511, SYNOPSYS_UNCONNECTED__1512, 
        SYNOPSYS_UNCONNECTED__1513, N65836, N65835, N65834, N65833, N65832, 
        N65831}) );
  hamming_N16000_CC2_DW01_add_264 add_2930_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62377, N62376, N62375, N62374, 
        N62373}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62390, 
        N62389, N62388, N62387, N62386}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1514, SYNOPSYS_UNCONNECTED__1515, 
        SYNOPSYS_UNCONNECTED__1516, SYNOPSYS_UNCONNECTED__1517, 
        SYNOPSYS_UNCONNECTED__1518, SYNOPSYS_UNCONNECTED__1519, 
        SYNOPSYS_UNCONNECTED__1520, N65823, N65822, N65821, N65820, N65819, 
        N65818}) );
  hamming_N16000_CC2_DW01_add_265 add_2931_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62351, N62350, N62349, N62348, 
        N62347}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62364, 
        N62363, N62362, N62361, N62360}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1521, SYNOPSYS_UNCONNECTED__1522, 
        SYNOPSYS_UNCONNECTED__1523, SYNOPSYS_UNCONNECTED__1524, 
        SYNOPSYS_UNCONNECTED__1525, SYNOPSYS_UNCONNECTED__1526, 
        SYNOPSYS_UNCONNECTED__1527, N65810, N65809, N65808, N65807, N65806, 
        N65805}) );
  hamming_N16000_CC2_DW01_add_266 add_2932_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62325, N62324, N62323, N62322, 
        N62321}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62338, 
        N62337, N62336, N62335, N62334}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1528, SYNOPSYS_UNCONNECTED__1529, 
        SYNOPSYS_UNCONNECTED__1530, SYNOPSYS_UNCONNECTED__1531, 
        SYNOPSYS_UNCONNECTED__1532, SYNOPSYS_UNCONNECTED__1533, 
        SYNOPSYS_UNCONNECTED__1534, N65797, N65796, N65795, N65794, N65793, 
        N65792}) );
  hamming_N16000_CC2_DW01_add_267 add_2933_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62299, N62298, N62297, N62296, 
        N62295}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62312, 
        N62311, N62310, N62309, N62308}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1535, SYNOPSYS_UNCONNECTED__1536, 
        SYNOPSYS_UNCONNECTED__1537, SYNOPSYS_UNCONNECTED__1538, 
        SYNOPSYS_UNCONNECTED__1539, SYNOPSYS_UNCONNECTED__1540, 
        SYNOPSYS_UNCONNECTED__1541, N65784, N65783, N65782, N65781, N65780, 
        N65779}) );
  hamming_N16000_CC2_DW01_add_268 add_2934_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62273, N62272, N62271, N62270, 
        N62269}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62286, 
        N62285, N62284, N62283, N62282}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1542, SYNOPSYS_UNCONNECTED__1543, 
        SYNOPSYS_UNCONNECTED__1544, SYNOPSYS_UNCONNECTED__1545, 
        SYNOPSYS_UNCONNECTED__1546, SYNOPSYS_UNCONNECTED__1547, 
        SYNOPSYS_UNCONNECTED__1548, N65771, N65770, N65769, N65768, N65767, 
        N65766}) );
  hamming_N16000_CC2_DW01_add_269 add_2935_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62247, N62246, N62245, N62244, 
        N62243}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62260, 
        N62259, N62258, N62257, N62256}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1549, SYNOPSYS_UNCONNECTED__1550, 
        SYNOPSYS_UNCONNECTED__1551, SYNOPSYS_UNCONNECTED__1552, 
        SYNOPSYS_UNCONNECTED__1553, SYNOPSYS_UNCONNECTED__1554, 
        SYNOPSYS_UNCONNECTED__1555, N65758, N65757, N65756, N65755, N65754, 
        N65753}) );
  hamming_N16000_CC2_DW01_add_270 add_2936_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62221, N62220, N62219, N62218, 
        N62217}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62234, 
        N62233, N62232, N62231, N62230}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1556, SYNOPSYS_UNCONNECTED__1557, 
        SYNOPSYS_UNCONNECTED__1558, SYNOPSYS_UNCONNECTED__1559, 
        SYNOPSYS_UNCONNECTED__1560, SYNOPSYS_UNCONNECTED__1561, 
        SYNOPSYS_UNCONNECTED__1562, N65745, N65744, N65743, N65742, N65741, 
        N65740}) );
  hamming_N16000_CC2_DW01_add_271 add_2937_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62195, N62194, N62193, N62192, 
        N62191}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62208, 
        N62207, N62206, N62205, N62204}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1563, SYNOPSYS_UNCONNECTED__1564, 
        SYNOPSYS_UNCONNECTED__1565, SYNOPSYS_UNCONNECTED__1566, 
        SYNOPSYS_UNCONNECTED__1567, SYNOPSYS_UNCONNECTED__1568, 
        SYNOPSYS_UNCONNECTED__1569, N65732, N65731, N65730, N65729, N65728, 
        N65727}) );
  hamming_N16000_CC2_DW01_add_272 add_2938_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62169, N62168, N62167, N62166, 
        N62165}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62182, 
        N62181, N62180, N62179, N62178}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1570, SYNOPSYS_UNCONNECTED__1571, 
        SYNOPSYS_UNCONNECTED__1572, SYNOPSYS_UNCONNECTED__1573, 
        SYNOPSYS_UNCONNECTED__1574, SYNOPSYS_UNCONNECTED__1575, 
        SYNOPSYS_UNCONNECTED__1576, N65719, N65718, N65717, N65716, N65715, 
        N65714}) );
  hamming_N16000_CC2_DW01_add_273 add_2939_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62143, N62142, N62141, N62140, 
        N62139}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62156, 
        N62155, N62154, N62153, N62152}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1577, SYNOPSYS_UNCONNECTED__1578, 
        SYNOPSYS_UNCONNECTED__1579, SYNOPSYS_UNCONNECTED__1580, 
        SYNOPSYS_UNCONNECTED__1581, SYNOPSYS_UNCONNECTED__1582, 
        SYNOPSYS_UNCONNECTED__1583, N65706, N65705, N65704, N65703, N65702, 
        N65701}) );
  hamming_N16000_CC2_DW01_add_274 add_2940_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62117, N62116, N62115, N62114, 
        N62113}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62130, 
        N62129, N62128, N62127, N62126}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1584, SYNOPSYS_UNCONNECTED__1585, 
        SYNOPSYS_UNCONNECTED__1586, SYNOPSYS_UNCONNECTED__1587, 
        SYNOPSYS_UNCONNECTED__1588, SYNOPSYS_UNCONNECTED__1589, 
        SYNOPSYS_UNCONNECTED__1590, N65693, N65692, N65691, N65690, N65689, 
        N65688}) );
  hamming_N16000_CC2_DW01_add_275 add_2941_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62091, N62090, N62089, N62088, 
        N62087}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62104, 
        N62103, N62102, N62101, N62100}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1591, SYNOPSYS_UNCONNECTED__1592, 
        SYNOPSYS_UNCONNECTED__1593, SYNOPSYS_UNCONNECTED__1594, 
        SYNOPSYS_UNCONNECTED__1595, SYNOPSYS_UNCONNECTED__1596, 
        SYNOPSYS_UNCONNECTED__1597, N65680, N65679, N65678, N65677, N65676, 
        N65675}) );
  hamming_N16000_CC2_DW01_add_276 add_2942_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62065, N62064, N62063, N62062, 
        N62061}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62078, 
        N62077, N62076, N62075, N62074}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1598, SYNOPSYS_UNCONNECTED__1599, 
        SYNOPSYS_UNCONNECTED__1600, SYNOPSYS_UNCONNECTED__1601, 
        SYNOPSYS_UNCONNECTED__1602, SYNOPSYS_UNCONNECTED__1603, 
        SYNOPSYS_UNCONNECTED__1604, N65667, N65666, N65665, N65664, N65663, 
        N65662}) );
  hamming_N16000_CC2_DW01_add_277 add_2943_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62039, N62038, N62037, N62036, 
        N62035}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62052, 
        N62051, N62050, N62049, N62048}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1605, SYNOPSYS_UNCONNECTED__1606, 
        SYNOPSYS_UNCONNECTED__1607, SYNOPSYS_UNCONNECTED__1608, 
        SYNOPSYS_UNCONNECTED__1609, SYNOPSYS_UNCONNECTED__1610, 
        SYNOPSYS_UNCONNECTED__1611, N65654, N65653, N65652, N65651, N65650, 
        N65649}) );
  hamming_N16000_CC2_DW01_add_278 add_2944_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62013, N62012, N62011, N62010, 
        N62009}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62026, 
        N62025, N62024, N62023, N62022}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1612, SYNOPSYS_UNCONNECTED__1613, 
        SYNOPSYS_UNCONNECTED__1614, SYNOPSYS_UNCONNECTED__1615, 
        SYNOPSYS_UNCONNECTED__1616, SYNOPSYS_UNCONNECTED__1617, 
        SYNOPSYS_UNCONNECTED__1618, N65641, N65640, N65639, N65638, N65637, 
        N65636}) );
  hamming_N16000_CC2_DW01_add_279 add_2945_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61987, N61986, N61985, N61984, 
        N61983}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N62000, 
        N61999, N61998, N61997, N61996}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1619, SYNOPSYS_UNCONNECTED__1620, 
        SYNOPSYS_UNCONNECTED__1621, SYNOPSYS_UNCONNECTED__1622, 
        SYNOPSYS_UNCONNECTED__1623, SYNOPSYS_UNCONNECTED__1624, 
        SYNOPSYS_UNCONNECTED__1625, N65628, N65627, N65626, N65625, N65624, 
        N65623}) );
  hamming_N16000_CC2_DW01_add_280 add_2946_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61961, N61960, N61959, N61958, 
        N61957}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61974, 
        N61973, N61972, N61971, N61970}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1626, SYNOPSYS_UNCONNECTED__1627, 
        SYNOPSYS_UNCONNECTED__1628, SYNOPSYS_UNCONNECTED__1629, 
        SYNOPSYS_UNCONNECTED__1630, SYNOPSYS_UNCONNECTED__1631, 
        SYNOPSYS_UNCONNECTED__1632, N65615, N65614, N65613, N65612, N65611, 
        N65610}) );
  hamming_N16000_CC2_DW01_add_281 add_2947_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61935, N61934, N61933, N61932, 
        N61931}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61948, 
        N61947, N61946, N61945, N61944}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1633, SYNOPSYS_UNCONNECTED__1634, 
        SYNOPSYS_UNCONNECTED__1635, SYNOPSYS_UNCONNECTED__1636, 
        SYNOPSYS_UNCONNECTED__1637, SYNOPSYS_UNCONNECTED__1638, 
        SYNOPSYS_UNCONNECTED__1639, N65602, N65601, N65600, N65599, N65598, 
        N65597}) );
  hamming_N16000_CC2_DW01_add_282 add_2948_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61909, N61908, N61907, N61906, 
        N61905}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61922, 
        N61921, N61920, N61919, N61918}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1640, SYNOPSYS_UNCONNECTED__1641, 
        SYNOPSYS_UNCONNECTED__1642, SYNOPSYS_UNCONNECTED__1643, 
        SYNOPSYS_UNCONNECTED__1644, SYNOPSYS_UNCONNECTED__1645, 
        SYNOPSYS_UNCONNECTED__1646, N65589, N65588, N65587, N65586, N65585, 
        N65584}) );
  hamming_N16000_CC2_DW01_add_283 add_2949_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61883, N61882, N61881, N61880, 
        N61879}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61896, 
        N61895, N61894, N61893, N61892}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1647, SYNOPSYS_UNCONNECTED__1648, 
        SYNOPSYS_UNCONNECTED__1649, SYNOPSYS_UNCONNECTED__1650, 
        SYNOPSYS_UNCONNECTED__1651, SYNOPSYS_UNCONNECTED__1652, 
        SYNOPSYS_UNCONNECTED__1653, N65576, N65575, N65574, N65573, N65572, 
        N65571}) );
  hamming_N16000_CC2_DW01_add_284 add_2950_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61857, N61856, N61855, N61854, 
        N61853}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61870, 
        N61869, N61868, N61867, N61866}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1654, SYNOPSYS_UNCONNECTED__1655, 
        SYNOPSYS_UNCONNECTED__1656, SYNOPSYS_UNCONNECTED__1657, 
        SYNOPSYS_UNCONNECTED__1658, SYNOPSYS_UNCONNECTED__1659, 
        SYNOPSYS_UNCONNECTED__1660, N65563, N65562, N65561, N65560, N65559, 
        N65558}) );
  hamming_N16000_CC2_DW01_add_285 add_2951_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61831, N61830, N61829, N61828, 
        N61827}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61844, 
        N61843, N61842, N61841, N61840}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1661, SYNOPSYS_UNCONNECTED__1662, 
        SYNOPSYS_UNCONNECTED__1663, SYNOPSYS_UNCONNECTED__1664, 
        SYNOPSYS_UNCONNECTED__1665, SYNOPSYS_UNCONNECTED__1666, 
        SYNOPSYS_UNCONNECTED__1667, N65550, N65549, N65548, N65547, N65546, 
        N65545}) );
  hamming_N16000_CC2_DW01_add_286 add_2952_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61805, N61804, N61803, N61802, 
        N61801}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61818, 
        N61817, N61816, N61815, N61814}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1668, SYNOPSYS_UNCONNECTED__1669, 
        SYNOPSYS_UNCONNECTED__1670, SYNOPSYS_UNCONNECTED__1671, 
        SYNOPSYS_UNCONNECTED__1672, SYNOPSYS_UNCONNECTED__1673, 
        SYNOPSYS_UNCONNECTED__1674, N65537, N65536, N65535, N65534, N65533, 
        N65532}) );
  hamming_N16000_CC2_DW01_add_287 add_2953_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61779, N61778, N61777, N61776, 
        N61775}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61792, 
        N61791, N61790, N61789, N61788}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1675, SYNOPSYS_UNCONNECTED__1676, 
        SYNOPSYS_UNCONNECTED__1677, SYNOPSYS_UNCONNECTED__1678, 
        SYNOPSYS_UNCONNECTED__1679, SYNOPSYS_UNCONNECTED__1680, 
        SYNOPSYS_UNCONNECTED__1681, N65524, N65523, N65522, N65521, N65520, 
        N65519}) );
  hamming_N16000_CC2_DW01_add_288 add_2954_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61753, N61752, N61751, N61750, 
        N61749}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61766, 
        N61765, N61764, N61763, N61762}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1682, SYNOPSYS_UNCONNECTED__1683, 
        SYNOPSYS_UNCONNECTED__1684, SYNOPSYS_UNCONNECTED__1685, 
        SYNOPSYS_UNCONNECTED__1686, SYNOPSYS_UNCONNECTED__1687, 
        SYNOPSYS_UNCONNECTED__1688, N65511, N65510, N65509, N65508, N65507, 
        N65506}) );
  hamming_N16000_CC2_DW01_add_289 add_2955_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61727, N61726, N61725, N61724, 
        N61723}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61740, 
        N61739, N61738, N61737, N61736}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1689, SYNOPSYS_UNCONNECTED__1690, 
        SYNOPSYS_UNCONNECTED__1691, SYNOPSYS_UNCONNECTED__1692, 
        SYNOPSYS_UNCONNECTED__1693, SYNOPSYS_UNCONNECTED__1694, 
        SYNOPSYS_UNCONNECTED__1695, N65498, N65497, N65496, N65495, N65494, 
        N65493}) );
  hamming_N16000_CC2_DW01_add_290 add_2956_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61701, N61700, N61699, N61698, 
        N61697}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61714, 
        N61713, N61712, N61711, N61710}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1696, SYNOPSYS_UNCONNECTED__1697, 
        SYNOPSYS_UNCONNECTED__1698, SYNOPSYS_UNCONNECTED__1699, 
        SYNOPSYS_UNCONNECTED__1700, SYNOPSYS_UNCONNECTED__1701, 
        SYNOPSYS_UNCONNECTED__1702, N65485, N65484, N65483, N65482, N65481, 
        N65480}) );
  hamming_N16000_CC2_DW01_add_291 add_2957_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61675, N61674, N61673, N61672, 
        N61671}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61688, 
        N61687, N61686, N61685, N61684}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1703, SYNOPSYS_UNCONNECTED__1704, 
        SYNOPSYS_UNCONNECTED__1705, SYNOPSYS_UNCONNECTED__1706, 
        SYNOPSYS_UNCONNECTED__1707, SYNOPSYS_UNCONNECTED__1708, 
        SYNOPSYS_UNCONNECTED__1709, N65472, N65471, N65470, N65469, N65468, 
        N65467}) );
  hamming_N16000_CC2_DW01_add_292 add_2958_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61649, N61648, N61647, N61646, 
        N61645}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61662, 
        N61661, N61660, N61659, N61658}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1710, SYNOPSYS_UNCONNECTED__1711, 
        SYNOPSYS_UNCONNECTED__1712, SYNOPSYS_UNCONNECTED__1713, 
        SYNOPSYS_UNCONNECTED__1714, SYNOPSYS_UNCONNECTED__1715, 
        SYNOPSYS_UNCONNECTED__1716, N65459, N65458, N65457, N65456, N65455, 
        N65454}) );
  hamming_N16000_CC2_DW01_add_293 add_2959_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61623, N61622, N61621, N61620, 
        N61619}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61636, 
        N61635, N61634, N61633, N61632}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1717, SYNOPSYS_UNCONNECTED__1718, 
        SYNOPSYS_UNCONNECTED__1719, SYNOPSYS_UNCONNECTED__1720, 
        SYNOPSYS_UNCONNECTED__1721, SYNOPSYS_UNCONNECTED__1722, 
        SYNOPSYS_UNCONNECTED__1723, N65446, N65445, N65444, N65443, N65442, 
        N65441}) );
  hamming_N16000_CC2_DW01_add_294 add_2960_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61597, N61596, N61595, N61594, 
        N61593}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61610, 
        N61609, N61608, N61607, N61606}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1724, SYNOPSYS_UNCONNECTED__1725, 
        SYNOPSYS_UNCONNECTED__1726, SYNOPSYS_UNCONNECTED__1727, 
        SYNOPSYS_UNCONNECTED__1728, SYNOPSYS_UNCONNECTED__1729, 
        SYNOPSYS_UNCONNECTED__1730, N65433, N65432, N65431, N65430, N65429, 
        N65428}) );
  hamming_N16000_CC2_DW01_add_295 add_2961_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61571, N61570, N61569, N61568, 
        N61567}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61584, 
        N61583, N61582, N61581, N61580}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1731, SYNOPSYS_UNCONNECTED__1732, 
        SYNOPSYS_UNCONNECTED__1733, SYNOPSYS_UNCONNECTED__1734, 
        SYNOPSYS_UNCONNECTED__1735, SYNOPSYS_UNCONNECTED__1736, 
        SYNOPSYS_UNCONNECTED__1737, N65420, N65419, N65418, N65417, N65416, 
        N65415}) );
  hamming_N16000_CC2_DW01_add_296 add_2962_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61545, N61544, N61543, N61542, 
        N61541}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61558, 
        N61557, N61556, N61555, N61554}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1738, SYNOPSYS_UNCONNECTED__1739, 
        SYNOPSYS_UNCONNECTED__1740, SYNOPSYS_UNCONNECTED__1741, 
        SYNOPSYS_UNCONNECTED__1742, SYNOPSYS_UNCONNECTED__1743, 
        SYNOPSYS_UNCONNECTED__1744, N65407, N65406, N65405, N65404, N65403, 
        N65402}) );
  hamming_N16000_CC2_DW01_add_297 add_2963_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61519, N61518, N61517, N61516, 
        N61515}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61532, 
        N61531, N61530, N61529, N61528}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1745, SYNOPSYS_UNCONNECTED__1746, 
        SYNOPSYS_UNCONNECTED__1747, SYNOPSYS_UNCONNECTED__1748, 
        SYNOPSYS_UNCONNECTED__1749, SYNOPSYS_UNCONNECTED__1750, 
        SYNOPSYS_UNCONNECTED__1751, N65394, N65393, N65392, N65391, N65390, 
        N65389}) );
  hamming_N16000_CC2_DW01_add_298 add_2964_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61493, N61492, N61491, N61490, 
        N61489}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61506, 
        N61505, N61504, N61503, N61502}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1752, SYNOPSYS_UNCONNECTED__1753, 
        SYNOPSYS_UNCONNECTED__1754, SYNOPSYS_UNCONNECTED__1755, 
        SYNOPSYS_UNCONNECTED__1756, SYNOPSYS_UNCONNECTED__1757, 
        SYNOPSYS_UNCONNECTED__1758, N65381, N65380, N65379, N65378, N65377, 
        N65376}) );
  hamming_N16000_CC2_DW01_add_299 add_2965_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61467, N61466, N61465, N61464, 
        N61463}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61480, 
        N61479, N61478, N61477, N61476}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1759, SYNOPSYS_UNCONNECTED__1760, 
        SYNOPSYS_UNCONNECTED__1761, SYNOPSYS_UNCONNECTED__1762, 
        SYNOPSYS_UNCONNECTED__1763, SYNOPSYS_UNCONNECTED__1764, 
        SYNOPSYS_UNCONNECTED__1765, N65368, N65367, N65366, N65365, N65364, 
        N65363}) );
  hamming_N16000_CC2_DW01_add_300 add_2966_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61441, N61440, N61439, N61438, 
        N61437}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61454, 
        N61453, N61452, N61451, N61450}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1766, SYNOPSYS_UNCONNECTED__1767, 
        SYNOPSYS_UNCONNECTED__1768, SYNOPSYS_UNCONNECTED__1769, 
        SYNOPSYS_UNCONNECTED__1770, SYNOPSYS_UNCONNECTED__1771, 
        SYNOPSYS_UNCONNECTED__1772, N65355, N65354, N65353, N65352, N65351, 
        N65350}) );
  hamming_N16000_CC2_DW01_add_301 add_2967_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61415, N61414, N61413, N61412, 
        N61411}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61428, 
        N61427, N61426, N61425, N61424}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1773, SYNOPSYS_UNCONNECTED__1774, 
        SYNOPSYS_UNCONNECTED__1775, SYNOPSYS_UNCONNECTED__1776, 
        SYNOPSYS_UNCONNECTED__1777, SYNOPSYS_UNCONNECTED__1778, 
        SYNOPSYS_UNCONNECTED__1779, N65342, N65341, N65340, N65339, N65338, 
        N65337}) );
  hamming_N16000_CC2_DW01_add_302 add_2968_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61389, N61388, N61387, N61386, 
        N61385}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61402, 
        N61401, N61400, N61399, N61398}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1780, SYNOPSYS_UNCONNECTED__1781, 
        SYNOPSYS_UNCONNECTED__1782, SYNOPSYS_UNCONNECTED__1783, 
        SYNOPSYS_UNCONNECTED__1784, SYNOPSYS_UNCONNECTED__1785, 
        SYNOPSYS_UNCONNECTED__1786, N65329, N65328, N65327, N65326, N65325, 
        N65324}) );
  hamming_N16000_CC2_DW01_add_303 add_2969_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61363, N61362, N61361, N61360, 
        N61359}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61376, 
        N61375, N61374, N61373, N61372}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1787, SYNOPSYS_UNCONNECTED__1788, 
        SYNOPSYS_UNCONNECTED__1789, SYNOPSYS_UNCONNECTED__1790, 
        SYNOPSYS_UNCONNECTED__1791, SYNOPSYS_UNCONNECTED__1792, 
        SYNOPSYS_UNCONNECTED__1793, N65316, N65315, N65314, N65313, N65312, 
        N65311}) );
  hamming_N16000_CC2_DW01_add_304 add_2970_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61337, N61336, N61335, N61334, 
        N61333}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61350, 
        N61349, N61348, N61347, N61346}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1794, SYNOPSYS_UNCONNECTED__1795, 
        SYNOPSYS_UNCONNECTED__1796, SYNOPSYS_UNCONNECTED__1797, 
        SYNOPSYS_UNCONNECTED__1798, SYNOPSYS_UNCONNECTED__1799, 
        SYNOPSYS_UNCONNECTED__1800, N65303, N65302, N65301, N65300, N65299, 
        N65298}) );
  hamming_N16000_CC2_DW01_add_305 add_2971_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61311, N61310, N61309, N61308, 
        N61307}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61324, 
        N61323, N61322, N61321, N61320}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1801, SYNOPSYS_UNCONNECTED__1802, 
        SYNOPSYS_UNCONNECTED__1803, SYNOPSYS_UNCONNECTED__1804, 
        SYNOPSYS_UNCONNECTED__1805, SYNOPSYS_UNCONNECTED__1806, 
        SYNOPSYS_UNCONNECTED__1807, N65290, N65289, N65288, N65287, N65286, 
        N65285}) );
  hamming_N16000_CC2_DW01_add_306 add_2972_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61285, N61284, N61283, N61282, 
        N61281}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61298, 
        N61297, N61296, N61295, N61294}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1808, SYNOPSYS_UNCONNECTED__1809, 
        SYNOPSYS_UNCONNECTED__1810, SYNOPSYS_UNCONNECTED__1811, 
        SYNOPSYS_UNCONNECTED__1812, SYNOPSYS_UNCONNECTED__1813, 
        SYNOPSYS_UNCONNECTED__1814, N65277, N65276, N65275, N65274, N65273, 
        N65272}) );
  hamming_N16000_CC2_DW01_add_307 add_2973_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61259, N61258, N61257, N61256, 
        N61255}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61272, 
        N61271, N61270, N61269, N61268}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1815, SYNOPSYS_UNCONNECTED__1816, 
        SYNOPSYS_UNCONNECTED__1817, SYNOPSYS_UNCONNECTED__1818, 
        SYNOPSYS_UNCONNECTED__1819, SYNOPSYS_UNCONNECTED__1820, 
        SYNOPSYS_UNCONNECTED__1821, N65264, N65263, N65262, N65261, N65260, 
        N65259}) );
  hamming_N16000_CC2_DW01_add_308 add_2974_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61233, N61232, N61231, N61230, 
        N61229}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61246, 
        N61245, N61244, N61243, N61242}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1822, SYNOPSYS_UNCONNECTED__1823, 
        SYNOPSYS_UNCONNECTED__1824, SYNOPSYS_UNCONNECTED__1825, 
        SYNOPSYS_UNCONNECTED__1826, SYNOPSYS_UNCONNECTED__1827, 
        SYNOPSYS_UNCONNECTED__1828, N65251, N65250, N65249, N65248, N65247, 
        N65246}) );
  hamming_N16000_CC2_DW01_add_309 add_2975_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61207, N61206, N61205, N61204, 
        N61203}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61220, 
        N61219, N61218, N61217, N61216}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1829, SYNOPSYS_UNCONNECTED__1830, 
        SYNOPSYS_UNCONNECTED__1831, SYNOPSYS_UNCONNECTED__1832, 
        SYNOPSYS_UNCONNECTED__1833, SYNOPSYS_UNCONNECTED__1834, 
        SYNOPSYS_UNCONNECTED__1835, N65238, N65237, N65236, N65235, N65234, 
        N65233}) );
  hamming_N16000_CC2_DW01_add_310 add_2976_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61181, N61180, N61179, N61178, 
        N61177}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61194, 
        N61193, N61192, N61191, N61190}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1836, SYNOPSYS_UNCONNECTED__1837, 
        SYNOPSYS_UNCONNECTED__1838, SYNOPSYS_UNCONNECTED__1839, 
        SYNOPSYS_UNCONNECTED__1840, SYNOPSYS_UNCONNECTED__1841, 
        SYNOPSYS_UNCONNECTED__1842, N65225, N65224, N65223, N65222, N65221, 
        N65220}) );
  hamming_N16000_CC2_DW01_add_311 add_2977_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61155, N61154, N61153, N61152, 
        N61151}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61168, 
        N61167, N61166, N61165, N61164}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1843, SYNOPSYS_UNCONNECTED__1844, 
        SYNOPSYS_UNCONNECTED__1845, SYNOPSYS_UNCONNECTED__1846, 
        SYNOPSYS_UNCONNECTED__1847, SYNOPSYS_UNCONNECTED__1848, 
        SYNOPSYS_UNCONNECTED__1849, N65212, N65211, N65210, N65209, N65208, 
        N65207}) );
  hamming_N16000_CC2_DW01_add_312 add_2978_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61129, N61128, N61127, N61126, 
        N61125}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61142, 
        N61141, N61140, N61139, N61138}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1850, SYNOPSYS_UNCONNECTED__1851, 
        SYNOPSYS_UNCONNECTED__1852, SYNOPSYS_UNCONNECTED__1853, 
        SYNOPSYS_UNCONNECTED__1854, SYNOPSYS_UNCONNECTED__1855, 
        SYNOPSYS_UNCONNECTED__1856, N65199, N65198, N65197, N65196, N65195, 
        N65194}) );
  hamming_N16000_CC2_DW01_add_313 add_2979_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61103, N61102, N61101, N61100, 
        N61099}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61116, 
        N61115, N61114, N61113, N61112}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1857, SYNOPSYS_UNCONNECTED__1858, 
        SYNOPSYS_UNCONNECTED__1859, SYNOPSYS_UNCONNECTED__1860, 
        SYNOPSYS_UNCONNECTED__1861, SYNOPSYS_UNCONNECTED__1862, 
        SYNOPSYS_UNCONNECTED__1863, N65186, N65185, N65184, N65183, N65182, 
        N65181}) );
  hamming_N16000_CC2_DW01_add_314 add_2980_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61077, N61076, N61075, N61074, 
        N61073}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61090, 
        N61089, N61088, N61087, N61086}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1864, SYNOPSYS_UNCONNECTED__1865, 
        SYNOPSYS_UNCONNECTED__1866, SYNOPSYS_UNCONNECTED__1867, 
        SYNOPSYS_UNCONNECTED__1868, SYNOPSYS_UNCONNECTED__1869, 
        SYNOPSYS_UNCONNECTED__1870, N65173, N65172, N65171, N65170, N65169, 
        N65168}) );
  hamming_N16000_CC2_DW01_add_315 add_2981_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61051, N61050, N61049, N61048, 
        N61047}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61064, 
        N61063, N61062, N61061, N61060}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1871, SYNOPSYS_UNCONNECTED__1872, 
        SYNOPSYS_UNCONNECTED__1873, SYNOPSYS_UNCONNECTED__1874, 
        SYNOPSYS_UNCONNECTED__1875, SYNOPSYS_UNCONNECTED__1876, 
        SYNOPSYS_UNCONNECTED__1877, N65160, N65159, N65158, N65157, N65156, 
        N65155}) );
  hamming_N16000_CC2_DW01_add_316 add_2982_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61025, N61024, N61023, N61022, 
        N61021}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61038, 
        N61037, N61036, N61035, N61034}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1878, SYNOPSYS_UNCONNECTED__1879, 
        SYNOPSYS_UNCONNECTED__1880, SYNOPSYS_UNCONNECTED__1881, 
        SYNOPSYS_UNCONNECTED__1882, SYNOPSYS_UNCONNECTED__1883, 
        SYNOPSYS_UNCONNECTED__1884, N65147, N65146, N65145, N65144, N65143, 
        N65142}) );
  hamming_N16000_CC2_DW01_add_317 add_2983_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60999, N60998, N60997, N60996, 
        N60995}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N61012, 
        N61011, N61010, N61009, N61008}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1885, SYNOPSYS_UNCONNECTED__1886, 
        SYNOPSYS_UNCONNECTED__1887, SYNOPSYS_UNCONNECTED__1888, 
        SYNOPSYS_UNCONNECTED__1889, SYNOPSYS_UNCONNECTED__1890, 
        SYNOPSYS_UNCONNECTED__1891, N65134, N65133, N65132, N65131, N65130, 
        N65129}) );
  hamming_N16000_CC2_DW01_add_318 add_2984_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60973, N60972, N60971, N60970, 
        N60969}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60986, 
        N60985, N60984, N60983, N60982}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1892, SYNOPSYS_UNCONNECTED__1893, 
        SYNOPSYS_UNCONNECTED__1894, SYNOPSYS_UNCONNECTED__1895, 
        SYNOPSYS_UNCONNECTED__1896, SYNOPSYS_UNCONNECTED__1897, 
        SYNOPSYS_UNCONNECTED__1898, N65121, N65120, N65119, N65118, N65117, 
        N65116}) );
  hamming_N16000_CC2_DW01_add_319 add_2985_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60947, N60946, N60945, N60944, 
        N60943}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60960, 
        N60959, N60958, N60957, N60956}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1899, SYNOPSYS_UNCONNECTED__1900, 
        SYNOPSYS_UNCONNECTED__1901, SYNOPSYS_UNCONNECTED__1902, 
        SYNOPSYS_UNCONNECTED__1903, SYNOPSYS_UNCONNECTED__1904, 
        SYNOPSYS_UNCONNECTED__1905, N65108, N65107, N65106, N65105, N65104, 
        N65103}) );
  hamming_N16000_CC2_DW01_add_320 add_2986_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60921, N60920, N60919, N60918, 
        N60917}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60934, 
        N60933, N60932, N60931, N60930}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1906, SYNOPSYS_UNCONNECTED__1907, 
        SYNOPSYS_UNCONNECTED__1908, SYNOPSYS_UNCONNECTED__1909, 
        SYNOPSYS_UNCONNECTED__1910, SYNOPSYS_UNCONNECTED__1911, 
        SYNOPSYS_UNCONNECTED__1912, N65095, N65094, N65093, N65092, N65091, 
        N65090}) );
  hamming_N16000_CC2_DW01_add_321 add_2987_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60895, N60894, N60893, N60892, 
        N60891}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60908, 
        N60907, N60906, N60905, N60904}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1913, SYNOPSYS_UNCONNECTED__1914, 
        SYNOPSYS_UNCONNECTED__1915, SYNOPSYS_UNCONNECTED__1916, 
        SYNOPSYS_UNCONNECTED__1917, SYNOPSYS_UNCONNECTED__1918, 
        SYNOPSYS_UNCONNECTED__1919, N65082, N65081, N65080, N65079, N65078, 
        N65077}) );
  hamming_N16000_CC2_DW01_add_322 add_2988_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60869, N60868, N60867, N60866, 
        N60865}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60882, 
        N60881, N60880, N60879, N60878}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1920, SYNOPSYS_UNCONNECTED__1921, 
        SYNOPSYS_UNCONNECTED__1922, SYNOPSYS_UNCONNECTED__1923, 
        SYNOPSYS_UNCONNECTED__1924, SYNOPSYS_UNCONNECTED__1925, 
        SYNOPSYS_UNCONNECTED__1926, N65069, N65068, N65067, N65066, N65065, 
        N65064}) );
  hamming_N16000_CC2_DW01_add_323 add_2989_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60843, N60842, N60841, N60840, 
        N60839}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60856, 
        N60855, N60854, N60853, N60852}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1927, SYNOPSYS_UNCONNECTED__1928, 
        SYNOPSYS_UNCONNECTED__1929, SYNOPSYS_UNCONNECTED__1930, 
        SYNOPSYS_UNCONNECTED__1931, SYNOPSYS_UNCONNECTED__1932, 
        SYNOPSYS_UNCONNECTED__1933, N65056, N65055, N65054, N65053, N65052, 
        N65051}) );
  hamming_N16000_CC2_DW01_add_324 add_2990_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60817, N60816, N60815, N60814, 
        N60813}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60830, 
        N60829, N60828, N60827, N60826}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1934, SYNOPSYS_UNCONNECTED__1935, 
        SYNOPSYS_UNCONNECTED__1936, SYNOPSYS_UNCONNECTED__1937, 
        SYNOPSYS_UNCONNECTED__1938, SYNOPSYS_UNCONNECTED__1939, 
        SYNOPSYS_UNCONNECTED__1940, N65043, N65042, N65041, N65040, N65039, 
        N65038}) );
  hamming_N16000_CC2_DW01_add_325 add_2991_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60791, N60790, N60789, N60788, 
        N60787}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60804, 
        N60803, N60802, N60801, N60800}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1941, SYNOPSYS_UNCONNECTED__1942, 
        SYNOPSYS_UNCONNECTED__1943, SYNOPSYS_UNCONNECTED__1944, 
        SYNOPSYS_UNCONNECTED__1945, SYNOPSYS_UNCONNECTED__1946, 
        SYNOPSYS_UNCONNECTED__1947, N65030, N65029, N65028, N65027, N65026, 
        N65025}) );
  hamming_N16000_CC2_DW01_add_326 add_2992_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60765, N60764, N60763, N60762, 
        N60761}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60778, 
        N60777, N60776, N60775, N60774}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1948, SYNOPSYS_UNCONNECTED__1949, 
        SYNOPSYS_UNCONNECTED__1950, SYNOPSYS_UNCONNECTED__1951, 
        SYNOPSYS_UNCONNECTED__1952, SYNOPSYS_UNCONNECTED__1953, 
        SYNOPSYS_UNCONNECTED__1954, N65017, N65016, N65015, N65014, N65013, 
        N65012}) );
  hamming_N16000_CC2_DW01_add_327 add_2993_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60739, N60738, N60737, N60736, 
        N60735}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60752, 
        N60751, N60750, N60749, N60748}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1955, SYNOPSYS_UNCONNECTED__1956, 
        SYNOPSYS_UNCONNECTED__1957, SYNOPSYS_UNCONNECTED__1958, 
        SYNOPSYS_UNCONNECTED__1959, SYNOPSYS_UNCONNECTED__1960, 
        SYNOPSYS_UNCONNECTED__1961, N65004, N65003, N65002, N65001, N65000, 
        N64999}) );
  hamming_N16000_CC2_DW01_add_328 add_2994_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60713, N60712, N60711, N60710, 
        N60709}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60726, 
        N60725, N60724, N60723, N60722}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1962, SYNOPSYS_UNCONNECTED__1963, 
        SYNOPSYS_UNCONNECTED__1964, SYNOPSYS_UNCONNECTED__1965, 
        SYNOPSYS_UNCONNECTED__1966, SYNOPSYS_UNCONNECTED__1967, 
        SYNOPSYS_UNCONNECTED__1968, N64991, N64990, N64989, N64988, N64987, 
        N64986}) );
  hamming_N16000_CC2_DW01_add_329 add_2995_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60687, N60686, N60685, N60684, 
        N60683}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60700, 
        N60699, N60698, N60697, N60696}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1969, SYNOPSYS_UNCONNECTED__1970, 
        SYNOPSYS_UNCONNECTED__1971, SYNOPSYS_UNCONNECTED__1972, 
        SYNOPSYS_UNCONNECTED__1973, SYNOPSYS_UNCONNECTED__1974, 
        SYNOPSYS_UNCONNECTED__1975, N64978, N64977, N64976, N64975, N64974, 
        N64973}) );
  hamming_N16000_CC2_DW01_add_330 add_2996_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60661, N60660, N60659, N60658, 
        N60657}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60674, 
        N60673, N60672, N60671, N60670}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1976, SYNOPSYS_UNCONNECTED__1977, 
        SYNOPSYS_UNCONNECTED__1978, SYNOPSYS_UNCONNECTED__1979, 
        SYNOPSYS_UNCONNECTED__1980, SYNOPSYS_UNCONNECTED__1981, 
        SYNOPSYS_UNCONNECTED__1982, N64965, N64964, N64963, N64962, N64961, 
        N64960}) );
  hamming_N16000_CC2_DW01_add_331 add_2997_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60635, N60634, N60633, N60632, 
        N60631}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60648, 
        N60647, N60646, N60645, N60644}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1983, SYNOPSYS_UNCONNECTED__1984, 
        SYNOPSYS_UNCONNECTED__1985, SYNOPSYS_UNCONNECTED__1986, 
        SYNOPSYS_UNCONNECTED__1987, SYNOPSYS_UNCONNECTED__1988, 
        SYNOPSYS_UNCONNECTED__1989, N64952, N64951, N64950, N64949, N64948, 
        N64947}) );
  hamming_N16000_CC2_DW01_add_332 add_2998_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60609, N60608, N60607, N60606, 
        N60605}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60622, 
        N60621, N60620, N60619, N60618}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1990, SYNOPSYS_UNCONNECTED__1991, 
        SYNOPSYS_UNCONNECTED__1992, SYNOPSYS_UNCONNECTED__1993, 
        SYNOPSYS_UNCONNECTED__1994, SYNOPSYS_UNCONNECTED__1995, 
        SYNOPSYS_UNCONNECTED__1996, N64939, N64938, N64937, N64936, N64935, 
        N64934}) );
  hamming_N16000_CC2_DW01_add_333 add_2999_root_add_71_I832 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60582, N60581, N60580, 
        N60579}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, N60596, 
        N60595, N60594, N60593, N60592}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1997, SYNOPSYS_UNCONNECTED__1998, 
        SYNOPSYS_UNCONNECTED__1999, SYNOPSYS_UNCONNECTED__2000, 
        SYNOPSYS_UNCONNECTED__2001, SYNOPSYS_UNCONNECTED__2002, 
        SYNOPSYS_UNCONNECTED__2003, N64926, N64925, N64924, N64923, N64922, 
        N64921}) );
  NAND U13350 ( .A(n5351), .B(n5352), .Z(N64912) );
  NAND U13351 ( .A(n5353), .B(n5354), .Z(n5352) );
  NANDN U13352 ( .A(n5355), .B(n5356), .Z(n5354) );
  NANDN U13353 ( .A(n5356), .B(n5355), .Z(n5351) );
  XOR U13354 ( .A(n5355), .B(n5357), .Z(N64911) );
  XNOR U13355 ( .A(n5353), .B(n5356), .Z(n5357) );
  NAND U13356 ( .A(n5358), .B(n5359), .Z(n5356) );
  NAND U13357 ( .A(n5360), .B(n5361), .Z(n5359) );
  NANDN U13358 ( .A(n5362), .B(n5363), .Z(n5361) );
  NANDN U13359 ( .A(n5363), .B(n5362), .Z(n5358) );
  AND U13360 ( .A(n5364), .B(n5365), .Z(n5353) );
  NAND U13361 ( .A(n5366), .B(n5367), .Z(n5365) );
  NANDN U13362 ( .A(n5368), .B(n5369), .Z(n5367) );
  NANDN U13363 ( .A(n5369), .B(n5368), .Z(n5364) );
  IV U13364 ( .A(n5370), .Z(n5369) );
  AND U13365 ( .A(n5371), .B(n5372), .Z(n5355) );
  NAND U13366 ( .A(n5373), .B(n5374), .Z(n5372) );
  NANDN U13367 ( .A(n5375), .B(n5376), .Z(n5374) );
  NANDN U13368 ( .A(n5376), .B(n5375), .Z(n5371) );
  XOR U13369 ( .A(n5368), .B(n5377), .Z(N64910) );
  XNOR U13370 ( .A(n5366), .B(n5370), .Z(n5377) );
  XOR U13371 ( .A(n5363), .B(n5378), .Z(n5370) );
  XNOR U13372 ( .A(n5360), .B(n5362), .Z(n5378) );
  AND U13373 ( .A(n5379), .B(n5380), .Z(n5362) );
  NANDN U13374 ( .A(n5381), .B(n5382), .Z(n5380) );
  OR U13375 ( .A(n5383), .B(n5384), .Z(n5382) );
  IV U13376 ( .A(n5385), .Z(n5384) );
  NANDN U13377 ( .A(n5385), .B(n5383), .Z(n5379) );
  AND U13378 ( .A(n5386), .B(n5387), .Z(n5360) );
  NAND U13379 ( .A(n5388), .B(n5389), .Z(n5387) );
  NANDN U13380 ( .A(n5390), .B(n5391), .Z(n5389) );
  NANDN U13381 ( .A(n5391), .B(n5390), .Z(n5386) );
  IV U13382 ( .A(n5392), .Z(n5391) );
  NAND U13383 ( .A(n5393), .B(n5394), .Z(n5363) );
  NANDN U13384 ( .A(n5395), .B(n5396), .Z(n5394) );
  NANDN U13385 ( .A(n5397), .B(n5398), .Z(n5396) );
  NANDN U13386 ( .A(n5398), .B(n5397), .Z(n5393) );
  IV U13387 ( .A(n5399), .Z(n5397) );
  AND U13388 ( .A(n5400), .B(n5401), .Z(n5366) );
  NAND U13389 ( .A(n5402), .B(n5403), .Z(n5401) );
  NANDN U13390 ( .A(n5404), .B(n5405), .Z(n5403) );
  NANDN U13391 ( .A(n5405), .B(n5404), .Z(n5400) );
  XOR U13392 ( .A(n5376), .B(n5406), .Z(n5368) );
  XNOR U13393 ( .A(n5373), .B(n5375), .Z(n5406) );
  AND U13394 ( .A(n5407), .B(n5408), .Z(n5375) );
  NANDN U13395 ( .A(n5409), .B(n5410), .Z(n5408) );
  OR U13396 ( .A(n5411), .B(n5412), .Z(n5410) );
  IV U13397 ( .A(n5413), .Z(n5412) );
  NANDN U13398 ( .A(n5413), .B(n5411), .Z(n5407) );
  AND U13399 ( .A(n5414), .B(n5415), .Z(n5373) );
  NAND U13400 ( .A(n5416), .B(n5417), .Z(n5415) );
  NANDN U13401 ( .A(n5418), .B(n5419), .Z(n5417) );
  NANDN U13402 ( .A(n5419), .B(n5418), .Z(n5414) );
  IV U13403 ( .A(n5420), .Z(n5419) );
  NAND U13404 ( .A(n5421), .B(n5422), .Z(n5376) );
  NANDN U13405 ( .A(n5423), .B(n5424), .Z(n5422) );
  NANDN U13406 ( .A(n5425), .B(n5426), .Z(n5424) );
  NANDN U13407 ( .A(n5426), .B(n5425), .Z(n5421) );
  IV U13408 ( .A(n5427), .Z(n5425) );
  XOR U13409 ( .A(n5402), .B(n5428), .Z(N64909) );
  XNOR U13410 ( .A(n5405), .B(n5404), .Z(n5428) );
  XNOR U13411 ( .A(n5416), .B(n5429), .Z(n5404) );
  XNOR U13412 ( .A(n5420), .B(n5418), .Z(n5429) );
  XOR U13413 ( .A(n5426), .B(n5430), .Z(n5418) );
  XNOR U13414 ( .A(n5423), .B(n5427), .Z(n5430) );
  AND U13415 ( .A(n5431), .B(n5432), .Z(n5427) );
  NAND U13416 ( .A(n5433), .B(n5434), .Z(n5432) );
  NAND U13417 ( .A(n5435), .B(n5436), .Z(n5431) );
  AND U13418 ( .A(n5437), .B(n5438), .Z(n5423) );
  NAND U13419 ( .A(n5439), .B(n5440), .Z(n5438) );
  NAND U13420 ( .A(n5441), .B(n5442), .Z(n5437) );
  NANDN U13421 ( .A(n5443), .B(n5444), .Z(n5426) );
  ANDN U13422 ( .B(n5445), .A(n5446), .Z(n5420) );
  XNOR U13423 ( .A(n5411), .B(n5447), .Z(n5416) );
  XNOR U13424 ( .A(n5409), .B(n5413), .Z(n5447) );
  AND U13425 ( .A(n5448), .B(n5449), .Z(n5413) );
  NAND U13426 ( .A(n5450), .B(n5451), .Z(n5449) );
  NAND U13427 ( .A(n5452), .B(n5453), .Z(n5448) );
  AND U13428 ( .A(n5454), .B(n5455), .Z(n5409) );
  NAND U13429 ( .A(n5456), .B(n5457), .Z(n5455) );
  NAND U13430 ( .A(n5458), .B(n5459), .Z(n5454) );
  AND U13431 ( .A(n5460), .B(n5461), .Z(n5411) );
  NAND U13432 ( .A(n5462), .B(n5463), .Z(n5405) );
  XNOR U13433 ( .A(n5388), .B(n5464), .Z(n5402) );
  XNOR U13434 ( .A(n5392), .B(n5390), .Z(n5464) );
  XOR U13435 ( .A(n5398), .B(n5465), .Z(n5390) );
  XNOR U13436 ( .A(n5395), .B(n5399), .Z(n5465) );
  AND U13437 ( .A(n5466), .B(n5467), .Z(n5399) );
  NAND U13438 ( .A(n5468), .B(n5469), .Z(n5467) );
  NAND U13439 ( .A(n5470), .B(n5471), .Z(n5466) );
  AND U13440 ( .A(n5472), .B(n5473), .Z(n5395) );
  NAND U13441 ( .A(n5474), .B(n5475), .Z(n5473) );
  NAND U13442 ( .A(n5476), .B(n5477), .Z(n5472) );
  NANDN U13443 ( .A(n5478), .B(n5479), .Z(n5398) );
  ANDN U13444 ( .B(n5480), .A(n5481), .Z(n5392) );
  XNOR U13445 ( .A(n5383), .B(n5482), .Z(n5388) );
  XNOR U13446 ( .A(n5381), .B(n5385), .Z(n5482) );
  AND U13447 ( .A(n5483), .B(n5484), .Z(n5385) );
  NAND U13448 ( .A(n5485), .B(n5486), .Z(n5484) );
  NAND U13449 ( .A(n5487), .B(n5488), .Z(n5483) );
  AND U13450 ( .A(n5489), .B(n5490), .Z(n5381) );
  NAND U13451 ( .A(n5491), .B(n5492), .Z(n5490) );
  NAND U13452 ( .A(n5493), .B(n5494), .Z(n5489) );
  AND U13453 ( .A(n5495), .B(n5496), .Z(n5383) );
  XOR U13454 ( .A(n5463), .B(n5462), .Z(N64908) );
  XNOR U13455 ( .A(n5480), .B(n5481), .Z(n5462) );
  XNOR U13456 ( .A(n5495), .B(n5496), .Z(n5481) );
  XOR U13457 ( .A(n5492), .B(n5491), .Z(n5496) );
  XOR U13458 ( .A(y[7980]), .B(x[7980]), .Z(n5491) );
  XOR U13459 ( .A(n5494), .B(n5493), .Z(n5492) );
  XOR U13460 ( .A(y[7982]), .B(x[7982]), .Z(n5493) );
  XOR U13461 ( .A(y[7981]), .B(x[7981]), .Z(n5494) );
  XOR U13462 ( .A(n5486), .B(n5485), .Z(n5495) );
  XOR U13463 ( .A(n5488), .B(n5487), .Z(n5485) );
  XOR U13464 ( .A(y[7979]), .B(x[7979]), .Z(n5487) );
  XOR U13465 ( .A(y[7978]), .B(x[7978]), .Z(n5488) );
  XOR U13466 ( .A(y[7977]), .B(x[7977]), .Z(n5486) );
  XNOR U13467 ( .A(n5479), .B(n5478), .Z(n5480) );
  XNOR U13468 ( .A(n5475), .B(n5474), .Z(n5478) );
  XOR U13469 ( .A(n5477), .B(n5476), .Z(n5474) );
  XOR U13470 ( .A(y[7976]), .B(x[7976]), .Z(n5476) );
  XOR U13471 ( .A(y[7975]), .B(x[7975]), .Z(n5477) );
  XOR U13472 ( .A(y[7974]), .B(x[7974]), .Z(n5475) );
  XOR U13473 ( .A(n5469), .B(n5468), .Z(n5479) );
  XOR U13474 ( .A(n5471), .B(n5470), .Z(n5468) );
  XOR U13475 ( .A(y[7973]), .B(x[7973]), .Z(n5470) );
  XOR U13476 ( .A(y[7972]), .B(x[7972]), .Z(n5471) );
  XOR U13477 ( .A(y[7971]), .B(x[7971]), .Z(n5469) );
  XNOR U13478 ( .A(n5445), .B(n5446), .Z(n5463) );
  XNOR U13479 ( .A(n5460), .B(n5461), .Z(n5446) );
  XOR U13480 ( .A(n5457), .B(n5456), .Z(n5461) );
  XOR U13481 ( .A(y[7968]), .B(x[7968]), .Z(n5456) );
  XOR U13482 ( .A(n5459), .B(n5458), .Z(n5457) );
  XOR U13483 ( .A(y[7970]), .B(x[7970]), .Z(n5458) );
  XOR U13484 ( .A(y[7969]), .B(x[7969]), .Z(n5459) );
  XOR U13485 ( .A(n5451), .B(n5450), .Z(n5460) );
  XOR U13486 ( .A(n5453), .B(n5452), .Z(n5450) );
  XOR U13487 ( .A(y[7967]), .B(x[7967]), .Z(n5452) );
  XOR U13488 ( .A(y[7966]), .B(x[7966]), .Z(n5453) );
  XOR U13489 ( .A(y[7965]), .B(x[7965]), .Z(n5451) );
  XNOR U13490 ( .A(n5444), .B(n5443), .Z(n5445) );
  XNOR U13491 ( .A(n5440), .B(n5439), .Z(n5443) );
  XOR U13492 ( .A(n5442), .B(n5441), .Z(n5439) );
  XOR U13493 ( .A(y[7964]), .B(x[7964]), .Z(n5441) );
  XOR U13494 ( .A(y[7963]), .B(x[7963]), .Z(n5442) );
  XOR U13495 ( .A(y[7962]), .B(x[7962]), .Z(n5440) );
  XOR U13496 ( .A(n5434), .B(n5433), .Z(n5444) );
  XOR U13497 ( .A(n5436), .B(n5435), .Z(n5433) );
  XOR U13498 ( .A(y[7961]), .B(x[7961]), .Z(n5435) );
  XOR U13499 ( .A(y[7960]), .B(x[7960]), .Z(n5436) );
  XOR U13500 ( .A(y[7959]), .B(x[7959]), .Z(n5434) );
  NAND U13501 ( .A(n5497), .B(n5498), .Z(N64899) );
  NAND U13502 ( .A(n5499), .B(n5500), .Z(n5498) );
  NANDN U13503 ( .A(n5501), .B(n5502), .Z(n5500) );
  NANDN U13504 ( .A(n5502), .B(n5501), .Z(n5497) );
  XOR U13505 ( .A(n5501), .B(n5503), .Z(N64898) );
  XNOR U13506 ( .A(n5499), .B(n5502), .Z(n5503) );
  NAND U13507 ( .A(n5504), .B(n5505), .Z(n5502) );
  NAND U13508 ( .A(n5506), .B(n5507), .Z(n5505) );
  NANDN U13509 ( .A(n5508), .B(n5509), .Z(n5507) );
  NANDN U13510 ( .A(n5509), .B(n5508), .Z(n5504) );
  AND U13511 ( .A(n5510), .B(n5511), .Z(n5499) );
  NAND U13512 ( .A(n5512), .B(n5513), .Z(n5511) );
  NANDN U13513 ( .A(n5514), .B(n5515), .Z(n5513) );
  NANDN U13514 ( .A(n5515), .B(n5514), .Z(n5510) );
  IV U13515 ( .A(n5516), .Z(n5515) );
  AND U13516 ( .A(n5517), .B(n5518), .Z(n5501) );
  NAND U13517 ( .A(n5519), .B(n5520), .Z(n5518) );
  NANDN U13518 ( .A(n5521), .B(n5522), .Z(n5520) );
  NANDN U13519 ( .A(n5522), .B(n5521), .Z(n5517) );
  XOR U13520 ( .A(n5514), .B(n5523), .Z(N64897) );
  XNOR U13521 ( .A(n5512), .B(n5516), .Z(n5523) );
  XOR U13522 ( .A(n5509), .B(n5524), .Z(n5516) );
  XNOR U13523 ( .A(n5506), .B(n5508), .Z(n5524) );
  AND U13524 ( .A(n5525), .B(n5526), .Z(n5508) );
  NANDN U13525 ( .A(n5527), .B(n5528), .Z(n5526) );
  OR U13526 ( .A(n5529), .B(n5530), .Z(n5528) );
  IV U13527 ( .A(n5531), .Z(n5530) );
  NANDN U13528 ( .A(n5531), .B(n5529), .Z(n5525) );
  AND U13529 ( .A(n5532), .B(n5533), .Z(n5506) );
  NAND U13530 ( .A(n5534), .B(n5535), .Z(n5533) );
  NANDN U13531 ( .A(n5536), .B(n5537), .Z(n5535) );
  NANDN U13532 ( .A(n5537), .B(n5536), .Z(n5532) );
  IV U13533 ( .A(n5538), .Z(n5537) );
  NAND U13534 ( .A(n5539), .B(n5540), .Z(n5509) );
  NANDN U13535 ( .A(n5541), .B(n5542), .Z(n5540) );
  NANDN U13536 ( .A(n5543), .B(n5544), .Z(n5542) );
  NANDN U13537 ( .A(n5544), .B(n5543), .Z(n5539) );
  IV U13538 ( .A(n5545), .Z(n5543) );
  AND U13539 ( .A(n5546), .B(n5547), .Z(n5512) );
  NAND U13540 ( .A(n5548), .B(n5549), .Z(n5547) );
  NANDN U13541 ( .A(n5550), .B(n5551), .Z(n5549) );
  NANDN U13542 ( .A(n5551), .B(n5550), .Z(n5546) );
  XOR U13543 ( .A(n5522), .B(n5552), .Z(n5514) );
  XNOR U13544 ( .A(n5519), .B(n5521), .Z(n5552) );
  AND U13545 ( .A(n5553), .B(n5554), .Z(n5521) );
  NANDN U13546 ( .A(n5555), .B(n5556), .Z(n5554) );
  OR U13547 ( .A(n5557), .B(n5558), .Z(n5556) );
  IV U13548 ( .A(n5559), .Z(n5558) );
  NANDN U13549 ( .A(n5559), .B(n5557), .Z(n5553) );
  AND U13550 ( .A(n5560), .B(n5561), .Z(n5519) );
  NAND U13551 ( .A(n5562), .B(n5563), .Z(n5561) );
  NANDN U13552 ( .A(n5564), .B(n5565), .Z(n5563) );
  NANDN U13553 ( .A(n5565), .B(n5564), .Z(n5560) );
  IV U13554 ( .A(n5566), .Z(n5565) );
  NAND U13555 ( .A(n5567), .B(n5568), .Z(n5522) );
  NANDN U13556 ( .A(n5569), .B(n5570), .Z(n5568) );
  NANDN U13557 ( .A(n5571), .B(n5572), .Z(n5570) );
  NANDN U13558 ( .A(n5572), .B(n5571), .Z(n5567) );
  IV U13559 ( .A(n5573), .Z(n5571) );
  XOR U13560 ( .A(n5548), .B(n5574), .Z(N64896) );
  XNOR U13561 ( .A(n5551), .B(n5550), .Z(n5574) );
  XNOR U13562 ( .A(n5562), .B(n5575), .Z(n5550) );
  XNOR U13563 ( .A(n5566), .B(n5564), .Z(n5575) );
  XOR U13564 ( .A(n5572), .B(n5576), .Z(n5564) );
  XNOR U13565 ( .A(n5569), .B(n5573), .Z(n5576) );
  AND U13566 ( .A(n5577), .B(n5578), .Z(n5573) );
  NAND U13567 ( .A(n5579), .B(n5580), .Z(n5578) );
  NAND U13568 ( .A(n5581), .B(n5582), .Z(n5577) );
  AND U13569 ( .A(n5583), .B(n5584), .Z(n5569) );
  NAND U13570 ( .A(n5585), .B(n5586), .Z(n5584) );
  NAND U13571 ( .A(n5587), .B(n5588), .Z(n5583) );
  NANDN U13572 ( .A(n5589), .B(n5590), .Z(n5572) );
  ANDN U13573 ( .B(n5591), .A(n5592), .Z(n5566) );
  XNOR U13574 ( .A(n5557), .B(n5593), .Z(n5562) );
  XNOR U13575 ( .A(n5555), .B(n5559), .Z(n5593) );
  AND U13576 ( .A(n5594), .B(n5595), .Z(n5559) );
  NAND U13577 ( .A(n5596), .B(n5597), .Z(n5595) );
  NAND U13578 ( .A(n5598), .B(n5599), .Z(n5594) );
  AND U13579 ( .A(n5600), .B(n5601), .Z(n5555) );
  NAND U13580 ( .A(n5602), .B(n5603), .Z(n5601) );
  NAND U13581 ( .A(n5604), .B(n5605), .Z(n5600) );
  AND U13582 ( .A(n5606), .B(n5607), .Z(n5557) );
  NAND U13583 ( .A(n5608), .B(n5609), .Z(n5551) );
  XNOR U13584 ( .A(n5534), .B(n5610), .Z(n5548) );
  XNOR U13585 ( .A(n5538), .B(n5536), .Z(n5610) );
  XOR U13586 ( .A(n5544), .B(n5611), .Z(n5536) );
  XNOR U13587 ( .A(n5541), .B(n5545), .Z(n5611) );
  AND U13588 ( .A(n5612), .B(n5613), .Z(n5545) );
  NAND U13589 ( .A(n5614), .B(n5615), .Z(n5613) );
  NAND U13590 ( .A(n5616), .B(n5617), .Z(n5612) );
  AND U13591 ( .A(n5618), .B(n5619), .Z(n5541) );
  NAND U13592 ( .A(n5620), .B(n5621), .Z(n5619) );
  NAND U13593 ( .A(n5622), .B(n5623), .Z(n5618) );
  NANDN U13594 ( .A(n5624), .B(n5625), .Z(n5544) );
  ANDN U13595 ( .B(n5626), .A(n5627), .Z(n5538) );
  XNOR U13596 ( .A(n5529), .B(n5628), .Z(n5534) );
  XNOR U13597 ( .A(n5527), .B(n5531), .Z(n5628) );
  AND U13598 ( .A(n5629), .B(n5630), .Z(n5531) );
  NAND U13599 ( .A(n5631), .B(n5632), .Z(n5630) );
  NAND U13600 ( .A(n5633), .B(n5634), .Z(n5629) );
  AND U13601 ( .A(n5635), .B(n5636), .Z(n5527) );
  NAND U13602 ( .A(n5637), .B(n5638), .Z(n5636) );
  NAND U13603 ( .A(n5639), .B(n5640), .Z(n5635) );
  AND U13604 ( .A(n5641), .B(n5642), .Z(n5529) );
  XOR U13605 ( .A(n5609), .B(n5608), .Z(N64895) );
  XNOR U13606 ( .A(n5626), .B(n5627), .Z(n5608) );
  XNOR U13607 ( .A(n5641), .B(n5642), .Z(n5627) );
  XOR U13608 ( .A(n5638), .B(n5637), .Z(n5642) );
  XOR U13609 ( .A(y[7956]), .B(x[7956]), .Z(n5637) );
  XOR U13610 ( .A(n5640), .B(n5639), .Z(n5638) );
  XOR U13611 ( .A(y[7958]), .B(x[7958]), .Z(n5639) );
  XOR U13612 ( .A(y[7957]), .B(x[7957]), .Z(n5640) );
  XOR U13613 ( .A(n5632), .B(n5631), .Z(n5641) );
  XOR U13614 ( .A(n5634), .B(n5633), .Z(n5631) );
  XOR U13615 ( .A(y[7955]), .B(x[7955]), .Z(n5633) );
  XOR U13616 ( .A(y[7954]), .B(x[7954]), .Z(n5634) );
  XOR U13617 ( .A(y[7953]), .B(x[7953]), .Z(n5632) );
  XNOR U13618 ( .A(n5625), .B(n5624), .Z(n5626) );
  XNOR U13619 ( .A(n5621), .B(n5620), .Z(n5624) );
  XOR U13620 ( .A(n5623), .B(n5622), .Z(n5620) );
  XOR U13621 ( .A(y[7952]), .B(x[7952]), .Z(n5622) );
  XOR U13622 ( .A(y[7951]), .B(x[7951]), .Z(n5623) );
  XOR U13623 ( .A(y[7950]), .B(x[7950]), .Z(n5621) );
  XOR U13624 ( .A(n5615), .B(n5614), .Z(n5625) );
  XOR U13625 ( .A(n5617), .B(n5616), .Z(n5614) );
  XOR U13626 ( .A(y[7949]), .B(x[7949]), .Z(n5616) );
  XOR U13627 ( .A(y[7948]), .B(x[7948]), .Z(n5617) );
  XOR U13628 ( .A(y[7947]), .B(x[7947]), .Z(n5615) );
  XNOR U13629 ( .A(n5591), .B(n5592), .Z(n5609) );
  XNOR U13630 ( .A(n5606), .B(n5607), .Z(n5592) );
  XOR U13631 ( .A(n5603), .B(n5602), .Z(n5607) );
  XOR U13632 ( .A(y[7944]), .B(x[7944]), .Z(n5602) );
  XOR U13633 ( .A(n5605), .B(n5604), .Z(n5603) );
  XOR U13634 ( .A(y[7946]), .B(x[7946]), .Z(n5604) );
  XOR U13635 ( .A(y[7945]), .B(x[7945]), .Z(n5605) );
  XOR U13636 ( .A(n5597), .B(n5596), .Z(n5606) );
  XOR U13637 ( .A(n5599), .B(n5598), .Z(n5596) );
  XOR U13638 ( .A(y[7943]), .B(x[7943]), .Z(n5598) );
  XOR U13639 ( .A(y[7942]), .B(x[7942]), .Z(n5599) );
  XOR U13640 ( .A(y[7941]), .B(x[7941]), .Z(n5597) );
  XNOR U13641 ( .A(n5590), .B(n5589), .Z(n5591) );
  XNOR U13642 ( .A(n5586), .B(n5585), .Z(n5589) );
  XOR U13643 ( .A(n5588), .B(n5587), .Z(n5585) );
  XOR U13644 ( .A(y[7940]), .B(x[7940]), .Z(n5587) );
  XOR U13645 ( .A(y[7939]), .B(x[7939]), .Z(n5588) );
  XOR U13646 ( .A(y[7938]), .B(x[7938]), .Z(n5586) );
  XOR U13647 ( .A(n5580), .B(n5579), .Z(n5590) );
  XOR U13648 ( .A(n5582), .B(n5581), .Z(n5579) );
  XOR U13649 ( .A(y[7937]), .B(x[7937]), .Z(n5581) );
  XOR U13650 ( .A(y[7936]), .B(x[7936]), .Z(n5582) );
  XOR U13651 ( .A(y[7935]), .B(x[7935]), .Z(n5580) );
  NAND U13652 ( .A(n5643), .B(n5644), .Z(N64886) );
  NAND U13653 ( .A(n5645), .B(n5646), .Z(n5644) );
  NANDN U13654 ( .A(n5647), .B(n5648), .Z(n5646) );
  NANDN U13655 ( .A(n5648), .B(n5647), .Z(n5643) );
  XOR U13656 ( .A(n5647), .B(n5649), .Z(N64885) );
  XNOR U13657 ( .A(n5645), .B(n5648), .Z(n5649) );
  NAND U13658 ( .A(n5650), .B(n5651), .Z(n5648) );
  NAND U13659 ( .A(n5652), .B(n5653), .Z(n5651) );
  NANDN U13660 ( .A(n5654), .B(n5655), .Z(n5653) );
  NANDN U13661 ( .A(n5655), .B(n5654), .Z(n5650) );
  AND U13662 ( .A(n5656), .B(n5657), .Z(n5645) );
  NAND U13663 ( .A(n5658), .B(n5659), .Z(n5657) );
  NANDN U13664 ( .A(n5660), .B(n5661), .Z(n5659) );
  NANDN U13665 ( .A(n5661), .B(n5660), .Z(n5656) );
  IV U13666 ( .A(n5662), .Z(n5661) );
  AND U13667 ( .A(n5663), .B(n5664), .Z(n5647) );
  NAND U13668 ( .A(n5665), .B(n5666), .Z(n5664) );
  NANDN U13669 ( .A(n5667), .B(n5668), .Z(n5666) );
  NANDN U13670 ( .A(n5668), .B(n5667), .Z(n5663) );
  XOR U13671 ( .A(n5660), .B(n5669), .Z(N64884) );
  XNOR U13672 ( .A(n5658), .B(n5662), .Z(n5669) );
  XOR U13673 ( .A(n5655), .B(n5670), .Z(n5662) );
  XNOR U13674 ( .A(n5652), .B(n5654), .Z(n5670) );
  AND U13675 ( .A(n5671), .B(n5672), .Z(n5654) );
  NANDN U13676 ( .A(n5673), .B(n5674), .Z(n5672) );
  OR U13677 ( .A(n5675), .B(n5676), .Z(n5674) );
  IV U13678 ( .A(n5677), .Z(n5676) );
  NANDN U13679 ( .A(n5677), .B(n5675), .Z(n5671) );
  AND U13680 ( .A(n5678), .B(n5679), .Z(n5652) );
  NAND U13681 ( .A(n5680), .B(n5681), .Z(n5679) );
  NANDN U13682 ( .A(n5682), .B(n5683), .Z(n5681) );
  NANDN U13683 ( .A(n5683), .B(n5682), .Z(n5678) );
  IV U13684 ( .A(n5684), .Z(n5683) );
  NAND U13685 ( .A(n5685), .B(n5686), .Z(n5655) );
  NANDN U13686 ( .A(n5687), .B(n5688), .Z(n5686) );
  NANDN U13687 ( .A(n5689), .B(n5690), .Z(n5688) );
  NANDN U13688 ( .A(n5690), .B(n5689), .Z(n5685) );
  IV U13689 ( .A(n5691), .Z(n5689) );
  AND U13690 ( .A(n5692), .B(n5693), .Z(n5658) );
  NAND U13691 ( .A(n5694), .B(n5695), .Z(n5693) );
  NANDN U13692 ( .A(n5696), .B(n5697), .Z(n5695) );
  NANDN U13693 ( .A(n5697), .B(n5696), .Z(n5692) );
  XOR U13694 ( .A(n5668), .B(n5698), .Z(n5660) );
  XNOR U13695 ( .A(n5665), .B(n5667), .Z(n5698) );
  AND U13696 ( .A(n5699), .B(n5700), .Z(n5667) );
  NANDN U13697 ( .A(n5701), .B(n5702), .Z(n5700) );
  OR U13698 ( .A(n5703), .B(n5704), .Z(n5702) );
  IV U13699 ( .A(n5705), .Z(n5704) );
  NANDN U13700 ( .A(n5705), .B(n5703), .Z(n5699) );
  AND U13701 ( .A(n5706), .B(n5707), .Z(n5665) );
  NAND U13702 ( .A(n5708), .B(n5709), .Z(n5707) );
  NANDN U13703 ( .A(n5710), .B(n5711), .Z(n5709) );
  NANDN U13704 ( .A(n5711), .B(n5710), .Z(n5706) );
  IV U13705 ( .A(n5712), .Z(n5711) );
  NAND U13706 ( .A(n5713), .B(n5714), .Z(n5668) );
  NANDN U13707 ( .A(n5715), .B(n5716), .Z(n5714) );
  NANDN U13708 ( .A(n5717), .B(n5718), .Z(n5716) );
  NANDN U13709 ( .A(n5718), .B(n5717), .Z(n5713) );
  IV U13710 ( .A(n5719), .Z(n5717) );
  XOR U13711 ( .A(n5694), .B(n5720), .Z(N64883) );
  XNOR U13712 ( .A(n5697), .B(n5696), .Z(n5720) );
  XNOR U13713 ( .A(n5708), .B(n5721), .Z(n5696) );
  XNOR U13714 ( .A(n5712), .B(n5710), .Z(n5721) );
  XOR U13715 ( .A(n5718), .B(n5722), .Z(n5710) );
  XNOR U13716 ( .A(n5715), .B(n5719), .Z(n5722) );
  AND U13717 ( .A(n5723), .B(n5724), .Z(n5719) );
  NAND U13718 ( .A(n5725), .B(n5726), .Z(n5724) );
  NAND U13719 ( .A(n5727), .B(n5728), .Z(n5723) );
  AND U13720 ( .A(n5729), .B(n5730), .Z(n5715) );
  NAND U13721 ( .A(n5731), .B(n5732), .Z(n5730) );
  NAND U13722 ( .A(n5733), .B(n5734), .Z(n5729) );
  NANDN U13723 ( .A(n5735), .B(n5736), .Z(n5718) );
  ANDN U13724 ( .B(n5737), .A(n5738), .Z(n5712) );
  XNOR U13725 ( .A(n5703), .B(n5739), .Z(n5708) );
  XNOR U13726 ( .A(n5701), .B(n5705), .Z(n5739) );
  AND U13727 ( .A(n5740), .B(n5741), .Z(n5705) );
  NAND U13728 ( .A(n5742), .B(n5743), .Z(n5741) );
  NAND U13729 ( .A(n5744), .B(n5745), .Z(n5740) );
  AND U13730 ( .A(n5746), .B(n5747), .Z(n5701) );
  NAND U13731 ( .A(n5748), .B(n5749), .Z(n5747) );
  NAND U13732 ( .A(n5750), .B(n5751), .Z(n5746) );
  AND U13733 ( .A(n5752), .B(n5753), .Z(n5703) );
  NAND U13734 ( .A(n5754), .B(n5755), .Z(n5697) );
  XNOR U13735 ( .A(n5680), .B(n5756), .Z(n5694) );
  XNOR U13736 ( .A(n5684), .B(n5682), .Z(n5756) );
  XOR U13737 ( .A(n5690), .B(n5757), .Z(n5682) );
  XNOR U13738 ( .A(n5687), .B(n5691), .Z(n5757) );
  AND U13739 ( .A(n5758), .B(n5759), .Z(n5691) );
  NAND U13740 ( .A(n5760), .B(n5761), .Z(n5759) );
  NAND U13741 ( .A(n5762), .B(n5763), .Z(n5758) );
  AND U13742 ( .A(n5764), .B(n5765), .Z(n5687) );
  NAND U13743 ( .A(n5766), .B(n5767), .Z(n5765) );
  NAND U13744 ( .A(n5768), .B(n5769), .Z(n5764) );
  NANDN U13745 ( .A(n5770), .B(n5771), .Z(n5690) );
  ANDN U13746 ( .B(n5772), .A(n5773), .Z(n5684) );
  XNOR U13747 ( .A(n5675), .B(n5774), .Z(n5680) );
  XNOR U13748 ( .A(n5673), .B(n5677), .Z(n5774) );
  AND U13749 ( .A(n5775), .B(n5776), .Z(n5677) );
  NAND U13750 ( .A(n5777), .B(n5778), .Z(n5776) );
  NAND U13751 ( .A(n5779), .B(n5780), .Z(n5775) );
  AND U13752 ( .A(n5781), .B(n5782), .Z(n5673) );
  NAND U13753 ( .A(n5783), .B(n5784), .Z(n5782) );
  NAND U13754 ( .A(n5785), .B(n5786), .Z(n5781) );
  AND U13755 ( .A(n5787), .B(n5788), .Z(n5675) );
  XOR U13756 ( .A(n5755), .B(n5754), .Z(N64882) );
  XNOR U13757 ( .A(n5772), .B(n5773), .Z(n5754) );
  XNOR U13758 ( .A(n5787), .B(n5788), .Z(n5773) );
  XOR U13759 ( .A(n5784), .B(n5783), .Z(n5788) );
  XOR U13760 ( .A(y[7932]), .B(x[7932]), .Z(n5783) );
  XOR U13761 ( .A(n5786), .B(n5785), .Z(n5784) );
  XOR U13762 ( .A(y[7934]), .B(x[7934]), .Z(n5785) );
  XOR U13763 ( .A(y[7933]), .B(x[7933]), .Z(n5786) );
  XOR U13764 ( .A(n5778), .B(n5777), .Z(n5787) );
  XOR U13765 ( .A(n5780), .B(n5779), .Z(n5777) );
  XOR U13766 ( .A(y[7931]), .B(x[7931]), .Z(n5779) );
  XOR U13767 ( .A(y[7930]), .B(x[7930]), .Z(n5780) );
  XOR U13768 ( .A(y[7929]), .B(x[7929]), .Z(n5778) );
  XNOR U13769 ( .A(n5771), .B(n5770), .Z(n5772) );
  XNOR U13770 ( .A(n5767), .B(n5766), .Z(n5770) );
  XOR U13771 ( .A(n5769), .B(n5768), .Z(n5766) );
  XOR U13772 ( .A(y[7928]), .B(x[7928]), .Z(n5768) );
  XOR U13773 ( .A(y[7927]), .B(x[7927]), .Z(n5769) );
  XOR U13774 ( .A(y[7926]), .B(x[7926]), .Z(n5767) );
  XOR U13775 ( .A(n5761), .B(n5760), .Z(n5771) );
  XOR U13776 ( .A(n5763), .B(n5762), .Z(n5760) );
  XOR U13777 ( .A(y[7925]), .B(x[7925]), .Z(n5762) );
  XOR U13778 ( .A(y[7924]), .B(x[7924]), .Z(n5763) );
  XOR U13779 ( .A(y[7923]), .B(x[7923]), .Z(n5761) );
  XNOR U13780 ( .A(n5737), .B(n5738), .Z(n5755) );
  XNOR U13781 ( .A(n5752), .B(n5753), .Z(n5738) );
  XOR U13782 ( .A(n5749), .B(n5748), .Z(n5753) );
  XOR U13783 ( .A(y[7920]), .B(x[7920]), .Z(n5748) );
  XOR U13784 ( .A(n5751), .B(n5750), .Z(n5749) );
  XOR U13785 ( .A(y[7922]), .B(x[7922]), .Z(n5750) );
  XOR U13786 ( .A(y[7921]), .B(x[7921]), .Z(n5751) );
  XOR U13787 ( .A(n5743), .B(n5742), .Z(n5752) );
  XOR U13788 ( .A(n5745), .B(n5744), .Z(n5742) );
  XOR U13789 ( .A(y[7919]), .B(x[7919]), .Z(n5744) );
  XOR U13790 ( .A(y[7918]), .B(x[7918]), .Z(n5745) );
  XOR U13791 ( .A(y[7917]), .B(x[7917]), .Z(n5743) );
  XNOR U13792 ( .A(n5736), .B(n5735), .Z(n5737) );
  XNOR U13793 ( .A(n5732), .B(n5731), .Z(n5735) );
  XOR U13794 ( .A(n5734), .B(n5733), .Z(n5731) );
  XOR U13795 ( .A(y[7916]), .B(x[7916]), .Z(n5733) );
  XOR U13796 ( .A(y[7915]), .B(x[7915]), .Z(n5734) );
  XOR U13797 ( .A(y[7914]), .B(x[7914]), .Z(n5732) );
  XOR U13798 ( .A(n5726), .B(n5725), .Z(n5736) );
  XOR U13799 ( .A(n5728), .B(n5727), .Z(n5725) );
  XOR U13800 ( .A(y[7913]), .B(x[7913]), .Z(n5727) );
  XOR U13801 ( .A(y[7912]), .B(x[7912]), .Z(n5728) );
  XOR U13802 ( .A(y[7911]), .B(x[7911]), .Z(n5726) );
  NAND U13803 ( .A(n5789), .B(n5790), .Z(N64873) );
  NAND U13804 ( .A(n5791), .B(n5792), .Z(n5790) );
  NANDN U13805 ( .A(n5793), .B(n5794), .Z(n5792) );
  NANDN U13806 ( .A(n5794), .B(n5793), .Z(n5789) );
  XOR U13807 ( .A(n5793), .B(n5795), .Z(N64872) );
  XNOR U13808 ( .A(n5791), .B(n5794), .Z(n5795) );
  NAND U13809 ( .A(n5796), .B(n5797), .Z(n5794) );
  NAND U13810 ( .A(n5798), .B(n5799), .Z(n5797) );
  NANDN U13811 ( .A(n5800), .B(n5801), .Z(n5799) );
  NANDN U13812 ( .A(n5801), .B(n5800), .Z(n5796) );
  AND U13813 ( .A(n5802), .B(n5803), .Z(n5791) );
  NAND U13814 ( .A(n5804), .B(n5805), .Z(n5803) );
  NANDN U13815 ( .A(n5806), .B(n5807), .Z(n5805) );
  NANDN U13816 ( .A(n5807), .B(n5806), .Z(n5802) );
  IV U13817 ( .A(n5808), .Z(n5807) );
  AND U13818 ( .A(n5809), .B(n5810), .Z(n5793) );
  NAND U13819 ( .A(n5811), .B(n5812), .Z(n5810) );
  NANDN U13820 ( .A(n5813), .B(n5814), .Z(n5812) );
  NANDN U13821 ( .A(n5814), .B(n5813), .Z(n5809) );
  XOR U13822 ( .A(n5806), .B(n5815), .Z(N64871) );
  XNOR U13823 ( .A(n5804), .B(n5808), .Z(n5815) );
  XOR U13824 ( .A(n5801), .B(n5816), .Z(n5808) );
  XNOR U13825 ( .A(n5798), .B(n5800), .Z(n5816) );
  AND U13826 ( .A(n5817), .B(n5818), .Z(n5800) );
  NANDN U13827 ( .A(n5819), .B(n5820), .Z(n5818) );
  OR U13828 ( .A(n5821), .B(n5822), .Z(n5820) );
  IV U13829 ( .A(n5823), .Z(n5822) );
  NANDN U13830 ( .A(n5823), .B(n5821), .Z(n5817) );
  AND U13831 ( .A(n5824), .B(n5825), .Z(n5798) );
  NAND U13832 ( .A(n5826), .B(n5827), .Z(n5825) );
  NANDN U13833 ( .A(n5828), .B(n5829), .Z(n5827) );
  NANDN U13834 ( .A(n5829), .B(n5828), .Z(n5824) );
  IV U13835 ( .A(n5830), .Z(n5829) );
  NAND U13836 ( .A(n5831), .B(n5832), .Z(n5801) );
  NANDN U13837 ( .A(n5833), .B(n5834), .Z(n5832) );
  NANDN U13838 ( .A(n5835), .B(n5836), .Z(n5834) );
  NANDN U13839 ( .A(n5836), .B(n5835), .Z(n5831) );
  IV U13840 ( .A(n5837), .Z(n5835) );
  AND U13841 ( .A(n5838), .B(n5839), .Z(n5804) );
  NAND U13842 ( .A(n5840), .B(n5841), .Z(n5839) );
  NANDN U13843 ( .A(n5842), .B(n5843), .Z(n5841) );
  NANDN U13844 ( .A(n5843), .B(n5842), .Z(n5838) );
  XOR U13845 ( .A(n5814), .B(n5844), .Z(n5806) );
  XNOR U13846 ( .A(n5811), .B(n5813), .Z(n5844) );
  AND U13847 ( .A(n5845), .B(n5846), .Z(n5813) );
  NANDN U13848 ( .A(n5847), .B(n5848), .Z(n5846) );
  OR U13849 ( .A(n5849), .B(n5850), .Z(n5848) );
  IV U13850 ( .A(n5851), .Z(n5850) );
  NANDN U13851 ( .A(n5851), .B(n5849), .Z(n5845) );
  AND U13852 ( .A(n5852), .B(n5853), .Z(n5811) );
  NAND U13853 ( .A(n5854), .B(n5855), .Z(n5853) );
  NANDN U13854 ( .A(n5856), .B(n5857), .Z(n5855) );
  NANDN U13855 ( .A(n5857), .B(n5856), .Z(n5852) );
  IV U13856 ( .A(n5858), .Z(n5857) );
  NAND U13857 ( .A(n5859), .B(n5860), .Z(n5814) );
  NANDN U13858 ( .A(n5861), .B(n5862), .Z(n5860) );
  NANDN U13859 ( .A(n5863), .B(n5864), .Z(n5862) );
  NANDN U13860 ( .A(n5864), .B(n5863), .Z(n5859) );
  IV U13861 ( .A(n5865), .Z(n5863) );
  XOR U13862 ( .A(n5840), .B(n5866), .Z(N64870) );
  XNOR U13863 ( .A(n5843), .B(n5842), .Z(n5866) );
  XNOR U13864 ( .A(n5854), .B(n5867), .Z(n5842) );
  XNOR U13865 ( .A(n5858), .B(n5856), .Z(n5867) );
  XOR U13866 ( .A(n5864), .B(n5868), .Z(n5856) );
  XNOR U13867 ( .A(n5861), .B(n5865), .Z(n5868) );
  AND U13868 ( .A(n5869), .B(n5870), .Z(n5865) );
  NAND U13869 ( .A(n5871), .B(n5872), .Z(n5870) );
  NAND U13870 ( .A(n5873), .B(n5874), .Z(n5869) );
  AND U13871 ( .A(n5875), .B(n5876), .Z(n5861) );
  NAND U13872 ( .A(n5877), .B(n5878), .Z(n5876) );
  NAND U13873 ( .A(n5879), .B(n5880), .Z(n5875) );
  NANDN U13874 ( .A(n5881), .B(n5882), .Z(n5864) );
  ANDN U13875 ( .B(n5883), .A(n5884), .Z(n5858) );
  XNOR U13876 ( .A(n5849), .B(n5885), .Z(n5854) );
  XNOR U13877 ( .A(n5847), .B(n5851), .Z(n5885) );
  AND U13878 ( .A(n5886), .B(n5887), .Z(n5851) );
  NAND U13879 ( .A(n5888), .B(n5889), .Z(n5887) );
  NAND U13880 ( .A(n5890), .B(n5891), .Z(n5886) );
  AND U13881 ( .A(n5892), .B(n5893), .Z(n5847) );
  NAND U13882 ( .A(n5894), .B(n5895), .Z(n5893) );
  NAND U13883 ( .A(n5896), .B(n5897), .Z(n5892) );
  AND U13884 ( .A(n5898), .B(n5899), .Z(n5849) );
  NAND U13885 ( .A(n5900), .B(n5901), .Z(n5843) );
  XNOR U13886 ( .A(n5826), .B(n5902), .Z(n5840) );
  XNOR U13887 ( .A(n5830), .B(n5828), .Z(n5902) );
  XOR U13888 ( .A(n5836), .B(n5903), .Z(n5828) );
  XNOR U13889 ( .A(n5833), .B(n5837), .Z(n5903) );
  AND U13890 ( .A(n5904), .B(n5905), .Z(n5837) );
  NAND U13891 ( .A(n5906), .B(n5907), .Z(n5905) );
  NAND U13892 ( .A(n5908), .B(n5909), .Z(n5904) );
  AND U13893 ( .A(n5910), .B(n5911), .Z(n5833) );
  NAND U13894 ( .A(n5912), .B(n5913), .Z(n5911) );
  NAND U13895 ( .A(n5914), .B(n5915), .Z(n5910) );
  NANDN U13896 ( .A(n5916), .B(n5917), .Z(n5836) );
  ANDN U13897 ( .B(n5918), .A(n5919), .Z(n5830) );
  XNOR U13898 ( .A(n5821), .B(n5920), .Z(n5826) );
  XNOR U13899 ( .A(n5819), .B(n5823), .Z(n5920) );
  AND U13900 ( .A(n5921), .B(n5922), .Z(n5823) );
  NAND U13901 ( .A(n5923), .B(n5924), .Z(n5922) );
  NAND U13902 ( .A(n5925), .B(n5926), .Z(n5921) );
  AND U13903 ( .A(n5927), .B(n5928), .Z(n5819) );
  NAND U13904 ( .A(n5929), .B(n5930), .Z(n5928) );
  NAND U13905 ( .A(n5931), .B(n5932), .Z(n5927) );
  AND U13906 ( .A(n5933), .B(n5934), .Z(n5821) );
  XOR U13907 ( .A(n5901), .B(n5900), .Z(N64869) );
  XNOR U13908 ( .A(n5918), .B(n5919), .Z(n5900) );
  XNOR U13909 ( .A(n5933), .B(n5934), .Z(n5919) );
  XOR U13910 ( .A(n5930), .B(n5929), .Z(n5934) );
  XOR U13911 ( .A(y[7908]), .B(x[7908]), .Z(n5929) );
  XOR U13912 ( .A(n5932), .B(n5931), .Z(n5930) );
  XOR U13913 ( .A(y[7910]), .B(x[7910]), .Z(n5931) );
  XOR U13914 ( .A(y[7909]), .B(x[7909]), .Z(n5932) );
  XOR U13915 ( .A(n5924), .B(n5923), .Z(n5933) );
  XOR U13916 ( .A(n5926), .B(n5925), .Z(n5923) );
  XOR U13917 ( .A(y[7907]), .B(x[7907]), .Z(n5925) );
  XOR U13918 ( .A(y[7906]), .B(x[7906]), .Z(n5926) );
  XOR U13919 ( .A(y[7905]), .B(x[7905]), .Z(n5924) );
  XNOR U13920 ( .A(n5917), .B(n5916), .Z(n5918) );
  XNOR U13921 ( .A(n5913), .B(n5912), .Z(n5916) );
  XOR U13922 ( .A(n5915), .B(n5914), .Z(n5912) );
  XOR U13923 ( .A(y[7904]), .B(x[7904]), .Z(n5914) );
  XOR U13924 ( .A(y[7903]), .B(x[7903]), .Z(n5915) );
  XOR U13925 ( .A(y[7902]), .B(x[7902]), .Z(n5913) );
  XOR U13926 ( .A(n5907), .B(n5906), .Z(n5917) );
  XOR U13927 ( .A(n5909), .B(n5908), .Z(n5906) );
  XOR U13928 ( .A(y[7901]), .B(x[7901]), .Z(n5908) );
  XOR U13929 ( .A(y[7900]), .B(x[7900]), .Z(n5909) );
  XOR U13930 ( .A(y[7899]), .B(x[7899]), .Z(n5907) );
  XNOR U13931 ( .A(n5883), .B(n5884), .Z(n5901) );
  XNOR U13932 ( .A(n5898), .B(n5899), .Z(n5884) );
  XOR U13933 ( .A(n5895), .B(n5894), .Z(n5899) );
  XOR U13934 ( .A(y[7896]), .B(x[7896]), .Z(n5894) );
  XOR U13935 ( .A(n5897), .B(n5896), .Z(n5895) );
  XOR U13936 ( .A(y[7898]), .B(x[7898]), .Z(n5896) );
  XOR U13937 ( .A(y[7897]), .B(x[7897]), .Z(n5897) );
  XOR U13938 ( .A(n5889), .B(n5888), .Z(n5898) );
  XOR U13939 ( .A(n5891), .B(n5890), .Z(n5888) );
  XOR U13940 ( .A(y[7895]), .B(x[7895]), .Z(n5890) );
  XOR U13941 ( .A(y[7894]), .B(x[7894]), .Z(n5891) );
  XOR U13942 ( .A(y[7893]), .B(x[7893]), .Z(n5889) );
  XNOR U13943 ( .A(n5882), .B(n5881), .Z(n5883) );
  XNOR U13944 ( .A(n5878), .B(n5877), .Z(n5881) );
  XOR U13945 ( .A(n5880), .B(n5879), .Z(n5877) );
  XOR U13946 ( .A(y[7892]), .B(x[7892]), .Z(n5879) );
  XOR U13947 ( .A(y[7891]), .B(x[7891]), .Z(n5880) );
  XOR U13948 ( .A(y[7890]), .B(x[7890]), .Z(n5878) );
  XOR U13949 ( .A(n5872), .B(n5871), .Z(n5882) );
  XOR U13950 ( .A(n5874), .B(n5873), .Z(n5871) );
  XOR U13951 ( .A(y[7889]), .B(x[7889]), .Z(n5873) );
  XOR U13952 ( .A(y[7888]), .B(x[7888]), .Z(n5874) );
  XOR U13953 ( .A(y[7887]), .B(x[7887]), .Z(n5872) );
  NAND U13954 ( .A(n5935), .B(n5936), .Z(N64860) );
  NAND U13955 ( .A(n5937), .B(n5938), .Z(n5936) );
  NANDN U13956 ( .A(n5939), .B(n5940), .Z(n5938) );
  NANDN U13957 ( .A(n5940), .B(n5939), .Z(n5935) );
  XOR U13958 ( .A(n5939), .B(n5941), .Z(N64859) );
  XNOR U13959 ( .A(n5937), .B(n5940), .Z(n5941) );
  NAND U13960 ( .A(n5942), .B(n5943), .Z(n5940) );
  NAND U13961 ( .A(n5944), .B(n5945), .Z(n5943) );
  NANDN U13962 ( .A(n5946), .B(n5947), .Z(n5945) );
  NANDN U13963 ( .A(n5947), .B(n5946), .Z(n5942) );
  AND U13964 ( .A(n5948), .B(n5949), .Z(n5937) );
  NAND U13965 ( .A(n5950), .B(n5951), .Z(n5949) );
  NANDN U13966 ( .A(n5952), .B(n5953), .Z(n5951) );
  NANDN U13967 ( .A(n5953), .B(n5952), .Z(n5948) );
  IV U13968 ( .A(n5954), .Z(n5953) );
  AND U13969 ( .A(n5955), .B(n5956), .Z(n5939) );
  NAND U13970 ( .A(n5957), .B(n5958), .Z(n5956) );
  NANDN U13971 ( .A(n5959), .B(n5960), .Z(n5958) );
  NANDN U13972 ( .A(n5960), .B(n5959), .Z(n5955) );
  XOR U13973 ( .A(n5952), .B(n5961), .Z(N64858) );
  XNOR U13974 ( .A(n5950), .B(n5954), .Z(n5961) );
  XOR U13975 ( .A(n5947), .B(n5962), .Z(n5954) );
  XNOR U13976 ( .A(n5944), .B(n5946), .Z(n5962) );
  AND U13977 ( .A(n5963), .B(n5964), .Z(n5946) );
  NANDN U13978 ( .A(n5965), .B(n5966), .Z(n5964) );
  OR U13979 ( .A(n5967), .B(n5968), .Z(n5966) );
  IV U13980 ( .A(n5969), .Z(n5968) );
  NANDN U13981 ( .A(n5969), .B(n5967), .Z(n5963) );
  AND U13982 ( .A(n5970), .B(n5971), .Z(n5944) );
  NAND U13983 ( .A(n5972), .B(n5973), .Z(n5971) );
  NANDN U13984 ( .A(n5974), .B(n5975), .Z(n5973) );
  NANDN U13985 ( .A(n5975), .B(n5974), .Z(n5970) );
  IV U13986 ( .A(n5976), .Z(n5975) );
  NAND U13987 ( .A(n5977), .B(n5978), .Z(n5947) );
  NANDN U13988 ( .A(n5979), .B(n5980), .Z(n5978) );
  NANDN U13989 ( .A(n5981), .B(n5982), .Z(n5980) );
  NANDN U13990 ( .A(n5982), .B(n5981), .Z(n5977) );
  IV U13991 ( .A(n5983), .Z(n5981) );
  AND U13992 ( .A(n5984), .B(n5985), .Z(n5950) );
  NAND U13993 ( .A(n5986), .B(n5987), .Z(n5985) );
  NANDN U13994 ( .A(n5988), .B(n5989), .Z(n5987) );
  NANDN U13995 ( .A(n5989), .B(n5988), .Z(n5984) );
  XOR U13996 ( .A(n5960), .B(n5990), .Z(n5952) );
  XNOR U13997 ( .A(n5957), .B(n5959), .Z(n5990) );
  AND U13998 ( .A(n5991), .B(n5992), .Z(n5959) );
  NANDN U13999 ( .A(n5993), .B(n5994), .Z(n5992) );
  OR U14000 ( .A(n5995), .B(n5996), .Z(n5994) );
  IV U14001 ( .A(n5997), .Z(n5996) );
  NANDN U14002 ( .A(n5997), .B(n5995), .Z(n5991) );
  AND U14003 ( .A(n5998), .B(n5999), .Z(n5957) );
  NAND U14004 ( .A(n6000), .B(n6001), .Z(n5999) );
  NANDN U14005 ( .A(n6002), .B(n6003), .Z(n6001) );
  NANDN U14006 ( .A(n6003), .B(n6002), .Z(n5998) );
  IV U14007 ( .A(n6004), .Z(n6003) );
  NAND U14008 ( .A(n6005), .B(n6006), .Z(n5960) );
  NANDN U14009 ( .A(n6007), .B(n6008), .Z(n6006) );
  NANDN U14010 ( .A(n6009), .B(n6010), .Z(n6008) );
  NANDN U14011 ( .A(n6010), .B(n6009), .Z(n6005) );
  IV U14012 ( .A(n6011), .Z(n6009) );
  XOR U14013 ( .A(n5986), .B(n6012), .Z(N64857) );
  XNOR U14014 ( .A(n5989), .B(n5988), .Z(n6012) );
  XNOR U14015 ( .A(n6000), .B(n6013), .Z(n5988) );
  XNOR U14016 ( .A(n6004), .B(n6002), .Z(n6013) );
  XOR U14017 ( .A(n6010), .B(n6014), .Z(n6002) );
  XNOR U14018 ( .A(n6007), .B(n6011), .Z(n6014) );
  AND U14019 ( .A(n6015), .B(n6016), .Z(n6011) );
  NAND U14020 ( .A(n6017), .B(n6018), .Z(n6016) );
  NAND U14021 ( .A(n6019), .B(n6020), .Z(n6015) );
  AND U14022 ( .A(n6021), .B(n6022), .Z(n6007) );
  NAND U14023 ( .A(n6023), .B(n6024), .Z(n6022) );
  NAND U14024 ( .A(n6025), .B(n6026), .Z(n6021) );
  NANDN U14025 ( .A(n6027), .B(n6028), .Z(n6010) );
  ANDN U14026 ( .B(n6029), .A(n6030), .Z(n6004) );
  XNOR U14027 ( .A(n5995), .B(n6031), .Z(n6000) );
  XNOR U14028 ( .A(n5993), .B(n5997), .Z(n6031) );
  AND U14029 ( .A(n6032), .B(n6033), .Z(n5997) );
  NAND U14030 ( .A(n6034), .B(n6035), .Z(n6033) );
  NAND U14031 ( .A(n6036), .B(n6037), .Z(n6032) );
  AND U14032 ( .A(n6038), .B(n6039), .Z(n5993) );
  NAND U14033 ( .A(n6040), .B(n6041), .Z(n6039) );
  NAND U14034 ( .A(n6042), .B(n6043), .Z(n6038) );
  AND U14035 ( .A(n6044), .B(n6045), .Z(n5995) );
  NAND U14036 ( .A(n6046), .B(n6047), .Z(n5989) );
  XNOR U14037 ( .A(n5972), .B(n6048), .Z(n5986) );
  XNOR U14038 ( .A(n5976), .B(n5974), .Z(n6048) );
  XOR U14039 ( .A(n5982), .B(n6049), .Z(n5974) );
  XNOR U14040 ( .A(n5979), .B(n5983), .Z(n6049) );
  AND U14041 ( .A(n6050), .B(n6051), .Z(n5983) );
  NAND U14042 ( .A(n6052), .B(n6053), .Z(n6051) );
  NAND U14043 ( .A(n6054), .B(n6055), .Z(n6050) );
  AND U14044 ( .A(n6056), .B(n6057), .Z(n5979) );
  NAND U14045 ( .A(n6058), .B(n6059), .Z(n6057) );
  NAND U14046 ( .A(n6060), .B(n6061), .Z(n6056) );
  NANDN U14047 ( .A(n6062), .B(n6063), .Z(n5982) );
  ANDN U14048 ( .B(n6064), .A(n6065), .Z(n5976) );
  XNOR U14049 ( .A(n5967), .B(n6066), .Z(n5972) );
  XNOR U14050 ( .A(n5965), .B(n5969), .Z(n6066) );
  AND U14051 ( .A(n6067), .B(n6068), .Z(n5969) );
  NAND U14052 ( .A(n6069), .B(n6070), .Z(n6068) );
  NAND U14053 ( .A(n6071), .B(n6072), .Z(n6067) );
  AND U14054 ( .A(n6073), .B(n6074), .Z(n5965) );
  NAND U14055 ( .A(n6075), .B(n6076), .Z(n6074) );
  NAND U14056 ( .A(n6077), .B(n6078), .Z(n6073) );
  AND U14057 ( .A(n6079), .B(n6080), .Z(n5967) );
  XOR U14058 ( .A(n6047), .B(n6046), .Z(N64856) );
  XNOR U14059 ( .A(n6064), .B(n6065), .Z(n6046) );
  XNOR U14060 ( .A(n6079), .B(n6080), .Z(n6065) );
  XOR U14061 ( .A(n6076), .B(n6075), .Z(n6080) );
  XOR U14062 ( .A(y[7884]), .B(x[7884]), .Z(n6075) );
  XOR U14063 ( .A(n6078), .B(n6077), .Z(n6076) );
  XOR U14064 ( .A(y[7886]), .B(x[7886]), .Z(n6077) );
  XOR U14065 ( .A(y[7885]), .B(x[7885]), .Z(n6078) );
  XOR U14066 ( .A(n6070), .B(n6069), .Z(n6079) );
  XOR U14067 ( .A(n6072), .B(n6071), .Z(n6069) );
  XOR U14068 ( .A(y[7883]), .B(x[7883]), .Z(n6071) );
  XOR U14069 ( .A(y[7882]), .B(x[7882]), .Z(n6072) );
  XOR U14070 ( .A(y[7881]), .B(x[7881]), .Z(n6070) );
  XNOR U14071 ( .A(n6063), .B(n6062), .Z(n6064) );
  XNOR U14072 ( .A(n6059), .B(n6058), .Z(n6062) );
  XOR U14073 ( .A(n6061), .B(n6060), .Z(n6058) );
  XOR U14074 ( .A(y[7880]), .B(x[7880]), .Z(n6060) );
  XOR U14075 ( .A(y[7879]), .B(x[7879]), .Z(n6061) );
  XOR U14076 ( .A(y[7878]), .B(x[7878]), .Z(n6059) );
  XOR U14077 ( .A(n6053), .B(n6052), .Z(n6063) );
  XOR U14078 ( .A(n6055), .B(n6054), .Z(n6052) );
  XOR U14079 ( .A(y[7877]), .B(x[7877]), .Z(n6054) );
  XOR U14080 ( .A(y[7876]), .B(x[7876]), .Z(n6055) );
  XOR U14081 ( .A(y[7875]), .B(x[7875]), .Z(n6053) );
  XNOR U14082 ( .A(n6029), .B(n6030), .Z(n6047) );
  XNOR U14083 ( .A(n6044), .B(n6045), .Z(n6030) );
  XOR U14084 ( .A(n6041), .B(n6040), .Z(n6045) );
  XOR U14085 ( .A(y[7872]), .B(x[7872]), .Z(n6040) );
  XOR U14086 ( .A(n6043), .B(n6042), .Z(n6041) );
  XOR U14087 ( .A(y[7874]), .B(x[7874]), .Z(n6042) );
  XOR U14088 ( .A(y[7873]), .B(x[7873]), .Z(n6043) );
  XOR U14089 ( .A(n6035), .B(n6034), .Z(n6044) );
  XOR U14090 ( .A(n6037), .B(n6036), .Z(n6034) );
  XOR U14091 ( .A(y[7871]), .B(x[7871]), .Z(n6036) );
  XOR U14092 ( .A(y[7870]), .B(x[7870]), .Z(n6037) );
  XOR U14093 ( .A(y[7869]), .B(x[7869]), .Z(n6035) );
  XNOR U14094 ( .A(n6028), .B(n6027), .Z(n6029) );
  XNOR U14095 ( .A(n6024), .B(n6023), .Z(n6027) );
  XOR U14096 ( .A(n6026), .B(n6025), .Z(n6023) );
  XOR U14097 ( .A(y[7868]), .B(x[7868]), .Z(n6025) );
  XOR U14098 ( .A(y[7867]), .B(x[7867]), .Z(n6026) );
  XOR U14099 ( .A(y[7866]), .B(x[7866]), .Z(n6024) );
  XOR U14100 ( .A(n6018), .B(n6017), .Z(n6028) );
  XOR U14101 ( .A(n6020), .B(n6019), .Z(n6017) );
  XOR U14102 ( .A(y[7865]), .B(x[7865]), .Z(n6019) );
  XOR U14103 ( .A(y[7864]), .B(x[7864]), .Z(n6020) );
  XOR U14104 ( .A(y[7863]), .B(x[7863]), .Z(n6018) );
  NAND U14105 ( .A(n6081), .B(n6082), .Z(N64847) );
  NAND U14106 ( .A(n6083), .B(n6084), .Z(n6082) );
  NANDN U14107 ( .A(n6085), .B(n6086), .Z(n6084) );
  NANDN U14108 ( .A(n6086), .B(n6085), .Z(n6081) );
  XOR U14109 ( .A(n6085), .B(n6087), .Z(N64846) );
  XNOR U14110 ( .A(n6083), .B(n6086), .Z(n6087) );
  NAND U14111 ( .A(n6088), .B(n6089), .Z(n6086) );
  NAND U14112 ( .A(n6090), .B(n6091), .Z(n6089) );
  NANDN U14113 ( .A(n6092), .B(n6093), .Z(n6091) );
  NANDN U14114 ( .A(n6093), .B(n6092), .Z(n6088) );
  AND U14115 ( .A(n6094), .B(n6095), .Z(n6083) );
  NAND U14116 ( .A(n6096), .B(n6097), .Z(n6095) );
  NANDN U14117 ( .A(n6098), .B(n6099), .Z(n6097) );
  NANDN U14118 ( .A(n6099), .B(n6098), .Z(n6094) );
  IV U14119 ( .A(n6100), .Z(n6099) );
  AND U14120 ( .A(n6101), .B(n6102), .Z(n6085) );
  NAND U14121 ( .A(n6103), .B(n6104), .Z(n6102) );
  NANDN U14122 ( .A(n6105), .B(n6106), .Z(n6104) );
  NANDN U14123 ( .A(n6106), .B(n6105), .Z(n6101) );
  XOR U14124 ( .A(n6098), .B(n6107), .Z(N64845) );
  XNOR U14125 ( .A(n6096), .B(n6100), .Z(n6107) );
  XOR U14126 ( .A(n6093), .B(n6108), .Z(n6100) );
  XNOR U14127 ( .A(n6090), .B(n6092), .Z(n6108) );
  AND U14128 ( .A(n6109), .B(n6110), .Z(n6092) );
  NANDN U14129 ( .A(n6111), .B(n6112), .Z(n6110) );
  OR U14130 ( .A(n6113), .B(n6114), .Z(n6112) );
  IV U14131 ( .A(n6115), .Z(n6114) );
  NANDN U14132 ( .A(n6115), .B(n6113), .Z(n6109) );
  AND U14133 ( .A(n6116), .B(n6117), .Z(n6090) );
  NAND U14134 ( .A(n6118), .B(n6119), .Z(n6117) );
  NANDN U14135 ( .A(n6120), .B(n6121), .Z(n6119) );
  NANDN U14136 ( .A(n6121), .B(n6120), .Z(n6116) );
  IV U14137 ( .A(n6122), .Z(n6121) );
  NAND U14138 ( .A(n6123), .B(n6124), .Z(n6093) );
  NANDN U14139 ( .A(n6125), .B(n6126), .Z(n6124) );
  NANDN U14140 ( .A(n6127), .B(n6128), .Z(n6126) );
  NANDN U14141 ( .A(n6128), .B(n6127), .Z(n6123) );
  IV U14142 ( .A(n6129), .Z(n6127) );
  AND U14143 ( .A(n6130), .B(n6131), .Z(n6096) );
  NAND U14144 ( .A(n6132), .B(n6133), .Z(n6131) );
  NANDN U14145 ( .A(n6134), .B(n6135), .Z(n6133) );
  NANDN U14146 ( .A(n6135), .B(n6134), .Z(n6130) );
  XOR U14147 ( .A(n6106), .B(n6136), .Z(n6098) );
  XNOR U14148 ( .A(n6103), .B(n6105), .Z(n6136) );
  AND U14149 ( .A(n6137), .B(n6138), .Z(n6105) );
  NANDN U14150 ( .A(n6139), .B(n6140), .Z(n6138) );
  OR U14151 ( .A(n6141), .B(n6142), .Z(n6140) );
  IV U14152 ( .A(n6143), .Z(n6142) );
  NANDN U14153 ( .A(n6143), .B(n6141), .Z(n6137) );
  AND U14154 ( .A(n6144), .B(n6145), .Z(n6103) );
  NAND U14155 ( .A(n6146), .B(n6147), .Z(n6145) );
  NANDN U14156 ( .A(n6148), .B(n6149), .Z(n6147) );
  NANDN U14157 ( .A(n6149), .B(n6148), .Z(n6144) );
  IV U14158 ( .A(n6150), .Z(n6149) );
  NAND U14159 ( .A(n6151), .B(n6152), .Z(n6106) );
  NANDN U14160 ( .A(n6153), .B(n6154), .Z(n6152) );
  NANDN U14161 ( .A(n6155), .B(n6156), .Z(n6154) );
  NANDN U14162 ( .A(n6156), .B(n6155), .Z(n6151) );
  IV U14163 ( .A(n6157), .Z(n6155) );
  XOR U14164 ( .A(n6132), .B(n6158), .Z(N64844) );
  XNOR U14165 ( .A(n6135), .B(n6134), .Z(n6158) );
  XNOR U14166 ( .A(n6146), .B(n6159), .Z(n6134) );
  XNOR U14167 ( .A(n6150), .B(n6148), .Z(n6159) );
  XOR U14168 ( .A(n6156), .B(n6160), .Z(n6148) );
  XNOR U14169 ( .A(n6153), .B(n6157), .Z(n6160) );
  AND U14170 ( .A(n6161), .B(n6162), .Z(n6157) );
  NAND U14171 ( .A(n6163), .B(n6164), .Z(n6162) );
  NAND U14172 ( .A(n6165), .B(n6166), .Z(n6161) );
  AND U14173 ( .A(n6167), .B(n6168), .Z(n6153) );
  NAND U14174 ( .A(n6169), .B(n6170), .Z(n6168) );
  NAND U14175 ( .A(n6171), .B(n6172), .Z(n6167) );
  NANDN U14176 ( .A(n6173), .B(n6174), .Z(n6156) );
  ANDN U14177 ( .B(n6175), .A(n6176), .Z(n6150) );
  XNOR U14178 ( .A(n6141), .B(n6177), .Z(n6146) );
  XNOR U14179 ( .A(n6139), .B(n6143), .Z(n6177) );
  AND U14180 ( .A(n6178), .B(n6179), .Z(n6143) );
  NAND U14181 ( .A(n6180), .B(n6181), .Z(n6179) );
  NAND U14182 ( .A(n6182), .B(n6183), .Z(n6178) );
  AND U14183 ( .A(n6184), .B(n6185), .Z(n6139) );
  NAND U14184 ( .A(n6186), .B(n6187), .Z(n6185) );
  NAND U14185 ( .A(n6188), .B(n6189), .Z(n6184) );
  AND U14186 ( .A(n6190), .B(n6191), .Z(n6141) );
  NAND U14187 ( .A(n6192), .B(n6193), .Z(n6135) );
  XNOR U14188 ( .A(n6118), .B(n6194), .Z(n6132) );
  XNOR U14189 ( .A(n6122), .B(n6120), .Z(n6194) );
  XOR U14190 ( .A(n6128), .B(n6195), .Z(n6120) );
  XNOR U14191 ( .A(n6125), .B(n6129), .Z(n6195) );
  AND U14192 ( .A(n6196), .B(n6197), .Z(n6129) );
  NAND U14193 ( .A(n6198), .B(n6199), .Z(n6197) );
  NAND U14194 ( .A(n6200), .B(n6201), .Z(n6196) );
  AND U14195 ( .A(n6202), .B(n6203), .Z(n6125) );
  NAND U14196 ( .A(n6204), .B(n6205), .Z(n6203) );
  NAND U14197 ( .A(n6206), .B(n6207), .Z(n6202) );
  NANDN U14198 ( .A(n6208), .B(n6209), .Z(n6128) );
  ANDN U14199 ( .B(n6210), .A(n6211), .Z(n6122) );
  XNOR U14200 ( .A(n6113), .B(n6212), .Z(n6118) );
  XNOR U14201 ( .A(n6111), .B(n6115), .Z(n6212) );
  AND U14202 ( .A(n6213), .B(n6214), .Z(n6115) );
  NAND U14203 ( .A(n6215), .B(n6216), .Z(n6214) );
  NAND U14204 ( .A(n6217), .B(n6218), .Z(n6213) );
  AND U14205 ( .A(n6219), .B(n6220), .Z(n6111) );
  NAND U14206 ( .A(n6221), .B(n6222), .Z(n6220) );
  NAND U14207 ( .A(n6223), .B(n6224), .Z(n6219) );
  AND U14208 ( .A(n6225), .B(n6226), .Z(n6113) );
  XOR U14209 ( .A(n6193), .B(n6192), .Z(N64843) );
  XNOR U14210 ( .A(n6210), .B(n6211), .Z(n6192) );
  XNOR U14211 ( .A(n6225), .B(n6226), .Z(n6211) );
  XOR U14212 ( .A(n6222), .B(n6221), .Z(n6226) );
  XOR U14213 ( .A(y[7860]), .B(x[7860]), .Z(n6221) );
  XOR U14214 ( .A(n6224), .B(n6223), .Z(n6222) );
  XOR U14215 ( .A(y[7862]), .B(x[7862]), .Z(n6223) );
  XOR U14216 ( .A(y[7861]), .B(x[7861]), .Z(n6224) );
  XOR U14217 ( .A(n6216), .B(n6215), .Z(n6225) );
  XOR U14218 ( .A(n6218), .B(n6217), .Z(n6215) );
  XOR U14219 ( .A(y[7859]), .B(x[7859]), .Z(n6217) );
  XOR U14220 ( .A(y[7858]), .B(x[7858]), .Z(n6218) );
  XOR U14221 ( .A(y[7857]), .B(x[7857]), .Z(n6216) );
  XNOR U14222 ( .A(n6209), .B(n6208), .Z(n6210) );
  XNOR U14223 ( .A(n6205), .B(n6204), .Z(n6208) );
  XOR U14224 ( .A(n6207), .B(n6206), .Z(n6204) );
  XOR U14225 ( .A(y[7856]), .B(x[7856]), .Z(n6206) );
  XOR U14226 ( .A(y[7855]), .B(x[7855]), .Z(n6207) );
  XOR U14227 ( .A(y[7854]), .B(x[7854]), .Z(n6205) );
  XOR U14228 ( .A(n6199), .B(n6198), .Z(n6209) );
  XOR U14229 ( .A(n6201), .B(n6200), .Z(n6198) );
  XOR U14230 ( .A(y[7853]), .B(x[7853]), .Z(n6200) );
  XOR U14231 ( .A(y[7852]), .B(x[7852]), .Z(n6201) );
  XOR U14232 ( .A(y[7851]), .B(x[7851]), .Z(n6199) );
  XNOR U14233 ( .A(n6175), .B(n6176), .Z(n6193) );
  XNOR U14234 ( .A(n6190), .B(n6191), .Z(n6176) );
  XOR U14235 ( .A(n6187), .B(n6186), .Z(n6191) );
  XOR U14236 ( .A(y[7848]), .B(x[7848]), .Z(n6186) );
  XOR U14237 ( .A(n6189), .B(n6188), .Z(n6187) );
  XOR U14238 ( .A(y[7850]), .B(x[7850]), .Z(n6188) );
  XOR U14239 ( .A(y[7849]), .B(x[7849]), .Z(n6189) );
  XOR U14240 ( .A(n6181), .B(n6180), .Z(n6190) );
  XOR U14241 ( .A(n6183), .B(n6182), .Z(n6180) );
  XOR U14242 ( .A(y[7847]), .B(x[7847]), .Z(n6182) );
  XOR U14243 ( .A(y[7846]), .B(x[7846]), .Z(n6183) );
  XOR U14244 ( .A(y[7845]), .B(x[7845]), .Z(n6181) );
  XNOR U14245 ( .A(n6174), .B(n6173), .Z(n6175) );
  XNOR U14246 ( .A(n6170), .B(n6169), .Z(n6173) );
  XOR U14247 ( .A(n6172), .B(n6171), .Z(n6169) );
  XOR U14248 ( .A(y[7844]), .B(x[7844]), .Z(n6171) );
  XOR U14249 ( .A(y[7843]), .B(x[7843]), .Z(n6172) );
  XOR U14250 ( .A(y[7842]), .B(x[7842]), .Z(n6170) );
  XOR U14251 ( .A(n6164), .B(n6163), .Z(n6174) );
  XOR U14252 ( .A(n6166), .B(n6165), .Z(n6163) );
  XOR U14253 ( .A(y[7841]), .B(x[7841]), .Z(n6165) );
  XOR U14254 ( .A(y[7840]), .B(x[7840]), .Z(n6166) );
  XOR U14255 ( .A(y[7839]), .B(x[7839]), .Z(n6164) );
  NAND U14256 ( .A(n6227), .B(n6228), .Z(N64834) );
  NAND U14257 ( .A(n6229), .B(n6230), .Z(n6228) );
  NANDN U14258 ( .A(n6231), .B(n6232), .Z(n6230) );
  NANDN U14259 ( .A(n6232), .B(n6231), .Z(n6227) );
  XOR U14260 ( .A(n6231), .B(n6233), .Z(N64833) );
  XNOR U14261 ( .A(n6229), .B(n6232), .Z(n6233) );
  NAND U14262 ( .A(n6234), .B(n6235), .Z(n6232) );
  NAND U14263 ( .A(n6236), .B(n6237), .Z(n6235) );
  NANDN U14264 ( .A(n6238), .B(n6239), .Z(n6237) );
  NANDN U14265 ( .A(n6239), .B(n6238), .Z(n6234) );
  AND U14266 ( .A(n6240), .B(n6241), .Z(n6229) );
  NAND U14267 ( .A(n6242), .B(n6243), .Z(n6241) );
  NANDN U14268 ( .A(n6244), .B(n6245), .Z(n6243) );
  NANDN U14269 ( .A(n6245), .B(n6244), .Z(n6240) );
  IV U14270 ( .A(n6246), .Z(n6245) );
  AND U14271 ( .A(n6247), .B(n6248), .Z(n6231) );
  NAND U14272 ( .A(n6249), .B(n6250), .Z(n6248) );
  NANDN U14273 ( .A(n6251), .B(n6252), .Z(n6250) );
  NANDN U14274 ( .A(n6252), .B(n6251), .Z(n6247) );
  XOR U14275 ( .A(n6244), .B(n6253), .Z(N64832) );
  XNOR U14276 ( .A(n6242), .B(n6246), .Z(n6253) );
  XOR U14277 ( .A(n6239), .B(n6254), .Z(n6246) );
  XNOR U14278 ( .A(n6236), .B(n6238), .Z(n6254) );
  AND U14279 ( .A(n6255), .B(n6256), .Z(n6238) );
  NANDN U14280 ( .A(n6257), .B(n6258), .Z(n6256) );
  OR U14281 ( .A(n6259), .B(n6260), .Z(n6258) );
  IV U14282 ( .A(n6261), .Z(n6260) );
  NANDN U14283 ( .A(n6261), .B(n6259), .Z(n6255) );
  AND U14284 ( .A(n6262), .B(n6263), .Z(n6236) );
  NAND U14285 ( .A(n6264), .B(n6265), .Z(n6263) );
  NANDN U14286 ( .A(n6266), .B(n6267), .Z(n6265) );
  NANDN U14287 ( .A(n6267), .B(n6266), .Z(n6262) );
  IV U14288 ( .A(n6268), .Z(n6267) );
  NAND U14289 ( .A(n6269), .B(n6270), .Z(n6239) );
  NANDN U14290 ( .A(n6271), .B(n6272), .Z(n6270) );
  NANDN U14291 ( .A(n6273), .B(n6274), .Z(n6272) );
  NANDN U14292 ( .A(n6274), .B(n6273), .Z(n6269) );
  IV U14293 ( .A(n6275), .Z(n6273) );
  AND U14294 ( .A(n6276), .B(n6277), .Z(n6242) );
  NAND U14295 ( .A(n6278), .B(n6279), .Z(n6277) );
  NANDN U14296 ( .A(n6280), .B(n6281), .Z(n6279) );
  NANDN U14297 ( .A(n6281), .B(n6280), .Z(n6276) );
  XOR U14298 ( .A(n6252), .B(n6282), .Z(n6244) );
  XNOR U14299 ( .A(n6249), .B(n6251), .Z(n6282) );
  AND U14300 ( .A(n6283), .B(n6284), .Z(n6251) );
  NANDN U14301 ( .A(n6285), .B(n6286), .Z(n6284) );
  OR U14302 ( .A(n6287), .B(n6288), .Z(n6286) );
  IV U14303 ( .A(n6289), .Z(n6288) );
  NANDN U14304 ( .A(n6289), .B(n6287), .Z(n6283) );
  AND U14305 ( .A(n6290), .B(n6291), .Z(n6249) );
  NAND U14306 ( .A(n6292), .B(n6293), .Z(n6291) );
  NANDN U14307 ( .A(n6294), .B(n6295), .Z(n6293) );
  NANDN U14308 ( .A(n6295), .B(n6294), .Z(n6290) );
  IV U14309 ( .A(n6296), .Z(n6295) );
  NAND U14310 ( .A(n6297), .B(n6298), .Z(n6252) );
  NANDN U14311 ( .A(n6299), .B(n6300), .Z(n6298) );
  NANDN U14312 ( .A(n6301), .B(n6302), .Z(n6300) );
  NANDN U14313 ( .A(n6302), .B(n6301), .Z(n6297) );
  IV U14314 ( .A(n6303), .Z(n6301) );
  XOR U14315 ( .A(n6278), .B(n6304), .Z(N64831) );
  XNOR U14316 ( .A(n6281), .B(n6280), .Z(n6304) );
  XNOR U14317 ( .A(n6292), .B(n6305), .Z(n6280) );
  XNOR U14318 ( .A(n6296), .B(n6294), .Z(n6305) );
  XOR U14319 ( .A(n6302), .B(n6306), .Z(n6294) );
  XNOR U14320 ( .A(n6299), .B(n6303), .Z(n6306) );
  AND U14321 ( .A(n6307), .B(n6308), .Z(n6303) );
  NAND U14322 ( .A(n6309), .B(n6310), .Z(n6308) );
  NAND U14323 ( .A(n6311), .B(n6312), .Z(n6307) );
  AND U14324 ( .A(n6313), .B(n6314), .Z(n6299) );
  NAND U14325 ( .A(n6315), .B(n6316), .Z(n6314) );
  NAND U14326 ( .A(n6317), .B(n6318), .Z(n6313) );
  NANDN U14327 ( .A(n6319), .B(n6320), .Z(n6302) );
  ANDN U14328 ( .B(n6321), .A(n6322), .Z(n6296) );
  XNOR U14329 ( .A(n6287), .B(n6323), .Z(n6292) );
  XNOR U14330 ( .A(n6285), .B(n6289), .Z(n6323) );
  AND U14331 ( .A(n6324), .B(n6325), .Z(n6289) );
  NAND U14332 ( .A(n6326), .B(n6327), .Z(n6325) );
  NAND U14333 ( .A(n6328), .B(n6329), .Z(n6324) );
  AND U14334 ( .A(n6330), .B(n6331), .Z(n6285) );
  NAND U14335 ( .A(n6332), .B(n6333), .Z(n6331) );
  NAND U14336 ( .A(n6334), .B(n6335), .Z(n6330) );
  AND U14337 ( .A(n6336), .B(n6337), .Z(n6287) );
  NAND U14338 ( .A(n6338), .B(n6339), .Z(n6281) );
  XNOR U14339 ( .A(n6264), .B(n6340), .Z(n6278) );
  XNOR U14340 ( .A(n6268), .B(n6266), .Z(n6340) );
  XOR U14341 ( .A(n6274), .B(n6341), .Z(n6266) );
  XNOR U14342 ( .A(n6271), .B(n6275), .Z(n6341) );
  AND U14343 ( .A(n6342), .B(n6343), .Z(n6275) );
  NAND U14344 ( .A(n6344), .B(n6345), .Z(n6343) );
  NAND U14345 ( .A(n6346), .B(n6347), .Z(n6342) );
  AND U14346 ( .A(n6348), .B(n6349), .Z(n6271) );
  NAND U14347 ( .A(n6350), .B(n6351), .Z(n6349) );
  NAND U14348 ( .A(n6352), .B(n6353), .Z(n6348) );
  NANDN U14349 ( .A(n6354), .B(n6355), .Z(n6274) );
  ANDN U14350 ( .B(n6356), .A(n6357), .Z(n6268) );
  XNOR U14351 ( .A(n6259), .B(n6358), .Z(n6264) );
  XNOR U14352 ( .A(n6257), .B(n6261), .Z(n6358) );
  AND U14353 ( .A(n6359), .B(n6360), .Z(n6261) );
  NAND U14354 ( .A(n6361), .B(n6362), .Z(n6360) );
  NAND U14355 ( .A(n6363), .B(n6364), .Z(n6359) );
  AND U14356 ( .A(n6365), .B(n6366), .Z(n6257) );
  NAND U14357 ( .A(n6367), .B(n6368), .Z(n6366) );
  NAND U14358 ( .A(n6369), .B(n6370), .Z(n6365) );
  AND U14359 ( .A(n6371), .B(n6372), .Z(n6259) );
  XOR U14360 ( .A(n6339), .B(n6338), .Z(N64830) );
  XNOR U14361 ( .A(n6356), .B(n6357), .Z(n6338) );
  XNOR U14362 ( .A(n6371), .B(n6372), .Z(n6357) );
  XOR U14363 ( .A(n6368), .B(n6367), .Z(n6372) );
  XOR U14364 ( .A(y[7836]), .B(x[7836]), .Z(n6367) );
  XOR U14365 ( .A(n6370), .B(n6369), .Z(n6368) );
  XOR U14366 ( .A(y[7838]), .B(x[7838]), .Z(n6369) );
  XOR U14367 ( .A(y[7837]), .B(x[7837]), .Z(n6370) );
  XOR U14368 ( .A(n6362), .B(n6361), .Z(n6371) );
  XOR U14369 ( .A(n6364), .B(n6363), .Z(n6361) );
  XOR U14370 ( .A(y[7835]), .B(x[7835]), .Z(n6363) );
  XOR U14371 ( .A(y[7834]), .B(x[7834]), .Z(n6364) );
  XOR U14372 ( .A(y[7833]), .B(x[7833]), .Z(n6362) );
  XNOR U14373 ( .A(n6355), .B(n6354), .Z(n6356) );
  XNOR U14374 ( .A(n6351), .B(n6350), .Z(n6354) );
  XOR U14375 ( .A(n6353), .B(n6352), .Z(n6350) );
  XOR U14376 ( .A(y[7832]), .B(x[7832]), .Z(n6352) );
  XOR U14377 ( .A(y[7831]), .B(x[7831]), .Z(n6353) );
  XOR U14378 ( .A(y[7830]), .B(x[7830]), .Z(n6351) );
  XOR U14379 ( .A(n6345), .B(n6344), .Z(n6355) );
  XOR U14380 ( .A(n6347), .B(n6346), .Z(n6344) );
  XOR U14381 ( .A(y[7829]), .B(x[7829]), .Z(n6346) );
  XOR U14382 ( .A(y[7828]), .B(x[7828]), .Z(n6347) );
  XOR U14383 ( .A(y[7827]), .B(x[7827]), .Z(n6345) );
  XNOR U14384 ( .A(n6321), .B(n6322), .Z(n6339) );
  XNOR U14385 ( .A(n6336), .B(n6337), .Z(n6322) );
  XOR U14386 ( .A(n6333), .B(n6332), .Z(n6337) );
  XOR U14387 ( .A(y[7824]), .B(x[7824]), .Z(n6332) );
  XOR U14388 ( .A(n6335), .B(n6334), .Z(n6333) );
  XOR U14389 ( .A(y[7826]), .B(x[7826]), .Z(n6334) );
  XOR U14390 ( .A(y[7825]), .B(x[7825]), .Z(n6335) );
  XOR U14391 ( .A(n6327), .B(n6326), .Z(n6336) );
  XOR U14392 ( .A(n6329), .B(n6328), .Z(n6326) );
  XOR U14393 ( .A(y[7823]), .B(x[7823]), .Z(n6328) );
  XOR U14394 ( .A(y[7822]), .B(x[7822]), .Z(n6329) );
  XOR U14395 ( .A(y[7821]), .B(x[7821]), .Z(n6327) );
  XNOR U14396 ( .A(n6320), .B(n6319), .Z(n6321) );
  XNOR U14397 ( .A(n6316), .B(n6315), .Z(n6319) );
  XOR U14398 ( .A(n6318), .B(n6317), .Z(n6315) );
  XOR U14399 ( .A(y[7820]), .B(x[7820]), .Z(n6317) );
  XOR U14400 ( .A(y[7819]), .B(x[7819]), .Z(n6318) );
  XOR U14401 ( .A(y[7818]), .B(x[7818]), .Z(n6316) );
  XOR U14402 ( .A(n6310), .B(n6309), .Z(n6320) );
  XOR U14403 ( .A(n6312), .B(n6311), .Z(n6309) );
  XOR U14404 ( .A(y[7817]), .B(x[7817]), .Z(n6311) );
  XOR U14405 ( .A(y[7816]), .B(x[7816]), .Z(n6312) );
  XOR U14406 ( .A(y[7815]), .B(x[7815]), .Z(n6310) );
  NAND U14407 ( .A(n6373), .B(n6374), .Z(N64821) );
  NAND U14408 ( .A(n6375), .B(n6376), .Z(n6374) );
  NANDN U14409 ( .A(n6377), .B(n6378), .Z(n6376) );
  NANDN U14410 ( .A(n6378), .B(n6377), .Z(n6373) );
  XOR U14411 ( .A(n6377), .B(n6379), .Z(N64820) );
  XNOR U14412 ( .A(n6375), .B(n6378), .Z(n6379) );
  NAND U14413 ( .A(n6380), .B(n6381), .Z(n6378) );
  NAND U14414 ( .A(n6382), .B(n6383), .Z(n6381) );
  NANDN U14415 ( .A(n6384), .B(n6385), .Z(n6383) );
  NANDN U14416 ( .A(n6385), .B(n6384), .Z(n6380) );
  AND U14417 ( .A(n6386), .B(n6387), .Z(n6375) );
  NAND U14418 ( .A(n6388), .B(n6389), .Z(n6387) );
  NANDN U14419 ( .A(n6390), .B(n6391), .Z(n6389) );
  NANDN U14420 ( .A(n6391), .B(n6390), .Z(n6386) );
  IV U14421 ( .A(n6392), .Z(n6391) );
  AND U14422 ( .A(n6393), .B(n6394), .Z(n6377) );
  NAND U14423 ( .A(n6395), .B(n6396), .Z(n6394) );
  NANDN U14424 ( .A(n6397), .B(n6398), .Z(n6396) );
  NANDN U14425 ( .A(n6398), .B(n6397), .Z(n6393) );
  XOR U14426 ( .A(n6390), .B(n6399), .Z(N64819) );
  XNOR U14427 ( .A(n6388), .B(n6392), .Z(n6399) );
  XOR U14428 ( .A(n6385), .B(n6400), .Z(n6392) );
  XNOR U14429 ( .A(n6382), .B(n6384), .Z(n6400) );
  AND U14430 ( .A(n6401), .B(n6402), .Z(n6384) );
  NANDN U14431 ( .A(n6403), .B(n6404), .Z(n6402) );
  OR U14432 ( .A(n6405), .B(n6406), .Z(n6404) );
  IV U14433 ( .A(n6407), .Z(n6406) );
  NANDN U14434 ( .A(n6407), .B(n6405), .Z(n6401) );
  AND U14435 ( .A(n6408), .B(n6409), .Z(n6382) );
  NAND U14436 ( .A(n6410), .B(n6411), .Z(n6409) );
  NANDN U14437 ( .A(n6412), .B(n6413), .Z(n6411) );
  NANDN U14438 ( .A(n6413), .B(n6412), .Z(n6408) );
  IV U14439 ( .A(n6414), .Z(n6413) );
  NAND U14440 ( .A(n6415), .B(n6416), .Z(n6385) );
  NANDN U14441 ( .A(n6417), .B(n6418), .Z(n6416) );
  NANDN U14442 ( .A(n6419), .B(n6420), .Z(n6418) );
  NANDN U14443 ( .A(n6420), .B(n6419), .Z(n6415) );
  IV U14444 ( .A(n6421), .Z(n6419) );
  AND U14445 ( .A(n6422), .B(n6423), .Z(n6388) );
  NAND U14446 ( .A(n6424), .B(n6425), .Z(n6423) );
  NANDN U14447 ( .A(n6426), .B(n6427), .Z(n6425) );
  NANDN U14448 ( .A(n6427), .B(n6426), .Z(n6422) );
  XOR U14449 ( .A(n6398), .B(n6428), .Z(n6390) );
  XNOR U14450 ( .A(n6395), .B(n6397), .Z(n6428) );
  AND U14451 ( .A(n6429), .B(n6430), .Z(n6397) );
  NANDN U14452 ( .A(n6431), .B(n6432), .Z(n6430) );
  OR U14453 ( .A(n6433), .B(n6434), .Z(n6432) );
  IV U14454 ( .A(n6435), .Z(n6434) );
  NANDN U14455 ( .A(n6435), .B(n6433), .Z(n6429) );
  AND U14456 ( .A(n6436), .B(n6437), .Z(n6395) );
  NAND U14457 ( .A(n6438), .B(n6439), .Z(n6437) );
  NANDN U14458 ( .A(n6440), .B(n6441), .Z(n6439) );
  NANDN U14459 ( .A(n6441), .B(n6440), .Z(n6436) );
  IV U14460 ( .A(n6442), .Z(n6441) );
  NAND U14461 ( .A(n6443), .B(n6444), .Z(n6398) );
  NANDN U14462 ( .A(n6445), .B(n6446), .Z(n6444) );
  NANDN U14463 ( .A(n6447), .B(n6448), .Z(n6446) );
  NANDN U14464 ( .A(n6448), .B(n6447), .Z(n6443) );
  IV U14465 ( .A(n6449), .Z(n6447) );
  XOR U14466 ( .A(n6424), .B(n6450), .Z(N64818) );
  XNOR U14467 ( .A(n6427), .B(n6426), .Z(n6450) );
  XNOR U14468 ( .A(n6438), .B(n6451), .Z(n6426) );
  XNOR U14469 ( .A(n6442), .B(n6440), .Z(n6451) );
  XOR U14470 ( .A(n6448), .B(n6452), .Z(n6440) );
  XNOR U14471 ( .A(n6445), .B(n6449), .Z(n6452) );
  AND U14472 ( .A(n6453), .B(n6454), .Z(n6449) );
  NAND U14473 ( .A(n6455), .B(n6456), .Z(n6454) );
  NAND U14474 ( .A(n6457), .B(n6458), .Z(n6453) );
  AND U14475 ( .A(n6459), .B(n6460), .Z(n6445) );
  NAND U14476 ( .A(n6461), .B(n6462), .Z(n6460) );
  NAND U14477 ( .A(n6463), .B(n6464), .Z(n6459) );
  NANDN U14478 ( .A(n6465), .B(n6466), .Z(n6448) );
  ANDN U14479 ( .B(n6467), .A(n6468), .Z(n6442) );
  XNOR U14480 ( .A(n6433), .B(n6469), .Z(n6438) );
  XNOR U14481 ( .A(n6431), .B(n6435), .Z(n6469) );
  AND U14482 ( .A(n6470), .B(n6471), .Z(n6435) );
  NAND U14483 ( .A(n6472), .B(n6473), .Z(n6471) );
  NAND U14484 ( .A(n6474), .B(n6475), .Z(n6470) );
  AND U14485 ( .A(n6476), .B(n6477), .Z(n6431) );
  NAND U14486 ( .A(n6478), .B(n6479), .Z(n6477) );
  NAND U14487 ( .A(n6480), .B(n6481), .Z(n6476) );
  AND U14488 ( .A(n6482), .B(n6483), .Z(n6433) );
  NAND U14489 ( .A(n6484), .B(n6485), .Z(n6427) );
  XNOR U14490 ( .A(n6410), .B(n6486), .Z(n6424) );
  XNOR U14491 ( .A(n6414), .B(n6412), .Z(n6486) );
  XOR U14492 ( .A(n6420), .B(n6487), .Z(n6412) );
  XNOR U14493 ( .A(n6417), .B(n6421), .Z(n6487) );
  AND U14494 ( .A(n6488), .B(n6489), .Z(n6421) );
  NAND U14495 ( .A(n6490), .B(n6491), .Z(n6489) );
  NAND U14496 ( .A(n6492), .B(n6493), .Z(n6488) );
  AND U14497 ( .A(n6494), .B(n6495), .Z(n6417) );
  NAND U14498 ( .A(n6496), .B(n6497), .Z(n6495) );
  NAND U14499 ( .A(n6498), .B(n6499), .Z(n6494) );
  NANDN U14500 ( .A(n6500), .B(n6501), .Z(n6420) );
  ANDN U14501 ( .B(n6502), .A(n6503), .Z(n6414) );
  XNOR U14502 ( .A(n6405), .B(n6504), .Z(n6410) );
  XNOR U14503 ( .A(n6403), .B(n6407), .Z(n6504) );
  AND U14504 ( .A(n6505), .B(n6506), .Z(n6407) );
  NAND U14505 ( .A(n6507), .B(n6508), .Z(n6506) );
  NAND U14506 ( .A(n6509), .B(n6510), .Z(n6505) );
  AND U14507 ( .A(n6511), .B(n6512), .Z(n6403) );
  NAND U14508 ( .A(n6513), .B(n6514), .Z(n6512) );
  NAND U14509 ( .A(n6515), .B(n6516), .Z(n6511) );
  AND U14510 ( .A(n6517), .B(n6518), .Z(n6405) );
  XOR U14511 ( .A(n6485), .B(n6484), .Z(N64817) );
  XNOR U14512 ( .A(n6502), .B(n6503), .Z(n6484) );
  XNOR U14513 ( .A(n6517), .B(n6518), .Z(n6503) );
  XOR U14514 ( .A(n6514), .B(n6513), .Z(n6518) );
  XOR U14515 ( .A(y[7812]), .B(x[7812]), .Z(n6513) );
  XOR U14516 ( .A(n6516), .B(n6515), .Z(n6514) );
  XOR U14517 ( .A(y[7814]), .B(x[7814]), .Z(n6515) );
  XOR U14518 ( .A(y[7813]), .B(x[7813]), .Z(n6516) );
  XOR U14519 ( .A(n6508), .B(n6507), .Z(n6517) );
  XOR U14520 ( .A(n6510), .B(n6509), .Z(n6507) );
  XOR U14521 ( .A(y[7811]), .B(x[7811]), .Z(n6509) );
  XOR U14522 ( .A(y[7810]), .B(x[7810]), .Z(n6510) );
  XOR U14523 ( .A(y[7809]), .B(x[7809]), .Z(n6508) );
  XNOR U14524 ( .A(n6501), .B(n6500), .Z(n6502) );
  XNOR U14525 ( .A(n6497), .B(n6496), .Z(n6500) );
  XOR U14526 ( .A(n6499), .B(n6498), .Z(n6496) );
  XOR U14527 ( .A(y[7808]), .B(x[7808]), .Z(n6498) );
  XOR U14528 ( .A(y[7807]), .B(x[7807]), .Z(n6499) );
  XOR U14529 ( .A(y[7806]), .B(x[7806]), .Z(n6497) );
  XOR U14530 ( .A(n6491), .B(n6490), .Z(n6501) );
  XOR U14531 ( .A(n6493), .B(n6492), .Z(n6490) );
  XOR U14532 ( .A(y[7805]), .B(x[7805]), .Z(n6492) );
  XOR U14533 ( .A(y[7804]), .B(x[7804]), .Z(n6493) );
  XOR U14534 ( .A(y[7803]), .B(x[7803]), .Z(n6491) );
  XNOR U14535 ( .A(n6467), .B(n6468), .Z(n6485) );
  XNOR U14536 ( .A(n6482), .B(n6483), .Z(n6468) );
  XOR U14537 ( .A(n6479), .B(n6478), .Z(n6483) );
  XOR U14538 ( .A(y[7800]), .B(x[7800]), .Z(n6478) );
  XOR U14539 ( .A(n6481), .B(n6480), .Z(n6479) );
  XOR U14540 ( .A(y[7802]), .B(x[7802]), .Z(n6480) );
  XOR U14541 ( .A(y[7801]), .B(x[7801]), .Z(n6481) );
  XOR U14542 ( .A(n6473), .B(n6472), .Z(n6482) );
  XOR U14543 ( .A(n6475), .B(n6474), .Z(n6472) );
  XOR U14544 ( .A(y[7799]), .B(x[7799]), .Z(n6474) );
  XOR U14545 ( .A(y[7798]), .B(x[7798]), .Z(n6475) );
  XOR U14546 ( .A(y[7797]), .B(x[7797]), .Z(n6473) );
  XNOR U14547 ( .A(n6466), .B(n6465), .Z(n6467) );
  XNOR U14548 ( .A(n6462), .B(n6461), .Z(n6465) );
  XOR U14549 ( .A(n6464), .B(n6463), .Z(n6461) );
  XOR U14550 ( .A(y[7796]), .B(x[7796]), .Z(n6463) );
  XOR U14551 ( .A(y[7795]), .B(x[7795]), .Z(n6464) );
  XOR U14552 ( .A(y[7794]), .B(x[7794]), .Z(n6462) );
  XOR U14553 ( .A(n6456), .B(n6455), .Z(n6466) );
  XOR U14554 ( .A(n6458), .B(n6457), .Z(n6455) );
  XOR U14555 ( .A(y[7793]), .B(x[7793]), .Z(n6457) );
  XOR U14556 ( .A(y[7792]), .B(x[7792]), .Z(n6458) );
  XOR U14557 ( .A(y[7791]), .B(x[7791]), .Z(n6456) );
  NAND U14558 ( .A(n6519), .B(n6520), .Z(N64808) );
  NAND U14559 ( .A(n6521), .B(n6522), .Z(n6520) );
  NANDN U14560 ( .A(n6523), .B(n6524), .Z(n6522) );
  NANDN U14561 ( .A(n6524), .B(n6523), .Z(n6519) );
  XOR U14562 ( .A(n6523), .B(n6525), .Z(N64807) );
  XNOR U14563 ( .A(n6521), .B(n6524), .Z(n6525) );
  NAND U14564 ( .A(n6526), .B(n6527), .Z(n6524) );
  NAND U14565 ( .A(n6528), .B(n6529), .Z(n6527) );
  NANDN U14566 ( .A(n6530), .B(n6531), .Z(n6529) );
  NANDN U14567 ( .A(n6531), .B(n6530), .Z(n6526) );
  AND U14568 ( .A(n6532), .B(n6533), .Z(n6521) );
  NAND U14569 ( .A(n6534), .B(n6535), .Z(n6533) );
  NANDN U14570 ( .A(n6536), .B(n6537), .Z(n6535) );
  NANDN U14571 ( .A(n6537), .B(n6536), .Z(n6532) );
  IV U14572 ( .A(n6538), .Z(n6537) );
  AND U14573 ( .A(n6539), .B(n6540), .Z(n6523) );
  NAND U14574 ( .A(n6541), .B(n6542), .Z(n6540) );
  NANDN U14575 ( .A(n6543), .B(n6544), .Z(n6542) );
  NANDN U14576 ( .A(n6544), .B(n6543), .Z(n6539) );
  XOR U14577 ( .A(n6536), .B(n6545), .Z(N64806) );
  XNOR U14578 ( .A(n6534), .B(n6538), .Z(n6545) );
  XOR U14579 ( .A(n6531), .B(n6546), .Z(n6538) );
  XNOR U14580 ( .A(n6528), .B(n6530), .Z(n6546) );
  AND U14581 ( .A(n6547), .B(n6548), .Z(n6530) );
  NANDN U14582 ( .A(n6549), .B(n6550), .Z(n6548) );
  OR U14583 ( .A(n6551), .B(n6552), .Z(n6550) );
  IV U14584 ( .A(n6553), .Z(n6552) );
  NANDN U14585 ( .A(n6553), .B(n6551), .Z(n6547) );
  AND U14586 ( .A(n6554), .B(n6555), .Z(n6528) );
  NAND U14587 ( .A(n6556), .B(n6557), .Z(n6555) );
  NANDN U14588 ( .A(n6558), .B(n6559), .Z(n6557) );
  NANDN U14589 ( .A(n6559), .B(n6558), .Z(n6554) );
  IV U14590 ( .A(n6560), .Z(n6559) );
  NAND U14591 ( .A(n6561), .B(n6562), .Z(n6531) );
  NANDN U14592 ( .A(n6563), .B(n6564), .Z(n6562) );
  NANDN U14593 ( .A(n6565), .B(n6566), .Z(n6564) );
  NANDN U14594 ( .A(n6566), .B(n6565), .Z(n6561) );
  IV U14595 ( .A(n6567), .Z(n6565) );
  AND U14596 ( .A(n6568), .B(n6569), .Z(n6534) );
  NAND U14597 ( .A(n6570), .B(n6571), .Z(n6569) );
  NANDN U14598 ( .A(n6572), .B(n6573), .Z(n6571) );
  NANDN U14599 ( .A(n6573), .B(n6572), .Z(n6568) );
  XOR U14600 ( .A(n6544), .B(n6574), .Z(n6536) );
  XNOR U14601 ( .A(n6541), .B(n6543), .Z(n6574) );
  AND U14602 ( .A(n6575), .B(n6576), .Z(n6543) );
  NANDN U14603 ( .A(n6577), .B(n6578), .Z(n6576) );
  OR U14604 ( .A(n6579), .B(n6580), .Z(n6578) );
  IV U14605 ( .A(n6581), .Z(n6580) );
  NANDN U14606 ( .A(n6581), .B(n6579), .Z(n6575) );
  AND U14607 ( .A(n6582), .B(n6583), .Z(n6541) );
  NAND U14608 ( .A(n6584), .B(n6585), .Z(n6583) );
  NANDN U14609 ( .A(n6586), .B(n6587), .Z(n6585) );
  NANDN U14610 ( .A(n6587), .B(n6586), .Z(n6582) );
  IV U14611 ( .A(n6588), .Z(n6587) );
  NAND U14612 ( .A(n6589), .B(n6590), .Z(n6544) );
  NANDN U14613 ( .A(n6591), .B(n6592), .Z(n6590) );
  NANDN U14614 ( .A(n6593), .B(n6594), .Z(n6592) );
  NANDN U14615 ( .A(n6594), .B(n6593), .Z(n6589) );
  IV U14616 ( .A(n6595), .Z(n6593) );
  XOR U14617 ( .A(n6570), .B(n6596), .Z(N64805) );
  XNOR U14618 ( .A(n6573), .B(n6572), .Z(n6596) );
  XNOR U14619 ( .A(n6584), .B(n6597), .Z(n6572) );
  XNOR U14620 ( .A(n6588), .B(n6586), .Z(n6597) );
  XOR U14621 ( .A(n6594), .B(n6598), .Z(n6586) );
  XNOR U14622 ( .A(n6591), .B(n6595), .Z(n6598) );
  AND U14623 ( .A(n6599), .B(n6600), .Z(n6595) );
  NAND U14624 ( .A(n6601), .B(n6602), .Z(n6600) );
  NAND U14625 ( .A(n6603), .B(n6604), .Z(n6599) );
  AND U14626 ( .A(n6605), .B(n6606), .Z(n6591) );
  NAND U14627 ( .A(n6607), .B(n6608), .Z(n6606) );
  NAND U14628 ( .A(n6609), .B(n6610), .Z(n6605) );
  NANDN U14629 ( .A(n6611), .B(n6612), .Z(n6594) );
  ANDN U14630 ( .B(n6613), .A(n6614), .Z(n6588) );
  XNOR U14631 ( .A(n6579), .B(n6615), .Z(n6584) );
  XNOR U14632 ( .A(n6577), .B(n6581), .Z(n6615) );
  AND U14633 ( .A(n6616), .B(n6617), .Z(n6581) );
  NAND U14634 ( .A(n6618), .B(n6619), .Z(n6617) );
  NAND U14635 ( .A(n6620), .B(n6621), .Z(n6616) );
  AND U14636 ( .A(n6622), .B(n6623), .Z(n6577) );
  NAND U14637 ( .A(n6624), .B(n6625), .Z(n6623) );
  NAND U14638 ( .A(n6626), .B(n6627), .Z(n6622) );
  AND U14639 ( .A(n6628), .B(n6629), .Z(n6579) );
  NAND U14640 ( .A(n6630), .B(n6631), .Z(n6573) );
  XNOR U14641 ( .A(n6556), .B(n6632), .Z(n6570) );
  XNOR U14642 ( .A(n6560), .B(n6558), .Z(n6632) );
  XOR U14643 ( .A(n6566), .B(n6633), .Z(n6558) );
  XNOR U14644 ( .A(n6563), .B(n6567), .Z(n6633) );
  AND U14645 ( .A(n6634), .B(n6635), .Z(n6567) );
  NAND U14646 ( .A(n6636), .B(n6637), .Z(n6635) );
  NAND U14647 ( .A(n6638), .B(n6639), .Z(n6634) );
  AND U14648 ( .A(n6640), .B(n6641), .Z(n6563) );
  NAND U14649 ( .A(n6642), .B(n6643), .Z(n6641) );
  NAND U14650 ( .A(n6644), .B(n6645), .Z(n6640) );
  NANDN U14651 ( .A(n6646), .B(n6647), .Z(n6566) );
  ANDN U14652 ( .B(n6648), .A(n6649), .Z(n6560) );
  XNOR U14653 ( .A(n6551), .B(n6650), .Z(n6556) );
  XNOR U14654 ( .A(n6549), .B(n6553), .Z(n6650) );
  AND U14655 ( .A(n6651), .B(n6652), .Z(n6553) );
  NAND U14656 ( .A(n6653), .B(n6654), .Z(n6652) );
  NAND U14657 ( .A(n6655), .B(n6656), .Z(n6651) );
  AND U14658 ( .A(n6657), .B(n6658), .Z(n6549) );
  NAND U14659 ( .A(n6659), .B(n6660), .Z(n6658) );
  NAND U14660 ( .A(n6661), .B(n6662), .Z(n6657) );
  AND U14661 ( .A(n6663), .B(n6664), .Z(n6551) );
  XOR U14662 ( .A(n6631), .B(n6630), .Z(N64804) );
  XNOR U14663 ( .A(n6648), .B(n6649), .Z(n6630) );
  XNOR U14664 ( .A(n6663), .B(n6664), .Z(n6649) );
  XOR U14665 ( .A(n6660), .B(n6659), .Z(n6664) );
  XOR U14666 ( .A(y[7788]), .B(x[7788]), .Z(n6659) );
  XOR U14667 ( .A(n6662), .B(n6661), .Z(n6660) );
  XOR U14668 ( .A(y[7790]), .B(x[7790]), .Z(n6661) );
  XOR U14669 ( .A(y[7789]), .B(x[7789]), .Z(n6662) );
  XOR U14670 ( .A(n6654), .B(n6653), .Z(n6663) );
  XOR U14671 ( .A(n6656), .B(n6655), .Z(n6653) );
  XOR U14672 ( .A(y[7787]), .B(x[7787]), .Z(n6655) );
  XOR U14673 ( .A(y[7786]), .B(x[7786]), .Z(n6656) );
  XOR U14674 ( .A(y[7785]), .B(x[7785]), .Z(n6654) );
  XNOR U14675 ( .A(n6647), .B(n6646), .Z(n6648) );
  XNOR U14676 ( .A(n6643), .B(n6642), .Z(n6646) );
  XOR U14677 ( .A(n6645), .B(n6644), .Z(n6642) );
  XOR U14678 ( .A(y[7784]), .B(x[7784]), .Z(n6644) );
  XOR U14679 ( .A(y[7783]), .B(x[7783]), .Z(n6645) );
  XOR U14680 ( .A(y[7782]), .B(x[7782]), .Z(n6643) );
  XOR U14681 ( .A(n6637), .B(n6636), .Z(n6647) );
  XOR U14682 ( .A(n6639), .B(n6638), .Z(n6636) );
  XOR U14683 ( .A(y[7781]), .B(x[7781]), .Z(n6638) );
  XOR U14684 ( .A(y[7780]), .B(x[7780]), .Z(n6639) );
  XOR U14685 ( .A(y[7779]), .B(x[7779]), .Z(n6637) );
  XNOR U14686 ( .A(n6613), .B(n6614), .Z(n6631) );
  XNOR U14687 ( .A(n6628), .B(n6629), .Z(n6614) );
  XOR U14688 ( .A(n6625), .B(n6624), .Z(n6629) );
  XOR U14689 ( .A(y[7776]), .B(x[7776]), .Z(n6624) );
  XOR U14690 ( .A(n6627), .B(n6626), .Z(n6625) );
  XOR U14691 ( .A(y[7778]), .B(x[7778]), .Z(n6626) );
  XOR U14692 ( .A(y[7777]), .B(x[7777]), .Z(n6627) );
  XOR U14693 ( .A(n6619), .B(n6618), .Z(n6628) );
  XOR U14694 ( .A(n6621), .B(n6620), .Z(n6618) );
  XOR U14695 ( .A(y[7775]), .B(x[7775]), .Z(n6620) );
  XOR U14696 ( .A(y[7774]), .B(x[7774]), .Z(n6621) );
  XOR U14697 ( .A(y[7773]), .B(x[7773]), .Z(n6619) );
  XNOR U14698 ( .A(n6612), .B(n6611), .Z(n6613) );
  XNOR U14699 ( .A(n6608), .B(n6607), .Z(n6611) );
  XOR U14700 ( .A(n6610), .B(n6609), .Z(n6607) );
  XOR U14701 ( .A(y[7772]), .B(x[7772]), .Z(n6609) );
  XOR U14702 ( .A(y[7771]), .B(x[7771]), .Z(n6610) );
  XOR U14703 ( .A(y[7770]), .B(x[7770]), .Z(n6608) );
  XOR U14704 ( .A(n6602), .B(n6601), .Z(n6612) );
  XOR U14705 ( .A(n6604), .B(n6603), .Z(n6601) );
  XOR U14706 ( .A(y[7769]), .B(x[7769]), .Z(n6603) );
  XOR U14707 ( .A(y[7768]), .B(x[7768]), .Z(n6604) );
  XOR U14708 ( .A(y[7767]), .B(x[7767]), .Z(n6602) );
  NAND U14709 ( .A(n6665), .B(n6666), .Z(N64795) );
  NAND U14710 ( .A(n6667), .B(n6668), .Z(n6666) );
  NANDN U14711 ( .A(n6669), .B(n6670), .Z(n6668) );
  NANDN U14712 ( .A(n6670), .B(n6669), .Z(n6665) );
  XOR U14713 ( .A(n6669), .B(n6671), .Z(N64794) );
  XNOR U14714 ( .A(n6667), .B(n6670), .Z(n6671) );
  NAND U14715 ( .A(n6672), .B(n6673), .Z(n6670) );
  NAND U14716 ( .A(n6674), .B(n6675), .Z(n6673) );
  NANDN U14717 ( .A(n6676), .B(n6677), .Z(n6675) );
  NANDN U14718 ( .A(n6677), .B(n6676), .Z(n6672) );
  AND U14719 ( .A(n6678), .B(n6679), .Z(n6667) );
  NAND U14720 ( .A(n6680), .B(n6681), .Z(n6679) );
  NANDN U14721 ( .A(n6682), .B(n6683), .Z(n6681) );
  NANDN U14722 ( .A(n6683), .B(n6682), .Z(n6678) );
  IV U14723 ( .A(n6684), .Z(n6683) );
  AND U14724 ( .A(n6685), .B(n6686), .Z(n6669) );
  NAND U14725 ( .A(n6687), .B(n6688), .Z(n6686) );
  NANDN U14726 ( .A(n6689), .B(n6690), .Z(n6688) );
  NANDN U14727 ( .A(n6690), .B(n6689), .Z(n6685) );
  XOR U14728 ( .A(n6682), .B(n6691), .Z(N64793) );
  XNOR U14729 ( .A(n6680), .B(n6684), .Z(n6691) );
  XOR U14730 ( .A(n6677), .B(n6692), .Z(n6684) );
  XNOR U14731 ( .A(n6674), .B(n6676), .Z(n6692) );
  AND U14732 ( .A(n6693), .B(n6694), .Z(n6676) );
  NANDN U14733 ( .A(n6695), .B(n6696), .Z(n6694) );
  OR U14734 ( .A(n6697), .B(n6698), .Z(n6696) );
  IV U14735 ( .A(n6699), .Z(n6698) );
  NANDN U14736 ( .A(n6699), .B(n6697), .Z(n6693) );
  AND U14737 ( .A(n6700), .B(n6701), .Z(n6674) );
  NAND U14738 ( .A(n6702), .B(n6703), .Z(n6701) );
  NANDN U14739 ( .A(n6704), .B(n6705), .Z(n6703) );
  NANDN U14740 ( .A(n6705), .B(n6704), .Z(n6700) );
  IV U14741 ( .A(n6706), .Z(n6705) );
  NAND U14742 ( .A(n6707), .B(n6708), .Z(n6677) );
  NANDN U14743 ( .A(n6709), .B(n6710), .Z(n6708) );
  NANDN U14744 ( .A(n6711), .B(n6712), .Z(n6710) );
  NANDN U14745 ( .A(n6712), .B(n6711), .Z(n6707) );
  IV U14746 ( .A(n6713), .Z(n6711) );
  AND U14747 ( .A(n6714), .B(n6715), .Z(n6680) );
  NAND U14748 ( .A(n6716), .B(n6717), .Z(n6715) );
  NANDN U14749 ( .A(n6718), .B(n6719), .Z(n6717) );
  NANDN U14750 ( .A(n6719), .B(n6718), .Z(n6714) );
  XOR U14751 ( .A(n6690), .B(n6720), .Z(n6682) );
  XNOR U14752 ( .A(n6687), .B(n6689), .Z(n6720) );
  AND U14753 ( .A(n6721), .B(n6722), .Z(n6689) );
  NANDN U14754 ( .A(n6723), .B(n6724), .Z(n6722) );
  OR U14755 ( .A(n6725), .B(n6726), .Z(n6724) );
  IV U14756 ( .A(n6727), .Z(n6726) );
  NANDN U14757 ( .A(n6727), .B(n6725), .Z(n6721) );
  AND U14758 ( .A(n6728), .B(n6729), .Z(n6687) );
  NAND U14759 ( .A(n6730), .B(n6731), .Z(n6729) );
  NANDN U14760 ( .A(n6732), .B(n6733), .Z(n6731) );
  NANDN U14761 ( .A(n6733), .B(n6732), .Z(n6728) );
  IV U14762 ( .A(n6734), .Z(n6733) );
  NAND U14763 ( .A(n6735), .B(n6736), .Z(n6690) );
  NANDN U14764 ( .A(n6737), .B(n6738), .Z(n6736) );
  NANDN U14765 ( .A(n6739), .B(n6740), .Z(n6738) );
  NANDN U14766 ( .A(n6740), .B(n6739), .Z(n6735) );
  IV U14767 ( .A(n6741), .Z(n6739) );
  XOR U14768 ( .A(n6716), .B(n6742), .Z(N64792) );
  XNOR U14769 ( .A(n6719), .B(n6718), .Z(n6742) );
  XNOR U14770 ( .A(n6730), .B(n6743), .Z(n6718) );
  XNOR U14771 ( .A(n6734), .B(n6732), .Z(n6743) );
  XOR U14772 ( .A(n6740), .B(n6744), .Z(n6732) );
  XNOR U14773 ( .A(n6737), .B(n6741), .Z(n6744) );
  AND U14774 ( .A(n6745), .B(n6746), .Z(n6741) );
  NAND U14775 ( .A(n6747), .B(n6748), .Z(n6746) );
  NAND U14776 ( .A(n6749), .B(n6750), .Z(n6745) );
  AND U14777 ( .A(n6751), .B(n6752), .Z(n6737) );
  NAND U14778 ( .A(n6753), .B(n6754), .Z(n6752) );
  NAND U14779 ( .A(n6755), .B(n6756), .Z(n6751) );
  NANDN U14780 ( .A(n6757), .B(n6758), .Z(n6740) );
  ANDN U14781 ( .B(n6759), .A(n6760), .Z(n6734) );
  XNOR U14782 ( .A(n6725), .B(n6761), .Z(n6730) );
  XNOR U14783 ( .A(n6723), .B(n6727), .Z(n6761) );
  AND U14784 ( .A(n6762), .B(n6763), .Z(n6727) );
  NAND U14785 ( .A(n6764), .B(n6765), .Z(n6763) );
  NAND U14786 ( .A(n6766), .B(n6767), .Z(n6762) );
  AND U14787 ( .A(n6768), .B(n6769), .Z(n6723) );
  NAND U14788 ( .A(n6770), .B(n6771), .Z(n6769) );
  NAND U14789 ( .A(n6772), .B(n6773), .Z(n6768) );
  AND U14790 ( .A(n6774), .B(n6775), .Z(n6725) );
  NAND U14791 ( .A(n6776), .B(n6777), .Z(n6719) );
  XNOR U14792 ( .A(n6702), .B(n6778), .Z(n6716) );
  XNOR U14793 ( .A(n6706), .B(n6704), .Z(n6778) );
  XOR U14794 ( .A(n6712), .B(n6779), .Z(n6704) );
  XNOR U14795 ( .A(n6709), .B(n6713), .Z(n6779) );
  AND U14796 ( .A(n6780), .B(n6781), .Z(n6713) );
  NAND U14797 ( .A(n6782), .B(n6783), .Z(n6781) );
  NAND U14798 ( .A(n6784), .B(n6785), .Z(n6780) );
  AND U14799 ( .A(n6786), .B(n6787), .Z(n6709) );
  NAND U14800 ( .A(n6788), .B(n6789), .Z(n6787) );
  NAND U14801 ( .A(n6790), .B(n6791), .Z(n6786) );
  NANDN U14802 ( .A(n6792), .B(n6793), .Z(n6712) );
  ANDN U14803 ( .B(n6794), .A(n6795), .Z(n6706) );
  XNOR U14804 ( .A(n6697), .B(n6796), .Z(n6702) );
  XNOR U14805 ( .A(n6695), .B(n6699), .Z(n6796) );
  AND U14806 ( .A(n6797), .B(n6798), .Z(n6699) );
  NAND U14807 ( .A(n6799), .B(n6800), .Z(n6798) );
  NAND U14808 ( .A(n6801), .B(n6802), .Z(n6797) );
  AND U14809 ( .A(n6803), .B(n6804), .Z(n6695) );
  NAND U14810 ( .A(n6805), .B(n6806), .Z(n6804) );
  NAND U14811 ( .A(n6807), .B(n6808), .Z(n6803) );
  AND U14812 ( .A(n6809), .B(n6810), .Z(n6697) );
  XOR U14813 ( .A(n6777), .B(n6776), .Z(N64791) );
  XNOR U14814 ( .A(n6794), .B(n6795), .Z(n6776) );
  XNOR U14815 ( .A(n6809), .B(n6810), .Z(n6795) );
  XOR U14816 ( .A(n6806), .B(n6805), .Z(n6810) );
  XOR U14817 ( .A(y[7764]), .B(x[7764]), .Z(n6805) );
  XOR U14818 ( .A(n6808), .B(n6807), .Z(n6806) );
  XOR U14819 ( .A(y[7766]), .B(x[7766]), .Z(n6807) );
  XOR U14820 ( .A(y[7765]), .B(x[7765]), .Z(n6808) );
  XOR U14821 ( .A(n6800), .B(n6799), .Z(n6809) );
  XOR U14822 ( .A(n6802), .B(n6801), .Z(n6799) );
  XOR U14823 ( .A(y[7763]), .B(x[7763]), .Z(n6801) );
  XOR U14824 ( .A(y[7762]), .B(x[7762]), .Z(n6802) );
  XOR U14825 ( .A(y[7761]), .B(x[7761]), .Z(n6800) );
  XNOR U14826 ( .A(n6793), .B(n6792), .Z(n6794) );
  XNOR U14827 ( .A(n6789), .B(n6788), .Z(n6792) );
  XOR U14828 ( .A(n6791), .B(n6790), .Z(n6788) );
  XOR U14829 ( .A(y[7760]), .B(x[7760]), .Z(n6790) );
  XOR U14830 ( .A(y[7759]), .B(x[7759]), .Z(n6791) );
  XOR U14831 ( .A(y[7758]), .B(x[7758]), .Z(n6789) );
  XOR U14832 ( .A(n6783), .B(n6782), .Z(n6793) );
  XOR U14833 ( .A(n6785), .B(n6784), .Z(n6782) );
  XOR U14834 ( .A(y[7757]), .B(x[7757]), .Z(n6784) );
  XOR U14835 ( .A(y[7756]), .B(x[7756]), .Z(n6785) );
  XOR U14836 ( .A(y[7755]), .B(x[7755]), .Z(n6783) );
  XNOR U14837 ( .A(n6759), .B(n6760), .Z(n6777) );
  XNOR U14838 ( .A(n6774), .B(n6775), .Z(n6760) );
  XOR U14839 ( .A(n6771), .B(n6770), .Z(n6775) );
  XOR U14840 ( .A(y[7752]), .B(x[7752]), .Z(n6770) );
  XOR U14841 ( .A(n6773), .B(n6772), .Z(n6771) );
  XOR U14842 ( .A(y[7754]), .B(x[7754]), .Z(n6772) );
  XOR U14843 ( .A(y[7753]), .B(x[7753]), .Z(n6773) );
  XOR U14844 ( .A(n6765), .B(n6764), .Z(n6774) );
  XOR U14845 ( .A(n6767), .B(n6766), .Z(n6764) );
  XOR U14846 ( .A(y[7751]), .B(x[7751]), .Z(n6766) );
  XOR U14847 ( .A(y[7750]), .B(x[7750]), .Z(n6767) );
  XOR U14848 ( .A(y[7749]), .B(x[7749]), .Z(n6765) );
  XNOR U14849 ( .A(n6758), .B(n6757), .Z(n6759) );
  XNOR U14850 ( .A(n6754), .B(n6753), .Z(n6757) );
  XOR U14851 ( .A(n6756), .B(n6755), .Z(n6753) );
  XOR U14852 ( .A(y[7748]), .B(x[7748]), .Z(n6755) );
  XOR U14853 ( .A(y[7747]), .B(x[7747]), .Z(n6756) );
  XOR U14854 ( .A(y[7746]), .B(x[7746]), .Z(n6754) );
  XOR U14855 ( .A(n6748), .B(n6747), .Z(n6758) );
  XOR U14856 ( .A(n6750), .B(n6749), .Z(n6747) );
  XOR U14857 ( .A(y[7745]), .B(x[7745]), .Z(n6749) );
  XOR U14858 ( .A(y[7744]), .B(x[7744]), .Z(n6750) );
  XOR U14859 ( .A(y[7743]), .B(x[7743]), .Z(n6748) );
  NAND U14860 ( .A(n6811), .B(n6812), .Z(N64782) );
  NAND U14861 ( .A(n6813), .B(n6814), .Z(n6812) );
  NANDN U14862 ( .A(n6815), .B(n6816), .Z(n6814) );
  NANDN U14863 ( .A(n6816), .B(n6815), .Z(n6811) );
  XOR U14864 ( .A(n6815), .B(n6817), .Z(N64781) );
  XNOR U14865 ( .A(n6813), .B(n6816), .Z(n6817) );
  NAND U14866 ( .A(n6818), .B(n6819), .Z(n6816) );
  NAND U14867 ( .A(n6820), .B(n6821), .Z(n6819) );
  NANDN U14868 ( .A(n6822), .B(n6823), .Z(n6821) );
  NANDN U14869 ( .A(n6823), .B(n6822), .Z(n6818) );
  AND U14870 ( .A(n6824), .B(n6825), .Z(n6813) );
  NAND U14871 ( .A(n6826), .B(n6827), .Z(n6825) );
  NANDN U14872 ( .A(n6828), .B(n6829), .Z(n6827) );
  NANDN U14873 ( .A(n6829), .B(n6828), .Z(n6824) );
  IV U14874 ( .A(n6830), .Z(n6829) );
  AND U14875 ( .A(n6831), .B(n6832), .Z(n6815) );
  NAND U14876 ( .A(n6833), .B(n6834), .Z(n6832) );
  NANDN U14877 ( .A(n6835), .B(n6836), .Z(n6834) );
  NANDN U14878 ( .A(n6836), .B(n6835), .Z(n6831) );
  XOR U14879 ( .A(n6828), .B(n6837), .Z(N64780) );
  XNOR U14880 ( .A(n6826), .B(n6830), .Z(n6837) );
  XOR U14881 ( .A(n6823), .B(n6838), .Z(n6830) );
  XNOR U14882 ( .A(n6820), .B(n6822), .Z(n6838) );
  AND U14883 ( .A(n6839), .B(n6840), .Z(n6822) );
  NANDN U14884 ( .A(n6841), .B(n6842), .Z(n6840) );
  OR U14885 ( .A(n6843), .B(n6844), .Z(n6842) );
  IV U14886 ( .A(n6845), .Z(n6844) );
  NANDN U14887 ( .A(n6845), .B(n6843), .Z(n6839) );
  AND U14888 ( .A(n6846), .B(n6847), .Z(n6820) );
  NAND U14889 ( .A(n6848), .B(n6849), .Z(n6847) );
  NANDN U14890 ( .A(n6850), .B(n6851), .Z(n6849) );
  NANDN U14891 ( .A(n6851), .B(n6850), .Z(n6846) );
  IV U14892 ( .A(n6852), .Z(n6851) );
  NAND U14893 ( .A(n6853), .B(n6854), .Z(n6823) );
  NANDN U14894 ( .A(n6855), .B(n6856), .Z(n6854) );
  NANDN U14895 ( .A(n6857), .B(n6858), .Z(n6856) );
  NANDN U14896 ( .A(n6858), .B(n6857), .Z(n6853) );
  IV U14897 ( .A(n6859), .Z(n6857) );
  AND U14898 ( .A(n6860), .B(n6861), .Z(n6826) );
  NAND U14899 ( .A(n6862), .B(n6863), .Z(n6861) );
  NANDN U14900 ( .A(n6864), .B(n6865), .Z(n6863) );
  NANDN U14901 ( .A(n6865), .B(n6864), .Z(n6860) );
  XOR U14902 ( .A(n6836), .B(n6866), .Z(n6828) );
  XNOR U14903 ( .A(n6833), .B(n6835), .Z(n6866) );
  AND U14904 ( .A(n6867), .B(n6868), .Z(n6835) );
  NANDN U14905 ( .A(n6869), .B(n6870), .Z(n6868) );
  OR U14906 ( .A(n6871), .B(n6872), .Z(n6870) );
  IV U14907 ( .A(n6873), .Z(n6872) );
  NANDN U14908 ( .A(n6873), .B(n6871), .Z(n6867) );
  AND U14909 ( .A(n6874), .B(n6875), .Z(n6833) );
  NAND U14910 ( .A(n6876), .B(n6877), .Z(n6875) );
  NANDN U14911 ( .A(n6878), .B(n6879), .Z(n6877) );
  NANDN U14912 ( .A(n6879), .B(n6878), .Z(n6874) );
  IV U14913 ( .A(n6880), .Z(n6879) );
  NAND U14914 ( .A(n6881), .B(n6882), .Z(n6836) );
  NANDN U14915 ( .A(n6883), .B(n6884), .Z(n6882) );
  NANDN U14916 ( .A(n6885), .B(n6886), .Z(n6884) );
  NANDN U14917 ( .A(n6886), .B(n6885), .Z(n6881) );
  IV U14918 ( .A(n6887), .Z(n6885) );
  XOR U14919 ( .A(n6862), .B(n6888), .Z(N64779) );
  XNOR U14920 ( .A(n6865), .B(n6864), .Z(n6888) );
  XNOR U14921 ( .A(n6876), .B(n6889), .Z(n6864) );
  XNOR U14922 ( .A(n6880), .B(n6878), .Z(n6889) );
  XOR U14923 ( .A(n6886), .B(n6890), .Z(n6878) );
  XNOR U14924 ( .A(n6883), .B(n6887), .Z(n6890) );
  AND U14925 ( .A(n6891), .B(n6892), .Z(n6887) );
  NAND U14926 ( .A(n6893), .B(n6894), .Z(n6892) );
  NAND U14927 ( .A(n6895), .B(n6896), .Z(n6891) );
  AND U14928 ( .A(n6897), .B(n6898), .Z(n6883) );
  NAND U14929 ( .A(n6899), .B(n6900), .Z(n6898) );
  NAND U14930 ( .A(n6901), .B(n6902), .Z(n6897) );
  NANDN U14931 ( .A(n6903), .B(n6904), .Z(n6886) );
  ANDN U14932 ( .B(n6905), .A(n6906), .Z(n6880) );
  XNOR U14933 ( .A(n6871), .B(n6907), .Z(n6876) );
  XNOR U14934 ( .A(n6869), .B(n6873), .Z(n6907) );
  AND U14935 ( .A(n6908), .B(n6909), .Z(n6873) );
  NAND U14936 ( .A(n6910), .B(n6911), .Z(n6909) );
  NAND U14937 ( .A(n6912), .B(n6913), .Z(n6908) );
  AND U14938 ( .A(n6914), .B(n6915), .Z(n6869) );
  NAND U14939 ( .A(n6916), .B(n6917), .Z(n6915) );
  NAND U14940 ( .A(n6918), .B(n6919), .Z(n6914) );
  AND U14941 ( .A(n6920), .B(n6921), .Z(n6871) );
  NAND U14942 ( .A(n6922), .B(n6923), .Z(n6865) );
  XNOR U14943 ( .A(n6848), .B(n6924), .Z(n6862) );
  XNOR U14944 ( .A(n6852), .B(n6850), .Z(n6924) );
  XOR U14945 ( .A(n6858), .B(n6925), .Z(n6850) );
  XNOR U14946 ( .A(n6855), .B(n6859), .Z(n6925) );
  AND U14947 ( .A(n6926), .B(n6927), .Z(n6859) );
  NAND U14948 ( .A(n6928), .B(n6929), .Z(n6927) );
  NAND U14949 ( .A(n6930), .B(n6931), .Z(n6926) );
  AND U14950 ( .A(n6932), .B(n6933), .Z(n6855) );
  NAND U14951 ( .A(n6934), .B(n6935), .Z(n6933) );
  NAND U14952 ( .A(n6936), .B(n6937), .Z(n6932) );
  NANDN U14953 ( .A(n6938), .B(n6939), .Z(n6858) );
  ANDN U14954 ( .B(n6940), .A(n6941), .Z(n6852) );
  XNOR U14955 ( .A(n6843), .B(n6942), .Z(n6848) );
  XNOR U14956 ( .A(n6841), .B(n6845), .Z(n6942) );
  AND U14957 ( .A(n6943), .B(n6944), .Z(n6845) );
  NAND U14958 ( .A(n6945), .B(n6946), .Z(n6944) );
  NAND U14959 ( .A(n6947), .B(n6948), .Z(n6943) );
  AND U14960 ( .A(n6949), .B(n6950), .Z(n6841) );
  NAND U14961 ( .A(n6951), .B(n6952), .Z(n6950) );
  NAND U14962 ( .A(n6953), .B(n6954), .Z(n6949) );
  AND U14963 ( .A(n6955), .B(n6956), .Z(n6843) );
  XOR U14964 ( .A(n6923), .B(n6922), .Z(N64778) );
  XNOR U14965 ( .A(n6940), .B(n6941), .Z(n6922) );
  XNOR U14966 ( .A(n6955), .B(n6956), .Z(n6941) );
  XOR U14967 ( .A(n6952), .B(n6951), .Z(n6956) );
  XOR U14968 ( .A(y[7740]), .B(x[7740]), .Z(n6951) );
  XOR U14969 ( .A(n6954), .B(n6953), .Z(n6952) );
  XOR U14970 ( .A(y[7742]), .B(x[7742]), .Z(n6953) );
  XOR U14971 ( .A(y[7741]), .B(x[7741]), .Z(n6954) );
  XOR U14972 ( .A(n6946), .B(n6945), .Z(n6955) );
  XOR U14973 ( .A(n6948), .B(n6947), .Z(n6945) );
  XOR U14974 ( .A(y[7739]), .B(x[7739]), .Z(n6947) );
  XOR U14975 ( .A(y[7738]), .B(x[7738]), .Z(n6948) );
  XOR U14976 ( .A(y[7737]), .B(x[7737]), .Z(n6946) );
  XNOR U14977 ( .A(n6939), .B(n6938), .Z(n6940) );
  XNOR U14978 ( .A(n6935), .B(n6934), .Z(n6938) );
  XOR U14979 ( .A(n6937), .B(n6936), .Z(n6934) );
  XOR U14980 ( .A(y[7736]), .B(x[7736]), .Z(n6936) );
  XOR U14981 ( .A(y[7735]), .B(x[7735]), .Z(n6937) );
  XOR U14982 ( .A(y[7734]), .B(x[7734]), .Z(n6935) );
  XOR U14983 ( .A(n6929), .B(n6928), .Z(n6939) );
  XOR U14984 ( .A(n6931), .B(n6930), .Z(n6928) );
  XOR U14985 ( .A(y[7733]), .B(x[7733]), .Z(n6930) );
  XOR U14986 ( .A(y[7732]), .B(x[7732]), .Z(n6931) );
  XOR U14987 ( .A(y[7731]), .B(x[7731]), .Z(n6929) );
  XNOR U14988 ( .A(n6905), .B(n6906), .Z(n6923) );
  XNOR U14989 ( .A(n6920), .B(n6921), .Z(n6906) );
  XOR U14990 ( .A(n6917), .B(n6916), .Z(n6921) );
  XOR U14991 ( .A(y[7728]), .B(x[7728]), .Z(n6916) );
  XOR U14992 ( .A(n6919), .B(n6918), .Z(n6917) );
  XOR U14993 ( .A(y[7730]), .B(x[7730]), .Z(n6918) );
  XOR U14994 ( .A(y[7729]), .B(x[7729]), .Z(n6919) );
  XOR U14995 ( .A(n6911), .B(n6910), .Z(n6920) );
  XOR U14996 ( .A(n6913), .B(n6912), .Z(n6910) );
  XOR U14997 ( .A(y[7727]), .B(x[7727]), .Z(n6912) );
  XOR U14998 ( .A(y[7726]), .B(x[7726]), .Z(n6913) );
  XOR U14999 ( .A(y[7725]), .B(x[7725]), .Z(n6911) );
  XNOR U15000 ( .A(n6904), .B(n6903), .Z(n6905) );
  XNOR U15001 ( .A(n6900), .B(n6899), .Z(n6903) );
  XOR U15002 ( .A(n6902), .B(n6901), .Z(n6899) );
  XOR U15003 ( .A(y[7724]), .B(x[7724]), .Z(n6901) );
  XOR U15004 ( .A(y[7723]), .B(x[7723]), .Z(n6902) );
  XOR U15005 ( .A(y[7722]), .B(x[7722]), .Z(n6900) );
  XOR U15006 ( .A(n6894), .B(n6893), .Z(n6904) );
  XOR U15007 ( .A(n6896), .B(n6895), .Z(n6893) );
  XOR U15008 ( .A(y[7721]), .B(x[7721]), .Z(n6895) );
  XOR U15009 ( .A(y[7720]), .B(x[7720]), .Z(n6896) );
  XOR U15010 ( .A(y[7719]), .B(x[7719]), .Z(n6894) );
  NAND U15011 ( .A(n6957), .B(n6958), .Z(N64769) );
  NAND U15012 ( .A(n6959), .B(n6960), .Z(n6958) );
  NANDN U15013 ( .A(n6961), .B(n6962), .Z(n6960) );
  NANDN U15014 ( .A(n6962), .B(n6961), .Z(n6957) );
  XOR U15015 ( .A(n6961), .B(n6963), .Z(N64768) );
  XNOR U15016 ( .A(n6959), .B(n6962), .Z(n6963) );
  NAND U15017 ( .A(n6964), .B(n6965), .Z(n6962) );
  NAND U15018 ( .A(n6966), .B(n6967), .Z(n6965) );
  NANDN U15019 ( .A(n6968), .B(n6969), .Z(n6967) );
  NANDN U15020 ( .A(n6969), .B(n6968), .Z(n6964) );
  AND U15021 ( .A(n6970), .B(n6971), .Z(n6959) );
  NAND U15022 ( .A(n6972), .B(n6973), .Z(n6971) );
  NANDN U15023 ( .A(n6974), .B(n6975), .Z(n6973) );
  NANDN U15024 ( .A(n6975), .B(n6974), .Z(n6970) );
  IV U15025 ( .A(n6976), .Z(n6975) );
  AND U15026 ( .A(n6977), .B(n6978), .Z(n6961) );
  NAND U15027 ( .A(n6979), .B(n6980), .Z(n6978) );
  NANDN U15028 ( .A(n6981), .B(n6982), .Z(n6980) );
  NANDN U15029 ( .A(n6982), .B(n6981), .Z(n6977) );
  XOR U15030 ( .A(n6974), .B(n6983), .Z(N64767) );
  XNOR U15031 ( .A(n6972), .B(n6976), .Z(n6983) );
  XOR U15032 ( .A(n6969), .B(n6984), .Z(n6976) );
  XNOR U15033 ( .A(n6966), .B(n6968), .Z(n6984) );
  AND U15034 ( .A(n6985), .B(n6986), .Z(n6968) );
  NANDN U15035 ( .A(n6987), .B(n6988), .Z(n6986) );
  OR U15036 ( .A(n6989), .B(n6990), .Z(n6988) );
  IV U15037 ( .A(n6991), .Z(n6990) );
  NANDN U15038 ( .A(n6991), .B(n6989), .Z(n6985) );
  AND U15039 ( .A(n6992), .B(n6993), .Z(n6966) );
  NAND U15040 ( .A(n6994), .B(n6995), .Z(n6993) );
  NANDN U15041 ( .A(n6996), .B(n6997), .Z(n6995) );
  NANDN U15042 ( .A(n6997), .B(n6996), .Z(n6992) );
  IV U15043 ( .A(n6998), .Z(n6997) );
  NAND U15044 ( .A(n6999), .B(n7000), .Z(n6969) );
  NANDN U15045 ( .A(n7001), .B(n7002), .Z(n7000) );
  NANDN U15046 ( .A(n7003), .B(n7004), .Z(n7002) );
  NANDN U15047 ( .A(n7004), .B(n7003), .Z(n6999) );
  IV U15048 ( .A(n7005), .Z(n7003) );
  AND U15049 ( .A(n7006), .B(n7007), .Z(n6972) );
  NAND U15050 ( .A(n7008), .B(n7009), .Z(n7007) );
  NANDN U15051 ( .A(n7010), .B(n7011), .Z(n7009) );
  NANDN U15052 ( .A(n7011), .B(n7010), .Z(n7006) );
  XOR U15053 ( .A(n6982), .B(n7012), .Z(n6974) );
  XNOR U15054 ( .A(n6979), .B(n6981), .Z(n7012) );
  AND U15055 ( .A(n7013), .B(n7014), .Z(n6981) );
  NANDN U15056 ( .A(n7015), .B(n7016), .Z(n7014) );
  OR U15057 ( .A(n7017), .B(n7018), .Z(n7016) );
  IV U15058 ( .A(n7019), .Z(n7018) );
  NANDN U15059 ( .A(n7019), .B(n7017), .Z(n7013) );
  AND U15060 ( .A(n7020), .B(n7021), .Z(n6979) );
  NAND U15061 ( .A(n7022), .B(n7023), .Z(n7021) );
  NANDN U15062 ( .A(n7024), .B(n7025), .Z(n7023) );
  NANDN U15063 ( .A(n7025), .B(n7024), .Z(n7020) );
  IV U15064 ( .A(n7026), .Z(n7025) );
  NAND U15065 ( .A(n7027), .B(n7028), .Z(n6982) );
  NANDN U15066 ( .A(n7029), .B(n7030), .Z(n7028) );
  NANDN U15067 ( .A(n7031), .B(n7032), .Z(n7030) );
  NANDN U15068 ( .A(n7032), .B(n7031), .Z(n7027) );
  IV U15069 ( .A(n7033), .Z(n7031) );
  XOR U15070 ( .A(n7008), .B(n7034), .Z(N64766) );
  XNOR U15071 ( .A(n7011), .B(n7010), .Z(n7034) );
  XNOR U15072 ( .A(n7022), .B(n7035), .Z(n7010) );
  XNOR U15073 ( .A(n7026), .B(n7024), .Z(n7035) );
  XOR U15074 ( .A(n7032), .B(n7036), .Z(n7024) );
  XNOR U15075 ( .A(n7029), .B(n7033), .Z(n7036) );
  AND U15076 ( .A(n7037), .B(n7038), .Z(n7033) );
  NAND U15077 ( .A(n7039), .B(n7040), .Z(n7038) );
  NAND U15078 ( .A(n7041), .B(n7042), .Z(n7037) );
  AND U15079 ( .A(n7043), .B(n7044), .Z(n7029) );
  NAND U15080 ( .A(n7045), .B(n7046), .Z(n7044) );
  NAND U15081 ( .A(n7047), .B(n7048), .Z(n7043) );
  NANDN U15082 ( .A(n7049), .B(n7050), .Z(n7032) );
  ANDN U15083 ( .B(n7051), .A(n7052), .Z(n7026) );
  XNOR U15084 ( .A(n7017), .B(n7053), .Z(n7022) );
  XNOR U15085 ( .A(n7015), .B(n7019), .Z(n7053) );
  AND U15086 ( .A(n7054), .B(n7055), .Z(n7019) );
  NAND U15087 ( .A(n7056), .B(n7057), .Z(n7055) );
  NAND U15088 ( .A(n7058), .B(n7059), .Z(n7054) );
  AND U15089 ( .A(n7060), .B(n7061), .Z(n7015) );
  NAND U15090 ( .A(n7062), .B(n7063), .Z(n7061) );
  NAND U15091 ( .A(n7064), .B(n7065), .Z(n7060) );
  AND U15092 ( .A(n7066), .B(n7067), .Z(n7017) );
  NAND U15093 ( .A(n7068), .B(n7069), .Z(n7011) );
  XNOR U15094 ( .A(n6994), .B(n7070), .Z(n7008) );
  XNOR U15095 ( .A(n6998), .B(n6996), .Z(n7070) );
  XOR U15096 ( .A(n7004), .B(n7071), .Z(n6996) );
  XNOR U15097 ( .A(n7001), .B(n7005), .Z(n7071) );
  AND U15098 ( .A(n7072), .B(n7073), .Z(n7005) );
  NAND U15099 ( .A(n7074), .B(n7075), .Z(n7073) );
  NAND U15100 ( .A(n7076), .B(n7077), .Z(n7072) );
  AND U15101 ( .A(n7078), .B(n7079), .Z(n7001) );
  NAND U15102 ( .A(n7080), .B(n7081), .Z(n7079) );
  NAND U15103 ( .A(n7082), .B(n7083), .Z(n7078) );
  NANDN U15104 ( .A(n7084), .B(n7085), .Z(n7004) );
  ANDN U15105 ( .B(n7086), .A(n7087), .Z(n6998) );
  XNOR U15106 ( .A(n6989), .B(n7088), .Z(n6994) );
  XNOR U15107 ( .A(n6987), .B(n6991), .Z(n7088) );
  AND U15108 ( .A(n7089), .B(n7090), .Z(n6991) );
  NAND U15109 ( .A(n7091), .B(n7092), .Z(n7090) );
  NAND U15110 ( .A(n7093), .B(n7094), .Z(n7089) );
  AND U15111 ( .A(n7095), .B(n7096), .Z(n6987) );
  NAND U15112 ( .A(n7097), .B(n7098), .Z(n7096) );
  NAND U15113 ( .A(n7099), .B(n7100), .Z(n7095) );
  AND U15114 ( .A(n7101), .B(n7102), .Z(n6989) );
  XOR U15115 ( .A(n7069), .B(n7068), .Z(N64765) );
  XNOR U15116 ( .A(n7086), .B(n7087), .Z(n7068) );
  XNOR U15117 ( .A(n7101), .B(n7102), .Z(n7087) );
  XOR U15118 ( .A(n7098), .B(n7097), .Z(n7102) );
  XOR U15119 ( .A(y[7716]), .B(x[7716]), .Z(n7097) );
  XOR U15120 ( .A(n7100), .B(n7099), .Z(n7098) );
  XOR U15121 ( .A(y[7718]), .B(x[7718]), .Z(n7099) );
  XOR U15122 ( .A(y[7717]), .B(x[7717]), .Z(n7100) );
  XOR U15123 ( .A(n7092), .B(n7091), .Z(n7101) );
  XOR U15124 ( .A(n7094), .B(n7093), .Z(n7091) );
  XOR U15125 ( .A(y[7715]), .B(x[7715]), .Z(n7093) );
  XOR U15126 ( .A(y[7714]), .B(x[7714]), .Z(n7094) );
  XOR U15127 ( .A(y[7713]), .B(x[7713]), .Z(n7092) );
  XNOR U15128 ( .A(n7085), .B(n7084), .Z(n7086) );
  XNOR U15129 ( .A(n7081), .B(n7080), .Z(n7084) );
  XOR U15130 ( .A(n7083), .B(n7082), .Z(n7080) );
  XOR U15131 ( .A(y[7712]), .B(x[7712]), .Z(n7082) );
  XOR U15132 ( .A(y[7711]), .B(x[7711]), .Z(n7083) );
  XOR U15133 ( .A(y[7710]), .B(x[7710]), .Z(n7081) );
  XOR U15134 ( .A(n7075), .B(n7074), .Z(n7085) );
  XOR U15135 ( .A(n7077), .B(n7076), .Z(n7074) );
  XOR U15136 ( .A(y[7709]), .B(x[7709]), .Z(n7076) );
  XOR U15137 ( .A(y[7708]), .B(x[7708]), .Z(n7077) );
  XOR U15138 ( .A(y[7707]), .B(x[7707]), .Z(n7075) );
  XNOR U15139 ( .A(n7051), .B(n7052), .Z(n7069) );
  XNOR U15140 ( .A(n7066), .B(n7067), .Z(n7052) );
  XOR U15141 ( .A(n7063), .B(n7062), .Z(n7067) );
  XOR U15142 ( .A(y[7704]), .B(x[7704]), .Z(n7062) );
  XOR U15143 ( .A(n7065), .B(n7064), .Z(n7063) );
  XOR U15144 ( .A(y[7706]), .B(x[7706]), .Z(n7064) );
  XOR U15145 ( .A(y[7705]), .B(x[7705]), .Z(n7065) );
  XOR U15146 ( .A(n7057), .B(n7056), .Z(n7066) );
  XOR U15147 ( .A(n7059), .B(n7058), .Z(n7056) );
  XOR U15148 ( .A(y[7703]), .B(x[7703]), .Z(n7058) );
  XOR U15149 ( .A(y[7702]), .B(x[7702]), .Z(n7059) );
  XOR U15150 ( .A(y[7701]), .B(x[7701]), .Z(n7057) );
  XNOR U15151 ( .A(n7050), .B(n7049), .Z(n7051) );
  XNOR U15152 ( .A(n7046), .B(n7045), .Z(n7049) );
  XOR U15153 ( .A(n7048), .B(n7047), .Z(n7045) );
  XOR U15154 ( .A(y[7700]), .B(x[7700]), .Z(n7047) );
  XOR U15155 ( .A(y[7699]), .B(x[7699]), .Z(n7048) );
  XOR U15156 ( .A(y[7698]), .B(x[7698]), .Z(n7046) );
  XOR U15157 ( .A(n7040), .B(n7039), .Z(n7050) );
  XOR U15158 ( .A(n7042), .B(n7041), .Z(n7039) );
  XOR U15159 ( .A(y[7697]), .B(x[7697]), .Z(n7041) );
  XOR U15160 ( .A(y[7696]), .B(x[7696]), .Z(n7042) );
  XOR U15161 ( .A(y[7695]), .B(x[7695]), .Z(n7040) );
  NAND U15162 ( .A(n7103), .B(n7104), .Z(N64756) );
  NAND U15163 ( .A(n7105), .B(n7106), .Z(n7104) );
  NANDN U15164 ( .A(n7107), .B(n7108), .Z(n7106) );
  NANDN U15165 ( .A(n7108), .B(n7107), .Z(n7103) );
  XOR U15166 ( .A(n7107), .B(n7109), .Z(N64755) );
  XNOR U15167 ( .A(n7105), .B(n7108), .Z(n7109) );
  NAND U15168 ( .A(n7110), .B(n7111), .Z(n7108) );
  NAND U15169 ( .A(n7112), .B(n7113), .Z(n7111) );
  NANDN U15170 ( .A(n7114), .B(n7115), .Z(n7113) );
  NANDN U15171 ( .A(n7115), .B(n7114), .Z(n7110) );
  AND U15172 ( .A(n7116), .B(n7117), .Z(n7105) );
  NAND U15173 ( .A(n7118), .B(n7119), .Z(n7117) );
  NANDN U15174 ( .A(n7120), .B(n7121), .Z(n7119) );
  NANDN U15175 ( .A(n7121), .B(n7120), .Z(n7116) );
  IV U15176 ( .A(n7122), .Z(n7121) );
  AND U15177 ( .A(n7123), .B(n7124), .Z(n7107) );
  NAND U15178 ( .A(n7125), .B(n7126), .Z(n7124) );
  NANDN U15179 ( .A(n7127), .B(n7128), .Z(n7126) );
  NANDN U15180 ( .A(n7128), .B(n7127), .Z(n7123) );
  XOR U15181 ( .A(n7120), .B(n7129), .Z(N64754) );
  XNOR U15182 ( .A(n7118), .B(n7122), .Z(n7129) );
  XOR U15183 ( .A(n7115), .B(n7130), .Z(n7122) );
  XNOR U15184 ( .A(n7112), .B(n7114), .Z(n7130) );
  AND U15185 ( .A(n7131), .B(n7132), .Z(n7114) );
  NANDN U15186 ( .A(n7133), .B(n7134), .Z(n7132) );
  OR U15187 ( .A(n7135), .B(n7136), .Z(n7134) );
  IV U15188 ( .A(n7137), .Z(n7136) );
  NANDN U15189 ( .A(n7137), .B(n7135), .Z(n7131) );
  AND U15190 ( .A(n7138), .B(n7139), .Z(n7112) );
  NAND U15191 ( .A(n7140), .B(n7141), .Z(n7139) );
  NANDN U15192 ( .A(n7142), .B(n7143), .Z(n7141) );
  NANDN U15193 ( .A(n7143), .B(n7142), .Z(n7138) );
  IV U15194 ( .A(n7144), .Z(n7143) );
  NAND U15195 ( .A(n7145), .B(n7146), .Z(n7115) );
  NANDN U15196 ( .A(n7147), .B(n7148), .Z(n7146) );
  NANDN U15197 ( .A(n7149), .B(n7150), .Z(n7148) );
  NANDN U15198 ( .A(n7150), .B(n7149), .Z(n7145) );
  IV U15199 ( .A(n7151), .Z(n7149) );
  AND U15200 ( .A(n7152), .B(n7153), .Z(n7118) );
  NAND U15201 ( .A(n7154), .B(n7155), .Z(n7153) );
  NANDN U15202 ( .A(n7156), .B(n7157), .Z(n7155) );
  NANDN U15203 ( .A(n7157), .B(n7156), .Z(n7152) );
  XOR U15204 ( .A(n7128), .B(n7158), .Z(n7120) );
  XNOR U15205 ( .A(n7125), .B(n7127), .Z(n7158) );
  AND U15206 ( .A(n7159), .B(n7160), .Z(n7127) );
  NANDN U15207 ( .A(n7161), .B(n7162), .Z(n7160) );
  OR U15208 ( .A(n7163), .B(n7164), .Z(n7162) );
  IV U15209 ( .A(n7165), .Z(n7164) );
  NANDN U15210 ( .A(n7165), .B(n7163), .Z(n7159) );
  AND U15211 ( .A(n7166), .B(n7167), .Z(n7125) );
  NAND U15212 ( .A(n7168), .B(n7169), .Z(n7167) );
  NANDN U15213 ( .A(n7170), .B(n7171), .Z(n7169) );
  NANDN U15214 ( .A(n7171), .B(n7170), .Z(n7166) );
  IV U15215 ( .A(n7172), .Z(n7171) );
  NAND U15216 ( .A(n7173), .B(n7174), .Z(n7128) );
  NANDN U15217 ( .A(n7175), .B(n7176), .Z(n7174) );
  NANDN U15218 ( .A(n7177), .B(n7178), .Z(n7176) );
  NANDN U15219 ( .A(n7178), .B(n7177), .Z(n7173) );
  IV U15220 ( .A(n7179), .Z(n7177) );
  XOR U15221 ( .A(n7154), .B(n7180), .Z(N64753) );
  XNOR U15222 ( .A(n7157), .B(n7156), .Z(n7180) );
  XNOR U15223 ( .A(n7168), .B(n7181), .Z(n7156) );
  XNOR U15224 ( .A(n7172), .B(n7170), .Z(n7181) );
  XOR U15225 ( .A(n7178), .B(n7182), .Z(n7170) );
  XNOR U15226 ( .A(n7175), .B(n7179), .Z(n7182) );
  AND U15227 ( .A(n7183), .B(n7184), .Z(n7179) );
  NAND U15228 ( .A(n7185), .B(n7186), .Z(n7184) );
  NAND U15229 ( .A(n7187), .B(n7188), .Z(n7183) );
  AND U15230 ( .A(n7189), .B(n7190), .Z(n7175) );
  NAND U15231 ( .A(n7191), .B(n7192), .Z(n7190) );
  NAND U15232 ( .A(n7193), .B(n7194), .Z(n7189) );
  NANDN U15233 ( .A(n7195), .B(n7196), .Z(n7178) );
  ANDN U15234 ( .B(n7197), .A(n7198), .Z(n7172) );
  XNOR U15235 ( .A(n7163), .B(n7199), .Z(n7168) );
  XNOR U15236 ( .A(n7161), .B(n7165), .Z(n7199) );
  AND U15237 ( .A(n7200), .B(n7201), .Z(n7165) );
  NAND U15238 ( .A(n7202), .B(n7203), .Z(n7201) );
  NAND U15239 ( .A(n7204), .B(n7205), .Z(n7200) );
  AND U15240 ( .A(n7206), .B(n7207), .Z(n7161) );
  NAND U15241 ( .A(n7208), .B(n7209), .Z(n7207) );
  NAND U15242 ( .A(n7210), .B(n7211), .Z(n7206) );
  AND U15243 ( .A(n7212), .B(n7213), .Z(n7163) );
  NAND U15244 ( .A(n7214), .B(n7215), .Z(n7157) );
  XNOR U15245 ( .A(n7140), .B(n7216), .Z(n7154) );
  XNOR U15246 ( .A(n7144), .B(n7142), .Z(n7216) );
  XOR U15247 ( .A(n7150), .B(n7217), .Z(n7142) );
  XNOR U15248 ( .A(n7147), .B(n7151), .Z(n7217) );
  AND U15249 ( .A(n7218), .B(n7219), .Z(n7151) );
  NAND U15250 ( .A(n7220), .B(n7221), .Z(n7219) );
  NAND U15251 ( .A(n7222), .B(n7223), .Z(n7218) );
  AND U15252 ( .A(n7224), .B(n7225), .Z(n7147) );
  NAND U15253 ( .A(n7226), .B(n7227), .Z(n7225) );
  NAND U15254 ( .A(n7228), .B(n7229), .Z(n7224) );
  NANDN U15255 ( .A(n7230), .B(n7231), .Z(n7150) );
  ANDN U15256 ( .B(n7232), .A(n7233), .Z(n7144) );
  XNOR U15257 ( .A(n7135), .B(n7234), .Z(n7140) );
  XNOR U15258 ( .A(n7133), .B(n7137), .Z(n7234) );
  AND U15259 ( .A(n7235), .B(n7236), .Z(n7137) );
  NAND U15260 ( .A(n7237), .B(n7238), .Z(n7236) );
  NAND U15261 ( .A(n7239), .B(n7240), .Z(n7235) );
  AND U15262 ( .A(n7241), .B(n7242), .Z(n7133) );
  NAND U15263 ( .A(n7243), .B(n7244), .Z(n7242) );
  NAND U15264 ( .A(n7245), .B(n7246), .Z(n7241) );
  AND U15265 ( .A(n7247), .B(n7248), .Z(n7135) );
  XOR U15266 ( .A(n7215), .B(n7214), .Z(N64752) );
  XNOR U15267 ( .A(n7232), .B(n7233), .Z(n7214) );
  XNOR U15268 ( .A(n7247), .B(n7248), .Z(n7233) );
  XOR U15269 ( .A(n7244), .B(n7243), .Z(n7248) );
  XOR U15270 ( .A(y[7692]), .B(x[7692]), .Z(n7243) );
  XOR U15271 ( .A(n7246), .B(n7245), .Z(n7244) );
  XOR U15272 ( .A(y[7694]), .B(x[7694]), .Z(n7245) );
  XOR U15273 ( .A(y[7693]), .B(x[7693]), .Z(n7246) );
  XOR U15274 ( .A(n7238), .B(n7237), .Z(n7247) );
  XOR U15275 ( .A(n7240), .B(n7239), .Z(n7237) );
  XOR U15276 ( .A(y[7691]), .B(x[7691]), .Z(n7239) );
  XOR U15277 ( .A(y[7690]), .B(x[7690]), .Z(n7240) );
  XOR U15278 ( .A(y[7689]), .B(x[7689]), .Z(n7238) );
  XNOR U15279 ( .A(n7231), .B(n7230), .Z(n7232) );
  XNOR U15280 ( .A(n7227), .B(n7226), .Z(n7230) );
  XOR U15281 ( .A(n7229), .B(n7228), .Z(n7226) );
  XOR U15282 ( .A(y[7688]), .B(x[7688]), .Z(n7228) );
  XOR U15283 ( .A(y[7687]), .B(x[7687]), .Z(n7229) );
  XOR U15284 ( .A(y[7686]), .B(x[7686]), .Z(n7227) );
  XOR U15285 ( .A(n7221), .B(n7220), .Z(n7231) );
  XOR U15286 ( .A(n7223), .B(n7222), .Z(n7220) );
  XOR U15287 ( .A(y[7685]), .B(x[7685]), .Z(n7222) );
  XOR U15288 ( .A(y[7684]), .B(x[7684]), .Z(n7223) );
  XOR U15289 ( .A(y[7683]), .B(x[7683]), .Z(n7221) );
  XNOR U15290 ( .A(n7197), .B(n7198), .Z(n7215) );
  XNOR U15291 ( .A(n7212), .B(n7213), .Z(n7198) );
  XOR U15292 ( .A(n7209), .B(n7208), .Z(n7213) );
  XOR U15293 ( .A(y[7680]), .B(x[7680]), .Z(n7208) );
  XOR U15294 ( .A(n7211), .B(n7210), .Z(n7209) );
  XOR U15295 ( .A(y[7682]), .B(x[7682]), .Z(n7210) );
  XOR U15296 ( .A(y[7681]), .B(x[7681]), .Z(n7211) );
  XOR U15297 ( .A(n7203), .B(n7202), .Z(n7212) );
  XOR U15298 ( .A(n7205), .B(n7204), .Z(n7202) );
  XOR U15299 ( .A(y[7679]), .B(x[7679]), .Z(n7204) );
  XOR U15300 ( .A(y[7678]), .B(x[7678]), .Z(n7205) );
  XOR U15301 ( .A(y[7677]), .B(x[7677]), .Z(n7203) );
  XNOR U15302 ( .A(n7196), .B(n7195), .Z(n7197) );
  XNOR U15303 ( .A(n7192), .B(n7191), .Z(n7195) );
  XOR U15304 ( .A(n7194), .B(n7193), .Z(n7191) );
  XOR U15305 ( .A(y[7676]), .B(x[7676]), .Z(n7193) );
  XOR U15306 ( .A(y[7675]), .B(x[7675]), .Z(n7194) );
  XOR U15307 ( .A(y[7674]), .B(x[7674]), .Z(n7192) );
  XOR U15308 ( .A(n7186), .B(n7185), .Z(n7196) );
  XOR U15309 ( .A(n7188), .B(n7187), .Z(n7185) );
  XOR U15310 ( .A(y[7673]), .B(x[7673]), .Z(n7187) );
  XOR U15311 ( .A(y[7672]), .B(x[7672]), .Z(n7188) );
  XOR U15312 ( .A(y[7671]), .B(x[7671]), .Z(n7186) );
  NAND U15313 ( .A(n7249), .B(n7250), .Z(N64743) );
  NAND U15314 ( .A(n7251), .B(n7252), .Z(n7250) );
  NANDN U15315 ( .A(n7253), .B(n7254), .Z(n7252) );
  NANDN U15316 ( .A(n7254), .B(n7253), .Z(n7249) );
  XOR U15317 ( .A(n7253), .B(n7255), .Z(N64742) );
  XNOR U15318 ( .A(n7251), .B(n7254), .Z(n7255) );
  NAND U15319 ( .A(n7256), .B(n7257), .Z(n7254) );
  NAND U15320 ( .A(n7258), .B(n7259), .Z(n7257) );
  NANDN U15321 ( .A(n7260), .B(n7261), .Z(n7259) );
  NANDN U15322 ( .A(n7261), .B(n7260), .Z(n7256) );
  AND U15323 ( .A(n7262), .B(n7263), .Z(n7251) );
  NAND U15324 ( .A(n7264), .B(n7265), .Z(n7263) );
  NANDN U15325 ( .A(n7266), .B(n7267), .Z(n7265) );
  NANDN U15326 ( .A(n7267), .B(n7266), .Z(n7262) );
  IV U15327 ( .A(n7268), .Z(n7267) );
  AND U15328 ( .A(n7269), .B(n7270), .Z(n7253) );
  NAND U15329 ( .A(n7271), .B(n7272), .Z(n7270) );
  NANDN U15330 ( .A(n7273), .B(n7274), .Z(n7272) );
  NANDN U15331 ( .A(n7274), .B(n7273), .Z(n7269) );
  XOR U15332 ( .A(n7266), .B(n7275), .Z(N64741) );
  XNOR U15333 ( .A(n7264), .B(n7268), .Z(n7275) );
  XOR U15334 ( .A(n7261), .B(n7276), .Z(n7268) );
  XNOR U15335 ( .A(n7258), .B(n7260), .Z(n7276) );
  AND U15336 ( .A(n7277), .B(n7278), .Z(n7260) );
  NANDN U15337 ( .A(n7279), .B(n7280), .Z(n7278) );
  OR U15338 ( .A(n7281), .B(n7282), .Z(n7280) );
  IV U15339 ( .A(n7283), .Z(n7282) );
  NANDN U15340 ( .A(n7283), .B(n7281), .Z(n7277) );
  AND U15341 ( .A(n7284), .B(n7285), .Z(n7258) );
  NAND U15342 ( .A(n7286), .B(n7287), .Z(n7285) );
  NANDN U15343 ( .A(n7288), .B(n7289), .Z(n7287) );
  NANDN U15344 ( .A(n7289), .B(n7288), .Z(n7284) );
  IV U15345 ( .A(n7290), .Z(n7289) );
  NAND U15346 ( .A(n7291), .B(n7292), .Z(n7261) );
  NANDN U15347 ( .A(n7293), .B(n7294), .Z(n7292) );
  NANDN U15348 ( .A(n7295), .B(n7296), .Z(n7294) );
  NANDN U15349 ( .A(n7296), .B(n7295), .Z(n7291) );
  IV U15350 ( .A(n7297), .Z(n7295) );
  AND U15351 ( .A(n7298), .B(n7299), .Z(n7264) );
  NAND U15352 ( .A(n7300), .B(n7301), .Z(n7299) );
  NANDN U15353 ( .A(n7302), .B(n7303), .Z(n7301) );
  NANDN U15354 ( .A(n7303), .B(n7302), .Z(n7298) );
  XOR U15355 ( .A(n7274), .B(n7304), .Z(n7266) );
  XNOR U15356 ( .A(n7271), .B(n7273), .Z(n7304) );
  AND U15357 ( .A(n7305), .B(n7306), .Z(n7273) );
  NANDN U15358 ( .A(n7307), .B(n7308), .Z(n7306) );
  OR U15359 ( .A(n7309), .B(n7310), .Z(n7308) );
  IV U15360 ( .A(n7311), .Z(n7310) );
  NANDN U15361 ( .A(n7311), .B(n7309), .Z(n7305) );
  AND U15362 ( .A(n7312), .B(n7313), .Z(n7271) );
  NAND U15363 ( .A(n7314), .B(n7315), .Z(n7313) );
  NANDN U15364 ( .A(n7316), .B(n7317), .Z(n7315) );
  NANDN U15365 ( .A(n7317), .B(n7316), .Z(n7312) );
  IV U15366 ( .A(n7318), .Z(n7317) );
  NAND U15367 ( .A(n7319), .B(n7320), .Z(n7274) );
  NANDN U15368 ( .A(n7321), .B(n7322), .Z(n7320) );
  NANDN U15369 ( .A(n7323), .B(n7324), .Z(n7322) );
  NANDN U15370 ( .A(n7324), .B(n7323), .Z(n7319) );
  IV U15371 ( .A(n7325), .Z(n7323) );
  XOR U15372 ( .A(n7300), .B(n7326), .Z(N64740) );
  XNOR U15373 ( .A(n7303), .B(n7302), .Z(n7326) );
  XNOR U15374 ( .A(n7314), .B(n7327), .Z(n7302) );
  XNOR U15375 ( .A(n7318), .B(n7316), .Z(n7327) );
  XOR U15376 ( .A(n7324), .B(n7328), .Z(n7316) );
  XNOR U15377 ( .A(n7321), .B(n7325), .Z(n7328) );
  AND U15378 ( .A(n7329), .B(n7330), .Z(n7325) );
  NAND U15379 ( .A(n7331), .B(n7332), .Z(n7330) );
  NAND U15380 ( .A(n7333), .B(n7334), .Z(n7329) );
  AND U15381 ( .A(n7335), .B(n7336), .Z(n7321) );
  NAND U15382 ( .A(n7337), .B(n7338), .Z(n7336) );
  NAND U15383 ( .A(n7339), .B(n7340), .Z(n7335) );
  NANDN U15384 ( .A(n7341), .B(n7342), .Z(n7324) );
  ANDN U15385 ( .B(n7343), .A(n7344), .Z(n7318) );
  XNOR U15386 ( .A(n7309), .B(n7345), .Z(n7314) );
  XNOR U15387 ( .A(n7307), .B(n7311), .Z(n7345) );
  AND U15388 ( .A(n7346), .B(n7347), .Z(n7311) );
  NAND U15389 ( .A(n7348), .B(n7349), .Z(n7347) );
  NAND U15390 ( .A(n7350), .B(n7351), .Z(n7346) );
  AND U15391 ( .A(n7352), .B(n7353), .Z(n7307) );
  NAND U15392 ( .A(n7354), .B(n7355), .Z(n7353) );
  NAND U15393 ( .A(n7356), .B(n7357), .Z(n7352) );
  AND U15394 ( .A(n7358), .B(n7359), .Z(n7309) );
  NAND U15395 ( .A(n7360), .B(n7361), .Z(n7303) );
  XNOR U15396 ( .A(n7286), .B(n7362), .Z(n7300) );
  XNOR U15397 ( .A(n7290), .B(n7288), .Z(n7362) );
  XOR U15398 ( .A(n7296), .B(n7363), .Z(n7288) );
  XNOR U15399 ( .A(n7293), .B(n7297), .Z(n7363) );
  AND U15400 ( .A(n7364), .B(n7365), .Z(n7297) );
  NAND U15401 ( .A(n7366), .B(n7367), .Z(n7365) );
  NAND U15402 ( .A(n7368), .B(n7369), .Z(n7364) );
  AND U15403 ( .A(n7370), .B(n7371), .Z(n7293) );
  NAND U15404 ( .A(n7372), .B(n7373), .Z(n7371) );
  NAND U15405 ( .A(n7374), .B(n7375), .Z(n7370) );
  NANDN U15406 ( .A(n7376), .B(n7377), .Z(n7296) );
  ANDN U15407 ( .B(n7378), .A(n7379), .Z(n7290) );
  XNOR U15408 ( .A(n7281), .B(n7380), .Z(n7286) );
  XNOR U15409 ( .A(n7279), .B(n7283), .Z(n7380) );
  AND U15410 ( .A(n7381), .B(n7382), .Z(n7283) );
  NAND U15411 ( .A(n7383), .B(n7384), .Z(n7382) );
  NAND U15412 ( .A(n7385), .B(n7386), .Z(n7381) );
  AND U15413 ( .A(n7387), .B(n7388), .Z(n7279) );
  NAND U15414 ( .A(n7389), .B(n7390), .Z(n7388) );
  NAND U15415 ( .A(n7391), .B(n7392), .Z(n7387) );
  AND U15416 ( .A(n7393), .B(n7394), .Z(n7281) );
  XOR U15417 ( .A(n7361), .B(n7360), .Z(N64739) );
  XNOR U15418 ( .A(n7378), .B(n7379), .Z(n7360) );
  XNOR U15419 ( .A(n7393), .B(n7394), .Z(n7379) );
  XOR U15420 ( .A(n7390), .B(n7389), .Z(n7394) );
  XOR U15421 ( .A(y[7668]), .B(x[7668]), .Z(n7389) );
  XOR U15422 ( .A(n7392), .B(n7391), .Z(n7390) );
  XOR U15423 ( .A(y[7670]), .B(x[7670]), .Z(n7391) );
  XOR U15424 ( .A(y[7669]), .B(x[7669]), .Z(n7392) );
  XOR U15425 ( .A(n7384), .B(n7383), .Z(n7393) );
  XOR U15426 ( .A(n7386), .B(n7385), .Z(n7383) );
  XOR U15427 ( .A(y[7667]), .B(x[7667]), .Z(n7385) );
  XOR U15428 ( .A(y[7666]), .B(x[7666]), .Z(n7386) );
  XOR U15429 ( .A(y[7665]), .B(x[7665]), .Z(n7384) );
  XNOR U15430 ( .A(n7377), .B(n7376), .Z(n7378) );
  XNOR U15431 ( .A(n7373), .B(n7372), .Z(n7376) );
  XOR U15432 ( .A(n7375), .B(n7374), .Z(n7372) );
  XOR U15433 ( .A(y[7664]), .B(x[7664]), .Z(n7374) );
  XOR U15434 ( .A(y[7663]), .B(x[7663]), .Z(n7375) );
  XOR U15435 ( .A(y[7662]), .B(x[7662]), .Z(n7373) );
  XOR U15436 ( .A(n7367), .B(n7366), .Z(n7377) );
  XOR U15437 ( .A(n7369), .B(n7368), .Z(n7366) );
  XOR U15438 ( .A(y[7661]), .B(x[7661]), .Z(n7368) );
  XOR U15439 ( .A(y[7660]), .B(x[7660]), .Z(n7369) );
  XOR U15440 ( .A(y[7659]), .B(x[7659]), .Z(n7367) );
  XNOR U15441 ( .A(n7343), .B(n7344), .Z(n7361) );
  XNOR U15442 ( .A(n7358), .B(n7359), .Z(n7344) );
  XOR U15443 ( .A(n7355), .B(n7354), .Z(n7359) );
  XOR U15444 ( .A(y[7656]), .B(x[7656]), .Z(n7354) );
  XOR U15445 ( .A(n7357), .B(n7356), .Z(n7355) );
  XOR U15446 ( .A(y[7658]), .B(x[7658]), .Z(n7356) );
  XOR U15447 ( .A(y[7657]), .B(x[7657]), .Z(n7357) );
  XOR U15448 ( .A(n7349), .B(n7348), .Z(n7358) );
  XOR U15449 ( .A(n7351), .B(n7350), .Z(n7348) );
  XOR U15450 ( .A(y[7655]), .B(x[7655]), .Z(n7350) );
  XOR U15451 ( .A(y[7654]), .B(x[7654]), .Z(n7351) );
  XOR U15452 ( .A(y[7653]), .B(x[7653]), .Z(n7349) );
  XNOR U15453 ( .A(n7342), .B(n7341), .Z(n7343) );
  XNOR U15454 ( .A(n7338), .B(n7337), .Z(n7341) );
  XOR U15455 ( .A(n7340), .B(n7339), .Z(n7337) );
  XOR U15456 ( .A(y[7652]), .B(x[7652]), .Z(n7339) );
  XOR U15457 ( .A(y[7651]), .B(x[7651]), .Z(n7340) );
  XOR U15458 ( .A(y[7650]), .B(x[7650]), .Z(n7338) );
  XOR U15459 ( .A(n7332), .B(n7331), .Z(n7342) );
  XOR U15460 ( .A(n7334), .B(n7333), .Z(n7331) );
  XOR U15461 ( .A(y[7649]), .B(x[7649]), .Z(n7333) );
  XOR U15462 ( .A(y[7648]), .B(x[7648]), .Z(n7334) );
  XOR U15463 ( .A(y[7647]), .B(x[7647]), .Z(n7332) );
  NAND U15464 ( .A(n7395), .B(n7396), .Z(N64730) );
  NAND U15465 ( .A(n7397), .B(n7398), .Z(n7396) );
  NANDN U15466 ( .A(n7399), .B(n7400), .Z(n7398) );
  NANDN U15467 ( .A(n7400), .B(n7399), .Z(n7395) );
  XOR U15468 ( .A(n7399), .B(n7401), .Z(N64729) );
  XNOR U15469 ( .A(n7397), .B(n7400), .Z(n7401) );
  NAND U15470 ( .A(n7402), .B(n7403), .Z(n7400) );
  NAND U15471 ( .A(n7404), .B(n7405), .Z(n7403) );
  NANDN U15472 ( .A(n7406), .B(n7407), .Z(n7405) );
  NANDN U15473 ( .A(n7407), .B(n7406), .Z(n7402) );
  AND U15474 ( .A(n7408), .B(n7409), .Z(n7397) );
  NAND U15475 ( .A(n7410), .B(n7411), .Z(n7409) );
  NANDN U15476 ( .A(n7412), .B(n7413), .Z(n7411) );
  NANDN U15477 ( .A(n7413), .B(n7412), .Z(n7408) );
  IV U15478 ( .A(n7414), .Z(n7413) );
  AND U15479 ( .A(n7415), .B(n7416), .Z(n7399) );
  NAND U15480 ( .A(n7417), .B(n7418), .Z(n7416) );
  NANDN U15481 ( .A(n7419), .B(n7420), .Z(n7418) );
  NANDN U15482 ( .A(n7420), .B(n7419), .Z(n7415) );
  XOR U15483 ( .A(n7412), .B(n7421), .Z(N64728) );
  XNOR U15484 ( .A(n7410), .B(n7414), .Z(n7421) );
  XOR U15485 ( .A(n7407), .B(n7422), .Z(n7414) );
  XNOR U15486 ( .A(n7404), .B(n7406), .Z(n7422) );
  AND U15487 ( .A(n7423), .B(n7424), .Z(n7406) );
  NANDN U15488 ( .A(n7425), .B(n7426), .Z(n7424) );
  OR U15489 ( .A(n7427), .B(n7428), .Z(n7426) );
  IV U15490 ( .A(n7429), .Z(n7428) );
  NANDN U15491 ( .A(n7429), .B(n7427), .Z(n7423) );
  AND U15492 ( .A(n7430), .B(n7431), .Z(n7404) );
  NAND U15493 ( .A(n7432), .B(n7433), .Z(n7431) );
  NANDN U15494 ( .A(n7434), .B(n7435), .Z(n7433) );
  NANDN U15495 ( .A(n7435), .B(n7434), .Z(n7430) );
  IV U15496 ( .A(n7436), .Z(n7435) );
  NAND U15497 ( .A(n7437), .B(n7438), .Z(n7407) );
  NANDN U15498 ( .A(n7439), .B(n7440), .Z(n7438) );
  NANDN U15499 ( .A(n7441), .B(n7442), .Z(n7440) );
  NANDN U15500 ( .A(n7442), .B(n7441), .Z(n7437) );
  IV U15501 ( .A(n7443), .Z(n7441) );
  AND U15502 ( .A(n7444), .B(n7445), .Z(n7410) );
  NAND U15503 ( .A(n7446), .B(n7447), .Z(n7445) );
  NANDN U15504 ( .A(n7448), .B(n7449), .Z(n7447) );
  NANDN U15505 ( .A(n7449), .B(n7448), .Z(n7444) );
  XOR U15506 ( .A(n7420), .B(n7450), .Z(n7412) );
  XNOR U15507 ( .A(n7417), .B(n7419), .Z(n7450) );
  AND U15508 ( .A(n7451), .B(n7452), .Z(n7419) );
  NANDN U15509 ( .A(n7453), .B(n7454), .Z(n7452) );
  OR U15510 ( .A(n7455), .B(n7456), .Z(n7454) );
  IV U15511 ( .A(n7457), .Z(n7456) );
  NANDN U15512 ( .A(n7457), .B(n7455), .Z(n7451) );
  AND U15513 ( .A(n7458), .B(n7459), .Z(n7417) );
  NAND U15514 ( .A(n7460), .B(n7461), .Z(n7459) );
  NANDN U15515 ( .A(n7462), .B(n7463), .Z(n7461) );
  NANDN U15516 ( .A(n7463), .B(n7462), .Z(n7458) );
  IV U15517 ( .A(n7464), .Z(n7463) );
  NAND U15518 ( .A(n7465), .B(n7466), .Z(n7420) );
  NANDN U15519 ( .A(n7467), .B(n7468), .Z(n7466) );
  NANDN U15520 ( .A(n7469), .B(n7470), .Z(n7468) );
  NANDN U15521 ( .A(n7470), .B(n7469), .Z(n7465) );
  IV U15522 ( .A(n7471), .Z(n7469) );
  XOR U15523 ( .A(n7446), .B(n7472), .Z(N64727) );
  XNOR U15524 ( .A(n7449), .B(n7448), .Z(n7472) );
  XNOR U15525 ( .A(n7460), .B(n7473), .Z(n7448) );
  XNOR U15526 ( .A(n7464), .B(n7462), .Z(n7473) );
  XOR U15527 ( .A(n7470), .B(n7474), .Z(n7462) );
  XNOR U15528 ( .A(n7467), .B(n7471), .Z(n7474) );
  AND U15529 ( .A(n7475), .B(n7476), .Z(n7471) );
  NAND U15530 ( .A(n7477), .B(n7478), .Z(n7476) );
  NAND U15531 ( .A(n7479), .B(n7480), .Z(n7475) );
  AND U15532 ( .A(n7481), .B(n7482), .Z(n7467) );
  NAND U15533 ( .A(n7483), .B(n7484), .Z(n7482) );
  NAND U15534 ( .A(n7485), .B(n7486), .Z(n7481) );
  NANDN U15535 ( .A(n7487), .B(n7488), .Z(n7470) );
  ANDN U15536 ( .B(n7489), .A(n7490), .Z(n7464) );
  XNOR U15537 ( .A(n7455), .B(n7491), .Z(n7460) );
  XNOR U15538 ( .A(n7453), .B(n7457), .Z(n7491) );
  AND U15539 ( .A(n7492), .B(n7493), .Z(n7457) );
  NAND U15540 ( .A(n7494), .B(n7495), .Z(n7493) );
  NAND U15541 ( .A(n7496), .B(n7497), .Z(n7492) );
  AND U15542 ( .A(n7498), .B(n7499), .Z(n7453) );
  NAND U15543 ( .A(n7500), .B(n7501), .Z(n7499) );
  NAND U15544 ( .A(n7502), .B(n7503), .Z(n7498) );
  AND U15545 ( .A(n7504), .B(n7505), .Z(n7455) );
  NAND U15546 ( .A(n7506), .B(n7507), .Z(n7449) );
  XNOR U15547 ( .A(n7432), .B(n7508), .Z(n7446) );
  XNOR U15548 ( .A(n7436), .B(n7434), .Z(n7508) );
  XOR U15549 ( .A(n7442), .B(n7509), .Z(n7434) );
  XNOR U15550 ( .A(n7439), .B(n7443), .Z(n7509) );
  AND U15551 ( .A(n7510), .B(n7511), .Z(n7443) );
  NAND U15552 ( .A(n7512), .B(n7513), .Z(n7511) );
  NAND U15553 ( .A(n7514), .B(n7515), .Z(n7510) );
  AND U15554 ( .A(n7516), .B(n7517), .Z(n7439) );
  NAND U15555 ( .A(n7518), .B(n7519), .Z(n7517) );
  NAND U15556 ( .A(n7520), .B(n7521), .Z(n7516) );
  NANDN U15557 ( .A(n7522), .B(n7523), .Z(n7442) );
  ANDN U15558 ( .B(n7524), .A(n7525), .Z(n7436) );
  XNOR U15559 ( .A(n7427), .B(n7526), .Z(n7432) );
  XNOR U15560 ( .A(n7425), .B(n7429), .Z(n7526) );
  AND U15561 ( .A(n7527), .B(n7528), .Z(n7429) );
  NAND U15562 ( .A(n7529), .B(n7530), .Z(n7528) );
  NAND U15563 ( .A(n7531), .B(n7532), .Z(n7527) );
  AND U15564 ( .A(n7533), .B(n7534), .Z(n7425) );
  NAND U15565 ( .A(n7535), .B(n7536), .Z(n7534) );
  NAND U15566 ( .A(n7537), .B(n7538), .Z(n7533) );
  AND U15567 ( .A(n7539), .B(n7540), .Z(n7427) );
  XOR U15568 ( .A(n7507), .B(n7506), .Z(N64726) );
  XNOR U15569 ( .A(n7524), .B(n7525), .Z(n7506) );
  XNOR U15570 ( .A(n7539), .B(n7540), .Z(n7525) );
  XOR U15571 ( .A(n7536), .B(n7535), .Z(n7540) );
  XOR U15572 ( .A(y[7644]), .B(x[7644]), .Z(n7535) );
  XOR U15573 ( .A(n7538), .B(n7537), .Z(n7536) );
  XOR U15574 ( .A(y[7646]), .B(x[7646]), .Z(n7537) );
  XOR U15575 ( .A(y[7645]), .B(x[7645]), .Z(n7538) );
  XOR U15576 ( .A(n7530), .B(n7529), .Z(n7539) );
  XOR U15577 ( .A(n7532), .B(n7531), .Z(n7529) );
  XOR U15578 ( .A(y[7643]), .B(x[7643]), .Z(n7531) );
  XOR U15579 ( .A(y[7642]), .B(x[7642]), .Z(n7532) );
  XOR U15580 ( .A(y[7641]), .B(x[7641]), .Z(n7530) );
  XNOR U15581 ( .A(n7523), .B(n7522), .Z(n7524) );
  XNOR U15582 ( .A(n7519), .B(n7518), .Z(n7522) );
  XOR U15583 ( .A(n7521), .B(n7520), .Z(n7518) );
  XOR U15584 ( .A(y[7640]), .B(x[7640]), .Z(n7520) );
  XOR U15585 ( .A(y[7639]), .B(x[7639]), .Z(n7521) );
  XOR U15586 ( .A(y[7638]), .B(x[7638]), .Z(n7519) );
  XOR U15587 ( .A(n7513), .B(n7512), .Z(n7523) );
  XOR U15588 ( .A(n7515), .B(n7514), .Z(n7512) );
  XOR U15589 ( .A(y[7637]), .B(x[7637]), .Z(n7514) );
  XOR U15590 ( .A(y[7636]), .B(x[7636]), .Z(n7515) );
  XOR U15591 ( .A(y[7635]), .B(x[7635]), .Z(n7513) );
  XNOR U15592 ( .A(n7489), .B(n7490), .Z(n7507) );
  XNOR U15593 ( .A(n7504), .B(n7505), .Z(n7490) );
  XOR U15594 ( .A(n7501), .B(n7500), .Z(n7505) );
  XOR U15595 ( .A(y[7632]), .B(x[7632]), .Z(n7500) );
  XOR U15596 ( .A(n7503), .B(n7502), .Z(n7501) );
  XOR U15597 ( .A(y[7634]), .B(x[7634]), .Z(n7502) );
  XOR U15598 ( .A(y[7633]), .B(x[7633]), .Z(n7503) );
  XOR U15599 ( .A(n7495), .B(n7494), .Z(n7504) );
  XOR U15600 ( .A(n7497), .B(n7496), .Z(n7494) );
  XOR U15601 ( .A(y[7631]), .B(x[7631]), .Z(n7496) );
  XOR U15602 ( .A(y[7630]), .B(x[7630]), .Z(n7497) );
  XOR U15603 ( .A(y[7629]), .B(x[7629]), .Z(n7495) );
  XNOR U15604 ( .A(n7488), .B(n7487), .Z(n7489) );
  XNOR U15605 ( .A(n7484), .B(n7483), .Z(n7487) );
  XOR U15606 ( .A(n7486), .B(n7485), .Z(n7483) );
  XOR U15607 ( .A(y[7628]), .B(x[7628]), .Z(n7485) );
  XOR U15608 ( .A(y[7627]), .B(x[7627]), .Z(n7486) );
  XOR U15609 ( .A(y[7626]), .B(x[7626]), .Z(n7484) );
  XOR U15610 ( .A(n7478), .B(n7477), .Z(n7488) );
  XOR U15611 ( .A(n7480), .B(n7479), .Z(n7477) );
  XOR U15612 ( .A(y[7625]), .B(x[7625]), .Z(n7479) );
  XOR U15613 ( .A(y[7624]), .B(x[7624]), .Z(n7480) );
  XOR U15614 ( .A(y[7623]), .B(x[7623]), .Z(n7478) );
  NAND U15615 ( .A(n7541), .B(n7542), .Z(N64717) );
  NAND U15616 ( .A(n7543), .B(n7544), .Z(n7542) );
  NANDN U15617 ( .A(n7545), .B(n7546), .Z(n7544) );
  NANDN U15618 ( .A(n7546), .B(n7545), .Z(n7541) );
  XOR U15619 ( .A(n7545), .B(n7547), .Z(N64716) );
  XNOR U15620 ( .A(n7543), .B(n7546), .Z(n7547) );
  NAND U15621 ( .A(n7548), .B(n7549), .Z(n7546) );
  NAND U15622 ( .A(n7550), .B(n7551), .Z(n7549) );
  NANDN U15623 ( .A(n7552), .B(n7553), .Z(n7551) );
  NANDN U15624 ( .A(n7553), .B(n7552), .Z(n7548) );
  AND U15625 ( .A(n7554), .B(n7555), .Z(n7543) );
  NAND U15626 ( .A(n7556), .B(n7557), .Z(n7555) );
  NANDN U15627 ( .A(n7558), .B(n7559), .Z(n7557) );
  NANDN U15628 ( .A(n7559), .B(n7558), .Z(n7554) );
  IV U15629 ( .A(n7560), .Z(n7559) );
  AND U15630 ( .A(n7561), .B(n7562), .Z(n7545) );
  NAND U15631 ( .A(n7563), .B(n7564), .Z(n7562) );
  NANDN U15632 ( .A(n7565), .B(n7566), .Z(n7564) );
  NANDN U15633 ( .A(n7566), .B(n7565), .Z(n7561) );
  XOR U15634 ( .A(n7558), .B(n7567), .Z(N64715) );
  XNOR U15635 ( .A(n7556), .B(n7560), .Z(n7567) );
  XOR U15636 ( .A(n7553), .B(n7568), .Z(n7560) );
  XNOR U15637 ( .A(n7550), .B(n7552), .Z(n7568) );
  AND U15638 ( .A(n7569), .B(n7570), .Z(n7552) );
  NANDN U15639 ( .A(n7571), .B(n7572), .Z(n7570) );
  OR U15640 ( .A(n7573), .B(n7574), .Z(n7572) );
  IV U15641 ( .A(n7575), .Z(n7574) );
  NANDN U15642 ( .A(n7575), .B(n7573), .Z(n7569) );
  AND U15643 ( .A(n7576), .B(n7577), .Z(n7550) );
  NAND U15644 ( .A(n7578), .B(n7579), .Z(n7577) );
  NANDN U15645 ( .A(n7580), .B(n7581), .Z(n7579) );
  NANDN U15646 ( .A(n7581), .B(n7580), .Z(n7576) );
  IV U15647 ( .A(n7582), .Z(n7581) );
  NAND U15648 ( .A(n7583), .B(n7584), .Z(n7553) );
  NANDN U15649 ( .A(n7585), .B(n7586), .Z(n7584) );
  NANDN U15650 ( .A(n7587), .B(n7588), .Z(n7586) );
  NANDN U15651 ( .A(n7588), .B(n7587), .Z(n7583) );
  IV U15652 ( .A(n7589), .Z(n7587) );
  AND U15653 ( .A(n7590), .B(n7591), .Z(n7556) );
  NAND U15654 ( .A(n7592), .B(n7593), .Z(n7591) );
  NANDN U15655 ( .A(n7594), .B(n7595), .Z(n7593) );
  NANDN U15656 ( .A(n7595), .B(n7594), .Z(n7590) );
  XOR U15657 ( .A(n7566), .B(n7596), .Z(n7558) );
  XNOR U15658 ( .A(n7563), .B(n7565), .Z(n7596) );
  AND U15659 ( .A(n7597), .B(n7598), .Z(n7565) );
  NANDN U15660 ( .A(n7599), .B(n7600), .Z(n7598) );
  OR U15661 ( .A(n7601), .B(n7602), .Z(n7600) );
  IV U15662 ( .A(n7603), .Z(n7602) );
  NANDN U15663 ( .A(n7603), .B(n7601), .Z(n7597) );
  AND U15664 ( .A(n7604), .B(n7605), .Z(n7563) );
  NAND U15665 ( .A(n7606), .B(n7607), .Z(n7605) );
  NANDN U15666 ( .A(n7608), .B(n7609), .Z(n7607) );
  NANDN U15667 ( .A(n7609), .B(n7608), .Z(n7604) );
  IV U15668 ( .A(n7610), .Z(n7609) );
  NAND U15669 ( .A(n7611), .B(n7612), .Z(n7566) );
  NANDN U15670 ( .A(n7613), .B(n7614), .Z(n7612) );
  NANDN U15671 ( .A(n7615), .B(n7616), .Z(n7614) );
  NANDN U15672 ( .A(n7616), .B(n7615), .Z(n7611) );
  IV U15673 ( .A(n7617), .Z(n7615) );
  XOR U15674 ( .A(n7592), .B(n7618), .Z(N64714) );
  XNOR U15675 ( .A(n7595), .B(n7594), .Z(n7618) );
  XNOR U15676 ( .A(n7606), .B(n7619), .Z(n7594) );
  XNOR U15677 ( .A(n7610), .B(n7608), .Z(n7619) );
  XOR U15678 ( .A(n7616), .B(n7620), .Z(n7608) );
  XNOR U15679 ( .A(n7613), .B(n7617), .Z(n7620) );
  AND U15680 ( .A(n7621), .B(n7622), .Z(n7617) );
  NAND U15681 ( .A(n7623), .B(n7624), .Z(n7622) );
  NAND U15682 ( .A(n7625), .B(n7626), .Z(n7621) );
  AND U15683 ( .A(n7627), .B(n7628), .Z(n7613) );
  NAND U15684 ( .A(n7629), .B(n7630), .Z(n7628) );
  NAND U15685 ( .A(n7631), .B(n7632), .Z(n7627) );
  NANDN U15686 ( .A(n7633), .B(n7634), .Z(n7616) );
  ANDN U15687 ( .B(n7635), .A(n7636), .Z(n7610) );
  XNOR U15688 ( .A(n7601), .B(n7637), .Z(n7606) );
  XNOR U15689 ( .A(n7599), .B(n7603), .Z(n7637) );
  AND U15690 ( .A(n7638), .B(n7639), .Z(n7603) );
  NAND U15691 ( .A(n7640), .B(n7641), .Z(n7639) );
  NAND U15692 ( .A(n7642), .B(n7643), .Z(n7638) );
  AND U15693 ( .A(n7644), .B(n7645), .Z(n7599) );
  NAND U15694 ( .A(n7646), .B(n7647), .Z(n7645) );
  NAND U15695 ( .A(n7648), .B(n7649), .Z(n7644) );
  AND U15696 ( .A(n7650), .B(n7651), .Z(n7601) );
  NAND U15697 ( .A(n7652), .B(n7653), .Z(n7595) );
  XNOR U15698 ( .A(n7578), .B(n7654), .Z(n7592) );
  XNOR U15699 ( .A(n7582), .B(n7580), .Z(n7654) );
  XOR U15700 ( .A(n7588), .B(n7655), .Z(n7580) );
  XNOR U15701 ( .A(n7585), .B(n7589), .Z(n7655) );
  AND U15702 ( .A(n7656), .B(n7657), .Z(n7589) );
  NAND U15703 ( .A(n7658), .B(n7659), .Z(n7657) );
  NAND U15704 ( .A(n7660), .B(n7661), .Z(n7656) );
  AND U15705 ( .A(n7662), .B(n7663), .Z(n7585) );
  NAND U15706 ( .A(n7664), .B(n7665), .Z(n7663) );
  NAND U15707 ( .A(n7666), .B(n7667), .Z(n7662) );
  NANDN U15708 ( .A(n7668), .B(n7669), .Z(n7588) );
  ANDN U15709 ( .B(n7670), .A(n7671), .Z(n7582) );
  XNOR U15710 ( .A(n7573), .B(n7672), .Z(n7578) );
  XNOR U15711 ( .A(n7571), .B(n7575), .Z(n7672) );
  AND U15712 ( .A(n7673), .B(n7674), .Z(n7575) );
  NAND U15713 ( .A(n7675), .B(n7676), .Z(n7674) );
  NAND U15714 ( .A(n7677), .B(n7678), .Z(n7673) );
  AND U15715 ( .A(n7679), .B(n7680), .Z(n7571) );
  NAND U15716 ( .A(n7681), .B(n7682), .Z(n7680) );
  NAND U15717 ( .A(n7683), .B(n7684), .Z(n7679) );
  AND U15718 ( .A(n7685), .B(n7686), .Z(n7573) );
  XOR U15719 ( .A(n7653), .B(n7652), .Z(N64713) );
  XNOR U15720 ( .A(n7670), .B(n7671), .Z(n7652) );
  XNOR U15721 ( .A(n7685), .B(n7686), .Z(n7671) );
  XOR U15722 ( .A(n7682), .B(n7681), .Z(n7686) );
  XOR U15723 ( .A(y[7620]), .B(x[7620]), .Z(n7681) );
  XOR U15724 ( .A(n7684), .B(n7683), .Z(n7682) );
  XOR U15725 ( .A(y[7622]), .B(x[7622]), .Z(n7683) );
  XOR U15726 ( .A(y[7621]), .B(x[7621]), .Z(n7684) );
  XOR U15727 ( .A(n7676), .B(n7675), .Z(n7685) );
  XOR U15728 ( .A(n7678), .B(n7677), .Z(n7675) );
  XOR U15729 ( .A(y[7619]), .B(x[7619]), .Z(n7677) );
  XOR U15730 ( .A(y[7618]), .B(x[7618]), .Z(n7678) );
  XOR U15731 ( .A(y[7617]), .B(x[7617]), .Z(n7676) );
  XNOR U15732 ( .A(n7669), .B(n7668), .Z(n7670) );
  XNOR U15733 ( .A(n7665), .B(n7664), .Z(n7668) );
  XOR U15734 ( .A(n7667), .B(n7666), .Z(n7664) );
  XOR U15735 ( .A(y[7616]), .B(x[7616]), .Z(n7666) );
  XOR U15736 ( .A(y[7615]), .B(x[7615]), .Z(n7667) );
  XOR U15737 ( .A(y[7614]), .B(x[7614]), .Z(n7665) );
  XOR U15738 ( .A(n7659), .B(n7658), .Z(n7669) );
  XOR U15739 ( .A(n7661), .B(n7660), .Z(n7658) );
  XOR U15740 ( .A(y[7613]), .B(x[7613]), .Z(n7660) );
  XOR U15741 ( .A(y[7612]), .B(x[7612]), .Z(n7661) );
  XOR U15742 ( .A(y[7611]), .B(x[7611]), .Z(n7659) );
  XNOR U15743 ( .A(n7635), .B(n7636), .Z(n7653) );
  XNOR U15744 ( .A(n7650), .B(n7651), .Z(n7636) );
  XOR U15745 ( .A(n7647), .B(n7646), .Z(n7651) );
  XOR U15746 ( .A(y[7608]), .B(x[7608]), .Z(n7646) );
  XOR U15747 ( .A(n7649), .B(n7648), .Z(n7647) );
  XOR U15748 ( .A(y[7610]), .B(x[7610]), .Z(n7648) );
  XOR U15749 ( .A(y[7609]), .B(x[7609]), .Z(n7649) );
  XOR U15750 ( .A(n7641), .B(n7640), .Z(n7650) );
  XOR U15751 ( .A(n7643), .B(n7642), .Z(n7640) );
  XOR U15752 ( .A(y[7607]), .B(x[7607]), .Z(n7642) );
  XOR U15753 ( .A(y[7606]), .B(x[7606]), .Z(n7643) );
  XOR U15754 ( .A(y[7605]), .B(x[7605]), .Z(n7641) );
  XNOR U15755 ( .A(n7634), .B(n7633), .Z(n7635) );
  XNOR U15756 ( .A(n7630), .B(n7629), .Z(n7633) );
  XOR U15757 ( .A(n7632), .B(n7631), .Z(n7629) );
  XOR U15758 ( .A(y[7604]), .B(x[7604]), .Z(n7631) );
  XOR U15759 ( .A(y[7603]), .B(x[7603]), .Z(n7632) );
  XOR U15760 ( .A(y[7602]), .B(x[7602]), .Z(n7630) );
  XOR U15761 ( .A(n7624), .B(n7623), .Z(n7634) );
  XOR U15762 ( .A(n7626), .B(n7625), .Z(n7623) );
  XOR U15763 ( .A(y[7601]), .B(x[7601]), .Z(n7625) );
  XOR U15764 ( .A(y[7600]), .B(x[7600]), .Z(n7626) );
  XOR U15765 ( .A(y[7599]), .B(x[7599]), .Z(n7624) );
  NAND U15766 ( .A(n7687), .B(n7688), .Z(N64704) );
  NAND U15767 ( .A(n7689), .B(n7690), .Z(n7688) );
  NANDN U15768 ( .A(n7691), .B(n7692), .Z(n7690) );
  NANDN U15769 ( .A(n7692), .B(n7691), .Z(n7687) );
  XOR U15770 ( .A(n7691), .B(n7693), .Z(N64703) );
  XNOR U15771 ( .A(n7689), .B(n7692), .Z(n7693) );
  NAND U15772 ( .A(n7694), .B(n7695), .Z(n7692) );
  NAND U15773 ( .A(n7696), .B(n7697), .Z(n7695) );
  NANDN U15774 ( .A(n7698), .B(n7699), .Z(n7697) );
  NANDN U15775 ( .A(n7699), .B(n7698), .Z(n7694) );
  AND U15776 ( .A(n7700), .B(n7701), .Z(n7689) );
  NAND U15777 ( .A(n7702), .B(n7703), .Z(n7701) );
  NANDN U15778 ( .A(n7704), .B(n7705), .Z(n7703) );
  NANDN U15779 ( .A(n7705), .B(n7704), .Z(n7700) );
  IV U15780 ( .A(n7706), .Z(n7705) );
  AND U15781 ( .A(n7707), .B(n7708), .Z(n7691) );
  NAND U15782 ( .A(n7709), .B(n7710), .Z(n7708) );
  NANDN U15783 ( .A(n7711), .B(n7712), .Z(n7710) );
  NANDN U15784 ( .A(n7712), .B(n7711), .Z(n7707) );
  XOR U15785 ( .A(n7704), .B(n7713), .Z(N64702) );
  XNOR U15786 ( .A(n7702), .B(n7706), .Z(n7713) );
  XOR U15787 ( .A(n7699), .B(n7714), .Z(n7706) );
  XNOR U15788 ( .A(n7696), .B(n7698), .Z(n7714) );
  AND U15789 ( .A(n7715), .B(n7716), .Z(n7698) );
  NANDN U15790 ( .A(n7717), .B(n7718), .Z(n7716) );
  OR U15791 ( .A(n7719), .B(n7720), .Z(n7718) );
  IV U15792 ( .A(n7721), .Z(n7720) );
  NANDN U15793 ( .A(n7721), .B(n7719), .Z(n7715) );
  AND U15794 ( .A(n7722), .B(n7723), .Z(n7696) );
  NAND U15795 ( .A(n7724), .B(n7725), .Z(n7723) );
  NANDN U15796 ( .A(n7726), .B(n7727), .Z(n7725) );
  NANDN U15797 ( .A(n7727), .B(n7726), .Z(n7722) );
  IV U15798 ( .A(n7728), .Z(n7727) );
  NAND U15799 ( .A(n7729), .B(n7730), .Z(n7699) );
  NANDN U15800 ( .A(n7731), .B(n7732), .Z(n7730) );
  NANDN U15801 ( .A(n7733), .B(n7734), .Z(n7732) );
  NANDN U15802 ( .A(n7734), .B(n7733), .Z(n7729) );
  IV U15803 ( .A(n7735), .Z(n7733) );
  AND U15804 ( .A(n7736), .B(n7737), .Z(n7702) );
  NAND U15805 ( .A(n7738), .B(n7739), .Z(n7737) );
  NANDN U15806 ( .A(n7740), .B(n7741), .Z(n7739) );
  NANDN U15807 ( .A(n7741), .B(n7740), .Z(n7736) );
  XOR U15808 ( .A(n7712), .B(n7742), .Z(n7704) );
  XNOR U15809 ( .A(n7709), .B(n7711), .Z(n7742) );
  AND U15810 ( .A(n7743), .B(n7744), .Z(n7711) );
  NANDN U15811 ( .A(n7745), .B(n7746), .Z(n7744) );
  OR U15812 ( .A(n7747), .B(n7748), .Z(n7746) );
  IV U15813 ( .A(n7749), .Z(n7748) );
  NANDN U15814 ( .A(n7749), .B(n7747), .Z(n7743) );
  AND U15815 ( .A(n7750), .B(n7751), .Z(n7709) );
  NAND U15816 ( .A(n7752), .B(n7753), .Z(n7751) );
  NANDN U15817 ( .A(n7754), .B(n7755), .Z(n7753) );
  NANDN U15818 ( .A(n7755), .B(n7754), .Z(n7750) );
  IV U15819 ( .A(n7756), .Z(n7755) );
  NAND U15820 ( .A(n7757), .B(n7758), .Z(n7712) );
  NANDN U15821 ( .A(n7759), .B(n7760), .Z(n7758) );
  NANDN U15822 ( .A(n7761), .B(n7762), .Z(n7760) );
  NANDN U15823 ( .A(n7762), .B(n7761), .Z(n7757) );
  IV U15824 ( .A(n7763), .Z(n7761) );
  XOR U15825 ( .A(n7738), .B(n7764), .Z(N64701) );
  XNOR U15826 ( .A(n7741), .B(n7740), .Z(n7764) );
  XNOR U15827 ( .A(n7752), .B(n7765), .Z(n7740) );
  XNOR U15828 ( .A(n7756), .B(n7754), .Z(n7765) );
  XOR U15829 ( .A(n7762), .B(n7766), .Z(n7754) );
  XNOR U15830 ( .A(n7759), .B(n7763), .Z(n7766) );
  AND U15831 ( .A(n7767), .B(n7768), .Z(n7763) );
  NAND U15832 ( .A(n7769), .B(n7770), .Z(n7768) );
  NAND U15833 ( .A(n7771), .B(n7772), .Z(n7767) );
  AND U15834 ( .A(n7773), .B(n7774), .Z(n7759) );
  NAND U15835 ( .A(n7775), .B(n7776), .Z(n7774) );
  NAND U15836 ( .A(n7777), .B(n7778), .Z(n7773) );
  NANDN U15837 ( .A(n7779), .B(n7780), .Z(n7762) );
  ANDN U15838 ( .B(n7781), .A(n7782), .Z(n7756) );
  XNOR U15839 ( .A(n7747), .B(n7783), .Z(n7752) );
  XNOR U15840 ( .A(n7745), .B(n7749), .Z(n7783) );
  AND U15841 ( .A(n7784), .B(n7785), .Z(n7749) );
  NAND U15842 ( .A(n7786), .B(n7787), .Z(n7785) );
  NAND U15843 ( .A(n7788), .B(n7789), .Z(n7784) );
  AND U15844 ( .A(n7790), .B(n7791), .Z(n7745) );
  NAND U15845 ( .A(n7792), .B(n7793), .Z(n7791) );
  NAND U15846 ( .A(n7794), .B(n7795), .Z(n7790) );
  AND U15847 ( .A(n7796), .B(n7797), .Z(n7747) );
  NAND U15848 ( .A(n7798), .B(n7799), .Z(n7741) );
  XNOR U15849 ( .A(n7724), .B(n7800), .Z(n7738) );
  XNOR U15850 ( .A(n7728), .B(n7726), .Z(n7800) );
  XOR U15851 ( .A(n7734), .B(n7801), .Z(n7726) );
  XNOR U15852 ( .A(n7731), .B(n7735), .Z(n7801) );
  AND U15853 ( .A(n7802), .B(n7803), .Z(n7735) );
  NAND U15854 ( .A(n7804), .B(n7805), .Z(n7803) );
  NAND U15855 ( .A(n7806), .B(n7807), .Z(n7802) );
  AND U15856 ( .A(n7808), .B(n7809), .Z(n7731) );
  NAND U15857 ( .A(n7810), .B(n7811), .Z(n7809) );
  NAND U15858 ( .A(n7812), .B(n7813), .Z(n7808) );
  NANDN U15859 ( .A(n7814), .B(n7815), .Z(n7734) );
  ANDN U15860 ( .B(n7816), .A(n7817), .Z(n7728) );
  XNOR U15861 ( .A(n7719), .B(n7818), .Z(n7724) );
  XNOR U15862 ( .A(n7717), .B(n7721), .Z(n7818) );
  AND U15863 ( .A(n7819), .B(n7820), .Z(n7721) );
  NAND U15864 ( .A(n7821), .B(n7822), .Z(n7820) );
  NAND U15865 ( .A(n7823), .B(n7824), .Z(n7819) );
  AND U15866 ( .A(n7825), .B(n7826), .Z(n7717) );
  NAND U15867 ( .A(n7827), .B(n7828), .Z(n7826) );
  NAND U15868 ( .A(n7829), .B(n7830), .Z(n7825) );
  AND U15869 ( .A(n7831), .B(n7832), .Z(n7719) );
  XOR U15870 ( .A(n7799), .B(n7798), .Z(N64700) );
  XNOR U15871 ( .A(n7816), .B(n7817), .Z(n7798) );
  XNOR U15872 ( .A(n7831), .B(n7832), .Z(n7817) );
  XOR U15873 ( .A(n7828), .B(n7827), .Z(n7832) );
  XOR U15874 ( .A(y[7596]), .B(x[7596]), .Z(n7827) );
  XOR U15875 ( .A(n7830), .B(n7829), .Z(n7828) );
  XOR U15876 ( .A(y[7598]), .B(x[7598]), .Z(n7829) );
  XOR U15877 ( .A(y[7597]), .B(x[7597]), .Z(n7830) );
  XOR U15878 ( .A(n7822), .B(n7821), .Z(n7831) );
  XOR U15879 ( .A(n7824), .B(n7823), .Z(n7821) );
  XOR U15880 ( .A(y[7595]), .B(x[7595]), .Z(n7823) );
  XOR U15881 ( .A(y[7594]), .B(x[7594]), .Z(n7824) );
  XOR U15882 ( .A(y[7593]), .B(x[7593]), .Z(n7822) );
  XNOR U15883 ( .A(n7815), .B(n7814), .Z(n7816) );
  XNOR U15884 ( .A(n7811), .B(n7810), .Z(n7814) );
  XOR U15885 ( .A(n7813), .B(n7812), .Z(n7810) );
  XOR U15886 ( .A(y[7592]), .B(x[7592]), .Z(n7812) );
  XOR U15887 ( .A(y[7591]), .B(x[7591]), .Z(n7813) );
  XOR U15888 ( .A(y[7590]), .B(x[7590]), .Z(n7811) );
  XOR U15889 ( .A(n7805), .B(n7804), .Z(n7815) );
  XOR U15890 ( .A(n7807), .B(n7806), .Z(n7804) );
  XOR U15891 ( .A(y[7589]), .B(x[7589]), .Z(n7806) );
  XOR U15892 ( .A(y[7588]), .B(x[7588]), .Z(n7807) );
  XOR U15893 ( .A(y[7587]), .B(x[7587]), .Z(n7805) );
  XNOR U15894 ( .A(n7781), .B(n7782), .Z(n7799) );
  XNOR U15895 ( .A(n7796), .B(n7797), .Z(n7782) );
  XOR U15896 ( .A(n7793), .B(n7792), .Z(n7797) );
  XOR U15897 ( .A(y[7584]), .B(x[7584]), .Z(n7792) );
  XOR U15898 ( .A(n7795), .B(n7794), .Z(n7793) );
  XOR U15899 ( .A(y[7586]), .B(x[7586]), .Z(n7794) );
  XOR U15900 ( .A(y[7585]), .B(x[7585]), .Z(n7795) );
  XOR U15901 ( .A(n7787), .B(n7786), .Z(n7796) );
  XOR U15902 ( .A(n7789), .B(n7788), .Z(n7786) );
  XOR U15903 ( .A(y[7583]), .B(x[7583]), .Z(n7788) );
  XOR U15904 ( .A(y[7582]), .B(x[7582]), .Z(n7789) );
  XOR U15905 ( .A(y[7581]), .B(x[7581]), .Z(n7787) );
  XNOR U15906 ( .A(n7780), .B(n7779), .Z(n7781) );
  XNOR U15907 ( .A(n7776), .B(n7775), .Z(n7779) );
  XOR U15908 ( .A(n7778), .B(n7777), .Z(n7775) );
  XOR U15909 ( .A(y[7580]), .B(x[7580]), .Z(n7777) );
  XOR U15910 ( .A(y[7579]), .B(x[7579]), .Z(n7778) );
  XOR U15911 ( .A(y[7578]), .B(x[7578]), .Z(n7776) );
  XOR U15912 ( .A(n7770), .B(n7769), .Z(n7780) );
  XOR U15913 ( .A(n7772), .B(n7771), .Z(n7769) );
  XOR U15914 ( .A(y[7577]), .B(x[7577]), .Z(n7771) );
  XOR U15915 ( .A(y[7576]), .B(x[7576]), .Z(n7772) );
  XOR U15916 ( .A(y[7575]), .B(x[7575]), .Z(n7770) );
  NAND U15917 ( .A(n7833), .B(n7834), .Z(N64691) );
  NAND U15918 ( .A(n7835), .B(n7836), .Z(n7834) );
  NANDN U15919 ( .A(n7837), .B(n7838), .Z(n7836) );
  NANDN U15920 ( .A(n7838), .B(n7837), .Z(n7833) );
  XOR U15921 ( .A(n7837), .B(n7839), .Z(N64690) );
  XNOR U15922 ( .A(n7835), .B(n7838), .Z(n7839) );
  NAND U15923 ( .A(n7840), .B(n7841), .Z(n7838) );
  NAND U15924 ( .A(n7842), .B(n7843), .Z(n7841) );
  NANDN U15925 ( .A(n7844), .B(n7845), .Z(n7843) );
  NANDN U15926 ( .A(n7845), .B(n7844), .Z(n7840) );
  AND U15927 ( .A(n7846), .B(n7847), .Z(n7835) );
  NAND U15928 ( .A(n7848), .B(n7849), .Z(n7847) );
  NANDN U15929 ( .A(n7850), .B(n7851), .Z(n7849) );
  NANDN U15930 ( .A(n7851), .B(n7850), .Z(n7846) );
  IV U15931 ( .A(n7852), .Z(n7851) );
  AND U15932 ( .A(n7853), .B(n7854), .Z(n7837) );
  NAND U15933 ( .A(n7855), .B(n7856), .Z(n7854) );
  NANDN U15934 ( .A(n7857), .B(n7858), .Z(n7856) );
  NANDN U15935 ( .A(n7858), .B(n7857), .Z(n7853) );
  XOR U15936 ( .A(n7850), .B(n7859), .Z(N64689) );
  XNOR U15937 ( .A(n7848), .B(n7852), .Z(n7859) );
  XOR U15938 ( .A(n7845), .B(n7860), .Z(n7852) );
  XNOR U15939 ( .A(n7842), .B(n7844), .Z(n7860) );
  AND U15940 ( .A(n7861), .B(n7862), .Z(n7844) );
  NANDN U15941 ( .A(n7863), .B(n7864), .Z(n7862) );
  OR U15942 ( .A(n7865), .B(n7866), .Z(n7864) );
  IV U15943 ( .A(n7867), .Z(n7866) );
  NANDN U15944 ( .A(n7867), .B(n7865), .Z(n7861) );
  AND U15945 ( .A(n7868), .B(n7869), .Z(n7842) );
  NAND U15946 ( .A(n7870), .B(n7871), .Z(n7869) );
  NANDN U15947 ( .A(n7872), .B(n7873), .Z(n7871) );
  NANDN U15948 ( .A(n7873), .B(n7872), .Z(n7868) );
  IV U15949 ( .A(n7874), .Z(n7873) );
  NAND U15950 ( .A(n7875), .B(n7876), .Z(n7845) );
  NANDN U15951 ( .A(n7877), .B(n7878), .Z(n7876) );
  NANDN U15952 ( .A(n7879), .B(n7880), .Z(n7878) );
  NANDN U15953 ( .A(n7880), .B(n7879), .Z(n7875) );
  IV U15954 ( .A(n7881), .Z(n7879) );
  AND U15955 ( .A(n7882), .B(n7883), .Z(n7848) );
  NAND U15956 ( .A(n7884), .B(n7885), .Z(n7883) );
  NANDN U15957 ( .A(n7886), .B(n7887), .Z(n7885) );
  NANDN U15958 ( .A(n7887), .B(n7886), .Z(n7882) );
  XOR U15959 ( .A(n7858), .B(n7888), .Z(n7850) );
  XNOR U15960 ( .A(n7855), .B(n7857), .Z(n7888) );
  AND U15961 ( .A(n7889), .B(n7890), .Z(n7857) );
  NANDN U15962 ( .A(n7891), .B(n7892), .Z(n7890) );
  OR U15963 ( .A(n7893), .B(n7894), .Z(n7892) );
  IV U15964 ( .A(n7895), .Z(n7894) );
  NANDN U15965 ( .A(n7895), .B(n7893), .Z(n7889) );
  AND U15966 ( .A(n7896), .B(n7897), .Z(n7855) );
  NAND U15967 ( .A(n7898), .B(n7899), .Z(n7897) );
  NANDN U15968 ( .A(n7900), .B(n7901), .Z(n7899) );
  NANDN U15969 ( .A(n7901), .B(n7900), .Z(n7896) );
  IV U15970 ( .A(n7902), .Z(n7901) );
  NAND U15971 ( .A(n7903), .B(n7904), .Z(n7858) );
  NANDN U15972 ( .A(n7905), .B(n7906), .Z(n7904) );
  NANDN U15973 ( .A(n7907), .B(n7908), .Z(n7906) );
  NANDN U15974 ( .A(n7908), .B(n7907), .Z(n7903) );
  IV U15975 ( .A(n7909), .Z(n7907) );
  XOR U15976 ( .A(n7884), .B(n7910), .Z(N64688) );
  XNOR U15977 ( .A(n7887), .B(n7886), .Z(n7910) );
  XNOR U15978 ( .A(n7898), .B(n7911), .Z(n7886) );
  XNOR U15979 ( .A(n7902), .B(n7900), .Z(n7911) );
  XOR U15980 ( .A(n7908), .B(n7912), .Z(n7900) );
  XNOR U15981 ( .A(n7905), .B(n7909), .Z(n7912) );
  AND U15982 ( .A(n7913), .B(n7914), .Z(n7909) );
  NAND U15983 ( .A(n7915), .B(n7916), .Z(n7914) );
  NAND U15984 ( .A(n7917), .B(n7918), .Z(n7913) );
  AND U15985 ( .A(n7919), .B(n7920), .Z(n7905) );
  NAND U15986 ( .A(n7921), .B(n7922), .Z(n7920) );
  NAND U15987 ( .A(n7923), .B(n7924), .Z(n7919) );
  NANDN U15988 ( .A(n7925), .B(n7926), .Z(n7908) );
  ANDN U15989 ( .B(n7927), .A(n7928), .Z(n7902) );
  XNOR U15990 ( .A(n7893), .B(n7929), .Z(n7898) );
  XNOR U15991 ( .A(n7891), .B(n7895), .Z(n7929) );
  AND U15992 ( .A(n7930), .B(n7931), .Z(n7895) );
  NAND U15993 ( .A(n7932), .B(n7933), .Z(n7931) );
  NAND U15994 ( .A(n7934), .B(n7935), .Z(n7930) );
  AND U15995 ( .A(n7936), .B(n7937), .Z(n7891) );
  NAND U15996 ( .A(n7938), .B(n7939), .Z(n7937) );
  NAND U15997 ( .A(n7940), .B(n7941), .Z(n7936) );
  AND U15998 ( .A(n7942), .B(n7943), .Z(n7893) );
  NAND U15999 ( .A(n7944), .B(n7945), .Z(n7887) );
  XNOR U16000 ( .A(n7870), .B(n7946), .Z(n7884) );
  XNOR U16001 ( .A(n7874), .B(n7872), .Z(n7946) );
  XOR U16002 ( .A(n7880), .B(n7947), .Z(n7872) );
  XNOR U16003 ( .A(n7877), .B(n7881), .Z(n7947) );
  AND U16004 ( .A(n7948), .B(n7949), .Z(n7881) );
  NAND U16005 ( .A(n7950), .B(n7951), .Z(n7949) );
  NAND U16006 ( .A(n7952), .B(n7953), .Z(n7948) );
  AND U16007 ( .A(n7954), .B(n7955), .Z(n7877) );
  NAND U16008 ( .A(n7956), .B(n7957), .Z(n7955) );
  NAND U16009 ( .A(n7958), .B(n7959), .Z(n7954) );
  NANDN U16010 ( .A(n7960), .B(n7961), .Z(n7880) );
  ANDN U16011 ( .B(n7962), .A(n7963), .Z(n7874) );
  XNOR U16012 ( .A(n7865), .B(n7964), .Z(n7870) );
  XNOR U16013 ( .A(n7863), .B(n7867), .Z(n7964) );
  AND U16014 ( .A(n7965), .B(n7966), .Z(n7867) );
  NAND U16015 ( .A(n7967), .B(n7968), .Z(n7966) );
  NAND U16016 ( .A(n7969), .B(n7970), .Z(n7965) );
  AND U16017 ( .A(n7971), .B(n7972), .Z(n7863) );
  NAND U16018 ( .A(n7973), .B(n7974), .Z(n7972) );
  NAND U16019 ( .A(n7975), .B(n7976), .Z(n7971) );
  AND U16020 ( .A(n7977), .B(n7978), .Z(n7865) );
  XOR U16021 ( .A(n7945), .B(n7944), .Z(N64687) );
  XNOR U16022 ( .A(n7962), .B(n7963), .Z(n7944) );
  XNOR U16023 ( .A(n7977), .B(n7978), .Z(n7963) );
  XOR U16024 ( .A(n7974), .B(n7973), .Z(n7978) );
  XOR U16025 ( .A(y[7572]), .B(x[7572]), .Z(n7973) );
  XOR U16026 ( .A(n7976), .B(n7975), .Z(n7974) );
  XOR U16027 ( .A(y[7574]), .B(x[7574]), .Z(n7975) );
  XOR U16028 ( .A(y[7573]), .B(x[7573]), .Z(n7976) );
  XOR U16029 ( .A(n7968), .B(n7967), .Z(n7977) );
  XOR U16030 ( .A(n7970), .B(n7969), .Z(n7967) );
  XOR U16031 ( .A(y[7571]), .B(x[7571]), .Z(n7969) );
  XOR U16032 ( .A(y[7570]), .B(x[7570]), .Z(n7970) );
  XOR U16033 ( .A(y[7569]), .B(x[7569]), .Z(n7968) );
  XNOR U16034 ( .A(n7961), .B(n7960), .Z(n7962) );
  XNOR U16035 ( .A(n7957), .B(n7956), .Z(n7960) );
  XOR U16036 ( .A(n7959), .B(n7958), .Z(n7956) );
  XOR U16037 ( .A(y[7568]), .B(x[7568]), .Z(n7958) );
  XOR U16038 ( .A(y[7567]), .B(x[7567]), .Z(n7959) );
  XOR U16039 ( .A(y[7566]), .B(x[7566]), .Z(n7957) );
  XOR U16040 ( .A(n7951), .B(n7950), .Z(n7961) );
  XOR U16041 ( .A(n7953), .B(n7952), .Z(n7950) );
  XOR U16042 ( .A(y[7565]), .B(x[7565]), .Z(n7952) );
  XOR U16043 ( .A(y[7564]), .B(x[7564]), .Z(n7953) );
  XOR U16044 ( .A(y[7563]), .B(x[7563]), .Z(n7951) );
  XNOR U16045 ( .A(n7927), .B(n7928), .Z(n7945) );
  XNOR U16046 ( .A(n7942), .B(n7943), .Z(n7928) );
  XOR U16047 ( .A(n7939), .B(n7938), .Z(n7943) );
  XOR U16048 ( .A(y[7560]), .B(x[7560]), .Z(n7938) );
  XOR U16049 ( .A(n7941), .B(n7940), .Z(n7939) );
  XOR U16050 ( .A(y[7562]), .B(x[7562]), .Z(n7940) );
  XOR U16051 ( .A(y[7561]), .B(x[7561]), .Z(n7941) );
  XOR U16052 ( .A(n7933), .B(n7932), .Z(n7942) );
  XOR U16053 ( .A(n7935), .B(n7934), .Z(n7932) );
  XOR U16054 ( .A(y[7559]), .B(x[7559]), .Z(n7934) );
  XOR U16055 ( .A(y[7558]), .B(x[7558]), .Z(n7935) );
  XOR U16056 ( .A(y[7557]), .B(x[7557]), .Z(n7933) );
  XNOR U16057 ( .A(n7926), .B(n7925), .Z(n7927) );
  XNOR U16058 ( .A(n7922), .B(n7921), .Z(n7925) );
  XOR U16059 ( .A(n7924), .B(n7923), .Z(n7921) );
  XOR U16060 ( .A(y[7556]), .B(x[7556]), .Z(n7923) );
  XOR U16061 ( .A(y[7555]), .B(x[7555]), .Z(n7924) );
  XOR U16062 ( .A(y[7554]), .B(x[7554]), .Z(n7922) );
  XOR U16063 ( .A(n7916), .B(n7915), .Z(n7926) );
  XOR U16064 ( .A(n7918), .B(n7917), .Z(n7915) );
  XOR U16065 ( .A(y[7553]), .B(x[7553]), .Z(n7917) );
  XOR U16066 ( .A(y[7552]), .B(x[7552]), .Z(n7918) );
  XOR U16067 ( .A(y[7551]), .B(x[7551]), .Z(n7916) );
  NAND U16068 ( .A(n7979), .B(n7980), .Z(N64678) );
  NAND U16069 ( .A(n7981), .B(n7982), .Z(n7980) );
  NANDN U16070 ( .A(n7983), .B(n7984), .Z(n7982) );
  NANDN U16071 ( .A(n7984), .B(n7983), .Z(n7979) );
  XOR U16072 ( .A(n7983), .B(n7985), .Z(N64677) );
  XNOR U16073 ( .A(n7981), .B(n7984), .Z(n7985) );
  NAND U16074 ( .A(n7986), .B(n7987), .Z(n7984) );
  NAND U16075 ( .A(n7988), .B(n7989), .Z(n7987) );
  NANDN U16076 ( .A(n7990), .B(n7991), .Z(n7989) );
  NANDN U16077 ( .A(n7991), .B(n7990), .Z(n7986) );
  AND U16078 ( .A(n7992), .B(n7993), .Z(n7981) );
  NAND U16079 ( .A(n7994), .B(n7995), .Z(n7993) );
  NANDN U16080 ( .A(n7996), .B(n7997), .Z(n7995) );
  NANDN U16081 ( .A(n7997), .B(n7996), .Z(n7992) );
  IV U16082 ( .A(n7998), .Z(n7997) );
  AND U16083 ( .A(n7999), .B(n8000), .Z(n7983) );
  NAND U16084 ( .A(n8001), .B(n8002), .Z(n8000) );
  NANDN U16085 ( .A(n8003), .B(n8004), .Z(n8002) );
  NANDN U16086 ( .A(n8004), .B(n8003), .Z(n7999) );
  XOR U16087 ( .A(n7996), .B(n8005), .Z(N64676) );
  XNOR U16088 ( .A(n7994), .B(n7998), .Z(n8005) );
  XOR U16089 ( .A(n7991), .B(n8006), .Z(n7998) );
  XNOR U16090 ( .A(n7988), .B(n7990), .Z(n8006) );
  AND U16091 ( .A(n8007), .B(n8008), .Z(n7990) );
  NANDN U16092 ( .A(n8009), .B(n8010), .Z(n8008) );
  OR U16093 ( .A(n8011), .B(n8012), .Z(n8010) );
  IV U16094 ( .A(n8013), .Z(n8012) );
  NANDN U16095 ( .A(n8013), .B(n8011), .Z(n8007) );
  AND U16096 ( .A(n8014), .B(n8015), .Z(n7988) );
  NAND U16097 ( .A(n8016), .B(n8017), .Z(n8015) );
  NANDN U16098 ( .A(n8018), .B(n8019), .Z(n8017) );
  NANDN U16099 ( .A(n8019), .B(n8018), .Z(n8014) );
  IV U16100 ( .A(n8020), .Z(n8019) );
  NAND U16101 ( .A(n8021), .B(n8022), .Z(n7991) );
  NANDN U16102 ( .A(n8023), .B(n8024), .Z(n8022) );
  NANDN U16103 ( .A(n8025), .B(n8026), .Z(n8024) );
  NANDN U16104 ( .A(n8026), .B(n8025), .Z(n8021) );
  IV U16105 ( .A(n8027), .Z(n8025) );
  AND U16106 ( .A(n8028), .B(n8029), .Z(n7994) );
  NAND U16107 ( .A(n8030), .B(n8031), .Z(n8029) );
  NANDN U16108 ( .A(n8032), .B(n8033), .Z(n8031) );
  NANDN U16109 ( .A(n8033), .B(n8032), .Z(n8028) );
  XOR U16110 ( .A(n8004), .B(n8034), .Z(n7996) );
  XNOR U16111 ( .A(n8001), .B(n8003), .Z(n8034) );
  AND U16112 ( .A(n8035), .B(n8036), .Z(n8003) );
  NANDN U16113 ( .A(n8037), .B(n8038), .Z(n8036) );
  OR U16114 ( .A(n8039), .B(n8040), .Z(n8038) );
  IV U16115 ( .A(n8041), .Z(n8040) );
  NANDN U16116 ( .A(n8041), .B(n8039), .Z(n8035) );
  AND U16117 ( .A(n8042), .B(n8043), .Z(n8001) );
  NAND U16118 ( .A(n8044), .B(n8045), .Z(n8043) );
  NANDN U16119 ( .A(n8046), .B(n8047), .Z(n8045) );
  NANDN U16120 ( .A(n8047), .B(n8046), .Z(n8042) );
  IV U16121 ( .A(n8048), .Z(n8047) );
  NAND U16122 ( .A(n8049), .B(n8050), .Z(n8004) );
  NANDN U16123 ( .A(n8051), .B(n8052), .Z(n8050) );
  NANDN U16124 ( .A(n8053), .B(n8054), .Z(n8052) );
  NANDN U16125 ( .A(n8054), .B(n8053), .Z(n8049) );
  IV U16126 ( .A(n8055), .Z(n8053) );
  XOR U16127 ( .A(n8030), .B(n8056), .Z(N64675) );
  XNOR U16128 ( .A(n8033), .B(n8032), .Z(n8056) );
  XNOR U16129 ( .A(n8044), .B(n8057), .Z(n8032) );
  XNOR U16130 ( .A(n8048), .B(n8046), .Z(n8057) );
  XOR U16131 ( .A(n8054), .B(n8058), .Z(n8046) );
  XNOR U16132 ( .A(n8051), .B(n8055), .Z(n8058) );
  AND U16133 ( .A(n8059), .B(n8060), .Z(n8055) );
  NAND U16134 ( .A(n8061), .B(n8062), .Z(n8060) );
  NAND U16135 ( .A(n8063), .B(n8064), .Z(n8059) );
  AND U16136 ( .A(n8065), .B(n8066), .Z(n8051) );
  NAND U16137 ( .A(n8067), .B(n8068), .Z(n8066) );
  NAND U16138 ( .A(n8069), .B(n8070), .Z(n8065) );
  NANDN U16139 ( .A(n8071), .B(n8072), .Z(n8054) );
  ANDN U16140 ( .B(n8073), .A(n8074), .Z(n8048) );
  XNOR U16141 ( .A(n8039), .B(n8075), .Z(n8044) );
  XNOR U16142 ( .A(n8037), .B(n8041), .Z(n8075) );
  AND U16143 ( .A(n8076), .B(n8077), .Z(n8041) );
  NAND U16144 ( .A(n8078), .B(n8079), .Z(n8077) );
  NAND U16145 ( .A(n8080), .B(n8081), .Z(n8076) );
  AND U16146 ( .A(n8082), .B(n8083), .Z(n8037) );
  NAND U16147 ( .A(n8084), .B(n8085), .Z(n8083) );
  NAND U16148 ( .A(n8086), .B(n8087), .Z(n8082) );
  AND U16149 ( .A(n8088), .B(n8089), .Z(n8039) );
  NAND U16150 ( .A(n8090), .B(n8091), .Z(n8033) );
  XNOR U16151 ( .A(n8016), .B(n8092), .Z(n8030) );
  XNOR U16152 ( .A(n8020), .B(n8018), .Z(n8092) );
  XOR U16153 ( .A(n8026), .B(n8093), .Z(n8018) );
  XNOR U16154 ( .A(n8023), .B(n8027), .Z(n8093) );
  AND U16155 ( .A(n8094), .B(n8095), .Z(n8027) );
  NAND U16156 ( .A(n8096), .B(n8097), .Z(n8095) );
  NAND U16157 ( .A(n8098), .B(n8099), .Z(n8094) );
  AND U16158 ( .A(n8100), .B(n8101), .Z(n8023) );
  NAND U16159 ( .A(n8102), .B(n8103), .Z(n8101) );
  NAND U16160 ( .A(n8104), .B(n8105), .Z(n8100) );
  NANDN U16161 ( .A(n8106), .B(n8107), .Z(n8026) );
  ANDN U16162 ( .B(n8108), .A(n8109), .Z(n8020) );
  XNOR U16163 ( .A(n8011), .B(n8110), .Z(n8016) );
  XNOR U16164 ( .A(n8009), .B(n8013), .Z(n8110) );
  AND U16165 ( .A(n8111), .B(n8112), .Z(n8013) );
  NAND U16166 ( .A(n8113), .B(n8114), .Z(n8112) );
  NAND U16167 ( .A(n8115), .B(n8116), .Z(n8111) );
  AND U16168 ( .A(n8117), .B(n8118), .Z(n8009) );
  NAND U16169 ( .A(n8119), .B(n8120), .Z(n8118) );
  NAND U16170 ( .A(n8121), .B(n8122), .Z(n8117) );
  AND U16171 ( .A(n8123), .B(n8124), .Z(n8011) );
  XOR U16172 ( .A(n8091), .B(n8090), .Z(N64674) );
  XNOR U16173 ( .A(n8108), .B(n8109), .Z(n8090) );
  XNOR U16174 ( .A(n8123), .B(n8124), .Z(n8109) );
  XOR U16175 ( .A(n8120), .B(n8119), .Z(n8124) );
  XOR U16176 ( .A(y[7548]), .B(x[7548]), .Z(n8119) );
  XOR U16177 ( .A(n8122), .B(n8121), .Z(n8120) );
  XOR U16178 ( .A(y[7550]), .B(x[7550]), .Z(n8121) );
  XOR U16179 ( .A(y[7549]), .B(x[7549]), .Z(n8122) );
  XOR U16180 ( .A(n8114), .B(n8113), .Z(n8123) );
  XOR U16181 ( .A(n8116), .B(n8115), .Z(n8113) );
  XOR U16182 ( .A(y[7547]), .B(x[7547]), .Z(n8115) );
  XOR U16183 ( .A(y[7546]), .B(x[7546]), .Z(n8116) );
  XOR U16184 ( .A(y[7545]), .B(x[7545]), .Z(n8114) );
  XNOR U16185 ( .A(n8107), .B(n8106), .Z(n8108) );
  XNOR U16186 ( .A(n8103), .B(n8102), .Z(n8106) );
  XOR U16187 ( .A(n8105), .B(n8104), .Z(n8102) );
  XOR U16188 ( .A(y[7544]), .B(x[7544]), .Z(n8104) );
  XOR U16189 ( .A(y[7543]), .B(x[7543]), .Z(n8105) );
  XOR U16190 ( .A(y[7542]), .B(x[7542]), .Z(n8103) );
  XOR U16191 ( .A(n8097), .B(n8096), .Z(n8107) );
  XOR U16192 ( .A(n8099), .B(n8098), .Z(n8096) );
  XOR U16193 ( .A(y[7541]), .B(x[7541]), .Z(n8098) );
  XOR U16194 ( .A(y[7540]), .B(x[7540]), .Z(n8099) );
  XOR U16195 ( .A(y[7539]), .B(x[7539]), .Z(n8097) );
  XNOR U16196 ( .A(n8073), .B(n8074), .Z(n8091) );
  XNOR U16197 ( .A(n8088), .B(n8089), .Z(n8074) );
  XOR U16198 ( .A(n8085), .B(n8084), .Z(n8089) );
  XOR U16199 ( .A(y[7536]), .B(x[7536]), .Z(n8084) );
  XOR U16200 ( .A(n8087), .B(n8086), .Z(n8085) );
  XOR U16201 ( .A(y[7538]), .B(x[7538]), .Z(n8086) );
  XOR U16202 ( .A(y[7537]), .B(x[7537]), .Z(n8087) );
  XOR U16203 ( .A(n8079), .B(n8078), .Z(n8088) );
  XOR U16204 ( .A(n8081), .B(n8080), .Z(n8078) );
  XOR U16205 ( .A(y[7535]), .B(x[7535]), .Z(n8080) );
  XOR U16206 ( .A(y[7534]), .B(x[7534]), .Z(n8081) );
  XOR U16207 ( .A(y[7533]), .B(x[7533]), .Z(n8079) );
  XNOR U16208 ( .A(n8072), .B(n8071), .Z(n8073) );
  XNOR U16209 ( .A(n8068), .B(n8067), .Z(n8071) );
  XOR U16210 ( .A(n8070), .B(n8069), .Z(n8067) );
  XOR U16211 ( .A(y[7532]), .B(x[7532]), .Z(n8069) );
  XOR U16212 ( .A(y[7531]), .B(x[7531]), .Z(n8070) );
  XOR U16213 ( .A(y[7530]), .B(x[7530]), .Z(n8068) );
  XOR U16214 ( .A(n8062), .B(n8061), .Z(n8072) );
  XOR U16215 ( .A(n8064), .B(n8063), .Z(n8061) );
  XOR U16216 ( .A(y[7529]), .B(x[7529]), .Z(n8063) );
  XOR U16217 ( .A(y[7528]), .B(x[7528]), .Z(n8064) );
  XOR U16218 ( .A(y[7527]), .B(x[7527]), .Z(n8062) );
  NAND U16219 ( .A(n8125), .B(n8126), .Z(N64665) );
  NAND U16220 ( .A(n8127), .B(n8128), .Z(n8126) );
  NANDN U16221 ( .A(n8129), .B(n8130), .Z(n8128) );
  NANDN U16222 ( .A(n8130), .B(n8129), .Z(n8125) );
  XOR U16223 ( .A(n8129), .B(n8131), .Z(N64664) );
  XNOR U16224 ( .A(n8127), .B(n8130), .Z(n8131) );
  NAND U16225 ( .A(n8132), .B(n8133), .Z(n8130) );
  NAND U16226 ( .A(n8134), .B(n8135), .Z(n8133) );
  NANDN U16227 ( .A(n8136), .B(n8137), .Z(n8135) );
  NANDN U16228 ( .A(n8137), .B(n8136), .Z(n8132) );
  AND U16229 ( .A(n8138), .B(n8139), .Z(n8127) );
  NAND U16230 ( .A(n8140), .B(n8141), .Z(n8139) );
  NANDN U16231 ( .A(n8142), .B(n8143), .Z(n8141) );
  NANDN U16232 ( .A(n8143), .B(n8142), .Z(n8138) );
  IV U16233 ( .A(n8144), .Z(n8143) );
  AND U16234 ( .A(n8145), .B(n8146), .Z(n8129) );
  NAND U16235 ( .A(n8147), .B(n8148), .Z(n8146) );
  NANDN U16236 ( .A(n8149), .B(n8150), .Z(n8148) );
  NANDN U16237 ( .A(n8150), .B(n8149), .Z(n8145) );
  XOR U16238 ( .A(n8142), .B(n8151), .Z(N64663) );
  XNOR U16239 ( .A(n8140), .B(n8144), .Z(n8151) );
  XOR U16240 ( .A(n8137), .B(n8152), .Z(n8144) );
  XNOR U16241 ( .A(n8134), .B(n8136), .Z(n8152) );
  AND U16242 ( .A(n8153), .B(n8154), .Z(n8136) );
  NANDN U16243 ( .A(n8155), .B(n8156), .Z(n8154) );
  OR U16244 ( .A(n8157), .B(n8158), .Z(n8156) );
  IV U16245 ( .A(n8159), .Z(n8158) );
  NANDN U16246 ( .A(n8159), .B(n8157), .Z(n8153) );
  AND U16247 ( .A(n8160), .B(n8161), .Z(n8134) );
  NAND U16248 ( .A(n8162), .B(n8163), .Z(n8161) );
  NANDN U16249 ( .A(n8164), .B(n8165), .Z(n8163) );
  NANDN U16250 ( .A(n8165), .B(n8164), .Z(n8160) );
  IV U16251 ( .A(n8166), .Z(n8165) );
  NAND U16252 ( .A(n8167), .B(n8168), .Z(n8137) );
  NANDN U16253 ( .A(n8169), .B(n8170), .Z(n8168) );
  NANDN U16254 ( .A(n8171), .B(n8172), .Z(n8170) );
  NANDN U16255 ( .A(n8172), .B(n8171), .Z(n8167) );
  IV U16256 ( .A(n8173), .Z(n8171) );
  AND U16257 ( .A(n8174), .B(n8175), .Z(n8140) );
  NAND U16258 ( .A(n8176), .B(n8177), .Z(n8175) );
  NANDN U16259 ( .A(n8178), .B(n8179), .Z(n8177) );
  NANDN U16260 ( .A(n8179), .B(n8178), .Z(n8174) );
  XOR U16261 ( .A(n8150), .B(n8180), .Z(n8142) );
  XNOR U16262 ( .A(n8147), .B(n8149), .Z(n8180) );
  AND U16263 ( .A(n8181), .B(n8182), .Z(n8149) );
  NANDN U16264 ( .A(n8183), .B(n8184), .Z(n8182) );
  OR U16265 ( .A(n8185), .B(n8186), .Z(n8184) );
  IV U16266 ( .A(n8187), .Z(n8186) );
  NANDN U16267 ( .A(n8187), .B(n8185), .Z(n8181) );
  AND U16268 ( .A(n8188), .B(n8189), .Z(n8147) );
  NAND U16269 ( .A(n8190), .B(n8191), .Z(n8189) );
  NANDN U16270 ( .A(n8192), .B(n8193), .Z(n8191) );
  NANDN U16271 ( .A(n8193), .B(n8192), .Z(n8188) );
  IV U16272 ( .A(n8194), .Z(n8193) );
  NAND U16273 ( .A(n8195), .B(n8196), .Z(n8150) );
  NANDN U16274 ( .A(n8197), .B(n8198), .Z(n8196) );
  NANDN U16275 ( .A(n8199), .B(n8200), .Z(n8198) );
  NANDN U16276 ( .A(n8200), .B(n8199), .Z(n8195) );
  IV U16277 ( .A(n8201), .Z(n8199) );
  XOR U16278 ( .A(n8176), .B(n8202), .Z(N64662) );
  XNOR U16279 ( .A(n8179), .B(n8178), .Z(n8202) );
  XNOR U16280 ( .A(n8190), .B(n8203), .Z(n8178) );
  XNOR U16281 ( .A(n8194), .B(n8192), .Z(n8203) );
  XOR U16282 ( .A(n8200), .B(n8204), .Z(n8192) );
  XNOR U16283 ( .A(n8197), .B(n8201), .Z(n8204) );
  AND U16284 ( .A(n8205), .B(n8206), .Z(n8201) );
  NAND U16285 ( .A(n8207), .B(n8208), .Z(n8206) );
  NAND U16286 ( .A(n8209), .B(n8210), .Z(n8205) );
  AND U16287 ( .A(n8211), .B(n8212), .Z(n8197) );
  NAND U16288 ( .A(n8213), .B(n8214), .Z(n8212) );
  NAND U16289 ( .A(n8215), .B(n8216), .Z(n8211) );
  NANDN U16290 ( .A(n8217), .B(n8218), .Z(n8200) );
  ANDN U16291 ( .B(n8219), .A(n8220), .Z(n8194) );
  XNOR U16292 ( .A(n8185), .B(n8221), .Z(n8190) );
  XNOR U16293 ( .A(n8183), .B(n8187), .Z(n8221) );
  AND U16294 ( .A(n8222), .B(n8223), .Z(n8187) );
  NAND U16295 ( .A(n8224), .B(n8225), .Z(n8223) );
  NAND U16296 ( .A(n8226), .B(n8227), .Z(n8222) );
  AND U16297 ( .A(n8228), .B(n8229), .Z(n8183) );
  NAND U16298 ( .A(n8230), .B(n8231), .Z(n8229) );
  NAND U16299 ( .A(n8232), .B(n8233), .Z(n8228) );
  AND U16300 ( .A(n8234), .B(n8235), .Z(n8185) );
  NAND U16301 ( .A(n8236), .B(n8237), .Z(n8179) );
  XNOR U16302 ( .A(n8162), .B(n8238), .Z(n8176) );
  XNOR U16303 ( .A(n8166), .B(n8164), .Z(n8238) );
  XOR U16304 ( .A(n8172), .B(n8239), .Z(n8164) );
  XNOR U16305 ( .A(n8169), .B(n8173), .Z(n8239) );
  AND U16306 ( .A(n8240), .B(n8241), .Z(n8173) );
  NAND U16307 ( .A(n8242), .B(n8243), .Z(n8241) );
  NAND U16308 ( .A(n8244), .B(n8245), .Z(n8240) );
  AND U16309 ( .A(n8246), .B(n8247), .Z(n8169) );
  NAND U16310 ( .A(n8248), .B(n8249), .Z(n8247) );
  NAND U16311 ( .A(n8250), .B(n8251), .Z(n8246) );
  NANDN U16312 ( .A(n8252), .B(n8253), .Z(n8172) );
  ANDN U16313 ( .B(n8254), .A(n8255), .Z(n8166) );
  XNOR U16314 ( .A(n8157), .B(n8256), .Z(n8162) );
  XNOR U16315 ( .A(n8155), .B(n8159), .Z(n8256) );
  AND U16316 ( .A(n8257), .B(n8258), .Z(n8159) );
  NAND U16317 ( .A(n8259), .B(n8260), .Z(n8258) );
  NAND U16318 ( .A(n8261), .B(n8262), .Z(n8257) );
  AND U16319 ( .A(n8263), .B(n8264), .Z(n8155) );
  NAND U16320 ( .A(n8265), .B(n8266), .Z(n8264) );
  NAND U16321 ( .A(n8267), .B(n8268), .Z(n8263) );
  AND U16322 ( .A(n8269), .B(n8270), .Z(n8157) );
  XOR U16323 ( .A(n8237), .B(n8236), .Z(N64661) );
  XNOR U16324 ( .A(n8254), .B(n8255), .Z(n8236) );
  XNOR U16325 ( .A(n8269), .B(n8270), .Z(n8255) );
  XOR U16326 ( .A(n8266), .B(n8265), .Z(n8270) );
  XOR U16327 ( .A(y[7524]), .B(x[7524]), .Z(n8265) );
  XOR U16328 ( .A(n8268), .B(n8267), .Z(n8266) );
  XOR U16329 ( .A(y[7526]), .B(x[7526]), .Z(n8267) );
  XOR U16330 ( .A(y[7525]), .B(x[7525]), .Z(n8268) );
  XOR U16331 ( .A(n8260), .B(n8259), .Z(n8269) );
  XOR U16332 ( .A(n8262), .B(n8261), .Z(n8259) );
  XOR U16333 ( .A(y[7523]), .B(x[7523]), .Z(n8261) );
  XOR U16334 ( .A(y[7522]), .B(x[7522]), .Z(n8262) );
  XOR U16335 ( .A(y[7521]), .B(x[7521]), .Z(n8260) );
  XNOR U16336 ( .A(n8253), .B(n8252), .Z(n8254) );
  XNOR U16337 ( .A(n8249), .B(n8248), .Z(n8252) );
  XOR U16338 ( .A(n8251), .B(n8250), .Z(n8248) );
  XOR U16339 ( .A(y[7520]), .B(x[7520]), .Z(n8250) );
  XOR U16340 ( .A(y[7519]), .B(x[7519]), .Z(n8251) );
  XOR U16341 ( .A(y[7518]), .B(x[7518]), .Z(n8249) );
  XOR U16342 ( .A(n8243), .B(n8242), .Z(n8253) );
  XOR U16343 ( .A(n8245), .B(n8244), .Z(n8242) );
  XOR U16344 ( .A(y[7517]), .B(x[7517]), .Z(n8244) );
  XOR U16345 ( .A(y[7516]), .B(x[7516]), .Z(n8245) );
  XOR U16346 ( .A(y[7515]), .B(x[7515]), .Z(n8243) );
  XNOR U16347 ( .A(n8219), .B(n8220), .Z(n8237) );
  XNOR U16348 ( .A(n8234), .B(n8235), .Z(n8220) );
  XOR U16349 ( .A(n8231), .B(n8230), .Z(n8235) );
  XOR U16350 ( .A(y[7512]), .B(x[7512]), .Z(n8230) );
  XOR U16351 ( .A(n8233), .B(n8232), .Z(n8231) );
  XOR U16352 ( .A(y[7514]), .B(x[7514]), .Z(n8232) );
  XOR U16353 ( .A(y[7513]), .B(x[7513]), .Z(n8233) );
  XOR U16354 ( .A(n8225), .B(n8224), .Z(n8234) );
  XOR U16355 ( .A(n8227), .B(n8226), .Z(n8224) );
  XOR U16356 ( .A(y[7511]), .B(x[7511]), .Z(n8226) );
  XOR U16357 ( .A(y[7510]), .B(x[7510]), .Z(n8227) );
  XOR U16358 ( .A(y[7509]), .B(x[7509]), .Z(n8225) );
  XNOR U16359 ( .A(n8218), .B(n8217), .Z(n8219) );
  XNOR U16360 ( .A(n8214), .B(n8213), .Z(n8217) );
  XOR U16361 ( .A(n8216), .B(n8215), .Z(n8213) );
  XOR U16362 ( .A(y[7508]), .B(x[7508]), .Z(n8215) );
  XOR U16363 ( .A(y[7507]), .B(x[7507]), .Z(n8216) );
  XOR U16364 ( .A(y[7506]), .B(x[7506]), .Z(n8214) );
  XOR U16365 ( .A(n8208), .B(n8207), .Z(n8218) );
  XOR U16366 ( .A(n8210), .B(n8209), .Z(n8207) );
  XOR U16367 ( .A(y[7505]), .B(x[7505]), .Z(n8209) );
  XOR U16368 ( .A(y[7504]), .B(x[7504]), .Z(n8210) );
  XOR U16369 ( .A(y[7503]), .B(x[7503]), .Z(n8208) );
  NAND U16370 ( .A(n8271), .B(n8272), .Z(N64652) );
  NAND U16371 ( .A(n8273), .B(n8274), .Z(n8272) );
  NANDN U16372 ( .A(n8275), .B(n8276), .Z(n8274) );
  NANDN U16373 ( .A(n8276), .B(n8275), .Z(n8271) );
  XOR U16374 ( .A(n8275), .B(n8277), .Z(N64651) );
  XNOR U16375 ( .A(n8273), .B(n8276), .Z(n8277) );
  NAND U16376 ( .A(n8278), .B(n8279), .Z(n8276) );
  NAND U16377 ( .A(n8280), .B(n8281), .Z(n8279) );
  NANDN U16378 ( .A(n8282), .B(n8283), .Z(n8281) );
  NANDN U16379 ( .A(n8283), .B(n8282), .Z(n8278) );
  AND U16380 ( .A(n8284), .B(n8285), .Z(n8273) );
  NAND U16381 ( .A(n8286), .B(n8287), .Z(n8285) );
  NANDN U16382 ( .A(n8288), .B(n8289), .Z(n8287) );
  NANDN U16383 ( .A(n8289), .B(n8288), .Z(n8284) );
  IV U16384 ( .A(n8290), .Z(n8289) );
  AND U16385 ( .A(n8291), .B(n8292), .Z(n8275) );
  NAND U16386 ( .A(n8293), .B(n8294), .Z(n8292) );
  NANDN U16387 ( .A(n8295), .B(n8296), .Z(n8294) );
  NANDN U16388 ( .A(n8296), .B(n8295), .Z(n8291) );
  XOR U16389 ( .A(n8288), .B(n8297), .Z(N64650) );
  XNOR U16390 ( .A(n8286), .B(n8290), .Z(n8297) );
  XOR U16391 ( .A(n8283), .B(n8298), .Z(n8290) );
  XNOR U16392 ( .A(n8280), .B(n8282), .Z(n8298) );
  AND U16393 ( .A(n8299), .B(n8300), .Z(n8282) );
  NANDN U16394 ( .A(n8301), .B(n8302), .Z(n8300) );
  OR U16395 ( .A(n8303), .B(n8304), .Z(n8302) );
  IV U16396 ( .A(n8305), .Z(n8304) );
  NANDN U16397 ( .A(n8305), .B(n8303), .Z(n8299) );
  AND U16398 ( .A(n8306), .B(n8307), .Z(n8280) );
  NAND U16399 ( .A(n8308), .B(n8309), .Z(n8307) );
  NANDN U16400 ( .A(n8310), .B(n8311), .Z(n8309) );
  NANDN U16401 ( .A(n8311), .B(n8310), .Z(n8306) );
  IV U16402 ( .A(n8312), .Z(n8311) );
  NAND U16403 ( .A(n8313), .B(n8314), .Z(n8283) );
  NANDN U16404 ( .A(n8315), .B(n8316), .Z(n8314) );
  NANDN U16405 ( .A(n8317), .B(n8318), .Z(n8316) );
  NANDN U16406 ( .A(n8318), .B(n8317), .Z(n8313) );
  IV U16407 ( .A(n8319), .Z(n8317) );
  AND U16408 ( .A(n8320), .B(n8321), .Z(n8286) );
  NAND U16409 ( .A(n8322), .B(n8323), .Z(n8321) );
  NANDN U16410 ( .A(n8324), .B(n8325), .Z(n8323) );
  NANDN U16411 ( .A(n8325), .B(n8324), .Z(n8320) );
  XOR U16412 ( .A(n8296), .B(n8326), .Z(n8288) );
  XNOR U16413 ( .A(n8293), .B(n8295), .Z(n8326) );
  AND U16414 ( .A(n8327), .B(n8328), .Z(n8295) );
  NANDN U16415 ( .A(n8329), .B(n8330), .Z(n8328) );
  OR U16416 ( .A(n8331), .B(n8332), .Z(n8330) );
  IV U16417 ( .A(n8333), .Z(n8332) );
  NANDN U16418 ( .A(n8333), .B(n8331), .Z(n8327) );
  AND U16419 ( .A(n8334), .B(n8335), .Z(n8293) );
  NAND U16420 ( .A(n8336), .B(n8337), .Z(n8335) );
  NANDN U16421 ( .A(n8338), .B(n8339), .Z(n8337) );
  NANDN U16422 ( .A(n8339), .B(n8338), .Z(n8334) );
  IV U16423 ( .A(n8340), .Z(n8339) );
  NAND U16424 ( .A(n8341), .B(n8342), .Z(n8296) );
  NANDN U16425 ( .A(n8343), .B(n8344), .Z(n8342) );
  NANDN U16426 ( .A(n8345), .B(n8346), .Z(n8344) );
  NANDN U16427 ( .A(n8346), .B(n8345), .Z(n8341) );
  IV U16428 ( .A(n8347), .Z(n8345) );
  XOR U16429 ( .A(n8322), .B(n8348), .Z(N64649) );
  XNOR U16430 ( .A(n8325), .B(n8324), .Z(n8348) );
  XNOR U16431 ( .A(n8336), .B(n8349), .Z(n8324) );
  XNOR U16432 ( .A(n8340), .B(n8338), .Z(n8349) );
  XOR U16433 ( .A(n8346), .B(n8350), .Z(n8338) );
  XNOR U16434 ( .A(n8343), .B(n8347), .Z(n8350) );
  AND U16435 ( .A(n8351), .B(n8352), .Z(n8347) );
  NAND U16436 ( .A(n8353), .B(n8354), .Z(n8352) );
  NAND U16437 ( .A(n8355), .B(n8356), .Z(n8351) );
  AND U16438 ( .A(n8357), .B(n8358), .Z(n8343) );
  NAND U16439 ( .A(n8359), .B(n8360), .Z(n8358) );
  NAND U16440 ( .A(n8361), .B(n8362), .Z(n8357) );
  NANDN U16441 ( .A(n8363), .B(n8364), .Z(n8346) );
  ANDN U16442 ( .B(n8365), .A(n8366), .Z(n8340) );
  XNOR U16443 ( .A(n8331), .B(n8367), .Z(n8336) );
  XNOR U16444 ( .A(n8329), .B(n8333), .Z(n8367) );
  AND U16445 ( .A(n8368), .B(n8369), .Z(n8333) );
  NAND U16446 ( .A(n8370), .B(n8371), .Z(n8369) );
  NAND U16447 ( .A(n8372), .B(n8373), .Z(n8368) );
  AND U16448 ( .A(n8374), .B(n8375), .Z(n8329) );
  NAND U16449 ( .A(n8376), .B(n8377), .Z(n8375) );
  NAND U16450 ( .A(n8378), .B(n8379), .Z(n8374) );
  AND U16451 ( .A(n8380), .B(n8381), .Z(n8331) );
  NAND U16452 ( .A(n8382), .B(n8383), .Z(n8325) );
  XNOR U16453 ( .A(n8308), .B(n8384), .Z(n8322) );
  XNOR U16454 ( .A(n8312), .B(n8310), .Z(n8384) );
  XOR U16455 ( .A(n8318), .B(n8385), .Z(n8310) );
  XNOR U16456 ( .A(n8315), .B(n8319), .Z(n8385) );
  AND U16457 ( .A(n8386), .B(n8387), .Z(n8319) );
  NAND U16458 ( .A(n8388), .B(n8389), .Z(n8387) );
  NAND U16459 ( .A(n8390), .B(n8391), .Z(n8386) );
  AND U16460 ( .A(n8392), .B(n8393), .Z(n8315) );
  NAND U16461 ( .A(n8394), .B(n8395), .Z(n8393) );
  NAND U16462 ( .A(n8396), .B(n8397), .Z(n8392) );
  NANDN U16463 ( .A(n8398), .B(n8399), .Z(n8318) );
  ANDN U16464 ( .B(n8400), .A(n8401), .Z(n8312) );
  XNOR U16465 ( .A(n8303), .B(n8402), .Z(n8308) );
  XNOR U16466 ( .A(n8301), .B(n8305), .Z(n8402) );
  AND U16467 ( .A(n8403), .B(n8404), .Z(n8305) );
  NAND U16468 ( .A(n8405), .B(n8406), .Z(n8404) );
  NAND U16469 ( .A(n8407), .B(n8408), .Z(n8403) );
  AND U16470 ( .A(n8409), .B(n8410), .Z(n8301) );
  NAND U16471 ( .A(n8411), .B(n8412), .Z(n8410) );
  NAND U16472 ( .A(n8413), .B(n8414), .Z(n8409) );
  AND U16473 ( .A(n8415), .B(n8416), .Z(n8303) );
  XOR U16474 ( .A(n8383), .B(n8382), .Z(N64648) );
  XNOR U16475 ( .A(n8400), .B(n8401), .Z(n8382) );
  XNOR U16476 ( .A(n8415), .B(n8416), .Z(n8401) );
  XOR U16477 ( .A(n8412), .B(n8411), .Z(n8416) );
  XOR U16478 ( .A(y[7500]), .B(x[7500]), .Z(n8411) );
  XOR U16479 ( .A(n8414), .B(n8413), .Z(n8412) );
  XOR U16480 ( .A(y[7502]), .B(x[7502]), .Z(n8413) );
  XOR U16481 ( .A(y[7501]), .B(x[7501]), .Z(n8414) );
  XOR U16482 ( .A(n8406), .B(n8405), .Z(n8415) );
  XOR U16483 ( .A(n8408), .B(n8407), .Z(n8405) );
  XOR U16484 ( .A(y[7499]), .B(x[7499]), .Z(n8407) );
  XOR U16485 ( .A(y[7498]), .B(x[7498]), .Z(n8408) );
  XOR U16486 ( .A(y[7497]), .B(x[7497]), .Z(n8406) );
  XNOR U16487 ( .A(n8399), .B(n8398), .Z(n8400) );
  XNOR U16488 ( .A(n8395), .B(n8394), .Z(n8398) );
  XOR U16489 ( .A(n8397), .B(n8396), .Z(n8394) );
  XOR U16490 ( .A(y[7496]), .B(x[7496]), .Z(n8396) );
  XOR U16491 ( .A(y[7495]), .B(x[7495]), .Z(n8397) );
  XOR U16492 ( .A(y[7494]), .B(x[7494]), .Z(n8395) );
  XOR U16493 ( .A(n8389), .B(n8388), .Z(n8399) );
  XOR U16494 ( .A(n8391), .B(n8390), .Z(n8388) );
  XOR U16495 ( .A(y[7493]), .B(x[7493]), .Z(n8390) );
  XOR U16496 ( .A(y[7492]), .B(x[7492]), .Z(n8391) );
  XOR U16497 ( .A(y[7491]), .B(x[7491]), .Z(n8389) );
  XNOR U16498 ( .A(n8365), .B(n8366), .Z(n8383) );
  XNOR U16499 ( .A(n8380), .B(n8381), .Z(n8366) );
  XOR U16500 ( .A(n8377), .B(n8376), .Z(n8381) );
  XOR U16501 ( .A(y[7488]), .B(x[7488]), .Z(n8376) );
  XOR U16502 ( .A(n8379), .B(n8378), .Z(n8377) );
  XOR U16503 ( .A(y[7490]), .B(x[7490]), .Z(n8378) );
  XOR U16504 ( .A(y[7489]), .B(x[7489]), .Z(n8379) );
  XOR U16505 ( .A(n8371), .B(n8370), .Z(n8380) );
  XOR U16506 ( .A(n8373), .B(n8372), .Z(n8370) );
  XOR U16507 ( .A(y[7487]), .B(x[7487]), .Z(n8372) );
  XOR U16508 ( .A(y[7486]), .B(x[7486]), .Z(n8373) );
  XOR U16509 ( .A(y[7485]), .B(x[7485]), .Z(n8371) );
  XNOR U16510 ( .A(n8364), .B(n8363), .Z(n8365) );
  XNOR U16511 ( .A(n8360), .B(n8359), .Z(n8363) );
  XOR U16512 ( .A(n8362), .B(n8361), .Z(n8359) );
  XOR U16513 ( .A(y[7484]), .B(x[7484]), .Z(n8361) );
  XOR U16514 ( .A(y[7483]), .B(x[7483]), .Z(n8362) );
  XOR U16515 ( .A(y[7482]), .B(x[7482]), .Z(n8360) );
  XOR U16516 ( .A(n8354), .B(n8353), .Z(n8364) );
  XOR U16517 ( .A(n8356), .B(n8355), .Z(n8353) );
  XOR U16518 ( .A(y[7481]), .B(x[7481]), .Z(n8355) );
  XOR U16519 ( .A(y[7480]), .B(x[7480]), .Z(n8356) );
  XOR U16520 ( .A(y[7479]), .B(x[7479]), .Z(n8354) );
  NAND U16521 ( .A(n8417), .B(n8418), .Z(N64639) );
  NAND U16522 ( .A(n8419), .B(n8420), .Z(n8418) );
  NANDN U16523 ( .A(n8421), .B(n8422), .Z(n8420) );
  NANDN U16524 ( .A(n8422), .B(n8421), .Z(n8417) );
  XOR U16525 ( .A(n8421), .B(n8423), .Z(N64638) );
  XNOR U16526 ( .A(n8419), .B(n8422), .Z(n8423) );
  NAND U16527 ( .A(n8424), .B(n8425), .Z(n8422) );
  NAND U16528 ( .A(n8426), .B(n8427), .Z(n8425) );
  NANDN U16529 ( .A(n8428), .B(n8429), .Z(n8427) );
  NANDN U16530 ( .A(n8429), .B(n8428), .Z(n8424) );
  AND U16531 ( .A(n8430), .B(n8431), .Z(n8419) );
  NAND U16532 ( .A(n8432), .B(n8433), .Z(n8431) );
  NANDN U16533 ( .A(n8434), .B(n8435), .Z(n8433) );
  NANDN U16534 ( .A(n8435), .B(n8434), .Z(n8430) );
  IV U16535 ( .A(n8436), .Z(n8435) );
  AND U16536 ( .A(n8437), .B(n8438), .Z(n8421) );
  NAND U16537 ( .A(n8439), .B(n8440), .Z(n8438) );
  NANDN U16538 ( .A(n8441), .B(n8442), .Z(n8440) );
  NANDN U16539 ( .A(n8442), .B(n8441), .Z(n8437) );
  XOR U16540 ( .A(n8434), .B(n8443), .Z(N64637) );
  XNOR U16541 ( .A(n8432), .B(n8436), .Z(n8443) );
  XOR U16542 ( .A(n8429), .B(n8444), .Z(n8436) );
  XNOR U16543 ( .A(n8426), .B(n8428), .Z(n8444) );
  AND U16544 ( .A(n8445), .B(n8446), .Z(n8428) );
  NANDN U16545 ( .A(n8447), .B(n8448), .Z(n8446) );
  OR U16546 ( .A(n8449), .B(n8450), .Z(n8448) );
  IV U16547 ( .A(n8451), .Z(n8450) );
  NANDN U16548 ( .A(n8451), .B(n8449), .Z(n8445) );
  AND U16549 ( .A(n8452), .B(n8453), .Z(n8426) );
  NAND U16550 ( .A(n8454), .B(n8455), .Z(n8453) );
  NANDN U16551 ( .A(n8456), .B(n8457), .Z(n8455) );
  NANDN U16552 ( .A(n8457), .B(n8456), .Z(n8452) );
  IV U16553 ( .A(n8458), .Z(n8457) );
  NAND U16554 ( .A(n8459), .B(n8460), .Z(n8429) );
  NANDN U16555 ( .A(n8461), .B(n8462), .Z(n8460) );
  NANDN U16556 ( .A(n8463), .B(n8464), .Z(n8462) );
  NANDN U16557 ( .A(n8464), .B(n8463), .Z(n8459) );
  IV U16558 ( .A(n8465), .Z(n8463) );
  AND U16559 ( .A(n8466), .B(n8467), .Z(n8432) );
  NAND U16560 ( .A(n8468), .B(n8469), .Z(n8467) );
  NANDN U16561 ( .A(n8470), .B(n8471), .Z(n8469) );
  NANDN U16562 ( .A(n8471), .B(n8470), .Z(n8466) );
  XOR U16563 ( .A(n8442), .B(n8472), .Z(n8434) );
  XNOR U16564 ( .A(n8439), .B(n8441), .Z(n8472) );
  AND U16565 ( .A(n8473), .B(n8474), .Z(n8441) );
  NANDN U16566 ( .A(n8475), .B(n8476), .Z(n8474) );
  OR U16567 ( .A(n8477), .B(n8478), .Z(n8476) );
  IV U16568 ( .A(n8479), .Z(n8478) );
  NANDN U16569 ( .A(n8479), .B(n8477), .Z(n8473) );
  AND U16570 ( .A(n8480), .B(n8481), .Z(n8439) );
  NAND U16571 ( .A(n8482), .B(n8483), .Z(n8481) );
  NANDN U16572 ( .A(n8484), .B(n8485), .Z(n8483) );
  NANDN U16573 ( .A(n8485), .B(n8484), .Z(n8480) );
  IV U16574 ( .A(n8486), .Z(n8485) );
  NAND U16575 ( .A(n8487), .B(n8488), .Z(n8442) );
  NANDN U16576 ( .A(n8489), .B(n8490), .Z(n8488) );
  NANDN U16577 ( .A(n8491), .B(n8492), .Z(n8490) );
  NANDN U16578 ( .A(n8492), .B(n8491), .Z(n8487) );
  IV U16579 ( .A(n8493), .Z(n8491) );
  XOR U16580 ( .A(n8468), .B(n8494), .Z(N64636) );
  XNOR U16581 ( .A(n8471), .B(n8470), .Z(n8494) );
  XNOR U16582 ( .A(n8482), .B(n8495), .Z(n8470) );
  XNOR U16583 ( .A(n8486), .B(n8484), .Z(n8495) );
  XOR U16584 ( .A(n8492), .B(n8496), .Z(n8484) );
  XNOR U16585 ( .A(n8489), .B(n8493), .Z(n8496) );
  AND U16586 ( .A(n8497), .B(n8498), .Z(n8493) );
  NAND U16587 ( .A(n8499), .B(n8500), .Z(n8498) );
  NAND U16588 ( .A(n8501), .B(n8502), .Z(n8497) );
  AND U16589 ( .A(n8503), .B(n8504), .Z(n8489) );
  NAND U16590 ( .A(n8505), .B(n8506), .Z(n8504) );
  NAND U16591 ( .A(n8507), .B(n8508), .Z(n8503) );
  NANDN U16592 ( .A(n8509), .B(n8510), .Z(n8492) );
  ANDN U16593 ( .B(n8511), .A(n8512), .Z(n8486) );
  XNOR U16594 ( .A(n8477), .B(n8513), .Z(n8482) );
  XNOR U16595 ( .A(n8475), .B(n8479), .Z(n8513) );
  AND U16596 ( .A(n8514), .B(n8515), .Z(n8479) );
  NAND U16597 ( .A(n8516), .B(n8517), .Z(n8515) );
  NAND U16598 ( .A(n8518), .B(n8519), .Z(n8514) );
  AND U16599 ( .A(n8520), .B(n8521), .Z(n8475) );
  NAND U16600 ( .A(n8522), .B(n8523), .Z(n8521) );
  NAND U16601 ( .A(n8524), .B(n8525), .Z(n8520) );
  AND U16602 ( .A(n8526), .B(n8527), .Z(n8477) );
  NAND U16603 ( .A(n8528), .B(n8529), .Z(n8471) );
  XNOR U16604 ( .A(n8454), .B(n8530), .Z(n8468) );
  XNOR U16605 ( .A(n8458), .B(n8456), .Z(n8530) );
  XOR U16606 ( .A(n8464), .B(n8531), .Z(n8456) );
  XNOR U16607 ( .A(n8461), .B(n8465), .Z(n8531) );
  AND U16608 ( .A(n8532), .B(n8533), .Z(n8465) );
  NAND U16609 ( .A(n8534), .B(n8535), .Z(n8533) );
  NAND U16610 ( .A(n8536), .B(n8537), .Z(n8532) );
  AND U16611 ( .A(n8538), .B(n8539), .Z(n8461) );
  NAND U16612 ( .A(n8540), .B(n8541), .Z(n8539) );
  NAND U16613 ( .A(n8542), .B(n8543), .Z(n8538) );
  NANDN U16614 ( .A(n8544), .B(n8545), .Z(n8464) );
  ANDN U16615 ( .B(n8546), .A(n8547), .Z(n8458) );
  XNOR U16616 ( .A(n8449), .B(n8548), .Z(n8454) );
  XNOR U16617 ( .A(n8447), .B(n8451), .Z(n8548) );
  AND U16618 ( .A(n8549), .B(n8550), .Z(n8451) );
  NAND U16619 ( .A(n8551), .B(n8552), .Z(n8550) );
  NAND U16620 ( .A(n8553), .B(n8554), .Z(n8549) );
  AND U16621 ( .A(n8555), .B(n8556), .Z(n8447) );
  NAND U16622 ( .A(n8557), .B(n8558), .Z(n8556) );
  NAND U16623 ( .A(n8559), .B(n8560), .Z(n8555) );
  AND U16624 ( .A(n8561), .B(n8562), .Z(n8449) );
  XOR U16625 ( .A(n8529), .B(n8528), .Z(N64635) );
  XNOR U16626 ( .A(n8546), .B(n8547), .Z(n8528) );
  XNOR U16627 ( .A(n8561), .B(n8562), .Z(n8547) );
  XOR U16628 ( .A(n8558), .B(n8557), .Z(n8562) );
  XOR U16629 ( .A(y[7476]), .B(x[7476]), .Z(n8557) );
  XOR U16630 ( .A(n8560), .B(n8559), .Z(n8558) );
  XOR U16631 ( .A(y[7478]), .B(x[7478]), .Z(n8559) );
  XOR U16632 ( .A(y[7477]), .B(x[7477]), .Z(n8560) );
  XOR U16633 ( .A(n8552), .B(n8551), .Z(n8561) );
  XOR U16634 ( .A(n8554), .B(n8553), .Z(n8551) );
  XOR U16635 ( .A(y[7475]), .B(x[7475]), .Z(n8553) );
  XOR U16636 ( .A(y[7474]), .B(x[7474]), .Z(n8554) );
  XOR U16637 ( .A(y[7473]), .B(x[7473]), .Z(n8552) );
  XNOR U16638 ( .A(n8545), .B(n8544), .Z(n8546) );
  XNOR U16639 ( .A(n8541), .B(n8540), .Z(n8544) );
  XOR U16640 ( .A(n8543), .B(n8542), .Z(n8540) );
  XOR U16641 ( .A(y[7472]), .B(x[7472]), .Z(n8542) );
  XOR U16642 ( .A(y[7471]), .B(x[7471]), .Z(n8543) );
  XOR U16643 ( .A(y[7470]), .B(x[7470]), .Z(n8541) );
  XOR U16644 ( .A(n8535), .B(n8534), .Z(n8545) );
  XOR U16645 ( .A(n8537), .B(n8536), .Z(n8534) );
  XOR U16646 ( .A(y[7469]), .B(x[7469]), .Z(n8536) );
  XOR U16647 ( .A(y[7468]), .B(x[7468]), .Z(n8537) );
  XOR U16648 ( .A(y[7467]), .B(x[7467]), .Z(n8535) );
  XNOR U16649 ( .A(n8511), .B(n8512), .Z(n8529) );
  XNOR U16650 ( .A(n8526), .B(n8527), .Z(n8512) );
  XOR U16651 ( .A(n8523), .B(n8522), .Z(n8527) );
  XOR U16652 ( .A(y[7464]), .B(x[7464]), .Z(n8522) );
  XOR U16653 ( .A(n8525), .B(n8524), .Z(n8523) );
  XOR U16654 ( .A(y[7466]), .B(x[7466]), .Z(n8524) );
  XOR U16655 ( .A(y[7465]), .B(x[7465]), .Z(n8525) );
  XOR U16656 ( .A(n8517), .B(n8516), .Z(n8526) );
  XOR U16657 ( .A(n8519), .B(n8518), .Z(n8516) );
  XOR U16658 ( .A(y[7463]), .B(x[7463]), .Z(n8518) );
  XOR U16659 ( .A(y[7462]), .B(x[7462]), .Z(n8519) );
  XOR U16660 ( .A(y[7461]), .B(x[7461]), .Z(n8517) );
  XNOR U16661 ( .A(n8510), .B(n8509), .Z(n8511) );
  XNOR U16662 ( .A(n8506), .B(n8505), .Z(n8509) );
  XOR U16663 ( .A(n8508), .B(n8507), .Z(n8505) );
  XOR U16664 ( .A(y[7460]), .B(x[7460]), .Z(n8507) );
  XOR U16665 ( .A(y[7459]), .B(x[7459]), .Z(n8508) );
  XOR U16666 ( .A(y[7458]), .B(x[7458]), .Z(n8506) );
  XOR U16667 ( .A(n8500), .B(n8499), .Z(n8510) );
  XOR U16668 ( .A(n8502), .B(n8501), .Z(n8499) );
  XOR U16669 ( .A(y[7457]), .B(x[7457]), .Z(n8501) );
  XOR U16670 ( .A(y[7456]), .B(x[7456]), .Z(n8502) );
  XOR U16671 ( .A(y[7455]), .B(x[7455]), .Z(n8500) );
  NAND U16672 ( .A(n8563), .B(n8564), .Z(N64626) );
  NAND U16673 ( .A(n8565), .B(n8566), .Z(n8564) );
  NANDN U16674 ( .A(n8567), .B(n8568), .Z(n8566) );
  NANDN U16675 ( .A(n8568), .B(n8567), .Z(n8563) );
  XOR U16676 ( .A(n8567), .B(n8569), .Z(N64625) );
  XNOR U16677 ( .A(n8565), .B(n8568), .Z(n8569) );
  NAND U16678 ( .A(n8570), .B(n8571), .Z(n8568) );
  NAND U16679 ( .A(n8572), .B(n8573), .Z(n8571) );
  NANDN U16680 ( .A(n8574), .B(n8575), .Z(n8573) );
  NANDN U16681 ( .A(n8575), .B(n8574), .Z(n8570) );
  AND U16682 ( .A(n8576), .B(n8577), .Z(n8565) );
  NAND U16683 ( .A(n8578), .B(n8579), .Z(n8577) );
  NANDN U16684 ( .A(n8580), .B(n8581), .Z(n8579) );
  NANDN U16685 ( .A(n8581), .B(n8580), .Z(n8576) );
  IV U16686 ( .A(n8582), .Z(n8581) );
  AND U16687 ( .A(n8583), .B(n8584), .Z(n8567) );
  NAND U16688 ( .A(n8585), .B(n8586), .Z(n8584) );
  NANDN U16689 ( .A(n8587), .B(n8588), .Z(n8586) );
  NANDN U16690 ( .A(n8588), .B(n8587), .Z(n8583) );
  XOR U16691 ( .A(n8580), .B(n8589), .Z(N64624) );
  XNOR U16692 ( .A(n8578), .B(n8582), .Z(n8589) );
  XOR U16693 ( .A(n8575), .B(n8590), .Z(n8582) );
  XNOR U16694 ( .A(n8572), .B(n8574), .Z(n8590) );
  AND U16695 ( .A(n8591), .B(n8592), .Z(n8574) );
  NANDN U16696 ( .A(n8593), .B(n8594), .Z(n8592) );
  OR U16697 ( .A(n8595), .B(n8596), .Z(n8594) );
  IV U16698 ( .A(n8597), .Z(n8596) );
  NANDN U16699 ( .A(n8597), .B(n8595), .Z(n8591) );
  AND U16700 ( .A(n8598), .B(n8599), .Z(n8572) );
  NAND U16701 ( .A(n8600), .B(n8601), .Z(n8599) );
  NANDN U16702 ( .A(n8602), .B(n8603), .Z(n8601) );
  NANDN U16703 ( .A(n8603), .B(n8602), .Z(n8598) );
  IV U16704 ( .A(n8604), .Z(n8603) );
  NAND U16705 ( .A(n8605), .B(n8606), .Z(n8575) );
  NANDN U16706 ( .A(n8607), .B(n8608), .Z(n8606) );
  NANDN U16707 ( .A(n8609), .B(n8610), .Z(n8608) );
  NANDN U16708 ( .A(n8610), .B(n8609), .Z(n8605) );
  IV U16709 ( .A(n8611), .Z(n8609) );
  AND U16710 ( .A(n8612), .B(n8613), .Z(n8578) );
  NAND U16711 ( .A(n8614), .B(n8615), .Z(n8613) );
  NANDN U16712 ( .A(n8616), .B(n8617), .Z(n8615) );
  NANDN U16713 ( .A(n8617), .B(n8616), .Z(n8612) );
  XOR U16714 ( .A(n8588), .B(n8618), .Z(n8580) );
  XNOR U16715 ( .A(n8585), .B(n8587), .Z(n8618) );
  AND U16716 ( .A(n8619), .B(n8620), .Z(n8587) );
  NANDN U16717 ( .A(n8621), .B(n8622), .Z(n8620) );
  OR U16718 ( .A(n8623), .B(n8624), .Z(n8622) );
  IV U16719 ( .A(n8625), .Z(n8624) );
  NANDN U16720 ( .A(n8625), .B(n8623), .Z(n8619) );
  AND U16721 ( .A(n8626), .B(n8627), .Z(n8585) );
  NAND U16722 ( .A(n8628), .B(n8629), .Z(n8627) );
  NANDN U16723 ( .A(n8630), .B(n8631), .Z(n8629) );
  NANDN U16724 ( .A(n8631), .B(n8630), .Z(n8626) );
  IV U16725 ( .A(n8632), .Z(n8631) );
  NAND U16726 ( .A(n8633), .B(n8634), .Z(n8588) );
  NANDN U16727 ( .A(n8635), .B(n8636), .Z(n8634) );
  NANDN U16728 ( .A(n8637), .B(n8638), .Z(n8636) );
  NANDN U16729 ( .A(n8638), .B(n8637), .Z(n8633) );
  IV U16730 ( .A(n8639), .Z(n8637) );
  XOR U16731 ( .A(n8614), .B(n8640), .Z(N64623) );
  XNOR U16732 ( .A(n8617), .B(n8616), .Z(n8640) );
  XNOR U16733 ( .A(n8628), .B(n8641), .Z(n8616) );
  XNOR U16734 ( .A(n8632), .B(n8630), .Z(n8641) );
  XOR U16735 ( .A(n8638), .B(n8642), .Z(n8630) );
  XNOR U16736 ( .A(n8635), .B(n8639), .Z(n8642) );
  AND U16737 ( .A(n8643), .B(n8644), .Z(n8639) );
  NAND U16738 ( .A(n8645), .B(n8646), .Z(n8644) );
  NAND U16739 ( .A(n8647), .B(n8648), .Z(n8643) );
  AND U16740 ( .A(n8649), .B(n8650), .Z(n8635) );
  NAND U16741 ( .A(n8651), .B(n8652), .Z(n8650) );
  NAND U16742 ( .A(n8653), .B(n8654), .Z(n8649) );
  NANDN U16743 ( .A(n8655), .B(n8656), .Z(n8638) );
  ANDN U16744 ( .B(n8657), .A(n8658), .Z(n8632) );
  XNOR U16745 ( .A(n8623), .B(n8659), .Z(n8628) );
  XNOR U16746 ( .A(n8621), .B(n8625), .Z(n8659) );
  AND U16747 ( .A(n8660), .B(n8661), .Z(n8625) );
  NAND U16748 ( .A(n8662), .B(n8663), .Z(n8661) );
  NAND U16749 ( .A(n8664), .B(n8665), .Z(n8660) );
  AND U16750 ( .A(n8666), .B(n8667), .Z(n8621) );
  NAND U16751 ( .A(n8668), .B(n8669), .Z(n8667) );
  NAND U16752 ( .A(n8670), .B(n8671), .Z(n8666) );
  AND U16753 ( .A(n8672), .B(n8673), .Z(n8623) );
  NAND U16754 ( .A(n8674), .B(n8675), .Z(n8617) );
  XNOR U16755 ( .A(n8600), .B(n8676), .Z(n8614) );
  XNOR U16756 ( .A(n8604), .B(n8602), .Z(n8676) );
  XOR U16757 ( .A(n8610), .B(n8677), .Z(n8602) );
  XNOR U16758 ( .A(n8607), .B(n8611), .Z(n8677) );
  AND U16759 ( .A(n8678), .B(n8679), .Z(n8611) );
  NAND U16760 ( .A(n8680), .B(n8681), .Z(n8679) );
  NAND U16761 ( .A(n8682), .B(n8683), .Z(n8678) );
  AND U16762 ( .A(n8684), .B(n8685), .Z(n8607) );
  NAND U16763 ( .A(n8686), .B(n8687), .Z(n8685) );
  NAND U16764 ( .A(n8688), .B(n8689), .Z(n8684) );
  NANDN U16765 ( .A(n8690), .B(n8691), .Z(n8610) );
  ANDN U16766 ( .B(n8692), .A(n8693), .Z(n8604) );
  XNOR U16767 ( .A(n8595), .B(n8694), .Z(n8600) );
  XNOR U16768 ( .A(n8593), .B(n8597), .Z(n8694) );
  AND U16769 ( .A(n8695), .B(n8696), .Z(n8597) );
  NAND U16770 ( .A(n8697), .B(n8698), .Z(n8696) );
  NAND U16771 ( .A(n8699), .B(n8700), .Z(n8695) );
  AND U16772 ( .A(n8701), .B(n8702), .Z(n8593) );
  NAND U16773 ( .A(n8703), .B(n8704), .Z(n8702) );
  NAND U16774 ( .A(n8705), .B(n8706), .Z(n8701) );
  AND U16775 ( .A(n8707), .B(n8708), .Z(n8595) );
  XOR U16776 ( .A(n8675), .B(n8674), .Z(N64622) );
  XNOR U16777 ( .A(n8692), .B(n8693), .Z(n8674) );
  XNOR U16778 ( .A(n8707), .B(n8708), .Z(n8693) );
  XOR U16779 ( .A(n8704), .B(n8703), .Z(n8708) );
  XOR U16780 ( .A(y[7452]), .B(x[7452]), .Z(n8703) );
  XOR U16781 ( .A(n8706), .B(n8705), .Z(n8704) );
  XOR U16782 ( .A(y[7454]), .B(x[7454]), .Z(n8705) );
  XOR U16783 ( .A(y[7453]), .B(x[7453]), .Z(n8706) );
  XOR U16784 ( .A(n8698), .B(n8697), .Z(n8707) );
  XOR U16785 ( .A(n8700), .B(n8699), .Z(n8697) );
  XOR U16786 ( .A(y[7451]), .B(x[7451]), .Z(n8699) );
  XOR U16787 ( .A(y[7450]), .B(x[7450]), .Z(n8700) );
  XOR U16788 ( .A(y[7449]), .B(x[7449]), .Z(n8698) );
  XNOR U16789 ( .A(n8691), .B(n8690), .Z(n8692) );
  XNOR U16790 ( .A(n8687), .B(n8686), .Z(n8690) );
  XOR U16791 ( .A(n8689), .B(n8688), .Z(n8686) );
  XOR U16792 ( .A(y[7448]), .B(x[7448]), .Z(n8688) );
  XOR U16793 ( .A(y[7447]), .B(x[7447]), .Z(n8689) );
  XOR U16794 ( .A(y[7446]), .B(x[7446]), .Z(n8687) );
  XOR U16795 ( .A(n8681), .B(n8680), .Z(n8691) );
  XOR U16796 ( .A(n8683), .B(n8682), .Z(n8680) );
  XOR U16797 ( .A(y[7445]), .B(x[7445]), .Z(n8682) );
  XOR U16798 ( .A(y[7444]), .B(x[7444]), .Z(n8683) );
  XOR U16799 ( .A(y[7443]), .B(x[7443]), .Z(n8681) );
  XNOR U16800 ( .A(n8657), .B(n8658), .Z(n8675) );
  XNOR U16801 ( .A(n8672), .B(n8673), .Z(n8658) );
  XOR U16802 ( .A(n8669), .B(n8668), .Z(n8673) );
  XOR U16803 ( .A(y[7440]), .B(x[7440]), .Z(n8668) );
  XOR U16804 ( .A(n8671), .B(n8670), .Z(n8669) );
  XOR U16805 ( .A(y[7442]), .B(x[7442]), .Z(n8670) );
  XOR U16806 ( .A(y[7441]), .B(x[7441]), .Z(n8671) );
  XOR U16807 ( .A(n8663), .B(n8662), .Z(n8672) );
  XOR U16808 ( .A(n8665), .B(n8664), .Z(n8662) );
  XOR U16809 ( .A(y[7439]), .B(x[7439]), .Z(n8664) );
  XOR U16810 ( .A(y[7438]), .B(x[7438]), .Z(n8665) );
  XOR U16811 ( .A(y[7437]), .B(x[7437]), .Z(n8663) );
  XNOR U16812 ( .A(n8656), .B(n8655), .Z(n8657) );
  XNOR U16813 ( .A(n8652), .B(n8651), .Z(n8655) );
  XOR U16814 ( .A(n8654), .B(n8653), .Z(n8651) );
  XOR U16815 ( .A(y[7436]), .B(x[7436]), .Z(n8653) );
  XOR U16816 ( .A(y[7435]), .B(x[7435]), .Z(n8654) );
  XOR U16817 ( .A(y[7434]), .B(x[7434]), .Z(n8652) );
  XOR U16818 ( .A(n8646), .B(n8645), .Z(n8656) );
  XOR U16819 ( .A(n8648), .B(n8647), .Z(n8645) );
  XOR U16820 ( .A(y[7433]), .B(x[7433]), .Z(n8647) );
  XOR U16821 ( .A(y[7432]), .B(x[7432]), .Z(n8648) );
  XOR U16822 ( .A(y[7431]), .B(x[7431]), .Z(n8646) );
  NAND U16823 ( .A(n8709), .B(n8710), .Z(N64613) );
  NAND U16824 ( .A(n8711), .B(n8712), .Z(n8710) );
  NANDN U16825 ( .A(n8713), .B(n8714), .Z(n8712) );
  NANDN U16826 ( .A(n8714), .B(n8713), .Z(n8709) );
  XOR U16827 ( .A(n8713), .B(n8715), .Z(N64612) );
  XNOR U16828 ( .A(n8711), .B(n8714), .Z(n8715) );
  NAND U16829 ( .A(n8716), .B(n8717), .Z(n8714) );
  NAND U16830 ( .A(n8718), .B(n8719), .Z(n8717) );
  NANDN U16831 ( .A(n8720), .B(n8721), .Z(n8719) );
  NANDN U16832 ( .A(n8721), .B(n8720), .Z(n8716) );
  AND U16833 ( .A(n8722), .B(n8723), .Z(n8711) );
  NAND U16834 ( .A(n8724), .B(n8725), .Z(n8723) );
  NANDN U16835 ( .A(n8726), .B(n8727), .Z(n8725) );
  NANDN U16836 ( .A(n8727), .B(n8726), .Z(n8722) );
  IV U16837 ( .A(n8728), .Z(n8727) );
  AND U16838 ( .A(n8729), .B(n8730), .Z(n8713) );
  NAND U16839 ( .A(n8731), .B(n8732), .Z(n8730) );
  NANDN U16840 ( .A(n8733), .B(n8734), .Z(n8732) );
  NANDN U16841 ( .A(n8734), .B(n8733), .Z(n8729) );
  XOR U16842 ( .A(n8726), .B(n8735), .Z(N64611) );
  XNOR U16843 ( .A(n8724), .B(n8728), .Z(n8735) );
  XOR U16844 ( .A(n8721), .B(n8736), .Z(n8728) );
  XNOR U16845 ( .A(n8718), .B(n8720), .Z(n8736) );
  AND U16846 ( .A(n8737), .B(n8738), .Z(n8720) );
  NANDN U16847 ( .A(n8739), .B(n8740), .Z(n8738) );
  OR U16848 ( .A(n8741), .B(n8742), .Z(n8740) );
  IV U16849 ( .A(n8743), .Z(n8742) );
  NANDN U16850 ( .A(n8743), .B(n8741), .Z(n8737) );
  AND U16851 ( .A(n8744), .B(n8745), .Z(n8718) );
  NAND U16852 ( .A(n8746), .B(n8747), .Z(n8745) );
  NANDN U16853 ( .A(n8748), .B(n8749), .Z(n8747) );
  NANDN U16854 ( .A(n8749), .B(n8748), .Z(n8744) );
  IV U16855 ( .A(n8750), .Z(n8749) );
  NAND U16856 ( .A(n8751), .B(n8752), .Z(n8721) );
  NANDN U16857 ( .A(n8753), .B(n8754), .Z(n8752) );
  NANDN U16858 ( .A(n8755), .B(n8756), .Z(n8754) );
  NANDN U16859 ( .A(n8756), .B(n8755), .Z(n8751) );
  IV U16860 ( .A(n8757), .Z(n8755) );
  AND U16861 ( .A(n8758), .B(n8759), .Z(n8724) );
  NAND U16862 ( .A(n8760), .B(n8761), .Z(n8759) );
  NANDN U16863 ( .A(n8762), .B(n8763), .Z(n8761) );
  NANDN U16864 ( .A(n8763), .B(n8762), .Z(n8758) );
  XOR U16865 ( .A(n8734), .B(n8764), .Z(n8726) );
  XNOR U16866 ( .A(n8731), .B(n8733), .Z(n8764) );
  AND U16867 ( .A(n8765), .B(n8766), .Z(n8733) );
  NANDN U16868 ( .A(n8767), .B(n8768), .Z(n8766) );
  OR U16869 ( .A(n8769), .B(n8770), .Z(n8768) );
  IV U16870 ( .A(n8771), .Z(n8770) );
  NANDN U16871 ( .A(n8771), .B(n8769), .Z(n8765) );
  AND U16872 ( .A(n8772), .B(n8773), .Z(n8731) );
  NAND U16873 ( .A(n8774), .B(n8775), .Z(n8773) );
  NANDN U16874 ( .A(n8776), .B(n8777), .Z(n8775) );
  NANDN U16875 ( .A(n8777), .B(n8776), .Z(n8772) );
  IV U16876 ( .A(n8778), .Z(n8777) );
  NAND U16877 ( .A(n8779), .B(n8780), .Z(n8734) );
  NANDN U16878 ( .A(n8781), .B(n8782), .Z(n8780) );
  NANDN U16879 ( .A(n8783), .B(n8784), .Z(n8782) );
  NANDN U16880 ( .A(n8784), .B(n8783), .Z(n8779) );
  IV U16881 ( .A(n8785), .Z(n8783) );
  XOR U16882 ( .A(n8760), .B(n8786), .Z(N64610) );
  XNOR U16883 ( .A(n8763), .B(n8762), .Z(n8786) );
  XNOR U16884 ( .A(n8774), .B(n8787), .Z(n8762) );
  XNOR U16885 ( .A(n8778), .B(n8776), .Z(n8787) );
  XOR U16886 ( .A(n8784), .B(n8788), .Z(n8776) );
  XNOR U16887 ( .A(n8781), .B(n8785), .Z(n8788) );
  AND U16888 ( .A(n8789), .B(n8790), .Z(n8785) );
  NAND U16889 ( .A(n8791), .B(n8792), .Z(n8790) );
  NAND U16890 ( .A(n8793), .B(n8794), .Z(n8789) );
  AND U16891 ( .A(n8795), .B(n8796), .Z(n8781) );
  NAND U16892 ( .A(n8797), .B(n8798), .Z(n8796) );
  NAND U16893 ( .A(n8799), .B(n8800), .Z(n8795) );
  NANDN U16894 ( .A(n8801), .B(n8802), .Z(n8784) );
  ANDN U16895 ( .B(n8803), .A(n8804), .Z(n8778) );
  XNOR U16896 ( .A(n8769), .B(n8805), .Z(n8774) );
  XNOR U16897 ( .A(n8767), .B(n8771), .Z(n8805) );
  AND U16898 ( .A(n8806), .B(n8807), .Z(n8771) );
  NAND U16899 ( .A(n8808), .B(n8809), .Z(n8807) );
  NAND U16900 ( .A(n8810), .B(n8811), .Z(n8806) );
  AND U16901 ( .A(n8812), .B(n8813), .Z(n8767) );
  NAND U16902 ( .A(n8814), .B(n8815), .Z(n8813) );
  NAND U16903 ( .A(n8816), .B(n8817), .Z(n8812) );
  AND U16904 ( .A(n8818), .B(n8819), .Z(n8769) );
  NAND U16905 ( .A(n8820), .B(n8821), .Z(n8763) );
  XNOR U16906 ( .A(n8746), .B(n8822), .Z(n8760) );
  XNOR U16907 ( .A(n8750), .B(n8748), .Z(n8822) );
  XOR U16908 ( .A(n8756), .B(n8823), .Z(n8748) );
  XNOR U16909 ( .A(n8753), .B(n8757), .Z(n8823) );
  AND U16910 ( .A(n8824), .B(n8825), .Z(n8757) );
  NAND U16911 ( .A(n8826), .B(n8827), .Z(n8825) );
  NAND U16912 ( .A(n8828), .B(n8829), .Z(n8824) );
  AND U16913 ( .A(n8830), .B(n8831), .Z(n8753) );
  NAND U16914 ( .A(n8832), .B(n8833), .Z(n8831) );
  NAND U16915 ( .A(n8834), .B(n8835), .Z(n8830) );
  NANDN U16916 ( .A(n8836), .B(n8837), .Z(n8756) );
  ANDN U16917 ( .B(n8838), .A(n8839), .Z(n8750) );
  XNOR U16918 ( .A(n8741), .B(n8840), .Z(n8746) );
  XNOR U16919 ( .A(n8739), .B(n8743), .Z(n8840) );
  AND U16920 ( .A(n8841), .B(n8842), .Z(n8743) );
  NAND U16921 ( .A(n8843), .B(n8844), .Z(n8842) );
  NAND U16922 ( .A(n8845), .B(n8846), .Z(n8841) );
  AND U16923 ( .A(n8847), .B(n8848), .Z(n8739) );
  NAND U16924 ( .A(n8849), .B(n8850), .Z(n8848) );
  NAND U16925 ( .A(n8851), .B(n8852), .Z(n8847) );
  AND U16926 ( .A(n8853), .B(n8854), .Z(n8741) );
  XOR U16927 ( .A(n8821), .B(n8820), .Z(N64609) );
  XNOR U16928 ( .A(n8838), .B(n8839), .Z(n8820) );
  XNOR U16929 ( .A(n8853), .B(n8854), .Z(n8839) );
  XOR U16930 ( .A(n8850), .B(n8849), .Z(n8854) );
  XOR U16931 ( .A(y[7428]), .B(x[7428]), .Z(n8849) );
  XOR U16932 ( .A(n8852), .B(n8851), .Z(n8850) );
  XOR U16933 ( .A(y[7430]), .B(x[7430]), .Z(n8851) );
  XOR U16934 ( .A(y[7429]), .B(x[7429]), .Z(n8852) );
  XOR U16935 ( .A(n8844), .B(n8843), .Z(n8853) );
  XOR U16936 ( .A(n8846), .B(n8845), .Z(n8843) );
  XOR U16937 ( .A(y[7427]), .B(x[7427]), .Z(n8845) );
  XOR U16938 ( .A(y[7426]), .B(x[7426]), .Z(n8846) );
  XOR U16939 ( .A(y[7425]), .B(x[7425]), .Z(n8844) );
  XNOR U16940 ( .A(n8837), .B(n8836), .Z(n8838) );
  XNOR U16941 ( .A(n8833), .B(n8832), .Z(n8836) );
  XOR U16942 ( .A(n8835), .B(n8834), .Z(n8832) );
  XOR U16943 ( .A(y[7424]), .B(x[7424]), .Z(n8834) );
  XOR U16944 ( .A(y[7423]), .B(x[7423]), .Z(n8835) );
  XOR U16945 ( .A(y[7422]), .B(x[7422]), .Z(n8833) );
  XOR U16946 ( .A(n8827), .B(n8826), .Z(n8837) );
  XOR U16947 ( .A(n8829), .B(n8828), .Z(n8826) );
  XOR U16948 ( .A(y[7421]), .B(x[7421]), .Z(n8828) );
  XOR U16949 ( .A(y[7420]), .B(x[7420]), .Z(n8829) );
  XOR U16950 ( .A(y[7419]), .B(x[7419]), .Z(n8827) );
  XNOR U16951 ( .A(n8803), .B(n8804), .Z(n8821) );
  XNOR U16952 ( .A(n8818), .B(n8819), .Z(n8804) );
  XOR U16953 ( .A(n8815), .B(n8814), .Z(n8819) );
  XOR U16954 ( .A(y[7416]), .B(x[7416]), .Z(n8814) );
  XOR U16955 ( .A(n8817), .B(n8816), .Z(n8815) );
  XOR U16956 ( .A(y[7418]), .B(x[7418]), .Z(n8816) );
  XOR U16957 ( .A(y[7417]), .B(x[7417]), .Z(n8817) );
  XOR U16958 ( .A(n8809), .B(n8808), .Z(n8818) );
  XOR U16959 ( .A(n8811), .B(n8810), .Z(n8808) );
  XOR U16960 ( .A(y[7415]), .B(x[7415]), .Z(n8810) );
  XOR U16961 ( .A(y[7414]), .B(x[7414]), .Z(n8811) );
  XOR U16962 ( .A(y[7413]), .B(x[7413]), .Z(n8809) );
  XNOR U16963 ( .A(n8802), .B(n8801), .Z(n8803) );
  XNOR U16964 ( .A(n8798), .B(n8797), .Z(n8801) );
  XOR U16965 ( .A(n8800), .B(n8799), .Z(n8797) );
  XOR U16966 ( .A(y[7412]), .B(x[7412]), .Z(n8799) );
  XOR U16967 ( .A(y[7411]), .B(x[7411]), .Z(n8800) );
  XOR U16968 ( .A(y[7410]), .B(x[7410]), .Z(n8798) );
  XOR U16969 ( .A(n8792), .B(n8791), .Z(n8802) );
  XOR U16970 ( .A(n8794), .B(n8793), .Z(n8791) );
  XOR U16971 ( .A(y[7409]), .B(x[7409]), .Z(n8793) );
  XOR U16972 ( .A(y[7408]), .B(x[7408]), .Z(n8794) );
  XOR U16973 ( .A(y[7407]), .B(x[7407]), .Z(n8792) );
  NAND U16974 ( .A(n8855), .B(n8856), .Z(N64600) );
  NAND U16975 ( .A(n8857), .B(n8858), .Z(n8856) );
  NANDN U16976 ( .A(n8859), .B(n8860), .Z(n8858) );
  NANDN U16977 ( .A(n8860), .B(n8859), .Z(n8855) );
  XOR U16978 ( .A(n8859), .B(n8861), .Z(N64599) );
  XNOR U16979 ( .A(n8857), .B(n8860), .Z(n8861) );
  NAND U16980 ( .A(n8862), .B(n8863), .Z(n8860) );
  NAND U16981 ( .A(n8864), .B(n8865), .Z(n8863) );
  NANDN U16982 ( .A(n8866), .B(n8867), .Z(n8865) );
  NANDN U16983 ( .A(n8867), .B(n8866), .Z(n8862) );
  AND U16984 ( .A(n8868), .B(n8869), .Z(n8857) );
  NAND U16985 ( .A(n8870), .B(n8871), .Z(n8869) );
  NANDN U16986 ( .A(n8872), .B(n8873), .Z(n8871) );
  NANDN U16987 ( .A(n8873), .B(n8872), .Z(n8868) );
  IV U16988 ( .A(n8874), .Z(n8873) );
  AND U16989 ( .A(n8875), .B(n8876), .Z(n8859) );
  NAND U16990 ( .A(n8877), .B(n8878), .Z(n8876) );
  NANDN U16991 ( .A(n8879), .B(n8880), .Z(n8878) );
  NANDN U16992 ( .A(n8880), .B(n8879), .Z(n8875) );
  XOR U16993 ( .A(n8872), .B(n8881), .Z(N64598) );
  XNOR U16994 ( .A(n8870), .B(n8874), .Z(n8881) );
  XOR U16995 ( .A(n8867), .B(n8882), .Z(n8874) );
  XNOR U16996 ( .A(n8864), .B(n8866), .Z(n8882) );
  AND U16997 ( .A(n8883), .B(n8884), .Z(n8866) );
  NANDN U16998 ( .A(n8885), .B(n8886), .Z(n8884) );
  OR U16999 ( .A(n8887), .B(n8888), .Z(n8886) );
  IV U17000 ( .A(n8889), .Z(n8888) );
  NANDN U17001 ( .A(n8889), .B(n8887), .Z(n8883) );
  AND U17002 ( .A(n8890), .B(n8891), .Z(n8864) );
  NAND U17003 ( .A(n8892), .B(n8893), .Z(n8891) );
  NANDN U17004 ( .A(n8894), .B(n8895), .Z(n8893) );
  NANDN U17005 ( .A(n8895), .B(n8894), .Z(n8890) );
  IV U17006 ( .A(n8896), .Z(n8895) );
  NAND U17007 ( .A(n8897), .B(n8898), .Z(n8867) );
  NANDN U17008 ( .A(n8899), .B(n8900), .Z(n8898) );
  NANDN U17009 ( .A(n8901), .B(n8902), .Z(n8900) );
  NANDN U17010 ( .A(n8902), .B(n8901), .Z(n8897) );
  IV U17011 ( .A(n8903), .Z(n8901) );
  AND U17012 ( .A(n8904), .B(n8905), .Z(n8870) );
  NAND U17013 ( .A(n8906), .B(n8907), .Z(n8905) );
  NANDN U17014 ( .A(n8908), .B(n8909), .Z(n8907) );
  NANDN U17015 ( .A(n8909), .B(n8908), .Z(n8904) );
  XOR U17016 ( .A(n8880), .B(n8910), .Z(n8872) );
  XNOR U17017 ( .A(n8877), .B(n8879), .Z(n8910) );
  AND U17018 ( .A(n8911), .B(n8912), .Z(n8879) );
  NANDN U17019 ( .A(n8913), .B(n8914), .Z(n8912) );
  OR U17020 ( .A(n8915), .B(n8916), .Z(n8914) );
  IV U17021 ( .A(n8917), .Z(n8916) );
  NANDN U17022 ( .A(n8917), .B(n8915), .Z(n8911) );
  AND U17023 ( .A(n8918), .B(n8919), .Z(n8877) );
  NAND U17024 ( .A(n8920), .B(n8921), .Z(n8919) );
  NANDN U17025 ( .A(n8922), .B(n8923), .Z(n8921) );
  NANDN U17026 ( .A(n8923), .B(n8922), .Z(n8918) );
  IV U17027 ( .A(n8924), .Z(n8923) );
  NAND U17028 ( .A(n8925), .B(n8926), .Z(n8880) );
  NANDN U17029 ( .A(n8927), .B(n8928), .Z(n8926) );
  NANDN U17030 ( .A(n8929), .B(n8930), .Z(n8928) );
  NANDN U17031 ( .A(n8930), .B(n8929), .Z(n8925) );
  IV U17032 ( .A(n8931), .Z(n8929) );
  XOR U17033 ( .A(n8906), .B(n8932), .Z(N64597) );
  XNOR U17034 ( .A(n8909), .B(n8908), .Z(n8932) );
  XNOR U17035 ( .A(n8920), .B(n8933), .Z(n8908) );
  XNOR U17036 ( .A(n8924), .B(n8922), .Z(n8933) );
  XOR U17037 ( .A(n8930), .B(n8934), .Z(n8922) );
  XNOR U17038 ( .A(n8927), .B(n8931), .Z(n8934) );
  AND U17039 ( .A(n8935), .B(n8936), .Z(n8931) );
  NAND U17040 ( .A(n8937), .B(n8938), .Z(n8936) );
  NAND U17041 ( .A(n8939), .B(n8940), .Z(n8935) );
  AND U17042 ( .A(n8941), .B(n8942), .Z(n8927) );
  NAND U17043 ( .A(n8943), .B(n8944), .Z(n8942) );
  NAND U17044 ( .A(n8945), .B(n8946), .Z(n8941) );
  NANDN U17045 ( .A(n8947), .B(n8948), .Z(n8930) );
  ANDN U17046 ( .B(n8949), .A(n8950), .Z(n8924) );
  XNOR U17047 ( .A(n8915), .B(n8951), .Z(n8920) );
  XNOR U17048 ( .A(n8913), .B(n8917), .Z(n8951) );
  AND U17049 ( .A(n8952), .B(n8953), .Z(n8917) );
  NAND U17050 ( .A(n8954), .B(n8955), .Z(n8953) );
  NAND U17051 ( .A(n8956), .B(n8957), .Z(n8952) );
  AND U17052 ( .A(n8958), .B(n8959), .Z(n8913) );
  NAND U17053 ( .A(n8960), .B(n8961), .Z(n8959) );
  NAND U17054 ( .A(n8962), .B(n8963), .Z(n8958) );
  AND U17055 ( .A(n8964), .B(n8965), .Z(n8915) );
  NAND U17056 ( .A(n8966), .B(n8967), .Z(n8909) );
  XNOR U17057 ( .A(n8892), .B(n8968), .Z(n8906) );
  XNOR U17058 ( .A(n8896), .B(n8894), .Z(n8968) );
  XOR U17059 ( .A(n8902), .B(n8969), .Z(n8894) );
  XNOR U17060 ( .A(n8899), .B(n8903), .Z(n8969) );
  AND U17061 ( .A(n8970), .B(n8971), .Z(n8903) );
  NAND U17062 ( .A(n8972), .B(n8973), .Z(n8971) );
  NAND U17063 ( .A(n8974), .B(n8975), .Z(n8970) );
  AND U17064 ( .A(n8976), .B(n8977), .Z(n8899) );
  NAND U17065 ( .A(n8978), .B(n8979), .Z(n8977) );
  NAND U17066 ( .A(n8980), .B(n8981), .Z(n8976) );
  NANDN U17067 ( .A(n8982), .B(n8983), .Z(n8902) );
  ANDN U17068 ( .B(n8984), .A(n8985), .Z(n8896) );
  XNOR U17069 ( .A(n8887), .B(n8986), .Z(n8892) );
  XNOR U17070 ( .A(n8885), .B(n8889), .Z(n8986) );
  AND U17071 ( .A(n8987), .B(n8988), .Z(n8889) );
  NAND U17072 ( .A(n8989), .B(n8990), .Z(n8988) );
  NAND U17073 ( .A(n8991), .B(n8992), .Z(n8987) );
  AND U17074 ( .A(n8993), .B(n8994), .Z(n8885) );
  NAND U17075 ( .A(n8995), .B(n8996), .Z(n8994) );
  NAND U17076 ( .A(n8997), .B(n8998), .Z(n8993) );
  AND U17077 ( .A(n8999), .B(n9000), .Z(n8887) );
  XOR U17078 ( .A(n8967), .B(n8966), .Z(N64596) );
  XNOR U17079 ( .A(n8984), .B(n8985), .Z(n8966) );
  XNOR U17080 ( .A(n8999), .B(n9000), .Z(n8985) );
  XOR U17081 ( .A(n8996), .B(n8995), .Z(n9000) );
  XOR U17082 ( .A(y[7404]), .B(x[7404]), .Z(n8995) );
  XOR U17083 ( .A(n8998), .B(n8997), .Z(n8996) );
  XOR U17084 ( .A(y[7406]), .B(x[7406]), .Z(n8997) );
  XOR U17085 ( .A(y[7405]), .B(x[7405]), .Z(n8998) );
  XOR U17086 ( .A(n8990), .B(n8989), .Z(n8999) );
  XOR U17087 ( .A(n8992), .B(n8991), .Z(n8989) );
  XOR U17088 ( .A(y[7403]), .B(x[7403]), .Z(n8991) );
  XOR U17089 ( .A(y[7402]), .B(x[7402]), .Z(n8992) );
  XOR U17090 ( .A(y[7401]), .B(x[7401]), .Z(n8990) );
  XNOR U17091 ( .A(n8983), .B(n8982), .Z(n8984) );
  XNOR U17092 ( .A(n8979), .B(n8978), .Z(n8982) );
  XOR U17093 ( .A(n8981), .B(n8980), .Z(n8978) );
  XOR U17094 ( .A(y[7400]), .B(x[7400]), .Z(n8980) );
  XOR U17095 ( .A(y[7399]), .B(x[7399]), .Z(n8981) );
  XOR U17096 ( .A(y[7398]), .B(x[7398]), .Z(n8979) );
  XOR U17097 ( .A(n8973), .B(n8972), .Z(n8983) );
  XOR U17098 ( .A(n8975), .B(n8974), .Z(n8972) );
  XOR U17099 ( .A(y[7397]), .B(x[7397]), .Z(n8974) );
  XOR U17100 ( .A(y[7396]), .B(x[7396]), .Z(n8975) );
  XOR U17101 ( .A(y[7395]), .B(x[7395]), .Z(n8973) );
  XNOR U17102 ( .A(n8949), .B(n8950), .Z(n8967) );
  XNOR U17103 ( .A(n8964), .B(n8965), .Z(n8950) );
  XOR U17104 ( .A(n8961), .B(n8960), .Z(n8965) );
  XOR U17105 ( .A(y[7392]), .B(x[7392]), .Z(n8960) );
  XOR U17106 ( .A(n8963), .B(n8962), .Z(n8961) );
  XOR U17107 ( .A(y[7394]), .B(x[7394]), .Z(n8962) );
  XOR U17108 ( .A(y[7393]), .B(x[7393]), .Z(n8963) );
  XOR U17109 ( .A(n8955), .B(n8954), .Z(n8964) );
  XOR U17110 ( .A(n8957), .B(n8956), .Z(n8954) );
  XOR U17111 ( .A(y[7391]), .B(x[7391]), .Z(n8956) );
  XOR U17112 ( .A(y[7390]), .B(x[7390]), .Z(n8957) );
  XOR U17113 ( .A(y[7389]), .B(x[7389]), .Z(n8955) );
  XNOR U17114 ( .A(n8948), .B(n8947), .Z(n8949) );
  XNOR U17115 ( .A(n8944), .B(n8943), .Z(n8947) );
  XOR U17116 ( .A(n8946), .B(n8945), .Z(n8943) );
  XOR U17117 ( .A(y[7388]), .B(x[7388]), .Z(n8945) );
  XOR U17118 ( .A(y[7387]), .B(x[7387]), .Z(n8946) );
  XOR U17119 ( .A(y[7386]), .B(x[7386]), .Z(n8944) );
  XOR U17120 ( .A(n8938), .B(n8937), .Z(n8948) );
  XOR U17121 ( .A(n8940), .B(n8939), .Z(n8937) );
  XOR U17122 ( .A(y[7385]), .B(x[7385]), .Z(n8939) );
  XOR U17123 ( .A(y[7384]), .B(x[7384]), .Z(n8940) );
  XOR U17124 ( .A(y[7383]), .B(x[7383]), .Z(n8938) );
  NAND U17125 ( .A(n9001), .B(n9002), .Z(N64587) );
  NAND U17126 ( .A(n9003), .B(n9004), .Z(n9002) );
  NANDN U17127 ( .A(n9005), .B(n9006), .Z(n9004) );
  NANDN U17128 ( .A(n9006), .B(n9005), .Z(n9001) );
  XOR U17129 ( .A(n9005), .B(n9007), .Z(N64586) );
  XNOR U17130 ( .A(n9003), .B(n9006), .Z(n9007) );
  NAND U17131 ( .A(n9008), .B(n9009), .Z(n9006) );
  NAND U17132 ( .A(n9010), .B(n9011), .Z(n9009) );
  NANDN U17133 ( .A(n9012), .B(n9013), .Z(n9011) );
  NANDN U17134 ( .A(n9013), .B(n9012), .Z(n9008) );
  AND U17135 ( .A(n9014), .B(n9015), .Z(n9003) );
  NAND U17136 ( .A(n9016), .B(n9017), .Z(n9015) );
  NANDN U17137 ( .A(n9018), .B(n9019), .Z(n9017) );
  NANDN U17138 ( .A(n9019), .B(n9018), .Z(n9014) );
  IV U17139 ( .A(n9020), .Z(n9019) );
  AND U17140 ( .A(n9021), .B(n9022), .Z(n9005) );
  NAND U17141 ( .A(n9023), .B(n9024), .Z(n9022) );
  NANDN U17142 ( .A(n9025), .B(n9026), .Z(n9024) );
  NANDN U17143 ( .A(n9026), .B(n9025), .Z(n9021) );
  XOR U17144 ( .A(n9018), .B(n9027), .Z(N64585) );
  XNOR U17145 ( .A(n9016), .B(n9020), .Z(n9027) );
  XOR U17146 ( .A(n9013), .B(n9028), .Z(n9020) );
  XNOR U17147 ( .A(n9010), .B(n9012), .Z(n9028) );
  AND U17148 ( .A(n9029), .B(n9030), .Z(n9012) );
  NANDN U17149 ( .A(n9031), .B(n9032), .Z(n9030) );
  OR U17150 ( .A(n9033), .B(n9034), .Z(n9032) );
  IV U17151 ( .A(n9035), .Z(n9034) );
  NANDN U17152 ( .A(n9035), .B(n9033), .Z(n9029) );
  AND U17153 ( .A(n9036), .B(n9037), .Z(n9010) );
  NAND U17154 ( .A(n9038), .B(n9039), .Z(n9037) );
  NANDN U17155 ( .A(n9040), .B(n9041), .Z(n9039) );
  NANDN U17156 ( .A(n9041), .B(n9040), .Z(n9036) );
  IV U17157 ( .A(n9042), .Z(n9041) );
  NAND U17158 ( .A(n9043), .B(n9044), .Z(n9013) );
  NANDN U17159 ( .A(n9045), .B(n9046), .Z(n9044) );
  NANDN U17160 ( .A(n9047), .B(n9048), .Z(n9046) );
  NANDN U17161 ( .A(n9048), .B(n9047), .Z(n9043) );
  IV U17162 ( .A(n9049), .Z(n9047) );
  AND U17163 ( .A(n9050), .B(n9051), .Z(n9016) );
  NAND U17164 ( .A(n9052), .B(n9053), .Z(n9051) );
  NANDN U17165 ( .A(n9054), .B(n9055), .Z(n9053) );
  NANDN U17166 ( .A(n9055), .B(n9054), .Z(n9050) );
  XOR U17167 ( .A(n9026), .B(n9056), .Z(n9018) );
  XNOR U17168 ( .A(n9023), .B(n9025), .Z(n9056) );
  AND U17169 ( .A(n9057), .B(n9058), .Z(n9025) );
  NANDN U17170 ( .A(n9059), .B(n9060), .Z(n9058) );
  OR U17171 ( .A(n9061), .B(n9062), .Z(n9060) );
  IV U17172 ( .A(n9063), .Z(n9062) );
  NANDN U17173 ( .A(n9063), .B(n9061), .Z(n9057) );
  AND U17174 ( .A(n9064), .B(n9065), .Z(n9023) );
  NAND U17175 ( .A(n9066), .B(n9067), .Z(n9065) );
  NANDN U17176 ( .A(n9068), .B(n9069), .Z(n9067) );
  NANDN U17177 ( .A(n9069), .B(n9068), .Z(n9064) );
  IV U17178 ( .A(n9070), .Z(n9069) );
  NAND U17179 ( .A(n9071), .B(n9072), .Z(n9026) );
  NANDN U17180 ( .A(n9073), .B(n9074), .Z(n9072) );
  NANDN U17181 ( .A(n9075), .B(n9076), .Z(n9074) );
  NANDN U17182 ( .A(n9076), .B(n9075), .Z(n9071) );
  IV U17183 ( .A(n9077), .Z(n9075) );
  XOR U17184 ( .A(n9052), .B(n9078), .Z(N64584) );
  XNOR U17185 ( .A(n9055), .B(n9054), .Z(n9078) );
  XNOR U17186 ( .A(n9066), .B(n9079), .Z(n9054) );
  XNOR U17187 ( .A(n9070), .B(n9068), .Z(n9079) );
  XOR U17188 ( .A(n9076), .B(n9080), .Z(n9068) );
  XNOR U17189 ( .A(n9073), .B(n9077), .Z(n9080) );
  AND U17190 ( .A(n9081), .B(n9082), .Z(n9077) );
  NAND U17191 ( .A(n9083), .B(n9084), .Z(n9082) );
  NAND U17192 ( .A(n9085), .B(n9086), .Z(n9081) );
  AND U17193 ( .A(n9087), .B(n9088), .Z(n9073) );
  NAND U17194 ( .A(n9089), .B(n9090), .Z(n9088) );
  NAND U17195 ( .A(n9091), .B(n9092), .Z(n9087) );
  NANDN U17196 ( .A(n9093), .B(n9094), .Z(n9076) );
  ANDN U17197 ( .B(n9095), .A(n9096), .Z(n9070) );
  XNOR U17198 ( .A(n9061), .B(n9097), .Z(n9066) );
  XNOR U17199 ( .A(n9059), .B(n9063), .Z(n9097) );
  AND U17200 ( .A(n9098), .B(n9099), .Z(n9063) );
  NAND U17201 ( .A(n9100), .B(n9101), .Z(n9099) );
  NAND U17202 ( .A(n9102), .B(n9103), .Z(n9098) );
  AND U17203 ( .A(n9104), .B(n9105), .Z(n9059) );
  NAND U17204 ( .A(n9106), .B(n9107), .Z(n9105) );
  NAND U17205 ( .A(n9108), .B(n9109), .Z(n9104) );
  AND U17206 ( .A(n9110), .B(n9111), .Z(n9061) );
  NAND U17207 ( .A(n9112), .B(n9113), .Z(n9055) );
  XNOR U17208 ( .A(n9038), .B(n9114), .Z(n9052) );
  XNOR U17209 ( .A(n9042), .B(n9040), .Z(n9114) );
  XOR U17210 ( .A(n9048), .B(n9115), .Z(n9040) );
  XNOR U17211 ( .A(n9045), .B(n9049), .Z(n9115) );
  AND U17212 ( .A(n9116), .B(n9117), .Z(n9049) );
  NAND U17213 ( .A(n9118), .B(n9119), .Z(n9117) );
  NAND U17214 ( .A(n9120), .B(n9121), .Z(n9116) );
  AND U17215 ( .A(n9122), .B(n9123), .Z(n9045) );
  NAND U17216 ( .A(n9124), .B(n9125), .Z(n9123) );
  NAND U17217 ( .A(n9126), .B(n9127), .Z(n9122) );
  NANDN U17218 ( .A(n9128), .B(n9129), .Z(n9048) );
  ANDN U17219 ( .B(n9130), .A(n9131), .Z(n9042) );
  XNOR U17220 ( .A(n9033), .B(n9132), .Z(n9038) );
  XNOR U17221 ( .A(n9031), .B(n9035), .Z(n9132) );
  AND U17222 ( .A(n9133), .B(n9134), .Z(n9035) );
  NAND U17223 ( .A(n9135), .B(n9136), .Z(n9134) );
  NAND U17224 ( .A(n9137), .B(n9138), .Z(n9133) );
  AND U17225 ( .A(n9139), .B(n9140), .Z(n9031) );
  NAND U17226 ( .A(n9141), .B(n9142), .Z(n9140) );
  NAND U17227 ( .A(n9143), .B(n9144), .Z(n9139) );
  AND U17228 ( .A(n9145), .B(n9146), .Z(n9033) );
  XOR U17229 ( .A(n9113), .B(n9112), .Z(N64583) );
  XNOR U17230 ( .A(n9130), .B(n9131), .Z(n9112) );
  XNOR U17231 ( .A(n9145), .B(n9146), .Z(n9131) );
  XOR U17232 ( .A(n9142), .B(n9141), .Z(n9146) );
  XOR U17233 ( .A(y[7380]), .B(x[7380]), .Z(n9141) );
  XOR U17234 ( .A(n9144), .B(n9143), .Z(n9142) );
  XOR U17235 ( .A(y[7382]), .B(x[7382]), .Z(n9143) );
  XOR U17236 ( .A(y[7381]), .B(x[7381]), .Z(n9144) );
  XOR U17237 ( .A(n9136), .B(n9135), .Z(n9145) );
  XOR U17238 ( .A(n9138), .B(n9137), .Z(n9135) );
  XOR U17239 ( .A(y[7379]), .B(x[7379]), .Z(n9137) );
  XOR U17240 ( .A(y[7378]), .B(x[7378]), .Z(n9138) );
  XOR U17241 ( .A(y[7377]), .B(x[7377]), .Z(n9136) );
  XNOR U17242 ( .A(n9129), .B(n9128), .Z(n9130) );
  XNOR U17243 ( .A(n9125), .B(n9124), .Z(n9128) );
  XOR U17244 ( .A(n9127), .B(n9126), .Z(n9124) );
  XOR U17245 ( .A(y[7376]), .B(x[7376]), .Z(n9126) );
  XOR U17246 ( .A(y[7375]), .B(x[7375]), .Z(n9127) );
  XOR U17247 ( .A(y[7374]), .B(x[7374]), .Z(n9125) );
  XOR U17248 ( .A(n9119), .B(n9118), .Z(n9129) );
  XOR U17249 ( .A(n9121), .B(n9120), .Z(n9118) );
  XOR U17250 ( .A(y[7373]), .B(x[7373]), .Z(n9120) );
  XOR U17251 ( .A(y[7372]), .B(x[7372]), .Z(n9121) );
  XOR U17252 ( .A(y[7371]), .B(x[7371]), .Z(n9119) );
  XNOR U17253 ( .A(n9095), .B(n9096), .Z(n9113) );
  XNOR U17254 ( .A(n9110), .B(n9111), .Z(n9096) );
  XOR U17255 ( .A(n9107), .B(n9106), .Z(n9111) );
  XOR U17256 ( .A(y[7368]), .B(x[7368]), .Z(n9106) );
  XOR U17257 ( .A(n9109), .B(n9108), .Z(n9107) );
  XOR U17258 ( .A(y[7370]), .B(x[7370]), .Z(n9108) );
  XOR U17259 ( .A(y[7369]), .B(x[7369]), .Z(n9109) );
  XOR U17260 ( .A(n9101), .B(n9100), .Z(n9110) );
  XOR U17261 ( .A(n9103), .B(n9102), .Z(n9100) );
  XOR U17262 ( .A(y[7367]), .B(x[7367]), .Z(n9102) );
  XOR U17263 ( .A(y[7366]), .B(x[7366]), .Z(n9103) );
  XOR U17264 ( .A(y[7365]), .B(x[7365]), .Z(n9101) );
  XNOR U17265 ( .A(n9094), .B(n9093), .Z(n9095) );
  XNOR U17266 ( .A(n9090), .B(n9089), .Z(n9093) );
  XOR U17267 ( .A(n9092), .B(n9091), .Z(n9089) );
  XOR U17268 ( .A(y[7364]), .B(x[7364]), .Z(n9091) );
  XOR U17269 ( .A(y[7363]), .B(x[7363]), .Z(n9092) );
  XOR U17270 ( .A(y[7362]), .B(x[7362]), .Z(n9090) );
  XOR U17271 ( .A(n9084), .B(n9083), .Z(n9094) );
  XOR U17272 ( .A(n9086), .B(n9085), .Z(n9083) );
  XOR U17273 ( .A(y[7361]), .B(x[7361]), .Z(n9085) );
  XOR U17274 ( .A(y[7360]), .B(x[7360]), .Z(n9086) );
  XOR U17275 ( .A(y[7359]), .B(x[7359]), .Z(n9084) );
  NAND U17276 ( .A(n9147), .B(n9148), .Z(N64574) );
  NAND U17277 ( .A(n9149), .B(n9150), .Z(n9148) );
  NANDN U17278 ( .A(n9151), .B(n9152), .Z(n9150) );
  NANDN U17279 ( .A(n9152), .B(n9151), .Z(n9147) );
  XOR U17280 ( .A(n9151), .B(n9153), .Z(N64573) );
  XNOR U17281 ( .A(n9149), .B(n9152), .Z(n9153) );
  NAND U17282 ( .A(n9154), .B(n9155), .Z(n9152) );
  NAND U17283 ( .A(n9156), .B(n9157), .Z(n9155) );
  NANDN U17284 ( .A(n9158), .B(n9159), .Z(n9157) );
  NANDN U17285 ( .A(n9159), .B(n9158), .Z(n9154) );
  AND U17286 ( .A(n9160), .B(n9161), .Z(n9149) );
  NAND U17287 ( .A(n9162), .B(n9163), .Z(n9161) );
  NANDN U17288 ( .A(n9164), .B(n9165), .Z(n9163) );
  NANDN U17289 ( .A(n9165), .B(n9164), .Z(n9160) );
  IV U17290 ( .A(n9166), .Z(n9165) );
  AND U17291 ( .A(n9167), .B(n9168), .Z(n9151) );
  NAND U17292 ( .A(n9169), .B(n9170), .Z(n9168) );
  NANDN U17293 ( .A(n9171), .B(n9172), .Z(n9170) );
  NANDN U17294 ( .A(n9172), .B(n9171), .Z(n9167) );
  XOR U17295 ( .A(n9164), .B(n9173), .Z(N64572) );
  XNOR U17296 ( .A(n9162), .B(n9166), .Z(n9173) );
  XOR U17297 ( .A(n9159), .B(n9174), .Z(n9166) );
  XNOR U17298 ( .A(n9156), .B(n9158), .Z(n9174) );
  AND U17299 ( .A(n9175), .B(n9176), .Z(n9158) );
  NANDN U17300 ( .A(n9177), .B(n9178), .Z(n9176) );
  OR U17301 ( .A(n9179), .B(n9180), .Z(n9178) );
  IV U17302 ( .A(n9181), .Z(n9180) );
  NANDN U17303 ( .A(n9181), .B(n9179), .Z(n9175) );
  AND U17304 ( .A(n9182), .B(n9183), .Z(n9156) );
  NAND U17305 ( .A(n9184), .B(n9185), .Z(n9183) );
  NANDN U17306 ( .A(n9186), .B(n9187), .Z(n9185) );
  NANDN U17307 ( .A(n9187), .B(n9186), .Z(n9182) );
  IV U17308 ( .A(n9188), .Z(n9187) );
  NAND U17309 ( .A(n9189), .B(n9190), .Z(n9159) );
  NANDN U17310 ( .A(n9191), .B(n9192), .Z(n9190) );
  NANDN U17311 ( .A(n9193), .B(n9194), .Z(n9192) );
  NANDN U17312 ( .A(n9194), .B(n9193), .Z(n9189) );
  IV U17313 ( .A(n9195), .Z(n9193) );
  AND U17314 ( .A(n9196), .B(n9197), .Z(n9162) );
  NAND U17315 ( .A(n9198), .B(n9199), .Z(n9197) );
  NANDN U17316 ( .A(n9200), .B(n9201), .Z(n9199) );
  NANDN U17317 ( .A(n9201), .B(n9200), .Z(n9196) );
  XOR U17318 ( .A(n9172), .B(n9202), .Z(n9164) );
  XNOR U17319 ( .A(n9169), .B(n9171), .Z(n9202) );
  AND U17320 ( .A(n9203), .B(n9204), .Z(n9171) );
  NANDN U17321 ( .A(n9205), .B(n9206), .Z(n9204) );
  OR U17322 ( .A(n9207), .B(n9208), .Z(n9206) );
  IV U17323 ( .A(n9209), .Z(n9208) );
  NANDN U17324 ( .A(n9209), .B(n9207), .Z(n9203) );
  AND U17325 ( .A(n9210), .B(n9211), .Z(n9169) );
  NAND U17326 ( .A(n9212), .B(n9213), .Z(n9211) );
  NANDN U17327 ( .A(n9214), .B(n9215), .Z(n9213) );
  NANDN U17328 ( .A(n9215), .B(n9214), .Z(n9210) );
  IV U17329 ( .A(n9216), .Z(n9215) );
  NAND U17330 ( .A(n9217), .B(n9218), .Z(n9172) );
  NANDN U17331 ( .A(n9219), .B(n9220), .Z(n9218) );
  NANDN U17332 ( .A(n9221), .B(n9222), .Z(n9220) );
  NANDN U17333 ( .A(n9222), .B(n9221), .Z(n9217) );
  IV U17334 ( .A(n9223), .Z(n9221) );
  XOR U17335 ( .A(n9198), .B(n9224), .Z(N64571) );
  XNOR U17336 ( .A(n9201), .B(n9200), .Z(n9224) );
  XNOR U17337 ( .A(n9212), .B(n9225), .Z(n9200) );
  XNOR U17338 ( .A(n9216), .B(n9214), .Z(n9225) );
  XOR U17339 ( .A(n9222), .B(n9226), .Z(n9214) );
  XNOR U17340 ( .A(n9219), .B(n9223), .Z(n9226) );
  AND U17341 ( .A(n9227), .B(n9228), .Z(n9223) );
  NAND U17342 ( .A(n9229), .B(n9230), .Z(n9228) );
  NAND U17343 ( .A(n9231), .B(n9232), .Z(n9227) );
  AND U17344 ( .A(n9233), .B(n9234), .Z(n9219) );
  NAND U17345 ( .A(n9235), .B(n9236), .Z(n9234) );
  NAND U17346 ( .A(n9237), .B(n9238), .Z(n9233) );
  NANDN U17347 ( .A(n9239), .B(n9240), .Z(n9222) );
  ANDN U17348 ( .B(n9241), .A(n9242), .Z(n9216) );
  XNOR U17349 ( .A(n9207), .B(n9243), .Z(n9212) );
  XNOR U17350 ( .A(n9205), .B(n9209), .Z(n9243) );
  AND U17351 ( .A(n9244), .B(n9245), .Z(n9209) );
  NAND U17352 ( .A(n9246), .B(n9247), .Z(n9245) );
  NAND U17353 ( .A(n9248), .B(n9249), .Z(n9244) );
  AND U17354 ( .A(n9250), .B(n9251), .Z(n9205) );
  NAND U17355 ( .A(n9252), .B(n9253), .Z(n9251) );
  NAND U17356 ( .A(n9254), .B(n9255), .Z(n9250) );
  AND U17357 ( .A(n9256), .B(n9257), .Z(n9207) );
  NAND U17358 ( .A(n9258), .B(n9259), .Z(n9201) );
  XNOR U17359 ( .A(n9184), .B(n9260), .Z(n9198) );
  XNOR U17360 ( .A(n9188), .B(n9186), .Z(n9260) );
  XOR U17361 ( .A(n9194), .B(n9261), .Z(n9186) );
  XNOR U17362 ( .A(n9191), .B(n9195), .Z(n9261) );
  AND U17363 ( .A(n9262), .B(n9263), .Z(n9195) );
  NAND U17364 ( .A(n9264), .B(n9265), .Z(n9263) );
  NAND U17365 ( .A(n9266), .B(n9267), .Z(n9262) );
  AND U17366 ( .A(n9268), .B(n9269), .Z(n9191) );
  NAND U17367 ( .A(n9270), .B(n9271), .Z(n9269) );
  NAND U17368 ( .A(n9272), .B(n9273), .Z(n9268) );
  NANDN U17369 ( .A(n9274), .B(n9275), .Z(n9194) );
  ANDN U17370 ( .B(n9276), .A(n9277), .Z(n9188) );
  XNOR U17371 ( .A(n9179), .B(n9278), .Z(n9184) );
  XNOR U17372 ( .A(n9177), .B(n9181), .Z(n9278) );
  AND U17373 ( .A(n9279), .B(n9280), .Z(n9181) );
  NAND U17374 ( .A(n9281), .B(n9282), .Z(n9280) );
  NAND U17375 ( .A(n9283), .B(n9284), .Z(n9279) );
  AND U17376 ( .A(n9285), .B(n9286), .Z(n9177) );
  NAND U17377 ( .A(n9287), .B(n9288), .Z(n9286) );
  NAND U17378 ( .A(n9289), .B(n9290), .Z(n9285) );
  AND U17379 ( .A(n9291), .B(n9292), .Z(n9179) );
  XOR U17380 ( .A(n9259), .B(n9258), .Z(N64570) );
  XNOR U17381 ( .A(n9276), .B(n9277), .Z(n9258) );
  XNOR U17382 ( .A(n9291), .B(n9292), .Z(n9277) );
  XOR U17383 ( .A(n9288), .B(n9287), .Z(n9292) );
  XOR U17384 ( .A(y[7356]), .B(x[7356]), .Z(n9287) );
  XOR U17385 ( .A(n9290), .B(n9289), .Z(n9288) );
  XOR U17386 ( .A(y[7358]), .B(x[7358]), .Z(n9289) );
  XOR U17387 ( .A(y[7357]), .B(x[7357]), .Z(n9290) );
  XOR U17388 ( .A(n9282), .B(n9281), .Z(n9291) );
  XOR U17389 ( .A(n9284), .B(n9283), .Z(n9281) );
  XOR U17390 ( .A(y[7355]), .B(x[7355]), .Z(n9283) );
  XOR U17391 ( .A(y[7354]), .B(x[7354]), .Z(n9284) );
  XOR U17392 ( .A(y[7353]), .B(x[7353]), .Z(n9282) );
  XNOR U17393 ( .A(n9275), .B(n9274), .Z(n9276) );
  XNOR U17394 ( .A(n9271), .B(n9270), .Z(n9274) );
  XOR U17395 ( .A(n9273), .B(n9272), .Z(n9270) );
  XOR U17396 ( .A(y[7352]), .B(x[7352]), .Z(n9272) );
  XOR U17397 ( .A(y[7351]), .B(x[7351]), .Z(n9273) );
  XOR U17398 ( .A(y[7350]), .B(x[7350]), .Z(n9271) );
  XOR U17399 ( .A(n9265), .B(n9264), .Z(n9275) );
  XOR U17400 ( .A(n9267), .B(n9266), .Z(n9264) );
  XOR U17401 ( .A(y[7349]), .B(x[7349]), .Z(n9266) );
  XOR U17402 ( .A(y[7348]), .B(x[7348]), .Z(n9267) );
  XOR U17403 ( .A(y[7347]), .B(x[7347]), .Z(n9265) );
  XNOR U17404 ( .A(n9241), .B(n9242), .Z(n9259) );
  XNOR U17405 ( .A(n9256), .B(n9257), .Z(n9242) );
  XOR U17406 ( .A(n9253), .B(n9252), .Z(n9257) );
  XOR U17407 ( .A(y[7344]), .B(x[7344]), .Z(n9252) );
  XOR U17408 ( .A(n9255), .B(n9254), .Z(n9253) );
  XOR U17409 ( .A(y[7346]), .B(x[7346]), .Z(n9254) );
  XOR U17410 ( .A(y[7345]), .B(x[7345]), .Z(n9255) );
  XOR U17411 ( .A(n9247), .B(n9246), .Z(n9256) );
  XOR U17412 ( .A(n9249), .B(n9248), .Z(n9246) );
  XOR U17413 ( .A(y[7343]), .B(x[7343]), .Z(n9248) );
  XOR U17414 ( .A(y[7342]), .B(x[7342]), .Z(n9249) );
  XOR U17415 ( .A(y[7341]), .B(x[7341]), .Z(n9247) );
  XNOR U17416 ( .A(n9240), .B(n9239), .Z(n9241) );
  XNOR U17417 ( .A(n9236), .B(n9235), .Z(n9239) );
  XOR U17418 ( .A(n9238), .B(n9237), .Z(n9235) );
  XOR U17419 ( .A(y[7340]), .B(x[7340]), .Z(n9237) );
  XOR U17420 ( .A(y[7339]), .B(x[7339]), .Z(n9238) );
  XOR U17421 ( .A(y[7338]), .B(x[7338]), .Z(n9236) );
  XOR U17422 ( .A(n9230), .B(n9229), .Z(n9240) );
  XOR U17423 ( .A(n9232), .B(n9231), .Z(n9229) );
  XOR U17424 ( .A(y[7337]), .B(x[7337]), .Z(n9231) );
  XOR U17425 ( .A(y[7336]), .B(x[7336]), .Z(n9232) );
  XOR U17426 ( .A(y[7335]), .B(x[7335]), .Z(n9230) );
  NAND U17427 ( .A(n9293), .B(n9294), .Z(N64561) );
  NAND U17428 ( .A(n9295), .B(n9296), .Z(n9294) );
  NANDN U17429 ( .A(n9297), .B(n9298), .Z(n9296) );
  NANDN U17430 ( .A(n9298), .B(n9297), .Z(n9293) );
  XOR U17431 ( .A(n9297), .B(n9299), .Z(N64560) );
  XNOR U17432 ( .A(n9295), .B(n9298), .Z(n9299) );
  NAND U17433 ( .A(n9300), .B(n9301), .Z(n9298) );
  NAND U17434 ( .A(n9302), .B(n9303), .Z(n9301) );
  NANDN U17435 ( .A(n9304), .B(n9305), .Z(n9303) );
  NANDN U17436 ( .A(n9305), .B(n9304), .Z(n9300) );
  AND U17437 ( .A(n9306), .B(n9307), .Z(n9295) );
  NAND U17438 ( .A(n9308), .B(n9309), .Z(n9307) );
  NANDN U17439 ( .A(n9310), .B(n9311), .Z(n9309) );
  NANDN U17440 ( .A(n9311), .B(n9310), .Z(n9306) );
  IV U17441 ( .A(n9312), .Z(n9311) );
  AND U17442 ( .A(n9313), .B(n9314), .Z(n9297) );
  NAND U17443 ( .A(n9315), .B(n9316), .Z(n9314) );
  NANDN U17444 ( .A(n9317), .B(n9318), .Z(n9316) );
  NANDN U17445 ( .A(n9318), .B(n9317), .Z(n9313) );
  XOR U17446 ( .A(n9310), .B(n9319), .Z(N64559) );
  XNOR U17447 ( .A(n9308), .B(n9312), .Z(n9319) );
  XOR U17448 ( .A(n9305), .B(n9320), .Z(n9312) );
  XNOR U17449 ( .A(n9302), .B(n9304), .Z(n9320) );
  AND U17450 ( .A(n9321), .B(n9322), .Z(n9304) );
  NANDN U17451 ( .A(n9323), .B(n9324), .Z(n9322) );
  OR U17452 ( .A(n9325), .B(n9326), .Z(n9324) );
  IV U17453 ( .A(n9327), .Z(n9326) );
  NANDN U17454 ( .A(n9327), .B(n9325), .Z(n9321) );
  AND U17455 ( .A(n9328), .B(n9329), .Z(n9302) );
  NAND U17456 ( .A(n9330), .B(n9331), .Z(n9329) );
  NANDN U17457 ( .A(n9332), .B(n9333), .Z(n9331) );
  NANDN U17458 ( .A(n9333), .B(n9332), .Z(n9328) );
  IV U17459 ( .A(n9334), .Z(n9333) );
  NAND U17460 ( .A(n9335), .B(n9336), .Z(n9305) );
  NANDN U17461 ( .A(n9337), .B(n9338), .Z(n9336) );
  NANDN U17462 ( .A(n9339), .B(n9340), .Z(n9338) );
  NANDN U17463 ( .A(n9340), .B(n9339), .Z(n9335) );
  IV U17464 ( .A(n9341), .Z(n9339) );
  AND U17465 ( .A(n9342), .B(n9343), .Z(n9308) );
  NAND U17466 ( .A(n9344), .B(n9345), .Z(n9343) );
  NANDN U17467 ( .A(n9346), .B(n9347), .Z(n9345) );
  NANDN U17468 ( .A(n9347), .B(n9346), .Z(n9342) );
  XOR U17469 ( .A(n9318), .B(n9348), .Z(n9310) );
  XNOR U17470 ( .A(n9315), .B(n9317), .Z(n9348) );
  AND U17471 ( .A(n9349), .B(n9350), .Z(n9317) );
  NANDN U17472 ( .A(n9351), .B(n9352), .Z(n9350) );
  OR U17473 ( .A(n9353), .B(n9354), .Z(n9352) );
  IV U17474 ( .A(n9355), .Z(n9354) );
  NANDN U17475 ( .A(n9355), .B(n9353), .Z(n9349) );
  AND U17476 ( .A(n9356), .B(n9357), .Z(n9315) );
  NAND U17477 ( .A(n9358), .B(n9359), .Z(n9357) );
  NANDN U17478 ( .A(n9360), .B(n9361), .Z(n9359) );
  NANDN U17479 ( .A(n9361), .B(n9360), .Z(n9356) );
  IV U17480 ( .A(n9362), .Z(n9361) );
  NAND U17481 ( .A(n9363), .B(n9364), .Z(n9318) );
  NANDN U17482 ( .A(n9365), .B(n9366), .Z(n9364) );
  NANDN U17483 ( .A(n9367), .B(n9368), .Z(n9366) );
  NANDN U17484 ( .A(n9368), .B(n9367), .Z(n9363) );
  IV U17485 ( .A(n9369), .Z(n9367) );
  XOR U17486 ( .A(n9344), .B(n9370), .Z(N64558) );
  XNOR U17487 ( .A(n9347), .B(n9346), .Z(n9370) );
  XNOR U17488 ( .A(n9358), .B(n9371), .Z(n9346) );
  XNOR U17489 ( .A(n9362), .B(n9360), .Z(n9371) );
  XOR U17490 ( .A(n9368), .B(n9372), .Z(n9360) );
  XNOR U17491 ( .A(n9365), .B(n9369), .Z(n9372) );
  AND U17492 ( .A(n9373), .B(n9374), .Z(n9369) );
  NAND U17493 ( .A(n9375), .B(n9376), .Z(n9374) );
  NAND U17494 ( .A(n9377), .B(n9378), .Z(n9373) );
  AND U17495 ( .A(n9379), .B(n9380), .Z(n9365) );
  NAND U17496 ( .A(n9381), .B(n9382), .Z(n9380) );
  NAND U17497 ( .A(n9383), .B(n9384), .Z(n9379) );
  NANDN U17498 ( .A(n9385), .B(n9386), .Z(n9368) );
  ANDN U17499 ( .B(n9387), .A(n9388), .Z(n9362) );
  XNOR U17500 ( .A(n9353), .B(n9389), .Z(n9358) );
  XNOR U17501 ( .A(n9351), .B(n9355), .Z(n9389) );
  AND U17502 ( .A(n9390), .B(n9391), .Z(n9355) );
  NAND U17503 ( .A(n9392), .B(n9393), .Z(n9391) );
  NAND U17504 ( .A(n9394), .B(n9395), .Z(n9390) );
  AND U17505 ( .A(n9396), .B(n9397), .Z(n9351) );
  NAND U17506 ( .A(n9398), .B(n9399), .Z(n9397) );
  NAND U17507 ( .A(n9400), .B(n9401), .Z(n9396) );
  AND U17508 ( .A(n9402), .B(n9403), .Z(n9353) );
  NAND U17509 ( .A(n9404), .B(n9405), .Z(n9347) );
  XNOR U17510 ( .A(n9330), .B(n9406), .Z(n9344) );
  XNOR U17511 ( .A(n9334), .B(n9332), .Z(n9406) );
  XOR U17512 ( .A(n9340), .B(n9407), .Z(n9332) );
  XNOR U17513 ( .A(n9337), .B(n9341), .Z(n9407) );
  AND U17514 ( .A(n9408), .B(n9409), .Z(n9341) );
  NAND U17515 ( .A(n9410), .B(n9411), .Z(n9409) );
  NAND U17516 ( .A(n9412), .B(n9413), .Z(n9408) );
  AND U17517 ( .A(n9414), .B(n9415), .Z(n9337) );
  NAND U17518 ( .A(n9416), .B(n9417), .Z(n9415) );
  NAND U17519 ( .A(n9418), .B(n9419), .Z(n9414) );
  NANDN U17520 ( .A(n9420), .B(n9421), .Z(n9340) );
  ANDN U17521 ( .B(n9422), .A(n9423), .Z(n9334) );
  XNOR U17522 ( .A(n9325), .B(n9424), .Z(n9330) );
  XNOR U17523 ( .A(n9323), .B(n9327), .Z(n9424) );
  AND U17524 ( .A(n9425), .B(n9426), .Z(n9327) );
  NAND U17525 ( .A(n9427), .B(n9428), .Z(n9426) );
  NAND U17526 ( .A(n9429), .B(n9430), .Z(n9425) );
  AND U17527 ( .A(n9431), .B(n9432), .Z(n9323) );
  NAND U17528 ( .A(n9433), .B(n9434), .Z(n9432) );
  NAND U17529 ( .A(n9435), .B(n9436), .Z(n9431) );
  AND U17530 ( .A(n9437), .B(n9438), .Z(n9325) );
  XOR U17531 ( .A(n9405), .B(n9404), .Z(N64557) );
  XNOR U17532 ( .A(n9422), .B(n9423), .Z(n9404) );
  XNOR U17533 ( .A(n9437), .B(n9438), .Z(n9423) );
  XOR U17534 ( .A(n9434), .B(n9433), .Z(n9438) );
  XOR U17535 ( .A(y[7332]), .B(x[7332]), .Z(n9433) );
  XOR U17536 ( .A(n9436), .B(n9435), .Z(n9434) );
  XOR U17537 ( .A(y[7334]), .B(x[7334]), .Z(n9435) );
  XOR U17538 ( .A(y[7333]), .B(x[7333]), .Z(n9436) );
  XOR U17539 ( .A(n9428), .B(n9427), .Z(n9437) );
  XOR U17540 ( .A(n9430), .B(n9429), .Z(n9427) );
  XOR U17541 ( .A(y[7331]), .B(x[7331]), .Z(n9429) );
  XOR U17542 ( .A(y[7330]), .B(x[7330]), .Z(n9430) );
  XOR U17543 ( .A(y[7329]), .B(x[7329]), .Z(n9428) );
  XNOR U17544 ( .A(n9421), .B(n9420), .Z(n9422) );
  XNOR U17545 ( .A(n9417), .B(n9416), .Z(n9420) );
  XOR U17546 ( .A(n9419), .B(n9418), .Z(n9416) );
  XOR U17547 ( .A(y[7328]), .B(x[7328]), .Z(n9418) );
  XOR U17548 ( .A(y[7327]), .B(x[7327]), .Z(n9419) );
  XOR U17549 ( .A(y[7326]), .B(x[7326]), .Z(n9417) );
  XOR U17550 ( .A(n9411), .B(n9410), .Z(n9421) );
  XOR U17551 ( .A(n9413), .B(n9412), .Z(n9410) );
  XOR U17552 ( .A(y[7325]), .B(x[7325]), .Z(n9412) );
  XOR U17553 ( .A(y[7324]), .B(x[7324]), .Z(n9413) );
  XOR U17554 ( .A(y[7323]), .B(x[7323]), .Z(n9411) );
  XNOR U17555 ( .A(n9387), .B(n9388), .Z(n9405) );
  XNOR U17556 ( .A(n9402), .B(n9403), .Z(n9388) );
  XOR U17557 ( .A(n9399), .B(n9398), .Z(n9403) );
  XOR U17558 ( .A(y[7320]), .B(x[7320]), .Z(n9398) );
  XOR U17559 ( .A(n9401), .B(n9400), .Z(n9399) );
  XOR U17560 ( .A(y[7322]), .B(x[7322]), .Z(n9400) );
  XOR U17561 ( .A(y[7321]), .B(x[7321]), .Z(n9401) );
  XOR U17562 ( .A(n9393), .B(n9392), .Z(n9402) );
  XOR U17563 ( .A(n9395), .B(n9394), .Z(n9392) );
  XOR U17564 ( .A(y[7319]), .B(x[7319]), .Z(n9394) );
  XOR U17565 ( .A(y[7318]), .B(x[7318]), .Z(n9395) );
  XOR U17566 ( .A(y[7317]), .B(x[7317]), .Z(n9393) );
  XNOR U17567 ( .A(n9386), .B(n9385), .Z(n9387) );
  XNOR U17568 ( .A(n9382), .B(n9381), .Z(n9385) );
  XOR U17569 ( .A(n9384), .B(n9383), .Z(n9381) );
  XOR U17570 ( .A(y[7316]), .B(x[7316]), .Z(n9383) );
  XOR U17571 ( .A(y[7315]), .B(x[7315]), .Z(n9384) );
  XOR U17572 ( .A(y[7314]), .B(x[7314]), .Z(n9382) );
  XOR U17573 ( .A(n9376), .B(n9375), .Z(n9386) );
  XOR U17574 ( .A(n9378), .B(n9377), .Z(n9375) );
  XOR U17575 ( .A(y[7313]), .B(x[7313]), .Z(n9377) );
  XOR U17576 ( .A(y[7312]), .B(x[7312]), .Z(n9378) );
  XOR U17577 ( .A(y[7311]), .B(x[7311]), .Z(n9376) );
  NAND U17578 ( .A(n9439), .B(n9440), .Z(N64548) );
  NAND U17579 ( .A(n9441), .B(n9442), .Z(n9440) );
  NANDN U17580 ( .A(n9443), .B(n9444), .Z(n9442) );
  NANDN U17581 ( .A(n9444), .B(n9443), .Z(n9439) );
  XOR U17582 ( .A(n9443), .B(n9445), .Z(N64547) );
  XNOR U17583 ( .A(n9441), .B(n9444), .Z(n9445) );
  NAND U17584 ( .A(n9446), .B(n9447), .Z(n9444) );
  NAND U17585 ( .A(n9448), .B(n9449), .Z(n9447) );
  NANDN U17586 ( .A(n9450), .B(n9451), .Z(n9449) );
  NANDN U17587 ( .A(n9451), .B(n9450), .Z(n9446) );
  AND U17588 ( .A(n9452), .B(n9453), .Z(n9441) );
  NAND U17589 ( .A(n9454), .B(n9455), .Z(n9453) );
  NANDN U17590 ( .A(n9456), .B(n9457), .Z(n9455) );
  NANDN U17591 ( .A(n9457), .B(n9456), .Z(n9452) );
  IV U17592 ( .A(n9458), .Z(n9457) );
  AND U17593 ( .A(n9459), .B(n9460), .Z(n9443) );
  NAND U17594 ( .A(n9461), .B(n9462), .Z(n9460) );
  NANDN U17595 ( .A(n9463), .B(n9464), .Z(n9462) );
  NANDN U17596 ( .A(n9464), .B(n9463), .Z(n9459) );
  XOR U17597 ( .A(n9456), .B(n9465), .Z(N64546) );
  XNOR U17598 ( .A(n9454), .B(n9458), .Z(n9465) );
  XOR U17599 ( .A(n9451), .B(n9466), .Z(n9458) );
  XNOR U17600 ( .A(n9448), .B(n9450), .Z(n9466) );
  AND U17601 ( .A(n9467), .B(n9468), .Z(n9450) );
  NANDN U17602 ( .A(n9469), .B(n9470), .Z(n9468) );
  OR U17603 ( .A(n9471), .B(n9472), .Z(n9470) );
  IV U17604 ( .A(n9473), .Z(n9472) );
  NANDN U17605 ( .A(n9473), .B(n9471), .Z(n9467) );
  AND U17606 ( .A(n9474), .B(n9475), .Z(n9448) );
  NAND U17607 ( .A(n9476), .B(n9477), .Z(n9475) );
  NANDN U17608 ( .A(n9478), .B(n9479), .Z(n9477) );
  NANDN U17609 ( .A(n9479), .B(n9478), .Z(n9474) );
  IV U17610 ( .A(n9480), .Z(n9479) );
  NAND U17611 ( .A(n9481), .B(n9482), .Z(n9451) );
  NANDN U17612 ( .A(n9483), .B(n9484), .Z(n9482) );
  NANDN U17613 ( .A(n9485), .B(n9486), .Z(n9484) );
  NANDN U17614 ( .A(n9486), .B(n9485), .Z(n9481) );
  IV U17615 ( .A(n9487), .Z(n9485) );
  AND U17616 ( .A(n9488), .B(n9489), .Z(n9454) );
  NAND U17617 ( .A(n9490), .B(n9491), .Z(n9489) );
  NANDN U17618 ( .A(n9492), .B(n9493), .Z(n9491) );
  NANDN U17619 ( .A(n9493), .B(n9492), .Z(n9488) );
  XOR U17620 ( .A(n9464), .B(n9494), .Z(n9456) );
  XNOR U17621 ( .A(n9461), .B(n9463), .Z(n9494) );
  AND U17622 ( .A(n9495), .B(n9496), .Z(n9463) );
  NANDN U17623 ( .A(n9497), .B(n9498), .Z(n9496) );
  OR U17624 ( .A(n9499), .B(n9500), .Z(n9498) );
  IV U17625 ( .A(n9501), .Z(n9500) );
  NANDN U17626 ( .A(n9501), .B(n9499), .Z(n9495) );
  AND U17627 ( .A(n9502), .B(n9503), .Z(n9461) );
  NAND U17628 ( .A(n9504), .B(n9505), .Z(n9503) );
  NANDN U17629 ( .A(n9506), .B(n9507), .Z(n9505) );
  NANDN U17630 ( .A(n9507), .B(n9506), .Z(n9502) );
  IV U17631 ( .A(n9508), .Z(n9507) );
  NAND U17632 ( .A(n9509), .B(n9510), .Z(n9464) );
  NANDN U17633 ( .A(n9511), .B(n9512), .Z(n9510) );
  NANDN U17634 ( .A(n9513), .B(n9514), .Z(n9512) );
  NANDN U17635 ( .A(n9514), .B(n9513), .Z(n9509) );
  IV U17636 ( .A(n9515), .Z(n9513) );
  XOR U17637 ( .A(n9490), .B(n9516), .Z(N64545) );
  XNOR U17638 ( .A(n9493), .B(n9492), .Z(n9516) );
  XNOR U17639 ( .A(n9504), .B(n9517), .Z(n9492) );
  XNOR U17640 ( .A(n9508), .B(n9506), .Z(n9517) );
  XOR U17641 ( .A(n9514), .B(n9518), .Z(n9506) );
  XNOR U17642 ( .A(n9511), .B(n9515), .Z(n9518) );
  AND U17643 ( .A(n9519), .B(n9520), .Z(n9515) );
  NAND U17644 ( .A(n9521), .B(n9522), .Z(n9520) );
  NAND U17645 ( .A(n9523), .B(n9524), .Z(n9519) );
  AND U17646 ( .A(n9525), .B(n9526), .Z(n9511) );
  NAND U17647 ( .A(n9527), .B(n9528), .Z(n9526) );
  NAND U17648 ( .A(n9529), .B(n9530), .Z(n9525) );
  NANDN U17649 ( .A(n9531), .B(n9532), .Z(n9514) );
  ANDN U17650 ( .B(n9533), .A(n9534), .Z(n9508) );
  XNOR U17651 ( .A(n9499), .B(n9535), .Z(n9504) );
  XNOR U17652 ( .A(n9497), .B(n9501), .Z(n9535) );
  AND U17653 ( .A(n9536), .B(n9537), .Z(n9501) );
  NAND U17654 ( .A(n9538), .B(n9539), .Z(n9537) );
  NAND U17655 ( .A(n9540), .B(n9541), .Z(n9536) );
  AND U17656 ( .A(n9542), .B(n9543), .Z(n9497) );
  NAND U17657 ( .A(n9544), .B(n9545), .Z(n9543) );
  NAND U17658 ( .A(n9546), .B(n9547), .Z(n9542) );
  AND U17659 ( .A(n9548), .B(n9549), .Z(n9499) );
  NAND U17660 ( .A(n9550), .B(n9551), .Z(n9493) );
  XNOR U17661 ( .A(n9476), .B(n9552), .Z(n9490) );
  XNOR U17662 ( .A(n9480), .B(n9478), .Z(n9552) );
  XOR U17663 ( .A(n9486), .B(n9553), .Z(n9478) );
  XNOR U17664 ( .A(n9483), .B(n9487), .Z(n9553) );
  AND U17665 ( .A(n9554), .B(n9555), .Z(n9487) );
  NAND U17666 ( .A(n9556), .B(n9557), .Z(n9555) );
  NAND U17667 ( .A(n9558), .B(n9559), .Z(n9554) );
  AND U17668 ( .A(n9560), .B(n9561), .Z(n9483) );
  NAND U17669 ( .A(n9562), .B(n9563), .Z(n9561) );
  NAND U17670 ( .A(n9564), .B(n9565), .Z(n9560) );
  NANDN U17671 ( .A(n9566), .B(n9567), .Z(n9486) );
  ANDN U17672 ( .B(n9568), .A(n9569), .Z(n9480) );
  XNOR U17673 ( .A(n9471), .B(n9570), .Z(n9476) );
  XNOR U17674 ( .A(n9469), .B(n9473), .Z(n9570) );
  AND U17675 ( .A(n9571), .B(n9572), .Z(n9473) );
  NAND U17676 ( .A(n9573), .B(n9574), .Z(n9572) );
  NAND U17677 ( .A(n9575), .B(n9576), .Z(n9571) );
  AND U17678 ( .A(n9577), .B(n9578), .Z(n9469) );
  NAND U17679 ( .A(n9579), .B(n9580), .Z(n9578) );
  NAND U17680 ( .A(n9581), .B(n9582), .Z(n9577) );
  AND U17681 ( .A(n9583), .B(n9584), .Z(n9471) );
  XOR U17682 ( .A(n9551), .B(n9550), .Z(N64544) );
  XNOR U17683 ( .A(n9568), .B(n9569), .Z(n9550) );
  XNOR U17684 ( .A(n9583), .B(n9584), .Z(n9569) );
  XOR U17685 ( .A(n9580), .B(n9579), .Z(n9584) );
  XOR U17686 ( .A(y[7308]), .B(x[7308]), .Z(n9579) );
  XOR U17687 ( .A(n9582), .B(n9581), .Z(n9580) );
  XOR U17688 ( .A(y[7310]), .B(x[7310]), .Z(n9581) );
  XOR U17689 ( .A(y[7309]), .B(x[7309]), .Z(n9582) );
  XOR U17690 ( .A(n9574), .B(n9573), .Z(n9583) );
  XOR U17691 ( .A(n9576), .B(n9575), .Z(n9573) );
  XOR U17692 ( .A(y[7307]), .B(x[7307]), .Z(n9575) );
  XOR U17693 ( .A(y[7306]), .B(x[7306]), .Z(n9576) );
  XOR U17694 ( .A(y[7305]), .B(x[7305]), .Z(n9574) );
  XNOR U17695 ( .A(n9567), .B(n9566), .Z(n9568) );
  XNOR U17696 ( .A(n9563), .B(n9562), .Z(n9566) );
  XOR U17697 ( .A(n9565), .B(n9564), .Z(n9562) );
  XOR U17698 ( .A(y[7304]), .B(x[7304]), .Z(n9564) );
  XOR U17699 ( .A(y[7303]), .B(x[7303]), .Z(n9565) );
  XOR U17700 ( .A(y[7302]), .B(x[7302]), .Z(n9563) );
  XOR U17701 ( .A(n9557), .B(n9556), .Z(n9567) );
  XOR U17702 ( .A(n9559), .B(n9558), .Z(n9556) );
  XOR U17703 ( .A(y[7301]), .B(x[7301]), .Z(n9558) );
  XOR U17704 ( .A(y[7300]), .B(x[7300]), .Z(n9559) );
  XOR U17705 ( .A(y[7299]), .B(x[7299]), .Z(n9557) );
  XNOR U17706 ( .A(n9533), .B(n9534), .Z(n9551) );
  XNOR U17707 ( .A(n9548), .B(n9549), .Z(n9534) );
  XOR U17708 ( .A(n9545), .B(n9544), .Z(n9549) );
  XOR U17709 ( .A(y[7296]), .B(x[7296]), .Z(n9544) );
  XOR U17710 ( .A(n9547), .B(n9546), .Z(n9545) );
  XOR U17711 ( .A(y[7298]), .B(x[7298]), .Z(n9546) );
  XOR U17712 ( .A(y[7297]), .B(x[7297]), .Z(n9547) );
  XOR U17713 ( .A(n9539), .B(n9538), .Z(n9548) );
  XOR U17714 ( .A(n9541), .B(n9540), .Z(n9538) );
  XOR U17715 ( .A(y[7295]), .B(x[7295]), .Z(n9540) );
  XOR U17716 ( .A(y[7294]), .B(x[7294]), .Z(n9541) );
  XOR U17717 ( .A(y[7293]), .B(x[7293]), .Z(n9539) );
  XNOR U17718 ( .A(n9532), .B(n9531), .Z(n9533) );
  XNOR U17719 ( .A(n9528), .B(n9527), .Z(n9531) );
  XOR U17720 ( .A(n9530), .B(n9529), .Z(n9527) );
  XOR U17721 ( .A(y[7292]), .B(x[7292]), .Z(n9529) );
  XOR U17722 ( .A(y[7291]), .B(x[7291]), .Z(n9530) );
  XOR U17723 ( .A(y[7290]), .B(x[7290]), .Z(n9528) );
  XOR U17724 ( .A(n9522), .B(n9521), .Z(n9532) );
  XOR U17725 ( .A(n9524), .B(n9523), .Z(n9521) );
  XOR U17726 ( .A(y[7289]), .B(x[7289]), .Z(n9523) );
  XOR U17727 ( .A(y[7288]), .B(x[7288]), .Z(n9524) );
  XOR U17728 ( .A(y[7287]), .B(x[7287]), .Z(n9522) );
  NAND U17729 ( .A(n9585), .B(n9586), .Z(N64535) );
  NAND U17730 ( .A(n9587), .B(n9588), .Z(n9586) );
  NANDN U17731 ( .A(n9589), .B(n9590), .Z(n9588) );
  NANDN U17732 ( .A(n9590), .B(n9589), .Z(n9585) );
  XOR U17733 ( .A(n9589), .B(n9591), .Z(N64534) );
  XNOR U17734 ( .A(n9587), .B(n9590), .Z(n9591) );
  NAND U17735 ( .A(n9592), .B(n9593), .Z(n9590) );
  NAND U17736 ( .A(n9594), .B(n9595), .Z(n9593) );
  NANDN U17737 ( .A(n9596), .B(n9597), .Z(n9595) );
  NANDN U17738 ( .A(n9597), .B(n9596), .Z(n9592) );
  AND U17739 ( .A(n9598), .B(n9599), .Z(n9587) );
  NAND U17740 ( .A(n9600), .B(n9601), .Z(n9599) );
  NANDN U17741 ( .A(n9602), .B(n9603), .Z(n9601) );
  NANDN U17742 ( .A(n9603), .B(n9602), .Z(n9598) );
  IV U17743 ( .A(n9604), .Z(n9603) );
  AND U17744 ( .A(n9605), .B(n9606), .Z(n9589) );
  NAND U17745 ( .A(n9607), .B(n9608), .Z(n9606) );
  NANDN U17746 ( .A(n9609), .B(n9610), .Z(n9608) );
  NANDN U17747 ( .A(n9610), .B(n9609), .Z(n9605) );
  XOR U17748 ( .A(n9602), .B(n9611), .Z(N64533) );
  XNOR U17749 ( .A(n9600), .B(n9604), .Z(n9611) );
  XOR U17750 ( .A(n9597), .B(n9612), .Z(n9604) );
  XNOR U17751 ( .A(n9594), .B(n9596), .Z(n9612) );
  AND U17752 ( .A(n9613), .B(n9614), .Z(n9596) );
  NANDN U17753 ( .A(n9615), .B(n9616), .Z(n9614) );
  OR U17754 ( .A(n9617), .B(n9618), .Z(n9616) );
  IV U17755 ( .A(n9619), .Z(n9618) );
  NANDN U17756 ( .A(n9619), .B(n9617), .Z(n9613) );
  AND U17757 ( .A(n9620), .B(n9621), .Z(n9594) );
  NAND U17758 ( .A(n9622), .B(n9623), .Z(n9621) );
  NANDN U17759 ( .A(n9624), .B(n9625), .Z(n9623) );
  NANDN U17760 ( .A(n9625), .B(n9624), .Z(n9620) );
  IV U17761 ( .A(n9626), .Z(n9625) );
  NAND U17762 ( .A(n9627), .B(n9628), .Z(n9597) );
  NANDN U17763 ( .A(n9629), .B(n9630), .Z(n9628) );
  NANDN U17764 ( .A(n9631), .B(n9632), .Z(n9630) );
  NANDN U17765 ( .A(n9632), .B(n9631), .Z(n9627) );
  IV U17766 ( .A(n9633), .Z(n9631) );
  AND U17767 ( .A(n9634), .B(n9635), .Z(n9600) );
  NAND U17768 ( .A(n9636), .B(n9637), .Z(n9635) );
  NANDN U17769 ( .A(n9638), .B(n9639), .Z(n9637) );
  NANDN U17770 ( .A(n9639), .B(n9638), .Z(n9634) );
  XOR U17771 ( .A(n9610), .B(n9640), .Z(n9602) );
  XNOR U17772 ( .A(n9607), .B(n9609), .Z(n9640) );
  AND U17773 ( .A(n9641), .B(n9642), .Z(n9609) );
  NANDN U17774 ( .A(n9643), .B(n9644), .Z(n9642) );
  OR U17775 ( .A(n9645), .B(n9646), .Z(n9644) );
  IV U17776 ( .A(n9647), .Z(n9646) );
  NANDN U17777 ( .A(n9647), .B(n9645), .Z(n9641) );
  AND U17778 ( .A(n9648), .B(n9649), .Z(n9607) );
  NAND U17779 ( .A(n9650), .B(n9651), .Z(n9649) );
  NANDN U17780 ( .A(n9652), .B(n9653), .Z(n9651) );
  NANDN U17781 ( .A(n9653), .B(n9652), .Z(n9648) );
  IV U17782 ( .A(n9654), .Z(n9653) );
  NAND U17783 ( .A(n9655), .B(n9656), .Z(n9610) );
  NANDN U17784 ( .A(n9657), .B(n9658), .Z(n9656) );
  NANDN U17785 ( .A(n9659), .B(n9660), .Z(n9658) );
  NANDN U17786 ( .A(n9660), .B(n9659), .Z(n9655) );
  IV U17787 ( .A(n9661), .Z(n9659) );
  XOR U17788 ( .A(n9636), .B(n9662), .Z(N64532) );
  XNOR U17789 ( .A(n9639), .B(n9638), .Z(n9662) );
  XNOR U17790 ( .A(n9650), .B(n9663), .Z(n9638) );
  XNOR U17791 ( .A(n9654), .B(n9652), .Z(n9663) );
  XOR U17792 ( .A(n9660), .B(n9664), .Z(n9652) );
  XNOR U17793 ( .A(n9657), .B(n9661), .Z(n9664) );
  AND U17794 ( .A(n9665), .B(n9666), .Z(n9661) );
  NAND U17795 ( .A(n9667), .B(n9668), .Z(n9666) );
  NAND U17796 ( .A(n9669), .B(n9670), .Z(n9665) );
  AND U17797 ( .A(n9671), .B(n9672), .Z(n9657) );
  NAND U17798 ( .A(n9673), .B(n9674), .Z(n9672) );
  NAND U17799 ( .A(n9675), .B(n9676), .Z(n9671) );
  NANDN U17800 ( .A(n9677), .B(n9678), .Z(n9660) );
  ANDN U17801 ( .B(n9679), .A(n9680), .Z(n9654) );
  XNOR U17802 ( .A(n9645), .B(n9681), .Z(n9650) );
  XNOR U17803 ( .A(n9643), .B(n9647), .Z(n9681) );
  AND U17804 ( .A(n9682), .B(n9683), .Z(n9647) );
  NAND U17805 ( .A(n9684), .B(n9685), .Z(n9683) );
  NAND U17806 ( .A(n9686), .B(n9687), .Z(n9682) );
  AND U17807 ( .A(n9688), .B(n9689), .Z(n9643) );
  NAND U17808 ( .A(n9690), .B(n9691), .Z(n9689) );
  NAND U17809 ( .A(n9692), .B(n9693), .Z(n9688) );
  AND U17810 ( .A(n9694), .B(n9695), .Z(n9645) );
  NAND U17811 ( .A(n9696), .B(n9697), .Z(n9639) );
  XNOR U17812 ( .A(n9622), .B(n9698), .Z(n9636) );
  XNOR U17813 ( .A(n9626), .B(n9624), .Z(n9698) );
  XOR U17814 ( .A(n9632), .B(n9699), .Z(n9624) );
  XNOR U17815 ( .A(n9629), .B(n9633), .Z(n9699) );
  AND U17816 ( .A(n9700), .B(n9701), .Z(n9633) );
  NAND U17817 ( .A(n9702), .B(n9703), .Z(n9701) );
  NAND U17818 ( .A(n9704), .B(n9705), .Z(n9700) );
  AND U17819 ( .A(n9706), .B(n9707), .Z(n9629) );
  NAND U17820 ( .A(n9708), .B(n9709), .Z(n9707) );
  NAND U17821 ( .A(n9710), .B(n9711), .Z(n9706) );
  NANDN U17822 ( .A(n9712), .B(n9713), .Z(n9632) );
  ANDN U17823 ( .B(n9714), .A(n9715), .Z(n9626) );
  XNOR U17824 ( .A(n9617), .B(n9716), .Z(n9622) );
  XNOR U17825 ( .A(n9615), .B(n9619), .Z(n9716) );
  AND U17826 ( .A(n9717), .B(n9718), .Z(n9619) );
  NAND U17827 ( .A(n9719), .B(n9720), .Z(n9718) );
  NAND U17828 ( .A(n9721), .B(n9722), .Z(n9717) );
  AND U17829 ( .A(n9723), .B(n9724), .Z(n9615) );
  NAND U17830 ( .A(n9725), .B(n9726), .Z(n9724) );
  NAND U17831 ( .A(n9727), .B(n9728), .Z(n9723) );
  AND U17832 ( .A(n9729), .B(n9730), .Z(n9617) );
  XOR U17833 ( .A(n9697), .B(n9696), .Z(N64531) );
  XNOR U17834 ( .A(n9714), .B(n9715), .Z(n9696) );
  XNOR U17835 ( .A(n9729), .B(n9730), .Z(n9715) );
  XOR U17836 ( .A(n9726), .B(n9725), .Z(n9730) );
  XOR U17837 ( .A(y[7284]), .B(x[7284]), .Z(n9725) );
  XOR U17838 ( .A(n9728), .B(n9727), .Z(n9726) );
  XOR U17839 ( .A(y[7286]), .B(x[7286]), .Z(n9727) );
  XOR U17840 ( .A(y[7285]), .B(x[7285]), .Z(n9728) );
  XOR U17841 ( .A(n9720), .B(n9719), .Z(n9729) );
  XOR U17842 ( .A(n9722), .B(n9721), .Z(n9719) );
  XOR U17843 ( .A(y[7283]), .B(x[7283]), .Z(n9721) );
  XOR U17844 ( .A(y[7282]), .B(x[7282]), .Z(n9722) );
  XOR U17845 ( .A(y[7281]), .B(x[7281]), .Z(n9720) );
  XNOR U17846 ( .A(n9713), .B(n9712), .Z(n9714) );
  XNOR U17847 ( .A(n9709), .B(n9708), .Z(n9712) );
  XOR U17848 ( .A(n9711), .B(n9710), .Z(n9708) );
  XOR U17849 ( .A(y[7280]), .B(x[7280]), .Z(n9710) );
  XOR U17850 ( .A(y[7279]), .B(x[7279]), .Z(n9711) );
  XOR U17851 ( .A(y[7278]), .B(x[7278]), .Z(n9709) );
  XOR U17852 ( .A(n9703), .B(n9702), .Z(n9713) );
  XOR U17853 ( .A(n9705), .B(n9704), .Z(n9702) );
  XOR U17854 ( .A(y[7277]), .B(x[7277]), .Z(n9704) );
  XOR U17855 ( .A(y[7276]), .B(x[7276]), .Z(n9705) );
  XOR U17856 ( .A(y[7275]), .B(x[7275]), .Z(n9703) );
  XNOR U17857 ( .A(n9679), .B(n9680), .Z(n9697) );
  XNOR U17858 ( .A(n9694), .B(n9695), .Z(n9680) );
  XOR U17859 ( .A(n9691), .B(n9690), .Z(n9695) );
  XOR U17860 ( .A(y[7272]), .B(x[7272]), .Z(n9690) );
  XOR U17861 ( .A(n9693), .B(n9692), .Z(n9691) );
  XOR U17862 ( .A(y[7274]), .B(x[7274]), .Z(n9692) );
  XOR U17863 ( .A(y[7273]), .B(x[7273]), .Z(n9693) );
  XOR U17864 ( .A(n9685), .B(n9684), .Z(n9694) );
  XOR U17865 ( .A(n9687), .B(n9686), .Z(n9684) );
  XOR U17866 ( .A(y[7271]), .B(x[7271]), .Z(n9686) );
  XOR U17867 ( .A(y[7270]), .B(x[7270]), .Z(n9687) );
  XOR U17868 ( .A(y[7269]), .B(x[7269]), .Z(n9685) );
  XNOR U17869 ( .A(n9678), .B(n9677), .Z(n9679) );
  XNOR U17870 ( .A(n9674), .B(n9673), .Z(n9677) );
  XOR U17871 ( .A(n9676), .B(n9675), .Z(n9673) );
  XOR U17872 ( .A(y[7268]), .B(x[7268]), .Z(n9675) );
  XOR U17873 ( .A(y[7267]), .B(x[7267]), .Z(n9676) );
  XOR U17874 ( .A(y[7266]), .B(x[7266]), .Z(n9674) );
  XOR U17875 ( .A(n9668), .B(n9667), .Z(n9678) );
  XOR U17876 ( .A(n9670), .B(n9669), .Z(n9667) );
  XOR U17877 ( .A(y[7265]), .B(x[7265]), .Z(n9669) );
  XOR U17878 ( .A(y[7264]), .B(x[7264]), .Z(n9670) );
  XOR U17879 ( .A(y[7263]), .B(x[7263]), .Z(n9668) );
  NAND U17880 ( .A(n9731), .B(n9732), .Z(N64522) );
  NAND U17881 ( .A(n9733), .B(n9734), .Z(n9732) );
  NANDN U17882 ( .A(n9735), .B(n9736), .Z(n9734) );
  NANDN U17883 ( .A(n9736), .B(n9735), .Z(n9731) );
  XOR U17884 ( .A(n9735), .B(n9737), .Z(N64521) );
  XNOR U17885 ( .A(n9733), .B(n9736), .Z(n9737) );
  NAND U17886 ( .A(n9738), .B(n9739), .Z(n9736) );
  NAND U17887 ( .A(n9740), .B(n9741), .Z(n9739) );
  NANDN U17888 ( .A(n9742), .B(n9743), .Z(n9741) );
  NANDN U17889 ( .A(n9743), .B(n9742), .Z(n9738) );
  AND U17890 ( .A(n9744), .B(n9745), .Z(n9733) );
  NAND U17891 ( .A(n9746), .B(n9747), .Z(n9745) );
  NANDN U17892 ( .A(n9748), .B(n9749), .Z(n9747) );
  NANDN U17893 ( .A(n9749), .B(n9748), .Z(n9744) );
  IV U17894 ( .A(n9750), .Z(n9749) );
  AND U17895 ( .A(n9751), .B(n9752), .Z(n9735) );
  NAND U17896 ( .A(n9753), .B(n9754), .Z(n9752) );
  NANDN U17897 ( .A(n9755), .B(n9756), .Z(n9754) );
  NANDN U17898 ( .A(n9756), .B(n9755), .Z(n9751) );
  XOR U17899 ( .A(n9748), .B(n9757), .Z(N64520) );
  XNOR U17900 ( .A(n9746), .B(n9750), .Z(n9757) );
  XOR U17901 ( .A(n9743), .B(n9758), .Z(n9750) );
  XNOR U17902 ( .A(n9740), .B(n9742), .Z(n9758) );
  AND U17903 ( .A(n9759), .B(n9760), .Z(n9742) );
  NANDN U17904 ( .A(n9761), .B(n9762), .Z(n9760) );
  OR U17905 ( .A(n9763), .B(n9764), .Z(n9762) );
  IV U17906 ( .A(n9765), .Z(n9764) );
  NANDN U17907 ( .A(n9765), .B(n9763), .Z(n9759) );
  AND U17908 ( .A(n9766), .B(n9767), .Z(n9740) );
  NAND U17909 ( .A(n9768), .B(n9769), .Z(n9767) );
  NANDN U17910 ( .A(n9770), .B(n9771), .Z(n9769) );
  NANDN U17911 ( .A(n9771), .B(n9770), .Z(n9766) );
  IV U17912 ( .A(n9772), .Z(n9771) );
  NAND U17913 ( .A(n9773), .B(n9774), .Z(n9743) );
  NANDN U17914 ( .A(n9775), .B(n9776), .Z(n9774) );
  NANDN U17915 ( .A(n9777), .B(n9778), .Z(n9776) );
  NANDN U17916 ( .A(n9778), .B(n9777), .Z(n9773) );
  IV U17917 ( .A(n9779), .Z(n9777) );
  AND U17918 ( .A(n9780), .B(n9781), .Z(n9746) );
  NAND U17919 ( .A(n9782), .B(n9783), .Z(n9781) );
  NANDN U17920 ( .A(n9784), .B(n9785), .Z(n9783) );
  NANDN U17921 ( .A(n9785), .B(n9784), .Z(n9780) );
  XOR U17922 ( .A(n9756), .B(n9786), .Z(n9748) );
  XNOR U17923 ( .A(n9753), .B(n9755), .Z(n9786) );
  AND U17924 ( .A(n9787), .B(n9788), .Z(n9755) );
  NANDN U17925 ( .A(n9789), .B(n9790), .Z(n9788) );
  OR U17926 ( .A(n9791), .B(n9792), .Z(n9790) );
  IV U17927 ( .A(n9793), .Z(n9792) );
  NANDN U17928 ( .A(n9793), .B(n9791), .Z(n9787) );
  AND U17929 ( .A(n9794), .B(n9795), .Z(n9753) );
  NAND U17930 ( .A(n9796), .B(n9797), .Z(n9795) );
  NANDN U17931 ( .A(n9798), .B(n9799), .Z(n9797) );
  NANDN U17932 ( .A(n9799), .B(n9798), .Z(n9794) );
  IV U17933 ( .A(n9800), .Z(n9799) );
  NAND U17934 ( .A(n9801), .B(n9802), .Z(n9756) );
  NANDN U17935 ( .A(n9803), .B(n9804), .Z(n9802) );
  NANDN U17936 ( .A(n9805), .B(n9806), .Z(n9804) );
  NANDN U17937 ( .A(n9806), .B(n9805), .Z(n9801) );
  IV U17938 ( .A(n9807), .Z(n9805) );
  XOR U17939 ( .A(n9782), .B(n9808), .Z(N64519) );
  XNOR U17940 ( .A(n9785), .B(n9784), .Z(n9808) );
  XNOR U17941 ( .A(n9796), .B(n9809), .Z(n9784) );
  XNOR U17942 ( .A(n9800), .B(n9798), .Z(n9809) );
  XOR U17943 ( .A(n9806), .B(n9810), .Z(n9798) );
  XNOR U17944 ( .A(n9803), .B(n9807), .Z(n9810) );
  AND U17945 ( .A(n9811), .B(n9812), .Z(n9807) );
  NAND U17946 ( .A(n9813), .B(n9814), .Z(n9812) );
  NAND U17947 ( .A(n9815), .B(n9816), .Z(n9811) );
  AND U17948 ( .A(n9817), .B(n9818), .Z(n9803) );
  NAND U17949 ( .A(n9819), .B(n9820), .Z(n9818) );
  NAND U17950 ( .A(n9821), .B(n9822), .Z(n9817) );
  NANDN U17951 ( .A(n9823), .B(n9824), .Z(n9806) );
  ANDN U17952 ( .B(n9825), .A(n9826), .Z(n9800) );
  XNOR U17953 ( .A(n9791), .B(n9827), .Z(n9796) );
  XNOR U17954 ( .A(n9789), .B(n9793), .Z(n9827) );
  AND U17955 ( .A(n9828), .B(n9829), .Z(n9793) );
  NAND U17956 ( .A(n9830), .B(n9831), .Z(n9829) );
  NAND U17957 ( .A(n9832), .B(n9833), .Z(n9828) );
  AND U17958 ( .A(n9834), .B(n9835), .Z(n9789) );
  NAND U17959 ( .A(n9836), .B(n9837), .Z(n9835) );
  NAND U17960 ( .A(n9838), .B(n9839), .Z(n9834) );
  AND U17961 ( .A(n9840), .B(n9841), .Z(n9791) );
  NAND U17962 ( .A(n9842), .B(n9843), .Z(n9785) );
  XNOR U17963 ( .A(n9768), .B(n9844), .Z(n9782) );
  XNOR U17964 ( .A(n9772), .B(n9770), .Z(n9844) );
  XOR U17965 ( .A(n9778), .B(n9845), .Z(n9770) );
  XNOR U17966 ( .A(n9775), .B(n9779), .Z(n9845) );
  AND U17967 ( .A(n9846), .B(n9847), .Z(n9779) );
  NAND U17968 ( .A(n9848), .B(n9849), .Z(n9847) );
  NAND U17969 ( .A(n9850), .B(n9851), .Z(n9846) );
  AND U17970 ( .A(n9852), .B(n9853), .Z(n9775) );
  NAND U17971 ( .A(n9854), .B(n9855), .Z(n9853) );
  NAND U17972 ( .A(n9856), .B(n9857), .Z(n9852) );
  NANDN U17973 ( .A(n9858), .B(n9859), .Z(n9778) );
  ANDN U17974 ( .B(n9860), .A(n9861), .Z(n9772) );
  XNOR U17975 ( .A(n9763), .B(n9862), .Z(n9768) );
  XNOR U17976 ( .A(n9761), .B(n9765), .Z(n9862) );
  AND U17977 ( .A(n9863), .B(n9864), .Z(n9765) );
  NAND U17978 ( .A(n9865), .B(n9866), .Z(n9864) );
  NAND U17979 ( .A(n9867), .B(n9868), .Z(n9863) );
  AND U17980 ( .A(n9869), .B(n9870), .Z(n9761) );
  NAND U17981 ( .A(n9871), .B(n9872), .Z(n9870) );
  NAND U17982 ( .A(n9873), .B(n9874), .Z(n9869) );
  AND U17983 ( .A(n9875), .B(n9876), .Z(n9763) );
  XOR U17984 ( .A(n9843), .B(n9842), .Z(N64518) );
  XNOR U17985 ( .A(n9860), .B(n9861), .Z(n9842) );
  XNOR U17986 ( .A(n9875), .B(n9876), .Z(n9861) );
  XOR U17987 ( .A(n9872), .B(n9871), .Z(n9876) );
  XOR U17988 ( .A(y[7260]), .B(x[7260]), .Z(n9871) );
  XOR U17989 ( .A(n9874), .B(n9873), .Z(n9872) );
  XOR U17990 ( .A(y[7262]), .B(x[7262]), .Z(n9873) );
  XOR U17991 ( .A(y[7261]), .B(x[7261]), .Z(n9874) );
  XOR U17992 ( .A(n9866), .B(n9865), .Z(n9875) );
  XOR U17993 ( .A(n9868), .B(n9867), .Z(n9865) );
  XOR U17994 ( .A(y[7259]), .B(x[7259]), .Z(n9867) );
  XOR U17995 ( .A(y[7258]), .B(x[7258]), .Z(n9868) );
  XOR U17996 ( .A(y[7257]), .B(x[7257]), .Z(n9866) );
  XNOR U17997 ( .A(n9859), .B(n9858), .Z(n9860) );
  XNOR U17998 ( .A(n9855), .B(n9854), .Z(n9858) );
  XOR U17999 ( .A(n9857), .B(n9856), .Z(n9854) );
  XOR U18000 ( .A(y[7256]), .B(x[7256]), .Z(n9856) );
  XOR U18001 ( .A(y[7255]), .B(x[7255]), .Z(n9857) );
  XOR U18002 ( .A(y[7254]), .B(x[7254]), .Z(n9855) );
  XOR U18003 ( .A(n9849), .B(n9848), .Z(n9859) );
  XOR U18004 ( .A(n9851), .B(n9850), .Z(n9848) );
  XOR U18005 ( .A(y[7253]), .B(x[7253]), .Z(n9850) );
  XOR U18006 ( .A(y[7252]), .B(x[7252]), .Z(n9851) );
  XOR U18007 ( .A(y[7251]), .B(x[7251]), .Z(n9849) );
  XNOR U18008 ( .A(n9825), .B(n9826), .Z(n9843) );
  XNOR U18009 ( .A(n9840), .B(n9841), .Z(n9826) );
  XOR U18010 ( .A(n9837), .B(n9836), .Z(n9841) );
  XOR U18011 ( .A(y[7248]), .B(x[7248]), .Z(n9836) );
  XOR U18012 ( .A(n9839), .B(n9838), .Z(n9837) );
  XOR U18013 ( .A(y[7250]), .B(x[7250]), .Z(n9838) );
  XOR U18014 ( .A(y[7249]), .B(x[7249]), .Z(n9839) );
  XOR U18015 ( .A(n9831), .B(n9830), .Z(n9840) );
  XOR U18016 ( .A(n9833), .B(n9832), .Z(n9830) );
  XOR U18017 ( .A(y[7247]), .B(x[7247]), .Z(n9832) );
  XOR U18018 ( .A(y[7246]), .B(x[7246]), .Z(n9833) );
  XOR U18019 ( .A(y[7245]), .B(x[7245]), .Z(n9831) );
  XNOR U18020 ( .A(n9824), .B(n9823), .Z(n9825) );
  XNOR U18021 ( .A(n9820), .B(n9819), .Z(n9823) );
  XOR U18022 ( .A(n9822), .B(n9821), .Z(n9819) );
  XOR U18023 ( .A(y[7244]), .B(x[7244]), .Z(n9821) );
  XOR U18024 ( .A(y[7243]), .B(x[7243]), .Z(n9822) );
  XOR U18025 ( .A(y[7242]), .B(x[7242]), .Z(n9820) );
  XOR U18026 ( .A(n9814), .B(n9813), .Z(n9824) );
  XOR U18027 ( .A(n9816), .B(n9815), .Z(n9813) );
  XOR U18028 ( .A(y[7241]), .B(x[7241]), .Z(n9815) );
  XOR U18029 ( .A(y[7240]), .B(x[7240]), .Z(n9816) );
  XOR U18030 ( .A(y[7239]), .B(x[7239]), .Z(n9814) );
  NAND U18031 ( .A(n9877), .B(n9878), .Z(N64509) );
  NAND U18032 ( .A(n9879), .B(n9880), .Z(n9878) );
  NANDN U18033 ( .A(n9881), .B(n9882), .Z(n9880) );
  NANDN U18034 ( .A(n9882), .B(n9881), .Z(n9877) );
  XOR U18035 ( .A(n9881), .B(n9883), .Z(N64508) );
  XNOR U18036 ( .A(n9879), .B(n9882), .Z(n9883) );
  NAND U18037 ( .A(n9884), .B(n9885), .Z(n9882) );
  NAND U18038 ( .A(n9886), .B(n9887), .Z(n9885) );
  NANDN U18039 ( .A(n9888), .B(n9889), .Z(n9887) );
  NANDN U18040 ( .A(n9889), .B(n9888), .Z(n9884) );
  AND U18041 ( .A(n9890), .B(n9891), .Z(n9879) );
  NAND U18042 ( .A(n9892), .B(n9893), .Z(n9891) );
  NANDN U18043 ( .A(n9894), .B(n9895), .Z(n9893) );
  NANDN U18044 ( .A(n9895), .B(n9894), .Z(n9890) );
  IV U18045 ( .A(n9896), .Z(n9895) );
  AND U18046 ( .A(n9897), .B(n9898), .Z(n9881) );
  NAND U18047 ( .A(n9899), .B(n9900), .Z(n9898) );
  NANDN U18048 ( .A(n9901), .B(n9902), .Z(n9900) );
  NANDN U18049 ( .A(n9902), .B(n9901), .Z(n9897) );
  XOR U18050 ( .A(n9894), .B(n9903), .Z(N64507) );
  XNOR U18051 ( .A(n9892), .B(n9896), .Z(n9903) );
  XOR U18052 ( .A(n9889), .B(n9904), .Z(n9896) );
  XNOR U18053 ( .A(n9886), .B(n9888), .Z(n9904) );
  AND U18054 ( .A(n9905), .B(n9906), .Z(n9888) );
  NANDN U18055 ( .A(n9907), .B(n9908), .Z(n9906) );
  OR U18056 ( .A(n9909), .B(n9910), .Z(n9908) );
  IV U18057 ( .A(n9911), .Z(n9910) );
  NANDN U18058 ( .A(n9911), .B(n9909), .Z(n9905) );
  AND U18059 ( .A(n9912), .B(n9913), .Z(n9886) );
  NAND U18060 ( .A(n9914), .B(n9915), .Z(n9913) );
  NANDN U18061 ( .A(n9916), .B(n9917), .Z(n9915) );
  NANDN U18062 ( .A(n9917), .B(n9916), .Z(n9912) );
  IV U18063 ( .A(n9918), .Z(n9917) );
  NAND U18064 ( .A(n9919), .B(n9920), .Z(n9889) );
  NANDN U18065 ( .A(n9921), .B(n9922), .Z(n9920) );
  NANDN U18066 ( .A(n9923), .B(n9924), .Z(n9922) );
  NANDN U18067 ( .A(n9924), .B(n9923), .Z(n9919) );
  IV U18068 ( .A(n9925), .Z(n9923) );
  AND U18069 ( .A(n9926), .B(n9927), .Z(n9892) );
  NAND U18070 ( .A(n9928), .B(n9929), .Z(n9927) );
  NANDN U18071 ( .A(n9930), .B(n9931), .Z(n9929) );
  NANDN U18072 ( .A(n9931), .B(n9930), .Z(n9926) );
  XOR U18073 ( .A(n9902), .B(n9932), .Z(n9894) );
  XNOR U18074 ( .A(n9899), .B(n9901), .Z(n9932) );
  AND U18075 ( .A(n9933), .B(n9934), .Z(n9901) );
  NANDN U18076 ( .A(n9935), .B(n9936), .Z(n9934) );
  OR U18077 ( .A(n9937), .B(n9938), .Z(n9936) );
  IV U18078 ( .A(n9939), .Z(n9938) );
  NANDN U18079 ( .A(n9939), .B(n9937), .Z(n9933) );
  AND U18080 ( .A(n9940), .B(n9941), .Z(n9899) );
  NAND U18081 ( .A(n9942), .B(n9943), .Z(n9941) );
  NANDN U18082 ( .A(n9944), .B(n9945), .Z(n9943) );
  NANDN U18083 ( .A(n9945), .B(n9944), .Z(n9940) );
  IV U18084 ( .A(n9946), .Z(n9945) );
  NAND U18085 ( .A(n9947), .B(n9948), .Z(n9902) );
  NANDN U18086 ( .A(n9949), .B(n9950), .Z(n9948) );
  NANDN U18087 ( .A(n9951), .B(n9952), .Z(n9950) );
  NANDN U18088 ( .A(n9952), .B(n9951), .Z(n9947) );
  IV U18089 ( .A(n9953), .Z(n9951) );
  XOR U18090 ( .A(n9928), .B(n9954), .Z(N64506) );
  XNOR U18091 ( .A(n9931), .B(n9930), .Z(n9954) );
  XNOR U18092 ( .A(n9942), .B(n9955), .Z(n9930) );
  XNOR U18093 ( .A(n9946), .B(n9944), .Z(n9955) );
  XOR U18094 ( .A(n9952), .B(n9956), .Z(n9944) );
  XNOR U18095 ( .A(n9949), .B(n9953), .Z(n9956) );
  AND U18096 ( .A(n9957), .B(n9958), .Z(n9953) );
  NAND U18097 ( .A(n9959), .B(n9960), .Z(n9958) );
  NAND U18098 ( .A(n9961), .B(n9962), .Z(n9957) );
  AND U18099 ( .A(n9963), .B(n9964), .Z(n9949) );
  NAND U18100 ( .A(n9965), .B(n9966), .Z(n9964) );
  NAND U18101 ( .A(n9967), .B(n9968), .Z(n9963) );
  NANDN U18102 ( .A(n9969), .B(n9970), .Z(n9952) );
  ANDN U18103 ( .B(n9971), .A(n9972), .Z(n9946) );
  XNOR U18104 ( .A(n9937), .B(n9973), .Z(n9942) );
  XNOR U18105 ( .A(n9935), .B(n9939), .Z(n9973) );
  AND U18106 ( .A(n9974), .B(n9975), .Z(n9939) );
  NAND U18107 ( .A(n9976), .B(n9977), .Z(n9975) );
  NAND U18108 ( .A(n9978), .B(n9979), .Z(n9974) );
  AND U18109 ( .A(n9980), .B(n9981), .Z(n9935) );
  NAND U18110 ( .A(n9982), .B(n9983), .Z(n9981) );
  NAND U18111 ( .A(n9984), .B(n9985), .Z(n9980) );
  AND U18112 ( .A(n9986), .B(n9987), .Z(n9937) );
  NAND U18113 ( .A(n9988), .B(n9989), .Z(n9931) );
  XNOR U18114 ( .A(n9914), .B(n9990), .Z(n9928) );
  XNOR U18115 ( .A(n9918), .B(n9916), .Z(n9990) );
  XOR U18116 ( .A(n9924), .B(n9991), .Z(n9916) );
  XNOR U18117 ( .A(n9921), .B(n9925), .Z(n9991) );
  AND U18118 ( .A(n9992), .B(n9993), .Z(n9925) );
  NAND U18119 ( .A(n9994), .B(n9995), .Z(n9993) );
  NAND U18120 ( .A(n9996), .B(n9997), .Z(n9992) );
  AND U18121 ( .A(n9998), .B(n9999), .Z(n9921) );
  NAND U18122 ( .A(n10000), .B(n10001), .Z(n9999) );
  NAND U18123 ( .A(n10002), .B(n10003), .Z(n9998) );
  NANDN U18124 ( .A(n10004), .B(n10005), .Z(n9924) );
  ANDN U18125 ( .B(n10006), .A(n10007), .Z(n9918) );
  XNOR U18126 ( .A(n9909), .B(n10008), .Z(n9914) );
  XNOR U18127 ( .A(n9907), .B(n9911), .Z(n10008) );
  AND U18128 ( .A(n10009), .B(n10010), .Z(n9911) );
  NAND U18129 ( .A(n10011), .B(n10012), .Z(n10010) );
  NAND U18130 ( .A(n10013), .B(n10014), .Z(n10009) );
  AND U18131 ( .A(n10015), .B(n10016), .Z(n9907) );
  NAND U18132 ( .A(n10017), .B(n10018), .Z(n10016) );
  NAND U18133 ( .A(n10019), .B(n10020), .Z(n10015) );
  AND U18134 ( .A(n10021), .B(n10022), .Z(n9909) );
  XOR U18135 ( .A(n9989), .B(n9988), .Z(N64505) );
  XNOR U18136 ( .A(n10006), .B(n10007), .Z(n9988) );
  XNOR U18137 ( .A(n10021), .B(n10022), .Z(n10007) );
  XOR U18138 ( .A(n10018), .B(n10017), .Z(n10022) );
  XOR U18139 ( .A(y[7236]), .B(x[7236]), .Z(n10017) );
  XOR U18140 ( .A(n10020), .B(n10019), .Z(n10018) );
  XOR U18141 ( .A(y[7238]), .B(x[7238]), .Z(n10019) );
  XOR U18142 ( .A(y[7237]), .B(x[7237]), .Z(n10020) );
  XOR U18143 ( .A(n10012), .B(n10011), .Z(n10021) );
  XOR U18144 ( .A(n10014), .B(n10013), .Z(n10011) );
  XOR U18145 ( .A(y[7235]), .B(x[7235]), .Z(n10013) );
  XOR U18146 ( .A(y[7234]), .B(x[7234]), .Z(n10014) );
  XOR U18147 ( .A(y[7233]), .B(x[7233]), .Z(n10012) );
  XNOR U18148 ( .A(n10005), .B(n10004), .Z(n10006) );
  XNOR U18149 ( .A(n10001), .B(n10000), .Z(n10004) );
  XOR U18150 ( .A(n10003), .B(n10002), .Z(n10000) );
  XOR U18151 ( .A(y[7232]), .B(x[7232]), .Z(n10002) );
  XOR U18152 ( .A(y[7231]), .B(x[7231]), .Z(n10003) );
  XOR U18153 ( .A(y[7230]), .B(x[7230]), .Z(n10001) );
  XOR U18154 ( .A(n9995), .B(n9994), .Z(n10005) );
  XOR U18155 ( .A(n9997), .B(n9996), .Z(n9994) );
  XOR U18156 ( .A(y[7229]), .B(x[7229]), .Z(n9996) );
  XOR U18157 ( .A(y[7228]), .B(x[7228]), .Z(n9997) );
  XOR U18158 ( .A(y[7227]), .B(x[7227]), .Z(n9995) );
  XNOR U18159 ( .A(n9971), .B(n9972), .Z(n9989) );
  XNOR U18160 ( .A(n9986), .B(n9987), .Z(n9972) );
  XOR U18161 ( .A(n9983), .B(n9982), .Z(n9987) );
  XOR U18162 ( .A(y[7224]), .B(x[7224]), .Z(n9982) );
  XOR U18163 ( .A(n9985), .B(n9984), .Z(n9983) );
  XOR U18164 ( .A(y[7226]), .B(x[7226]), .Z(n9984) );
  XOR U18165 ( .A(y[7225]), .B(x[7225]), .Z(n9985) );
  XOR U18166 ( .A(n9977), .B(n9976), .Z(n9986) );
  XOR U18167 ( .A(n9979), .B(n9978), .Z(n9976) );
  XOR U18168 ( .A(y[7223]), .B(x[7223]), .Z(n9978) );
  XOR U18169 ( .A(y[7222]), .B(x[7222]), .Z(n9979) );
  XOR U18170 ( .A(y[7221]), .B(x[7221]), .Z(n9977) );
  XNOR U18171 ( .A(n9970), .B(n9969), .Z(n9971) );
  XNOR U18172 ( .A(n9966), .B(n9965), .Z(n9969) );
  XOR U18173 ( .A(n9968), .B(n9967), .Z(n9965) );
  XOR U18174 ( .A(y[7220]), .B(x[7220]), .Z(n9967) );
  XOR U18175 ( .A(y[7219]), .B(x[7219]), .Z(n9968) );
  XOR U18176 ( .A(y[7218]), .B(x[7218]), .Z(n9966) );
  XOR U18177 ( .A(n9960), .B(n9959), .Z(n9970) );
  XOR U18178 ( .A(n9962), .B(n9961), .Z(n9959) );
  XOR U18179 ( .A(y[7217]), .B(x[7217]), .Z(n9961) );
  XOR U18180 ( .A(y[7216]), .B(x[7216]), .Z(n9962) );
  XOR U18181 ( .A(y[7215]), .B(x[7215]), .Z(n9960) );
  NAND U18182 ( .A(n10023), .B(n10024), .Z(N64496) );
  NAND U18183 ( .A(n10025), .B(n10026), .Z(n10024) );
  NANDN U18184 ( .A(n10027), .B(n10028), .Z(n10026) );
  NANDN U18185 ( .A(n10028), .B(n10027), .Z(n10023) );
  XOR U18186 ( .A(n10027), .B(n10029), .Z(N64495) );
  XNOR U18187 ( .A(n10025), .B(n10028), .Z(n10029) );
  NAND U18188 ( .A(n10030), .B(n10031), .Z(n10028) );
  NAND U18189 ( .A(n10032), .B(n10033), .Z(n10031) );
  NANDN U18190 ( .A(n10034), .B(n10035), .Z(n10033) );
  NANDN U18191 ( .A(n10035), .B(n10034), .Z(n10030) );
  AND U18192 ( .A(n10036), .B(n10037), .Z(n10025) );
  NAND U18193 ( .A(n10038), .B(n10039), .Z(n10037) );
  NANDN U18194 ( .A(n10040), .B(n10041), .Z(n10039) );
  NANDN U18195 ( .A(n10041), .B(n10040), .Z(n10036) );
  IV U18196 ( .A(n10042), .Z(n10041) );
  AND U18197 ( .A(n10043), .B(n10044), .Z(n10027) );
  NAND U18198 ( .A(n10045), .B(n10046), .Z(n10044) );
  NANDN U18199 ( .A(n10047), .B(n10048), .Z(n10046) );
  NANDN U18200 ( .A(n10048), .B(n10047), .Z(n10043) );
  XOR U18201 ( .A(n10040), .B(n10049), .Z(N64494) );
  XNOR U18202 ( .A(n10038), .B(n10042), .Z(n10049) );
  XOR U18203 ( .A(n10035), .B(n10050), .Z(n10042) );
  XNOR U18204 ( .A(n10032), .B(n10034), .Z(n10050) );
  AND U18205 ( .A(n10051), .B(n10052), .Z(n10034) );
  NANDN U18206 ( .A(n10053), .B(n10054), .Z(n10052) );
  OR U18207 ( .A(n10055), .B(n10056), .Z(n10054) );
  IV U18208 ( .A(n10057), .Z(n10056) );
  NANDN U18209 ( .A(n10057), .B(n10055), .Z(n10051) );
  AND U18210 ( .A(n10058), .B(n10059), .Z(n10032) );
  NAND U18211 ( .A(n10060), .B(n10061), .Z(n10059) );
  NANDN U18212 ( .A(n10062), .B(n10063), .Z(n10061) );
  NANDN U18213 ( .A(n10063), .B(n10062), .Z(n10058) );
  IV U18214 ( .A(n10064), .Z(n10063) );
  NAND U18215 ( .A(n10065), .B(n10066), .Z(n10035) );
  NANDN U18216 ( .A(n10067), .B(n10068), .Z(n10066) );
  NANDN U18217 ( .A(n10069), .B(n10070), .Z(n10068) );
  NANDN U18218 ( .A(n10070), .B(n10069), .Z(n10065) );
  IV U18219 ( .A(n10071), .Z(n10069) );
  AND U18220 ( .A(n10072), .B(n10073), .Z(n10038) );
  NAND U18221 ( .A(n10074), .B(n10075), .Z(n10073) );
  NANDN U18222 ( .A(n10076), .B(n10077), .Z(n10075) );
  NANDN U18223 ( .A(n10077), .B(n10076), .Z(n10072) );
  XOR U18224 ( .A(n10048), .B(n10078), .Z(n10040) );
  XNOR U18225 ( .A(n10045), .B(n10047), .Z(n10078) );
  AND U18226 ( .A(n10079), .B(n10080), .Z(n10047) );
  NANDN U18227 ( .A(n10081), .B(n10082), .Z(n10080) );
  OR U18228 ( .A(n10083), .B(n10084), .Z(n10082) );
  IV U18229 ( .A(n10085), .Z(n10084) );
  NANDN U18230 ( .A(n10085), .B(n10083), .Z(n10079) );
  AND U18231 ( .A(n10086), .B(n10087), .Z(n10045) );
  NAND U18232 ( .A(n10088), .B(n10089), .Z(n10087) );
  NANDN U18233 ( .A(n10090), .B(n10091), .Z(n10089) );
  NANDN U18234 ( .A(n10091), .B(n10090), .Z(n10086) );
  IV U18235 ( .A(n10092), .Z(n10091) );
  NAND U18236 ( .A(n10093), .B(n10094), .Z(n10048) );
  NANDN U18237 ( .A(n10095), .B(n10096), .Z(n10094) );
  NANDN U18238 ( .A(n10097), .B(n10098), .Z(n10096) );
  NANDN U18239 ( .A(n10098), .B(n10097), .Z(n10093) );
  IV U18240 ( .A(n10099), .Z(n10097) );
  XOR U18241 ( .A(n10074), .B(n10100), .Z(N64493) );
  XNOR U18242 ( .A(n10077), .B(n10076), .Z(n10100) );
  XNOR U18243 ( .A(n10088), .B(n10101), .Z(n10076) );
  XNOR U18244 ( .A(n10092), .B(n10090), .Z(n10101) );
  XOR U18245 ( .A(n10098), .B(n10102), .Z(n10090) );
  XNOR U18246 ( .A(n10095), .B(n10099), .Z(n10102) );
  AND U18247 ( .A(n10103), .B(n10104), .Z(n10099) );
  NAND U18248 ( .A(n10105), .B(n10106), .Z(n10104) );
  NAND U18249 ( .A(n10107), .B(n10108), .Z(n10103) );
  AND U18250 ( .A(n10109), .B(n10110), .Z(n10095) );
  NAND U18251 ( .A(n10111), .B(n10112), .Z(n10110) );
  NAND U18252 ( .A(n10113), .B(n10114), .Z(n10109) );
  NANDN U18253 ( .A(n10115), .B(n10116), .Z(n10098) );
  ANDN U18254 ( .B(n10117), .A(n10118), .Z(n10092) );
  XNOR U18255 ( .A(n10083), .B(n10119), .Z(n10088) );
  XNOR U18256 ( .A(n10081), .B(n10085), .Z(n10119) );
  AND U18257 ( .A(n10120), .B(n10121), .Z(n10085) );
  NAND U18258 ( .A(n10122), .B(n10123), .Z(n10121) );
  NAND U18259 ( .A(n10124), .B(n10125), .Z(n10120) );
  AND U18260 ( .A(n10126), .B(n10127), .Z(n10081) );
  NAND U18261 ( .A(n10128), .B(n10129), .Z(n10127) );
  NAND U18262 ( .A(n10130), .B(n10131), .Z(n10126) );
  AND U18263 ( .A(n10132), .B(n10133), .Z(n10083) );
  NAND U18264 ( .A(n10134), .B(n10135), .Z(n10077) );
  XNOR U18265 ( .A(n10060), .B(n10136), .Z(n10074) );
  XNOR U18266 ( .A(n10064), .B(n10062), .Z(n10136) );
  XOR U18267 ( .A(n10070), .B(n10137), .Z(n10062) );
  XNOR U18268 ( .A(n10067), .B(n10071), .Z(n10137) );
  AND U18269 ( .A(n10138), .B(n10139), .Z(n10071) );
  NAND U18270 ( .A(n10140), .B(n10141), .Z(n10139) );
  NAND U18271 ( .A(n10142), .B(n10143), .Z(n10138) );
  AND U18272 ( .A(n10144), .B(n10145), .Z(n10067) );
  NAND U18273 ( .A(n10146), .B(n10147), .Z(n10145) );
  NAND U18274 ( .A(n10148), .B(n10149), .Z(n10144) );
  NANDN U18275 ( .A(n10150), .B(n10151), .Z(n10070) );
  ANDN U18276 ( .B(n10152), .A(n10153), .Z(n10064) );
  XNOR U18277 ( .A(n10055), .B(n10154), .Z(n10060) );
  XNOR U18278 ( .A(n10053), .B(n10057), .Z(n10154) );
  AND U18279 ( .A(n10155), .B(n10156), .Z(n10057) );
  NAND U18280 ( .A(n10157), .B(n10158), .Z(n10156) );
  NAND U18281 ( .A(n10159), .B(n10160), .Z(n10155) );
  AND U18282 ( .A(n10161), .B(n10162), .Z(n10053) );
  NAND U18283 ( .A(n10163), .B(n10164), .Z(n10162) );
  NAND U18284 ( .A(n10165), .B(n10166), .Z(n10161) );
  AND U18285 ( .A(n10167), .B(n10168), .Z(n10055) );
  XOR U18286 ( .A(n10135), .B(n10134), .Z(N64492) );
  XNOR U18287 ( .A(n10152), .B(n10153), .Z(n10134) );
  XNOR U18288 ( .A(n10167), .B(n10168), .Z(n10153) );
  XOR U18289 ( .A(n10164), .B(n10163), .Z(n10168) );
  XOR U18290 ( .A(y[7212]), .B(x[7212]), .Z(n10163) );
  XOR U18291 ( .A(n10166), .B(n10165), .Z(n10164) );
  XOR U18292 ( .A(y[7214]), .B(x[7214]), .Z(n10165) );
  XOR U18293 ( .A(y[7213]), .B(x[7213]), .Z(n10166) );
  XOR U18294 ( .A(n10158), .B(n10157), .Z(n10167) );
  XOR U18295 ( .A(n10160), .B(n10159), .Z(n10157) );
  XOR U18296 ( .A(y[7211]), .B(x[7211]), .Z(n10159) );
  XOR U18297 ( .A(y[7210]), .B(x[7210]), .Z(n10160) );
  XOR U18298 ( .A(y[7209]), .B(x[7209]), .Z(n10158) );
  XNOR U18299 ( .A(n10151), .B(n10150), .Z(n10152) );
  XNOR U18300 ( .A(n10147), .B(n10146), .Z(n10150) );
  XOR U18301 ( .A(n10149), .B(n10148), .Z(n10146) );
  XOR U18302 ( .A(y[7208]), .B(x[7208]), .Z(n10148) );
  XOR U18303 ( .A(y[7207]), .B(x[7207]), .Z(n10149) );
  XOR U18304 ( .A(y[7206]), .B(x[7206]), .Z(n10147) );
  XOR U18305 ( .A(n10141), .B(n10140), .Z(n10151) );
  XOR U18306 ( .A(n10143), .B(n10142), .Z(n10140) );
  XOR U18307 ( .A(y[7205]), .B(x[7205]), .Z(n10142) );
  XOR U18308 ( .A(y[7204]), .B(x[7204]), .Z(n10143) );
  XOR U18309 ( .A(y[7203]), .B(x[7203]), .Z(n10141) );
  XNOR U18310 ( .A(n10117), .B(n10118), .Z(n10135) );
  XNOR U18311 ( .A(n10132), .B(n10133), .Z(n10118) );
  XOR U18312 ( .A(n10129), .B(n10128), .Z(n10133) );
  XOR U18313 ( .A(y[7200]), .B(x[7200]), .Z(n10128) );
  XOR U18314 ( .A(n10131), .B(n10130), .Z(n10129) );
  XOR U18315 ( .A(y[7202]), .B(x[7202]), .Z(n10130) );
  XOR U18316 ( .A(y[7201]), .B(x[7201]), .Z(n10131) );
  XOR U18317 ( .A(n10123), .B(n10122), .Z(n10132) );
  XOR U18318 ( .A(n10125), .B(n10124), .Z(n10122) );
  XOR U18319 ( .A(y[7199]), .B(x[7199]), .Z(n10124) );
  XOR U18320 ( .A(y[7198]), .B(x[7198]), .Z(n10125) );
  XOR U18321 ( .A(y[7197]), .B(x[7197]), .Z(n10123) );
  XNOR U18322 ( .A(n10116), .B(n10115), .Z(n10117) );
  XNOR U18323 ( .A(n10112), .B(n10111), .Z(n10115) );
  XOR U18324 ( .A(n10114), .B(n10113), .Z(n10111) );
  XOR U18325 ( .A(y[7196]), .B(x[7196]), .Z(n10113) );
  XOR U18326 ( .A(y[7195]), .B(x[7195]), .Z(n10114) );
  XOR U18327 ( .A(y[7194]), .B(x[7194]), .Z(n10112) );
  XOR U18328 ( .A(n10106), .B(n10105), .Z(n10116) );
  XOR U18329 ( .A(n10108), .B(n10107), .Z(n10105) );
  XOR U18330 ( .A(y[7193]), .B(x[7193]), .Z(n10107) );
  XOR U18331 ( .A(y[7192]), .B(x[7192]), .Z(n10108) );
  XOR U18332 ( .A(y[7191]), .B(x[7191]), .Z(n10106) );
  NAND U18333 ( .A(n10169), .B(n10170), .Z(N64483) );
  NAND U18334 ( .A(n10171), .B(n10172), .Z(n10170) );
  NANDN U18335 ( .A(n10173), .B(n10174), .Z(n10172) );
  NANDN U18336 ( .A(n10174), .B(n10173), .Z(n10169) );
  XOR U18337 ( .A(n10173), .B(n10175), .Z(N64482) );
  XNOR U18338 ( .A(n10171), .B(n10174), .Z(n10175) );
  NAND U18339 ( .A(n10176), .B(n10177), .Z(n10174) );
  NAND U18340 ( .A(n10178), .B(n10179), .Z(n10177) );
  NANDN U18341 ( .A(n10180), .B(n10181), .Z(n10179) );
  NANDN U18342 ( .A(n10181), .B(n10180), .Z(n10176) );
  AND U18343 ( .A(n10182), .B(n10183), .Z(n10171) );
  NAND U18344 ( .A(n10184), .B(n10185), .Z(n10183) );
  NANDN U18345 ( .A(n10186), .B(n10187), .Z(n10185) );
  NANDN U18346 ( .A(n10187), .B(n10186), .Z(n10182) );
  IV U18347 ( .A(n10188), .Z(n10187) );
  AND U18348 ( .A(n10189), .B(n10190), .Z(n10173) );
  NAND U18349 ( .A(n10191), .B(n10192), .Z(n10190) );
  NANDN U18350 ( .A(n10193), .B(n10194), .Z(n10192) );
  NANDN U18351 ( .A(n10194), .B(n10193), .Z(n10189) );
  XOR U18352 ( .A(n10186), .B(n10195), .Z(N64481) );
  XNOR U18353 ( .A(n10184), .B(n10188), .Z(n10195) );
  XOR U18354 ( .A(n10181), .B(n10196), .Z(n10188) );
  XNOR U18355 ( .A(n10178), .B(n10180), .Z(n10196) );
  AND U18356 ( .A(n10197), .B(n10198), .Z(n10180) );
  NANDN U18357 ( .A(n10199), .B(n10200), .Z(n10198) );
  OR U18358 ( .A(n10201), .B(n10202), .Z(n10200) );
  IV U18359 ( .A(n10203), .Z(n10202) );
  NANDN U18360 ( .A(n10203), .B(n10201), .Z(n10197) );
  AND U18361 ( .A(n10204), .B(n10205), .Z(n10178) );
  NAND U18362 ( .A(n10206), .B(n10207), .Z(n10205) );
  NANDN U18363 ( .A(n10208), .B(n10209), .Z(n10207) );
  NANDN U18364 ( .A(n10209), .B(n10208), .Z(n10204) );
  IV U18365 ( .A(n10210), .Z(n10209) );
  NAND U18366 ( .A(n10211), .B(n10212), .Z(n10181) );
  NANDN U18367 ( .A(n10213), .B(n10214), .Z(n10212) );
  NANDN U18368 ( .A(n10215), .B(n10216), .Z(n10214) );
  NANDN U18369 ( .A(n10216), .B(n10215), .Z(n10211) );
  IV U18370 ( .A(n10217), .Z(n10215) );
  AND U18371 ( .A(n10218), .B(n10219), .Z(n10184) );
  NAND U18372 ( .A(n10220), .B(n10221), .Z(n10219) );
  NANDN U18373 ( .A(n10222), .B(n10223), .Z(n10221) );
  NANDN U18374 ( .A(n10223), .B(n10222), .Z(n10218) );
  XOR U18375 ( .A(n10194), .B(n10224), .Z(n10186) );
  XNOR U18376 ( .A(n10191), .B(n10193), .Z(n10224) );
  AND U18377 ( .A(n10225), .B(n10226), .Z(n10193) );
  NANDN U18378 ( .A(n10227), .B(n10228), .Z(n10226) );
  OR U18379 ( .A(n10229), .B(n10230), .Z(n10228) );
  IV U18380 ( .A(n10231), .Z(n10230) );
  NANDN U18381 ( .A(n10231), .B(n10229), .Z(n10225) );
  AND U18382 ( .A(n10232), .B(n10233), .Z(n10191) );
  NAND U18383 ( .A(n10234), .B(n10235), .Z(n10233) );
  NANDN U18384 ( .A(n10236), .B(n10237), .Z(n10235) );
  NANDN U18385 ( .A(n10237), .B(n10236), .Z(n10232) );
  IV U18386 ( .A(n10238), .Z(n10237) );
  NAND U18387 ( .A(n10239), .B(n10240), .Z(n10194) );
  NANDN U18388 ( .A(n10241), .B(n10242), .Z(n10240) );
  NANDN U18389 ( .A(n10243), .B(n10244), .Z(n10242) );
  NANDN U18390 ( .A(n10244), .B(n10243), .Z(n10239) );
  IV U18391 ( .A(n10245), .Z(n10243) );
  XOR U18392 ( .A(n10220), .B(n10246), .Z(N64480) );
  XNOR U18393 ( .A(n10223), .B(n10222), .Z(n10246) );
  XNOR U18394 ( .A(n10234), .B(n10247), .Z(n10222) );
  XNOR U18395 ( .A(n10238), .B(n10236), .Z(n10247) );
  XOR U18396 ( .A(n10244), .B(n10248), .Z(n10236) );
  XNOR U18397 ( .A(n10241), .B(n10245), .Z(n10248) );
  AND U18398 ( .A(n10249), .B(n10250), .Z(n10245) );
  NAND U18399 ( .A(n10251), .B(n10252), .Z(n10250) );
  NAND U18400 ( .A(n10253), .B(n10254), .Z(n10249) );
  AND U18401 ( .A(n10255), .B(n10256), .Z(n10241) );
  NAND U18402 ( .A(n10257), .B(n10258), .Z(n10256) );
  NAND U18403 ( .A(n10259), .B(n10260), .Z(n10255) );
  NANDN U18404 ( .A(n10261), .B(n10262), .Z(n10244) );
  ANDN U18405 ( .B(n10263), .A(n10264), .Z(n10238) );
  XNOR U18406 ( .A(n10229), .B(n10265), .Z(n10234) );
  XNOR U18407 ( .A(n10227), .B(n10231), .Z(n10265) );
  AND U18408 ( .A(n10266), .B(n10267), .Z(n10231) );
  NAND U18409 ( .A(n10268), .B(n10269), .Z(n10267) );
  NAND U18410 ( .A(n10270), .B(n10271), .Z(n10266) );
  AND U18411 ( .A(n10272), .B(n10273), .Z(n10227) );
  NAND U18412 ( .A(n10274), .B(n10275), .Z(n10273) );
  NAND U18413 ( .A(n10276), .B(n10277), .Z(n10272) );
  AND U18414 ( .A(n10278), .B(n10279), .Z(n10229) );
  NAND U18415 ( .A(n10280), .B(n10281), .Z(n10223) );
  XNOR U18416 ( .A(n10206), .B(n10282), .Z(n10220) );
  XNOR U18417 ( .A(n10210), .B(n10208), .Z(n10282) );
  XOR U18418 ( .A(n10216), .B(n10283), .Z(n10208) );
  XNOR U18419 ( .A(n10213), .B(n10217), .Z(n10283) );
  AND U18420 ( .A(n10284), .B(n10285), .Z(n10217) );
  NAND U18421 ( .A(n10286), .B(n10287), .Z(n10285) );
  NAND U18422 ( .A(n10288), .B(n10289), .Z(n10284) );
  AND U18423 ( .A(n10290), .B(n10291), .Z(n10213) );
  NAND U18424 ( .A(n10292), .B(n10293), .Z(n10291) );
  NAND U18425 ( .A(n10294), .B(n10295), .Z(n10290) );
  NANDN U18426 ( .A(n10296), .B(n10297), .Z(n10216) );
  ANDN U18427 ( .B(n10298), .A(n10299), .Z(n10210) );
  XNOR U18428 ( .A(n10201), .B(n10300), .Z(n10206) );
  XNOR U18429 ( .A(n10199), .B(n10203), .Z(n10300) );
  AND U18430 ( .A(n10301), .B(n10302), .Z(n10203) );
  NAND U18431 ( .A(n10303), .B(n10304), .Z(n10302) );
  NAND U18432 ( .A(n10305), .B(n10306), .Z(n10301) );
  AND U18433 ( .A(n10307), .B(n10308), .Z(n10199) );
  NAND U18434 ( .A(n10309), .B(n10310), .Z(n10308) );
  NAND U18435 ( .A(n10311), .B(n10312), .Z(n10307) );
  AND U18436 ( .A(n10313), .B(n10314), .Z(n10201) );
  XOR U18437 ( .A(n10281), .B(n10280), .Z(N64479) );
  XNOR U18438 ( .A(n10298), .B(n10299), .Z(n10280) );
  XNOR U18439 ( .A(n10313), .B(n10314), .Z(n10299) );
  XOR U18440 ( .A(n10310), .B(n10309), .Z(n10314) );
  XOR U18441 ( .A(y[7188]), .B(x[7188]), .Z(n10309) );
  XOR U18442 ( .A(n10312), .B(n10311), .Z(n10310) );
  XOR U18443 ( .A(y[7190]), .B(x[7190]), .Z(n10311) );
  XOR U18444 ( .A(y[7189]), .B(x[7189]), .Z(n10312) );
  XOR U18445 ( .A(n10304), .B(n10303), .Z(n10313) );
  XOR U18446 ( .A(n10306), .B(n10305), .Z(n10303) );
  XOR U18447 ( .A(y[7187]), .B(x[7187]), .Z(n10305) );
  XOR U18448 ( .A(y[7186]), .B(x[7186]), .Z(n10306) );
  XOR U18449 ( .A(y[7185]), .B(x[7185]), .Z(n10304) );
  XNOR U18450 ( .A(n10297), .B(n10296), .Z(n10298) );
  XNOR U18451 ( .A(n10293), .B(n10292), .Z(n10296) );
  XOR U18452 ( .A(n10295), .B(n10294), .Z(n10292) );
  XOR U18453 ( .A(y[7184]), .B(x[7184]), .Z(n10294) );
  XOR U18454 ( .A(y[7183]), .B(x[7183]), .Z(n10295) );
  XOR U18455 ( .A(y[7182]), .B(x[7182]), .Z(n10293) );
  XOR U18456 ( .A(n10287), .B(n10286), .Z(n10297) );
  XOR U18457 ( .A(n10289), .B(n10288), .Z(n10286) );
  XOR U18458 ( .A(y[7181]), .B(x[7181]), .Z(n10288) );
  XOR U18459 ( .A(y[7180]), .B(x[7180]), .Z(n10289) );
  XOR U18460 ( .A(y[7179]), .B(x[7179]), .Z(n10287) );
  XNOR U18461 ( .A(n10263), .B(n10264), .Z(n10281) );
  XNOR U18462 ( .A(n10278), .B(n10279), .Z(n10264) );
  XOR U18463 ( .A(n10275), .B(n10274), .Z(n10279) );
  XOR U18464 ( .A(y[7176]), .B(x[7176]), .Z(n10274) );
  XOR U18465 ( .A(n10277), .B(n10276), .Z(n10275) );
  XOR U18466 ( .A(y[7178]), .B(x[7178]), .Z(n10276) );
  XOR U18467 ( .A(y[7177]), .B(x[7177]), .Z(n10277) );
  XOR U18468 ( .A(n10269), .B(n10268), .Z(n10278) );
  XOR U18469 ( .A(n10271), .B(n10270), .Z(n10268) );
  XOR U18470 ( .A(y[7175]), .B(x[7175]), .Z(n10270) );
  XOR U18471 ( .A(y[7174]), .B(x[7174]), .Z(n10271) );
  XOR U18472 ( .A(y[7173]), .B(x[7173]), .Z(n10269) );
  XNOR U18473 ( .A(n10262), .B(n10261), .Z(n10263) );
  XNOR U18474 ( .A(n10258), .B(n10257), .Z(n10261) );
  XOR U18475 ( .A(n10260), .B(n10259), .Z(n10257) );
  XOR U18476 ( .A(y[7172]), .B(x[7172]), .Z(n10259) );
  XOR U18477 ( .A(y[7171]), .B(x[7171]), .Z(n10260) );
  XOR U18478 ( .A(y[7170]), .B(x[7170]), .Z(n10258) );
  XOR U18479 ( .A(n10252), .B(n10251), .Z(n10262) );
  XOR U18480 ( .A(n10254), .B(n10253), .Z(n10251) );
  XOR U18481 ( .A(y[7169]), .B(x[7169]), .Z(n10253) );
  XOR U18482 ( .A(y[7168]), .B(x[7168]), .Z(n10254) );
  XOR U18483 ( .A(y[7167]), .B(x[7167]), .Z(n10252) );
  NAND U18484 ( .A(n10315), .B(n10316), .Z(N64470) );
  NAND U18485 ( .A(n10317), .B(n10318), .Z(n10316) );
  NANDN U18486 ( .A(n10319), .B(n10320), .Z(n10318) );
  NANDN U18487 ( .A(n10320), .B(n10319), .Z(n10315) );
  XOR U18488 ( .A(n10319), .B(n10321), .Z(N64469) );
  XNOR U18489 ( .A(n10317), .B(n10320), .Z(n10321) );
  NAND U18490 ( .A(n10322), .B(n10323), .Z(n10320) );
  NAND U18491 ( .A(n10324), .B(n10325), .Z(n10323) );
  NANDN U18492 ( .A(n10326), .B(n10327), .Z(n10325) );
  NANDN U18493 ( .A(n10327), .B(n10326), .Z(n10322) );
  AND U18494 ( .A(n10328), .B(n10329), .Z(n10317) );
  NAND U18495 ( .A(n10330), .B(n10331), .Z(n10329) );
  NANDN U18496 ( .A(n10332), .B(n10333), .Z(n10331) );
  NANDN U18497 ( .A(n10333), .B(n10332), .Z(n10328) );
  IV U18498 ( .A(n10334), .Z(n10333) );
  AND U18499 ( .A(n10335), .B(n10336), .Z(n10319) );
  NAND U18500 ( .A(n10337), .B(n10338), .Z(n10336) );
  NANDN U18501 ( .A(n10339), .B(n10340), .Z(n10338) );
  NANDN U18502 ( .A(n10340), .B(n10339), .Z(n10335) );
  XOR U18503 ( .A(n10332), .B(n10341), .Z(N64468) );
  XNOR U18504 ( .A(n10330), .B(n10334), .Z(n10341) );
  XOR U18505 ( .A(n10327), .B(n10342), .Z(n10334) );
  XNOR U18506 ( .A(n10324), .B(n10326), .Z(n10342) );
  AND U18507 ( .A(n10343), .B(n10344), .Z(n10326) );
  NANDN U18508 ( .A(n10345), .B(n10346), .Z(n10344) );
  OR U18509 ( .A(n10347), .B(n10348), .Z(n10346) );
  IV U18510 ( .A(n10349), .Z(n10348) );
  NANDN U18511 ( .A(n10349), .B(n10347), .Z(n10343) );
  AND U18512 ( .A(n10350), .B(n10351), .Z(n10324) );
  NAND U18513 ( .A(n10352), .B(n10353), .Z(n10351) );
  NANDN U18514 ( .A(n10354), .B(n10355), .Z(n10353) );
  NANDN U18515 ( .A(n10355), .B(n10354), .Z(n10350) );
  IV U18516 ( .A(n10356), .Z(n10355) );
  NAND U18517 ( .A(n10357), .B(n10358), .Z(n10327) );
  NANDN U18518 ( .A(n10359), .B(n10360), .Z(n10358) );
  NANDN U18519 ( .A(n10361), .B(n10362), .Z(n10360) );
  NANDN U18520 ( .A(n10362), .B(n10361), .Z(n10357) );
  IV U18521 ( .A(n10363), .Z(n10361) );
  AND U18522 ( .A(n10364), .B(n10365), .Z(n10330) );
  NAND U18523 ( .A(n10366), .B(n10367), .Z(n10365) );
  NANDN U18524 ( .A(n10368), .B(n10369), .Z(n10367) );
  NANDN U18525 ( .A(n10369), .B(n10368), .Z(n10364) );
  XOR U18526 ( .A(n10340), .B(n10370), .Z(n10332) );
  XNOR U18527 ( .A(n10337), .B(n10339), .Z(n10370) );
  AND U18528 ( .A(n10371), .B(n10372), .Z(n10339) );
  NANDN U18529 ( .A(n10373), .B(n10374), .Z(n10372) );
  OR U18530 ( .A(n10375), .B(n10376), .Z(n10374) );
  IV U18531 ( .A(n10377), .Z(n10376) );
  NANDN U18532 ( .A(n10377), .B(n10375), .Z(n10371) );
  AND U18533 ( .A(n10378), .B(n10379), .Z(n10337) );
  NAND U18534 ( .A(n10380), .B(n10381), .Z(n10379) );
  NANDN U18535 ( .A(n10382), .B(n10383), .Z(n10381) );
  NANDN U18536 ( .A(n10383), .B(n10382), .Z(n10378) );
  IV U18537 ( .A(n10384), .Z(n10383) );
  NAND U18538 ( .A(n10385), .B(n10386), .Z(n10340) );
  NANDN U18539 ( .A(n10387), .B(n10388), .Z(n10386) );
  NANDN U18540 ( .A(n10389), .B(n10390), .Z(n10388) );
  NANDN U18541 ( .A(n10390), .B(n10389), .Z(n10385) );
  IV U18542 ( .A(n10391), .Z(n10389) );
  XOR U18543 ( .A(n10366), .B(n10392), .Z(N64467) );
  XNOR U18544 ( .A(n10369), .B(n10368), .Z(n10392) );
  XNOR U18545 ( .A(n10380), .B(n10393), .Z(n10368) );
  XNOR U18546 ( .A(n10384), .B(n10382), .Z(n10393) );
  XOR U18547 ( .A(n10390), .B(n10394), .Z(n10382) );
  XNOR U18548 ( .A(n10387), .B(n10391), .Z(n10394) );
  AND U18549 ( .A(n10395), .B(n10396), .Z(n10391) );
  NAND U18550 ( .A(n10397), .B(n10398), .Z(n10396) );
  NAND U18551 ( .A(n10399), .B(n10400), .Z(n10395) );
  AND U18552 ( .A(n10401), .B(n10402), .Z(n10387) );
  NAND U18553 ( .A(n10403), .B(n10404), .Z(n10402) );
  NAND U18554 ( .A(n10405), .B(n10406), .Z(n10401) );
  NANDN U18555 ( .A(n10407), .B(n10408), .Z(n10390) );
  ANDN U18556 ( .B(n10409), .A(n10410), .Z(n10384) );
  XNOR U18557 ( .A(n10375), .B(n10411), .Z(n10380) );
  XNOR U18558 ( .A(n10373), .B(n10377), .Z(n10411) );
  AND U18559 ( .A(n10412), .B(n10413), .Z(n10377) );
  NAND U18560 ( .A(n10414), .B(n10415), .Z(n10413) );
  NAND U18561 ( .A(n10416), .B(n10417), .Z(n10412) );
  AND U18562 ( .A(n10418), .B(n10419), .Z(n10373) );
  NAND U18563 ( .A(n10420), .B(n10421), .Z(n10419) );
  NAND U18564 ( .A(n10422), .B(n10423), .Z(n10418) );
  AND U18565 ( .A(n10424), .B(n10425), .Z(n10375) );
  NAND U18566 ( .A(n10426), .B(n10427), .Z(n10369) );
  XNOR U18567 ( .A(n10352), .B(n10428), .Z(n10366) );
  XNOR U18568 ( .A(n10356), .B(n10354), .Z(n10428) );
  XOR U18569 ( .A(n10362), .B(n10429), .Z(n10354) );
  XNOR U18570 ( .A(n10359), .B(n10363), .Z(n10429) );
  AND U18571 ( .A(n10430), .B(n10431), .Z(n10363) );
  NAND U18572 ( .A(n10432), .B(n10433), .Z(n10431) );
  NAND U18573 ( .A(n10434), .B(n10435), .Z(n10430) );
  AND U18574 ( .A(n10436), .B(n10437), .Z(n10359) );
  NAND U18575 ( .A(n10438), .B(n10439), .Z(n10437) );
  NAND U18576 ( .A(n10440), .B(n10441), .Z(n10436) );
  NANDN U18577 ( .A(n10442), .B(n10443), .Z(n10362) );
  ANDN U18578 ( .B(n10444), .A(n10445), .Z(n10356) );
  XNOR U18579 ( .A(n10347), .B(n10446), .Z(n10352) );
  XNOR U18580 ( .A(n10345), .B(n10349), .Z(n10446) );
  AND U18581 ( .A(n10447), .B(n10448), .Z(n10349) );
  NAND U18582 ( .A(n10449), .B(n10450), .Z(n10448) );
  NAND U18583 ( .A(n10451), .B(n10452), .Z(n10447) );
  AND U18584 ( .A(n10453), .B(n10454), .Z(n10345) );
  NAND U18585 ( .A(n10455), .B(n10456), .Z(n10454) );
  NAND U18586 ( .A(n10457), .B(n10458), .Z(n10453) );
  AND U18587 ( .A(n10459), .B(n10460), .Z(n10347) );
  XOR U18588 ( .A(n10427), .B(n10426), .Z(N64466) );
  XNOR U18589 ( .A(n10444), .B(n10445), .Z(n10426) );
  XNOR U18590 ( .A(n10459), .B(n10460), .Z(n10445) );
  XOR U18591 ( .A(n10456), .B(n10455), .Z(n10460) );
  XOR U18592 ( .A(y[7164]), .B(x[7164]), .Z(n10455) );
  XOR U18593 ( .A(n10458), .B(n10457), .Z(n10456) );
  XOR U18594 ( .A(y[7166]), .B(x[7166]), .Z(n10457) );
  XOR U18595 ( .A(y[7165]), .B(x[7165]), .Z(n10458) );
  XOR U18596 ( .A(n10450), .B(n10449), .Z(n10459) );
  XOR U18597 ( .A(n10452), .B(n10451), .Z(n10449) );
  XOR U18598 ( .A(y[7163]), .B(x[7163]), .Z(n10451) );
  XOR U18599 ( .A(y[7162]), .B(x[7162]), .Z(n10452) );
  XOR U18600 ( .A(y[7161]), .B(x[7161]), .Z(n10450) );
  XNOR U18601 ( .A(n10443), .B(n10442), .Z(n10444) );
  XNOR U18602 ( .A(n10439), .B(n10438), .Z(n10442) );
  XOR U18603 ( .A(n10441), .B(n10440), .Z(n10438) );
  XOR U18604 ( .A(y[7160]), .B(x[7160]), .Z(n10440) );
  XOR U18605 ( .A(y[7159]), .B(x[7159]), .Z(n10441) );
  XOR U18606 ( .A(y[7158]), .B(x[7158]), .Z(n10439) );
  XOR U18607 ( .A(n10433), .B(n10432), .Z(n10443) );
  XOR U18608 ( .A(n10435), .B(n10434), .Z(n10432) );
  XOR U18609 ( .A(y[7157]), .B(x[7157]), .Z(n10434) );
  XOR U18610 ( .A(y[7156]), .B(x[7156]), .Z(n10435) );
  XOR U18611 ( .A(y[7155]), .B(x[7155]), .Z(n10433) );
  XNOR U18612 ( .A(n10409), .B(n10410), .Z(n10427) );
  XNOR U18613 ( .A(n10424), .B(n10425), .Z(n10410) );
  XOR U18614 ( .A(n10421), .B(n10420), .Z(n10425) );
  XOR U18615 ( .A(y[7152]), .B(x[7152]), .Z(n10420) );
  XOR U18616 ( .A(n10423), .B(n10422), .Z(n10421) );
  XOR U18617 ( .A(y[7154]), .B(x[7154]), .Z(n10422) );
  XOR U18618 ( .A(y[7153]), .B(x[7153]), .Z(n10423) );
  XOR U18619 ( .A(n10415), .B(n10414), .Z(n10424) );
  XOR U18620 ( .A(n10417), .B(n10416), .Z(n10414) );
  XOR U18621 ( .A(y[7151]), .B(x[7151]), .Z(n10416) );
  XOR U18622 ( .A(y[7150]), .B(x[7150]), .Z(n10417) );
  XOR U18623 ( .A(y[7149]), .B(x[7149]), .Z(n10415) );
  XNOR U18624 ( .A(n10408), .B(n10407), .Z(n10409) );
  XNOR U18625 ( .A(n10404), .B(n10403), .Z(n10407) );
  XOR U18626 ( .A(n10406), .B(n10405), .Z(n10403) );
  XOR U18627 ( .A(y[7148]), .B(x[7148]), .Z(n10405) );
  XOR U18628 ( .A(y[7147]), .B(x[7147]), .Z(n10406) );
  XOR U18629 ( .A(y[7146]), .B(x[7146]), .Z(n10404) );
  XOR U18630 ( .A(n10398), .B(n10397), .Z(n10408) );
  XOR U18631 ( .A(n10400), .B(n10399), .Z(n10397) );
  XOR U18632 ( .A(y[7145]), .B(x[7145]), .Z(n10399) );
  XOR U18633 ( .A(y[7144]), .B(x[7144]), .Z(n10400) );
  XOR U18634 ( .A(y[7143]), .B(x[7143]), .Z(n10398) );
  NAND U18635 ( .A(n10461), .B(n10462), .Z(N64457) );
  NAND U18636 ( .A(n10463), .B(n10464), .Z(n10462) );
  NANDN U18637 ( .A(n10465), .B(n10466), .Z(n10464) );
  NANDN U18638 ( .A(n10466), .B(n10465), .Z(n10461) );
  XOR U18639 ( .A(n10465), .B(n10467), .Z(N64456) );
  XNOR U18640 ( .A(n10463), .B(n10466), .Z(n10467) );
  NAND U18641 ( .A(n10468), .B(n10469), .Z(n10466) );
  NAND U18642 ( .A(n10470), .B(n10471), .Z(n10469) );
  NANDN U18643 ( .A(n10472), .B(n10473), .Z(n10471) );
  NANDN U18644 ( .A(n10473), .B(n10472), .Z(n10468) );
  AND U18645 ( .A(n10474), .B(n10475), .Z(n10463) );
  NAND U18646 ( .A(n10476), .B(n10477), .Z(n10475) );
  NANDN U18647 ( .A(n10478), .B(n10479), .Z(n10477) );
  NANDN U18648 ( .A(n10479), .B(n10478), .Z(n10474) );
  IV U18649 ( .A(n10480), .Z(n10479) );
  AND U18650 ( .A(n10481), .B(n10482), .Z(n10465) );
  NAND U18651 ( .A(n10483), .B(n10484), .Z(n10482) );
  NANDN U18652 ( .A(n10485), .B(n10486), .Z(n10484) );
  NANDN U18653 ( .A(n10486), .B(n10485), .Z(n10481) );
  XOR U18654 ( .A(n10478), .B(n10487), .Z(N64455) );
  XNOR U18655 ( .A(n10476), .B(n10480), .Z(n10487) );
  XOR U18656 ( .A(n10473), .B(n10488), .Z(n10480) );
  XNOR U18657 ( .A(n10470), .B(n10472), .Z(n10488) );
  AND U18658 ( .A(n10489), .B(n10490), .Z(n10472) );
  NANDN U18659 ( .A(n10491), .B(n10492), .Z(n10490) );
  OR U18660 ( .A(n10493), .B(n10494), .Z(n10492) );
  IV U18661 ( .A(n10495), .Z(n10494) );
  NANDN U18662 ( .A(n10495), .B(n10493), .Z(n10489) );
  AND U18663 ( .A(n10496), .B(n10497), .Z(n10470) );
  NAND U18664 ( .A(n10498), .B(n10499), .Z(n10497) );
  NANDN U18665 ( .A(n10500), .B(n10501), .Z(n10499) );
  NANDN U18666 ( .A(n10501), .B(n10500), .Z(n10496) );
  IV U18667 ( .A(n10502), .Z(n10501) );
  NAND U18668 ( .A(n10503), .B(n10504), .Z(n10473) );
  NANDN U18669 ( .A(n10505), .B(n10506), .Z(n10504) );
  NANDN U18670 ( .A(n10507), .B(n10508), .Z(n10506) );
  NANDN U18671 ( .A(n10508), .B(n10507), .Z(n10503) );
  IV U18672 ( .A(n10509), .Z(n10507) );
  AND U18673 ( .A(n10510), .B(n10511), .Z(n10476) );
  NAND U18674 ( .A(n10512), .B(n10513), .Z(n10511) );
  NANDN U18675 ( .A(n10514), .B(n10515), .Z(n10513) );
  NANDN U18676 ( .A(n10515), .B(n10514), .Z(n10510) );
  XOR U18677 ( .A(n10486), .B(n10516), .Z(n10478) );
  XNOR U18678 ( .A(n10483), .B(n10485), .Z(n10516) );
  AND U18679 ( .A(n10517), .B(n10518), .Z(n10485) );
  NANDN U18680 ( .A(n10519), .B(n10520), .Z(n10518) );
  OR U18681 ( .A(n10521), .B(n10522), .Z(n10520) );
  IV U18682 ( .A(n10523), .Z(n10522) );
  NANDN U18683 ( .A(n10523), .B(n10521), .Z(n10517) );
  AND U18684 ( .A(n10524), .B(n10525), .Z(n10483) );
  NAND U18685 ( .A(n10526), .B(n10527), .Z(n10525) );
  NANDN U18686 ( .A(n10528), .B(n10529), .Z(n10527) );
  NANDN U18687 ( .A(n10529), .B(n10528), .Z(n10524) );
  IV U18688 ( .A(n10530), .Z(n10529) );
  NAND U18689 ( .A(n10531), .B(n10532), .Z(n10486) );
  NANDN U18690 ( .A(n10533), .B(n10534), .Z(n10532) );
  NANDN U18691 ( .A(n10535), .B(n10536), .Z(n10534) );
  NANDN U18692 ( .A(n10536), .B(n10535), .Z(n10531) );
  IV U18693 ( .A(n10537), .Z(n10535) );
  XOR U18694 ( .A(n10512), .B(n10538), .Z(N64454) );
  XNOR U18695 ( .A(n10515), .B(n10514), .Z(n10538) );
  XNOR U18696 ( .A(n10526), .B(n10539), .Z(n10514) );
  XNOR U18697 ( .A(n10530), .B(n10528), .Z(n10539) );
  XOR U18698 ( .A(n10536), .B(n10540), .Z(n10528) );
  XNOR U18699 ( .A(n10533), .B(n10537), .Z(n10540) );
  AND U18700 ( .A(n10541), .B(n10542), .Z(n10537) );
  NAND U18701 ( .A(n10543), .B(n10544), .Z(n10542) );
  NAND U18702 ( .A(n10545), .B(n10546), .Z(n10541) );
  AND U18703 ( .A(n10547), .B(n10548), .Z(n10533) );
  NAND U18704 ( .A(n10549), .B(n10550), .Z(n10548) );
  NAND U18705 ( .A(n10551), .B(n10552), .Z(n10547) );
  NANDN U18706 ( .A(n10553), .B(n10554), .Z(n10536) );
  ANDN U18707 ( .B(n10555), .A(n10556), .Z(n10530) );
  XNOR U18708 ( .A(n10521), .B(n10557), .Z(n10526) );
  XNOR U18709 ( .A(n10519), .B(n10523), .Z(n10557) );
  AND U18710 ( .A(n10558), .B(n10559), .Z(n10523) );
  NAND U18711 ( .A(n10560), .B(n10561), .Z(n10559) );
  NAND U18712 ( .A(n10562), .B(n10563), .Z(n10558) );
  AND U18713 ( .A(n10564), .B(n10565), .Z(n10519) );
  NAND U18714 ( .A(n10566), .B(n10567), .Z(n10565) );
  NAND U18715 ( .A(n10568), .B(n10569), .Z(n10564) );
  AND U18716 ( .A(n10570), .B(n10571), .Z(n10521) );
  NAND U18717 ( .A(n10572), .B(n10573), .Z(n10515) );
  XNOR U18718 ( .A(n10498), .B(n10574), .Z(n10512) );
  XNOR U18719 ( .A(n10502), .B(n10500), .Z(n10574) );
  XOR U18720 ( .A(n10508), .B(n10575), .Z(n10500) );
  XNOR U18721 ( .A(n10505), .B(n10509), .Z(n10575) );
  AND U18722 ( .A(n10576), .B(n10577), .Z(n10509) );
  NAND U18723 ( .A(n10578), .B(n10579), .Z(n10577) );
  NAND U18724 ( .A(n10580), .B(n10581), .Z(n10576) );
  AND U18725 ( .A(n10582), .B(n10583), .Z(n10505) );
  NAND U18726 ( .A(n10584), .B(n10585), .Z(n10583) );
  NAND U18727 ( .A(n10586), .B(n10587), .Z(n10582) );
  NANDN U18728 ( .A(n10588), .B(n10589), .Z(n10508) );
  ANDN U18729 ( .B(n10590), .A(n10591), .Z(n10502) );
  XNOR U18730 ( .A(n10493), .B(n10592), .Z(n10498) );
  XNOR U18731 ( .A(n10491), .B(n10495), .Z(n10592) );
  AND U18732 ( .A(n10593), .B(n10594), .Z(n10495) );
  NAND U18733 ( .A(n10595), .B(n10596), .Z(n10594) );
  NAND U18734 ( .A(n10597), .B(n10598), .Z(n10593) );
  AND U18735 ( .A(n10599), .B(n10600), .Z(n10491) );
  NAND U18736 ( .A(n10601), .B(n10602), .Z(n10600) );
  NAND U18737 ( .A(n10603), .B(n10604), .Z(n10599) );
  AND U18738 ( .A(n10605), .B(n10606), .Z(n10493) );
  XOR U18739 ( .A(n10573), .B(n10572), .Z(N64453) );
  XNOR U18740 ( .A(n10590), .B(n10591), .Z(n10572) );
  XNOR U18741 ( .A(n10605), .B(n10606), .Z(n10591) );
  XOR U18742 ( .A(n10602), .B(n10601), .Z(n10606) );
  XOR U18743 ( .A(y[7140]), .B(x[7140]), .Z(n10601) );
  XOR U18744 ( .A(n10604), .B(n10603), .Z(n10602) );
  XOR U18745 ( .A(y[7142]), .B(x[7142]), .Z(n10603) );
  XOR U18746 ( .A(y[7141]), .B(x[7141]), .Z(n10604) );
  XOR U18747 ( .A(n10596), .B(n10595), .Z(n10605) );
  XOR U18748 ( .A(n10598), .B(n10597), .Z(n10595) );
  XOR U18749 ( .A(y[7139]), .B(x[7139]), .Z(n10597) );
  XOR U18750 ( .A(y[7138]), .B(x[7138]), .Z(n10598) );
  XOR U18751 ( .A(y[7137]), .B(x[7137]), .Z(n10596) );
  XNOR U18752 ( .A(n10589), .B(n10588), .Z(n10590) );
  XNOR U18753 ( .A(n10585), .B(n10584), .Z(n10588) );
  XOR U18754 ( .A(n10587), .B(n10586), .Z(n10584) );
  XOR U18755 ( .A(y[7136]), .B(x[7136]), .Z(n10586) );
  XOR U18756 ( .A(y[7135]), .B(x[7135]), .Z(n10587) );
  XOR U18757 ( .A(y[7134]), .B(x[7134]), .Z(n10585) );
  XOR U18758 ( .A(n10579), .B(n10578), .Z(n10589) );
  XOR U18759 ( .A(n10581), .B(n10580), .Z(n10578) );
  XOR U18760 ( .A(y[7133]), .B(x[7133]), .Z(n10580) );
  XOR U18761 ( .A(y[7132]), .B(x[7132]), .Z(n10581) );
  XOR U18762 ( .A(y[7131]), .B(x[7131]), .Z(n10579) );
  XNOR U18763 ( .A(n10555), .B(n10556), .Z(n10573) );
  XNOR U18764 ( .A(n10570), .B(n10571), .Z(n10556) );
  XOR U18765 ( .A(n10567), .B(n10566), .Z(n10571) );
  XOR U18766 ( .A(y[7128]), .B(x[7128]), .Z(n10566) );
  XOR U18767 ( .A(n10569), .B(n10568), .Z(n10567) );
  XOR U18768 ( .A(y[7130]), .B(x[7130]), .Z(n10568) );
  XOR U18769 ( .A(y[7129]), .B(x[7129]), .Z(n10569) );
  XOR U18770 ( .A(n10561), .B(n10560), .Z(n10570) );
  XOR U18771 ( .A(n10563), .B(n10562), .Z(n10560) );
  XOR U18772 ( .A(y[7127]), .B(x[7127]), .Z(n10562) );
  XOR U18773 ( .A(y[7126]), .B(x[7126]), .Z(n10563) );
  XOR U18774 ( .A(y[7125]), .B(x[7125]), .Z(n10561) );
  XNOR U18775 ( .A(n10554), .B(n10553), .Z(n10555) );
  XNOR U18776 ( .A(n10550), .B(n10549), .Z(n10553) );
  XOR U18777 ( .A(n10552), .B(n10551), .Z(n10549) );
  XOR U18778 ( .A(y[7124]), .B(x[7124]), .Z(n10551) );
  XOR U18779 ( .A(y[7123]), .B(x[7123]), .Z(n10552) );
  XOR U18780 ( .A(y[7122]), .B(x[7122]), .Z(n10550) );
  XOR U18781 ( .A(n10544), .B(n10543), .Z(n10554) );
  XOR U18782 ( .A(n10546), .B(n10545), .Z(n10543) );
  XOR U18783 ( .A(y[7121]), .B(x[7121]), .Z(n10545) );
  XOR U18784 ( .A(y[7120]), .B(x[7120]), .Z(n10546) );
  XOR U18785 ( .A(y[7119]), .B(x[7119]), .Z(n10544) );
  NAND U18786 ( .A(n10607), .B(n10608), .Z(N64444) );
  NAND U18787 ( .A(n10609), .B(n10610), .Z(n10608) );
  NANDN U18788 ( .A(n10611), .B(n10612), .Z(n10610) );
  NANDN U18789 ( .A(n10612), .B(n10611), .Z(n10607) );
  XOR U18790 ( .A(n10611), .B(n10613), .Z(N64443) );
  XNOR U18791 ( .A(n10609), .B(n10612), .Z(n10613) );
  NAND U18792 ( .A(n10614), .B(n10615), .Z(n10612) );
  NAND U18793 ( .A(n10616), .B(n10617), .Z(n10615) );
  NANDN U18794 ( .A(n10618), .B(n10619), .Z(n10617) );
  NANDN U18795 ( .A(n10619), .B(n10618), .Z(n10614) );
  AND U18796 ( .A(n10620), .B(n10621), .Z(n10609) );
  NAND U18797 ( .A(n10622), .B(n10623), .Z(n10621) );
  NANDN U18798 ( .A(n10624), .B(n10625), .Z(n10623) );
  NANDN U18799 ( .A(n10625), .B(n10624), .Z(n10620) );
  IV U18800 ( .A(n10626), .Z(n10625) );
  AND U18801 ( .A(n10627), .B(n10628), .Z(n10611) );
  NAND U18802 ( .A(n10629), .B(n10630), .Z(n10628) );
  NANDN U18803 ( .A(n10631), .B(n10632), .Z(n10630) );
  NANDN U18804 ( .A(n10632), .B(n10631), .Z(n10627) );
  XOR U18805 ( .A(n10624), .B(n10633), .Z(N64442) );
  XNOR U18806 ( .A(n10622), .B(n10626), .Z(n10633) );
  XOR U18807 ( .A(n10619), .B(n10634), .Z(n10626) );
  XNOR U18808 ( .A(n10616), .B(n10618), .Z(n10634) );
  AND U18809 ( .A(n10635), .B(n10636), .Z(n10618) );
  NANDN U18810 ( .A(n10637), .B(n10638), .Z(n10636) );
  OR U18811 ( .A(n10639), .B(n10640), .Z(n10638) );
  IV U18812 ( .A(n10641), .Z(n10640) );
  NANDN U18813 ( .A(n10641), .B(n10639), .Z(n10635) );
  AND U18814 ( .A(n10642), .B(n10643), .Z(n10616) );
  NAND U18815 ( .A(n10644), .B(n10645), .Z(n10643) );
  NANDN U18816 ( .A(n10646), .B(n10647), .Z(n10645) );
  NANDN U18817 ( .A(n10647), .B(n10646), .Z(n10642) );
  IV U18818 ( .A(n10648), .Z(n10647) );
  NAND U18819 ( .A(n10649), .B(n10650), .Z(n10619) );
  NANDN U18820 ( .A(n10651), .B(n10652), .Z(n10650) );
  NANDN U18821 ( .A(n10653), .B(n10654), .Z(n10652) );
  NANDN U18822 ( .A(n10654), .B(n10653), .Z(n10649) );
  IV U18823 ( .A(n10655), .Z(n10653) );
  AND U18824 ( .A(n10656), .B(n10657), .Z(n10622) );
  NAND U18825 ( .A(n10658), .B(n10659), .Z(n10657) );
  NANDN U18826 ( .A(n10660), .B(n10661), .Z(n10659) );
  NANDN U18827 ( .A(n10661), .B(n10660), .Z(n10656) );
  XOR U18828 ( .A(n10632), .B(n10662), .Z(n10624) );
  XNOR U18829 ( .A(n10629), .B(n10631), .Z(n10662) );
  AND U18830 ( .A(n10663), .B(n10664), .Z(n10631) );
  NANDN U18831 ( .A(n10665), .B(n10666), .Z(n10664) );
  OR U18832 ( .A(n10667), .B(n10668), .Z(n10666) );
  IV U18833 ( .A(n10669), .Z(n10668) );
  NANDN U18834 ( .A(n10669), .B(n10667), .Z(n10663) );
  AND U18835 ( .A(n10670), .B(n10671), .Z(n10629) );
  NAND U18836 ( .A(n10672), .B(n10673), .Z(n10671) );
  NANDN U18837 ( .A(n10674), .B(n10675), .Z(n10673) );
  NANDN U18838 ( .A(n10675), .B(n10674), .Z(n10670) );
  IV U18839 ( .A(n10676), .Z(n10675) );
  NAND U18840 ( .A(n10677), .B(n10678), .Z(n10632) );
  NANDN U18841 ( .A(n10679), .B(n10680), .Z(n10678) );
  NANDN U18842 ( .A(n10681), .B(n10682), .Z(n10680) );
  NANDN U18843 ( .A(n10682), .B(n10681), .Z(n10677) );
  IV U18844 ( .A(n10683), .Z(n10681) );
  XOR U18845 ( .A(n10658), .B(n10684), .Z(N64441) );
  XNOR U18846 ( .A(n10661), .B(n10660), .Z(n10684) );
  XNOR U18847 ( .A(n10672), .B(n10685), .Z(n10660) );
  XNOR U18848 ( .A(n10676), .B(n10674), .Z(n10685) );
  XOR U18849 ( .A(n10682), .B(n10686), .Z(n10674) );
  XNOR U18850 ( .A(n10679), .B(n10683), .Z(n10686) );
  AND U18851 ( .A(n10687), .B(n10688), .Z(n10683) );
  NAND U18852 ( .A(n10689), .B(n10690), .Z(n10688) );
  NAND U18853 ( .A(n10691), .B(n10692), .Z(n10687) );
  AND U18854 ( .A(n10693), .B(n10694), .Z(n10679) );
  NAND U18855 ( .A(n10695), .B(n10696), .Z(n10694) );
  NAND U18856 ( .A(n10697), .B(n10698), .Z(n10693) );
  NANDN U18857 ( .A(n10699), .B(n10700), .Z(n10682) );
  ANDN U18858 ( .B(n10701), .A(n10702), .Z(n10676) );
  XNOR U18859 ( .A(n10667), .B(n10703), .Z(n10672) );
  XNOR U18860 ( .A(n10665), .B(n10669), .Z(n10703) );
  AND U18861 ( .A(n10704), .B(n10705), .Z(n10669) );
  NAND U18862 ( .A(n10706), .B(n10707), .Z(n10705) );
  NAND U18863 ( .A(n10708), .B(n10709), .Z(n10704) );
  AND U18864 ( .A(n10710), .B(n10711), .Z(n10665) );
  NAND U18865 ( .A(n10712), .B(n10713), .Z(n10711) );
  NAND U18866 ( .A(n10714), .B(n10715), .Z(n10710) );
  AND U18867 ( .A(n10716), .B(n10717), .Z(n10667) );
  NAND U18868 ( .A(n10718), .B(n10719), .Z(n10661) );
  XNOR U18869 ( .A(n10644), .B(n10720), .Z(n10658) );
  XNOR U18870 ( .A(n10648), .B(n10646), .Z(n10720) );
  XOR U18871 ( .A(n10654), .B(n10721), .Z(n10646) );
  XNOR U18872 ( .A(n10651), .B(n10655), .Z(n10721) );
  AND U18873 ( .A(n10722), .B(n10723), .Z(n10655) );
  NAND U18874 ( .A(n10724), .B(n10725), .Z(n10723) );
  NAND U18875 ( .A(n10726), .B(n10727), .Z(n10722) );
  AND U18876 ( .A(n10728), .B(n10729), .Z(n10651) );
  NAND U18877 ( .A(n10730), .B(n10731), .Z(n10729) );
  NAND U18878 ( .A(n10732), .B(n10733), .Z(n10728) );
  NANDN U18879 ( .A(n10734), .B(n10735), .Z(n10654) );
  ANDN U18880 ( .B(n10736), .A(n10737), .Z(n10648) );
  XNOR U18881 ( .A(n10639), .B(n10738), .Z(n10644) );
  XNOR U18882 ( .A(n10637), .B(n10641), .Z(n10738) );
  AND U18883 ( .A(n10739), .B(n10740), .Z(n10641) );
  NAND U18884 ( .A(n10741), .B(n10742), .Z(n10740) );
  NAND U18885 ( .A(n10743), .B(n10744), .Z(n10739) );
  AND U18886 ( .A(n10745), .B(n10746), .Z(n10637) );
  NAND U18887 ( .A(n10747), .B(n10748), .Z(n10746) );
  NAND U18888 ( .A(n10749), .B(n10750), .Z(n10745) );
  AND U18889 ( .A(n10751), .B(n10752), .Z(n10639) );
  XOR U18890 ( .A(n10719), .B(n10718), .Z(N64440) );
  XNOR U18891 ( .A(n10736), .B(n10737), .Z(n10718) );
  XNOR U18892 ( .A(n10751), .B(n10752), .Z(n10737) );
  XOR U18893 ( .A(n10748), .B(n10747), .Z(n10752) );
  XOR U18894 ( .A(y[7116]), .B(x[7116]), .Z(n10747) );
  XOR U18895 ( .A(n10750), .B(n10749), .Z(n10748) );
  XOR U18896 ( .A(y[7118]), .B(x[7118]), .Z(n10749) );
  XOR U18897 ( .A(y[7117]), .B(x[7117]), .Z(n10750) );
  XOR U18898 ( .A(n10742), .B(n10741), .Z(n10751) );
  XOR U18899 ( .A(n10744), .B(n10743), .Z(n10741) );
  XOR U18900 ( .A(y[7115]), .B(x[7115]), .Z(n10743) );
  XOR U18901 ( .A(y[7114]), .B(x[7114]), .Z(n10744) );
  XOR U18902 ( .A(y[7113]), .B(x[7113]), .Z(n10742) );
  XNOR U18903 ( .A(n10735), .B(n10734), .Z(n10736) );
  XNOR U18904 ( .A(n10731), .B(n10730), .Z(n10734) );
  XOR U18905 ( .A(n10733), .B(n10732), .Z(n10730) );
  XOR U18906 ( .A(y[7112]), .B(x[7112]), .Z(n10732) );
  XOR U18907 ( .A(y[7111]), .B(x[7111]), .Z(n10733) );
  XOR U18908 ( .A(y[7110]), .B(x[7110]), .Z(n10731) );
  XOR U18909 ( .A(n10725), .B(n10724), .Z(n10735) );
  XOR U18910 ( .A(n10727), .B(n10726), .Z(n10724) );
  XOR U18911 ( .A(y[7109]), .B(x[7109]), .Z(n10726) );
  XOR U18912 ( .A(y[7108]), .B(x[7108]), .Z(n10727) );
  XOR U18913 ( .A(y[7107]), .B(x[7107]), .Z(n10725) );
  XNOR U18914 ( .A(n10701), .B(n10702), .Z(n10719) );
  XNOR U18915 ( .A(n10716), .B(n10717), .Z(n10702) );
  XOR U18916 ( .A(n10713), .B(n10712), .Z(n10717) );
  XOR U18917 ( .A(y[7104]), .B(x[7104]), .Z(n10712) );
  XOR U18918 ( .A(n10715), .B(n10714), .Z(n10713) );
  XOR U18919 ( .A(y[7106]), .B(x[7106]), .Z(n10714) );
  XOR U18920 ( .A(y[7105]), .B(x[7105]), .Z(n10715) );
  XOR U18921 ( .A(n10707), .B(n10706), .Z(n10716) );
  XOR U18922 ( .A(n10709), .B(n10708), .Z(n10706) );
  XOR U18923 ( .A(y[7103]), .B(x[7103]), .Z(n10708) );
  XOR U18924 ( .A(y[7102]), .B(x[7102]), .Z(n10709) );
  XOR U18925 ( .A(y[7101]), .B(x[7101]), .Z(n10707) );
  XNOR U18926 ( .A(n10700), .B(n10699), .Z(n10701) );
  XNOR U18927 ( .A(n10696), .B(n10695), .Z(n10699) );
  XOR U18928 ( .A(n10698), .B(n10697), .Z(n10695) );
  XOR U18929 ( .A(y[7100]), .B(x[7100]), .Z(n10697) );
  XOR U18930 ( .A(y[7099]), .B(x[7099]), .Z(n10698) );
  XOR U18931 ( .A(y[7098]), .B(x[7098]), .Z(n10696) );
  XOR U18932 ( .A(n10690), .B(n10689), .Z(n10700) );
  XOR U18933 ( .A(n10692), .B(n10691), .Z(n10689) );
  XOR U18934 ( .A(y[7097]), .B(x[7097]), .Z(n10691) );
  XOR U18935 ( .A(y[7096]), .B(x[7096]), .Z(n10692) );
  XOR U18936 ( .A(y[7095]), .B(x[7095]), .Z(n10690) );
  NAND U18937 ( .A(n10753), .B(n10754), .Z(N64431) );
  NAND U18938 ( .A(n10755), .B(n10756), .Z(n10754) );
  NANDN U18939 ( .A(n10757), .B(n10758), .Z(n10756) );
  NANDN U18940 ( .A(n10758), .B(n10757), .Z(n10753) );
  XOR U18941 ( .A(n10757), .B(n10759), .Z(N64430) );
  XNOR U18942 ( .A(n10755), .B(n10758), .Z(n10759) );
  NAND U18943 ( .A(n10760), .B(n10761), .Z(n10758) );
  NAND U18944 ( .A(n10762), .B(n10763), .Z(n10761) );
  NANDN U18945 ( .A(n10764), .B(n10765), .Z(n10763) );
  NANDN U18946 ( .A(n10765), .B(n10764), .Z(n10760) );
  AND U18947 ( .A(n10766), .B(n10767), .Z(n10755) );
  NAND U18948 ( .A(n10768), .B(n10769), .Z(n10767) );
  NANDN U18949 ( .A(n10770), .B(n10771), .Z(n10769) );
  NANDN U18950 ( .A(n10771), .B(n10770), .Z(n10766) );
  IV U18951 ( .A(n10772), .Z(n10771) );
  AND U18952 ( .A(n10773), .B(n10774), .Z(n10757) );
  NAND U18953 ( .A(n10775), .B(n10776), .Z(n10774) );
  NANDN U18954 ( .A(n10777), .B(n10778), .Z(n10776) );
  NANDN U18955 ( .A(n10778), .B(n10777), .Z(n10773) );
  XOR U18956 ( .A(n10770), .B(n10779), .Z(N64429) );
  XNOR U18957 ( .A(n10768), .B(n10772), .Z(n10779) );
  XOR U18958 ( .A(n10765), .B(n10780), .Z(n10772) );
  XNOR U18959 ( .A(n10762), .B(n10764), .Z(n10780) );
  AND U18960 ( .A(n10781), .B(n10782), .Z(n10764) );
  NANDN U18961 ( .A(n10783), .B(n10784), .Z(n10782) );
  OR U18962 ( .A(n10785), .B(n10786), .Z(n10784) );
  IV U18963 ( .A(n10787), .Z(n10786) );
  NANDN U18964 ( .A(n10787), .B(n10785), .Z(n10781) );
  AND U18965 ( .A(n10788), .B(n10789), .Z(n10762) );
  NAND U18966 ( .A(n10790), .B(n10791), .Z(n10789) );
  NANDN U18967 ( .A(n10792), .B(n10793), .Z(n10791) );
  NANDN U18968 ( .A(n10793), .B(n10792), .Z(n10788) );
  IV U18969 ( .A(n10794), .Z(n10793) );
  NAND U18970 ( .A(n10795), .B(n10796), .Z(n10765) );
  NANDN U18971 ( .A(n10797), .B(n10798), .Z(n10796) );
  NANDN U18972 ( .A(n10799), .B(n10800), .Z(n10798) );
  NANDN U18973 ( .A(n10800), .B(n10799), .Z(n10795) );
  IV U18974 ( .A(n10801), .Z(n10799) );
  AND U18975 ( .A(n10802), .B(n10803), .Z(n10768) );
  NAND U18976 ( .A(n10804), .B(n10805), .Z(n10803) );
  NANDN U18977 ( .A(n10806), .B(n10807), .Z(n10805) );
  NANDN U18978 ( .A(n10807), .B(n10806), .Z(n10802) );
  XOR U18979 ( .A(n10778), .B(n10808), .Z(n10770) );
  XNOR U18980 ( .A(n10775), .B(n10777), .Z(n10808) );
  AND U18981 ( .A(n10809), .B(n10810), .Z(n10777) );
  NANDN U18982 ( .A(n10811), .B(n10812), .Z(n10810) );
  OR U18983 ( .A(n10813), .B(n10814), .Z(n10812) );
  IV U18984 ( .A(n10815), .Z(n10814) );
  NANDN U18985 ( .A(n10815), .B(n10813), .Z(n10809) );
  AND U18986 ( .A(n10816), .B(n10817), .Z(n10775) );
  NAND U18987 ( .A(n10818), .B(n10819), .Z(n10817) );
  NANDN U18988 ( .A(n10820), .B(n10821), .Z(n10819) );
  NANDN U18989 ( .A(n10821), .B(n10820), .Z(n10816) );
  IV U18990 ( .A(n10822), .Z(n10821) );
  NAND U18991 ( .A(n10823), .B(n10824), .Z(n10778) );
  NANDN U18992 ( .A(n10825), .B(n10826), .Z(n10824) );
  NANDN U18993 ( .A(n10827), .B(n10828), .Z(n10826) );
  NANDN U18994 ( .A(n10828), .B(n10827), .Z(n10823) );
  IV U18995 ( .A(n10829), .Z(n10827) );
  XOR U18996 ( .A(n10804), .B(n10830), .Z(N64428) );
  XNOR U18997 ( .A(n10807), .B(n10806), .Z(n10830) );
  XNOR U18998 ( .A(n10818), .B(n10831), .Z(n10806) );
  XNOR U18999 ( .A(n10822), .B(n10820), .Z(n10831) );
  XOR U19000 ( .A(n10828), .B(n10832), .Z(n10820) );
  XNOR U19001 ( .A(n10825), .B(n10829), .Z(n10832) );
  AND U19002 ( .A(n10833), .B(n10834), .Z(n10829) );
  NAND U19003 ( .A(n10835), .B(n10836), .Z(n10834) );
  NAND U19004 ( .A(n10837), .B(n10838), .Z(n10833) );
  AND U19005 ( .A(n10839), .B(n10840), .Z(n10825) );
  NAND U19006 ( .A(n10841), .B(n10842), .Z(n10840) );
  NAND U19007 ( .A(n10843), .B(n10844), .Z(n10839) );
  NANDN U19008 ( .A(n10845), .B(n10846), .Z(n10828) );
  ANDN U19009 ( .B(n10847), .A(n10848), .Z(n10822) );
  XNOR U19010 ( .A(n10813), .B(n10849), .Z(n10818) );
  XNOR U19011 ( .A(n10811), .B(n10815), .Z(n10849) );
  AND U19012 ( .A(n10850), .B(n10851), .Z(n10815) );
  NAND U19013 ( .A(n10852), .B(n10853), .Z(n10851) );
  NAND U19014 ( .A(n10854), .B(n10855), .Z(n10850) );
  AND U19015 ( .A(n10856), .B(n10857), .Z(n10811) );
  NAND U19016 ( .A(n10858), .B(n10859), .Z(n10857) );
  NAND U19017 ( .A(n10860), .B(n10861), .Z(n10856) );
  AND U19018 ( .A(n10862), .B(n10863), .Z(n10813) );
  NAND U19019 ( .A(n10864), .B(n10865), .Z(n10807) );
  XNOR U19020 ( .A(n10790), .B(n10866), .Z(n10804) );
  XNOR U19021 ( .A(n10794), .B(n10792), .Z(n10866) );
  XOR U19022 ( .A(n10800), .B(n10867), .Z(n10792) );
  XNOR U19023 ( .A(n10797), .B(n10801), .Z(n10867) );
  AND U19024 ( .A(n10868), .B(n10869), .Z(n10801) );
  NAND U19025 ( .A(n10870), .B(n10871), .Z(n10869) );
  NAND U19026 ( .A(n10872), .B(n10873), .Z(n10868) );
  AND U19027 ( .A(n10874), .B(n10875), .Z(n10797) );
  NAND U19028 ( .A(n10876), .B(n10877), .Z(n10875) );
  NAND U19029 ( .A(n10878), .B(n10879), .Z(n10874) );
  NANDN U19030 ( .A(n10880), .B(n10881), .Z(n10800) );
  ANDN U19031 ( .B(n10882), .A(n10883), .Z(n10794) );
  XNOR U19032 ( .A(n10785), .B(n10884), .Z(n10790) );
  XNOR U19033 ( .A(n10783), .B(n10787), .Z(n10884) );
  AND U19034 ( .A(n10885), .B(n10886), .Z(n10787) );
  NAND U19035 ( .A(n10887), .B(n10888), .Z(n10886) );
  NAND U19036 ( .A(n10889), .B(n10890), .Z(n10885) );
  AND U19037 ( .A(n10891), .B(n10892), .Z(n10783) );
  NAND U19038 ( .A(n10893), .B(n10894), .Z(n10892) );
  NAND U19039 ( .A(n10895), .B(n10896), .Z(n10891) );
  AND U19040 ( .A(n10897), .B(n10898), .Z(n10785) );
  XOR U19041 ( .A(n10865), .B(n10864), .Z(N64427) );
  XNOR U19042 ( .A(n10882), .B(n10883), .Z(n10864) );
  XNOR U19043 ( .A(n10897), .B(n10898), .Z(n10883) );
  XOR U19044 ( .A(n10894), .B(n10893), .Z(n10898) );
  XOR U19045 ( .A(y[7092]), .B(x[7092]), .Z(n10893) );
  XOR U19046 ( .A(n10896), .B(n10895), .Z(n10894) );
  XOR U19047 ( .A(y[7094]), .B(x[7094]), .Z(n10895) );
  XOR U19048 ( .A(y[7093]), .B(x[7093]), .Z(n10896) );
  XOR U19049 ( .A(n10888), .B(n10887), .Z(n10897) );
  XOR U19050 ( .A(n10890), .B(n10889), .Z(n10887) );
  XOR U19051 ( .A(y[7091]), .B(x[7091]), .Z(n10889) );
  XOR U19052 ( .A(y[7090]), .B(x[7090]), .Z(n10890) );
  XOR U19053 ( .A(y[7089]), .B(x[7089]), .Z(n10888) );
  XNOR U19054 ( .A(n10881), .B(n10880), .Z(n10882) );
  XNOR U19055 ( .A(n10877), .B(n10876), .Z(n10880) );
  XOR U19056 ( .A(n10879), .B(n10878), .Z(n10876) );
  XOR U19057 ( .A(y[7088]), .B(x[7088]), .Z(n10878) );
  XOR U19058 ( .A(y[7087]), .B(x[7087]), .Z(n10879) );
  XOR U19059 ( .A(y[7086]), .B(x[7086]), .Z(n10877) );
  XOR U19060 ( .A(n10871), .B(n10870), .Z(n10881) );
  XOR U19061 ( .A(n10873), .B(n10872), .Z(n10870) );
  XOR U19062 ( .A(y[7085]), .B(x[7085]), .Z(n10872) );
  XOR U19063 ( .A(y[7084]), .B(x[7084]), .Z(n10873) );
  XOR U19064 ( .A(y[7083]), .B(x[7083]), .Z(n10871) );
  XNOR U19065 ( .A(n10847), .B(n10848), .Z(n10865) );
  XNOR U19066 ( .A(n10862), .B(n10863), .Z(n10848) );
  XOR U19067 ( .A(n10859), .B(n10858), .Z(n10863) );
  XOR U19068 ( .A(y[7080]), .B(x[7080]), .Z(n10858) );
  XOR U19069 ( .A(n10861), .B(n10860), .Z(n10859) );
  XOR U19070 ( .A(y[7082]), .B(x[7082]), .Z(n10860) );
  XOR U19071 ( .A(y[7081]), .B(x[7081]), .Z(n10861) );
  XOR U19072 ( .A(n10853), .B(n10852), .Z(n10862) );
  XOR U19073 ( .A(n10855), .B(n10854), .Z(n10852) );
  XOR U19074 ( .A(y[7079]), .B(x[7079]), .Z(n10854) );
  XOR U19075 ( .A(y[7078]), .B(x[7078]), .Z(n10855) );
  XOR U19076 ( .A(y[7077]), .B(x[7077]), .Z(n10853) );
  XNOR U19077 ( .A(n10846), .B(n10845), .Z(n10847) );
  XNOR U19078 ( .A(n10842), .B(n10841), .Z(n10845) );
  XOR U19079 ( .A(n10844), .B(n10843), .Z(n10841) );
  XOR U19080 ( .A(y[7076]), .B(x[7076]), .Z(n10843) );
  XOR U19081 ( .A(y[7075]), .B(x[7075]), .Z(n10844) );
  XOR U19082 ( .A(y[7074]), .B(x[7074]), .Z(n10842) );
  XOR U19083 ( .A(n10836), .B(n10835), .Z(n10846) );
  XOR U19084 ( .A(n10838), .B(n10837), .Z(n10835) );
  XOR U19085 ( .A(y[7073]), .B(x[7073]), .Z(n10837) );
  XOR U19086 ( .A(y[7072]), .B(x[7072]), .Z(n10838) );
  XOR U19087 ( .A(y[7071]), .B(x[7071]), .Z(n10836) );
  NAND U19088 ( .A(n10899), .B(n10900), .Z(N64418) );
  NAND U19089 ( .A(n10901), .B(n10902), .Z(n10900) );
  NANDN U19090 ( .A(n10903), .B(n10904), .Z(n10902) );
  NANDN U19091 ( .A(n10904), .B(n10903), .Z(n10899) );
  XOR U19092 ( .A(n10903), .B(n10905), .Z(N64417) );
  XNOR U19093 ( .A(n10901), .B(n10904), .Z(n10905) );
  NAND U19094 ( .A(n10906), .B(n10907), .Z(n10904) );
  NAND U19095 ( .A(n10908), .B(n10909), .Z(n10907) );
  NANDN U19096 ( .A(n10910), .B(n10911), .Z(n10909) );
  NANDN U19097 ( .A(n10911), .B(n10910), .Z(n10906) );
  AND U19098 ( .A(n10912), .B(n10913), .Z(n10901) );
  NAND U19099 ( .A(n10914), .B(n10915), .Z(n10913) );
  NANDN U19100 ( .A(n10916), .B(n10917), .Z(n10915) );
  NANDN U19101 ( .A(n10917), .B(n10916), .Z(n10912) );
  IV U19102 ( .A(n10918), .Z(n10917) );
  AND U19103 ( .A(n10919), .B(n10920), .Z(n10903) );
  NAND U19104 ( .A(n10921), .B(n10922), .Z(n10920) );
  NANDN U19105 ( .A(n10923), .B(n10924), .Z(n10922) );
  NANDN U19106 ( .A(n10924), .B(n10923), .Z(n10919) );
  XOR U19107 ( .A(n10916), .B(n10925), .Z(N64416) );
  XNOR U19108 ( .A(n10914), .B(n10918), .Z(n10925) );
  XOR U19109 ( .A(n10911), .B(n10926), .Z(n10918) );
  XNOR U19110 ( .A(n10908), .B(n10910), .Z(n10926) );
  AND U19111 ( .A(n10927), .B(n10928), .Z(n10910) );
  NANDN U19112 ( .A(n10929), .B(n10930), .Z(n10928) );
  OR U19113 ( .A(n10931), .B(n10932), .Z(n10930) );
  IV U19114 ( .A(n10933), .Z(n10932) );
  NANDN U19115 ( .A(n10933), .B(n10931), .Z(n10927) );
  AND U19116 ( .A(n10934), .B(n10935), .Z(n10908) );
  NAND U19117 ( .A(n10936), .B(n10937), .Z(n10935) );
  NANDN U19118 ( .A(n10938), .B(n10939), .Z(n10937) );
  NANDN U19119 ( .A(n10939), .B(n10938), .Z(n10934) );
  IV U19120 ( .A(n10940), .Z(n10939) );
  NAND U19121 ( .A(n10941), .B(n10942), .Z(n10911) );
  NANDN U19122 ( .A(n10943), .B(n10944), .Z(n10942) );
  NANDN U19123 ( .A(n10945), .B(n10946), .Z(n10944) );
  NANDN U19124 ( .A(n10946), .B(n10945), .Z(n10941) );
  IV U19125 ( .A(n10947), .Z(n10945) );
  AND U19126 ( .A(n10948), .B(n10949), .Z(n10914) );
  NAND U19127 ( .A(n10950), .B(n10951), .Z(n10949) );
  NANDN U19128 ( .A(n10952), .B(n10953), .Z(n10951) );
  NANDN U19129 ( .A(n10953), .B(n10952), .Z(n10948) );
  XOR U19130 ( .A(n10924), .B(n10954), .Z(n10916) );
  XNOR U19131 ( .A(n10921), .B(n10923), .Z(n10954) );
  AND U19132 ( .A(n10955), .B(n10956), .Z(n10923) );
  NANDN U19133 ( .A(n10957), .B(n10958), .Z(n10956) );
  OR U19134 ( .A(n10959), .B(n10960), .Z(n10958) );
  IV U19135 ( .A(n10961), .Z(n10960) );
  NANDN U19136 ( .A(n10961), .B(n10959), .Z(n10955) );
  AND U19137 ( .A(n10962), .B(n10963), .Z(n10921) );
  NAND U19138 ( .A(n10964), .B(n10965), .Z(n10963) );
  NANDN U19139 ( .A(n10966), .B(n10967), .Z(n10965) );
  NANDN U19140 ( .A(n10967), .B(n10966), .Z(n10962) );
  IV U19141 ( .A(n10968), .Z(n10967) );
  NAND U19142 ( .A(n10969), .B(n10970), .Z(n10924) );
  NANDN U19143 ( .A(n10971), .B(n10972), .Z(n10970) );
  NANDN U19144 ( .A(n10973), .B(n10974), .Z(n10972) );
  NANDN U19145 ( .A(n10974), .B(n10973), .Z(n10969) );
  IV U19146 ( .A(n10975), .Z(n10973) );
  XOR U19147 ( .A(n10950), .B(n10976), .Z(N64415) );
  XNOR U19148 ( .A(n10953), .B(n10952), .Z(n10976) );
  XNOR U19149 ( .A(n10964), .B(n10977), .Z(n10952) );
  XNOR U19150 ( .A(n10968), .B(n10966), .Z(n10977) );
  XOR U19151 ( .A(n10974), .B(n10978), .Z(n10966) );
  XNOR U19152 ( .A(n10971), .B(n10975), .Z(n10978) );
  AND U19153 ( .A(n10979), .B(n10980), .Z(n10975) );
  NAND U19154 ( .A(n10981), .B(n10982), .Z(n10980) );
  NAND U19155 ( .A(n10983), .B(n10984), .Z(n10979) );
  AND U19156 ( .A(n10985), .B(n10986), .Z(n10971) );
  NAND U19157 ( .A(n10987), .B(n10988), .Z(n10986) );
  NAND U19158 ( .A(n10989), .B(n10990), .Z(n10985) );
  NANDN U19159 ( .A(n10991), .B(n10992), .Z(n10974) );
  ANDN U19160 ( .B(n10993), .A(n10994), .Z(n10968) );
  XNOR U19161 ( .A(n10959), .B(n10995), .Z(n10964) );
  XNOR U19162 ( .A(n10957), .B(n10961), .Z(n10995) );
  AND U19163 ( .A(n10996), .B(n10997), .Z(n10961) );
  NAND U19164 ( .A(n10998), .B(n10999), .Z(n10997) );
  NAND U19165 ( .A(n11000), .B(n11001), .Z(n10996) );
  AND U19166 ( .A(n11002), .B(n11003), .Z(n10957) );
  NAND U19167 ( .A(n11004), .B(n11005), .Z(n11003) );
  NAND U19168 ( .A(n11006), .B(n11007), .Z(n11002) );
  AND U19169 ( .A(n11008), .B(n11009), .Z(n10959) );
  NAND U19170 ( .A(n11010), .B(n11011), .Z(n10953) );
  XNOR U19171 ( .A(n10936), .B(n11012), .Z(n10950) );
  XNOR U19172 ( .A(n10940), .B(n10938), .Z(n11012) );
  XOR U19173 ( .A(n10946), .B(n11013), .Z(n10938) );
  XNOR U19174 ( .A(n10943), .B(n10947), .Z(n11013) );
  AND U19175 ( .A(n11014), .B(n11015), .Z(n10947) );
  NAND U19176 ( .A(n11016), .B(n11017), .Z(n11015) );
  NAND U19177 ( .A(n11018), .B(n11019), .Z(n11014) );
  AND U19178 ( .A(n11020), .B(n11021), .Z(n10943) );
  NAND U19179 ( .A(n11022), .B(n11023), .Z(n11021) );
  NAND U19180 ( .A(n11024), .B(n11025), .Z(n11020) );
  NANDN U19181 ( .A(n11026), .B(n11027), .Z(n10946) );
  ANDN U19182 ( .B(n11028), .A(n11029), .Z(n10940) );
  XNOR U19183 ( .A(n10931), .B(n11030), .Z(n10936) );
  XNOR U19184 ( .A(n10929), .B(n10933), .Z(n11030) );
  AND U19185 ( .A(n11031), .B(n11032), .Z(n10933) );
  NAND U19186 ( .A(n11033), .B(n11034), .Z(n11032) );
  NAND U19187 ( .A(n11035), .B(n11036), .Z(n11031) );
  AND U19188 ( .A(n11037), .B(n11038), .Z(n10929) );
  NAND U19189 ( .A(n11039), .B(n11040), .Z(n11038) );
  NAND U19190 ( .A(n11041), .B(n11042), .Z(n11037) );
  AND U19191 ( .A(n11043), .B(n11044), .Z(n10931) );
  XOR U19192 ( .A(n11011), .B(n11010), .Z(N64414) );
  XNOR U19193 ( .A(n11028), .B(n11029), .Z(n11010) );
  XNOR U19194 ( .A(n11043), .B(n11044), .Z(n11029) );
  XOR U19195 ( .A(n11040), .B(n11039), .Z(n11044) );
  XOR U19196 ( .A(y[7068]), .B(x[7068]), .Z(n11039) );
  XOR U19197 ( .A(n11042), .B(n11041), .Z(n11040) );
  XOR U19198 ( .A(y[7070]), .B(x[7070]), .Z(n11041) );
  XOR U19199 ( .A(y[7069]), .B(x[7069]), .Z(n11042) );
  XOR U19200 ( .A(n11034), .B(n11033), .Z(n11043) );
  XOR U19201 ( .A(n11036), .B(n11035), .Z(n11033) );
  XOR U19202 ( .A(y[7067]), .B(x[7067]), .Z(n11035) );
  XOR U19203 ( .A(y[7066]), .B(x[7066]), .Z(n11036) );
  XOR U19204 ( .A(y[7065]), .B(x[7065]), .Z(n11034) );
  XNOR U19205 ( .A(n11027), .B(n11026), .Z(n11028) );
  XNOR U19206 ( .A(n11023), .B(n11022), .Z(n11026) );
  XOR U19207 ( .A(n11025), .B(n11024), .Z(n11022) );
  XOR U19208 ( .A(y[7064]), .B(x[7064]), .Z(n11024) );
  XOR U19209 ( .A(y[7063]), .B(x[7063]), .Z(n11025) );
  XOR U19210 ( .A(y[7062]), .B(x[7062]), .Z(n11023) );
  XOR U19211 ( .A(n11017), .B(n11016), .Z(n11027) );
  XOR U19212 ( .A(n11019), .B(n11018), .Z(n11016) );
  XOR U19213 ( .A(y[7061]), .B(x[7061]), .Z(n11018) );
  XOR U19214 ( .A(y[7060]), .B(x[7060]), .Z(n11019) );
  XOR U19215 ( .A(y[7059]), .B(x[7059]), .Z(n11017) );
  XNOR U19216 ( .A(n10993), .B(n10994), .Z(n11011) );
  XNOR U19217 ( .A(n11008), .B(n11009), .Z(n10994) );
  XOR U19218 ( .A(n11005), .B(n11004), .Z(n11009) );
  XOR U19219 ( .A(y[7056]), .B(x[7056]), .Z(n11004) );
  XOR U19220 ( .A(n11007), .B(n11006), .Z(n11005) );
  XOR U19221 ( .A(y[7058]), .B(x[7058]), .Z(n11006) );
  XOR U19222 ( .A(y[7057]), .B(x[7057]), .Z(n11007) );
  XOR U19223 ( .A(n10999), .B(n10998), .Z(n11008) );
  XOR U19224 ( .A(n11001), .B(n11000), .Z(n10998) );
  XOR U19225 ( .A(y[7055]), .B(x[7055]), .Z(n11000) );
  XOR U19226 ( .A(y[7054]), .B(x[7054]), .Z(n11001) );
  XOR U19227 ( .A(y[7053]), .B(x[7053]), .Z(n10999) );
  XNOR U19228 ( .A(n10992), .B(n10991), .Z(n10993) );
  XNOR U19229 ( .A(n10988), .B(n10987), .Z(n10991) );
  XOR U19230 ( .A(n10990), .B(n10989), .Z(n10987) );
  XOR U19231 ( .A(y[7052]), .B(x[7052]), .Z(n10989) );
  XOR U19232 ( .A(y[7051]), .B(x[7051]), .Z(n10990) );
  XOR U19233 ( .A(y[7050]), .B(x[7050]), .Z(n10988) );
  XOR U19234 ( .A(n10982), .B(n10981), .Z(n10992) );
  XOR U19235 ( .A(n10984), .B(n10983), .Z(n10981) );
  XOR U19236 ( .A(y[7049]), .B(x[7049]), .Z(n10983) );
  XOR U19237 ( .A(y[7048]), .B(x[7048]), .Z(n10984) );
  XOR U19238 ( .A(y[7047]), .B(x[7047]), .Z(n10982) );
  NAND U19239 ( .A(n11045), .B(n11046), .Z(N64405) );
  NAND U19240 ( .A(n11047), .B(n11048), .Z(n11046) );
  NANDN U19241 ( .A(n11049), .B(n11050), .Z(n11048) );
  NANDN U19242 ( .A(n11050), .B(n11049), .Z(n11045) );
  XOR U19243 ( .A(n11049), .B(n11051), .Z(N64404) );
  XNOR U19244 ( .A(n11047), .B(n11050), .Z(n11051) );
  NAND U19245 ( .A(n11052), .B(n11053), .Z(n11050) );
  NAND U19246 ( .A(n11054), .B(n11055), .Z(n11053) );
  NANDN U19247 ( .A(n11056), .B(n11057), .Z(n11055) );
  NANDN U19248 ( .A(n11057), .B(n11056), .Z(n11052) );
  AND U19249 ( .A(n11058), .B(n11059), .Z(n11047) );
  NAND U19250 ( .A(n11060), .B(n11061), .Z(n11059) );
  NANDN U19251 ( .A(n11062), .B(n11063), .Z(n11061) );
  NANDN U19252 ( .A(n11063), .B(n11062), .Z(n11058) );
  IV U19253 ( .A(n11064), .Z(n11063) );
  AND U19254 ( .A(n11065), .B(n11066), .Z(n11049) );
  NAND U19255 ( .A(n11067), .B(n11068), .Z(n11066) );
  NANDN U19256 ( .A(n11069), .B(n11070), .Z(n11068) );
  NANDN U19257 ( .A(n11070), .B(n11069), .Z(n11065) );
  XOR U19258 ( .A(n11062), .B(n11071), .Z(N64403) );
  XNOR U19259 ( .A(n11060), .B(n11064), .Z(n11071) );
  XOR U19260 ( .A(n11057), .B(n11072), .Z(n11064) );
  XNOR U19261 ( .A(n11054), .B(n11056), .Z(n11072) );
  AND U19262 ( .A(n11073), .B(n11074), .Z(n11056) );
  NANDN U19263 ( .A(n11075), .B(n11076), .Z(n11074) );
  OR U19264 ( .A(n11077), .B(n11078), .Z(n11076) );
  IV U19265 ( .A(n11079), .Z(n11078) );
  NANDN U19266 ( .A(n11079), .B(n11077), .Z(n11073) );
  AND U19267 ( .A(n11080), .B(n11081), .Z(n11054) );
  NAND U19268 ( .A(n11082), .B(n11083), .Z(n11081) );
  NANDN U19269 ( .A(n11084), .B(n11085), .Z(n11083) );
  NANDN U19270 ( .A(n11085), .B(n11084), .Z(n11080) );
  IV U19271 ( .A(n11086), .Z(n11085) );
  NAND U19272 ( .A(n11087), .B(n11088), .Z(n11057) );
  NANDN U19273 ( .A(n11089), .B(n11090), .Z(n11088) );
  NANDN U19274 ( .A(n11091), .B(n11092), .Z(n11090) );
  NANDN U19275 ( .A(n11092), .B(n11091), .Z(n11087) );
  IV U19276 ( .A(n11093), .Z(n11091) );
  AND U19277 ( .A(n11094), .B(n11095), .Z(n11060) );
  NAND U19278 ( .A(n11096), .B(n11097), .Z(n11095) );
  NANDN U19279 ( .A(n11098), .B(n11099), .Z(n11097) );
  NANDN U19280 ( .A(n11099), .B(n11098), .Z(n11094) );
  XOR U19281 ( .A(n11070), .B(n11100), .Z(n11062) );
  XNOR U19282 ( .A(n11067), .B(n11069), .Z(n11100) );
  AND U19283 ( .A(n11101), .B(n11102), .Z(n11069) );
  NANDN U19284 ( .A(n11103), .B(n11104), .Z(n11102) );
  OR U19285 ( .A(n11105), .B(n11106), .Z(n11104) );
  IV U19286 ( .A(n11107), .Z(n11106) );
  NANDN U19287 ( .A(n11107), .B(n11105), .Z(n11101) );
  AND U19288 ( .A(n11108), .B(n11109), .Z(n11067) );
  NAND U19289 ( .A(n11110), .B(n11111), .Z(n11109) );
  NANDN U19290 ( .A(n11112), .B(n11113), .Z(n11111) );
  NANDN U19291 ( .A(n11113), .B(n11112), .Z(n11108) );
  IV U19292 ( .A(n11114), .Z(n11113) );
  NAND U19293 ( .A(n11115), .B(n11116), .Z(n11070) );
  NANDN U19294 ( .A(n11117), .B(n11118), .Z(n11116) );
  NANDN U19295 ( .A(n11119), .B(n11120), .Z(n11118) );
  NANDN U19296 ( .A(n11120), .B(n11119), .Z(n11115) );
  IV U19297 ( .A(n11121), .Z(n11119) );
  XOR U19298 ( .A(n11096), .B(n11122), .Z(N64402) );
  XNOR U19299 ( .A(n11099), .B(n11098), .Z(n11122) );
  XNOR U19300 ( .A(n11110), .B(n11123), .Z(n11098) );
  XNOR U19301 ( .A(n11114), .B(n11112), .Z(n11123) );
  XOR U19302 ( .A(n11120), .B(n11124), .Z(n11112) );
  XNOR U19303 ( .A(n11117), .B(n11121), .Z(n11124) );
  AND U19304 ( .A(n11125), .B(n11126), .Z(n11121) );
  NAND U19305 ( .A(n11127), .B(n11128), .Z(n11126) );
  NAND U19306 ( .A(n11129), .B(n11130), .Z(n11125) );
  AND U19307 ( .A(n11131), .B(n11132), .Z(n11117) );
  NAND U19308 ( .A(n11133), .B(n11134), .Z(n11132) );
  NAND U19309 ( .A(n11135), .B(n11136), .Z(n11131) );
  NANDN U19310 ( .A(n11137), .B(n11138), .Z(n11120) );
  ANDN U19311 ( .B(n11139), .A(n11140), .Z(n11114) );
  XNOR U19312 ( .A(n11105), .B(n11141), .Z(n11110) );
  XNOR U19313 ( .A(n11103), .B(n11107), .Z(n11141) );
  AND U19314 ( .A(n11142), .B(n11143), .Z(n11107) );
  NAND U19315 ( .A(n11144), .B(n11145), .Z(n11143) );
  NAND U19316 ( .A(n11146), .B(n11147), .Z(n11142) );
  AND U19317 ( .A(n11148), .B(n11149), .Z(n11103) );
  NAND U19318 ( .A(n11150), .B(n11151), .Z(n11149) );
  NAND U19319 ( .A(n11152), .B(n11153), .Z(n11148) );
  AND U19320 ( .A(n11154), .B(n11155), .Z(n11105) );
  NAND U19321 ( .A(n11156), .B(n11157), .Z(n11099) );
  XNOR U19322 ( .A(n11082), .B(n11158), .Z(n11096) );
  XNOR U19323 ( .A(n11086), .B(n11084), .Z(n11158) );
  XOR U19324 ( .A(n11092), .B(n11159), .Z(n11084) );
  XNOR U19325 ( .A(n11089), .B(n11093), .Z(n11159) );
  AND U19326 ( .A(n11160), .B(n11161), .Z(n11093) );
  NAND U19327 ( .A(n11162), .B(n11163), .Z(n11161) );
  NAND U19328 ( .A(n11164), .B(n11165), .Z(n11160) );
  AND U19329 ( .A(n11166), .B(n11167), .Z(n11089) );
  NAND U19330 ( .A(n11168), .B(n11169), .Z(n11167) );
  NAND U19331 ( .A(n11170), .B(n11171), .Z(n11166) );
  NANDN U19332 ( .A(n11172), .B(n11173), .Z(n11092) );
  ANDN U19333 ( .B(n11174), .A(n11175), .Z(n11086) );
  XNOR U19334 ( .A(n11077), .B(n11176), .Z(n11082) );
  XNOR U19335 ( .A(n11075), .B(n11079), .Z(n11176) );
  AND U19336 ( .A(n11177), .B(n11178), .Z(n11079) );
  NAND U19337 ( .A(n11179), .B(n11180), .Z(n11178) );
  NAND U19338 ( .A(n11181), .B(n11182), .Z(n11177) );
  AND U19339 ( .A(n11183), .B(n11184), .Z(n11075) );
  NAND U19340 ( .A(n11185), .B(n11186), .Z(n11184) );
  NAND U19341 ( .A(n11187), .B(n11188), .Z(n11183) );
  AND U19342 ( .A(n11189), .B(n11190), .Z(n11077) );
  XOR U19343 ( .A(n11157), .B(n11156), .Z(N64401) );
  XNOR U19344 ( .A(n11174), .B(n11175), .Z(n11156) );
  XNOR U19345 ( .A(n11189), .B(n11190), .Z(n11175) );
  XOR U19346 ( .A(n11186), .B(n11185), .Z(n11190) );
  XOR U19347 ( .A(y[7044]), .B(x[7044]), .Z(n11185) );
  XOR U19348 ( .A(n11188), .B(n11187), .Z(n11186) );
  XOR U19349 ( .A(y[7046]), .B(x[7046]), .Z(n11187) );
  XOR U19350 ( .A(y[7045]), .B(x[7045]), .Z(n11188) );
  XOR U19351 ( .A(n11180), .B(n11179), .Z(n11189) );
  XOR U19352 ( .A(n11182), .B(n11181), .Z(n11179) );
  XOR U19353 ( .A(y[7043]), .B(x[7043]), .Z(n11181) );
  XOR U19354 ( .A(y[7042]), .B(x[7042]), .Z(n11182) );
  XOR U19355 ( .A(y[7041]), .B(x[7041]), .Z(n11180) );
  XNOR U19356 ( .A(n11173), .B(n11172), .Z(n11174) );
  XNOR U19357 ( .A(n11169), .B(n11168), .Z(n11172) );
  XOR U19358 ( .A(n11171), .B(n11170), .Z(n11168) );
  XOR U19359 ( .A(y[7040]), .B(x[7040]), .Z(n11170) );
  XOR U19360 ( .A(y[7039]), .B(x[7039]), .Z(n11171) );
  XOR U19361 ( .A(y[7038]), .B(x[7038]), .Z(n11169) );
  XOR U19362 ( .A(n11163), .B(n11162), .Z(n11173) );
  XOR U19363 ( .A(n11165), .B(n11164), .Z(n11162) );
  XOR U19364 ( .A(y[7037]), .B(x[7037]), .Z(n11164) );
  XOR U19365 ( .A(y[7036]), .B(x[7036]), .Z(n11165) );
  XOR U19366 ( .A(y[7035]), .B(x[7035]), .Z(n11163) );
  XNOR U19367 ( .A(n11139), .B(n11140), .Z(n11157) );
  XNOR U19368 ( .A(n11154), .B(n11155), .Z(n11140) );
  XOR U19369 ( .A(n11151), .B(n11150), .Z(n11155) );
  XOR U19370 ( .A(y[7032]), .B(x[7032]), .Z(n11150) );
  XOR U19371 ( .A(n11153), .B(n11152), .Z(n11151) );
  XOR U19372 ( .A(y[7034]), .B(x[7034]), .Z(n11152) );
  XOR U19373 ( .A(y[7033]), .B(x[7033]), .Z(n11153) );
  XOR U19374 ( .A(n11145), .B(n11144), .Z(n11154) );
  XOR U19375 ( .A(n11147), .B(n11146), .Z(n11144) );
  XOR U19376 ( .A(y[7031]), .B(x[7031]), .Z(n11146) );
  XOR U19377 ( .A(y[7030]), .B(x[7030]), .Z(n11147) );
  XOR U19378 ( .A(y[7029]), .B(x[7029]), .Z(n11145) );
  XNOR U19379 ( .A(n11138), .B(n11137), .Z(n11139) );
  XNOR U19380 ( .A(n11134), .B(n11133), .Z(n11137) );
  XOR U19381 ( .A(n11136), .B(n11135), .Z(n11133) );
  XOR U19382 ( .A(y[7028]), .B(x[7028]), .Z(n11135) );
  XOR U19383 ( .A(y[7027]), .B(x[7027]), .Z(n11136) );
  XOR U19384 ( .A(y[7026]), .B(x[7026]), .Z(n11134) );
  XOR U19385 ( .A(n11128), .B(n11127), .Z(n11138) );
  XOR U19386 ( .A(n11130), .B(n11129), .Z(n11127) );
  XOR U19387 ( .A(y[7025]), .B(x[7025]), .Z(n11129) );
  XOR U19388 ( .A(y[7024]), .B(x[7024]), .Z(n11130) );
  XOR U19389 ( .A(y[7023]), .B(x[7023]), .Z(n11128) );
  NAND U19390 ( .A(n11191), .B(n11192), .Z(N64392) );
  NAND U19391 ( .A(n11193), .B(n11194), .Z(n11192) );
  NANDN U19392 ( .A(n11195), .B(n11196), .Z(n11194) );
  NANDN U19393 ( .A(n11196), .B(n11195), .Z(n11191) );
  XOR U19394 ( .A(n11195), .B(n11197), .Z(N64391) );
  XNOR U19395 ( .A(n11193), .B(n11196), .Z(n11197) );
  NAND U19396 ( .A(n11198), .B(n11199), .Z(n11196) );
  NAND U19397 ( .A(n11200), .B(n11201), .Z(n11199) );
  NANDN U19398 ( .A(n11202), .B(n11203), .Z(n11201) );
  NANDN U19399 ( .A(n11203), .B(n11202), .Z(n11198) );
  AND U19400 ( .A(n11204), .B(n11205), .Z(n11193) );
  NAND U19401 ( .A(n11206), .B(n11207), .Z(n11205) );
  NANDN U19402 ( .A(n11208), .B(n11209), .Z(n11207) );
  NANDN U19403 ( .A(n11209), .B(n11208), .Z(n11204) );
  IV U19404 ( .A(n11210), .Z(n11209) );
  AND U19405 ( .A(n11211), .B(n11212), .Z(n11195) );
  NAND U19406 ( .A(n11213), .B(n11214), .Z(n11212) );
  NANDN U19407 ( .A(n11215), .B(n11216), .Z(n11214) );
  NANDN U19408 ( .A(n11216), .B(n11215), .Z(n11211) );
  XOR U19409 ( .A(n11208), .B(n11217), .Z(N64390) );
  XNOR U19410 ( .A(n11206), .B(n11210), .Z(n11217) );
  XOR U19411 ( .A(n11203), .B(n11218), .Z(n11210) );
  XNOR U19412 ( .A(n11200), .B(n11202), .Z(n11218) );
  AND U19413 ( .A(n11219), .B(n11220), .Z(n11202) );
  NANDN U19414 ( .A(n11221), .B(n11222), .Z(n11220) );
  OR U19415 ( .A(n11223), .B(n11224), .Z(n11222) );
  IV U19416 ( .A(n11225), .Z(n11224) );
  NANDN U19417 ( .A(n11225), .B(n11223), .Z(n11219) );
  AND U19418 ( .A(n11226), .B(n11227), .Z(n11200) );
  NAND U19419 ( .A(n11228), .B(n11229), .Z(n11227) );
  NANDN U19420 ( .A(n11230), .B(n11231), .Z(n11229) );
  NANDN U19421 ( .A(n11231), .B(n11230), .Z(n11226) );
  IV U19422 ( .A(n11232), .Z(n11231) );
  NAND U19423 ( .A(n11233), .B(n11234), .Z(n11203) );
  NANDN U19424 ( .A(n11235), .B(n11236), .Z(n11234) );
  NANDN U19425 ( .A(n11237), .B(n11238), .Z(n11236) );
  NANDN U19426 ( .A(n11238), .B(n11237), .Z(n11233) );
  IV U19427 ( .A(n11239), .Z(n11237) );
  AND U19428 ( .A(n11240), .B(n11241), .Z(n11206) );
  NAND U19429 ( .A(n11242), .B(n11243), .Z(n11241) );
  NANDN U19430 ( .A(n11244), .B(n11245), .Z(n11243) );
  NANDN U19431 ( .A(n11245), .B(n11244), .Z(n11240) );
  XOR U19432 ( .A(n11216), .B(n11246), .Z(n11208) );
  XNOR U19433 ( .A(n11213), .B(n11215), .Z(n11246) );
  AND U19434 ( .A(n11247), .B(n11248), .Z(n11215) );
  NANDN U19435 ( .A(n11249), .B(n11250), .Z(n11248) );
  OR U19436 ( .A(n11251), .B(n11252), .Z(n11250) );
  IV U19437 ( .A(n11253), .Z(n11252) );
  NANDN U19438 ( .A(n11253), .B(n11251), .Z(n11247) );
  AND U19439 ( .A(n11254), .B(n11255), .Z(n11213) );
  NAND U19440 ( .A(n11256), .B(n11257), .Z(n11255) );
  NANDN U19441 ( .A(n11258), .B(n11259), .Z(n11257) );
  NANDN U19442 ( .A(n11259), .B(n11258), .Z(n11254) );
  IV U19443 ( .A(n11260), .Z(n11259) );
  NAND U19444 ( .A(n11261), .B(n11262), .Z(n11216) );
  NANDN U19445 ( .A(n11263), .B(n11264), .Z(n11262) );
  NANDN U19446 ( .A(n11265), .B(n11266), .Z(n11264) );
  NANDN U19447 ( .A(n11266), .B(n11265), .Z(n11261) );
  IV U19448 ( .A(n11267), .Z(n11265) );
  XOR U19449 ( .A(n11242), .B(n11268), .Z(N64389) );
  XNOR U19450 ( .A(n11245), .B(n11244), .Z(n11268) );
  XNOR U19451 ( .A(n11256), .B(n11269), .Z(n11244) );
  XNOR U19452 ( .A(n11260), .B(n11258), .Z(n11269) );
  XOR U19453 ( .A(n11266), .B(n11270), .Z(n11258) );
  XNOR U19454 ( .A(n11263), .B(n11267), .Z(n11270) );
  AND U19455 ( .A(n11271), .B(n11272), .Z(n11267) );
  NAND U19456 ( .A(n11273), .B(n11274), .Z(n11272) );
  NAND U19457 ( .A(n11275), .B(n11276), .Z(n11271) );
  AND U19458 ( .A(n11277), .B(n11278), .Z(n11263) );
  NAND U19459 ( .A(n11279), .B(n11280), .Z(n11278) );
  NAND U19460 ( .A(n11281), .B(n11282), .Z(n11277) );
  NANDN U19461 ( .A(n11283), .B(n11284), .Z(n11266) );
  ANDN U19462 ( .B(n11285), .A(n11286), .Z(n11260) );
  XNOR U19463 ( .A(n11251), .B(n11287), .Z(n11256) );
  XNOR U19464 ( .A(n11249), .B(n11253), .Z(n11287) );
  AND U19465 ( .A(n11288), .B(n11289), .Z(n11253) );
  NAND U19466 ( .A(n11290), .B(n11291), .Z(n11289) );
  NAND U19467 ( .A(n11292), .B(n11293), .Z(n11288) );
  AND U19468 ( .A(n11294), .B(n11295), .Z(n11249) );
  NAND U19469 ( .A(n11296), .B(n11297), .Z(n11295) );
  NAND U19470 ( .A(n11298), .B(n11299), .Z(n11294) );
  AND U19471 ( .A(n11300), .B(n11301), .Z(n11251) );
  NAND U19472 ( .A(n11302), .B(n11303), .Z(n11245) );
  XNOR U19473 ( .A(n11228), .B(n11304), .Z(n11242) );
  XNOR U19474 ( .A(n11232), .B(n11230), .Z(n11304) );
  XOR U19475 ( .A(n11238), .B(n11305), .Z(n11230) );
  XNOR U19476 ( .A(n11235), .B(n11239), .Z(n11305) );
  AND U19477 ( .A(n11306), .B(n11307), .Z(n11239) );
  NAND U19478 ( .A(n11308), .B(n11309), .Z(n11307) );
  NAND U19479 ( .A(n11310), .B(n11311), .Z(n11306) );
  AND U19480 ( .A(n11312), .B(n11313), .Z(n11235) );
  NAND U19481 ( .A(n11314), .B(n11315), .Z(n11313) );
  NAND U19482 ( .A(n11316), .B(n11317), .Z(n11312) );
  NANDN U19483 ( .A(n11318), .B(n11319), .Z(n11238) );
  ANDN U19484 ( .B(n11320), .A(n11321), .Z(n11232) );
  XNOR U19485 ( .A(n11223), .B(n11322), .Z(n11228) );
  XNOR U19486 ( .A(n11221), .B(n11225), .Z(n11322) );
  AND U19487 ( .A(n11323), .B(n11324), .Z(n11225) );
  NAND U19488 ( .A(n11325), .B(n11326), .Z(n11324) );
  NAND U19489 ( .A(n11327), .B(n11328), .Z(n11323) );
  AND U19490 ( .A(n11329), .B(n11330), .Z(n11221) );
  NAND U19491 ( .A(n11331), .B(n11332), .Z(n11330) );
  NAND U19492 ( .A(n11333), .B(n11334), .Z(n11329) );
  AND U19493 ( .A(n11335), .B(n11336), .Z(n11223) );
  XOR U19494 ( .A(n11303), .B(n11302), .Z(N64388) );
  XNOR U19495 ( .A(n11320), .B(n11321), .Z(n11302) );
  XNOR U19496 ( .A(n11335), .B(n11336), .Z(n11321) );
  XOR U19497 ( .A(n11332), .B(n11331), .Z(n11336) );
  XOR U19498 ( .A(y[7020]), .B(x[7020]), .Z(n11331) );
  XOR U19499 ( .A(n11334), .B(n11333), .Z(n11332) );
  XOR U19500 ( .A(y[7022]), .B(x[7022]), .Z(n11333) );
  XOR U19501 ( .A(y[7021]), .B(x[7021]), .Z(n11334) );
  XOR U19502 ( .A(n11326), .B(n11325), .Z(n11335) );
  XOR U19503 ( .A(n11328), .B(n11327), .Z(n11325) );
  XOR U19504 ( .A(y[7019]), .B(x[7019]), .Z(n11327) );
  XOR U19505 ( .A(y[7018]), .B(x[7018]), .Z(n11328) );
  XOR U19506 ( .A(y[7017]), .B(x[7017]), .Z(n11326) );
  XNOR U19507 ( .A(n11319), .B(n11318), .Z(n11320) );
  XNOR U19508 ( .A(n11315), .B(n11314), .Z(n11318) );
  XOR U19509 ( .A(n11317), .B(n11316), .Z(n11314) );
  XOR U19510 ( .A(y[7016]), .B(x[7016]), .Z(n11316) );
  XOR U19511 ( .A(y[7015]), .B(x[7015]), .Z(n11317) );
  XOR U19512 ( .A(y[7014]), .B(x[7014]), .Z(n11315) );
  XOR U19513 ( .A(n11309), .B(n11308), .Z(n11319) );
  XOR U19514 ( .A(n11311), .B(n11310), .Z(n11308) );
  XOR U19515 ( .A(y[7013]), .B(x[7013]), .Z(n11310) );
  XOR U19516 ( .A(y[7012]), .B(x[7012]), .Z(n11311) );
  XOR U19517 ( .A(y[7011]), .B(x[7011]), .Z(n11309) );
  XNOR U19518 ( .A(n11285), .B(n11286), .Z(n11303) );
  XNOR U19519 ( .A(n11300), .B(n11301), .Z(n11286) );
  XOR U19520 ( .A(n11297), .B(n11296), .Z(n11301) );
  XOR U19521 ( .A(y[7008]), .B(x[7008]), .Z(n11296) );
  XOR U19522 ( .A(n11299), .B(n11298), .Z(n11297) );
  XOR U19523 ( .A(y[7010]), .B(x[7010]), .Z(n11298) );
  XOR U19524 ( .A(y[7009]), .B(x[7009]), .Z(n11299) );
  XOR U19525 ( .A(n11291), .B(n11290), .Z(n11300) );
  XOR U19526 ( .A(n11293), .B(n11292), .Z(n11290) );
  XOR U19527 ( .A(y[7007]), .B(x[7007]), .Z(n11292) );
  XOR U19528 ( .A(y[7006]), .B(x[7006]), .Z(n11293) );
  XOR U19529 ( .A(y[7005]), .B(x[7005]), .Z(n11291) );
  XNOR U19530 ( .A(n11284), .B(n11283), .Z(n11285) );
  XNOR U19531 ( .A(n11280), .B(n11279), .Z(n11283) );
  XOR U19532 ( .A(n11282), .B(n11281), .Z(n11279) );
  XOR U19533 ( .A(y[7004]), .B(x[7004]), .Z(n11281) );
  XOR U19534 ( .A(y[7003]), .B(x[7003]), .Z(n11282) );
  XOR U19535 ( .A(y[7002]), .B(x[7002]), .Z(n11280) );
  XOR U19536 ( .A(n11274), .B(n11273), .Z(n11284) );
  XOR U19537 ( .A(n11276), .B(n11275), .Z(n11273) );
  XOR U19538 ( .A(y[7001]), .B(x[7001]), .Z(n11275) );
  XOR U19539 ( .A(y[7000]), .B(x[7000]), .Z(n11276) );
  XOR U19540 ( .A(y[6999]), .B(x[6999]), .Z(n11274) );
  NAND U19541 ( .A(n11337), .B(n11338), .Z(N64379) );
  NAND U19542 ( .A(n11339), .B(n11340), .Z(n11338) );
  NANDN U19543 ( .A(n11341), .B(n11342), .Z(n11340) );
  NANDN U19544 ( .A(n11342), .B(n11341), .Z(n11337) );
  XOR U19545 ( .A(n11341), .B(n11343), .Z(N64378) );
  XNOR U19546 ( .A(n11339), .B(n11342), .Z(n11343) );
  NAND U19547 ( .A(n11344), .B(n11345), .Z(n11342) );
  NAND U19548 ( .A(n11346), .B(n11347), .Z(n11345) );
  NANDN U19549 ( .A(n11348), .B(n11349), .Z(n11347) );
  NANDN U19550 ( .A(n11349), .B(n11348), .Z(n11344) );
  AND U19551 ( .A(n11350), .B(n11351), .Z(n11339) );
  NAND U19552 ( .A(n11352), .B(n11353), .Z(n11351) );
  NANDN U19553 ( .A(n11354), .B(n11355), .Z(n11353) );
  NANDN U19554 ( .A(n11355), .B(n11354), .Z(n11350) );
  IV U19555 ( .A(n11356), .Z(n11355) );
  AND U19556 ( .A(n11357), .B(n11358), .Z(n11341) );
  NAND U19557 ( .A(n11359), .B(n11360), .Z(n11358) );
  NANDN U19558 ( .A(n11361), .B(n11362), .Z(n11360) );
  NANDN U19559 ( .A(n11362), .B(n11361), .Z(n11357) );
  XOR U19560 ( .A(n11354), .B(n11363), .Z(N64377) );
  XNOR U19561 ( .A(n11352), .B(n11356), .Z(n11363) );
  XOR U19562 ( .A(n11349), .B(n11364), .Z(n11356) );
  XNOR U19563 ( .A(n11346), .B(n11348), .Z(n11364) );
  AND U19564 ( .A(n11365), .B(n11366), .Z(n11348) );
  NANDN U19565 ( .A(n11367), .B(n11368), .Z(n11366) );
  OR U19566 ( .A(n11369), .B(n11370), .Z(n11368) );
  IV U19567 ( .A(n11371), .Z(n11370) );
  NANDN U19568 ( .A(n11371), .B(n11369), .Z(n11365) );
  AND U19569 ( .A(n11372), .B(n11373), .Z(n11346) );
  NAND U19570 ( .A(n11374), .B(n11375), .Z(n11373) );
  NANDN U19571 ( .A(n11376), .B(n11377), .Z(n11375) );
  NANDN U19572 ( .A(n11377), .B(n11376), .Z(n11372) );
  IV U19573 ( .A(n11378), .Z(n11377) );
  NAND U19574 ( .A(n11379), .B(n11380), .Z(n11349) );
  NANDN U19575 ( .A(n11381), .B(n11382), .Z(n11380) );
  NANDN U19576 ( .A(n11383), .B(n11384), .Z(n11382) );
  NANDN U19577 ( .A(n11384), .B(n11383), .Z(n11379) );
  IV U19578 ( .A(n11385), .Z(n11383) );
  AND U19579 ( .A(n11386), .B(n11387), .Z(n11352) );
  NAND U19580 ( .A(n11388), .B(n11389), .Z(n11387) );
  NANDN U19581 ( .A(n11390), .B(n11391), .Z(n11389) );
  NANDN U19582 ( .A(n11391), .B(n11390), .Z(n11386) );
  XOR U19583 ( .A(n11362), .B(n11392), .Z(n11354) );
  XNOR U19584 ( .A(n11359), .B(n11361), .Z(n11392) );
  AND U19585 ( .A(n11393), .B(n11394), .Z(n11361) );
  NANDN U19586 ( .A(n11395), .B(n11396), .Z(n11394) );
  OR U19587 ( .A(n11397), .B(n11398), .Z(n11396) );
  IV U19588 ( .A(n11399), .Z(n11398) );
  NANDN U19589 ( .A(n11399), .B(n11397), .Z(n11393) );
  AND U19590 ( .A(n11400), .B(n11401), .Z(n11359) );
  NAND U19591 ( .A(n11402), .B(n11403), .Z(n11401) );
  NANDN U19592 ( .A(n11404), .B(n11405), .Z(n11403) );
  NANDN U19593 ( .A(n11405), .B(n11404), .Z(n11400) );
  IV U19594 ( .A(n11406), .Z(n11405) );
  NAND U19595 ( .A(n11407), .B(n11408), .Z(n11362) );
  NANDN U19596 ( .A(n11409), .B(n11410), .Z(n11408) );
  NANDN U19597 ( .A(n11411), .B(n11412), .Z(n11410) );
  NANDN U19598 ( .A(n11412), .B(n11411), .Z(n11407) );
  IV U19599 ( .A(n11413), .Z(n11411) );
  XOR U19600 ( .A(n11388), .B(n11414), .Z(N64376) );
  XNOR U19601 ( .A(n11391), .B(n11390), .Z(n11414) );
  XNOR U19602 ( .A(n11402), .B(n11415), .Z(n11390) );
  XNOR U19603 ( .A(n11406), .B(n11404), .Z(n11415) );
  XOR U19604 ( .A(n11412), .B(n11416), .Z(n11404) );
  XNOR U19605 ( .A(n11409), .B(n11413), .Z(n11416) );
  AND U19606 ( .A(n11417), .B(n11418), .Z(n11413) );
  NAND U19607 ( .A(n11419), .B(n11420), .Z(n11418) );
  NAND U19608 ( .A(n11421), .B(n11422), .Z(n11417) );
  AND U19609 ( .A(n11423), .B(n11424), .Z(n11409) );
  NAND U19610 ( .A(n11425), .B(n11426), .Z(n11424) );
  NAND U19611 ( .A(n11427), .B(n11428), .Z(n11423) );
  NANDN U19612 ( .A(n11429), .B(n11430), .Z(n11412) );
  ANDN U19613 ( .B(n11431), .A(n11432), .Z(n11406) );
  XNOR U19614 ( .A(n11397), .B(n11433), .Z(n11402) );
  XNOR U19615 ( .A(n11395), .B(n11399), .Z(n11433) );
  AND U19616 ( .A(n11434), .B(n11435), .Z(n11399) );
  NAND U19617 ( .A(n11436), .B(n11437), .Z(n11435) );
  NAND U19618 ( .A(n11438), .B(n11439), .Z(n11434) );
  AND U19619 ( .A(n11440), .B(n11441), .Z(n11395) );
  NAND U19620 ( .A(n11442), .B(n11443), .Z(n11441) );
  NAND U19621 ( .A(n11444), .B(n11445), .Z(n11440) );
  AND U19622 ( .A(n11446), .B(n11447), .Z(n11397) );
  NAND U19623 ( .A(n11448), .B(n11449), .Z(n11391) );
  XNOR U19624 ( .A(n11374), .B(n11450), .Z(n11388) );
  XNOR U19625 ( .A(n11378), .B(n11376), .Z(n11450) );
  XOR U19626 ( .A(n11384), .B(n11451), .Z(n11376) );
  XNOR U19627 ( .A(n11381), .B(n11385), .Z(n11451) );
  AND U19628 ( .A(n11452), .B(n11453), .Z(n11385) );
  NAND U19629 ( .A(n11454), .B(n11455), .Z(n11453) );
  NAND U19630 ( .A(n11456), .B(n11457), .Z(n11452) );
  AND U19631 ( .A(n11458), .B(n11459), .Z(n11381) );
  NAND U19632 ( .A(n11460), .B(n11461), .Z(n11459) );
  NAND U19633 ( .A(n11462), .B(n11463), .Z(n11458) );
  NANDN U19634 ( .A(n11464), .B(n11465), .Z(n11384) );
  ANDN U19635 ( .B(n11466), .A(n11467), .Z(n11378) );
  XNOR U19636 ( .A(n11369), .B(n11468), .Z(n11374) );
  XNOR U19637 ( .A(n11367), .B(n11371), .Z(n11468) );
  AND U19638 ( .A(n11469), .B(n11470), .Z(n11371) );
  NAND U19639 ( .A(n11471), .B(n11472), .Z(n11470) );
  NAND U19640 ( .A(n11473), .B(n11474), .Z(n11469) );
  AND U19641 ( .A(n11475), .B(n11476), .Z(n11367) );
  NAND U19642 ( .A(n11477), .B(n11478), .Z(n11476) );
  NAND U19643 ( .A(n11479), .B(n11480), .Z(n11475) );
  AND U19644 ( .A(n11481), .B(n11482), .Z(n11369) );
  XOR U19645 ( .A(n11449), .B(n11448), .Z(N64375) );
  XNOR U19646 ( .A(n11466), .B(n11467), .Z(n11448) );
  XNOR U19647 ( .A(n11481), .B(n11482), .Z(n11467) );
  XOR U19648 ( .A(n11478), .B(n11477), .Z(n11482) );
  XOR U19649 ( .A(y[6996]), .B(x[6996]), .Z(n11477) );
  XOR U19650 ( .A(n11480), .B(n11479), .Z(n11478) );
  XOR U19651 ( .A(y[6998]), .B(x[6998]), .Z(n11479) );
  XOR U19652 ( .A(y[6997]), .B(x[6997]), .Z(n11480) );
  XOR U19653 ( .A(n11472), .B(n11471), .Z(n11481) );
  XOR U19654 ( .A(n11474), .B(n11473), .Z(n11471) );
  XOR U19655 ( .A(y[6995]), .B(x[6995]), .Z(n11473) );
  XOR U19656 ( .A(y[6994]), .B(x[6994]), .Z(n11474) );
  XOR U19657 ( .A(y[6993]), .B(x[6993]), .Z(n11472) );
  XNOR U19658 ( .A(n11465), .B(n11464), .Z(n11466) );
  XNOR U19659 ( .A(n11461), .B(n11460), .Z(n11464) );
  XOR U19660 ( .A(n11463), .B(n11462), .Z(n11460) );
  XOR U19661 ( .A(y[6992]), .B(x[6992]), .Z(n11462) );
  XOR U19662 ( .A(y[6991]), .B(x[6991]), .Z(n11463) );
  XOR U19663 ( .A(y[6990]), .B(x[6990]), .Z(n11461) );
  XOR U19664 ( .A(n11455), .B(n11454), .Z(n11465) );
  XOR U19665 ( .A(n11457), .B(n11456), .Z(n11454) );
  XOR U19666 ( .A(y[6989]), .B(x[6989]), .Z(n11456) );
  XOR U19667 ( .A(y[6988]), .B(x[6988]), .Z(n11457) );
  XOR U19668 ( .A(y[6987]), .B(x[6987]), .Z(n11455) );
  XNOR U19669 ( .A(n11431), .B(n11432), .Z(n11449) );
  XNOR U19670 ( .A(n11446), .B(n11447), .Z(n11432) );
  XOR U19671 ( .A(n11443), .B(n11442), .Z(n11447) );
  XOR U19672 ( .A(y[6984]), .B(x[6984]), .Z(n11442) );
  XOR U19673 ( .A(n11445), .B(n11444), .Z(n11443) );
  XOR U19674 ( .A(y[6986]), .B(x[6986]), .Z(n11444) );
  XOR U19675 ( .A(y[6985]), .B(x[6985]), .Z(n11445) );
  XOR U19676 ( .A(n11437), .B(n11436), .Z(n11446) );
  XOR U19677 ( .A(n11439), .B(n11438), .Z(n11436) );
  XOR U19678 ( .A(y[6983]), .B(x[6983]), .Z(n11438) );
  XOR U19679 ( .A(y[6982]), .B(x[6982]), .Z(n11439) );
  XOR U19680 ( .A(y[6981]), .B(x[6981]), .Z(n11437) );
  XNOR U19681 ( .A(n11430), .B(n11429), .Z(n11431) );
  XNOR U19682 ( .A(n11426), .B(n11425), .Z(n11429) );
  XOR U19683 ( .A(n11428), .B(n11427), .Z(n11425) );
  XOR U19684 ( .A(y[6980]), .B(x[6980]), .Z(n11427) );
  XOR U19685 ( .A(y[6979]), .B(x[6979]), .Z(n11428) );
  XOR U19686 ( .A(y[6978]), .B(x[6978]), .Z(n11426) );
  XOR U19687 ( .A(n11420), .B(n11419), .Z(n11430) );
  XOR U19688 ( .A(n11422), .B(n11421), .Z(n11419) );
  XOR U19689 ( .A(y[6977]), .B(x[6977]), .Z(n11421) );
  XOR U19690 ( .A(y[6976]), .B(x[6976]), .Z(n11422) );
  XOR U19691 ( .A(y[6975]), .B(x[6975]), .Z(n11420) );
  NAND U19692 ( .A(n11483), .B(n11484), .Z(N64366) );
  NAND U19693 ( .A(n11485), .B(n11486), .Z(n11484) );
  NANDN U19694 ( .A(n11487), .B(n11488), .Z(n11486) );
  NANDN U19695 ( .A(n11488), .B(n11487), .Z(n11483) );
  XOR U19696 ( .A(n11487), .B(n11489), .Z(N64365) );
  XNOR U19697 ( .A(n11485), .B(n11488), .Z(n11489) );
  NAND U19698 ( .A(n11490), .B(n11491), .Z(n11488) );
  NAND U19699 ( .A(n11492), .B(n11493), .Z(n11491) );
  NANDN U19700 ( .A(n11494), .B(n11495), .Z(n11493) );
  NANDN U19701 ( .A(n11495), .B(n11494), .Z(n11490) );
  AND U19702 ( .A(n11496), .B(n11497), .Z(n11485) );
  NAND U19703 ( .A(n11498), .B(n11499), .Z(n11497) );
  NANDN U19704 ( .A(n11500), .B(n11501), .Z(n11499) );
  NANDN U19705 ( .A(n11501), .B(n11500), .Z(n11496) );
  IV U19706 ( .A(n11502), .Z(n11501) );
  AND U19707 ( .A(n11503), .B(n11504), .Z(n11487) );
  NAND U19708 ( .A(n11505), .B(n11506), .Z(n11504) );
  NANDN U19709 ( .A(n11507), .B(n11508), .Z(n11506) );
  NANDN U19710 ( .A(n11508), .B(n11507), .Z(n11503) );
  XOR U19711 ( .A(n11500), .B(n11509), .Z(N64364) );
  XNOR U19712 ( .A(n11498), .B(n11502), .Z(n11509) );
  XOR U19713 ( .A(n11495), .B(n11510), .Z(n11502) );
  XNOR U19714 ( .A(n11492), .B(n11494), .Z(n11510) );
  AND U19715 ( .A(n11511), .B(n11512), .Z(n11494) );
  NANDN U19716 ( .A(n11513), .B(n11514), .Z(n11512) );
  OR U19717 ( .A(n11515), .B(n11516), .Z(n11514) );
  IV U19718 ( .A(n11517), .Z(n11516) );
  NANDN U19719 ( .A(n11517), .B(n11515), .Z(n11511) );
  AND U19720 ( .A(n11518), .B(n11519), .Z(n11492) );
  NAND U19721 ( .A(n11520), .B(n11521), .Z(n11519) );
  NANDN U19722 ( .A(n11522), .B(n11523), .Z(n11521) );
  NANDN U19723 ( .A(n11523), .B(n11522), .Z(n11518) );
  IV U19724 ( .A(n11524), .Z(n11523) );
  NAND U19725 ( .A(n11525), .B(n11526), .Z(n11495) );
  NANDN U19726 ( .A(n11527), .B(n11528), .Z(n11526) );
  NANDN U19727 ( .A(n11529), .B(n11530), .Z(n11528) );
  NANDN U19728 ( .A(n11530), .B(n11529), .Z(n11525) );
  IV U19729 ( .A(n11531), .Z(n11529) );
  AND U19730 ( .A(n11532), .B(n11533), .Z(n11498) );
  NAND U19731 ( .A(n11534), .B(n11535), .Z(n11533) );
  NANDN U19732 ( .A(n11536), .B(n11537), .Z(n11535) );
  NANDN U19733 ( .A(n11537), .B(n11536), .Z(n11532) );
  XOR U19734 ( .A(n11508), .B(n11538), .Z(n11500) );
  XNOR U19735 ( .A(n11505), .B(n11507), .Z(n11538) );
  AND U19736 ( .A(n11539), .B(n11540), .Z(n11507) );
  NANDN U19737 ( .A(n11541), .B(n11542), .Z(n11540) );
  OR U19738 ( .A(n11543), .B(n11544), .Z(n11542) );
  IV U19739 ( .A(n11545), .Z(n11544) );
  NANDN U19740 ( .A(n11545), .B(n11543), .Z(n11539) );
  AND U19741 ( .A(n11546), .B(n11547), .Z(n11505) );
  NAND U19742 ( .A(n11548), .B(n11549), .Z(n11547) );
  NANDN U19743 ( .A(n11550), .B(n11551), .Z(n11549) );
  NANDN U19744 ( .A(n11551), .B(n11550), .Z(n11546) );
  IV U19745 ( .A(n11552), .Z(n11551) );
  NAND U19746 ( .A(n11553), .B(n11554), .Z(n11508) );
  NANDN U19747 ( .A(n11555), .B(n11556), .Z(n11554) );
  NANDN U19748 ( .A(n11557), .B(n11558), .Z(n11556) );
  NANDN U19749 ( .A(n11558), .B(n11557), .Z(n11553) );
  IV U19750 ( .A(n11559), .Z(n11557) );
  XOR U19751 ( .A(n11534), .B(n11560), .Z(N64363) );
  XNOR U19752 ( .A(n11537), .B(n11536), .Z(n11560) );
  XNOR U19753 ( .A(n11548), .B(n11561), .Z(n11536) );
  XNOR U19754 ( .A(n11552), .B(n11550), .Z(n11561) );
  XOR U19755 ( .A(n11558), .B(n11562), .Z(n11550) );
  XNOR U19756 ( .A(n11555), .B(n11559), .Z(n11562) );
  AND U19757 ( .A(n11563), .B(n11564), .Z(n11559) );
  NAND U19758 ( .A(n11565), .B(n11566), .Z(n11564) );
  NAND U19759 ( .A(n11567), .B(n11568), .Z(n11563) );
  AND U19760 ( .A(n11569), .B(n11570), .Z(n11555) );
  NAND U19761 ( .A(n11571), .B(n11572), .Z(n11570) );
  NAND U19762 ( .A(n11573), .B(n11574), .Z(n11569) );
  NANDN U19763 ( .A(n11575), .B(n11576), .Z(n11558) );
  ANDN U19764 ( .B(n11577), .A(n11578), .Z(n11552) );
  XNOR U19765 ( .A(n11543), .B(n11579), .Z(n11548) );
  XNOR U19766 ( .A(n11541), .B(n11545), .Z(n11579) );
  AND U19767 ( .A(n11580), .B(n11581), .Z(n11545) );
  NAND U19768 ( .A(n11582), .B(n11583), .Z(n11581) );
  NAND U19769 ( .A(n11584), .B(n11585), .Z(n11580) );
  AND U19770 ( .A(n11586), .B(n11587), .Z(n11541) );
  NAND U19771 ( .A(n11588), .B(n11589), .Z(n11587) );
  NAND U19772 ( .A(n11590), .B(n11591), .Z(n11586) );
  AND U19773 ( .A(n11592), .B(n11593), .Z(n11543) );
  NAND U19774 ( .A(n11594), .B(n11595), .Z(n11537) );
  XNOR U19775 ( .A(n11520), .B(n11596), .Z(n11534) );
  XNOR U19776 ( .A(n11524), .B(n11522), .Z(n11596) );
  XOR U19777 ( .A(n11530), .B(n11597), .Z(n11522) );
  XNOR U19778 ( .A(n11527), .B(n11531), .Z(n11597) );
  AND U19779 ( .A(n11598), .B(n11599), .Z(n11531) );
  NAND U19780 ( .A(n11600), .B(n11601), .Z(n11599) );
  NAND U19781 ( .A(n11602), .B(n11603), .Z(n11598) );
  AND U19782 ( .A(n11604), .B(n11605), .Z(n11527) );
  NAND U19783 ( .A(n11606), .B(n11607), .Z(n11605) );
  NAND U19784 ( .A(n11608), .B(n11609), .Z(n11604) );
  NANDN U19785 ( .A(n11610), .B(n11611), .Z(n11530) );
  ANDN U19786 ( .B(n11612), .A(n11613), .Z(n11524) );
  XNOR U19787 ( .A(n11515), .B(n11614), .Z(n11520) );
  XNOR U19788 ( .A(n11513), .B(n11517), .Z(n11614) );
  AND U19789 ( .A(n11615), .B(n11616), .Z(n11517) );
  NAND U19790 ( .A(n11617), .B(n11618), .Z(n11616) );
  NAND U19791 ( .A(n11619), .B(n11620), .Z(n11615) );
  AND U19792 ( .A(n11621), .B(n11622), .Z(n11513) );
  NAND U19793 ( .A(n11623), .B(n11624), .Z(n11622) );
  NAND U19794 ( .A(n11625), .B(n11626), .Z(n11621) );
  AND U19795 ( .A(n11627), .B(n11628), .Z(n11515) );
  XOR U19796 ( .A(n11595), .B(n11594), .Z(N64362) );
  XNOR U19797 ( .A(n11612), .B(n11613), .Z(n11594) );
  XNOR U19798 ( .A(n11627), .B(n11628), .Z(n11613) );
  XOR U19799 ( .A(n11624), .B(n11623), .Z(n11628) );
  XOR U19800 ( .A(y[6972]), .B(x[6972]), .Z(n11623) );
  XOR U19801 ( .A(n11626), .B(n11625), .Z(n11624) );
  XOR U19802 ( .A(y[6974]), .B(x[6974]), .Z(n11625) );
  XOR U19803 ( .A(y[6973]), .B(x[6973]), .Z(n11626) );
  XOR U19804 ( .A(n11618), .B(n11617), .Z(n11627) );
  XOR U19805 ( .A(n11620), .B(n11619), .Z(n11617) );
  XOR U19806 ( .A(y[6971]), .B(x[6971]), .Z(n11619) );
  XOR U19807 ( .A(y[6970]), .B(x[6970]), .Z(n11620) );
  XOR U19808 ( .A(y[6969]), .B(x[6969]), .Z(n11618) );
  XNOR U19809 ( .A(n11611), .B(n11610), .Z(n11612) );
  XNOR U19810 ( .A(n11607), .B(n11606), .Z(n11610) );
  XOR U19811 ( .A(n11609), .B(n11608), .Z(n11606) );
  XOR U19812 ( .A(y[6968]), .B(x[6968]), .Z(n11608) );
  XOR U19813 ( .A(y[6967]), .B(x[6967]), .Z(n11609) );
  XOR U19814 ( .A(y[6966]), .B(x[6966]), .Z(n11607) );
  XOR U19815 ( .A(n11601), .B(n11600), .Z(n11611) );
  XOR U19816 ( .A(n11603), .B(n11602), .Z(n11600) );
  XOR U19817 ( .A(y[6965]), .B(x[6965]), .Z(n11602) );
  XOR U19818 ( .A(y[6964]), .B(x[6964]), .Z(n11603) );
  XOR U19819 ( .A(y[6963]), .B(x[6963]), .Z(n11601) );
  XNOR U19820 ( .A(n11577), .B(n11578), .Z(n11595) );
  XNOR U19821 ( .A(n11592), .B(n11593), .Z(n11578) );
  XOR U19822 ( .A(n11589), .B(n11588), .Z(n11593) );
  XOR U19823 ( .A(y[6960]), .B(x[6960]), .Z(n11588) );
  XOR U19824 ( .A(n11591), .B(n11590), .Z(n11589) );
  XOR U19825 ( .A(y[6962]), .B(x[6962]), .Z(n11590) );
  XOR U19826 ( .A(y[6961]), .B(x[6961]), .Z(n11591) );
  XOR U19827 ( .A(n11583), .B(n11582), .Z(n11592) );
  XOR U19828 ( .A(n11585), .B(n11584), .Z(n11582) );
  XOR U19829 ( .A(y[6959]), .B(x[6959]), .Z(n11584) );
  XOR U19830 ( .A(y[6958]), .B(x[6958]), .Z(n11585) );
  XOR U19831 ( .A(y[6957]), .B(x[6957]), .Z(n11583) );
  XNOR U19832 ( .A(n11576), .B(n11575), .Z(n11577) );
  XNOR U19833 ( .A(n11572), .B(n11571), .Z(n11575) );
  XOR U19834 ( .A(n11574), .B(n11573), .Z(n11571) );
  XOR U19835 ( .A(y[6956]), .B(x[6956]), .Z(n11573) );
  XOR U19836 ( .A(y[6955]), .B(x[6955]), .Z(n11574) );
  XOR U19837 ( .A(y[6954]), .B(x[6954]), .Z(n11572) );
  XOR U19838 ( .A(n11566), .B(n11565), .Z(n11576) );
  XOR U19839 ( .A(n11568), .B(n11567), .Z(n11565) );
  XOR U19840 ( .A(y[6953]), .B(x[6953]), .Z(n11567) );
  XOR U19841 ( .A(y[6952]), .B(x[6952]), .Z(n11568) );
  XOR U19842 ( .A(y[6951]), .B(x[6951]), .Z(n11566) );
  NAND U19843 ( .A(n11629), .B(n11630), .Z(N64353) );
  NAND U19844 ( .A(n11631), .B(n11632), .Z(n11630) );
  NANDN U19845 ( .A(n11633), .B(n11634), .Z(n11632) );
  NANDN U19846 ( .A(n11634), .B(n11633), .Z(n11629) );
  XOR U19847 ( .A(n11633), .B(n11635), .Z(N64352) );
  XNOR U19848 ( .A(n11631), .B(n11634), .Z(n11635) );
  NAND U19849 ( .A(n11636), .B(n11637), .Z(n11634) );
  NAND U19850 ( .A(n11638), .B(n11639), .Z(n11637) );
  NANDN U19851 ( .A(n11640), .B(n11641), .Z(n11639) );
  NANDN U19852 ( .A(n11641), .B(n11640), .Z(n11636) );
  AND U19853 ( .A(n11642), .B(n11643), .Z(n11631) );
  NAND U19854 ( .A(n11644), .B(n11645), .Z(n11643) );
  NANDN U19855 ( .A(n11646), .B(n11647), .Z(n11645) );
  NANDN U19856 ( .A(n11647), .B(n11646), .Z(n11642) );
  IV U19857 ( .A(n11648), .Z(n11647) );
  AND U19858 ( .A(n11649), .B(n11650), .Z(n11633) );
  NAND U19859 ( .A(n11651), .B(n11652), .Z(n11650) );
  NANDN U19860 ( .A(n11653), .B(n11654), .Z(n11652) );
  NANDN U19861 ( .A(n11654), .B(n11653), .Z(n11649) );
  XOR U19862 ( .A(n11646), .B(n11655), .Z(N64351) );
  XNOR U19863 ( .A(n11644), .B(n11648), .Z(n11655) );
  XOR U19864 ( .A(n11641), .B(n11656), .Z(n11648) );
  XNOR U19865 ( .A(n11638), .B(n11640), .Z(n11656) );
  AND U19866 ( .A(n11657), .B(n11658), .Z(n11640) );
  NANDN U19867 ( .A(n11659), .B(n11660), .Z(n11658) );
  OR U19868 ( .A(n11661), .B(n11662), .Z(n11660) );
  IV U19869 ( .A(n11663), .Z(n11662) );
  NANDN U19870 ( .A(n11663), .B(n11661), .Z(n11657) );
  AND U19871 ( .A(n11664), .B(n11665), .Z(n11638) );
  NAND U19872 ( .A(n11666), .B(n11667), .Z(n11665) );
  NANDN U19873 ( .A(n11668), .B(n11669), .Z(n11667) );
  NANDN U19874 ( .A(n11669), .B(n11668), .Z(n11664) );
  IV U19875 ( .A(n11670), .Z(n11669) );
  NAND U19876 ( .A(n11671), .B(n11672), .Z(n11641) );
  NANDN U19877 ( .A(n11673), .B(n11674), .Z(n11672) );
  NANDN U19878 ( .A(n11675), .B(n11676), .Z(n11674) );
  NANDN U19879 ( .A(n11676), .B(n11675), .Z(n11671) );
  IV U19880 ( .A(n11677), .Z(n11675) );
  AND U19881 ( .A(n11678), .B(n11679), .Z(n11644) );
  NAND U19882 ( .A(n11680), .B(n11681), .Z(n11679) );
  NANDN U19883 ( .A(n11682), .B(n11683), .Z(n11681) );
  NANDN U19884 ( .A(n11683), .B(n11682), .Z(n11678) );
  XOR U19885 ( .A(n11654), .B(n11684), .Z(n11646) );
  XNOR U19886 ( .A(n11651), .B(n11653), .Z(n11684) );
  AND U19887 ( .A(n11685), .B(n11686), .Z(n11653) );
  NANDN U19888 ( .A(n11687), .B(n11688), .Z(n11686) );
  OR U19889 ( .A(n11689), .B(n11690), .Z(n11688) );
  IV U19890 ( .A(n11691), .Z(n11690) );
  NANDN U19891 ( .A(n11691), .B(n11689), .Z(n11685) );
  AND U19892 ( .A(n11692), .B(n11693), .Z(n11651) );
  NAND U19893 ( .A(n11694), .B(n11695), .Z(n11693) );
  NANDN U19894 ( .A(n11696), .B(n11697), .Z(n11695) );
  NANDN U19895 ( .A(n11697), .B(n11696), .Z(n11692) );
  IV U19896 ( .A(n11698), .Z(n11697) );
  NAND U19897 ( .A(n11699), .B(n11700), .Z(n11654) );
  NANDN U19898 ( .A(n11701), .B(n11702), .Z(n11700) );
  NANDN U19899 ( .A(n11703), .B(n11704), .Z(n11702) );
  NANDN U19900 ( .A(n11704), .B(n11703), .Z(n11699) );
  IV U19901 ( .A(n11705), .Z(n11703) );
  XOR U19902 ( .A(n11680), .B(n11706), .Z(N64350) );
  XNOR U19903 ( .A(n11683), .B(n11682), .Z(n11706) );
  XNOR U19904 ( .A(n11694), .B(n11707), .Z(n11682) );
  XNOR U19905 ( .A(n11698), .B(n11696), .Z(n11707) );
  XOR U19906 ( .A(n11704), .B(n11708), .Z(n11696) );
  XNOR U19907 ( .A(n11701), .B(n11705), .Z(n11708) );
  AND U19908 ( .A(n11709), .B(n11710), .Z(n11705) );
  NAND U19909 ( .A(n11711), .B(n11712), .Z(n11710) );
  NAND U19910 ( .A(n11713), .B(n11714), .Z(n11709) );
  AND U19911 ( .A(n11715), .B(n11716), .Z(n11701) );
  NAND U19912 ( .A(n11717), .B(n11718), .Z(n11716) );
  NAND U19913 ( .A(n11719), .B(n11720), .Z(n11715) );
  NANDN U19914 ( .A(n11721), .B(n11722), .Z(n11704) );
  ANDN U19915 ( .B(n11723), .A(n11724), .Z(n11698) );
  XNOR U19916 ( .A(n11689), .B(n11725), .Z(n11694) );
  XNOR U19917 ( .A(n11687), .B(n11691), .Z(n11725) );
  AND U19918 ( .A(n11726), .B(n11727), .Z(n11691) );
  NAND U19919 ( .A(n11728), .B(n11729), .Z(n11727) );
  NAND U19920 ( .A(n11730), .B(n11731), .Z(n11726) );
  AND U19921 ( .A(n11732), .B(n11733), .Z(n11687) );
  NAND U19922 ( .A(n11734), .B(n11735), .Z(n11733) );
  NAND U19923 ( .A(n11736), .B(n11737), .Z(n11732) );
  AND U19924 ( .A(n11738), .B(n11739), .Z(n11689) );
  NAND U19925 ( .A(n11740), .B(n11741), .Z(n11683) );
  XNOR U19926 ( .A(n11666), .B(n11742), .Z(n11680) );
  XNOR U19927 ( .A(n11670), .B(n11668), .Z(n11742) );
  XOR U19928 ( .A(n11676), .B(n11743), .Z(n11668) );
  XNOR U19929 ( .A(n11673), .B(n11677), .Z(n11743) );
  AND U19930 ( .A(n11744), .B(n11745), .Z(n11677) );
  NAND U19931 ( .A(n11746), .B(n11747), .Z(n11745) );
  NAND U19932 ( .A(n11748), .B(n11749), .Z(n11744) );
  AND U19933 ( .A(n11750), .B(n11751), .Z(n11673) );
  NAND U19934 ( .A(n11752), .B(n11753), .Z(n11751) );
  NAND U19935 ( .A(n11754), .B(n11755), .Z(n11750) );
  NANDN U19936 ( .A(n11756), .B(n11757), .Z(n11676) );
  ANDN U19937 ( .B(n11758), .A(n11759), .Z(n11670) );
  XNOR U19938 ( .A(n11661), .B(n11760), .Z(n11666) );
  XNOR U19939 ( .A(n11659), .B(n11663), .Z(n11760) );
  AND U19940 ( .A(n11761), .B(n11762), .Z(n11663) );
  NAND U19941 ( .A(n11763), .B(n11764), .Z(n11762) );
  NAND U19942 ( .A(n11765), .B(n11766), .Z(n11761) );
  AND U19943 ( .A(n11767), .B(n11768), .Z(n11659) );
  NAND U19944 ( .A(n11769), .B(n11770), .Z(n11768) );
  NAND U19945 ( .A(n11771), .B(n11772), .Z(n11767) );
  AND U19946 ( .A(n11773), .B(n11774), .Z(n11661) );
  XOR U19947 ( .A(n11741), .B(n11740), .Z(N64349) );
  XNOR U19948 ( .A(n11758), .B(n11759), .Z(n11740) );
  XNOR U19949 ( .A(n11773), .B(n11774), .Z(n11759) );
  XOR U19950 ( .A(n11770), .B(n11769), .Z(n11774) );
  XOR U19951 ( .A(y[6948]), .B(x[6948]), .Z(n11769) );
  XOR U19952 ( .A(n11772), .B(n11771), .Z(n11770) );
  XOR U19953 ( .A(y[6950]), .B(x[6950]), .Z(n11771) );
  XOR U19954 ( .A(y[6949]), .B(x[6949]), .Z(n11772) );
  XOR U19955 ( .A(n11764), .B(n11763), .Z(n11773) );
  XOR U19956 ( .A(n11766), .B(n11765), .Z(n11763) );
  XOR U19957 ( .A(y[6947]), .B(x[6947]), .Z(n11765) );
  XOR U19958 ( .A(y[6946]), .B(x[6946]), .Z(n11766) );
  XOR U19959 ( .A(y[6945]), .B(x[6945]), .Z(n11764) );
  XNOR U19960 ( .A(n11757), .B(n11756), .Z(n11758) );
  XNOR U19961 ( .A(n11753), .B(n11752), .Z(n11756) );
  XOR U19962 ( .A(n11755), .B(n11754), .Z(n11752) );
  XOR U19963 ( .A(y[6944]), .B(x[6944]), .Z(n11754) );
  XOR U19964 ( .A(y[6943]), .B(x[6943]), .Z(n11755) );
  XOR U19965 ( .A(y[6942]), .B(x[6942]), .Z(n11753) );
  XOR U19966 ( .A(n11747), .B(n11746), .Z(n11757) );
  XOR U19967 ( .A(n11749), .B(n11748), .Z(n11746) );
  XOR U19968 ( .A(y[6941]), .B(x[6941]), .Z(n11748) );
  XOR U19969 ( .A(y[6940]), .B(x[6940]), .Z(n11749) );
  XOR U19970 ( .A(y[6939]), .B(x[6939]), .Z(n11747) );
  XNOR U19971 ( .A(n11723), .B(n11724), .Z(n11741) );
  XNOR U19972 ( .A(n11738), .B(n11739), .Z(n11724) );
  XOR U19973 ( .A(n11735), .B(n11734), .Z(n11739) );
  XOR U19974 ( .A(y[6936]), .B(x[6936]), .Z(n11734) );
  XOR U19975 ( .A(n11737), .B(n11736), .Z(n11735) );
  XOR U19976 ( .A(y[6938]), .B(x[6938]), .Z(n11736) );
  XOR U19977 ( .A(y[6937]), .B(x[6937]), .Z(n11737) );
  XOR U19978 ( .A(n11729), .B(n11728), .Z(n11738) );
  XOR U19979 ( .A(n11731), .B(n11730), .Z(n11728) );
  XOR U19980 ( .A(y[6935]), .B(x[6935]), .Z(n11730) );
  XOR U19981 ( .A(y[6934]), .B(x[6934]), .Z(n11731) );
  XOR U19982 ( .A(y[6933]), .B(x[6933]), .Z(n11729) );
  XNOR U19983 ( .A(n11722), .B(n11721), .Z(n11723) );
  XNOR U19984 ( .A(n11718), .B(n11717), .Z(n11721) );
  XOR U19985 ( .A(n11720), .B(n11719), .Z(n11717) );
  XOR U19986 ( .A(y[6932]), .B(x[6932]), .Z(n11719) );
  XOR U19987 ( .A(y[6931]), .B(x[6931]), .Z(n11720) );
  XOR U19988 ( .A(y[6930]), .B(x[6930]), .Z(n11718) );
  XOR U19989 ( .A(n11712), .B(n11711), .Z(n11722) );
  XOR U19990 ( .A(n11714), .B(n11713), .Z(n11711) );
  XOR U19991 ( .A(y[6929]), .B(x[6929]), .Z(n11713) );
  XOR U19992 ( .A(y[6928]), .B(x[6928]), .Z(n11714) );
  XOR U19993 ( .A(y[6927]), .B(x[6927]), .Z(n11712) );
  NAND U19994 ( .A(n11775), .B(n11776), .Z(N64340) );
  NAND U19995 ( .A(n11777), .B(n11778), .Z(n11776) );
  NANDN U19996 ( .A(n11779), .B(n11780), .Z(n11778) );
  NANDN U19997 ( .A(n11780), .B(n11779), .Z(n11775) );
  XOR U19998 ( .A(n11779), .B(n11781), .Z(N64339) );
  XNOR U19999 ( .A(n11777), .B(n11780), .Z(n11781) );
  NAND U20000 ( .A(n11782), .B(n11783), .Z(n11780) );
  NAND U20001 ( .A(n11784), .B(n11785), .Z(n11783) );
  NANDN U20002 ( .A(n11786), .B(n11787), .Z(n11785) );
  NANDN U20003 ( .A(n11787), .B(n11786), .Z(n11782) );
  AND U20004 ( .A(n11788), .B(n11789), .Z(n11777) );
  NAND U20005 ( .A(n11790), .B(n11791), .Z(n11789) );
  NANDN U20006 ( .A(n11792), .B(n11793), .Z(n11791) );
  NANDN U20007 ( .A(n11793), .B(n11792), .Z(n11788) );
  IV U20008 ( .A(n11794), .Z(n11793) );
  AND U20009 ( .A(n11795), .B(n11796), .Z(n11779) );
  NAND U20010 ( .A(n11797), .B(n11798), .Z(n11796) );
  NANDN U20011 ( .A(n11799), .B(n11800), .Z(n11798) );
  NANDN U20012 ( .A(n11800), .B(n11799), .Z(n11795) );
  XOR U20013 ( .A(n11792), .B(n11801), .Z(N64338) );
  XNOR U20014 ( .A(n11790), .B(n11794), .Z(n11801) );
  XOR U20015 ( .A(n11787), .B(n11802), .Z(n11794) );
  XNOR U20016 ( .A(n11784), .B(n11786), .Z(n11802) );
  AND U20017 ( .A(n11803), .B(n11804), .Z(n11786) );
  NANDN U20018 ( .A(n11805), .B(n11806), .Z(n11804) );
  OR U20019 ( .A(n11807), .B(n11808), .Z(n11806) );
  IV U20020 ( .A(n11809), .Z(n11808) );
  NANDN U20021 ( .A(n11809), .B(n11807), .Z(n11803) );
  AND U20022 ( .A(n11810), .B(n11811), .Z(n11784) );
  NAND U20023 ( .A(n11812), .B(n11813), .Z(n11811) );
  NANDN U20024 ( .A(n11814), .B(n11815), .Z(n11813) );
  NANDN U20025 ( .A(n11815), .B(n11814), .Z(n11810) );
  IV U20026 ( .A(n11816), .Z(n11815) );
  NAND U20027 ( .A(n11817), .B(n11818), .Z(n11787) );
  NANDN U20028 ( .A(n11819), .B(n11820), .Z(n11818) );
  NANDN U20029 ( .A(n11821), .B(n11822), .Z(n11820) );
  NANDN U20030 ( .A(n11822), .B(n11821), .Z(n11817) );
  IV U20031 ( .A(n11823), .Z(n11821) );
  AND U20032 ( .A(n11824), .B(n11825), .Z(n11790) );
  NAND U20033 ( .A(n11826), .B(n11827), .Z(n11825) );
  NANDN U20034 ( .A(n11828), .B(n11829), .Z(n11827) );
  NANDN U20035 ( .A(n11829), .B(n11828), .Z(n11824) );
  XOR U20036 ( .A(n11800), .B(n11830), .Z(n11792) );
  XNOR U20037 ( .A(n11797), .B(n11799), .Z(n11830) );
  AND U20038 ( .A(n11831), .B(n11832), .Z(n11799) );
  NANDN U20039 ( .A(n11833), .B(n11834), .Z(n11832) );
  OR U20040 ( .A(n11835), .B(n11836), .Z(n11834) );
  IV U20041 ( .A(n11837), .Z(n11836) );
  NANDN U20042 ( .A(n11837), .B(n11835), .Z(n11831) );
  AND U20043 ( .A(n11838), .B(n11839), .Z(n11797) );
  NAND U20044 ( .A(n11840), .B(n11841), .Z(n11839) );
  NANDN U20045 ( .A(n11842), .B(n11843), .Z(n11841) );
  NANDN U20046 ( .A(n11843), .B(n11842), .Z(n11838) );
  IV U20047 ( .A(n11844), .Z(n11843) );
  NAND U20048 ( .A(n11845), .B(n11846), .Z(n11800) );
  NANDN U20049 ( .A(n11847), .B(n11848), .Z(n11846) );
  NANDN U20050 ( .A(n11849), .B(n11850), .Z(n11848) );
  NANDN U20051 ( .A(n11850), .B(n11849), .Z(n11845) );
  IV U20052 ( .A(n11851), .Z(n11849) );
  XOR U20053 ( .A(n11826), .B(n11852), .Z(N64337) );
  XNOR U20054 ( .A(n11829), .B(n11828), .Z(n11852) );
  XNOR U20055 ( .A(n11840), .B(n11853), .Z(n11828) );
  XNOR U20056 ( .A(n11844), .B(n11842), .Z(n11853) );
  XOR U20057 ( .A(n11850), .B(n11854), .Z(n11842) );
  XNOR U20058 ( .A(n11847), .B(n11851), .Z(n11854) );
  AND U20059 ( .A(n11855), .B(n11856), .Z(n11851) );
  NAND U20060 ( .A(n11857), .B(n11858), .Z(n11856) );
  NAND U20061 ( .A(n11859), .B(n11860), .Z(n11855) );
  AND U20062 ( .A(n11861), .B(n11862), .Z(n11847) );
  NAND U20063 ( .A(n11863), .B(n11864), .Z(n11862) );
  NAND U20064 ( .A(n11865), .B(n11866), .Z(n11861) );
  NANDN U20065 ( .A(n11867), .B(n11868), .Z(n11850) );
  ANDN U20066 ( .B(n11869), .A(n11870), .Z(n11844) );
  XNOR U20067 ( .A(n11835), .B(n11871), .Z(n11840) );
  XNOR U20068 ( .A(n11833), .B(n11837), .Z(n11871) );
  AND U20069 ( .A(n11872), .B(n11873), .Z(n11837) );
  NAND U20070 ( .A(n11874), .B(n11875), .Z(n11873) );
  NAND U20071 ( .A(n11876), .B(n11877), .Z(n11872) );
  AND U20072 ( .A(n11878), .B(n11879), .Z(n11833) );
  NAND U20073 ( .A(n11880), .B(n11881), .Z(n11879) );
  NAND U20074 ( .A(n11882), .B(n11883), .Z(n11878) );
  AND U20075 ( .A(n11884), .B(n11885), .Z(n11835) );
  NAND U20076 ( .A(n11886), .B(n11887), .Z(n11829) );
  XNOR U20077 ( .A(n11812), .B(n11888), .Z(n11826) );
  XNOR U20078 ( .A(n11816), .B(n11814), .Z(n11888) );
  XOR U20079 ( .A(n11822), .B(n11889), .Z(n11814) );
  XNOR U20080 ( .A(n11819), .B(n11823), .Z(n11889) );
  AND U20081 ( .A(n11890), .B(n11891), .Z(n11823) );
  NAND U20082 ( .A(n11892), .B(n11893), .Z(n11891) );
  NAND U20083 ( .A(n11894), .B(n11895), .Z(n11890) );
  AND U20084 ( .A(n11896), .B(n11897), .Z(n11819) );
  NAND U20085 ( .A(n11898), .B(n11899), .Z(n11897) );
  NAND U20086 ( .A(n11900), .B(n11901), .Z(n11896) );
  NANDN U20087 ( .A(n11902), .B(n11903), .Z(n11822) );
  ANDN U20088 ( .B(n11904), .A(n11905), .Z(n11816) );
  XNOR U20089 ( .A(n11807), .B(n11906), .Z(n11812) );
  XNOR U20090 ( .A(n11805), .B(n11809), .Z(n11906) );
  AND U20091 ( .A(n11907), .B(n11908), .Z(n11809) );
  NAND U20092 ( .A(n11909), .B(n11910), .Z(n11908) );
  NAND U20093 ( .A(n11911), .B(n11912), .Z(n11907) );
  AND U20094 ( .A(n11913), .B(n11914), .Z(n11805) );
  NAND U20095 ( .A(n11915), .B(n11916), .Z(n11914) );
  NAND U20096 ( .A(n11917), .B(n11918), .Z(n11913) );
  AND U20097 ( .A(n11919), .B(n11920), .Z(n11807) );
  XOR U20098 ( .A(n11887), .B(n11886), .Z(N64336) );
  XNOR U20099 ( .A(n11904), .B(n11905), .Z(n11886) );
  XNOR U20100 ( .A(n11919), .B(n11920), .Z(n11905) );
  XOR U20101 ( .A(n11916), .B(n11915), .Z(n11920) );
  XOR U20102 ( .A(y[6924]), .B(x[6924]), .Z(n11915) );
  XOR U20103 ( .A(n11918), .B(n11917), .Z(n11916) );
  XOR U20104 ( .A(y[6926]), .B(x[6926]), .Z(n11917) );
  XOR U20105 ( .A(y[6925]), .B(x[6925]), .Z(n11918) );
  XOR U20106 ( .A(n11910), .B(n11909), .Z(n11919) );
  XOR U20107 ( .A(n11912), .B(n11911), .Z(n11909) );
  XOR U20108 ( .A(y[6923]), .B(x[6923]), .Z(n11911) );
  XOR U20109 ( .A(y[6922]), .B(x[6922]), .Z(n11912) );
  XOR U20110 ( .A(y[6921]), .B(x[6921]), .Z(n11910) );
  XNOR U20111 ( .A(n11903), .B(n11902), .Z(n11904) );
  XNOR U20112 ( .A(n11899), .B(n11898), .Z(n11902) );
  XOR U20113 ( .A(n11901), .B(n11900), .Z(n11898) );
  XOR U20114 ( .A(y[6920]), .B(x[6920]), .Z(n11900) );
  XOR U20115 ( .A(y[6919]), .B(x[6919]), .Z(n11901) );
  XOR U20116 ( .A(y[6918]), .B(x[6918]), .Z(n11899) );
  XOR U20117 ( .A(n11893), .B(n11892), .Z(n11903) );
  XOR U20118 ( .A(n11895), .B(n11894), .Z(n11892) );
  XOR U20119 ( .A(y[6917]), .B(x[6917]), .Z(n11894) );
  XOR U20120 ( .A(y[6916]), .B(x[6916]), .Z(n11895) );
  XOR U20121 ( .A(y[6915]), .B(x[6915]), .Z(n11893) );
  XNOR U20122 ( .A(n11869), .B(n11870), .Z(n11887) );
  XNOR U20123 ( .A(n11884), .B(n11885), .Z(n11870) );
  XOR U20124 ( .A(n11881), .B(n11880), .Z(n11885) );
  XOR U20125 ( .A(y[6912]), .B(x[6912]), .Z(n11880) );
  XOR U20126 ( .A(n11883), .B(n11882), .Z(n11881) );
  XOR U20127 ( .A(y[6914]), .B(x[6914]), .Z(n11882) );
  XOR U20128 ( .A(y[6913]), .B(x[6913]), .Z(n11883) );
  XOR U20129 ( .A(n11875), .B(n11874), .Z(n11884) );
  XOR U20130 ( .A(n11877), .B(n11876), .Z(n11874) );
  XOR U20131 ( .A(y[6911]), .B(x[6911]), .Z(n11876) );
  XOR U20132 ( .A(y[6910]), .B(x[6910]), .Z(n11877) );
  XOR U20133 ( .A(y[6909]), .B(x[6909]), .Z(n11875) );
  XNOR U20134 ( .A(n11868), .B(n11867), .Z(n11869) );
  XNOR U20135 ( .A(n11864), .B(n11863), .Z(n11867) );
  XOR U20136 ( .A(n11866), .B(n11865), .Z(n11863) );
  XOR U20137 ( .A(y[6908]), .B(x[6908]), .Z(n11865) );
  XOR U20138 ( .A(y[6907]), .B(x[6907]), .Z(n11866) );
  XOR U20139 ( .A(y[6906]), .B(x[6906]), .Z(n11864) );
  XOR U20140 ( .A(n11858), .B(n11857), .Z(n11868) );
  XOR U20141 ( .A(n11860), .B(n11859), .Z(n11857) );
  XOR U20142 ( .A(y[6905]), .B(x[6905]), .Z(n11859) );
  XOR U20143 ( .A(y[6904]), .B(x[6904]), .Z(n11860) );
  XOR U20144 ( .A(y[6903]), .B(x[6903]), .Z(n11858) );
  NAND U20145 ( .A(n11921), .B(n11922), .Z(N64327) );
  NAND U20146 ( .A(n11923), .B(n11924), .Z(n11922) );
  NANDN U20147 ( .A(n11925), .B(n11926), .Z(n11924) );
  NANDN U20148 ( .A(n11926), .B(n11925), .Z(n11921) );
  XOR U20149 ( .A(n11925), .B(n11927), .Z(N64326) );
  XNOR U20150 ( .A(n11923), .B(n11926), .Z(n11927) );
  NAND U20151 ( .A(n11928), .B(n11929), .Z(n11926) );
  NAND U20152 ( .A(n11930), .B(n11931), .Z(n11929) );
  NANDN U20153 ( .A(n11932), .B(n11933), .Z(n11931) );
  NANDN U20154 ( .A(n11933), .B(n11932), .Z(n11928) );
  AND U20155 ( .A(n11934), .B(n11935), .Z(n11923) );
  NAND U20156 ( .A(n11936), .B(n11937), .Z(n11935) );
  NANDN U20157 ( .A(n11938), .B(n11939), .Z(n11937) );
  NANDN U20158 ( .A(n11939), .B(n11938), .Z(n11934) );
  IV U20159 ( .A(n11940), .Z(n11939) );
  AND U20160 ( .A(n11941), .B(n11942), .Z(n11925) );
  NAND U20161 ( .A(n11943), .B(n11944), .Z(n11942) );
  NANDN U20162 ( .A(n11945), .B(n11946), .Z(n11944) );
  NANDN U20163 ( .A(n11946), .B(n11945), .Z(n11941) );
  XOR U20164 ( .A(n11938), .B(n11947), .Z(N64325) );
  XNOR U20165 ( .A(n11936), .B(n11940), .Z(n11947) );
  XOR U20166 ( .A(n11933), .B(n11948), .Z(n11940) );
  XNOR U20167 ( .A(n11930), .B(n11932), .Z(n11948) );
  AND U20168 ( .A(n11949), .B(n11950), .Z(n11932) );
  NANDN U20169 ( .A(n11951), .B(n11952), .Z(n11950) );
  OR U20170 ( .A(n11953), .B(n11954), .Z(n11952) );
  IV U20171 ( .A(n11955), .Z(n11954) );
  NANDN U20172 ( .A(n11955), .B(n11953), .Z(n11949) );
  AND U20173 ( .A(n11956), .B(n11957), .Z(n11930) );
  NAND U20174 ( .A(n11958), .B(n11959), .Z(n11957) );
  NANDN U20175 ( .A(n11960), .B(n11961), .Z(n11959) );
  NANDN U20176 ( .A(n11961), .B(n11960), .Z(n11956) );
  IV U20177 ( .A(n11962), .Z(n11961) );
  NAND U20178 ( .A(n11963), .B(n11964), .Z(n11933) );
  NANDN U20179 ( .A(n11965), .B(n11966), .Z(n11964) );
  NANDN U20180 ( .A(n11967), .B(n11968), .Z(n11966) );
  NANDN U20181 ( .A(n11968), .B(n11967), .Z(n11963) );
  IV U20182 ( .A(n11969), .Z(n11967) );
  AND U20183 ( .A(n11970), .B(n11971), .Z(n11936) );
  NAND U20184 ( .A(n11972), .B(n11973), .Z(n11971) );
  NANDN U20185 ( .A(n11974), .B(n11975), .Z(n11973) );
  NANDN U20186 ( .A(n11975), .B(n11974), .Z(n11970) );
  XOR U20187 ( .A(n11946), .B(n11976), .Z(n11938) );
  XNOR U20188 ( .A(n11943), .B(n11945), .Z(n11976) );
  AND U20189 ( .A(n11977), .B(n11978), .Z(n11945) );
  NANDN U20190 ( .A(n11979), .B(n11980), .Z(n11978) );
  OR U20191 ( .A(n11981), .B(n11982), .Z(n11980) );
  IV U20192 ( .A(n11983), .Z(n11982) );
  NANDN U20193 ( .A(n11983), .B(n11981), .Z(n11977) );
  AND U20194 ( .A(n11984), .B(n11985), .Z(n11943) );
  NAND U20195 ( .A(n11986), .B(n11987), .Z(n11985) );
  NANDN U20196 ( .A(n11988), .B(n11989), .Z(n11987) );
  NANDN U20197 ( .A(n11989), .B(n11988), .Z(n11984) );
  IV U20198 ( .A(n11990), .Z(n11989) );
  NAND U20199 ( .A(n11991), .B(n11992), .Z(n11946) );
  NANDN U20200 ( .A(n11993), .B(n11994), .Z(n11992) );
  NANDN U20201 ( .A(n11995), .B(n11996), .Z(n11994) );
  NANDN U20202 ( .A(n11996), .B(n11995), .Z(n11991) );
  IV U20203 ( .A(n11997), .Z(n11995) );
  XOR U20204 ( .A(n11972), .B(n11998), .Z(N64324) );
  XNOR U20205 ( .A(n11975), .B(n11974), .Z(n11998) );
  XNOR U20206 ( .A(n11986), .B(n11999), .Z(n11974) );
  XNOR U20207 ( .A(n11990), .B(n11988), .Z(n11999) );
  XOR U20208 ( .A(n11996), .B(n12000), .Z(n11988) );
  XNOR U20209 ( .A(n11993), .B(n11997), .Z(n12000) );
  AND U20210 ( .A(n12001), .B(n12002), .Z(n11997) );
  NAND U20211 ( .A(n12003), .B(n12004), .Z(n12002) );
  NAND U20212 ( .A(n12005), .B(n12006), .Z(n12001) );
  AND U20213 ( .A(n12007), .B(n12008), .Z(n11993) );
  NAND U20214 ( .A(n12009), .B(n12010), .Z(n12008) );
  NAND U20215 ( .A(n12011), .B(n12012), .Z(n12007) );
  NANDN U20216 ( .A(n12013), .B(n12014), .Z(n11996) );
  ANDN U20217 ( .B(n12015), .A(n12016), .Z(n11990) );
  XNOR U20218 ( .A(n11981), .B(n12017), .Z(n11986) );
  XNOR U20219 ( .A(n11979), .B(n11983), .Z(n12017) );
  AND U20220 ( .A(n12018), .B(n12019), .Z(n11983) );
  NAND U20221 ( .A(n12020), .B(n12021), .Z(n12019) );
  NAND U20222 ( .A(n12022), .B(n12023), .Z(n12018) );
  AND U20223 ( .A(n12024), .B(n12025), .Z(n11979) );
  NAND U20224 ( .A(n12026), .B(n12027), .Z(n12025) );
  NAND U20225 ( .A(n12028), .B(n12029), .Z(n12024) );
  AND U20226 ( .A(n12030), .B(n12031), .Z(n11981) );
  NAND U20227 ( .A(n12032), .B(n12033), .Z(n11975) );
  XNOR U20228 ( .A(n11958), .B(n12034), .Z(n11972) );
  XNOR U20229 ( .A(n11962), .B(n11960), .Z(n12034) );
  XOR U20230 ( .A(n11968), .B(n12035), .Z(n11960) );
  XNOR U20231 ( .A(n11965), .B(n11969), .Z(n12035) );
  AND U20232 ( .A(n12036), .B(n12037), .Z(n11969) );
  NAND U20233 ( .A(n12038), .B(n12039), .Z(n12037) );
  NAND U20234 ( .A(n12040), .B(n12041), .Z(n12036) );
  AND U20235 ( .A(n12042), .B(n12043), .Z(n11965) );
  NAND U20236 ( .A(n12044), .B(n12045), .Z(n12043) );
  NAND U20237 ( .A(n12046), .B(n12047), .Z(n12042) );
  NANDN U20238 ( .A(n12048), .B(n12049), .Z(n11968) );
  ANDN U20239 ( .B(n12050), .A(n12051), .Z(n11962) );
  XNOR U20240 ( .A(n11953), .B(n12052), .Z(n11958) );
  XNOR U20241 ( .A(n11951), .B(n11955), .Z(n12052) );
  AND U20242 ( .A(n12053), .B(n12054), .Z(n11955) );
  NAND U20243 ( .A(n12055), .B(n12056), .Z(n12054) );
  NAND U20244 ( .A(n12057), .B(n12058), .Z(n12053) );
  AND U20245 ( .A(n12059), .B(n12060), .Z(n11951) );
  NAND U20246 ( .A(n12061), .B(n12062), .Z(n12060) );
  NAND U20247 ( .A(n12063), .B(n12064), .Z(n12059) );
  AND U20248 ( .A(n12065), .B(n12066), .Z(n11953) );
  XOR U20249 ( .A(n12033), .B(n12032), .Z(N64323) );
  XNOR U20250 ( .A(n12050), .B(n12051), .Z(n12032) );
  XNOR U20251 ( .A(n12065), .B(n12066), .Z(n12051) );
  XOR U20252 ( .A(n12062), .B(n12061), .Z(n12066) );
  XOR U20253 ( .A(y[6900]), .B(x[6900]), .Z(n12061) );
  XOR U20254 ( .A(n12064), .B(n12063), .Z(n12062) );
  XOR U20255 ( .A(y[6902]), .B(x[6902]), .Z(n12063) );
  XOR U20256 ( .A(y[6901]), .B(x[6901]), .Z(n12064) );
  XOR U20257 ( .A(n12056), .B(n12055), .Z(n12065) );
  XOR U20258 ( .A(n12058), .B(n12057), .Z(n12055) );
  XOR U20259 ( .A(y[6899]), .B(x[6899]), .Z(n12057) );
  XOR U20260 ( .A(y[6898]), .B(x[6898]), .Z(n12058) );
  XOR U20261 ( .A(y[6897]), .B(x[6897]), .Z(n12056) );
  XNOR U20262 ( .A(n12049), .B(n12048), .Z(n12050) );
  XNOR U20263 ( .A(n12045), .B(n12044), .Z(n12048) );
  XOR U20264 ( .A(n12047), .B(n12046), .Z(n12044) );
  XOR U20265 ( .A(y[6896]), .B(x[6896]), .Z(n12046) );
  XOR U20266 ( .A(y[6895]), .B(x[6895]), .Z(n12047) );
  XOR U20267 ( .A(y[6894]), .B(x[6894]), .Z(n12045) );
  XOR U20268 ( .A(n12039), .B(n12038), .Z(n12049) );
  XOR U20269 ( .A(n12041), .B(n12040), .Z(n12038) );
  XOR U20270 ( .A(y[6893]), .B(x[6893]), .Z(n12040) );
  XOR U20271 ( .A(y[6892]), .B(x[6892]), .Z(n12041) );
  XOR U20272 ( .A(y[6891]), .B(x[6891]), .Z(n12039) );
  XNOR U20273 ( .A(n12015), .B(n12016), .Z(n12033) );
  XNOR U20274 ( .A(n12030), .B(n12031), .Z(n12016) );
  XOR U20275 ( .A(n12027), .B(n12026), .Z(n12031) );
  XOR U20276 ( .A(y[6888]), .B(x[6888]), .Z(n12026) );
  XOR U20277 ( .A(n12029), .B(n12028), .Z(n12027) );
  XOR U20278 ( .A(y[6890]), .B(x[6890]), .Z(n12028) );
  XOR U20279 ( .A(y[6889]), .B(x[6889]), .Z(n12029) );
  XOR U20280 ( .A(n12021), .B(n12020), .Z(n12030) );
  XOR U20281 ( .A(n12023), .B(n12022), .Z(n12020) );
  XOR U20282 ( .A(y[6887]), .B(x[6887]), .Z(n12022) );
  XOR U20283 ( .A(y[6886]), .B(x[6886]), .Z(n12023) );
  XOR U20284 ( .A(y[6885]), .B(x[6885]), .Z(n12021) );
  XNOR U20285 ( .A(n12014), .B(n12013), .Z(n12015) );
  XNOR U20286 ( .A(n12010), .B(n12009), .Z(n12013) );
  XOR U20287 ( .A(n12012), .B(n12011), .Z(n12009) );
  XOR U20288 ( .A(y[6884]), .B(x[6884]), .Z(n12011) );
  XOR U20289 ( .A(y[6883]), .B(x[6883]), .Z(n12012) );
  XOR U20290 ( .A(y[6882]), .B(x[6882]), .Z(n12010) );
  XOR U20291 ( .A(n12004), .B(n12003), .Z(n12014) );
  XOR U20292 ( .A(n12006), .B(n12005), .Z(n12003) );
  XOR U20293 ( .A(y[6881]), .B(x[6881]), .Z(n12005) );
  XOR U20294 ( .A(y[6880]), .B(x[6880]), .Z(n12006) );
  XOR U20295 ( .A(y[6879]), .B(x[6879]), .Z(n12004) );
  NAND U20296 ( .A(n12067), .B(n12068), .Z(N64314) );
  NAND U20297 ( .A(n12069), .B(n12070), .Z(n12068) );
  NANDN U20298 ( .A(n12071), .B(n12072), .Z(n12070) );
  NANDN U20299 ( .A(n12072), .B(n12071), .Z(n12067) );
  XOR U20300 ( .A(n12071), .B(n12073), .Z(N64313) );
  XNOR U20301 ( .A(n12069), .B(n12072), .Z(n12073) );
  NAND U20302 ( .A(n12074), .B(n12075), .Z(n12072) );
  NAND U20303 ( .A(n12076), .B(n12077), .Z(n12075) );
  NANDN U20304 ( .A(n12078), .B(n12079), .Z(n12077) );
  NANDN U20305 ( .A(n12079), .B(n12078), .Z(n12074) );
  AND U20306 ( .A(n12080), .B(n12081), .Z(n12069) );
  NAND U20307 ( .A(n12082), .B(n12083), .Z(n12081) );
  NANDN U20308 ( .A(n12084), .B(n12085), .Z(n12083) );
  NANDN U20309 ( .A(n12085), .B(n12084), .Z(n12080) );
  IV U20310 ( .A(n12086), .Z(n12085) );
  AND U20311 ( .A(n12087), .B(n12088), .Z(n12071) );
  NAND U20312 ( .A(n12089), .B(n12090), .Z(n12088) );
  NANDN U20313 ( .A(n12091), .B(n12092), .Z(n12090) );
  NANDN U20314 ( .A(n12092), .B(n12091), .Z(n12087) );
  XOR U20315 ( .A(n12084), .B(n12093), .Z(N64312) );
  XNOR U20316 ( .A(n12082), .B(n12086), .Z(n12093) );
  XOR U20317 ( .A(n12079), .B(n12094), .Z(n12086) );
  XNOR U20318 ( .A(n12076), .B(n12078), .Z(n12094) );
  AND U20319 ( .A(n12095), .B(n12096), .Z(n12078) );
  NANDN U20320 ( .A(n12097), .B(n12098), .Z(n12096) );
  OR U20321 ( .A(n12099), .B(n12100), .Z(n12098) );
  IV U20322 ( .A(n12101), .Z(n12100) );
  NANDN U20323 ( .A(n12101), .B(n12099), .Z(n12095) );
  AND U20324 ( .A(n12102), .B(n12103), .Z(n12076) );
  NAND U20325 ( .A(n12104), .B(n12105), .Z(n12103) );
  NANDN U20326 ( .A(n12106), .B(n12107), .Z(n12105) );
  NANDN U20327 ( .A(n12107), .B(n12106), .Z(n12102) );
  IV U20328 ( .A(n12108), .Z(n12107) );
  NAND U20329 ( .A(n12109), .B(n12110), .Z(n12079) );
  NANDN U20330 ( .A(n12111), .B(n12112), .Z(n12110) );
  NANDN U20331 ( .A(n12113), .B(n12114), .Z(n12112) );
  NANDN U20332 ( .A(n12114), .B(n12113), .Z(n12109) );
  IV U20333 ( .A(n12115), .Z(n12113) );
  AND U20334 ( .A(n12116), .B(n12117), .Z(n12082) );
  NAND U20335 ( .A(n12118), .B(n12119), .Z(n12117) );
  NANDN U20336 ( .A(n12120), .B(n12121), .Z(n12119) );
  NANDN U20337 ( .A(n12121), .B(n12120), .Z(n12116) );
  XOR U20338 ( .A(n12092), .B(n12122), .Z(n12084) );
  XNOR U20339 ( .A(n12089), .B(n12091), .Z(n12122) );
  AND U20340 ( .A(n12123), .B(n12124), .Z(n12091) );
  NANDN U20341 ( .A(n12125), .B(n12126), .Z(n12124) );
  OR U20342 ( .A(n12127), .B(n12128), .Z(n12126) );
  IV U20343 ( .A(n12129), .Z(n12128) );
  NANDN U20344 ( .A(n12129), .B(n12127), .Z(n12123) );
  AND U20345 ( .A(n12130), .B(n12131), .Z(n12089) );
  NAND U20346 ( .A(n12132), .B(n12133), .Z(n12131) );
  NANDN U20347 ( .A(n12134), .B(n12135), .Z(n12133) );
  NANDN U20348 ( .A(n12135), .B(n12134), .Z(n12130) );
  IV U20349 ( .A(n12136), .Z(n12135) );
  NAND U20350 ( .A(n12137), .B(n12138), .Z(n12092) );
  NANDN U20351 ( .A(n12139), .B(n12140), .Z(n12138) );
  NANDN U20352 ( .A(n12141), .B(n12142), .Z(n12140) );
  NANDN U20353 ( .A(n12142), .B(n12141), .Z(n12137) );
  IV U20354 ( .A(n12143), .Z(n12141) );
  XOR U20355 ( .A(n12118), .B(n12144), .Z(N64311) );
  XNOR U20356 ( .A(n12121), .B(n12120), .Z(n12144) );
  XNOR U20357 ( .A(n12132), .B(n12145), .Z(n12120) );
  XNOR U20358 ( .A(n12136), .B(n12134), .Z(n12145) );
  XOR U20359 ( .A(n12142), .B(n12146), .Z(n12134) );
  XNOR U20360 ( .A(n12139), .B(n12143), .Z(n12146) );
  AND U20361 ( .A(n12147), .B(n12148), .Z(n12143) );
  NAND U20362 ( .A(n12149), .B(n12150), .Z(n12148) );
  NAND U20363 ( .A(n12151), .B(n12152), .Z(n12147) );
  AND U20364 ( .A(n12153), .B(n12154), .Z(n12139) );
  NAND U20365 ( .A(n12155), .B(n12156), .Z(n12154) );
  NAND U20366 ( .A(n12157), .B(n12158), .Z(n12153) );
  NANDN U20367 ( .A(n12159), .B(n12160), .Z(n12142) );
  ANDN U20368 ( .B(n12161), .A(n12162), .Z(n12136) );
  XNOR U20369 ( .A(n12127), .B(n12163), .Z(n12132) );
  XNOR U20370 ( .A(n12125), .B(n12129), .Z(n12163) );
  AND U20371 ( .A(n12164), .B(n12165), .Z(n12129) );
  NAND U20372 ( .A(n12166), .B(n12167), .Z(n12165) );
  NAND U20373 ( .A(n12168), .B(n12169), .Z(n12164) );
  AND U20374 ( .A(n12170), .B(n12171), .Z(n12125) );
  NAND U20375 ( .A(n12172), .B(n12173), .Z(n12171) );
  NAND U20376 ( .A(n12174), .B(n12175), .Z(n12170) );
  AND U20377 ( .A(n12176), .B(n12177), .Z(n12127) );
  NAND U20378 ( .A(n12178), .B(n12179), .Z(n12121) );
  XNOR U20379 ( .A(n12104), .B(n12180), .Z(n12118) );
  XNOR U20380 ( .A(n12108), .B(n12106), .Z(n12180) );
  XOR U20381 ( .A(n12114), .B(n12181), .Z(n12106) );
  XNOR U20382 ( .A(n12111), .B(n12115), .Z(n12181) );
  AND U20383 ( .A(n12182), .B(n12183), .Z(n12115) );
  NAND U20384 ( .A(n12184), .B(n12185), .Z(n12183) );
  NAND U20385 ( .A(n12186), .B(n12187), .Z(n12182) );
  AND U20386 ( .A(n12188), .B(n12189), .Z(n12111) );
  NAND U20387 ( .A(n12190), .B(n12191), .Z(n12189) );
  NAND U20388 ( .A(n12192), .B(n12193), .Z(n12188) );
  NANDN U20389 ( .A(n12194), .B(n12195), .Z(n12114) );
  ANDN U20390 ( .B(n12196), .A(n12197), .Z(n12108) );
  XNOR U20391 ( .A(n12099), .B(n12198), .Z(n12104) );
  XNOR U20392 ( .A(n12097), .B(n12101), .Z(n12198) );
  AND U20393 ( .A(n12199), .B(n12200), .Z(n12101) );
  NAND U20394 ( .A(n12201), .B(n12202), .Z(n12200) );
  NAND U20395 ( .A(n12203), .B(n12204), .Z(n12199) );
  AND U20396 ( .A(n12205), .B(n12206), .Z(n12097) );
  NAND U20397 ( .A(n12207), .B(n12208), .Z(n12206) );
  NAND U20398 ( .A(n12209), .B(n12210), .Z(n12205) );
  AND U20399 ( .A(n12211), .B(n12212), .Z(n12099) );
  XOR U20400 ( .A(n12179), .B(n12178), .Z(N64310) );
  XNOR U20401 ( .A(n12196), .B(n12197), .Z(n12178) );
  XNOR U20402 ( .A(n12211), .B(n12212), .Z(n12197) );
  XOR U20403 ( .A(n12208), .B(n12207), .Z(n12212) );
  XOR U20404 ( .A(y[6876]), .B(x[6876]), .Z(n12207) );
  XOR U20405 ( .A(n12210), .B(n12209), .Z(n12208) );
  XOR U20406 ( .A(y[6878]), .B(x[6878]), .Z(n12209) );
  XOR U20407 ( .A(y[6877]), .B(x[6877]), .Z(n12210) );
  XOR U20408 ( .A(n12202), .B(n12201), .Z(n12211) );
  XOR U20409 ( .A(n12204), .B(n12203), .Z(n12201) );
  XOR U20410 ( .A(y[6875]), .B(x[6875]), .Z(n12203) );
  XOR U20411 ( .A(y[6874]), .B(x[6874]), .Z(n12204) );
  XOR U20412 ( .A(y[6873]), .B(x[6873]), .Z(n12202) );
  XNOR U20413 ( .A(n12195), .B(n12194), .Z(n12196) );
  XNOR U20414 ( .A(n12191), .B(n12190), .Z(n12194) );
  XOR U20415 ( .A(n12193), .B(n12192), .Z(n12190) );
  XOR U20416 ( .A(y[6872]), .B(x[6872]), .Z(n12192) );
  XOR U20417 ( .A(y[6871]), .B(x[6871]), .Z(n12193) );
  XOR U20418 ( .A(y[6870]), .B(x[6870]), .Z(n12191) );
  XOR U20419 ( .A(n12185), .B(n12184), .Z(n12195) );
  XOR U20420 ( .A(n12187), .B(n12186), .Z(n12184) );
  XOR U20421 ( .A(y[6869]), .B(x[6869]), .Z(n12186) );
  XOR U20422 ( .A(y[6868]), .B(x[6868]), .Z(n12187) );
  XOR U20423 ( .A(y[6867]), .B(x[6867]), .Z(n12185) );
  XNOR U20424 ( .A(n12161), .B(n12162), .Z(n12179) );
  XNOR U20425 ( .A(n12176), .B(n12177), .Z(n12162) );
  XOR U20426 ( .A(n12173), .B(n12172), .Z(n12177) );
  XOR U20427 ( .A(y[6864]), .B(x[6864]), .Z(n12172) );
  XOR U20428 ( .A(n12175), .B(n12174), .Z(n12173) );
  XOR U20429 ( .A(y[6866]), .B(x[6866]), .Z(n12174) );
  XOR U20430 ( .A(y[6865]), .B(x[6865]), .Z(n12175) );
  XOR U20431 ( .A(n12167), .B(n12166), .Z(n12176) );
  XOR U20432 ( .A(n12169), .B(n12168), .Z(n12166) );
  XOR U20433 ( .A(y[6863]), .B(x[6863]), .Z(n12168) );
  XOR U20434 ( .A(y[6862]), .B(x[6862]), .Z(n12169) );
  XOR U20435 ( .A(y[6861]), .B(x[6861]), .Z(n12167) );
  XNOR U20436 ( .A(n12160), .B(n12159), .Z(n12161) );
  XNOR U20437 ( .A(n12156), .B(n12155), .Z(n12159) );
  XOR U20438 ( .A(n12158), .B(n12157), .Z(n12155) );
  XOR U20439 ( .A(y[6860]), .B(x[6860]), .Z(n12157) );
  XOR U20440 ( .A(y[6859]), .B(x[6859]), .Z(n12158) );
  XOR U20441 ( .A(y[6858]), .B(x[6858]), .Z(n12156) );
  XOR U20442 ( .A(n12150), .B(n12149), .Z(n12160) );
  XOR U20443 ( .A(n12152), .B(n12151), .Z(n12149) );
  XOR U20444 ( .A(y[6857]), .B(x[6857]), .Z(n12151) );
  XOR U20445 ( .A(y[6856]), .B(x[6856]), .Z(n12152) );
  XOR U20446 ( .A(y[6855]), .B(x[6855]), .Z(n12150) );
  NAND U20447 ( .A(n12213), .B(n12214), .Z(N64301) );
  NAND U20448 ( .A(n12215), .B(n12216), .Z(n12214) );
  NANDN U20449 ( .A(n12217), .B(n12218), .Z(n12216) );
  NANDN U20450 ( .A(n12218), .B(n12217), .Z(n12213) );
  XOR U20451 ( .A(n12217), .B(n12219), .Z(N64300) );
  XNOR U20452 ( .A(n12215), .B(n12218), .Z(n12219) );
  NAND U20453 ( .A(n12220), .B(n12221), .Z(n12218) );
  NAND U20454 ( .A(n12222), .B(n12223), .Z(n12221) );
  NANDN U20455 ( .A(n12224), .B(n12225), .Z(n12223) );
  NANDN U20456 ( .A(n12225), .B(n12224), .Z(n12220) );
  AND U20457 ( .A(n12226), .B(n12227), .Z(n12215) );
  NAND U20458 ( .A(n12228), .B(n12229), .Z(n12227) );
  NANDN U20459 ( .A(n12230), .B(n12231), .Z(n12229) );
  NANDN U20460 ( .A(n12231), .B(n12230), .Z(n12226) );
  IV U20461 ( .A(n12232), .Z(n12231) );
  AND U20462 ( .A(n12233), .B(n12234), .Z(n12217) );
  NAND U20463 ( .A(n12235), .B(n12236), .Z(n12234) );
  NANDN U20464 ( .A(n12237), .B(n12238), .Z(n12236) );
  NANDN U20465 ( .A(n12238), .B(n12237), .Z(n12233) );
  XOR U20466 ( .A(n12230), .B(n12239), .Z(N64299) );
  XNOR U20467 ( .A(n12228), .B(n12232), .Z(n12239) );
  XOR U20468 ( .A(n12225), .B(n12240), .Z(n12232) );
  XNOR U20469 ( .A(n12222), .B(n12224), .Z(n12240) );
  AND U20470 ( .A(n12241), .B(n12242), .Z(n12224) );
  NANDN U20471 ( .A(n12243), .B(n12244), .Z(n12242) );
  OR U20472 ( .A(n12245), .B(n12246), .Z(n12244) );
  IV U20473 ( .A(n12247), .Z(n12246) );
  NANDN U20474 ( .A(n12247), .B(n12245), .Z(n12241) );
  AND U20475 ( .A(n12248), .B(n12249), .Z(n12222) );
  NAND U20476 ( .A(n12250), .B(n12251), .Z(n12249) );
  NANDN U20477 ( .A(n12252), .B(n12253), .Z(n12251) );
  NANDN U20478 ( .A(n12253), .B(n12252), .Z(n12248) );
  IV U20479 ( .A(n12254), .Z(n12253) );
  NAND U20480 ( .A(n12255), .B(n12256), .Z(n12225) );
  NANDN U20481 ( .A(n12257), .B(n12258), .Z(n12256) );
  NANDN U20482 ( .A(n12259), .B(n12260), .Z(n12258) );
  NANDN U20483 ( .A(n12260), .B(n12259), .Z(n12255) );
  IV U20484 ( .A(n12261), .Z(n12259) );
  AND U20485 ( .A(n12262), .B(n12263), .Z(n12228) );
  NAND U20486 ( .A(n12264), .B(n12265), .Z(n12263) );
  NANDN U20487 ( .A(n12266), .B(n12267), .Z(n12265) );
  NANDN U20488 ( .A(n12267), .B(n12266), .Z(n12262) );
  XOR U20489 ( .A(n12238), .B(n12268), .Z(n12230) );
  XNOR U20490 ( .A(n12235), .B(n12237), .Z(n12268) );
  AND U20491 ( .A(n12269), .B(n12270), .Z(n12237) );
  NANDN U20492 ( .A(n12271), .B(n12272), .Z(n12270) );
  OR U20493 ( .A(n12273), .B(n12274), .Z(n12272) );
  IV U20494 ( .A(n12275), .Z(n12274) );
  NANDN U20495 ( .A(n12275), .B(n12273), .Z(n12269) );
  AND U20496 ( .A(n12276), .B(n12277), .Z(n12235) );
  NAND U20497 ( .A(n12278), .B(n12279), .Z(n12277) );
  NANDN U20498 ( .A(n12280), .B(n12281), .Z(n12279) );
  NANDN U20499 ( .A(n12281), .B(n12280), .Z(n12276) );
  IV U20500 ( .A(n12282), .Z(n12281) );
  NAND U20501 ( .A(n12283), .B(n12284), .Z(n12238) );
  NANDN U20502 ( .A(n12285), .B(n12286), .Z(n12284) );
  NANDN U20503 ( .A(n12287), .B(n12288), .Z(n12286) );
  NANDN U20504 ( .A(n12288), .B(n12287), .Z(n12283) );
  IV U20505 ( .A(n12289), .Z(n12287) );
  XOR U20506 ( .A(n12264), .B(n12290), .Z(N64298) );
  XNOR U20507 ( .A(n12267), .B(n12266), .Z(n12290) );
  XNOR U20508 ( .A(n12278), .B(n12291), .Z(n12266) );
  XNOR U20509 ( .A(n12282), .B(n12280), .Z(n12291) );
  XOR U20510 ( .A(n12288), .B(n12292), .Z(n12280) );
  XNOR U20511 ( .A(n12285), .B(n12289), .Z(n12292) );
  AND U20512 ( .A(n12293), .B(n12294), .Z(n12289) );
  NAND U20513 ( .A(n12295), .B(n12296), .Z(n12294) );
  NAND U20514 ( .A(n12297), .B(n12298), .Z(n12293) );
  AND U20515 ( .A(n12299), .B(n12300), .Z(n12285) );
  NAND U20516 ( .A(n12301), .B(n12302), .Z(n12300) );
  NAND U20517 ( .A(n12303), .B(n12304), .Z(n12299) );
  NANDN U20518 ( .A(n12305), .B(n12306), .Z(n12288) );
  ANDN U20519 ( .B(n12307), .A(n12308), .Z(n12282) );
  XNOR U20520 ( .A(n12273), .B(n12309), .Z(n12278) );
  XNOR U20521 ( .A(n12271), .B(n12275), .Z(n12309) );
  AND U20522 ( .A(n12310), .B(n12311), .Z(n12275) );
  NAND U20523 ( .A(n12312), .B(n12313), .Z(n12311) );
  NAND U20524 ( .A(n12314), .B(n12315), .Z(n12310) );
  AND U20525 ( .A(n12316), .B(n12317), .Z(n12271) );
  NAND U20526 ( .A(n12318), .B(n12319), .Z(n12317) );
  NAND U20527 ( .A(n12320), .B(n12321), .Z(n12316) );
  AND U20528 ( .A(n12322), .B(n12323), .Z(n12273) );
  NAND U20529 ( .A(n12324), .B(n12325), .Z(n12267) );
  XNOR U20530 ( .A(n12250), .B(n12326), .Z(n12264) );
  XNOR U20531 ( .A(n12254), .B(n12252), .Z(n12326) );
  XOR U20532 ( .A(n12260), .B(n12327), .Z(n12252) );
  XNOR U20533 ( .A(n12257), .B(n12261), .Z(n12327) );
  AND U20534 ( .A(n12328), .B(n12329), .Z(n12261) );
  NAND U20535 ( .A(n12330), .B(n12331), .Z(n12329) );
  NAND U20536 ( .A(n12332), .B(n12333), .Z(n12328) );
  AND U20537 ( .A(n12334), .B(n12335), .Z(n12257) );
  NAND U20538 ( .A(n12336), .B(n12337), .Z(n12335) );
  NAND U20539 ( .A(n12338), .B(n12339), .Z(n12334) );
  NANDN U20540 ( .A(n12340), .B(n12341), .Z(n12260) );
  ANDN U20541 ( .B(n12342), .A(n12343), .Z(n12254) );
  XNOR U20542 ( .A(n12245), .B(n12344), .Z(n12250) );
  XNOR U20543 ( .A(n12243), .B(n12247), .Z(n12344) );
  AND U20544 ( .A(n12345), .B(n12346), .Z(n12247) );
  NAND U20545 ( .A(n12347), .B(n12348), .Z(n12346) );
  NAND U20546 ( .A(n12349), .B(n12350), .Z(n12345) );
  AND U20547 ( .A(n12351), .B(n12352), .Z(n12243) );
  NAND U20548 ( .A(n12353), .B(n12354), .Z(n12352) );
  NAND U20549 ( .A(n12355), .B(n12356), .Z(n12351) );
  AND U20550 ( .A(n12357), .B(n12358), .Z(n12245) );
  XOR U20551 ( .A(n12325), .B(n12324), .Z(N64297) );
  XNOR U20552 ( .A(n12342), .B(n12343), .Z(n12324) );
  XNOR U20553 ( .A(n12357), .B(n12358), .Z(n12343) );
  XOR U20554 ( .A(n12354), .B(n12353), .Z(n12358) );
  XOR U20555 ( .A(y[6852]), .B(x[6852]), .Z(n12353) );
  XOR U20556 ( .A(n12356), .B(n12355), .Z(n12354) );
  XOR U20557 ( .A(y[6854]), .B(x[6854]), .Z(n12355) );
  XOR U20558 ( .A(y[6853]), .B(x[6853]), .Z(n12356) );
  XOR U20559 ( .A(n12348), .B(n12347), .Z(n12357) );
  XOR U20560 ( .A(n12350), .B(n12349), .Z(n12347) );
  XOR U20561 ( .A(y[6851]), .B(x[6851]), .Z(n12349) );
  XOR U20562 ( .A(y[6850]), .B(x[6850]), .Z(n12350) );
  XOR U20563 ( .A(y[6849]), .B(x[6849]), .Z(n12348) );
  XNOR U20564 ( .A(n12341), .B(n12340), .Z(n12342) );
  XNOR U20565 ( .A(n12337), .B(n12336), .Z(n12340) );
  XOR U20566 ( .A(n12339), .B(n12338), .Z(n12336) );
  XOR U20567 ( .A(y[6848]), .B(x[6848]), .Z(n12338) );
  XOR U20568 ( .A(y[6847]), .B(x[6847]), .Z(n12339) );
  XOR U20569 ( .A(y[6846]), .B(x[6846]), .Z(n12337) );
  XOR U20570 ( .A(n12331), .B(n12330), .Z(n12341) );
  XOR U20571 ( .A(n12333), .B(n12332), .Z(n12330) );
  XOR U20572 ( .A(y[6845]), .B(x[6845]), .Z(n12332) );
  XOR U20573 ( .A(y[6844]), .B(x[6844]), .Z(n12333) );
  XOR U20574 ( .A(y[6843]), .B(x[6843]), .Z(n12331) );
  XNOR U20575 ( .A(n12307), .B(n12308), .Z(n12325) );
  XNOR U20576 ( .A(n12322), .B(n12323), .Z(n12308) );
  XOR U20577 ( .A(n12319), .B(n12318), .Z(n12323) );
  XOR U20578 ( .A(y[6840]), .B(x[6840]), .Z(n12318) );
  XOR U20579 ( .A(n12321), .B(n12320), .Z(n12319) );
  XOR U20580 ( .A(y[6842]), .B(x[6842]), .Z(n12320) );
  XOR U20581 ( .A(y[6841]), .B(x[6841]), .Z(n12321) );
  XOR U20582 ( .A(n12313), .B(n12312), .Z(n12322) );
  XOR U20583 ( .A(n12315), .B(n12314), .Z(n12312) );
  XOR U20584 ( .A(y[6839]), .B(x[6839]), .Z(n12314) );
  XOR U20585 ( .A(y[6838]), .B(x[6838]), .Z(n12315) );
  XOR U20586 ( .A(y[6837]), .B(x[6837]), .Z(n12313) );
  XNOR U20587 ( .A(n12306), .B(n12305), .Z(n12307) );
  XNOR U20588 ( .A(n12302), .B(n12301), .Z(n12305) );
  XOR U20589 ( .A(n12304), .B(n12303), .Z(n12301) );
  XOR U20590 ( .A(y[6836]), .B(x[6836]), .Z(n12303) );
  XOR U20591 ( .A(y[6835]), .B(x[6835]), .Z(n12304) );
  XOR U20592 ( .A(y[6834]), .B(x[6834]), .Z(n12302) );
  XOR U20593 ( .A(n12296), .B(n12295), .Z(n12306) );
  XOR U20594 ( .A(n12298), .B(n12297), .Z(n12295) );
  XOR U20595 ( .A(y[6833]), .B(x[6833]), .Z(n12297) );
  XOR U20596 ( .A(y[6832]), .B(x[6832]), .Z(n12298) );
  XOR U20597 ( .A(y[6831]), .B(x[6831]), .Z(n12296) );
  NAND U20598 ( .A(n12359), .B(n12360), .Z(N64288) );
  NAND U20599 ( .A(n12361), .B(n12362), .Z(n12360) );
  NANDN U20600 ( .A(n12363), .B(n12364), .Z(n12362) );
  NANDN U20601 ( .A(n12364), .B(n12363), .Z(n12359) );
  XOR U20602 ( .A(n12363), .B(n12365), .Z(N64287) );
  XNOR U20603 ( .A(n12361), .B(n12364), .Z(n12365) );
  NAND U20604 ( .A(n12366), .B(n12367), .Z(n12364) );
  NAND U20605 ( .A(n12368), .B(n12369), .Z(n12367) );
  NANDN U20606 ( .A(n12370), .B(n12371), .Z(n12369) );
  NANDN U20607 ( .A(n12371), .B(n12370), .Z(n12366) );
  AND U20608 ( .A(n12372), .B(n12373), .Z(n12361) );
  NAND U20609 ( .A(n12374), .B(n12375), .Z(n12373) );
  NANDN U20610 ( .A(n12376), .B(n12377), .Z(n12375) );
  NANDN U20611 ( .A(n12377), .B(n12376), .Z(n12372) );
  IV U20612 ( .A(n12378), .Z(n12377) );
  AND U20613 ( .A(n12379), .B(n12380), .Z(n12363) );
  NAND U20614 ( .A(n12381), .B(n12382), .Z(n12380) );
  NANDN U20615 ( .A(n12383), .B(n12384), .Z(n12382) );
  NANDN U20616 ( .A(n12384), .B(n12383), .Z(n12379) );
  XOR U20617 ( .A(n12376), .B(n12385), .Z(N64286) );
  XNOR U20618 ( .A(n12374), .B(n12378), .Z(n12385) );
  XOR U20619 ( .A(n12371), .B(n12386), .Z(n12378) );
  XNOR U20620 ( .A(n12368), .B(n12370), .Z(n12386) );
  AND U20621 ( .A(n12387), .B(n12388), .Z(n12370) );
  NANDN U20622 ( .A(n12389), .B(n12390), .Z(n12388) );
  OR U20623 ( .A(n12391), .B(n12392), .Z(n12390) );
  IV U20624 ( .A(n12393), .Z(n12392) );
  NANDN U20625 ( .A(n12393), .B(n12391), .Z(n12387) );
  AND U20626 ( .A(n12394), .B(n12395), .Z(n12368) );
  NAND U20627 ( .A(n12396), .B(n12397), .Z(n12395) );
  NANDN U20628 ( .A(n12398), .B(n12399), .Z(n12397) );
  NANDN U20629 ( .A(n12399), .B(n12398), .Z(n12394) );
  IV U20630 ( .A(n12400), .Z(n12399) );
  NAND U20631 ( .A(n12401), .B(n12402), .Z(n12371) );
  NANDN U20632 ( .A(n12403), .B(n12404), .Z(n12402) );
  NANDN U20633 ( .A(n12405), .B(n12406), .Z(n12404) );
  NANDN U20634 ( .A(n12406), .B(n12405), .Z(n12401) );
  IV U20635 ( .A(n12407), .Z(n12405) );
  AND U20636 ( .A(n12408), .B(n12409), .Z(n12374) );
  NAND U20637 ( .A(n12410), .B(n12411), .Z(n12409) );
  NANDN U20638 ( .A(n12412), .B(n12413), .Z(n12411) );
  NANDN U20639 ( .A(n12413), .B(n12412), .Z(n12408) );
  XOR U20640 ( .A(n12384), .B(n12414), .Z(n12376) );
  XNOR U20641 ( .A(n12381), .B(n12383), .Z(n12414) );
  AND U20642 ( .A(n12415), .B(n12416), .Z(n12383) );
  NANDN U20643 ( .A(n12417), .B(n12418), .Z(n12416) );
  OR U20644 ( .A(n12419), .B(n12420), .Z(n12418) );
  IV U20645 ( .A(n12421), .Z(n12420) );
  NANDN U20646 ( .A(n12421), .B(n12419), .Z(n12415) );
  AND U20647 ( .A(n12422), .B(n12423), .Z(n12381) );
  NAND U20648 ( .A(n12424), .B(n12425), .Z(n12423) );
  NANDN U20649 ( .A(n12426), .B(n12427), .Z(n12425) );
  NANDN U20650 ( .A(n12427), .B(n12426), .Z(n12422) );
  IV U20651 ( .A(n12428), .Z(n12427) );
  NAND U20652 ( .A(n12429), .B(n12430), .Z(n12384) );
  NANDN U20653 ( .A(n12431), .B(n12432), .Z(n12430) );
  NANDN U20654 ( .A(n12433), .B(n12434), .Z(n12432) );
  NANDN U20655 ( .A(n12434), .B(n12433), .Z(n12429) );
  IV U20656 ( .A(n12435), .Z(n12433) );
  XOR U20657 ( .A(n12410), .B(n12436), .Z(N64285) );
  XNOR U20658 ( .A(n12413), .B(n12412), .Z(n12436) );
  XNOR U20659 ( .A(n12424), .B(n12437), .Z(n12412) );
  XNOR U20660 ( .A(n12428), .B(n12426), .Z(n12437) );
  XOR U20661 ( .A(n12434), .B(n12438), .Z(n12426) );
  XNOR U20662 ( .A(n12431), .B(n12435), .Z(n12438) );
  AND U20663 ( .A(n12439), .B(n12440), .Z(n12435) );
  NAND U20664 ( .A(n12441), .B(n12442), .Z(n12440) );
  NAND U20665 ( .A(n12443), .B(n12444), .Z(n12439) );
  AND U20666 ( .A(n12445), .B(n12446), .Z(n12431) );
  NAND U20667 ( .A(n12447), .B(n12448), .Z(n12446) );
  NAND U20668 ( .A(n12449), .B(n12450), .Z(n12445) );
  NANDN U20669 ( .A(n12451), .B(n12452), .Z(n12434) );
  ANDN U20670 ( .B(n12453), .A(n12454), .Z(n12428) );
  XNOR U20671 ( .A(n12419), .B(n12455), .Z(n12424) );
  XNOR U20672 ( .A(n12417), .B(n12421), .Z(n12455) );
  AND U20673 ( .A(n12456), .B(n12457), .Z(n12421) );
  NAND U20674 ( .A(n12458), .B(n12459), .Z(n12457) );
  NAND U20675 ( .A(n12460), .B(n12461), .Z(n12456) );
  AND U20676 ( .A(n12462), .B(n12463), .Z(n12417) );
  NAND U20677 ( .A(n12464), .B(n12465), .Z(n12463) );
  NAND U20678 ( .A(n12466), .B(n12467), .Z(n12462) );
  AND U20679 ( .A(n12468), .B(n12469), .Z(n12419) );
  NAND U20680 ( .A(n12470), .B(n12471), .Z(n12413) );
  XNOR U20681 ( .A(n12396), .B(n12472), .Z(n12410) );
  XNOR U20682 ( .A(n12400), .B(n12398), .Z(n12472) );
  XOR U20683 ( .A(n12406), .B(n12473), .Z(n12398) );
  XNOR U20684 ( .A(n12403), .B(n12407), .Z(n12473) );
  AND U20685 ( .A(n12474), .B(n12475), .Z(n12407) );
  NAND U20686 ( .A(n12476), .B(n12477), .Z(n12475) );
  NAND U20687 ( .A(n12478), .B(n12479), .Z(n12474) );
  AND U20688 ( .A(n12480), .B(n12481), .Z(n12403) );
  NAND U20689 ( .A(n12482), .B(n12483), .Z(n12481) );
  NAND U20690 ( .A(n12484), .B(n12485), .Z(n12480) );
  NANDN U20691 ( .A(n12486), .B(n12487), .Z(n12406) );
  ANDN U20692 ( .B(n12488), .A(n12489), .Z(n12400) );
  XNOR U20693 ( .A(n12391), .B(n12490), .Z(n12396) );
  XNOR U20694 ( .A(n12389), .B(n12393), .Z(n12490) );
  AND U20695 ( .A(n12491), .B(n12492), .Z(n12393) );
  NAND U20696 ( .A(n12493), .B(n12494), .Z(n12492) );
  NAND U20697 ( .A(n12495), .B(n12496), .Z(n12491) );
  AND U20698 ( .A(n12497), .B(n12498), .Z(n12389) );
  NAND U20699 ( .A(n12499), .B(n12500), .Z(n12498) );
  NAND U20700 ( .A(n12501), .B(n12502), .Z(n12497) );
  AND U20701 ( .A(n12503), .B(n12504), .Z(n12391) );
  XOR U20702 ( .A(n12471), .B(n12470), .Z(N64284) );
  XNOR U20703 ( .A(n12488), .B(n12489), .Z(n12470) );
  XNOR U20704 ( .A(n12503), .B(n12504), .Z(n12489) );
  XOR U20705 ( .A(n12500), .B(n12499), .Z(n12504) );
  XOR U20706 ( .A(y[6828]), .B(x[6828]), .Z(n12499) );
  XOR U20707 ( .A(n12502), .B(n12501), .Z(n12500) );
  XOR U20708 ( .A(y[6830]), .B(x[6830]), .Z(n12501) );
  XOR U20709 ( .A(y[6829]), .B(x[6829]), .Z(n12502) );
  XOR U20710 ( .A(n12494), .B(n12493), .Z(n12503) );
  XOR U20711 ( .A(n12496), .B(n12495), .Z(n12493) );
  XOR U20712 ( .A(y[6827]), .B(x[6827]), .Z(n12495) );
  XOR U20713 ( .A(y[6826]), .B(x[6826]), .Z(n12496) );
  XOR U20714 ( .A(y[6825]), .B(x[6825]), .Z(n12494) );
  XNOR U20715 ( .A(n12487), .B(n12486), .Z(n12488) );
  XNOR U20716 ( .A(n12483), .B(n12482), .Z(n12486) );
  XOR U20717 ( .A(n12485), .B(n12484), .Z(n12482) );
  XOR U20718 ( .A(y[6824]), .B(x[6824]), .Z(n12484) );
  XOR U20719 ( .A(y[6823]), .B(x[6823]), .Z(n12485) );
  XOR U20720 ( .A(y[6822]), .B(x[6822]), .Z(n12483) );
  XOR U20721 ( .A(n12477), .B(n12476), .Z(n12487) );
  XOR U20722 ( .A(n12479), .B(n12478), .Z(n12476) );
  XOR U20723 ( .A(y[6821]), .B(x[6821]), .Z(n12478) );
  XOR U20724 ( .A(y[6820]), .B(x[6820]), .Z(n12479) );
  XOR U20725 ( .A(y[6819]), .B(x[6819]), .Z(n12477) );
  XNOR U20726 ( .A(n12453), .B(n12454), .Z(n12471) );
  XNOR U20727 ( .A(n12468), .B(n12469), .Z(n12454) );
  XOR U20728 ( .A(n12465), .B(n12464), .Z(n12469) );
  XOR U20729 ( .A(y[6816]), .B(x[6816]), .Z(n12464) );
  XOR U20730 ( .A(n12467), .B(n12466), .Z(n12465) );
  XOR U20731 ( .A(y[6818]), .B(x[6818]), .Z(n12466) );
  XOR U20732 ( .A(y[6817]), .B(x[6817]), .Z(n12467) );
  XOR U20733 ( .A(n12459), .B(n12458), .Z(n12468) );
  XOR U20734 ( .A(n12461), .B(n12460), .Z(n12458) );
  XOR U20735 ( .A(y[6815]), .B(x[6815]), .Z(n12460) );
  XOR U20736 ( .A(y[6814]), .B(x[6814]), .Z(n12461) );
  XOR U20737 ( .A(y[6813]), .B(x[6813]), .Z(n12459) );
  XNOR U20738 ( .A(n12452), .B(n12451), .Z(n12453) );
  XNOR U20739 ( .A(n12448), .B(n12447), .Z(n12451) );
  XOR U20740 ( .A(n12450), .B(n12449), .Z(n12447) );
  XOR U20741 ( .A(y[6812]), .B(x[6812]), .Z(n12449) );
  XOR U20742 ( .A(y[6811]), .B(x[6811]), .Z(n12450) );
  XOR U20743 ( .A(y[6810]), .B(x[6810]), .Z(n12448) );
  XOR U20744 ( .A(n12442), .B(n12441), .Z(n12452) );
  XOR U20745 ( .A(n12444), .B(n12443), .Z(n12441) );
  XOR U20746 ( .A(y[6809]), .B(x[6809]), .Z(n12443) );
  XOR U20747 ( .A(y[6808]), .B(x[6808]), .Z(n12444) );
  XOR U20748 ( .A(y[6807]), .B(x[6807]), .Z(n12442) );
  NAND U20749 ( .A(n12505), .B(n12506), .Z(N64275) );
  NAND U20750 ( .A(n12507), .B(n12508), .Z(n12506) );
  NANDN U20751 ( .A(n12509), .B(n12510), .Z(n12508) );
  NANDN U20752 ( .A(n12510), .B(n12509), .Z(n12505) );
  XOR U20753 ( .A(n12509), .B(n12511), .Z(N64274) );
  XNOR U20754 ( .A(n12507), .B(n12510), .Z(n12511) );
  NAND U20755 ( .A(n12512), .B(n12513), .Z(n12510) );
  NAND U20756 ( .A(n12514), .B(n12515), .Z(n12513) );
  NANDN U20757 ( .A(n12516), .B(n12517), .Z(n12515) );
  NANDN U20758 ( .A(n12517), .B(n12516), .Z(n12512) );
  AND U20759 ( .A(n12518), .B(n12519), .Z(n12507) );
  NAND U20760 ( .A(n12520), .B(n12521), .Z(n12519) );
  NANDN U20761 ( .A(n12522), .B(n12523), .Z(n12521) );
  NANDN U20762 ( .A(n12523), .B(n12522), .Z(n12518) );
  IV U20763 ( .A(n12524), .Z(n12523) );
  AND U20764 ( .A(n12525), .B(n12526), .Z(n12509) );
  NAND U20765 ( .A(n12527), .B(n12528), .Z(n12526) );
  NANDN U20766 ( .A(n12529), .B(n12530), .Z(n12528) );
  NANDN U20767 ( .A(n12530), .B(n12529), .Z(n12525) );
  XOR U20768 ( .A(n12522), .B(n12531), .Z(N64273) );
  XNOR U20769 ( .A(n12520), .B(n12524), .Z(n12531) );
  XOR U20770 ( .A(n12517), .B(n12532), .Z(n12524) );
  XNOR U20771 ( .A(n12514), .B(n12516), .Z(n12532) );
  AND U20772 ( .A(n12533), .B(n12534), .Z(n12516) );
  NANDN U20773 ( .A(n12535), .B(n12536), .Z(n12534) );
  OR U20774 ( .A(n12537), .B(n12538), .Z(n12536) );
  IV U20775 ( .A(n12539), .Z(n12538) );
  NANDN U20776 ( .A(n12539), .B(n12537), .Z(n12533) );
  AND U20777 ( .A(n12540), .B(n12541), .Z(n12514) );
  NAND U20778 ( .A(n12542), .B(n12543), .Z(n12541) );
  NANDN U20779 ( .A(n12544), .B(n12545), .Z(n12543) );
  NANDN U20780 ( .A(n12545), .B(n12544), .Z(n12540) );
  IV U20781 ( .A(n12546), .Z(n12545) );
  NAND U20782 ( .A(n12547), .B(n12548), .Z(n12517) );
  NANDN U20783 ( .A(n12549), .B(n12550), .Z(n12548) );
  NANDN U20784 ( .A(n12551), .B(n12552), .Z(n12550) );
  NANDN U20785 ( .A(n12552), .B(n12551), .Z(n12547) );
  IV U20786 ( .A(n12553), .Z(n12551) );
  AND U20787 ( .A(n12554), .B(n12555), .Z(n12520) );
  NAND U20788 ( .A(n12556), .B(n12557), .Z(n12555) );
  NANDN U20789 ( .A(n12558), .B(n12559), .Z(n12557) );
  NANDN U20790 ( .A(n12559), .B(n12558), .Z(n12554) );
  XOR U20791 ( .A(n12530), .B(n12560), .Z(n12522) );
  XNOR U20792 ( .A(n12527), .B(n12529), .Z(n12560) );
  AND U20793 ( .A(n12561), .B(n12562), .Z(n12529) );
  NANDN U20794 ( .A(n12563), .B(n12564), .Z(n12562) );
  OR U20795 ( .A(n12565), .B(n12566), .Z(n12564) );
  IV U20796 ( .A(n12567), .Z(n12566) );
  NANDN U20797 ( .A(n12567), .B(n12565), .Z(n12561) );
  AND U20798 ( .A(n12568), .B(n12569), .Z(n12527) );
  NAND U20799 ( .A(n12570), .B(n12571), .Z(n12569) );
  NANDN U20800 ( .A(n12572), .B(n12573), .Z(n12571) );
  NANDN U20801 ( .A(n12573), .B(n12572), .Z(n12568) );
  IV U20802 ( .A(n12574), .Z(n12573) );
  NAND U20803 ( .A(n12575), .B(n12576), .Z(n12530) );
  NANDN U20804 ( .A(n12577), .B(n12578), .Z(n12576) );
  NANDN U20805 ( .A(n12579), .B(n12580), .Z(n12578) );
  NANDN U20806 ( .A(n12580), .B(n12579), .Z(n12575) );
  IV U20807 ( .A(n12581), .Z(n12579) );
  XOR U20808 ( .A(n12556), .B(n12582), .Z(N64272) );
  XNOR U20809 ( .A(n12559), .B(n12558), .Z(n12582) );
  XNOR U20810 ( .A(n12570), .B(n12583), .Z(n12558) );
  XNOR U20811 ( .A(n12574), .B(n12572), .Z(n12583) );
  XOR U20812 ( .A(n12580), .B(n12584), .Z(n12572) );
  XNOR U20813 ( .A(n12577), .B(n12581), .Z(n12584) );
  AND U20814 ( .A(n12585), .B(n12586), .Z(n12581) );
  NAND U20815 ( .A(n12587), .B(n12588), .Z(n12586) );
  NAND U20816 ( .A(n12589), .B(n12590), .Z(n12585) );
  AND U20817 ( .A(n12591), .B(n12592), .Z(n12577) );
  NAND U20818 ( .A(n12593), .B(n12594), .Z(n12592) );
  NAND U20819 ( .A(n12595), .B(n12596), .Z(n12591) );
  NANDN U20820 ( .A(n12597), .B(n12598), .Z(n12580) );
  ANDN U20821 ( .B(n12599), .A(n12600), .Z(n12574) );
  XNOR U20822 ( .A(n12565), .B(n12601), .Z(n12570) );
  XNOR U20823 ( .A(n12563), .B(n12567), .Z(n12601) );
  AND U20824 ( .A(n12602), .B(n12603), .Z(n12567) );
  NAND U20825 ( .A(n12604), .B(n12605), .Z(n12603) );
  NAND U20826 ( .A(n12606), .B(n12607), .Z(n12602) );
  AND U20827 ( .A(n12608), .B(n12609), .Z(n12563) );
  NAND U20828 ( .A(n12610), .B(n12611), .Z(n12609) );
  NAND U20829 ( .A(n12612), .B(n12613), .Z(n12608) );
  AND U20830 ( .A(n12614), .B(n12615), .Z(n12565) );
  NAND U20831 ( .A(n12616), .B(n12617), .Z(n12559) );
  XNOR U20832 ( .A(n12542), .B(n12618), .Z(n12556) );
  XNOR U20833 ( .A(n12546), .B(n12544), .Z(n12618) );
  XOR U20834 ( .A(n12552), .B(n12619), .Z(n12544) );
  XNOR U20835 ( .A(n12549), .B(n12553), .Z(n12619) );
  AND U20836 ( .A(n12620), .B(n12621), .Z(n12553) );
  NAND U20837 ( .A(n12622), .B(n12623), .Z(n12621) );
  NAND U20838 ( .A(n12624), .B(n12625), .Z(n12620) );
  AND U20839 ( .A(n12626), .B(n12627), .Z(n12549) );
  NAND U20840 ( .A(n12628), .B(n12629), .Z(n12627) );
  NAND U20841 ( .A(n12630), .B(n12631), .Z(n12626) );
  NANDN U20842 ( .A(n12632), .B(n12633), .Z(n12552) );
  ANDN U20843 ( .B(n12634), .A(n12635), .Z(n12546) );
  XNOR U20844 ( .A(n12537), .B(n12636), .Z(n12542) );
  XNOR U20845 ( .A(n12535), .B(n12539), .Z(n12636) );
  AND U20846 ( .A(n12637), .B(n12638), .Z(n12539) );
  NAND U20847 ( .A(n12639), .B(n12640), .Z(n12638) );
  NAND U20848 ( .A(n12641), .B(n12642), .Z(n12637) );
  AND U20849 ( .A(n12643), .B(n12644), .Z(n12535) );
  NAND U20850 ( .A(n12645), .B(n12646), .Z(n12644) );
  NAND U20851 ( .A(n12647), .B(n12648), .Z(n12643) );
  AND U20852 ( .A(n12649), .B(n12650), .Z(n12537) );
  XOR U20853 ( .A(n12617), .B(n12616), .Z(N64271) );
  XNOR U20854 ( .A(n12634), .B(n12635), .Z(n12616) );
  XNOR U20855 ( .A(n12649), .B(n12650), .Z(n12635) );
  XOR U20856 ( .A(n12646), .B(n12645), .Z(n12650) );
  XOR U20857 ( .A(y[6804]), .B(x[6804]), .Z(n12645) );
  XOR U20858 ( .A(n12648), .B(n12647), .Z(n12646) );
  XOR U20859 ( .A(y[6806]), .B(x[6806]), .Z(n12647) );
  XOR U20860 ( .A(y[6805]), .B(x[6805]), .Z(n12648) );
  XOR U20861 ( .A(n12640), .B(n12639), .Z(n12649) );
  XOR U20862 ( .A(n12642), .B(n12641), .Z(n12639) );
  XOR U20863 ( .A(y[6803]), .B(x[6803]), .Z(n12641) );
  XOR U20864 ( .A(y[6802]), .B(x[6802]), .Z(n12642) );
  XOR U20865 ( .A(y[6801]), .B(x[6801]), .Z(n12640) );
  XNOR U20866 ( .A(n12633), .B(n12632), .Z(n12634) );
  XNOR U20867 ( .A(n12629), .B(n12628), .Z(n12632) );
  XOR U20868 ( .A(n12631), .B(n12630), .Z(n12628) );
  XOR U20869 ( .A(y[6800]), .B(x[6800]), .Z(n12630) );
  XOR U20870 ( .A(y[6799]), .B(x[6799]), .Z(n12631) );
  XOR U20871 ( .A(y[6798]), .B(x[6798]), .Z(n12629) );
  XOR U20872 ( .A(n12623), .B(n12622), .Z(n12633) );
  XOR U20873 ( .A(n12625), .B(n12624), .Z(n12622) );
  XOR U20874 ( .A(y[6797]), .B(x[6797]), .Z(n12624) );
  XOR U20875 ( .A(y[6796]), .B(x[6796]), .Z(n12625) );
  XOR U20876 ( .A(y[6795]), .B(x[6795]), .Z(n12623) );
  XNOR U20877 ( .A(n12599), .B(n12600), .Z(n12617) );
  XNOR U20878 ( .A(n12614), .B(n12615), .Z(n12600) );
  XOR U20879 ( .A(n12611), .B(n12610), .Z(n12615) );
  XOR U20880 ( .A(y[6792]), .B(x[6792]), .Z(n12610) );
  XOR U20881 ( .A(n12613), .B(n12612), .Z(n12611) );
  XOR U20882 ( .A(y[6794]), .B(x[6794]), .Z(n12612) );
  XOR U20883 ( .A(y[6793]), .B(x[6793]), .Z(n12613) );
  XOR U20884 ( .A(n12605), .B(n12604), .Z(n12614) );
  XOR U20885 ( .A(n12607), .B(n12606), .Z(n12604) );
  XOR U20886 ( .A(y[6791]), .B(x[6791]), .Z(n12606) );
  XOR U20887 ( .A(y[6790]), .B(x[6790]), .Z(n12607) );
  XOR U20888 ( .A(y[6789]), .B(x[6789]), .Z(n12605) );
  XNOR U20889 ( .A(n12598), .B(n12597), .Z(n12599) );
  XNOR U20890 ( .A(n12594), .B(n12593), .Z(n12597) );
  XOR U20891 ( .A(n12596), .B(n12595), .Z(n12593) );
  XOR U20892 ( .A(y[6788]), .B(x[6788]), .Z(n12595) );
  XOR U20893 ( .A(y[6787]), .B(x[6787]), .Z(n12596) );
  XOR U20894 ( .A(y[6786]), .B(x[6786]), .Z(n12594) );
  XOR U20895 ( .A(n12588), .B(n12587), .Z(n12598) );
  XOR U20896 ( .A(n12590), .B(n12589), .Z(n12587) );
  XOR U20897 ( .A(y[6785]), .B(x[6785]), .Z(n12589) );
  XOR U20898 ( .A(y[6784]), .B(x[6784]), .Z(n12590) );
  XOR U20899 ( .A(y[6783]), .B(x[6783]), .Z(n12588) );
  NAND U20900 ( .A(n12651), .B(n12652), .Z(N64262) );
  NAND U20901 ( .A(n12653), .B(n12654), .Z(n12652) );
  NANDN U20902 ( .A(n12655), .B(n12656), .Z(n12654) );
  NANDN U20903 ( .A(n12656), .B(n12655), .Z(n12651) );
  XOR U20904 ( .A(n12655), .B(n12657), .Z(N64261) );
  XNOR U20905 ( .A(n12653), .B(n12656), .Z(n12657) );
  NAND U20906 ( .A(n12658), .B(n12659), .Z(n12656) );
  NAND U20907 ( .A(n12660), .B(n12661), .Z(n12659) );
  NANDN U20908 ( .A(n12662), .B(n12663), .Z(n12661) );
  NANDN U20909 ( .A(n12663), .B(n12662), .Z(n12658) );
  AND U20910 ( .A(n12664), .B(n12665), .Z(n12653) );
  NAND U20911 ( .A(n12666), .B(n12667), .Z(n12665) );
  NANDN U20912 ( .A(n12668), .B(n12669), .Z(n12667) );
  NANDN U20913 ( .A(n12669), .B(n12668), .Z(n12664) );
  IV U20914 ( .A(n12670), .Z(n12669) );
  AND U20915 ( .A(n12671), .B(n12672), .Z(n12655) );
  NAND U20916 ( .A(n12673), .B(n12674), .Z(n12672) );
  NANDN U20917 ( .A(n12675), .B(n12676), .Z(n12674) );
  NANDN U20918 ( .A(n12676), .B(n12675), .Z(n12671) );
  XOR U20919 ( .A(n12668), .B(n12677), .Z(N64260) );
  XNOR U20920 ( .A(n12666), .B(n12670), .Z(n12677) );
  XOR U20921 ( .A(n12663), .B(n12678), .Z(n12670) );
  XNOR U20922 ( .A(n12660), .B(n12662), .Z(n12678) );
  AND U20923 ( .A(n12679), .B(n12680), .Z(n12662) );
  NANDN U20924 ( .A(n12681), .B(n12682), .Z(n12680) );
  OR U20925 ( .A(n12683), .B(n12684), .Z(n12682) );
  IV U20926 ( .A(n12685), .Z(n12684) );
  NANDN U20927 ( .A(n12685), .B(n12683), .Z(n12679) );
  AND U20928 ( .A(n12686), .B(n12687), .Z(n12660) );
  NAND U20929 ( .A(n12688), .B(n12689), .Z(n12687) );
  NANDN U20930 ( .A(n12690), .B(n12691), .Z(n12689) );
  NANDN U20931 ( .A(n12691), .B(n12690), .Z(n12686) );
  IV U20932 ( .A(n12692), .Z(n12691) );
  NAND U20933 ( .A(n12693), .B(n12694), .Z(n12663) );
  NANDN U20934 ( .A(n12695), .B(n12696), .Z(n12694) );
  NANDN U20935 ( .A(n12697), .B(n12698), .Z(n12696) );
  NANDN U20936 ( .A(n12698), .B(n12697), .Z(n12693) );
  IV U20937 ( .A(n12699), .Z(n12697) );
  AND U20938 ( .A(n12700), .B(n12701), .Z(n12666) );
  NAND U20939 ( .A(n12702), .B(n12703), .Z(n12701) );
  NANDN U20940 ( .A(n12704), .B(n12705), .Z(n12703) );
  NANDN U20941 ( .A(n12705), .B(n12704), .Z(n12700) );
  XOR U20942 ( .A(n12676), .B(n12706), .Z(n12668) );
  XNOR U20943 ( .A(n12673), .B(n12675), .Z(n12706) );
  AND U20944 ( .A(n12707), .B(n12708), .Z(n12675) );
  NANDN U20945 ( .A(n12709), .B(n12710), .Z(n12708) );
  OR U20946 ( .A(n12711), .B(n12712), .Z(n12710) );
  IV U20947 ( .A(n12713), .Z(n12712) );
  NANDN U20948 ( .A(n12713), .B(n12711), .Z(n12707) );
  AND U20949 ( .A(n12714), .B(n12715), .Z(n12673) );
  NAND U20950 ( .A(n12716), .B(n12717), .Z(n12715) );
  NANDN U20951 ( .A(n12718), .B(n12719), .Z(n12717) );
  NANDN U20952 ( .A(n12719), .B(n12718), .Z(n12714) );
  IV U20953 ( .A(n12720), .Z(n12719) );
  NAND U20954 ( .A(n12721), .B(n12722), .Z(n12676) );
  NANDN U20955 ( .A(n12723), .B(n12724), .Z(n12722) );
  NANDN U20956 ( .A(n12725), .B(n12726), .Z(n12724) );
  NANDN U20957 ( .A(n12726), .B(n12725), .Z(n12721) );
  IV U20958 ( .A(n12727), .Z(n12725) );
  XOR U20959 ( .A(n12702), .B(n12728), .Z(N64259) );
  XNOR U20960 ( .A(n12705), .B(n12704), .Z(n12728) );
  XNOR U20961 ( .A(n12716), .B(n12729), .Z(n12704) );
  XNOR U20962 ( .A(n12720), .B(n12718), .Z(n12729) );
  XOR U20963 ( .A(n12726), .B(n12730), .Z(n12718) );
  XNOR U20964 ( .A(n12723), .B(n12727), .Z(n12730) );
  AND U20965 ( .A(n12731), .B(n12732), .Z(n12727) );
  NAND U20966 ( .A(n12733), .B(n12734), .Z(n12732) );
  NAND U20967 ( .A(n12735), .B(n12736), .Z(n12731) );
  AND U20968 ( .A(n12737), .B(n12738), .Z(n12723) );
  NAND U20969 ( .A(n12739), .B(n12740), .Z(n12738) );
  NAND U20970 ( .A(n12741), .B(n12742), .Z(n12737) );
  NANDN U20971 ( .A(n12743), .B(n12744), .Z(n12726) );
  ANDN U20972 ( .B(n12745), .A(n12746), .Z(n12720) );
  XNOR U20973 ( .A(n12711), .B(n12747), .Z(n12716) );
  XNOR U20974 ( .A(n12709), .B(n12713), .Z(n12747) );
  AND U20975 ( .A(n12748), .B(n12749), .Z(n12713) );
  NAND U20976 ( .A(n12750), .B(n12751), .Z(n12749) );
  NAND U20977 ( .A(n12752), .B(n12753), .Z(n12748) );
  AND U20978 ( .A(n12754), .B(n12755), .Z(n12709) );
  NAND U20979 ( .A(n12756), .B(n12757), .Z(n12755) );
  NAND U20980 ( .A(n12758), .B(n12759), .Z(n12754) );
  AND U20981 ( .A(n12760), .B(n12761), .Z(n12711) );
  NAND U20982 ( .A(n12762), .B(n12763), .Z(n12705) );
  XNOR U20983 ( .A(n12688), .B(n12764), .Z(n12702) );
  XNOR U20984 ( .A(n12692), .B(n12690), .Z(n12764) );
  XOR U20985 ( .A(n12698), .B(n12765), .Z(n12690) );
  XNOR U20986 ( .A(n12695), .B(n12699), .Z(n12765) );
  AND U20987 ( .A(n12766), .B(n12767), .Z(n12699) );
  NAND U20988 ( .A(n12768), .B(n12769), .Z(n12767) );
  NAND U20989 ( .A(n12770), .B(n12771), .Z(n12766) );
  AND U20990 ( .A(n12772), .B(n12773), .Z(n12695) );
  NAND U20991 ( .A(n12774), .B(n12775), .Z(n12773) );
  NAND U20992 ( .A(n12776), .B(n12777), .Z(n12772) );
  NANDN U20993 ( .A(n12778), .B(n12779), .Z(n12698) );
  ANDN U20994 ( .B(n12780), .A(n12781), .Z(n12692) );
  XNOR U20995 ( .A(n12683), .B(n12782), .Z(n12688) );
  XNOR U20996 ( .A(n12681), .B(n12685), .Z(n12782) );
  AND U20997 ( .A(n12783), .B(n12784), .Z(n12685) );
  NAND U20998 ( .A(n12785), .B(n12786), .Z(n12784) );
  NAND U20999 ( .A(n12787), .B(n12788), .Z(n12783) );
  AND U21000 ( .A(n12789), .B(n12790), .Z(n12681) );
  NAND U21001 ( .A(n12791), .B(n12792), .Z(n12790) );
  NAND U21002 ( .A(n12793), .B(n12794), .Z(n12789) );
  AND U21003 ( .A(n12795), .B(n12796), .Z(n12683) );
  XOR U21004 ( .A(n12763), .B(n12762), .Z(N64258) );
  XNOR U21005 ( .A(n12780), .B(n12781), .Z(n12762) );
  XNOR U21006 ( .A(n12795), .B(n12796), .Z(n12781) );
  XOR U21007 ( .A(n12792), .B(n12791), .Z(n12796) );
  XOR U21008 ( .A(y[6780]), .B(x[6780]), .Z(n12791) );
  XOR U21009 ( .A(n12794), .B(n12793), .Z(n12792) );
  XOR U21010 ( .A(y[6782]), .B(x[6782]), .Z(n12793) );
  XOR U21011 ( .A(y[6781]), .B(x[6781]), .Z(n12794) );
  XOR U21012 ( .A(n12786), .B(n12785), .Z(n12795) );
  XOR U21013 ( .A(n12788), .B(n12787), .Z(n12785) );
  XOR U21014 ( .A(y[6779]), .B(x[6779]), .Z(n12787) );
  XOR U21015 ( .A(y[6778]), .B(x[6778]), .Z(n12788) );
  XOR U21016 ( .A(y[6777]), .B(x[6777]), .Z(n12786) );
  XNOR U21017 ( .A(n12779), .B(n12778), .Z(n12780) );
  XNOR U21018 ( .A(n12775), .B(n12774), .Z(n12778) );
  XOR U21019 ( .A(n12777), .B(n12776), .Z(n12774) );
  XOR U21020 ( .A(y[6776]), .B(x[6776]), .Z(n12776) );
  XOR U21021 ( .A(y[6775]), .B(x[6775]), .Z(n12777) );
  XOR U21022 ( .A(y[6774]), .B(x[6774]), .Z(n12775) );
  XOR U21023 ( .A(n12769), .B(n12768), .Z(n12779) );
  XOR U21024 ( .A(n12771), .B(n12770), .Z(n12768) );
  XOR U21025 ( .A(y[6773]), .B(x[6773]), .Z(n12770) );
  XOR U21026 ( .A(y[6772]), .B(x[6772]), .Z(n12771) );
  XOR U21027 ( .A(y[6771]), .B(x[6771]), .Z(n12769) );
  XNOR U21028 ( .A(n12745), .B(n12746), .Z(n12763) );
  XNOR U21029 ( .A(n12760), .B(n12761), .Z(n12746) );
  XOR U21030 ( .A(n12757), .B(n12756), .Z(n12761) );
  XOR U21031 ( .A(y[6768]), .B(x[6768]), .Z(n12756) );
  XOR U21032 ( .A(n12759), .B(n12758), .Z(n12757) );
  XOR U21033 ( .A(y[6770]), .B(x[6770]), .Z(n12758) );
  XOR U21034 ( .A(y[6769]), .B(x[6769]), .Z(n12759) );
  XOR U21035 ( .A(n12751), .B(n12750), .Z(n12760) );
  XOR U21036 ( .A(n12753), .B(n12752), .Z(n12750) );
  XOR U21037 ( .A(y[6767]), .B(x[6767]), .Z(n12752) );
  XOR U21038 ( .A(y[6766]), .B(x[6766]), .Z(n12753) );
  XOR U21039 ( .A(y[6765]), .B(x[6765]), .Z(n12751) );
  XNOR U21040 ( .A(n12744), .B(n12743), .Z(n12745) );
  XNOR U21041 ( .A(n12740), .B(n12739), .Z(n12743) );
  XOR U21042 ( .A(n12742), .B(n12741), .Z(n12739) );
  XOR U21043 ( .A(y[6764]), .B(x[6764]), .Z(n12741) );
  XOR U21044 ( .A(y[6763]), .B(x[6763]), .Z(n12742) );
  XOR U21045 ( .A(y[6762]), .B(x[6762]), .Z(n12740) );
  XOR U21046 ( .A(n12734), .B(n12733), .Z(n12744) );
  XOR U21047 ( .A(n12736), .B(n12735), .Z(n12733) );
  XOR U21048 ( .A(y[6761]), .B(x[6761]), .Z(n12735) );
  XOR U21049 ( .A(y[6760]), .B(x[6760]), .Z(n12736) );
  XOR U21050 ( .A(y[6759]), .B(x[6759]), .Z(n12734) );
  NAND U21051 ( .A(n12797), .B(n12798), .Z(N64249) );
  NAND U21052 ( .A(n12799), .B(n12800), .Z(n12798) );
  NANDN U21053 ( .A(n12801), .B(n12802), .Z(n12800) );
  NANDN U21054 ( .A(n12802), .B(n12801), .Z(n12797) );
  XOR U21055 ( .A(n12801), .B(n12803), .Z(N64248) );
  XNOR U21056 ( .A(n12799), .B(n12802), .Z(n12803) );
  NAND U21057 ( .A(n12804), .B(n12805), .Z(n12802) );
  NAND U21058 ( .A(n12806), .B(n12807), .Z(n12805) );
  NANDN U21059 ( .A(n12808), .B(n12809), .Z(n12807) );
  NANDN U21060 ( .A(n12809), .B(n12808), .Z(n12804) );
  AND U21061 ( .A(n12810), .B(n12811), .Z(n12799) );
  NAND U21062 ( .A(n12812), .B(n12813), .Z(n12811) );
  NANDN U21063 ( .A(n12814), .B(n12815), .Z(n12813) );
  NANDN U21064 ( .A(n12815), .B(n12814), .Z(n12810) );
  IV U21065 ( .A(n12816), .Z(n12815) );
  AND U21066 ( .A(n12817), .B(n12818), .Z(n12801) );
  NAND U21067 ( .A(n12819), .B(n12820), .Z(n12818) );
  NANDN U21068 ( .A(n12821), .B(n12822), .Z(n12820) );
  NANDN U21069 ( .A(n12822), .B(n12821), .Z(n12817) );
  XOR U21070 ( .A(n12814), .B(n12823), .Z(N64247) );
  XNOR U21071 ( .A(n12812), .B(n12816), .Z(n12823) );
  XOR U21072 ( .A(n12809), .B(n12824), .Z(n12816) );
  XNOR U21073 ( .A(n12806), .B(n12808), .Z(n12824) );
  AND U21074 ( .A(n12825), .B(n12826), .Z(n12808) );
  NANDN U21075 ( .A(n12827), .B(n12828), .Z(n12826) );
  OR U21076 ( .A(n12829), .B(n12830), .Z(n12828) );
  IV U21077 ( .A(n12831), .Z(n12830) );
  NANDN U21078 ( .A(n12831), .B(n12829), .Z(n12825) );
  AND U21079 ( .A(n12832), .B(n12833), .Z(n12806) );
  NAND U21080 ( .A(n12834), .B(n12835), .Z(n12833) );
  NANDN U21081 ( .A(n12836), .B(n12837), .Z(n12835) );
  NANDN U21082 ( .A(n12837), .B(n12836), .Z(n12832) );
  IV U21083 ( .A(n12838), .Z(n12837) );
  NAND U21084 ( .A(n12839), .B(n12840), .Z(n12809) );
  NANDN U21085 ( .A(n12841), .B(n12842), .Z(n12840) );
  NANDN U21086 ( .A(n12843), .B(n12844), .Z(n12842) );
  NANDN U21087 ( .A(n12844), .B(n12843), .Z(n12839) );
  IV U21088 ( .A(n12845), .Z(n12843) );
  AND U21089 ( .A(n12846), .B(n12847), .Z(n12812) );
  NAND U21090 ( .A(n12848), .B(n12849), .Z(n12847) );
  NANDN U21091 ( .A(n12850), .B(n12851), .Z(n12849) );
  NANDN U21092 ( .A(n12851), .B(n12850), .Z(n12846) );
  XOR U21093 ( .A(n12822), .B(n12852), .Z(n12814) );
  XNOR U21094 ( .A(n12819), .B(n12821), .Z(n12852) );
  AND U21095 ( .A(n12853), .B(n12854), .Z(n12821) );
  NANDN U21096 ( .A(n12855), .B(n12856), .Z(n12854) );
  OR U21097 ( .A(n12857), .B(n12858), .Z(n12856) );
  IV U21098 ( .A(n12859), .Z(n12858) );
  NANDN U21099 ( .A(n12859), .B(n12857), .Z(n12853) );
  AND U21100 ( .A(n12860), .B(n12861), .Z(n12819) );
  NAND U21101 ( .A(n12862), .B(n12863), .Z(n12861) );
  NANDN U21102 ( .A(n12864), .B(n12865), .Z(n12863) );
  NANDN U21103 ( .A(n12865), .B(n12864), .Z(n12860) );
  IV U21104 ( .A(n12866), .Z(n12865) );
  NAND U21105 ( .A(n12867), .B(n12868), .Z(n12822) );
  NANDN U21106 ( .A(n12869), .B(n12870), .Z(n12868) );
  NANDN U21107 ( .A(n12871), .B(n12872), .Z(n12870) );
  NANDN U21108 ( .A(n12872), .B(n12871), .Z(n12867) );
  IV U21109 ( .A(n12873), .Z(n12871) );
  XOR U21110 ( .A(n12848), .B(n12874), .Z(N64246) );
  XNOR U21111 ( .A(n12851), .B(n12850), .Z(n12874) );
  XNOR U21112 ( .A(n12862), .B(n12875), .Z(n12850) );
  XNOR U21113 ( .A(n12866), .B(n12864), .Z(n12875) );
  XOR U21114 ( .A(n12872), .B(n12876), .Z(n12864) );
  XNOR U21115 ( .A(n12869), .B(n12873), .Z(n12876) );
  AND U21116 ( .A(n12877), .B(n12878), .Z(n12873) );
  NAND U21117 ( .A(n12879), .B(n12880), .Z(n12878) );
  NAND U21118 ( .A(n12881), .B(n12882), .Z(n12877) );
  AND U21119 ( .A(n12883), .B(n12884), .Z(n12869) );
  NAND U21120 ( .A(n12885), .B(n12886), .Z(n12884) );
  NAND U21121 ( .A(n12887), .B(n12888), .Z(n12883) );
  NANDN U21122 ( .A(n12889), .B(n12890), .Z(n12872) );
  ANDN U21123 ( .B(n12891), .A(n12892), .Z(n12866) );
  XNOR U21124 ( .A(n12857), .B(n12893), .Z(n12862) );
  XNOR U21125 ( .A(n12855), .B(n12859), .Z(n12893) );
  AND U21126 ( .A(n12894), .B(n12895), .Z(n12859) );
  NAND U21127 ( .A(n12896), .B(n12897), .Z(n12895) );
  NAND U21128 ( .A(n12898), .B(n12899), .Z(n12894) );
  AND U21129 ( .A(n12900), .B(n12901), .Z(n12855) );
  NAND U21130 ( .A(n12902), .B(n12903), .Z(n12901) );
  NAND U21131 ( .A(n12904), .B(n12905), .Z(n12900) );
  AND U21132 ( .A(n12906), .B(n12907), .Z(n12857) );
  NAND U21133 ( .A(n12908), .B(n12909), .Z(n12851) );
  XNOR U21134 ( .A(n12834), .B(n12910), .Z(n12848) );
  XNOR U21135 ( .A(n12838), .B(n12836), .Z(n12910) );
  XOR U21136 ( .A(n12844), .B(n12911), .Z(n12836) );
  XNOR U21137 ( .A(n12841), .B(n12845), .Z(n12911) );
  AND U21138 ( .A(n12912), .B(n12913), .Z(n12845) );
  NAND U21139 ( .A(n12914), .B(n12915), .Z(n12913) );
  NAND U21140 ( .A(n12916), .B(n12917), .Z(n12912) );
  AND U21141 ( .A(n12918), .B(n12919), .Z(n12841) );
  NAND U21142 ( .A(n12920), .B(n12921), .Z(n12919) );
  NAND U21143 ( .A(n12922), .B(n12923), .Z(n12918) );
  NANDN U21144 ( .A(n12924), .B(n12925), .Z(n12844) );
  ANDN U21145 ( .B(n12926), .A(n12927), .Z(n12838) );
  XNOR U21146 ( .A(n12829), .B(n12928), .Z(n12834) );
  XNOR U21147 ( .A(n12827), .B(n12831), .Z(n12928) );
  AND U21148 ( .A(n12929), .B(n12930), .Z(n12831) );
  NAND U21149 ( .A(n12931), .B(n12932), .Z(n12930) );
  NAND U21150 ( .A(n12933), .B(n12934), .Z(n12929) );
  AND U21151 ( .A(n12935), .B(n12936), .Z(n12827) );
  NAND U21152 ( .A(n12937), .B(n12938), .Z(n12936) );
  NAND U21153 ( .A(n12939), .B(n12940), .Z(n12935) );
  AND U21154 ( .A(n12941), .B(n12942), .Z(n12829) );
  XOR U21155 ( .A(n12909), .B(n12908), .Z(N64245) );
  XNOR U21156 ( .A(n12926), .B(n12927), .Z(n12908) );
  XNOR U21157 ( .A(n12941), .B(n12942), .Z(n12927) );
  XOR U21158 ( .A(n12938), .B(n12937), .Z(n12942) );
  XOR U21159 ( .A(y[6756]), .B(x[6756]), .Z(n12937) );
  XOR U21160 ( .A(n12940), .B(n12939), .Z(n12938) );
  XOR U21161 ( .A(y[6758]), .B(x[6758]), .Z(n12939) );
  XOR U21162 ( .A(y[6757]), .B(x[6757]), .Z(n12940) );
  XOR U21163 ( .A(n12932), .B(n12931), .Z(n12941) );
  XOR U21164 ( .A(n12934), .B(n12933), .Z(n12931) );
  XOR U21165 ( .A(y[6755]), .B(x[6755]), .Z(n12933) );
  XOR U21166 ( .A(y[6754]), .B(x[6754]), .Z(n12934) );
  XOR U21167 ( .A(y[6753]), .B(x[6753]), .Z(n12932) );
  XNOR U21168 ( .A(n12925), .B(n12924), .Z(n12926) );
  XNOR U21169 ( .A(n12921), .B(n12920), .Z(n12924) );
  XOR U21170 ( .A(n12923), .B(n12922), .Z(n12920) );
  XOR U21171 ( .A(y[6752]), .B(x[6752]), .Z(n12922) );
  XOR U21172 ( .A(y[6751]), .B(x[6751]), .Z(n12923) );
  XOR U21173 ( .A(y[6750]), .B(x[6750]), .Z(n12921) );
  XOR U21174 ( .A(n12915), .B(n12914), .Z(n12925) );
  XOR U21175 ( .A(n12917), .B(n12916), .Z(n12914) );
  XOR U21176 ( .A(y[6749]), .B(x[6749]), .Z(n12916) );
  XOR U21177 ( .A(y[6748]), .B(x[6748]), .Z(n12917) );
  XOR U21178 ( .A(y[6747]), .B(x[6747]), .Z(n12915) );
  XNOR U21179 ( .A(n12891), .B(n12892), .Z(n12909) );
  XNOR U21180 ( .A(n12906), .B(n12907), .Z(n12892) );
  XOR U21181 ( .A(n12903), .B(n12902), .Z(n12907) );
  XOR U21182 ( .A(y[6744]), .B(x[6744]), .Z(n12902) );
  XOR U21183 ( .A(n12905), .B(n12904), .Z(n12903) );
  XOR U21184 ( .A(y[6746]), .B(x[6746]), .Z(n12904) );
  XOR U21185 ( .A(y[6745]), .B(x[6745]), .Z(n12905) );
  XOR U21186 ( .A(n12897), .B(n12896), .Z(n12906) );
  XOR U21187 ( .A(n12899), .B(n12898), .Z(n12896) );
  XOR U21188 ( .A(y[6743]), .B(x[6743]), .Z(n12898) );
  XOR U21189 ( .A(y[6742]), .B(x[6742]), .Z(n12899) );
  XOR U21190 ( .A(y[6741]), .B(x[6741]), .Z(n12897) );
  XNOR U21191 ( .A(n12890), .B(n12889), .Z(n12891) );
  XNOR U21192 ( .A(n12886), .B(n12885), .Z(n12889) );
  XOR U21193 ( .A(n12888), .B(n12887), .Z(n12885) );
  XOR U21194 ( .A(y[6740]), .B(x[6740]), .Z(n12887) );
  XOR U21195 ( .A(y[6739]), .B(x[6739]), .Z(n12888) );
  XOR U21196 ( .A(y[6738]), .B(x[6738]), .Z(n12886) );
  XOR U21197 ( .A(n12880), .B(n12879), .Z(n12890) );
  XOR U21198 ( .A(n12882), .B(n12881), .Z(n12879) );
  XOR U21199 ( .A(y[6737]), .B(x[6737]), .Z(n12881) );
  XOR U21200 ( .A(y[6736]), .B(x[6736]), .Z(n12882) );
  XOR U21201 ( .A(y[6735]), .B(x[6735]), .Z(n12880) );
  NAND U21202 ( .A(n12943), .B(n12944), .Z(N64236) );
  NAND U21203 ( .A(n12945), .B(n12946), .Z(n12944) );
  NANDN U21204 ( .A(n12947), .B(n12948), .Z(n12946) );
  NANDN U21205 ( .A(n12948), .B(n12947), .Z(n12943) );
  XOR U21206 ( .A(n12947), .B(n12949), .Z(N64235) );
  XNOR U21207 ( .A(n12945), .B(n12948), .Z(n12949) );
  NAND U21208 ( .A(n12950), .B(n12951), .Z(n12948) );
  NAND U21209 ( .A(n12952), .B(n12953), .Z(n12951) );
  NANDN U21210 ( .A(n12954), .B(n12955), .Z(n12953) );
  NANDN U21211 ( .A(n12955), .B(n12954), .Z(n12950) );
  AND U21212 ( .A(n12956), .B(n12957), .Z(n12945) );
  NAND U21213 ( .A(n12958), .B(n12959), .Z(n12957) );
  NANDN U21214 ( .A(n12960), .B(n12961), .Z(n12959) );
  NANDN U21215 ( .A(n12961), .B(n12960), .Z(n12956) );
  IV U21216 ( .A(n12962), .Z(n12961) );
  AND U21217 ( .A(n12963), .B(n12964), .Z(n12947) );
  NAND U21218 ( .A(n12965), .B(n12966), .Z(n12964) );
  NANDN U21219 ( .A(n12967), .B(n12968), .Z(n12966) );
  NANDN U21220 ( .A(n12968), .B(n12967), .Z(n12963) );
  XOR U21221 ( .A(n12960), .B(n12969), .Z(N64234) );
  XNOR U21222 ( .A(n12958), .B(n12962), .Z(n12969) );
  XOR U21223 ( .A(n12955), .B(n12970), .Z(n12962) );
  XNOR U21224 ( .A(n12952), .B(n12954), .Z(n12970) );
  AND U21225 ( .A(n12971), .B(n12972), .Z(n12954) );
  NANDN U21226 ( .A(n12973), .B(n12974), .Z(n12972) );
  OR U21227 ( .A(n12975), .B(n12976), .Z(n12974) );
  IV U21228 ( .A(n12977), .Z(n12976) );
  NANDN U21229 ( .A(n12977), .B(n12975), .Z(n12971) );
  AND U21230 ( .A(n12978), .B(n12979), .Z(n12952) );
  NAND U21231 ( .A(n12980), .B(n12981), .Z(n12979) );
  NANDN U21232 ( .A(n12982), .B(n12983), .Z(n12981) );
  NANDN U21233 ( .A(n12983), .B(n12982), .Z(n12978) );
  IV U21234 ( .A(n12984), .Z(n12983) );
  NAND U21235 ( .A(n12985), .B(n12986), .Z(n12955) );
  NANDN U21236 ( .A(n12987), .B(n12988), .Z(n12986) );
  NANDN U21237 ( .A(n12989), .B(n12990), .Z(n12988) );
  NANDN U21238 ( .A(n12990), .B(n12989), .Z(n12985) );
  IV U21239 ( .A(n12991), .Z(n12989) );
  AND U21240 ( .A(n12992), .B(n12993), .Z(n12958) );
  NAND U21241 ( .A(n12994), .B(n12995), .Z(n12993) );
  NANDN U21242 ( .A(n12996), .B(n12997), .Z(n12995) );
  NANDN U21243 ( .A(n12997), .B(n12996), .Z(n12992) );
  XOR U21244 ( .A(n12968), .B(n12998), .Z(n12960) );
  XNOR U21245 ( .A(n12965), .B(n12967), .Z(n12998) );
  AND U21246 ( .A(n12999), .B(n13000), .Z(n12967) );
  NANDN U21247 ( .A(n13001), .B(n13002), .Z(n13000) );
  OR U21248 ( .A(n13003), .B(n13004), .Z(n13002) );
  IV U21249 ( .A(n13005), .Z(n13004) );
  NANDN U21250 ( .A(n13005), .B(n13003), .Z(n12999) );
  AND U21251 ( .A(n13006), .B(n13007), .Z(n12965) );
  NAND U21252 ( .A(n13008), .B(n13009), .Z(n13007) );
  NANDN U21253 ( .A(n13010), .B(n13011), .Z(n13009) );
  NANDN U21254 ( .A(n13011), .B(n13010), .Z(n13006) );
  IV U21255 ( .A(n13012), .Z(n13011) );
  NAND U21256 ( .A(n13013), .B(n13014), .Z(n12968) );
  NANDN U21257 ( .A(n13015), .B(n13016), .Z(n13014) );
  NANDN U21258 ( .A(n13017), .B(n13018), .Z(n13016) );
  NANDN U21259 ( .A(n13018), .B(n13017), .Z(n13013) );
  IV U21260 ( .A(n13019), .Z(n13017) );
  XOR U21261 ( .A(n12994), .B(n13020), .Z(N64233) );
  XNOR U21262 ( .A(n12997), .B(n12996), .Z(n13020) );
  XNOR U21263 ( .A(n13008), .B(n13021), .Z(n12996) );
  XNOR U21264 ( .A(n13012), .B(n13010), .Z(n13021) );
  XOR U21265 ( .A(n13018), .B(n13022), .Z(n13010) );
  XNOR U21266 ( .A(n13015), .B(n13019), .Z(n13022) );
  AND U21267 ( .A(n13023), .B(n13024), .Z(n13019) );
  NAND U21268 ( .A(n13025), .B(n13026), .Z(n13024) );
  NAND U21269 ( .A(n13027), .B(n13028), .Z(n13023) );
  AND U21270 ( .A(n13029), .B(n13030), .Z(n13015) );
  NAND U21271 ( .A(n13031), .B(n13032), .Z(n13030) );
  NAND U21272 ( .A(n13033), .B(n13034), .Z(n13029) );
  NANDN U21273 ( .A(n13035), .B(n13036), .Z(n13018) );
  ANDN U21274 ( .B(n13037), .A(n13038), .Z(n13012) );
  XNOR U21275 ( .A(n13003), .B(n13039), .Z(n13008) );
  XNOR U21276 ( .A(n13001), .B(n13005), .Z(n13039) );
  AND U21277 ( .A(n13040), .B(n13041), .Z(n13005) );
  NAND U21278 ( .A(n13042), .B(n13043), .Z(n13041) );
  NAND U21279 ( .A(n13044), .B(n13045), .Z(n13040) );
  AND U21280 ( .A(n13046), .B(n13047), .Z(n13001) );
  NAND U21281 ( .A(n13048), .B(n13049), .Z(n13047) );
  NAND U21282 ( .A(n13050), .B(n13051), .Z(n13046) );
  AND U21283 ( .A(n13052), .B(n13053), .Z(n13003) );
  NAND U21284 ( .A(n13054), .B(n13055), .Z(n12997) );
  XNOR U21285 ( .A(n12980), .B(n13056), .Z(n12994) );
  XNOR U21286 ( .A(n12984), .B(n12982), .Z(n13056) );
  XOR U21287 ( .A(n12990), .B(n13057), .Z(n12982) );
  XNOR U21288 ( .A(n12987), .B(n12991), .Z(n13057) );
  AND U21289 ( .A(n13058), .B(n13059), .Z(n12991) );
  NAND U21290 ( .A(n13060), .B(n13061), .Z(n13059) );
  NAND U21291 ( .A(n13062), .B(n13063), .Z(n13058) );
  AND U21292 ( .A(n13064), .B(n13065), .Z(n12987) );
  NAND U21293 ( .A(n13066), .B(n13067), .Z(n13065) );
  NAND U21294 ( .A(n13068), .B(n13069), .Z(n13064) );
  NANDN U21295 ( .A(n13070), .B(n13071), .Z(n12990) );
  ANDN U21296 ( .B(n13072), .A(n13073), .Z(n12984) );
  XNOR U21297 ( .A(n12975), .B(n13074), .Z(n12980) );
  XNOR U21298 ( .A(n12973), .B(n12977), .Z(n13074) );
  AND U21299 ( .A(n13075), .B(n13076), .Z(n12977) );
  NAND U21300 ( .A(n13077), .B(n13078), .Z(n13076) );
  NAND U21301 ( .A(n13079), .B(n13080), .Z(n13075) );
  AND U21302 ( .A(n13081), .B(n13082), .Z(n12973) );
  NAND U21303 ( .A(n13083), .B(n13084), .Z(n13082) );
  NAND U21304 ( .A(n13085), .B(n13086), .Z(n13081) );
  AND U21305 ( .A(n13087), .B(n13088), .Z(n12975) );
  XOR U21306 ( .A(n13055), .B(n13054), .Z(N64232) );
  XNOR U21307 ( .A(n13072), .B(n13073), .Z(n13054) );
  XNOR U21308 ( .A(n13087), .B(n13088), .Z(n13073) );
  XOR U21309 ( .A(n13084), .B(n13083), .Z(n13088) );
  XOR U21310 ( .A(y[6732]), .B(x[6732]), .Z(n13083) );
  XOR U21311 ( .A(n13086), .B(n13085), .Z(n13084) );
  XOR U21312 ( .A(y[6734]), .B(x[6734]), .Z(n13085) );
  XOR U21313 ( .A(y[6733]), .B(x[6733]), .Z(n13086) );
  XOR U21314 ( .A(n13078), .B(n13077), .Z(n13087) );
  XOR U21315 ( .A(n13080), .B(n13079), .Z(n13077) );
  XOR U21316 ( .A(y[6731]), .B(x[6731]), .Z(n13079) );
  XOR U21317 ( .A(y[6730]), .B(x[6730]), .Z(n13080) );
  XOR U21318 ( .A(y[6729]), .B(x[6729]), .Z(n13078) );
  XNOR U21319 ( .A(n13071), .B(n13070), .Z(n13072) );
  XNOR U21320 ( .A(n13067), .B(n13066), .Z(n13070) );
  XOR U21321 ( .A(n13069), .B(n13068), .Z(n13066) );
  XOR U21322 ( .A(y[6728]), .B(x[6728]), .Z(n13068) );
  XOR U21323 ( .A(y[6727]), .B(x[6727]), .Z(n13069) );
  XOR U21324 ( .A(y[6726]), .B(x[6726]), .Z(n13067) );
  XOR U21325 ( .A(n13061), .B(n13060), .Z(n13071) );
  XOR U21326 ( .A(n13063), .B(n13062), .Z(n13060) );
  XOR U21327 ( .A(y[6725]), .B(x[6725]), .Z(n13062) );
  XOR U21328 ( .A(y[6724]), .B(x[6724]), .Z(n13063) );
  XOR U21329 ( .A(y[6723]), .B(x[6723]), .Z(n13061) );
  XNOR U21330 ( .A(n13037), .B(n13038), .Z(n13055) );
  XNOR U21331 ( .A(n13052), .B(n13053), .Z(n13038) );
  XOR U21332 ( .A(n13049), .B(n13048), .Z(n13053) );
  XOR U21333 ( .A(y[6720]), .B(x[6720]), .Z(n13048) );
  XOR U21334 ( .A(n13051), .B(n13050), .Z(n13049) );
  XOR U21335 ( .A(y[6722]), .B(x[6722]), .Z(n13050) );
  XOR U21336 ( .A(y[6721]), .B(x[6721]), .Z(n13051) );
  XOR U21337 ( .A(n13043), .B(n13042), .Z(n13052) );
  XOR U21338 ( .A(n13045), .B(n13044), .Z(n13042) );
  XOR U21339 ( .A(y[6719]), .B(x[6719]), .Z(n13044) );
  XOR U21340 ( .A(y[6718]), .B(x[6718]), .Z(n13045) );
  XOR U21341 ( .A(y[6717]), .B(x[6717]), .Z(n13043) );
  XNOR U21342 ( .A(n13036), .B(n13035), .Z(n13037) );
  XNOR U21343 ( .A(n13032), .B(n13031), .Z(n13035) );
  XOR U21344 ( .A(n13034), .B(n13033), .Z(n13031) );
  XOR U21345 ( .A(y[6716]), .B(x[6716]), .Z(n13033) );
  XOR U21346 ( .A(y[6715]), .B(x[6715]), .Z(n13034) );
  XOR U21347 ( .A(y[6714]), .B(x[6714]), .Z(n13032) );
  XOR U21348 ( .A(n13026), .B(n13025), .Z(n13036) );
  XOR U21349 ( .A(n13028), .B(n13027), .Z(n13025) );
  XOR U21350 ( .A(y[6713]), .B(x[6713]), .Z(n13027) );
  XOR U21351 ( .A(y[6712]), .B(x[6712]), .Z(n13028) );
  XOR U21352 ( .A(y[6711]), .B(x[6711]), .Z(n13026) );
  NAND U21353 ( .A(n13089), .B(n13090), .Z(N64223) );
  NAND U21354 ( .A(n13091), .B(n13092), .Z(n13090) );
  NANDN U21355 ( .A(n13093), .B(n13094), .Z(n13092) );
  NANDN U21356 ( .A(n13094), .B(n13093), .Z(n13089) );
  XOR U21357 ( .A(n13093), .B(n13095), .Z(N64222) );
  XNOR U21358 ( .A(n13091), .B(n13094), .Z(n13095) );
  NAND U21359 ( .A(n13096), .B(n13097), .Z(n13094) );
  NAND U21360 ( .A(n13098), .B(n13099), .Z(n13097) );
  NANDN U21361 ( .A(n13100), .B(n13101), .Z(n13099) );
  NANDN U21362 ( .A(n13101), .B(n13100), .Z(n13096) );
  AND U21363 ( .A(n13102), .B(n13103), .Z(n13091) );
  NAND U21364 ( .A(n13104), .B(n13105), .Z(n13103) );
  NANDN U21365 ( .A(n13106), .B(n13107), .Z(n13105) );
  NANDN U21366 ( .A(n13107), .B(n13106), .Z(n13102) );
  IV U21367 ( .A(n13108), .Z(n13107) );
  AND U21368 ( .A(n13109), .B(n13110), .Z(n13093) );
  NAND U21369 ( .A(n13111), .B(n13112), .Z(n13110) );
  NANDN U21370 ( .A(n13113), .B(n13114), .Z(n13112) );
  NANDN U21371 ( .A(n13114), .B(n13113), .Z(n13109) );
  XOR U21372 ( .A(n13106), .B(n13115), .Z(N64221) );
  XNOR U21373 ( .A(n13104), .B(n13108), .Z(n13115) );
  XOR U21374 ( .A(n13101), .B(n13116), .Z(n13108) );
  XNOR U21375 ( .A(n13098), .B(n13100), .Z(n13116) );
  AND U21376 ( .A(n13117), .B(n13118), .Z(n13100) );
  NANDN U21377 ( .A(n13119), .B(n13120), .Z(n13118) );
  OR U21378 ( .A(n13121), .B(n13122), .Z(n13120) );
  IV U21379 ( .A(n13123), .Z(n13122) );
  NANDN U21380 ( .A(n13123), .B(n13121), .Z(n13117) );
  AND U21381 ( .A(n13124), .B(n13125), .Z(n13098) );
  NAND U21382 ( .A(n13126), .B(n13127), .Z(n13125) );
  NANDN U21383 ( .A(n13128), .B(n13129), .Z(n13127) );
  NANDN U21384 ( .A(n13129), .B(n13128), .Z(n13124) );
  IV U21385 ( .A(n13130), .Z(n13129) );
  NAND U21386 ( .A(n13131), .B(n13132), .Z(n13101) );
  NANDN U21387 ( .A(n13133), .B(n13134), .Z(n13132) );
  NANDN U21388 ( .A(n13135), .B(n13136), .Z(n13134) );
  NANDN U21389 ( .A(n13136), .B(n13135), .Z(n13131) );
  IV U21390 ( .A(n13137), .Z(n13135) );
  AND U21391 ( .A(n13138), .B(n13139), .Z(n13104) );
  NAND U21392 ( .A(n13140), .B(n13141), .Z(n13139) );
  NANDN U21393 ( .A(n13142), .B(n13143), .Z(n13141) );
  NANDN U21394 ( .A(n13143), .B(n13142), .Z(n13138) );
  XOR U21395 ( .A(n13114), .B(n13144), .Z(n13106) );
  XNOR U21396 ( .A(n13111), .B(n13113), .Z(n13144) );
  AND U21397 ( .A(n13145), .B(n13146), .Z(n13113) );
  NANDN U21398 ( .A(n13147), .B(n13148), .Z(n13146) );
  OR U21399 ( .A(n13149), .B(n13150), .Z(n13148) );
  IV U21400 ( .A(n13151), .Z(n13150) );
  NANDN U21401 ( .A(n13151), .B(n13149), .Z(n13145) );
  AND U21402 ( .A(n13152), .B(n13153), .Z(n13111) );
  NAND U21403 ( .A(n13154), .B(n13155), .Z(n13153) );
  NANDN U21404 ( .A(n13156), .B(n13157), .Z(n13155) );
  NANDN U21405 ( .A(n13157), .B(n13156), .Z(n13152) );
  IV U21406 ( .A(n13158), .Z(n13157) );
  NAND U21407 ( .A(n13159), .B(n13160), .Z(n13114) );
  NANDN U21408 ( .A(n13161), .B(n13162), .Z(n13160) );
  NANDN U21409 ( .A(n13163), .B(n13164), .Z(n13162) );
  NANDN U21410 ( .A(n13164), .B(n13163), .Z(n13159) );
  IV U21411 ( .A(n13165), .Z(n13163) );
  XOR U21412 ( .A(n13140), .B(n13166), .Z(N64220) );
  XNOR U21413 ( .A(n13143), .B(n13142), .Z(n13166) );
  XNOR U21414 ( .A(n13154), .B(n13167), .Z(n13142) );
  XNOR U21415 ( .A(n13158), .B(n13156), .Z(n13167) );
  XOR U21416 ( .A(n13164), .B(n13168), .Z(n13156) );
  XNOR U21417 ( .A(n13161), .B(n13165), .Z(n13168) );
  AND U21418 ( .A(n13169), .B(n13170), .Z(n13165) );
  NAND U21419 ( .A(n13171), .B(n13172), .Z(n13170) );
  NAND U21420 ( .A(n13173), .B(n13174), .Z(n13169) );
  AND U21421 ( .A(n13175), .B(n13176), .Z(n13161) );
  NAND U21422 ( .A(n13177), .B(n13178), .Z(n13176) );
  NAND U21423 ( .A(n13179), .B(n13180), .Z(n13175) );
  NANDN U21424 ( .A(n13181), .B(n13182), .Z(n13164) );
  ANDN U21425 ( .B(n13183), .A(n13184), .Z(n13158) );
  XNOR U21426 ( .A(n13149), .B(n13185), .Z(n13154) );
  XNOR U21427 ( .A(n13147), .B(n13151), .Z(n13185) );
  AND U21428 ( .A(n13186), .B(n13187), .Z(n13151) );
  NAND U21429 ( .A(n13188), .B(n13189), .Z(n13187) );
  NAND U21430 ( .A(n13190), .B(n13191), .Z(n13186) );
  AND U21431 ( .A(n13192), .B(n13193), .Z(n13147) );
  NAND U21432 ( .A(n13194), .B(n13195), .Z(n13193) );
  NAND U21433 ( .A(n13196), .B(n13197), .Z(n13192) );
  AND U21434 ( .A(n13198), .B(n13199), .Z(n13149) );
  NAND U21435 ( .A(n13200), .B(n13201), .Z(n13143) );
  XNOR U21436 ( .A(n13126), .B(n13202), .Z(n13140) );
  XNOR U21437 ( .A(n13130), .B(n13128), .Z(n13202) );
  XOR U21438 ( .A(n13136), .B(n13203), .Z(n13128) );
  XNOR U21439 ( .A(n13133), .B(n13137), .Z(n13203) );
  AND U21440 ( .A(n13204), .B(n13205), .Z(n13137) );
  NAND U21441 ( .A(n13206), .B(n13207), .Z(n13205) );
  NAND U21442 ( .A(n13208), .B(n13209), .Z(n13204) );
  AND U21443 ( .A(n13210), .B(n13211), .Z(n13133) );
  NAND U21444 ( .A(n13212), .B(n13213), .Z(n13211) );
  NAND U21445 ( .A(n13214), .B(n13215), .Z(n13210) );
  NANDN U21446 ( .A(n13216), .B(n13217), .Z(n13136) );
  ANDN U21447 ( .B(n13218), .A(n13219), .Z(n13130) );
  XNOR U21448 ( .A(n13121), .B(n13220), .Z(n13126) );
  XNOR U21449 ( .A(n13119), .B(n13123), .Z(n13220) );
  AND U21450 ( .A(n13221), .B(n13222), .Z(n13123) );
  NAND U21451 ( .A(n13223), .B(n13224), .Z(n13222) );
  NAND U21452 ( .A(n13225), .B(n13226), .Z(n13221) );
  AND U21453 ( .A(n13227), .B(n13228), .Z(n13119) );
  NAND U21454 ( .A(n13229), .B(n13230), .Z(n13228) );
  NAND U21455 ( .A(n13231), .B(n13232), .Z(n13227) );
  AND U21456 ( .A(n13233), .B(n13234), .Z(n13121) );
  XOR U21457 ( .A(n13201), .B(n13200), .Z(N64219) );
  XNOR U21458 ( .A(n13218), .B(n13219), .Z(n13200) );
  XNOR U21459 ( .A(n13233), .B(n13234), .Z(n13219) );
  XOR U21460 ( .A(n13230), .B(n13229), .Z(n13234) );
  XOR U21461 ( .A(y[6708]), .B(x[6708]), .Z(n13229) );
  XOR U21462 ( .A(n13232), .B(n13231), .Z(n13230) );
  XOR U21463 ( .A(y[6710]), .B(x[6710]), .Z(n13231) );
  XOR U21464 ( .A(y[6709]), .B(x[6709]), .Z(n13232) );
  XOR U21465 ( .A(n13224), .B(n13223), .Z(n13233) );
  XOR U21466 ( .A(n13226), .B(n13225), .Z(n13223) );
  XOR U21467 ( .A(y[6707]), .B(x[6707]), .Z(n13225) );
  XOR U21468 ( .A(y[6706]), .B(x[6706]), .Z(n13226) );
  XOR U21469 ( .A(y[6705]), .B(x[6705]), .Z(n13224) );
  XNOR U21470 ( .A(n13217), .B(n13216), .Z(n13218) );
  XNOR U21471 ( .A(n13213), .B(n13212), .Z(n13216) );
  XOR U21472 ( .A(n13215), .B(n13214), .Z(n13212) );
  XOR U21473 ( .A(y[6704]), .B(x[6704]), .Z(n13214) );
  XOR U21474 ( .A(y[6703]), .B(x[6703]), .Z(n13215) );
  XOR U21475 ( .A(y[6702]), .B(x[6702]), .Z(n13213) );
  XOR U21476 ( .A(n13207), .B(n13206), .Z(n13217) );
  XOR U21477 ( .A(n13209), .B(n13208), .Z(n13206) );
  XOR U21478 ( .A(y[6701]), .B(x[6701]), .Z(n13208) );
  XOR U21479 ( .A(y[6700]), .B(x[6700]), .Z(n13209) );
  XOR U21480 ( .A(y[6699]), .B(x[6699]), .Z(n13207) );
  XNOR U21481 ( .A(n13183), .B(n13184), .Z(n13201) );
  XNOR U21482 ( .A(n13198), .B(n13199), .Z(n13184) );
  XOR U21483 ( .A(n13195), .B(n13194), .Z(n13199) );
  XOR U21484 ( .A(y[6696]), .B(x[6696]), .Z(n13194) );
  XOR U21485 ( .A(n13197), .B(n13196), .Z(n13195) );
  XOR U21486 ( .A(y[6698]), .B(x[6698]), .Z(n13196) );
  XOR U21487 ( .A(y[6697]), .B(x[6697]), .Z(n13197) );
  XOR U21488 ( .A(n13189), .B(n13188), .Z(n13198) );
  XOR U21489 ( .A(n13191), .B(n13190), .Z(n13188) );
  XOR U21490 ( .A(y[6695]), .B(x[6695]), .Z(n13190) );
  XOR U21491 ( .A(y[6694]), .B(x[6694]), .Z(n13191) );
  XOR U21492 ( .A(y[6693]), .B(x[6693]), .Z(n13189) );
  XNOR U21493 ( .A(n13182), .B(n13181), .Z(n13183) );
  XNOR U21494 ( .A(n13178), .B(n13177), .Z(n13181) );
  XOR U21495 ( .A(n13180), .B(n13179), .Z(n13177) );
  XOR U21496 ( .A(y[6692]), .B(x[6692]), .Z(n13179) );
  XOR U21497 ( .A(y[6691]), .B(x[6691]), .Z(n13180) );
  XOR U21498 ( .A(y[6690]), .B(x[6690]), .Z(n13178) );
  XOR U21499 ( .A(n13172), .B(n13171), .Z(n13182) );
  XOR U21500 ( .A(n13174), .B(n13173), .Z(n13171) );
  XOR U21501 ( .A(y[6689]), .B(x[6689]), .Z(n13173) );
  XOR U21502 ( .A(y[6688]), .B(x[6688]), .Z(n13174) );
  XOR U21503 ( .A(y[6687]), .B(x[6687]), .Z(n13172) );
  NAND U21504 ( .A(n13235), .B(n13236), .Z(N64210) );
  NAND U21505 ( .A(n13237), .B(n13238), .Z(n13236) );
  NANDN U21506 ( .A(n13239), .B(n13240), .Z(n13238) );
  NANDN U21507 ( .A(n13240), .B(n13239), .Z(n13235) );
  XOR U21508 ( .A(n13239), .B(n13241), .Z(N64209) );
  XNOR U21509 ( .A(n13237), .B(n13240), .Z(n13241) );
  NAND U21510 ( .A(n13242), .B(n13243), .Z(n13240) );
  NAND U21511 ( .A(n13244), .B(n13245), .Z(n13243) );
  NANDN U21512 ( .A(n13246), .B(n13247), .Z(n13245) );
  NANDN U21513 ( .A(n13247), .B(n13246), .Z(n13242) );
  AND U21514 ( .A(n13248), .B(n13249), .Z(n13237) );
  NAND U21515 ( .A(n13250), .B(n13251), .Z(n13249) );
  NANDN U21516 ( .A(n13252), .B(n13253), .Z(n13251) );
  NANDN U21517 ( .A(n13253), .B(n13252), .Z(n13248) );
  IV U21518 ( .A(n13254), .Z(n13253) );
  AND U21519 ( .A(n13255), .B(n13256), .Z(n13239) );
  NAND U21520 ( .A(n13257), .B(n13258), .Z(n13256) );
  NANDN U21521 ( .A(n13259), .B(n13260), .Z(n13258) );
  NANDN U21522 ( .A(n13260), .B(n13259), .Z(n13255) );
  XOR U21523 ( .A(n13252), .B(n13261), .Z(N64208) );
  XNOR U21524 ( .A(n13250), .B(n13254), .Z(n13261) );
  XOR U21525 ( .A(n13247), .B(n13262), .Z(n13254) );
  XNOR U21526 ( .A(n13244), .B(n13246), .Z(n13262) );
  AND U21527 ( .A(n13263), .B(n13264), .Z(n13246) );
  NANDN U21528 ( .A(n13265), .B(n13266), .Z(n13264) );
  OR U21529 ( .A(n13267), .B(n13268), .Z(n13266) );
  IV U21530 ( .A(n13269), .Z(n13268) );
  NANDN U21531 ( .A(n13269), .B(n13267), .Z(n13263) );
  AND U21532 ( .A(n13270), .B(n13271), .Z(n13244) );
  NAND U21533 ( .A(n13272), .B(n13273), .Z(n13271) );
  NANDN U21534 ( .A(n13274), .B(n13275), .Z(n13273) );
  NANDN U21535 ( .A(n13275), .B(n13274), .Z(n13270) );
  IV U21536 ( .A(n13276), .Z(n13275) );
  NAND U21537 ( .A(n13277), .B(n13278), .Z(n13247) );
  NANDN U21538 ( .A(n13279), .B(n13280), .Z(n13278) );
  NANDN U21539 ( .A(n13281), .B(n13282), .Z(n13280) );
  NANDN U21540 ( .A(n13282), .B(n13281), .Z(n13277) );
  IV U21541 ( .A(n13283), .Z(n13281) );
  AND U21542 ( .A(n13284), .B(n13285), .Z(n13250) );
  NAND U21543 ( .A(n13286), .B(n13287), .Z(n13285) );
  NANDN U21544 ( .A(n13288), .B(n13289), .Z(n13287) );
  NANDN U21545 ( .A(n13289), .B(n13288), .Z(n13284) );
  XOR U21546 ( .A(n13260), .B(n13290), .Z(n13252) );
  XNOR U21547 ( .A(n13257), .B(n13259), .Z(n13290) );
  AND U21548 ( .A(n13291), .B(n13292), .Z(n13259) );
  NANDN U21549 ( .A(n13293), .B(n13294), .Z(n13292) );
  OR U21550 ( .A(n13295), .B(n13296), .Z(n13294) );
  IV U21551 ( .A(n13297), .Z(n13296) );
  NANDN U21552 ( .A(n13297), .B(n13295), .Z(n13291) );
  AND U21553 ( .A(n13298), .B(n13299), .Z(n13257) );
  NAND U21554 ( .A(n13300), .B(n13301), .Z(n13299) );
  NANDN U21555 ( .A(n13302), .B(n13303), .Z(n13301) );
  NANDN U21556 ( .A(n13303), .B(n13302), .Z(n13298) );
  IV U21557 ( .A(n13304), .Z(n13303) );
  NAND U21558 ( .A(n13305), .B(n13306), .Z(n13260) );
  NANDN U21559 ( .A(n13307), .B(n13308), .Z(n13306) );
  NANDN U21560 ( .A(n13309), .B(n13310), .Z(n13308) );
  NANDN U21561 ( .A(n13310), .B(n13309), .Z(n13305) );
  IV U21562 ( .A(n13311), .Z(n13309) );
  XOR U21563 ( .A(n13286), .B(n13312), .Z(N64207) );
  XNOR U21564 ( .A(n13289), .B(n13288), .Z(n13312) );
  XNOR U21565 ( .A(n13300), .B(n13313), .Z(n13288) );
  XNOR U21566 ( .A(n13304), .B(n13302), .Z(n13313) );
  XOR U21567 ( .A(n13310), .B(n13314), .Z(n13302) );
  XNOR U21568 ( .A(n13307), .B(n13311), .Z(n13314) );
  AND U21569 ( .A(n13315), .B(n13316), .Z(n13311) );
  NAND U21570 ( .A(n13317), .B(n13318), .Z(n13316) );
  NAND U21571 ( .A(n13319), .B(n13320), .Z(n13315) );
  AND U21572 ( .A(n13321), .B(n13322), .Z(n13307) );
  NAND U21573 ( .A(n13323), .B(n13324), .Z(n13322) );
  NAND U21574 ( .A(n13325), .B(n13326), .Z(n13321) );
  NANDN U21575 ( .A(n13327), .B(n13328), .Z(n13310) );
  ANDN U21576 ( .B(n13329), .A(n13330), .Z(n13304) );
  XNOR U21577 ( .A(n13295), .B(n13331), .Z(n13300) );
  XNOR U21578 ( .A(n13293), .B(n13297), .Z(n13331) );
  AND U21579 ( .A(n13332), .B(n13333), .Z(n13297) );
  NAND U21580 ( .A(n13334), .B(n13335), .Z(n13333) );
  NAND U21581 ( .A(n13336), .B(n13337), .Z(n13332) );
  AND U21582 ( .A(n13338), .B(n13339), .Z(n13293) );
  NAND U21583 ( .A(n13340), .B(n13341), .Z(n13339) );
  NAND U21584 ( .A(n13342), .B(n13343), .Z(n13338) );
  AND U21585 ( .A(n13344), .B(n13345), .Z(n13295) );
  NAND U21586 ( .A(n13346), .B(n13347), .Z(n13289) );
  XNOR U21587 ( .A(n13272), .B(n13348), .Z(n13286) );
  XNOR U21588 ( .A(n13276), .B(n13274), .Z(n13348) );
  XOR U21589 ( .A(n13282), .B(n13349), .Z(n13274) );
  XNOR U21590 ( .A(n13279), .B(n13283), .Z(n13349) );
  AND U21591 ( .A(n13350), .B(n13351), .Z(n13283) );
  NAND U21592 ( .A(n13352), .B(n13353), .Z(n13351) );
  NAND U21593 ( .A(n13354), .B(n13355), .Z(n13350) );
  AND U21594 ( .A(n13356), .B(n13357), .Z(n13279) );
  NAND U21595 ( .A(n13358), .B(n13359), .Z(n13357) );
  NAND U21596 ( .A(n13360), .B(n13361), .Z(n13356) );
  NANDN U21597 ( .A(n13362), .B(n13363), .Z(n13282) );
  ANDN U21598 ( .B(n13364), .A(n13365), .Z(n13276) );
  XNOR U21599 ( .A(n13267), .B(n13366), .Z(n13272) );
  XNOR U21600 ( .A(n13265), .B(n13269), .Z(n13366) );
  AND U21601 ( .A(n13367), .B(n13368), .Z(n13269) );
  NAND U21602 ( .A(n13369), .B(n13370), .Z(n13368) );
  NAND U21603 ( .A(n13371), .B(n13372), .Z(n13367) );
  AND U21604 ( .A(n13373), .B(n13374), .Z(n13265) );
  NAND U21605 ( .A(n13375), .B(n13376), .Z(n13374) );
  NAND U21606 ( .A(n13377), .B(n13378), .Z(n13373) );
  AND U21607 ( .A(n13379), .B(n13380), .Z(n13267) );
  XOR U21608 ( .A(n13347), .B(n13346), .Z(N64206) );
  XNOR U21609 ( .A(n13364), .B(n13365), .Z(n13346) );
  XNOR U21610 ( .A(n13379), .B(n13380), .Z(n13365) );
  XOR U21611 ( .A(n13376), .B(n13375), .Z(n13380) );
  XOR U21612 ( .A(y[6684]), .B(x[6684]), .Z(n13375) );
  XOR U21613 ( .A(n13378), .B(n13377), .Z(n13376) );
  XOR U21614 ( .A(y[6686]), .B(x[6686]), .Z(n13377) );
  XOR U21615 ( .A(y[6685]), .B(x[6685]), .Z(n13378) );
  XOR U21616 ( .A(n13370), .B(n13369), .Z(n13379) );
  XOR U21617 ( .A(n13372), .B(n13371), .Z(n13369) );
  XOR U21618 ( .A(y[6683]), .B(x[6683]), .Z(n13371) );
  XOR U21619 ( .A(y[6682]), .B(x[6682]), .Z(n13372) );
  XOR U21620 ( .A(y[6681]), .B(x[6681]), .Z(n13370) );
  XNOR U21621 ( .A(n13363), .B(n13362), .Z(n13364) );
  XNOR U21622 ( .A(n13359), .B(n13358), .Z(n13362) );
  XOR U21623 ( .A(n13361), .B(n13360), .Z(n13358) );
  XOR U21624 ( .A(y[6680]), .B(x[6680]), .Z(n13360) );
  XOR U21625 ( .A(y[6679]), .B(x[6679]), .Z(n13361) );
  XOR U21626 ( .A(y[6678]), .B(x[6678]), .Z(n13359) );
  XOR U21627 ( .A(n13353), .B(n13352), .Z(n13363) );
  XOR U21628 ( .A(n13355), .B(n13354), .Z(n13352) );
  XOR U21629 ( .A(y[6677]), .B(x[6677]), .Z(n13354) );
  XOR U21630 ( .A(y[6676]), .B(x[6676]), .Z(n13355) );
  XOR U21631 ( .A(y[6675]), .B(x[6675]), .Z(n13353) );
  XNOR U21632 ( .A(n13329), .B(n13330), .Z(n13347) );
  XNOR U21633 ( .A(n13344), .B(n13345), .Z(n13330) );
  XOR U21634 ( .A(n13341), .B(n13340), .Z(n13345) );
  XOR U21635 ( .A(y[6672]), .B(x[6672]), .Z(n13340) );
  XOR U21636 ( .A(n13343), .B(n13342), .Z(n13341) );
  XOR U21637 ( .A(y[6674]), .B(x[6674]), .Z(n13342) );
  XOR U21638 ( .A(y[6673]), .B(x[6673]), .Z(n13343) );
  XOR U21639 ( .A(n13335), .B(n13334), .Z(n13344) );
  XOR U21640 ( .A(n13337), .B(n13336), .Z(n13334) );
  XOR U21641 ( .A(y[6671]), .B(x[6671]), .Z(n13336) );
  XOR U21642 ( .A(y[6670]), .B(x[6670]), .Z(n13337) );
  XOR U21643 ( .A(y[6669]), .B(x[6669]), .Z(n13335) );
  XNOR U21644 ( .A(n13328), .B(n13327), .Z(n13329) );
  XNOR U21645 ( .A(n13324), .B(n13323), .Z(n13327) );
  XOR U21646 ( .A(n13326), .B(n13325), .Z(n13323) );
  XOR U21647 ( .A(y[6668]), .B(x[6668]), .Z(n13325) );
  XOR U21648 ( .A(y[6667]), .B(x[6667]), .Z(n13326) );
  XOR U21649 ( .A(y[6666]), .B(x[6666]), .Z(n13324) );
  XOR U21650 ( .A(n13318), .B(n13317), .Z(n13328) );
  XOR U21651 ( .A(n13320), .B(n13319), .Z(n13317) );
  XOR U21652 ( .A(y[6665]), .B(x[6665]), .Z(n13319) );
  XOR U21653 ( .A(y[6664]), .B(x[6664]), .Z(n13320) );
  XOR U21654 ( .A(y[6663]), .B(x[6663]), .Z(n13318) );
  NAND U21655 ( .A(n13381), .B(n13382), .Z(N64197) );
  NAND U21656 ( .A(n13383), .B(n13384), .Z(n13382) );
  NANDN U21657 ( .A(n13385), .B(n13386), .Z(n13384) );
  NANDN U21658 ( .A(n13386), .B(n13385), .Z(n13381) );
  XOR U21659 ( .A(n13385), .B(n13387), .Z(N64196) );
  XNOR U21660 ( .A(n13383), .B(n13386), .Z(n13387) );
  NAND U21661 ( .A(n13388), .B(n13389), .Z(n13386) );
  NAND U21662 ( .A(n13390), .B(n13391), .Z(n13389) );
  NANDN U21663 ( .A(n13392), .B(n13393), .Z(n13391) );
  NANDN U21664 ( .A(n13393), .B(n13392), .Z(n13388) );
  AND U21665 ( .A(n13394), .B(n13395), .Z(n13383) );
  NAND U21666 ( .A(n13396), .B(n13397), .Z(n13395) );
  NANDN U21667 ( .A(n13398), .B(n13399), .Z(n13397) );
  NANDN U21668 ( .A(n13399), .B(n13398), .Z(n13394) );
  IV U21669 ( .A(n13400), .Z(n13399) );
  AND U21670 ( .A(n13401), .B(n13402), .Z(n13385) );
  NAND U21671 ( .A(n13403), .B(n13404), .Z(n13402) );
  NANDN U21672 ( .A(n13405), .B(n13406), .Z(n13404) );
  NANDN U21673 ( .A(n13406), .B(n13405), .Z(n13401) );
  XOR U21674 ( .A(n13398), .B(n13407), .Z(N64195) );
  XNOR U21675 ( .A(n13396), .B(n13400), .Z(n13407) );
  XOR U21676 ( .A(n13393), .B(n13408), .Z(n13400) );
  XNOR U21677 ( .A(n13390), .B(n13392), .Z(n13408) );
  AND U21678 ( .A(n13409), .B(n13410), .Z(n13392) );
  NANDN U21679 ( .A(n13411), .B(n13412), .Z(n13410) );
  OR U21680 ( .A(n13413), .B(n13414), .Z(n13412) );
  IV U21681 ( .A(n13415), .Z(n13414) );
  NANDN U21682 ( .A(n13415), .B(n13413), .Z(n13409) );
  AND U21683 ( .A(n13416), .B(n13417), .Z(n13390) );
  NAND U21684 ( .A(n13418), .B(n13419), .Z(n13417) );
  NANDN U21685 ( .A(n13420), .B(n13421), .Z(n13419) );
  NANDN U21686 ( .A(n13421), .B(n13420), .Z(n13416) );
  IV U21687 ( .A(n13422), .Z(n13421) );
  NAND U21688 ( .A(n13423), .B(n13424), .Z(n13393) );
  NANDN U21689 ( .A(n13425), .B(n13426), .Z(n13424) );
  NANDN U21690 ( .A(n13427), .B(n13428), .Z(n13426) );
  NANDN U21691 ( .A(n13428), .B(n13427), .Z(n13423) );
  IV U21692 ( .A(n13429), .Z(n13427) );
  AND U21693 ( .A(n13430), .B(n13431), .Z(n13396) );
  NAND U21694 ( .A(n13432), .B(n13433), .Z(n13431) );
  NANDN U21695 ( .A(n13434), .B(n13435), .Z(n13433) );
  NANDN U21696 ( .A(n13435), .B(n13434), .Z(n13430) );
  XOR U21697 ( .A(n13406), .B(n13436), .Z(n13398) );
  XNOR U21698 ( .A(n13403), .B(n13405), .Z(n13436) );
  AND U21699 ( .A(n13437), .B(n13438), .Z(n13405) );
  NANDN U21700 ( .A(n13439), .B(n13440), .Z(n13438) );
  OR U21701 ( .A(n13441), .B(n13442), .Z(n13440) );
  IV U21702 ( .A(n13443), .Z(n13442) );
  NANDN U21703 ( .A(n13443), .B(n13441), .Z(n13437) );
  AND U21704 ( .A(n13444), .B(n13445), .Z(n13403) );
  NAND U21705 ( .A(n13446), .B(n13447), .Z(n13445) );
  NANDN U21706 ( .A(n13448), .B(n13449), .Z(n13447) );
  NANDN U21707 ( .A(n13449), .B(n13448), .Z(n13444) );
  IV U21708 ( .A(n13450), .Z(n13449) );
  NAND U21709 ( .A(n13451), .B(n13452), .Z(n13406) );
  NANDN U21710 ( .A(n13453), .B(n13454), .Z(n13452) );
  NANDN U21711 ( .A(n13455), .B(n13456), .Z(n13454) );
  NANDN U21712 ( .A(n13456), .B(n13455), .Z(n13451) );
  IV U21713 ( .A(n13457), .Z(n13455) );
  XOR U21714 ( .A(n13432), .B(n13458), .Z(N64194) );
  XNOR U21715 ( .A(n13435), .B(n13434), .Z(n13458) );
  XNOR U21716 ( .A(n13446), .B(n13459), .Z(n13434) );
  XNOR U21717 ( .A(n13450), .B(n13448), .Z(n13459) );
  XOR U21718 ( .A(n13456), .B(n13460), .Z(n13448) );
  XNOR U21719 ( .A(n13453), .B(n13457), .Z(n13460) );
  AND U21720 ( .A(n13461), .B(n13462), .Z(n13457) );
  NAND U21721 ( .A(n13463), .B(n13464), .Z(n13462) );
  NAND U21722 ( .A(n13465), .B(n13466), .Z(n13461) );
  AND U21723 ( .A(n13467), .B(n13468), .Z(n13453) );
  NAND U21724 ( .A(n13469), .B(n13470), .Z(n13468) );
  NAND U21725 ( .A(n13471), .B(n13472), .Z(n13467) );
  NANDN U21726 ( .A(n13473), .B(n13474), .Z(n13456) );
  ANDN U21727 ( .B(n13475), .A(n13476), .Z(n13450) );
  XNOR U21728 ( .A(n13441), .B(n13477), .Z(n13446) );
  XNOR U21729 ( .A(n13439), .B(n13443), .Z(n13477) );
  AND U21730 ( .A(n13478), .B(n13479), .Z(n13443) );
  NAND U21731 ( .A(n13480), .B(n13481), .Z(n13479) );
  NAND U21732 ( .A(n13482), .B(n13483), .Z(n13478) );
  AND U21733 ( .A(n13484), .B(n13485), .Z(n13439) );
  NAND U21734 ( .A(n13486), .B(n13487), .Z(n13485) );
  NAND U21735 ( .A(n13488), .B(n13489), .Z(n13484) );
  AND U21736 ( .A(n13490), .B(n13491), .Z(n13441) );
  NAND U21737 ( .A(n13492), .B(n13493), .Z(n13435) );
  XNOR U21738 ( .A(n13418), .B(n13494), .Z(n13432) );
  XNOR U21739 ( .A(n13422), .B(n13420), .Z(n13494) );
  XOR U21740 ( .A(n13428), .B(n13495), .Z(n13420) );
  XNOR U21741 ( .A(n13425), .B(n13429), .Z(n13495) );
  AND U21742 ( .A(n13496), .B(n13497), .Z(n13429) );
  NAND U21743 ( .A(n13498), .B(n13499), .Z(n13497) );
  NAND U21744 ( .A(n13500), .B(n13501), .Z(n13496) );
  AND U21745 ( .A(n13502), .B(n13503), .Z(n13425) );
  NAND U21746 ( .A(n13504), .B(n13505), .Z(n13503) );
  NAND U21747 ( .A(n13506), .B(n13507), .Z(n13502) );
  NANDN U21748 ( .A(n13508), .B(n13509), .Z(n13428) );
  ANDN U21749 ( .B(n13510), .A(n13511), .Z(n13422) );
  XNOR U21750 ( .A(n13413), .B(n13512), .Z(n13418) );
  XNOR U21751 ( .A(n13411), .B(n13415), .Z(n13512) );
  AND U21752 ( .A(n13513), .B(n13514), .Z(n13415) );
  NAND U21753 ( .A(n13515), .B(n13516), .Z(n13514) );
  NAND U21754 ( .A(n13517), .B(n13518), .Z(n13513) );
  AND U21755 ( .A(n13519), .B(n13520), .Z(n13411) );
  NAND U21756 ( .A(n13521), .B(n13522), .Z(n13520) );
  NAND U21757 ( .A(n13523), .B(n13524), .Z(n13519) );
  AND U21758 ( .A(n13525), .B(n13526), .Z(n13413) );
  XOR U21759 ( .A(n13493), .B(n13492), .Z(N64193) );
  XNOR U21760 ( .A(n13510), .B(n13511), .Z(n13492) );
  XNOR U21761 ( .A(n13525), .B(n13526), .Z(n13511) );
  XOR U21762 ( .A(n13522), .B(n13521), .Z(n13526) );
  XOR U21763 ( .A(y[6660]), .B(x[6660]), .Z(n13521) );
  XOR U21764 ( .A(n13524), .B(n13523), .Z(n13522) );
  XOR U21765 ( .A(y[6662]), .B(x[6662]), .Z(n13523) );
  XOR U21766 ( .A(y[6661]), .B(x[6661]), .Z(n13524) );
  XOR U21767 ( .A(n13516), .B(n13515), .Z(n13525) );
  XOR U21768 ( .A(n13518), .B(n13517), .Z(n13515) );
  XOR U21769 ( .A(y[6659]), .B(x[6659]), .Z(n13517) );
  XOR U21770 ( .A(y[6658]), .B(x[6658]), .Z(n13518) );
  XOR U21771 ( .A(y[6657]), .B(x[6657]), .Z(n13516) );
  XNOR U21772 ( .A(n13509), .B(n13508), .Z(n13510) );
  XNOR U21773 ( .A(n13505), .B(n13504), .Z(n13508) );
  XOR U21774 ( .A(n13507), .B(n13506), .Z(n13504) );
  XOR U21775 ( .A(y[6656]), .B(x[6656]), .Z(n13506) );
  XOR U21776 ( .A(y[6655]), .B(x[6655]), .Z(n13507) );
  XOR U21777 ( .A(y[6654]), .B(x[6654]), .Z(n13505) );
  XOR U21778 ( .A(n13499), .B(n13498), .Z(n13509) );
  XOR U21779 ( .A(n13501), .B(n13500), .Z(n13498) );
  XOR U21780 ( .A(y[6653]), .B(x[6653]), .Z(n13500) );
  XOR U21781 ( .A(y[6652]), .B(x[6652]), .Z(n13501) );
  XOR U21782 ( .A(y[6651]), .B(x[6651]), .Z(n13499) );
  XNOR U21783 ( .A(n13475), .B(n13476), .Z(n13493) );
  XNOR U21784 ( .A(n13490), .B(n13491), .Z(n13476) );
  XOR U21785 ( .A(n13487), .B(n13486), .Z(n13491) );
  XOR U21786 ( .A(y[6648]), .B(x[6648]), .Z(n13486) );
  XOR U21787 ( .A(n13489), .B(n13488), .Z(n13487) );
  XOR U21788 ( .A(y[6650]), .B(x[6650]), .Z(n13488) );
  XOR U21789 ( .A(y[6649]), .B(x[6649]), .Z(n13489) );
  XOR U21790 ( .A(n13481), .B(n13480), .Z(n13490) );
  XOR U21791 ( .A(n13483), .B(n13482), .Z(n13480) );
  XOR U21792 ( .A(y[6647]), .B(x[6647]), .Z(n13482) );
  XOR U21793 ( .A(y[6646]), .B(x[6646]), .Z(n13483) );
  XOR U21794 ( .A(y[6645]), .B(x[6645]), .Z(n13481) );
  XNOR U21795 ( .A(n13474), .B(n13473), .Z(n13475) );
  XNOR U21796 ( .A(n13470), .B(n13469), .Z(n13473) );
  XOR U21797 ( .A(n13472), .B(n13471), .Z(n13469) );
  XOR U21798 ( .A(y[6644]), .B(x[6644]), .Z(n13471) );
  XOR U21799 ( .A(y[6643]), .B(x[6643]), .Z(n13472) );
  XOR U21800 ( .A(y[6642]), .B(x[6642]), .Z(n13470) );
  XOR U21801 ( .A(n13464), .B(n13463), .Z(n13474) );
  XOR U21802 ( .A(n13466), .B(n13465), .Z(n13463) );
  XOR U21803 ( .A(y[6641]), .B(x[6641]), .Z(n13465) );
  XOR U21804 ( .A(y[6640]), .B(x[6640]), .Z(n13466) );
  XOR U21805 ( .A(y[6639]), .B(x[6639]), .Z(n13464) );
  NAND U21806 ( .A(n13527), .B(n13528), .Z(N64184) );
  NAND U21807 ( .A(n13529), .B(n13530), .Z(n13528) );
  NANDN U21808 ( .A(n13531), .B(n13532), .Z(n13530) );
  NANDN U21809 ( .A(n13532), .B(n13531), .Z(n13527) );
  XOR U21810 ( .A(n13531), .B(n13533), .Z(N64183) );
  XNOR U21811 ( .A(n13529), .B(n13532), .Z(n13533) );
  NAND U21812 ( .A(n13534), .B(n13535), .Z(n13532) );
  NAND U21813 ( .A(n13536), .B(n13537), .Z(n13535) );
  NANDN U21814 ( .A(n13538), .B(n13539), .Z(n13537) );
  NANDN U21815 ( .A(n13539), .B(n13538), .Z(n13534) );
  AND U21816 ( .A(n13540), .B(n13541), .Z(n13529) );
  NAND U21817 ( .A(n13542), .B(n13543), .Z(n13541) );
  NANDN U21818 ( .A(n13544), .B(n13545), .Z(n13543) );
  NANDN U21819 ( .A(n13545), .B(n13544), .Z(n13540) );
  IV U21820 ( .A(n13546), .Z(n13545) );
  AND U21821 ( .A(n13547), .B(n13548), .Z(n13531) );
  NAND U21822 ( .A(n13549), .B(n13550), .Z(n13548) );
  NANDN U21823 ( .A(n13551), .B(n13552), .Z(n13550) );
  NANDN U21824 ( .A(n13552), .B(n13551), .Z(n13547) );
  XOR U21825 ( .A(n13544), .B(n13553), .Z(N64182) );
  XNOR U21826 ( .A(n13542), .B(n13546), .Z(n13553) );
  XOR U21827 ( .A(n13539), .B(n13554), .Z(n13546) );
  XNOR U21828 ( .A(n13536), .B(n13538), .Z(n13554) );
  AND U21829 ( .A(n13555), .B(n13556), .Z(n13538) );
  NANDN U21830 ( .A(n13557), .B(n13558), .Z(n13556) );
  OR U21831 ( .A(n13559), .B(n13560), .Z(n13558) );
  IV U21832 ( .A(n13561), .Z(n13560) );
  NANDN U21833 ( .A(n13561), .B(n13559), .Z(n13555) );
  AND U21834 ( .A(n13562), .B(n13563), .Z(n13536) );
  NAND U21835 ( .A(n13564), .B(n13565), .Z(n13563) );
  NANDN U21836 ( .A(n13566), .B(n13567), .Z(n13565) );
  NANDN U21837 ( .A(n13567), .B(n13566), .Z(n13562) );
  IV U21838 ( .A(n13568), .Z(n13567) );
  NAND U21839 ( .A(n13569), .B(n13570), .Z(n13539) );
  NANDN U21840 ( .A(n13571), .B(n13572), .Z(n13570) );
  NANDN U21841 ( .A(n13573), .B(n13574), .Z(n13572) );
  NANDN U21842 ( .A(n13574), .B(n13573), .Z(n13569) );
  IV U21843 ( .A(n13575), .Z(n13573) );
  AND U21844 ( .A(n13576), .B(n13577), .Z(n13542) );
  NAND U21845 ( .A(n13578), .B(n13579), .Z(n13577) );
  NANDN U21846 ( .A(n13580), .B(n13581), .Z(n13579) );
  NANDN U21847 ( .A(n13581), .B(n13580), .Z(n13576) );
  XOR U21848 ( .A(n13552), .B(n13582), .Z(n13544) );
  XNOR U21849 ( .A(n13549), .B(n13551), .Z(n13582) );
  AND U21850 ( .A(n13583), .B(n13584), .Z(n13551) );
  NANDN U21851 ( .A(n13585), .B(n13586), .Z(n13584) );
  OR U21852 ( .A(n13587), .B(n13588), .Z(n13586) );
  IV U21853 ( .A(n13589), .Z(n13588) );
  NANDN U21854 ( .A(n13589), .B(n13587), .Z(n13583) );
  AND U21855 ( .A(n13590), .B(n13591), .Z(n13549) );
  NAND U21856 ( .A(n13592), .B(n13593), .Z(n13591) );
  NANDN U21857 ( .A(n13594), .B(n13595), .Z(n13593) );
  NANDN U21858 ( .A(n13595), .B(n13594), .Z(n13590) );
  IV U21859 ( .A(n13596), .Z(n13595) );
  NAND U21860 ( .A(n13597), .B(n13598), .Z(n13552) );
  NANDN U21861 ( .A(n13599), .B(n13600), .Z(n13598) );
  NANDN U21862 ( .A(n13601), .B(n13602), .Z(n13600) );
  NANDN U21863 ( .A(n13602), .B(n13601), .Z(n13597) );
  IV U21864 ( .A(n13603), .Z(n13601) );
  XOR U21865 ( .A(n13578), .B(n13604), .Z(N64181) );
  XNOR U21866 ( .A(n13581), .B(n13580), .Z(n13604) );
  XNOR U21867 ( .A(n13592), .B(n13605), .Z(n13580) );
  XNOR U21868 ( .A(n13596), .B(n13594), .Z(n13605) );
  XOR U21869 ( .A(n13602), .B(n13606), .Z(n13594) );
  XNOR U21870 ( .A(n13599), .B(n13603), .Z(n13606) );
  AND U21871 ( .A(n13607), .B(n13608), .Z(n13603) );
  NAND U21872 ( .A(n13609), .B(n13610), .Z(n13608) );
  NAND U21873 ( .A(n13611), .B(n13612), .Z(n13607) );
  AND U21874 ( .A(n13613), .B(n13614), .Z(n13599) );
  NAND U21875 ( .A(n13615), .B(n13616), .Z(n13614) );
  NAND U21876 ( .A(n13617), .B(n13618), .Z(n13613) );
  NANDN U21877 ( .A(n13619), .B(n13620), .Z(n13602) );
  ANDN U21878 ( .B(n13621), .A(n13622), .Z(n13596) );
  XNOR U21879 ( .A(n13587), .B(n13623), .Z(n13592) );
  XNOR U21880 ( .A(n13585), .B(n13589), .Z(n13623) );
  AND U21881 ( .A(n13624), .B(n13625), .Z(n13589) );
  NAND U21882 ( .A(n13626), .B(n13627), .Z(n13625) );
  NAND U21883 ( .A(n13628), .B(n13629), .Z(n13624) );
  AND U21884 ( .A(n13630), .B(n13631), .Z(n13585) );
  NAND U21885 ( .A(n13632), .B(n13633), .Z(n13631) );
  NAND U21886 ( .A(n13634), .B(n13635), .Z(n13630) );
  AND U21887 ( .A(n13636), .B(n13637), .Z(n13587) );
  NAND U21888 ( .A(n13638), .B(n13639), .Z(n13581) );
  XNOR U21889 ( .A(n13564), .B(n13640), .Z(n13578) );
  XNOR U21890 ( .A(n13568), .B(n13566), .Z(n13640) );
  XOR U21891 ( .A(n13574), .B(n13641), .Z(n13566) );
  XNOR U21892 ( .A(n13571), .B(n13575), .Z(n13641) );
  AND U21893 ( .A(n13642), .B(n13643), .Z(n13575) );
  NAND U21894 ( .A(n13644), .B(n13645), .Z(n13643) );
  NAND U21895 ( .A(n13646), .B(n13647), .Z(n13642) );
  AND U21896 ( .A(n13648), .B(n13649), .Z(n13571) );
  NAND U21897 ( .A(n13650), .B(n13651), .Z(n13649) );
  NAND U21898 ( .A(n13652), .B(n13653), .Z(n13648) );
  NANDN U21899 ( .A(n13654), .B(n13655), .Z(n13574) );
  ANDN U21900 ( .B(n13656), .A(n13657), .Z(n13568) );
  XNOR U21901 ( .A(n13559), .B(n13658), .Z(n13564) );
  XNOR U21902 ( .A(n13557), .B(n13561), .Z(n13658) );
  AND U21903 ( .A(n13659), .B(n13660), .Z(n13561) );
  NAND U21904 ( .A(n13661), .B(n13662), .Z(n13660) );
  NAND U21905 ( .A(n13663), .B(n13664), .Z(n13659) );
  AND U21906 ( .A(n13665), .B(n13666), .Z(n13557) );
  NAND U21907 ( .A(n13667), .B(n13668), .Z(n13666) );
  NAND U21908 ( .A(n13669), .B(n13670), .Z(n13665) );
  AND U21909 ( .A(n13671), .B(n13672), .Z(n13559) );
  XOR U21910 ( .A(n13639), .B(n13638), .Z(N64180) );
  XNOR U21911 ( .A(n13656), .B(n13657), .Z(n13638) );
  XNOR U21912 ( .A(n13671), .B(n13672), .Z(n13657) );
  XOR U21913 ( .A(n13668), .B(n13667), .Z(n13672) );
  XOR U21914 ( .A(y[6636]), .B(x[6636]), .Z(n13667) );
  XOR U21915 ( .A(n13670), .B(n13669), .Z(n13668) );
  XOR U21916 ( .A(y[6638]), .B(x[6638]), .Z(n13669) );
  XOR U21917 ( .A(y[6637]), .B(x[6637]), .Z(n13670) );
  XOR U21918 ( .A(n13662), .B(n13661), .Z(n13671) );
  XOR U21919 ( .A(n13664), .B(n13663), .Z(n13661) );
  XOR U21920 ( .A(y[6635]), .B(x[6635]), .Z(n13663) );
  XOR U21921 ( .A(y[6634]), .B(x[6634]), .Z(n13664) );
  XOR U21922 ( .A(y[6633]), .B(x[6633]), .Z(n13662) );
  XNOR U21923 ( .A(n13655), .B(n13654), .Z(n13656) );
  XNOR U21924 ( .A(n13651), .B(n13650), .Z(n13654) );
  XOR U21925 ( .A(n13653), .B(n13652), .Z(n13650) );
  XOR U21926 ( .A(y[6632]), .B(x[6632]), .Z(n13652) );
  XOR U21927 ( .A(y[6631]), .B(x[6631]), .Z(n13653) );
  XOR U21928 ( .A(y[6630]), .B(x[6630]), .Z(n13651) );
  XOR U21929 ( .A(n13645), .B(n13644), .Z(n13655) );
  XOR U21930 ( .A(n13647), .B(n13646), .Z(n13644) );
  XOR U21931 ( .A(y[6629]), .B(x[6629]), .Z(n13646) );
  XOR U21932 ( .A(y[6628]), .B(x[6628]), .Z(n13647) );
  XOR U21933 ( .A(y[6627]), .B(x[6627]), .Z(n13645) );
  XNOR U21934 ( .A(n13621), .B(n13622), .Z(n13639) );
  XNOR U21935 ( .A(n13636), .B(n13637), .Z(n13622) );
  XOR U21936 ( .A(n13633), .B(n13632), .Z(n13637) );
  XOR U21937 ( .A(y[6624]), .B(x[6624]), .Z(n13632) );
  XOR U21938 ( .A(n13635), .B(n13634), .Z(n13633) );
  XOR U21939 ( .A(y[6626]), .B(x[6626]), .Z(n13634) );
  XOR U21940 ( .A(y[6625]), .B(x[6625]), .Z(n13635) );
  XOR U21941 ( .A(n13627), .B(n13626), .Z(n13636) );
  XOR U21942 ( .A(n13629), .B(n13628), .Z(n13626) );
  XOR U21943 ( .A(y[6623]), .B(x[6623]), .Z(n13628) );
  XOR U21944 ( .A(y[6622]), .B(x[6622]), .Z(n13629) );
  XOR U21945 ( .A(y[6621]), .B(x[6621]), .Z(n13627) );
  XNOR U21946 ( .A(n13620), .B(n13619), .Z(n13621) );
  XNOR U21947 ( .A(n13616), .B(n13615), .Z(n13619) );
  XOR U21948 ( .A(n13618), .B(n13617), .Z(n13615) );
  XOR U21949 ( .A(y[6620]), .B(x[6620]), .Z(n13617) );
  XOR U21950 ( .A(y[6619]), .B(x[6619]), .Z(n13618) );
  XOR U21951 ( .A(y[6618]), .B(x[6618]), .Z(n13616) );
  XOR U21952 ( .A(n13610), .B(n13609), .Z(n13620) );
  XOR U21953 ( .A(n13612), .B(n13611), .Z(n13609) );
  XOR U21954 ( .A(y[6617]), .B(x[6617]), .Z(n13611) );
  XOR U21955 ( .A(y[6616]), .B(x[6616]), .Z(n13612) );
  XOR U21956 ( .A(y[6615]), .B(x[6615]), .Z(n13610) );
  NAND U21957 ( .A(n13673), .B(n13674), .Z(N64171) );
  NAND U21958 ( .A(n13675), .B(n13676), .Z(n13674) );
  NANDN U21959 ( .A(n13677), .B(n13678), .Z(n13676) );
  NANDN U21960 ( .A(n13678), .B(n13677), .Z(n13673) );
  XOR U21961 ( .A(n13677), .B(n13679), .Z(N64170) );
  XNOR U21962 ( .A(n13675), .B(n13678), .Z(n13679) );
  NAND U21963 ( .A(n13680), .B(n13681), .Z(n13678) );
  NAND U21964 ( .A(n13682), .B(n13683), .Z(n13681) );
  NANDN U21965 ( .A(n13684), .B(n13685), .Z(n13683) );
  NANDN U21966 ( .A(n13685), .B(n13684), .Z(n13680) );
  AND U21967 ( .A(n13686), .B(n13687), .Z(n13675) );
  NAND U21968 ( .A(n13688), .B(n13689), .Z(n13687) );
  NANDN U21969 ( .A(n13690), .B(n13691), .Z(n13689) );
  NANDN U21970 ( .A(n13691), .B(n13690), .Z(n13686) );
  IV U21971 ( .A(n13692), .Z(n13691) );
  AND U21972 ( .A(n13693), .B(n13694), .Z(n13677) );
  NAND U21973 ( .A(n13695), .B(n13696), .Z(n13694) );
  NANDN U21974 ( .A(n13697), .B(n13698), .Z(n13696) );
  NANDN U21975 ( .A(n13698), .B(n13697), .Z(n13693) );
  XOR U21976 ( .A(n13690), .B(n13699), .Z(N64169) );
  XNOR U21977 ( .A(n13688), .B(n13692), .Z(n13699) );
  XOR U21978 ( .A(n13685), .B(n13700), .Z(n13692) );
  XNOR U21979 ( .A(n13682), .B(n13684), .Z(n13700) );
  AND U21980 ( .A(n13701), .B(n13702), .Z(n13684) );
  NANDN U21981 ( .A(n13703), .B(n13704), .Z(n13702) );
  OR U21982 ( .A(n13705), .B(n13706), .Z(n13704) );
  IV U21983 ( .A(n13707), .Z(n13706) );
  NANDN U21984 ( .A(n13707), .B(n13705), .Z(n13701) );
  AND U21985 ( .A(n13708), .B(n13709), .Z(n13682) );
  NAND U21986 ( .A(n13710), .B(n13711), .Z(n13709) );
  NANDN U21987 ( .A(n13712), .B(n13713), .Z(n13711) );
  NANDN U21988 ( .A(n13713), .B(n13712), .Z(n13708) );
  IV U21989 ( .A(n13714), .Z(n13713) );
  NAND U21990 ( .A(n13715), .B(n13716), .Z(n13685) );
  NANDN U21991 ( .A(n13717), .B(n13718), .Z(n13716) );
  NANDN U21992 ( .A(n13719), .B(n13720), .Z(n13718) );
  NANDN U21993 ( .A(n13720), .B(n13719), .Z(n13715) );
  IV U21994 ( .A(n13721), .Z(n13719) );
  AND U21995 ( .A(n13722), .B(n13723), .Z(n13688) );
  NAND U21996 ( .A(n13724), .B(n13725), .Z(n13723) );
  NANDN U21997 ( .A(n13726), .B(n13727), .Z(n13725) );
  NANDN U21998 ( .A(n13727), .B(n13726), .Z(n13722) );
  XOR U21999 ( .A(n13698), .B(n13728), .Z(n13690) );
  XNOR U22000 ( .A(n13695), .B(n13697), .Z(n13728) );
  AND U22001 ( .A(n13729), .B(n13730), .Z(n13697) );
  NANDN U22002 ( .A(n13731), .B(n13732), .Z(n13730) );
  OR U22003 ( .A(n13733), .B(n13734), .Z(n13732) );
  IV U22004 ( .A(n13735), .Z(n13734) );
  NANDN U22005 ( .A(n13735), .B(n13733), .Z(n13729) );
  AND U22006 ( .A(n13736), .B(n13737), .Z(n13695) );
  NAND U22007 ( .A(n13738), .B(n13739), .Z(n13737) );
  NANDN U22008 ( .A(n13740), .B(n13741), .Z(n13739) );
  NANDN U22009 ( .A(n13741), .B(n13740), .Z(n13736) );
  IV U22010 ( .A(n13742), .Z(n13741) );
  NAND U22011 ( .A(n13743), .B(n13744), .Z(n13698) );
  NANDN U22012 ( .A(n13745), .B(n13746), .Z(n13744) );
  NANDN U22013 ( .A(n13747), .B(n13748), .Z(n13746) );
  NANDN U22014 ( .A(n13748), .B(n13747), .Z(n13743) );
  IV U22015 ( .A(n13749), .Z(n13747) );
  XOR U22016 ( .A(n13724), .B(n13750), .Z(N64168) );
  XNOR U22017 ( .A(n13727), .B(n13726), .Z(n13750) );
  XNOR U22018 ( .A(n13738), .B(n13751), .Z(n13726) );
  XNOR U22019 ( .A(n13742), .B(n13740), .Z(n13751) );
  XOR U22020 ( .A(n13748), .B(n13752), .Z(n13740) );
  XNOR U22021 ( .A(n13745), .B(n13749), .Z(n13752) );
  AND U22022 ( .A(n13753), .B(n13754), .Z(n13749) );
  NAND U22023 ( .A(n13755), .B(n13756), .Z(n13754) );
  NAND U22024 ( .A(n13757), .B(n13758), .Z(n13753) );
  AND U22025 ( .A(n13759), .B(n13760), .Z(n13745) );
  NAND U22026 ( .A(n13761), .B(n13762), .Z(n13760) );
  NAND U22027 ( .A(n13763), .B(n13764), .Z(n13759) );
  NANDN U22028 ( .A(n13765), .B(n13766), .Z(n13748) );
  ANDN U22029 ( .B(n13767), .A(n13768), .Z(n13742) );
  XNOR U22030 ( .A(n13733), .B(n13769), .Z(n13738) );
  XNOR U22031 ( .A(n13731), .B(n13735), .Z(n13769) );
  AND U22032 ( .A(n13770), .B(n13771), .Z(n13735) );
  NAND U22033 ( .A(n13772), .B(n13773), .Z(n13771) );
  NAND U22034 ( .A(n13774), .B(n13775), .Z(n13770) );
  AND U22035 ( .A(n13776), .B(n13777), .Z(n13731) );
  NAND U22036 ( .A(n13778), .B(n13779), .Z(n13777) );
  NAND U22037 ( .A(n13780), .B(n13781), .Z(n13776) );
  AND U22038 ( .A(n13782), .B(n13783), .Z(n13733) );
  NAND U22039 ( .A(n13784), .B(n13785), .Z(n13727) );
  XNOR U22040 ( .A(n13710), .B(n13786), .Z(n13724) );
  XNOR U22041 ( .A(n13714), .B(n13712), .Z(n13786) );
  XOR U22042 ( .A(n13720), .B(n13787), .Z(n13712) );
  XNOR U22043 ( .A(n13717), .B(n13721), .Z(n13787) );
  AND U22044 ( .A(n13788), .B(n13789), .Z(n13721) );
  NAND U22045 ( .A(n13790), .B(n13791), .Z(n13789) );
  NAND U22046 ( .A(n13792), .B(n13793), .Z(n13788) );
  AND U22047 ( .A(n13794), .B(n13795), .Z(n13717) );
  NAND U22048 ( .A(n13796), .B(n13797), .Z(n13795) );
  NAND U22049 ( .A(n13798), .B(n13799), .Z(n13794) );
  NANDN U22050 ( .A(n13800), .B(n13801), .Z(n13720) );
  ANDN U22051 ( .B(n13802), .A(n13803), .Z(n13714) );
  XNOR U22052 ( .A(n13705), .B(n13804), .Z(n13710) );
  XNOR U22053 ( .A(n13703), .B(n13707), .Z(n13804) );
  AND U22054 ( .A(n13805), .B(n13806), .Z(n13707) );
  NAND U22055 ( .A(n13807), .B(n13808), .Z(n13806) );
  NAND U22056 ( .A(n13809), .B(n13810), .Z(n13805) );
  AND U22057 ( .A(n13811), .B(n13812), .Z(n13703) );
  NAND U22058 ( .A(n13813), .B(n13814), .Z(n13812) );
  NAND U22059 ( .A(n13815), .B(n13816), .Z(n13811) );
  AND U22060 ( .A(n13817), .B(n13818), .Z(n13705) );
  XOR U22061 ( .A(n13785), .B(n13784), .Z(N64167) );
  XNOR U22062 ( .A(n13802), .B(n13803), .Z(n13784) );
  XNOR U22063 ( .A(n13817), .B(n13818), .Z(n13803) );
  XOR U22064 ( .A(n13814), .B(n13813), .Z(n13818) );
  XOR U22065 ( .A(y[6612]), .B(x[6612]), .Z(n13813) );
  XOR U22066 ( .A(n13816), .B(n13815), .Z(n13814) );
  XOR U22067 ( .A(y[6614]), .B(x[6614]), .Z(n13815) );
  XOR U22068 ( .A(y[6613]), .B(x[6613]), .Z(n13816) );
  XOR U22069 ( .A(n13808), .B(n13807), .Z(n13817) );
  XOR U22070 ( .A(n13810), .B(n13809), .Z(n13807) );
  XOR U22071 ( .A(y[6611]), .B(x[6611]), .Z(n13809) );
  XOR U22072 ( .A(y[6610]), .B(x[6610]), .Z(n13810) );
  XOR U22073 ( .A(y[6609]), .B(x[6609]), .Z(n13808) );
  XNOR U22074 ( .A(n13801), .B(n13800), .Z(n13802) );
  XNOR U22075 ( .A(n13797), .B(n13796), .Z(n13800) );
  XOR U22076 ( .A(n13799), .B(n13798), .Z(n13796) );
  XOR U22077 ( .A(y[6608]), .B(x[6608]), .Z(n13798) );
  XOR U22078 ( .A(y[6607]), .B(x[6607]), .Z(n13799) );
  XOR U22079 ( .A(y[6606]), .B(x[6606]), .Z(n13797) );
  XOR U22080 ( .A(n13791), .B(n13790), .Z(n13801) );
  XOR U22081 ( .A(n13793), .B(n13792), .Z(n13790) );
  XOR U22082 ( .A(y[6605]), .B(x[6605]), .Z(n13792) );
  XOR U22083 ( .A(y[6604]), .B(x[6604]), .Z(n13793) );
  XOR U22084 ( .A(y[6603]), .B(x[6603]), .Z(n13791) );
  XNOR U22085 ( .A(n13767), .B(n13768), .Z(n13785) );
  XNOR U22086 ( .A(n13782), .B(n13783), .Z(n13768) );
  XOR U22087 ( .A(n13779), .B(n13778), .Z(n13783) );
  XOR U22088 ( .A(y[6600]), .B(x[6600]), .Z(n13778) );
  XOR U22089 ( .A(n13781), .B(n13780), .Z(n13779) );
  XOR U22090 ( .A(y[6602]), .B(x[6602]), .Z(n13780) );
  XOR U22091 ( .A(y[6601]), .B(x[6601]), .Z(n13781) );
  XOR U22092 ( .A(n13773), .B(n13772), .Z(n13782) );
  XOR U22093 ( .A(n13775), .B(n13774), .Z(n13772) );
  XOR U22094 ( .A(y[6599]), .B(x[6599]), .Z(n13774) );
  XOR U22095 ( .A(y[6598]), .B(x[6598]), .Z(n13775) );
  XOR U22096 ( .A(y[6597]), .B(x[6597]), .Z(n13773) );
  XNOR U22097 ( .A(n13766), .B(n13765), .Z(n13767) );
  XNOR U22098 ( .A(n13762), .B(n13761), .Z(n13765) );
  XOR U22099 ( .A(n13764), .B(n13763), .Z(n13761) );
  XOR U22100 ( .A(y[6596]), .B(x[6596]), .Z(n13763) );
  XOR U22101 ( .A(y[6595]), .B(x[6595]), .Z(n13764) );
  XOR U22102 ( .A(y[6594]), .B(x[6594]), .Z(n13762) );
  XOR U22103 ( .A(n13756), .B(n13755), .Z(n13766) );
  XOR U22104 ( .A(n13758), .B(n13757), .Z(n13755) );
  XOR U22105 ( .A(y[6593]), .B(x[6593]), .Z(n13757) );
  XOR U22106 ( .A(y[6592]), .B(x[6592]), .Z(n13758) );
  XOR U22107 ( .A(y[6591]), .B(x[6591]), .Z(n13756) );
  NAND U22108 ( .A(n13819), .B(n13820), .Z(N64158) );
  NAND U22109 ( .A(n13821), .B(n13822), .Z(n13820) );
  NANDN U22110 ( .A(n13823), .B(n13824), .Z(n13822) );
  NANDN U22111 ( .A(n13824), .B(n13823), .Z(n13819) );
  XOR U22112 ( .A(n13823), .B(n13825), .Z(N64157) );
  XNOR U22113 ( .A(n13821), .B(n13824), .Z(n13825) );
  NAND U22114 ( .A(n13826), .B(n13827), .Z(n13824) );
  NAND U22115 ( .A(n13828), .B(n13829), .Z(n13827) );
  NANDN U22116 ( .A(n13830), .B(n13831), .Z(n13829) );
  NANDN U22117 ( .A(n13831), .B(n13830), .Z(n13826) );
  AND U22118 ( .A(n13832), .B(n13833), .Z(n13821) );
  NAND U22119 ( .A(n13834), .B(n13835), .Z(n13833) );
  NANDN U22120 ( .A(n13836), .B(n13837), .Z(n13835) );
  NANDN U22121 ( .A(n13837), .B(n13836), .Z(n13832) );
  IV U22122 ( .A(n13838), .Z(n13837) );
  AND U22123 ( .A(n13839), .B(n13840), .Z(n13823) );
  NAND U22124 ( .A(n13841), .B(n13842), .Z(n13840) );
  NANDN U22125 ( .A(n13843), .B(n13844), .Z(n13842) );
  NANDN U22126 ( .A(n13844), .B(n13843), .Z(n13839) );
  XOR U22127 ( .A(n13836), .B(n13845), .Z(N64156) );
  XNOR U22128 ( .A(n13834), .B(n13838), .Z(n13845) );
  XOR U22129 ( .A(n13831), .B(n13846), .Z(n13838) );
  XNOR U22130 ( .A(n13828), .B(n13830), .Z(n13846) );
  AND U22131 ( .A(n13847), .B(n13848), .Z(n13830) );
  NANDN U22132 ( .A(n13849), .B(n13850), .Z(n13848) );
  OR U22133 ( .A(n13851), .B(n13852), .Z(n13850) );
  IV U22134 ( .A(n13853), .Z(n13852) );
  NANDN U22135 ( .A(n13853), .B(n13851), .Z(n13847) );
  AND U22136 ( .A(n13854), .B(n13855), .Z(n13828) );
  NAND U22137 ( .A(n13856), .B(n13857), .Z(n13855) );
  NANDN U22138 ( .A(n13858), .B(n13859), .Z(n13857) );
  NANDN U22139 ( .A(n13859), .B(n13858), .Z(n13854) );
  IV U22140 ( .A(n13860), .Z(n13859) );
  NAND U22141 ( .A(n13861), .B(n13862), .Z(n13831) );
  NANDN U22142 ( .A(n13863), .B(n13864), .Z(n13862) );
  NANDN U22143 ( .A(n13865), .B(n13866), .Z(n13864) );
  NANDN U22144 ( .A(n13866), .B(n13865), .Z(n13861) );
  IV U22145 ( .A(n13867), .Z(n13865) );
  AND U22146 ( .A(n13868), .B(n13869), .Z(n13834) );
  NAND U22147 ( .A(n13870), .B(n13871), .Z(n13869) );
  NANDN U22148 ( .A(n13872), .B(n13873), .Z(n13871) );
  NANDN U22149 ( .A(n13873), .B(n13872), .Z(n13868) );
  XOR U22150 ( .A(n13844), .B(n13874), .Z(n13836) );
  XNOR U22151 ( .A(n13841), .B(n13843), .Z(n13874) );
  AND U22152 ( .A(n13875), .B(n13876), .Z(n13843) );
  NANDN U22153 ( .A(n13877), .B(n13878), .Z(n13876) );
  OR U22154 ( .A(n13879), .B(n13880), .Z(n13878) );
  IV U22155 ( .A(n13881), .Z(n13880) );
  NANDN U22156 ( .A(n13881), .B(n13879), .Z(n13875) );
  AND U22157 ( .A(n13882), .B(n13883), .Z(n13841) );
  NAND U22158 ( .A(n13884), .B(n13885), .Z(n13883) );
  NANDN U22159 ( .A(n13886), .B(n13887), .Z(n13885) );
  NANDN U22160 ( .A(n13887), .B(n13886), .Z(n13882) );
  IV U22161 ( .A(n13888), .Z(n13887) );
  NAND U22162 ( .A(n13889), .B(n13890), .Z(n13844) );
  NANDN U22163 ( .A(n13891), .B(n13892), .Z(n13890) );
  NANDN U22164 ( .A(n13893), .B(n13894), .Z(n13892) );
  NANDN U22165 ( .A(n13894), .B(n13893), .Z(n13889) );
  IV U22166 ( .A(n13895), .Z(n13893) );
  XOR U22167 ( .A(n13870), .B(n13896), .Z(N64155) );
  XNOR U22168 ( .A(n13873), .B(n13872), .Z(n13896) );
  XNOR U22169 ( .A(n13884), .B(n13897), .Z(n13872) );
  XNOR U22170 ( .A(n13888), .B(n13886), .Z(n13897) );
  XOR U22171 ( .A(n13894), .B(n13898), .Z(n13886) );
  XNOR U22172 ( .A(n13891), .B(n13895), .Z(n13898) );
  AND U22173 ( .A(n13899), .B(n13900), .Z(n13895) );
  NAND U22174 ( .A(n13901), .B(n13902), .Z(n13900) );
  NAND U22175 ( .A(n13903), .B(n13904), .Z(n13899) );
  AND U22176 ( .A(n13905), .B(n13906), .Z(n13891) );
  NAND U22177 ( .A(n13907), .B(n13908), .Z(n13906) );
  NAND U22178 ( .A(n13909), .B(n13910), .Z(n13905) );
  NANDN U22179 ( .A(n13911), .B(n13912), .Z(n13894) );
  ANDN U22180 ( .B(n13913), .A(n13914), .Z(n13888) );
  XNOR U22181 ( .A(n13879), .B(n13915), .Z(n13884) );
  XNOR U22182 ( .A(n13877), .B(n13881), .Z(n13915) );
  AND U22183 ( .A(n13916), .B(n13917), .Z(n13881) );
  NAND U22184 ( .A(n13918), .B(n13919), .Z(n13917) );
  NAND U22185 ( .A(n13920), .B(n13921), .Z(n13916) );
  AND U22186 ( .A(n13922), .B(n13923), .Z(n13877) );
  NAND U22187 ( .A(n13924), .B(n13925), .Z(n13923) );
  NAND U22188 ( .A(n13926), .B(n13927), .Z(n13922) );
  AND U22189 ( .A(n13928), .B(n13929), .Z(n13879) );
  NAND U22190 ( .A(n13930), .B(n13931), .Z(n13873) );
  XNOR U22191 ( .A(n13856), .B(n13932), .Z(n13870) );
  XNOR U22192 ( .A(n13860), .B(n13858), .Z(n13932) );
  XOR U22193 ( .A(n13866), .B(n13933), .Z(n13858) );
  XNOR U22194 ( .A(n13863), .B(n13867), .Z(n13933) );
  AND U22195 ( .A(n13934), .B(n13935), .Z(n13867) );
  NAND U22196 ( .A(n13936), .B(n13937), .Z(n13935) );
  NAND U22197 ( .A(n13938), .B(n13939), .Z(n13934) );
  AND U22198 ( .A(n13940), .B(n13941), .Z(n13863) );
  NAND U22199 ( .A(n13942), .B(n13943), .Z(n13941) );
  NAND U22200 ( .A(n13944), .B(n13945), .Z(n13940) );
  NANDN U22201 ( .A(n13946), .B(n13947), .Z(n13866) );
  ANDN U22202 ( .B(n13948), .A(n13949), .Z(n13860) );
  XNOR U22203 ( .A(n13851), .B(n13950), .Z(n13856) );
  XNOR U22204 ( .A(n13849), .B(n13853), .Z(n13950) );
  AND U22205 ( .A(n13951), .B(n13952), .Z(n13853) );
  NAND U22206 ( .A(n13953), .B(n13954), .Z(n13952) );
  NAND U22207 ( .A(n13955), .B(n13956), .Z(n13951) );
  AND U22208 ( .A(n13957), .B(n13958), .Z(n13849) );
  NAND U22209 ( .A(n13959), .B(n13960), .Z(n13958) );
  NAND U22210 ( .A(n13961), .B(n13962), .Z(n13957) );
  AND U22211 ( .A(n13963), .B(n13964), .Z(n13851) );
  XOR U22212 ( .A(n13931), .B(n13930), .Z(N64154) );
  XNOR U22213 ( .A(n13948), .B(n13949), .Z(n13930) );
  XNOR U22214 ( .A(n13963), .B(n13964), .Z(n13949) );
  XOR U22215 ( .A(n13960), .B(n13959), .Z(n13964) );
  XOR U22216 ( .A(y[6588]), .B(x[6588]), .Z(n13959) );
  XOR U22217 ( .A(n13962), .B(n13961), .Z(n13960) );
  XOR U22218 ( .A(y[6590]), .B(x[6590]), .Z(n13961) );
  XOR U22219 ( .A(y[6589]), .B(x[6589]), .Z(n13962) );
  XOR U22220 ( .A(n13954), .B(n13953), .Z(n13963) );
  XOR U22221 ( .A(n13956), .B(n13955), .Z(n13953) );
  XOR U22222 ( .A(y[6587]), .B(x[6587]), .Z(n13955) );
  XOR U22223 ( .A(y[6586]), .B(x[6586]), .Z(n13956) );
  XOR U22224 ( .A(y[6585]), .B(x[6585]), .Z(n13954) );
  XNOR U22225 ( .A(n13947), .B(n13946), .Z(n13948) );
  XNOR U22226 ( .A(n13943), .B(n13942), .Z(n13946) );
  XOR U22227 ( .A(n13945), .B(n13944), .Z(n13942) );
  XOR U22228 ( .A(y[6584]), .B(x[6584]), .Z(n13944) );
  XOR U22229 ( .A(y[6583]), .B(x[6583]), .Z(n13945) );
  XOR U22230 ( .A(y[6582]), .B(x[6582]), .Z(n13943) );
  XOR U22231 ( .A(n13937), .B(n13936), .Z(n13947) );
  XOR U22232 ( .A(n13939), .B(n13938), .Z(n13936) );
  XOR U22233 ( .A(y[6581]), .B(x[6581]), .Z(n13938) );
  XOR U22234 ( .A(y[6580]), .B(x[6580]), .Z(n13939) );
  XOR U22235 ( .A(y[6579]), .B(x[6579]), .Z(n13937) );
  XNOR U22236 ( .A(n13913), .B(n13914), .Z(n13931) );
  XNOR U22237 ( .A(n13928), .B(n13929), .Z(n13914) );
  XOR U22238 ( .A(n13925), .B(n13924), .Z(n13929) );
  XOR U22239 ( .A(y[6576]), .B(x[6576]), .Z(n13924) );
  XOR U22240 ( .A(n13927), .B(n13926), .Z(n13925) );
  XOR U22241 ( .A(y[6578]), .B(x[6578]), .Z(n13926) );
  XOR U22242 ( .A(y[6577]), .B(x[6577]), .Z(n13927) );
  XOR U22243 ( .A(n13919), .B(n13918), .Z(n13928) );
  XOR U22244 ( .A(n13921), .B(n13920), .Z(n13918) );
  XOR U22245 ( .A(y[6575]), .B(x[6575]), .Z(n13920) );
  XOR U22246 ( .A(y[6574]), .B(x[6574]), .Z(n13921) );
  XOR U22247 ( .A(y[6573]), .B(x[6573]), .Z(n13919) );
  XNOR U22248 ( .A(n13912), .B(n13911), .Z(n13913) );
  XNOR U22249 ( .A(n13908), .B(n13907), .Z(n13911) );
  XOR U22250 ( .A(n13910), .B(n13909), .Z(n13907) );
  XOR U22251 ( .A(y[6572]), .B(x[6572]), .Z(n13909) );
  XOR U22252 ( .A(y[6571]), .B(x[6571]), .Z(n13910) );
  XOR U22253 ( .A(y[6570]), .B(x[6570]), .Z(n13908) );
  XOR U22254 ( .A(n13902), .B(n13901), .Z(n13912) );
  XOR U22255 ( .A(n13904), .B(n13903), .Z(n13901) );
  XOR U22256 ( .A(y[6569]), .B(x[6569]), .Z(n13903) );
  XOR U22257 ( .A(y[6568]), .B(x[6568]), .Z(n13904) );
  XOR U22258 ( .A(y[6567]), .B(x[6567]), .Z(n13902) );
  NAND U22259 ( .A(n13965), .B(n13966), .Z(N64145) );
  NAND U22260 ( .A(n13967), .B(n13968), .Z(n13966) );
  NANDN U22261 ( .A(n13969), .B(n13970), .Z(n13968) );
  NANDN U22262 ( .A(n13970), .B(n13969), .Z(n13965) );
  XOR U22263 ( .A(n13969), .B(n13971), .Z(N64144) );
  XNOR U22264 ( .A(n13967), .B(n13970), .Z(n13971) );
  NAND U22265 ( .A(n13972), .B(n13973), .Z(n13970) );
  NAND U22266 ( .A(n13974), .B(n13975), .Z(n13973) );
  NANDN U22267 ( .A(n13976), .B(n13977), .Z(n13975) );
  NANDN U22268 ( .A(n13977), .B(n13976), .Z(n13972) );
  AND U22269 ( .A(n13978), .B(n13979), .Z(n13967) );
  NAND U22270 ( .A(n13980), .B(n13981), .Z(n13979) );
  NANDN U22271 ( .A(n13982), .B(n13983), .Z(n13981) );
  NANDN U22272 ( .A(n13983), .B(n13982), .Z(n13978) );
  IV U22273 ( .A(n13984), .Z(n13983) );
  AND U22274 ( .A(n13985), .B(n13986), .Z(n13969) );
  NAND U22275 ( .A(n13987), .B(n13988), .Z(n13986) );
  NANDN U22276 ( .A(n13989), .B(n13990), .Z(n13988) );
  NANDN U22277 ( .A(n13990), .B(n13989), .Z(n13985) );
  XOR U22278 ( .A(n13982), .B(n13991), .Z(N64143) );
  XNOR U22279 ( .A(n13980), .B(n13984), .Z(n13991) );
  XOR U22280 ( .A(n13977), .B(n13992), .Z(n13984) );
  XNOR U22281 ( .A(n13974), .B(n13976), .Z(n13992) );
  AND U22282 ( .A(n13993), .B(n13994), .Z(n13976) );
  NANDN U22283 ( .A(n13995), .B(n13996), .Z(n13994) );
  OR U22284 ( .A(n13997), .B(n13998), .Z(n13996) );
  IV U22285 ( .A(n13999), .Z(n13998) );
  NANDN U22286 ( .A(n13999), .B(n13997), .Z(n13993) );
  AND U22287 ( .A(n14000), .B(n14001), .Z(n13974) );
  NAND U22288 ( .A(n14002), .B(n14003), .Z(n14001) );
  NANDN U22289 ( .A(n14004), .B(n14005), .Z(n14003) );
  NANDN U22290 ( .A(n14005), .B(n14004), .Z(n14000) );
  IV U22291 ( .A(n14006), .Z(n14005) );
  NAND U22292 ( .A(n14007), .B(n14008), .Z(n13977) );
  NANDN U22293 ( .A(n14009), .B(n14010), .Z(n14008) );
  NANDN U22294 ( .A(n14011), .B(n14012), .Z(n14010) );
  NANDN U22295 ( .A(n14012), .B(n14011), .Z(n14007) );
  IV U22296 ( .A(n14013), .Z(n14011) );
  AND U22297 ( .A(n14014), .B(n14015), .Z(n13980) );
  NAND U22298 ( .A(n14016), .B(n14017), .Z(n14015) );
  NANDN U22299 ( .A(n14018), .B(n14019), .Z(n14017) );
  NANDN U22300 ( .A(n14019), .B(n14018), .Z(n14014) );
  XOR U22301 ( .A(n13990), .B(n14020), .Z(n13982) );
  XNOR U22302 ( .A(n13987), .B(n13989), .Z(n14020) );
  AND U22303 ( .A(n14021), .B(n14022), .Z(n13989) );
  NANDN U22304 ( .A(n14023), .B(n14024), .Z(n14022) );
  OR U22305 ( .A(n14025), .B(n14026), .Z(n14024) );
  IV U22306 ( .A(n14027), .Z(n14026) );
  NANDN U22307 ( .A(n14027), .B(n14025), .Z(n14021) );
  AND U22308 ( .A(n14028), .B(n14029), .Z(n13987) );
  NAND U22309 ( .A(n14030), .B(n14031), .Z(n14029) );
  NANDN U22310 ( .A(n14032), .B(n14033), .Z(n14031) );
  NANDN U22311 ( .A(n14033), .B(n14032), .Z(n14028) );
  IV U22312 ( .A(n14034), .Z(n14033) );
  NAND U22313 ( .A(n14035), .B(n14036), .Z(n13990) );
  NANDN U22314 ( .A(n14037), .B(n14038), .Z(n14036) );
  NANDN U22315 ( .A(n14039), .B(n14040), .Z(n14038) );
  NANDN U22316 ( .A(n14040), .B(n14039), .Z(n14035) );
  IV U22317 ( .A(n14041), .Z(n14039) );
  XOR U22318 ( .A(n14016), .B(n14042), .Z(N64142) );
  XNOR U22319 ( .A(n14019), .B(n14018), .Z(n14042) );
  XNOR U22320 ( .A(n14030), .B(n14043), .Z(n14018) );
  XNOR U22321 ( .A(n14034), .B(n14032), .Z(n14043) );
  XOR U22322 ( .A(n14040), .B(n14044), .Z(n14032) );
  XNOR U22323 ( .A(n14037), .B(n14041), .Z(n14044) );
  AND U22324 ( .A(n14045), .B(n14046), .Z(n14041) );
  NAND U22325 ( .A(n14047), .B(n14048), .Z(n14046) );
  NAND U22326 ( .A(n14049), .B(n14050), .Z(n14045) );
  AND U22327 ( .A(n14051), .B(n14052), .Z(n14037) );
  NAND U22328 ( .A(n14053), .B(n14054), .Z(n14052) );
  NAND U22329 ( .A(n14055), .B(n14056), .Z(n14051) );
  NANDN U22330 ( .A(n14057), .B(n14058), .Z(n14040) );
  ANDN U22331 ( .B(n14059), .A(n14060), .Z(n14034) );
  XNOR U22332 ( .A(n14025), .B(n14061), .Z(n14030) );
  XNOR U22333 ( .A(n14023), .B(n14027), .Z(n14061) );
  AND U22334 ( .A(n14062), .B(n14063), .Z(n14027) );
  NAND U22335 ( .A(n14064), .B(n14065), .Z(n14063) );
  NAND U22336 ( .A(n14066), .B(n14067), .Z(n14062) );
  AND U22337 ( .A(n14068), .B(n14069), .Z(n14023) );
  NAND U22338 ( .A(n14070), .B(n14071), .Z(n14069) );
  NAND U22339 ( .A(n14072), .B(n14073), .Z(n14068) );
  AND U22340 ( .A(n14074), .B(n14075), .Z(n14025) );
  NAND U22341 ( .A(n14076), .B(n14077), .Z(n14019) );
  XNOR U22342 ( .A(n14002), .B(n14078), .Z(n14016) );
  XNOR U22343 ( .A(n14006), .B(n14004), .Z(n14078) );
  XOR U22344 ( .A(n14012), .B(n14079), .Z(n14004) );
  XNOR U22345 ( .A(n14009), .B(n14013), .Z(n14079) );
  AND U22346 ( .A(n14080), .B(n14081), .Z(n14013) );
  NAND U22347 ( .A(n14082), .B(n14083), .Z(n14081) );
  NAND U22348 ( .A(n14084), .B(n14085), .Z(n14080) );
  AND U22349 ( .A(n14086), .B(n14087), .Z(n14009) );
  NAND U22350 ( .A(n14088), .B(n14089), .Z(n14087) );
  NAND U22351 ( .A(n14090), .B(n14091), .Z(n14086) );
  NANDN U22352 ( .A(n14092), .B(n14093), .Z(n14012) );
  ANDN U22353 ( .B(n14094), .A(n14095), .Z(n14006) );
  XNOR U22354 ( .A(n13997), .B(n14096), .Z(n14002) );
  XNOR U22355 ( .A(n13995), .B(n13999), .Z(n14096) );
  AND U22356 ( .A(n14097), .B(n14098), .Z(n13999) );
  NAND U22357 ( .A(n14099), .B(n14100), .Z(n14098) );
  NAND U22358 ( .A(n14101), .B(n14102), .Z(n14097) );
  AND U22359 ( .A(n14103), .B(n14104), .Z(n13995) );
  NAND U22360 ( .A(n14105), .B(n14106), .Z(n14104) );
  NAND U22361 ( .A(n14107), .B(n14108), .Z(n14103) );
  AND U22362 ( .A(n14109), .B(n14110), .Z(n13997) );
  XOR U22363 ( .A(n14077), .B(n14076), .Z(N64141) );
  XNOR U22364 ( .A(n14094), .B(n14095), .Z(n14076) );
  XNOR U22365 ( .A(n14109), .B(n14110), .Z(n14095) );
  XOR U22366 ( .A(n14106), .B(n14105), .Z(n14110) );
  XOR U22367 ( .A(y[6564]), .B(x[6564]), .Z(n14105) );
  XOR U22368 ( .A(n14108), .B(n14107), .Z(n14106) );
  XOR U22369 ( .A(y[6566]), .B(x[6566]), .Z(n14107) );
  XOR U22370 ( .A(y[6565]), .B(x[6565]), .Z(n14108) );
  XOR U22371 ( .A(n14100), .B(n14099), .Z(n14109) );
  XOR U22372 ( .A(n14102), .B(n14101), .Z(n14099) );
  XOR U22373 ( .A(y[6563]), .B(x[6563]), .Z(n14101) );
  XOR U22374 ( .A(y[6562]), .B(x[6562]), .Z(n14102) );
  XOR U22375 ( .A(y[6561]), .B(x[6561]), .Z(n14100) );
  XNOR U22376 ( .A(n14093), .B(n14092), .Z(n14094) );
  XNOR U22377 ( .A(n14089), .B(n14088), .Z(n14092) );
  XOR U22378 ( .A(n14091), .B(n14090), .Z(n14088) );
  XOR U22379 ( .A(y[6560]), .B(x[6560]), .Z(n14090) );
  XOR U22380 ( .A(y[6559]), .B(x[6559]), .Z(n14091) );
  XOR U22381 ( .A(y[6558]), .B(x[6558]), .Z(n14089) );
  XOR U22382 ( .A(n14083), .B(n14082), .Z(n14093) );
  XOR U22383 ( .A(n14085), .B(n14084), .Z(n14082) );
  XOR U22384 ( .A(y[6557]), .B(x[6557]), .Z(n14084) );
  XOR U22385 ( .A(y[6556]), .B(x[6556]), .Z(n14085) );
  XOR U22386 ( .A(y[6555]), .B(x[6555]), .Z(n14083) );
  XNOR U22387 ( .A(n14059), .B(n14060), .Z(n14077) );
  XNOR U22388 ( .A(n14074), .B(n14075), .Z(n14060) );
  XOR U22389 ( .A(n14071), .B(n14070), .Z(n14075) );
  XOR U22390 ( .A(y[6552]), .B(x[6552]), .Z(n14070) );
  XOR U22391 ( .A(n14073), .B(n14072), .Z(n14071) );
  XOR U22392 ( .A(y[6554]), .B(x[6554]), .Z(n14072) );
  XOR U22393 ( .A(y[6553]), .B(x[6553]), .Z(n14073) );
  XOR U22394 ( .A(n14065), .B(n14064), .Z(n14074) );
  XOR U22395 ( .A(n14067), .B(n14066), .Z(n14064) );
  XOR U22396 ( .A(y[6551]), .B(x[6551]), .Z(n14066) );
  XOR U22397 ( .A(y[6550]), .B(x[6550]), .Z(n14067) );
  XOR U22398 ( .A(y[6549]), .B(x[6549]), .Z(n14065) );
  XNOR U22399 ( .A(n14058), .B(n14057), .Z(n14059) );
  XNOR U22400 ( .A(n14054), .B(n14053), .Z(n14057) );
  XOR U22401 ( .A(n14056), .B(n14055), .Z(n14053) );
  XOR U22402 ( .A(y[6548]), .B(x[6548]), .Z(n14055) );
  XOR U22403 ( .A(y[6547]), .B(x[6547]), .Z(n14056) );
  XOR U22404 ( .A(y[6546]), .B(x[6546]), .Z(n14054) );
  XOR U22405 ( .A(n14048), .B(n14047), .Z(n14058) );
  XOR U22406 ( .A(n14050), .B(n14049), .Z(n14047) );
  XOR U22407 ( .A(y[6545]), .B(x[6545]), .Z(n14049) );
  XOR U22408 ( .A(y[6544]), .B(x[6544]), .Z(n14050) );
  XOR U22409 ( .A(y[6543]), .B(x[6543]), .Z(n14048) );
  NAND U22410 ( .A(n14111), .B(n14112), .Z(N64132) );
  NAND U22411 ( .A(n14113), .B(n14114), .Z(n14112) );
  NANDN U22412 ( .A(n14115), .B(n14116), .Z(n14114) );
  NANDN U22413 ( .A(n14116), .B(n14115), .Z(n14111) );
  XOR U22414 ( .A(n14115), .B(n14117), .Z(N64131) );
  XNOR U22415 ( .A(n14113), .B(n14116), .Z(n14117) );
  NAND U22416 ( .A(n14118), .B(n14119), .Z(n14116) );
  NAND U22417 ( .A(n14120), .B(n14121), .Z(n14119) );
  NANDN U22418 ( .A(n14122), .B(n14123), .Z(n14121) );
  NANDN U22419 ( .A(n14123), .B(n14122), .Z(n14118) );
  AND U22420 ( .A(n14124), .B(n14125), .Z(n14113) );
  NAND U22421 ( .A(n14126), .B(n14127), .Z(n14125) );
  NANDN U22422 ( .A(n14128), .B(n14129), .Z(n14127) );
  NANDN U22423 ( .A(n14129), .B(n14128), .Z(n14124) );
  IV U22424 ( .A(n14130), .Z(n14129) );
  AND U22425 ( .A(n14131), .B(n14132), .Z(n14115) );
  NAND U22426 ( .A(n14133), .B(n14134), .Z(n14132) );
  NANDN U22427 ( .A(n14135), .B(n14136), .Z(n14134) );
  NANDN U22428 ( .A(n14136), .B(n14135), .Z(n14131) );
  XOR U22429 ( .A(n14128), .B(n14137), .Z(N64130) );
  XNOR U22430 ( .A(n14126), .B(n14130), .Z(n14137) );
  XOR U22431 ( .A(n14123), .B(n14138), .Z(n14130) );
  XNOR U22432 ( .A(n14120), .B(n14122), .Z(n14138) );
  AND U22433 ( .A(n14139), .B(n14140), .Z(n14122) );
  NANDN U22434 ( .A(n14141), .B(n14142), .Z(n14140) );
  OR U22435 ( .A(n14143), .B(n14144), .Z(n14142) );
  IV U22436 ( .A(n14145), .Z(n14144) );
  NANDN U22437 ( .A(n14145), .B(n14143), .Z(n14139) );
  AND U22438 ( .A(n14146), .B(n14147), .Z(n14120) );
  NAND U22439 ( .A(n14148), .B(n14149), .Z(n14147) );
  NANDN U22440 ( .A(n14150), .B(n14151), .Z(n14149) );
  NANDN U22441 ( .A(n14151), .B(n14150), .Z(n14146) );
  IV U22442 ( .A(n14152), .Z(n14151) );
  NAND U22443 ( .A(n14153), .B(n14154), .Z(n14123) );
  NANDN U22444 ( .A(n14155), .B(n14156), .Z(n14154) );
  NANDN U22445 ( .A(n14157), .B(n14158), .Z(n14156) );
  NANDN U22446 ( .A(n14158), .B(n14157), .Z(n14153) );
  IV U22447 ( .A(n14159), .Z(n14157) );
  AND U22448 ( .A(n14160), .B(n14161), .Z(n14126) );
  NAND U22449 ( .A(n14162), .B(n14163), .Z(n14161) );
  NANDN U22450 ( .A(n14164), .B(n14165), .Z(n14163) );
  NANDN U22451 ( .A(n14165), .B(n14164), .Z(n14160) );
  XOR U22452 ( .A(n14136), .B(n14166), .Z(n14128) );
  XNOR U22453 ( .A(n14133), .B(n14135), .Z(n14166) );
  AND U22454 ( .A(n14167), .B(n14168), .Z(n14135) );
  NANDN U22455 ( .A(n14169), .B(n14170), .Z(n14168) );
  OR U22456 ( .A(n14171), .B(n14172), .Z(n14170) );
  IV U22457 ( .A(n14173), .Z(n14172) );
  NANDN U22458 ( .A(n14173), .B(n14171), .Z(n14167) );
  AND U22459 ( .A(n14174), .B(n14175), .Z(n14133) );
  NAND U22460 ( .A(n14176), .B(n14177), .Z(n14175) );
  NANDN U22461 ( .A(n14178), .B(n14179), .Z(n14177) );
  NANDN U22462 ( .A(n14179), .B(n14178), .Z(n14174) );
  IV U22463 ( .A(n14180), .Z(n14179) );
  NAND U22464 ( .A(n14181), .B(n14182), .Z(n14136) );
  NANDN U22465 ( .A(n14183), .B(n14184), .Z(n14182) );
  NANDN U22466 ( .A(n14185), .B(n14186), .Z(n14184) );
  NANDN U22467 ( .A(n14186), .B(n14185), .Z(n14181) );
  IV U22468 ( .A(n14187), .Z(n14185) );
  XOR U22469 ( .A(n14162), .B(n14188), .Z(N64129) );
  XNOR U22470 ( .A(n14165), .B(n14164), .Z(n14188) );
  XNOR U22471 ( .A(n14176), .B(n14189), .Z(n14164) );
  XNOR U22472 ( .A(n14180), .B(n14178), .Z(n14189) );
  XOR U22473 ( .A(n14186), .B(n14190), .Z(n14178) );
  XNOR U22474 ( .A(n14183), .B(n14187), .Z(n14190) );
  AND U22475 ( .A(n14191), .B(n14192), .Z(n14187) );
  NAND U22476 ( .A(n14193), .B(n14194), .Z(n14192) );
  NAND U22477 ( .A(n14195), .B(n14196), .Z(n14191) );
  AND U22478 ( .A(n14197), .B(n14198), .Z(n14183) );
  NAND U22479 ( .A(n14199), .B(n14200), .Z(n14198) );
  NAND U22480 ( .A(n14201), .B(n14202), .Z(n14197) );
  NANDN U22481 ( .A(n14203), .B(n14204), .Z(n14186) );
  ANDN U22482 ( .B(n14205), .A(n14206), .Z(n14180) );
  XNOR U22483 ( .A(n14171), .B(n14207), .Z(n14176) );
  XNOR U22484 ( .A(n14169), .B(n14173), .Z(n14207) );
  AND U22485 ( .A(n14208), .B(n14209), .Z(n14173) );
  NAND U22486 ( .A(n14210), .B(n14211), .Z(n14209) );
  NAND U22487 ( .A(n14212), .B(n14213), .Z(n14208) );
  AND U22488 ( .A(n14214), .B(n14215), .Z(n14169) );
  NAND U22489 ( .A(n14216), .B(n14217), .Z(n14215) );
  NAND U22490 ( .A(n14218), .B(n14219), .Z(n14214) );
  AND U22491 ( .A(n14220), .B(n14221), .Z(n14171) );
  NAND U22492 ( .A(n14222), .B(n14223), .Z(n14165) );
  XNOR U22493 ( .A(n14148), .B(n14224), .Z(n14162) );
  XNOR U22494 ( .A(n14152), .B(n14150), .Z(n14224) );
  XOR U22495 ( .A(n14158), .B(n14225), .Z(n14150) );
  XNOR U22496 ( .A(n14155), .B(n14159), .Z(n14225) );
  AND U22497 ( .A(n14226), .B(n14227), .Z(n14159) );
  NAND U22498 ( .A(n14228), .B(n14229), .Z(n14227) );
  NAND U22499 ( .A(n14230), .B(n14231), .Z(n14226) );
  AND U22500 ( .A(n14232), .B(n14233), .Z(n14155) );
  NAND U22501 ( .A(n14234), .B(n14235), .Z(n14233) );
  NAND U22502 ( .A(n14236), .B(n14237), .Z(n14232) );
  NANDN U22503 ( .A(n14238), .B(n14239), .Z(n14158) );
  ANDN U22504 ( .B(n14240), .A(n14241), .Z(n14152) );
  XNOR U22505 ( .A(n14143), .B(n14242), .Z(n14148) );
  XNOR U22506 ( .A(n14141), .B(n14145), .Z(n14242) );
  AND U22507 ( .A(n14243), .B(n14244), .Z(n14145) );
  NAND U22508 ( .A(n14245), .B(n14246), .Z(n14244) );
  NAND U22509 ( .A(n14247), .B(n14248), .Z(n14243) );
  AND U22510 ( .A(n14249), .B(n14250), .Z(n14141) );
  NAND U22511 ( .A(n14251), .B(n14252), .Z(n14250) );
  NAND U22512 ( .A(n14253), .B(n14254), .Z(n14249) );
  AND U22513 ( .A(n14255), .B(n14256), .Z(n14143) );
  XOR U22514 ( .A(n14223), .B(n14222), .Z(N64128) );
  XNOR U22515 ( .A(n14240), .B(n14241), .Z(n14222) );
  XNOR U22516 ( .A(n14255), .B(n14256), .Z(n14241) );
  XOR U22517 ( .A(n14252), .B(n14251), .Z(n14256) );
  XOR U22518 ( .A(y[6540]), .B(x[6540]), .Z(n14251) );
  XOR U22519 ( .A(n14254), .B(n14253), .Z(n14252) );
  XOR U22520 ( .A(y[6542]), .B(x[6542]), .Z(n14253) );
  XOR U22521 ( .A(y[6541]), .B(x[6541]), .Z(n14254) );
  XOR U22522 ( .A(n14246), .B(n14245), .Z(n14255) );
  XOR U22523 ( .A(n14248), .B(n14247), .Z(n14245) );
  XOR U22524 ( .A(y[6539]), .B(x[6539]), .Z(n14247) );
  XOR U22525 ( .A(y[6538]), .B(x[6538]), .Z(n14248) );
  XOR U22526 ( .A(y[6537]), .B(x[6537]), .Z(n14246) );
  XNOR U22527 ( .A(n14239), .B(n14238), .Z(n14240) );
  XNOR U22528 ( .A(n14235), .B(n14234), .Z(n14238) );
  XOR U22529 ( .A(n14237), .B(n14236), .Z(n14234) );
  XOR U22530 ( .A(y[6536]), .B(x[6536]), .Z(n14236) );
  XOR U22531 ( .A(y[6535]), .B(x[6535]), .Z(n14237) );
  XOR U22532 ( .A(y[6534]), .B(x[6534]), .Z(n14235) );
  XOR U22533 ( .A(n14229), .B(n14228), .Z(n14239) );
  XOR U22534 ( .A(n14231), .B(n14230), .Z(n14228) );
  XOR U22535 ( .A(y[6533]), .B(x[6533]), .Z(n14230) );
  XOR U22536 ( .A(y[6532]), .B(x[6532]), .Z(n14231) );
  XOR U22537 ( .A(y[6531]), .B(x[6531]), .Z(n14229) );
  XNOR U22538 ( .A(n14205), .B(n14206), .Z(n14223) );
  XNOR U22539 ( .A(n14220), .B(n14221), .Z(n14206) );
  XOR U22540 ( .A(n14217), .B(n14216), .Z(n14221) );
  XOR U22541 ( .A(y[6528]), .B(x[6528]), .Z(n14216) );
  XOR U22542 ( .A(n14219), .B(n14218), .Z(n14217) );
  XOR U22543 ( .A(y[6530]), .B(x[6530]), .Z(n14218) );
  XOR U22544 ( .A(y[6529]), .B(x[6529]), .Z(n14219) );
  XOR U22545 ( .A(n14211), .B(n14210), .Z(n14220) );
  XOR U22546 ( .A(n14213), .B(n14212), .Z(n14210) );
  XOR U22547 ( .A(y[6527]), .B(x[6527]), .Z(n14212) );
  XOR U22548 ( .A(y[6526]), .B(x[6526]), .Z(n14213) );
  XOR U22549 ( .A(y[6525]), .B(x[6525]), .Z(n14211) );
  XNOR U22550 ( .A(n14204), .B(n14203), .Z(n14205) );
  XNOR U22551 ( .A(n14200), .B(n14199), .Z(n14203) );
  XOR U22552 ( .A(n14202), .B(n14201), .Z(n14199) );
  XOR U22553 ( .A(y[6524]), .B(x[6524]), .Z(n14201) );
  XOR U22554 ( .A(y[6523]), .B(x[6523]), .Z(n14202) );
  XOR U22555 ( .A(y[6522]), .B(x[6522]), .Z(n14200) );
  XOR U22556 ( .A(n14194), .B(n14193), .Z(n14204) );
  XOR U22557 ( .A(n14196), .B(n14195), .Z(n14193) );
  XOR U22558 ( .A(y[6521]), .B(x[6521]), .Z(n14195) );
  XOR U22559 ( .A(y[6520]), .B(x[6520]), .Z(n14196) );
  XOR U22560 ( .A(y[6519]), .B(x[6519]), .Z(n14194) );
  NAND U22561 ( .A(n14257), .B(n14258), .Z(N64119) );
  NAND U22562 ( .A(n14259), .B(n14260), .Z(n14258) );
  NANDN U22563 ( .A(n14261), .B(n14262), .Z(n14260) );
  NANDN U22564 ( .A(n14262), .B(n14261), .Z(n14257) );
  XOR U22565 ( .A(n14261), .B(n14263), .Z(N64118) );
  XNOR U22566 ( .A(n14259), .B(n14262), .Z(n14263) );
  NAND U22567 ( .A(n14264), .B(n14265), .Z(n14262) );
  NAND U22568 ( .A(n14266), .B(n14267), .Z(n14265) );
  NANDN U22569 ( .A(n14268), .B(n14269), .Z(n14267) );
  NANDN U22570 ( .A(n14269), .B(n14268), .Z(n14264) );
  AND U22571 ( .A(n14270), .B(n14271), .Z(n14259) );
  NAND U22572 ( .A(n14272), .B(n14273), .Z(n14271) );
  NANDN U22573 ( .A(n14274), .B(n14275), .Z(n14273) );
  NANDN U22574 ( .A(n14275), .B(n14274), .Z(n14270) );
  IV U22575 ( .A(n14276), .Z(n14275) );
  AND U22576 ( .A(n14277), .B(n14278), .Z(n14261) );
  NAND U22577 ( .A(n14279), .B(n14280), .Z(n14278) );
  NANDN U22578 ( .A(n14281), .B(n14282), .Z(n14280) );
  NANDN U22579 ( .A(n14282), .B(n14281), .Z(n14277) );
  XOR U22580 ( .A(n14274), .B(n14283), .Z(N64117) );
  XNOR U22581 ( .A(n14272), .B(n14276), .Z(n14283) );
  XOR U22582 ( .A(n14269), .B(n14284), .Z(n14276) );
  XNOR U22583 ( .A(n14266), .B(n14268), .Z(n14284) );
  AND U22584 ( .A(n14285), .B(n14286), .Z(n14268) );
  NANDN U22585 ( .A(n14287), .B(n14288), .Z(n14286) );
  OR U22586 ( .A(n14289), .B(n14290), .Z(n14288) );
  IV U22587 ( .A(n14291), .Z(n14290) );
  NANDN U22588 ( .A(n14291), .B(n14289), .Z(n14285) );
  AND U22589 ( .A(n14292), .B(n14293), .Z(n14266) );
  NAND U22590 ( .A(n14294), .B(n14295), .Z(n14293) );
  NANDN U22591 ( .A(n14296), .B(n14297), .Z(n14295) );
  NANDN U22592 ( .A(n14297), .B(n14296), .Z(n14292) );
  IV U22593 ( .A(n14298), .Z(n14297) );
  NAND U22594 ( .A(n14299), .B(n14300), .Z(n14269) );
  NANDN U22595 ( .A(n14301), .B(n14302), .Z(n14300) );
  NANDN U22596 ( .A(n14303), .B(n14304), .Z(n14302) );
  NANDN U22597 ( .A(n14304), .B(n14303), .Z(n14299) );
  IV U22598 ( .A(n14305), .Z(n14303) );
  AND U22599 ( .A(n14306), .B(n14307), .Z(n14272) );
  NAND U22600 ( .A(n14308), .B(n14309), .Z(n14307) );
  NANDN U22601 ( .A(n14310), .B(n14311), .Z(n14309) );
  NANDN U22602 ( .A(n14311), .B(n14310), .Z(n14306) );
  XOR U22603 ( .A(n14282), .B(n14312), .Z(n14274) );
  XNOR U22604 ( .A(n14279), .B(n14281), .Z(n14312) );
  AND U22605 ( .A(n14313), .B(n14314), .Z(n14281) );
  NANDN U22606 ( .A(n14315), .B(n14316), .Z(n14314) );
  OR U22607 ( .A(n14317), .B(n14318), .Z(n14316) );
  IV U22608 ( .A(n14319), .Z(n14318) );
  NANDN U22609 ( .A(n14319), .B(n14317), .Z(n14313) );
  AND U22610 ( .A(n14320), .B(n14321), .Z(n14279) );
  NAND U22611 ( .A(n14322), .B(n14323), .Z(n14321) );
  NANDN U22612 ( .A(n14324), .B(n14325), .Z(n14323) );
  NANDN U22613 ( .A(n14325), .B(n14324), .Z(n14320) );
  IV U22614 ( .A(n14326), .Z(n14325) );
  NAND U22615 ( .A(n14327), .B(n14328), .Z(n14282) );
  NANDN U22616 ( .A(n14329), .B(n14330), .Z(n14328) );
  NANDN U22617 ( .A(n14331), .B(n14332), .Z(n14330) );
  NANDN U22618 ( .A(n14332), .B(n14331), .Z(n14327) );
  IV U22619 ( .A(n14333), .Z(n14331) );
  XOR U22620 ( .A(n14308), .B(n14334), .Z(N64116) );
  XNOR U22621 ( .A(n14311), .B(n14310), .Z(n14334) );
  XNOR U22622 ( .A(n14322), .B(n14335), .Z(n14310) );
  XNOR U22623 ( .A(n14326), .B(n14324), .Z(n14335) );
  XOR U22624 ( .A(n14332), .B(n14336), .Z(n14324) );
  XNOR U22625 ( .A(n14329), .B(n14333), .Z(n14336) );
  AND U22626 ( .A(n14337), .B(n14338), .Z(n14333) );
  NAND U22627 ( .A(n14339), .B(n14340), .Z(n14338) );
  NAND U22628 ( .A(n14341), .B(n14342), .Z(n14337) );
  AND U22629 ( .A(n14343), .B(n14344), .Z(n14329) );
  NAND U22630 ( .A(n14345), .B(n14346), .Z(n14344) );
  NAND U22631 ( .A(n14347), .B(n14348), .Z(n14343) );
  NANDN U22632 ( .A(n14349), .B(n14350), .Z(n14332) );
  ANDN U22633 ( .B(n14351), .A(n14352), .Z(n14326) );
  XNOR U22634 ( .A(n14317), .B(n14353), .Z(n14322) );
  XNOR U22635 ( .A(n14315), .B(n14319), .Z(n14353) );
  AND U22636 ( .A(n14354), .B(n14355), .Z(n14319) );
  NAND U22637 ( .A(n14356), .B(n14357), .Z(n14355) );
  NAND U22638 ( .A(n14358), .B(n14359), .Z(n14354) );
  AND U22639 ( .A(n14360), .B(n14361), .Z(n14315) );
  NAND U22640 ( .A(n14362), .B(n14363), .Z(n14361) );
  NAND U22641 ( .A(n14364), .B(n14365), .Z(n14360) );
  AND U22642 ( .A(n14366), .B(n14367), .Z(n14317) );
  NAND U22643 ( .A(n14368), .B(n14369), .Z(n14311) );
  XNOR U22644 ( .A(n14294), .B(n14370), .Z(n14308) );
  XNOR U22645 ( .A(n14298), .B(n14296), .Z(n14370) );
  XOR U22646 ( .A(n14304), .B(n14371), .Z(n14296) );
  XNOR U22647 ( .A(n14301), .B(n14305), .Z(n14371) );
  AND U22648 ( .A(n14372), .B(n14373), .Z(n14305) );
  NAND U22649 ( .A(n14374), .B(n14375), .Z(n14373) );
  NAND U22650 ( .A(n14376), .B(n14377), .Z(n14372) );
  AND U22651 ( .A(n14378), .B(n14379), .Z(n14301) );
  NAND U22652 ( .A(n14380), .B(n14381), .Z(n14379) );
  NAND U22653 ( .A(n14382), .B(n14383), .Z(n14378) );
  NANDN U22654 ( .A(n14384), .B(n14385), .Z(n14304) );
  ANDN U22655 ( .B(n14386), .A(n14387), .Z(n14298) );
  XNOR U22656 ( .A(n14289), .B(n14388), .Z(n14294) );
  XNOR U22657 ( .A(n14287), .B(n14291), .Z(n14388) );
  AND U22658 ( .A(n14389), .B(n14390), .Z(n14291) );
  NAND U22659 ( .A(n14391), .B(n14392), .Z(n14390) );
  NAND U22660 ( .A(n14393), .B(n14394), .Z(n14389) );
  AND U22661 ( .A(n14395), .B(n14396), .Z(n14287) );
  NAND U22662 ( .A(n14397), .B(n14398), .Z(n14396) );
  NAND U22663 ( .A(n14399), .B(n14400), .Z(n14395) );
  AND U22664 ( .A(n14401), .B(n14402), .Z(n14289) );
  XOR U22665 ( .A(n14369), .B(n14368), .Z(N64115) );
  XNOR U22666 ( .A(n14386), .B(n14387), .Z(n14368) );
  XNOR U22667 ( .A(n14401), .B(n14402), .Z(n14387) );
  XOR U22668 ( .A(n14398), .B(n14397), .Z(n14402) );
  XOR U22669 ( .A(y[6516]), .B(x[6516]), .Z(n14397) );
  XOR U22670 ( .A(n14400), .B(n14399), .Z(n14398) );
  XOR U22671 ( .A(y[6518]), .B(x[6518]), .Z(n14399) );
  XOR U22672 ( .A(y[6517]), .B(x[6517]), .Z(n14400) );
  XOR U22673 ( .A(n14392), .B(n14391), .Z(n14401) );
  XOR U22674 ( .A(n14394), .B(n14393), .Z(n14391) );
  XOR U22675 ( .A(y[6515]), .B(x[6515]), .Z(n14393) );
  XOR U22676 ( .A(y[6514]), .B(x[6514]), .Z(n14394) );
  XOR U22677 ( .A(y[6513]), .B(x[6513]), .Z(n14392) );
  XNOR U22678 ( .A(n14385), .B(n14384), .Z(n14386) );
  XNOR U22679 ( .A(n14381), .B(n14380), .Z(n14384) );
  XOR U22680 ( .A(n14383), .B(n14382), .Z(n14380) );
  XOR U22681 ( .A(y[6512]), .B(x[6512]), .Z(n14382) );
  XOR U22682 ( .A(y[6511]), .B(x[6511]), .Z(n14383) );
  XOR U22683 ( .A(y[6510]), .B(x[6510]), .Z(n14381) );
  XOR U22684 ( .A(n14375), .B(n14374), .Z(n14385) );
  XOR U22685 ( .A(n14377), .B(n14376), .Z(n14374) );
  XOR U22686 ( .A(y[6509]), .B(x[6509]), .Z(n14376) );
  XOR U22687 ( .A(y[6508]), .B(x[6508]), .Z(n14377) );
  XOR U22688 ( .A(y[6507]), .B(x[6507]), .Z(n14375) );
  XNOR U22689 ( .A(n14351), .B(n14352), .Z(n14369) );
  XNOR U22690 ( .A(n14366), .B(n14367), .Z(n14352) );
  XOR U22691 ( .A(n14363), .B(n14362), .Z(n14367) );
  XOR U22692 ( .A(y[6504]), .B(x[6504]), .Z(n14362) );
  XOR U22693 ( .A(n14365), .B(n14364), .Z(n14363) );
  XOR U22694 ( .A(y[6506]), .B(x[6506]), .Z(n14364) );
  XOR U22695 ( .A(y[6505]), .B(x[6505]), .Z(n14365) );
  XOR U22696 ( .A(n14357), .B(n14356), .Z(n14366) );
  XOR U22697 ( .A(n14359), .B(n14358), .Z(n14356) );
  XOR U22698 ( .A(y[6503]), .B(x[6503]), .Z(n14358) );
  XOR U22699 ( .A(y[6502]), .B(x[6502]), .Z(n14359) );
  XOR U22700 ( .A(y[6501]), .B(x[6501]), .Z(n14357) );
  XNOR U22701 ( .A(n14350), .B(n14349), .Z(n14351) );
  XNOR U22702 ( .A(n14346), .B(n14345), .Z(n14349) );
  XOR U22703 ( .A(n14348), .B(n14347), .Z(n14345) );
  XOR U22704 ( .A(y[6500]), .B(x[6500]), .Z(n14347) );
  XOR U22705 ( .A(y[6499]), .B(x[6499]), .Z(n14348) );
  XOR U22706 ( .A(y[6498]), .B(x[6498]), .Z(n14346) );
  XOR U22707 ( .A(n14340), .B(n14339), .Z(n14350) );
  XOR U22708 ( .A(n14342), .B(n14341), .Z(n14339) );
  XOR U22709 ( .A(y[6497]), .B(x[6497]), .Z(n14341) );
  XOR U22710 ( .A(y[6496]), .B(x[6496]), .Z(n14342) );
  XOR U22711 ( .A(y[6495]), .B(x[6495]), .Z(n14340) );
  NAND U22712 ( .A(n14403), .B(n14404), .Z(N64106) );
  NAND U22713 ( .A(n14405), .B(n14406), .Z(n14404) );
  NANDN U22714 ( .A(n14407), .B(n14408), .Z(n14406) );
  NANDN U22715 ( .A(n14408), .B(n14407), .Z(n14403) );
  XOR U22716 ( .A(n14407), .B(n14409), .Z(N64105) );
  XNOR U22717 ( .A(n14405), .B(n14408), .Z(n14409) );
  NAND U22718 ( .A(n14410), .B(n14411), .Z(n14408) );
  NAND U22719 ( .A(n14412), .B(n14413), .Z(n14411) );
  NANDN U22720 ( .A(n14414), .B(n14415), .Z(n14413) );
  NANDN U22721 ( .A(n14415), .B(n14414), .Z(n14410) );
  AND U22722 ( .A(n14416), .B(n14417), .Z(n14405) );
  NAND U22723 ( .A(n14418), .B(n14419), .Z(n14417) );
  NANDN U22724 ( .A(n14420), .B(n14421), .Z(n14419) );
  NANDN U22725 ( .A(n14421), .B(n14420), .Z(n14416) );
  IV U22726 ( .A(n14422), .Z(n14421) );
  AND U22727 ( .A(n14423), .B(n14424), .Z(n14407) );
  NAND U22728 ( .A(n14425), .B(n14426), .Z(n14424) );
  NANDN U22729 ( .A(n14427), .B(n14428), .Z(n14426) );
  NANDN U22730 ( .A(n14428), .B(n14427), .Z(n14423) );
  XOR U22731 ( .A(n14420), .B(n14429), .Z(N64104) );
  XNOR U22732 ( .A(n14418), .B(n14422), .Z(n14429) );
  XOR U22733 ( .A(n14415), .B(n14430), .Z(n14422) );
  XNOR U22734 ( .A(n14412), .B(n14414), .Z(n14430) );
  AND U22735 ( .A(n14431), .B(n14432), .Z(n14414) );
  NANDN U22736 ( .A(n14433), .B(n14434), .Z(n14432) );
  OR U22737 ( .A(n14435), .B(n14436), .Z(n14434) );
  IV U22738 ( .A(n14437), .Z(n14436) );
  NANDN U22739 ( .A(n14437), .B(n14435), .Z(n14431) );
  AND U22740 ( .A(n14438), .B(n14439), .Z(n14412) );
  NAND U22741 ( .A(n14440), .B(n14441), .Z(n14439) );
  NANDN U22742 ( .A(n14442), .B(n14443), .Z(n14441) );
  NANDN U22743 ( .A(n14443), .B(n14442), .Z(n14438) );
  IV U22744 ( .A(n14444), .Z(n14443) );
  NAND U22745 ( .A(n14445), .B(n14446), .Z(n14415) );
  NANDN U22746 ( .A(n14447), .B(n14448), .Z(n14446) );
  NANDN U22747 ( .A(n14449), .B(n14450), .Z(n14448) );
  NANDN U22748 ( .A(n14450), .B(n14449), .Z(n14445) );
  IV U22749 ( .A(n14451), .Z(n14449) );
  AND U22750 ( .A(n14452), .B(n14453), .Z(n14418) );
  NAND U22751 ( .A(n14454), .B(n14455), .Z(n14453) );
  NANDN U22752 ( .A(n14456), .B(n14457), .Z(n14455) );
  NANDN U22753 ( .A(n14457), .B(n14456), .Z(n14452) );
  XOR U22754 ( .A(n14428), .B(n14458), .Z(n14420) );
  XNOR U22755 ( .A(n14425), .B(n14427), .Z(n14458) );
  AND U22756 ( .A(n14459), .B(n14460), .Z(n14427) );
  NANDN U22757 ( .A(n14461), .B(n14462), .Z(n14460) );
  OR U22758 ( .A(n14463), .B(n14464), .Z(n14462) );
  IV U22759 ( .A(n14465), .Z(n14464) );
  NANDN U22760 ( .A(n14465), .B(n14463), .Z(n14459) );
  AND U22761 ( .A(n14466), .B(n14467), .Z(n14425) );
  NAND U22762 ( .A(n14468), .B(n14469), .Z(n14467) );
  NANDN U22763 ( .A(n14470), .B(n14471), .Z(n14469) );
  NANDN U22764 ( .A(n14471), .B(n14470), .Z(n14466) );
  IV U22765 ( .A(n14472), .Z(n14471) );
  NAND U22766 ( .A(n14473), .B(n14474), .Z(n14428) );
  NANDN U22767 ( .A(n14475), .B(n14476), .Z(n14474) );
  NANDN U22768 ( .A(n14477), .B(n14478), .Z(n14476) );
  NANDN U22769 ( .A(n14478), .B(n14477), .Z(n14473) );
  IV U22770 ( .A(n14479), .Z(n14477) );
  XOR U22771 ( .A(n14454), .B(n14480), .Z(N64103) );
  XNOR U22772 ( .A(n14457), .B(n14456), .Z(n14480) );
  XNOR U22773 ( .A(n14468), .B(n14481), .Z(n14456) );
  XNOR U22774 ( .A(n14472), .B(n14470), .Z(n14481) );
  XOR U22775 ( .A(n14478), .B(n14482), .Z(n14470) );
  XNOR U22776 ( .A(n14475), .B(n14479), .Z(n14482) );
  AND U22777 ( .A(n14483), .B(n14484), .Z(n14479) );
  NAND U22778 ( .A(n14485), .B(n14486), .Z(n14484) );
  NAND U22779 ( .A(n14487), .B(n14488), .Z(n14483) );
  AND U22780 ( .A(n14489), .B(n14490), .Z(n14475) );
  NAND U22781 ( .A(n14491), .B(n14492), .Z(n14490) );
  NAND U22782 ( .A(n14493), .B(n14494), .Z(n14489) );
  NANDN U22783 ( .A(n14495), .B(n14496), .Z(n14478) );
  ANDN U22784 ( .B(n14497), .A(n14498), .Z(n14472) );
  XNOR U22785 ( .A(n14463), .B(n14499), .Z(n14468) );
  XNOR U22786 ( .A(n14461), .B(n14465), .Z(n14499) );
  AND U22787 ( .A(n14500), .B(n14501), .Z(n14465) );
  NAND U22788 ( .A(n14502), .B(n14503), .Z(n14501) );
  NAND U22789 ( .A(n14504), .B(n14505), .Z(n14500) );
  AND U22790 ( .A(n14506), .B(n14507), .Z(n14461) );
  NAND U22791 ( .A(n14508), .B(n14509), .Z(n14507) );
  NAND U22792 ( .A(n14510), .B(n14511), .Z(n14506) );
  AND U22793 ( .A(n14512), .B(n14513), .Z(n14463) );
  NAND U22794 ( .A(n14514), .B(n14515), .Z(n14457) );
  XNOR U22795 ( .A(n14440), .B(n14516), .Z(n14454) );
  XNOR U22796 ( .A(n14444), .B(n14442), .Z(n14516) );
  XOR U22797 ( .A(n14450), .B(n14517), .Z(n14442) );
  XNOR U22798 ( .A(n14447), .B(n14451), .Z(n14517) );
  AND U22799 ( .A(n14518), .B(n14519), .Z(n14451) );
  NAND U22800 ( .A(n14520), .B(n14521), .Z(n14519) );
  NAND U22801 ( .A(n14522), .B(n14523), .Z(n14518) );
  AND U22802 ( .A(n14524), .B(n14525), .Z(n14447) );
  NAND U22803 ( .A(n14526), .B(n14527), .Z(n14525) );
  NAND U22804 ( .A(n14528), .B(n14529), .Z(n14524) );
  NANDN U22805 ( .A(n14530), .B(n14531), .Z(n14450) );
  ANDN U22806 ( .B(n14532), .A(n14533), .Z(n14444) );
  XNOR U22807 ( .A(n14435), .B(n14534), .Z(n14440) );
  XNOR U22808 ( .A(n14433), .B(n14437), .Z(n14534) );
  AND U22809 ( .A(n14535), .B(n14536), .Z(n14437) );
  NAND U22810 ( .A(n14537), .B(n14538), .Z(n14536) );
  NAND U22811 ( .A(n14539), .B(n14540), .Z(n14535) );
  AND U22812 ( .A(n14541), .B(n14542), .Z(n14433) );
  NAND U22813 ( .A(n14543), .B(n14544), .Z(n14542) );
  NAND U22814 ( .A(n14545), .B(n14546), .Z(n14541) );
  AND U22815 ( .A(n14547), .B(n14548), .Z(n14435) );
  XOR U22816 ( .A(n14515), .B(n14514), .Z(N64102) );
  XNOR U22817 ( .A(n14532), .B(n14533), .Z(n14514) );
  XNOR U22818 ( .A(n14547), .B(n14548), .Z(n14533) );
  XOR U22819 ( .A(n14544), .B(n14543), .Z(n14548) );
  XOR U22820 ( .A(y[6492]), .B(x[6492]), .Z(n14543) );
  XOR U22821 ( .A(n14546), .B(n14545), .Z(n14544) );
  XOR U22822 ( .A(y[6494]), .B(x[6494]), .Z(n14545) );
  XOR U22823 ( .A(y[6493]), .B(x[6493]), .Z(n14546) );
  XOR U22824 ( .A(n14538), .B(n14537), .Z(n14547) );
  XOR U22825 ( .A(n14540), .B(n14539), .Z(n14537) );
  XOR U22826 ( .A(y[6491]), .B(x[6491]), .Z(n14539) );
  XOR U22827 ( .A(y[6490]), .B(x[6490]), .Z(n14540) );
  XOR U22828 ( .A(y[6489]), .B(x[6489]), .Z(n14538) );
  XNOR U22829 ( .A(n14531), .B(n14530), .Z(n14532) );
  XNOR U22830 ( .A(n14527), .B(n14526), .Z(n14530) );
  XOR U22831 ( .A(n14529), .B(n14528), .Z(n14526) );
  XOR U22832 ( .A(y[6488]), .B(x[6488]), .Z(n14528) );
  XOR U22833 ( .A(y[6487]), .B(x[6487]), .Z(n14529) );
  XOR U22834 ( .A(y[6486]), .B(x[6486]), .Z(n14527) );
  XOR U22835 ( .A(n14521), .B(n14520), .Z(n14531) );
  XOR U22836 ( .A(n14523), .B(n14522), .Z(n14520) );
  XOR U22837 ( .A(y[6485]), .B(x[6485]), .Z(n14522) );
  XOR U22838 ( .A(y[6484]), .B(x[6484]), .Z(n14523) );
  XOR U22839 ( .A(y[6483]), .B(x[6483]), .Z(n14521) );
  XNOR U22840 ( .A(n14497), .B(n14498), .Z(n14515) );
  XNOR U22841 ( .A(n14512), .B(n14513), .Z(n14498) );
  XOR U22842 ( .A(n14509), .B(n14508), .Z(n14513) );
  XOR U22843 ( .A(y[6480]), .B(x[6480]), .Z(n14508) );
  XOR U22844 ( .A(n14511), .B(n14510), .Z(n14509) );
  XOR U22845 ( .A(y[6482]), .B(x[6482]), .Z(n14510) );
  XOR U22846 ( .A(y[6481]), .B(x[6481]), .Z(n14511) );
  XOR U22847 ( .A(n14503), .B(n14502), .Z(n14512) );
  XOR U22848 ( .A(n14505), .B(n14504), .Z(n14502) );
  XOR U22849 ( .A(y[6479]), .B(x[6479]), .Z(n14504) );
  XOR U22850 ( .A(y[6478]), .B(x[6478]), .Z(n14505) );
  XOR U22851 ( .A(y[6477]), .B(x[6477]), .Z(n14503) );
  XNOR U22852 ( .A(n14496), .B(n14495), .Z(n14497) );
  XNOR U22853 ( .A(n14492), .B(n14491), .Z(n14495) );
  XOR U22854 ( .A(n14494), .B(n14493), .Z(n14491) );
  XOR U22855 ( .A(y[6476]), .B(x[6476]), .Z(n14493) );
  XOR U22856 ( .A(y[6475]), .B(x[6475]), .Z(n14494) );
  XOR U22857 ( .A(y[6474]), .B(x[6474]), .Z(n14492) );
  XOR U22858 ( .A(n14486), .B(n14485), .Z(n14496) );
  XOR U22859 ( .A(n14488), .B(n14487), .Z(n14485) );
  XOR U22860 ( .A(y[6473]), .B(x[6473]), .Z(n14487) );
  XOR U22861 ( .A(y[6472]), .B(x[6472]), .Z(n14488) );
  XOR U22862 ( .A(y[6471]), .B(x[6471]), .Z(n14486) );
  NAND U22863 ( .A(n14549), .B(n14550), .Z(N64093) );
  NAND U22864 ( .A(n14551), .B(n14552), .Z(n14550) );
  NANDN U22865 ( .A(n14553), .B(n14554), .Z(n14552) );
  NANDN U22866 ( .A(n14554), .B(n14553), .Z(n14549) );
  XOR U22867 ( .A(n14553), .B(n14555), .Z(N64092) );
  XNOR U22868 ( .A(n14551), .B(n14554), .Z(n14555) );
  NAND U22869 ( .A(n14556), .B(n14557), .Z(n14554) );
  NAND U22870 ( .A(n14558), .B(n14559), .Z(n14557) );
  NANDN U22871 ( .A(n14560), .B(n14561), .Z(n14559) );
  NANDN U22872 ( .A(n14561), .B(n14560), .Z(n14556) );
  AND U22873 ( .A(n14562), .B(n14563), .Z(n14551) );
  NAND U22874 ( .A(n14564), .B(n14565), .Z(n14563) );
  NANDN U22875 ( .A(n14566), .B(n14567), .Z(n14565) );
  NANDN U22876 ( .A(n14567), .B(n14566), .Z(n14562) );
  IV U22877 ( .A(n14568), .Z(n14567) );
  AND U22878 ( .A(n14569), .B(n14570), .Z(n14553) );
  NAND U22879 ( .A(n14571), .B(n14572), .Z(n14570) );
  NANDN U22880 ( .A(n14573), .B(n14574), .Z(n14572) );
  NANDN U22881 ( .A(n14574), .B(n14573), .Z(n14569) );
  XOR U22882 ( .A(n14566), .B(n14575), .Z(N64091) );
  XNOR U22883 ( .A(n14564), .B(n14568), .Z(n14575) );
  XOR U22884 ( .A(n14561), .B(n14576), .Z(n14568) );
  XNOR U22885 ( .A(n14558), .B(n14560), .Z(n14576) );
  AND U22886 ( .A(n14577), .B(n14578), .Z(n14560) );
  NANDN U22887 ( .A(n14579), .B(n14580), .Z(n14578) );
  OR U22888 ( .A(n14581), .B(n14582), .Z(n14580) );
  IV U22889 ( .A(n14583), .Z(n14582) );
  NANDN U22890 ( .A(n14583), .B(n14581), .Z(n14577) );
  AND U22891 ( .A(n14584), .B(n14585), .Z(n14558) );
  NAND U22892 ( .A(n14586), .B(n14587), .Z(n14585) );
  NANDN U22893 ( .A(n14588), .B(n14589), .Z(n14587) );
  NANDN U22894 ( .A(n14589), .B(n14588), .Z(n14584) );
  IV U22895 ( .A(n14590), .Z(n14589) );
  NAND U22896 ( .A(n14591), .B(n14592), .Z(n14561) );
  NANDN U22897 ( .A(n14593), .B(n14594), .Z(n14592) );
  NANDN U22898 ( .A(n14595), .B(n14596), .Z(n14594) );
  NANDN U22899 ( .A(n14596), .B(n14595), .Z(n14591) );
  IV U22900 ( .A(n14597), .Z(n14595) );
  AND U22901 ( .A(n14598), .B(n14599), .Z(n14564) );
  NAND U22902 ( .A(n14600), .B(n14601), .Z(n14599) );
  NANDN U22903 ( .A(n14602), .B(n14603), .Z(n14601) );
  NANDN U22904 ( .A(n14603), .B(n14602), .Z(n14598) );
  XOR U22905 ( .A(n14574), .B(n14604), .Z(n14566) );
  XNOR U22906 ( .A(n14571), .B(n14573), .Z(n14604) );
  AND U22907 ( .A(n14605), .B(n14606), .Z(n14573) );
  NANDN U22908 ( .A(n14607), .B(n14608), .Z(n14606) );
  OR U22909 ( .A(n14609), .B(n14610), .Z(n14608) );
  IV U22910 ( .A(n14611), .Z(n14610) );
  NANDN U22911 ( .A(n14611), .B(n14609), .Z(n14605) );
  AND U22912 ( .A(n14612), .B(n14613), .Z(n14571) );
  NAND U22913 ( .A(n14614), .B(n14615), .Z(n14613) );
  NANDN U22914 ( .A(n14616), .B(n14617), .Z(n14615) );
  NANDN U22915 ( .A(n14617), .B(n14616), .Z(n14612) );
  IV U22916 ( .A(n14618), .Z(n14617) );
  NAND U22917 ( .A(n14619), .B(n14620), .Z(n14574) );
  NANDN U22918 ( .A(n14621), .B(n14622), .Z(n14620) );
  NANDN U22919 ( .A(n14623), .B(n14624), .Z(n14622) );
  NANDN U22920 ( .A(n14624), .B(n14623), .Z(n14619) );
  IV U22921 ( .A(n14625), .Z(n14623) );
  XOR U22922 ( .A(n14600), .B(n14626), .Z(N64090) );
  XNOR U22923 ( .A(n14603), .B(n14602), .Z(n14626) );
  XNOR U22924 ( .A(n14614), .B(n14627), .Z(n14602) );
  XNOR U22925 ( .A(n14618), .B(n14616), .Z(n14627) );
  XOR U22926 ( .A(n14624), .B(n14628), .Z(n14616) );
  XNOR U22927 ( .A(n14621), .B(n14625), .Z(n14628) );
  AND U22928 ( .A(n14629), .B(n14630), .Z(n14625) );
  NAND U22929 ( .A(n14631), .B(n14632), .Z(n14630) );
  NAND U22930 ( .A(n14633), .B(n14634), .Z(n14629) );
  AND U22931 ( .A(n14635), .B(n14636), .Z(n14621) );
  NAND U22932 ( .A(n14637), .B(n14638), .Z(n14636) );
  NAND U22933 ( .A(n14639), .B(n14640), .Z(n14635) );
  NANDN U22934 ( .A(n14641), .B(n14642), .Z(n14624) );
  ANDN U22935 ( .B(n14643), .A(n14644), .Z(n14618) );
  XNOR U22936 ( .A(n14609), .B(n14645), .Z(n14614) );
  XNOR U22937 ( .A(n14607), .B(n14611), .Z(n14645) );
  AND U22938 ( .A(n14646), .B(n14647), .Z(n14611) );
  NAND U22939 ( .A(n14648), .B(n14649), .Z(n14647) );
  NAND U22940 ( .A(n14650), .B(n14651), .Z(n14646) );
  AND U22941 ( .A(n14652), .B(n14653), .Z(n14607) );
  NAND U22942 ( .A(n14654), .B(n14655), .Z(n14653) );
  NAND U22943 ( .A(n14656), .B(n14657), .Z(n14652) );
  AND U22944 ( .A(n14658), .B(n14659), .Z(n14609) );
  NAND U22945 ( .A(n14660), .B(n14661), .Z(n14603) );
  XNOR U22946 ( .A(n14586), .B(n14662), .Z(n14600) );
  XNOR U22947 ( .A(n14590), .B(n14588), .Z(n14662) );
  XOR U22948 ( .A(n14596), .B(n14663), .Z(n14588) );
  XNOR U22949 ( .A(n14593), .B(n14597), .Z(n14663) );
  AND U22950 ( .A(n14664), .B(n14665), .Z(n14597) );
  NAND U22951 ( .A(n14666), .B(n14667), .Z(n14665) );
  NAND U22952 ( .A(n14668), .B(n14669), .Z(n14664) );
  AND U22953 ( .A(n14670), .B(n14671), .Z(n14593) );
  NAND U22954 ( .A(n14672), .B(n14673), .Z(n14671) );
  NAND U22955 ( .A(n14674), .B(n14675), .Z(n14670) );
  NANDN U22956 ( .A(n14676), .B(n14677), .Z(n14596) );
  ANDN U22957 ( .B(n14678), .A(n14679), .Z(n14590) );
  XNOR U22958 ( .A(n14581), .B(n14680), .Z(n14586) );
  XNOR U22959 ( .A(n14579), .B(n14583), .Z(n14680) );
  AND U22960 ( .A(n14681), .B(n14682), .Z(n14583) );
  NAND U22961 ( .A(n14683), .B(n14684), .Z(n14682) );
  NAND U22962 ( .A(n14685), .B(n14686), .Z(n14681) );
  AND U22963 ( .A(n14687), .B(n14688), .Z(n14579) );
  NAND U22964 ( .A(n14689), .B(n14690), .Z(n14688) );
  NAND U22965 ( .A(n14691), .B(n14692), .Z(n14687) );
  AND U22966 ( .A(n14693), .B(n14694), .Z(n14581) );
  XOR U22967 ( .A(n14661), .B(n14660), .Z(N64089) );
  XNOR U22968 ( .A(n14678), .B(n14679), .Z(n14660) );
  XNOR U22969 ( .A(n14693), .B(n14694), .Z(n14679) );
  XOR U22970 ( .A(n14690), .B(n14689), .Z(n14694) );
  XOR U22971 ( .A(y[6468]), .B(x[6468]), .Z(n14689) );
  XOR U22972 ( .A(n14692), .B(n14691), .Z(n14690) );
  XOR U22973 ( .A(y[6470]), .B(x[6470]), .Z(n14691) );
  XOR U22974 ( .A(y[6469]), .B(x[6469]), .Z(n14692) );
  XOR U22975 ( .A(n14684), .B(n14683), .Z(n14693) );
  XOR U22976 ( .A(n14686), .B(n14685), .Z(n14683) );
  XOR U22977 ( .A(y[6467]), .B(x[6467]), .Z(n14685) );
  XOR U22978 ( .A(y[6466]), .B(x[6466]), .Z(n14686) );
  XOR U22979 ( .A(y[6465]), .B(x[6465]), .Z(n14684) );
  XNOR U22980 ( .A(n14677), .B(n14676), .Z(n14678) );
  XNOR U22981 ( .A(n14673), .B(n14672), .Z(n14676) );
  XOR U22982 ( .A(n14675), .B(n14674), .Z(n14672) );
  XOR U22983 ( .A(y[6464]), .B(x[6464]), .Z(n14674) );
  XOR U22984 ( .A(y[6463]), .B(x[6463]), .Z(n14675) );
  XOR U22985 ( .A(y[6462]), .B(x[6462]), .Z(n14673) );
  XOR U22986 ( .A(n14667), .B(n14666), .Z(n14677) );
  XOR U22987 ( .A(n14669), .B(n14668), .Z(n14666) );
  XOR U22988 ( .A(y[6461]), .B(x[6461]), .Z(n14668) );
  XOR U22989 ( .A(y[6460]), .B(x[6460]), .Z(n14669) );
  XOR U22990 ( .A(y[6459]), .B(x[6459]), .Z(n14667) );
  XNOR U22991 ( .A(n14643), .B(n14644), .Z(n14661) );
  XNOR U22992 ( .A(n14658), .B(n14659), .Z(n14644) );
  XOR U22993 ( .A(n14655), .B(n14654), .Z(n14659) );
  XOR U22994 ( .A(y[6456]), .B(x[6456]), .Z(n14654) );
  XOR U22995 ( .A(n14657), .B(n14656), .Z(n14655) );
  XOR U22996 ( .A(y[6458]), .B(x[6458]), .Z(n14656) );
  XOR U22997 ( .A(y[6457]), .B(x[6457]), .Z(n14657) );
  XOR U22998 ( .A(n14649), .B(n14648), .Z(n14658) );
  XOR U22999 ( .A(n14651), .B(n14650), .Z(n14648) );
  XOR U23000 ( .A(y[6455]), .B(x[6455]), .Z(n14650) );
  XOR U23001 ( .A(y[6454]), .B(x[6454]), .Z(n14651) );
  XOR U23002 ( .A(y[6453]), .B(x[6453]), .Z(n14649) );
  XNOR U23003 ( .A(n14642), .B(n14641), .Z(n14643) );
  XNOR U23004 ( .A(n14638), .B(n14637), .Z(n14641) );
  XOR U23005 ( .A(n14640), .B(n14639), .Z(n14637) );
  XOR U23006 ( .A(y[6452]), .B(x[6452]), .Z(n14639) );
  XOR U23007 ( .A(y[6451]), .B(x[6451]), .Z(n14640) );
  XOR U23008 ( .A(y[6450]), .B(x[6450]), .Z(n14638) );
  XOR U23009 ( .A(n14632), .B(n14631), .Z(n14642) );
  XOR U23010 ( .A(n14634), .B(n14633), .Z(n14631) );
  XOR U23011 ( .A(y[6449]), .B(x[6449]), .Z(n14633) );
  XOR U23012 ( .A(y[6448]), .B(x[6448]), .Z(n14634) );
  XOR U23013 ( .A(y[6447]), .B(x[6447]), .Z(n14632) );
  NAND U23014 ( .A(n14695), .B(n14696), .Z(N64080) );
  NAND U23015 ( .A(n14697), .B(n14698), .Z(n14696) );
  NANDN U23016 ( .A(n14699), .B(n14700), .Z(n14698) );
  NANDN U23017 ( .A(n14700), .B(n14699), .Z(n14695) );
  XOR U23018 ( .A(n14699), .B(n14701), .Z(N64079) );
  XNOR U23019 ( .A(n14697), .B(n14700), .Z(n14701) );
  NAND U23020 ( .A(n14702), .B(n14703), .Z(n14700) );
  NAND U23021 ( .A(n14704), .B(n14705), .Z(n14703) );
  NANDN U23022 ( .A(n14706), .B(n14707), .Z(n14705) );
  NANDN U23023 ( .A(n14707), .B(n14706), .Z(n14702) );
  AND U23024 ( .A(n14708), .B(n14709), .Z(n14697) );
  NAND U23025 ( .A(n14710), .B(n14711), .Z(n14709) );
  NANDN U23026 ( .A(n14712), .B(n14713), .Z(n14711) );
  NANDN U23027 ( .A(n14713), .B(n14712), .Z(n14708) );
  IV U23028 ( .A(n14714), .Z(n14713) );
  AND U23029 ( .A(n14715), .B(n14716), .Z(n14699) );
  NAND U23030 ( .A(n14717), .B(n14718), .Z(n14716) );
  NANDN U23031 ( .A(n14719), .B(n14720), .Z(n14718) );
  NANDN U23032 ( .A(n14720), .B(n14719), .Z(n14715) );
  XOR U23033 ( .A(n14712), .B(n14721), .Z(N64078) );
  XNOR U23034 ( .A(n14710), .B(n14714), .Z(n14721) );
  XOR U23035 ( .A(n14707), .B(n14722), .Z(n14714) );
  XNOR U23036 ( .A(n14704), .B(n14706), .Z(n14722) );
  AND U23037 ( .A(n14723), .B(n14724), .Z(n14706) );
  NANDN U23038 ( .A(n14725), .B(n14726), .Z(n14724) );
  OR U23039 ( .A(n14727), .B(n14728), .Z(n14726) );
  IV U23040 ( .A(n14729), .Z(n14728) );
  NANDN U23041 ( .A(n14729), .B(n14727), .Z(n14723) );
  AND U23042 ( .A(n14730), .B(n14731), .Z(n14704) );
  NAND U23043 ( .A(n14732), .B(n14733), .Z(n14731) );
  NANDN U23044 ( .A(n14734), .B(n14735), .Z(n14733) );
  NANDN U23045 ( .A(n14735), .B(n14734), .Z(n14730) );
  IV U23046 ( .A(n14736), .Z(n14735) );
  NAND U23047 ( .A(n14737), .B(n14738), .Z(n14707) );
  NANDN U23048 ( .A(n14739), .B(n14740), .Z(n14738) );
  NANDN U23049 ( .A(n14741), .B(n14742), .Z(n14740) );
  NANDN U23050 ( .A(n14742), .B(n14741), .Z(n14737) );
  IV U23051 ( .A(n14743), .Z(n14741) );
  AND U23052 ( .A(n14744), .B(n14745), .Z(n14710) );
  NAND U23053 ( .A(n14746), .B(n14747), .Z(n14745) );
  NANDN U23054 ( .A(n14748), .B(n14749), .Z(n14747) );
  NANDN U23055 ( .A(n14749), .B(n14748), .Z(n14744) );
  XOR U23056 ( .A(n14720), .B(n14750), .Z(n14712) );
  XNOR U23057 ( .A(n14717), .B(n14719), .Z(n14750) );
  AND U23058 ( .A(n14751), .B(n14752), .Z(n14719) );
  NANDN U23059 ( .A(n14753), .B(n14754), .Z(n14752) );
  OR U23060 ( .A(n14755), .B(n14756), .Z(n14754) );
  IV U23061 ( .A(n14757), .Z(n14756) );
  NANDN U23062 ( .A(n14757), .B(n14755), .Z(n14751) );
  AND U23063 ( .A(n14758), .B(n14759), .Z(n14717) );
  NAND U23064 ( .A(n14760), .B(n14761), .Z(n14759) );
  NANDN U23065 ( .A(n14762), .B(n14763), .Z(n14761) );
  NANDN U23066 ( .A(n14763), .B(n14762), .Z(n14758) );
  IV U23067 ( .A(n14764), .Z(n14763) );
  NAND U23068 ( .A(n14765), .B(n14766), .Z(n14720) );
  NANDN U23069 ( .A(n14767), .B(n14768), .Z(n14766) );
  NANDN U23070 ( .A(n14769), .B(n14770), .Z(n14768) );
  NANDN U23071 ( .A(n14770), .B(n14769), .Z(n14765) );
  IV U23072 ( .A(n14771), .Z(n14769) );
  XOR U23073 ( .A(n14746), .B(n14772), .Z(N64077) );
  XNOR U23074 ( .A(n14749), .B(n14748), .Z(n14772) );
  XNOR U23075 ( .A(n14760), .B(n14773), .Z(n14748) );
  XNOR U23076 ( .A(n14764), .B(n14762), .Z(n14773) );
  XOR U23077 ( .A(n14770), .B(n14774), .Z(n14762) );
  XNOR U23078 ( .A(n14767), .B(n14771), .Z(n14774) );
  AND U23079 ( .A(n14775), .B(n14776), .Z(n14771) );
  NAND U23080 ( .A(n14777), .B(n14778), .Z(n14776) );
  NAND U23081 ( .A(n14779), .B(n14780), .Z(n14775) );
  AND U23082 ( .A(n14781), .B(n14782), .Z(n14767) );
  NAND U23083 ( .A(n14783), .B(n14784), .Z(n14782) );
  NAND U23084 ( .A(n14785), .B(n14786), .Z(n14781) );
  NANDN U23085 ( .A(n14787), .B(n14788), .Z(n14770) );
  ANDN U23086 ( .B(n14789), .A(n14790), .Z(n14764) );
  XNOR U23087 ( .A(n14755), .B(n14791), .Z(n14760) );
  XNOR U23088 ( .A(n14753), .B(n14757), .Z(n14791) );
  AND U23089 ( .A(n14792), .B(n14793), .Z(n14757) );
  NAND U23090 ( .A(n14794), .B(n14795), .Z(n14793) );
  NAND U23091 ( .A(n14796), .B(n14797), .Z(n14792) );
  AND U23092 ( .A(n14798), .B(n14799), .Z(n14753) );
  NAND U23093 ( .A(n14800), .B(n14801), .Z(n14799) );
  NAND U23094 ( .A(n14802), .B(n14803), .Z(n14798) );
  AND U23095 ( .A(n14804), .B(n14805), .Z(n14755) );
  NAND U23096 ( .A(n14806), .B(n14807), .Z(n14749) );
  XNOR U23097 ( .A(n14732), .B(n14808), .Z(n14746) );
  XNOR U23098 ( .A(n14736), .B(n14734), .Z(n14808) );
  XOR U23099 ( .A(n14742), .B(n14809), .Z(n14734) );
  XNOR U23100 ( .A(n14739), .B(n14743), .Z(n14809) );
  AND U23101 ( .A(n14810), .B(n14811), .Z(n14743) );
  NAND U23102 ( .A(n14812), .B(n14813), .Z(n14811) );
  NAND U23103 ( .A(n14814), .B(n14815), .Z(n14810) );
  AND U23104 ( .A(n14816), .B(n14817), .Z(n14739) );
  NAND U23105 ( .A(n14818), .B(n14819), .Z(n14817) );
  NAND U23106 ( .A(n14820), .B(n14821), .Z(n14816) );
  NANDN U23107 ( .A(n14822), .B(n14823), .Z(n14742) );
  ANDN U23108 ( .B(n14824), .A(n14825), .Z(n14736) );
  XNOR U23109 ( .A(n14727), .B(n14826), .Z(n14732) );
  XNOR U23110 ( .A(n14725), .B(n14729), .Z(n14826) );
  AND U23111 ( .A(n14827), .B(n14828), .Z(n14729) );
  NAND U23112 ( .A(n14829), .B(n14830), .Z(n14828) );
  NAND U23113 ( .A(n14831), .B(n14832), .Z(n14827) );
  AND U23114 ( .A(n14833), .B(n14834), .Z(n14725) );
  NAND U23115 ( .A(n14835), .B(n14836), .Z(n14834) );
  NAND U23116 ( .A(n14837), .B(n14838), .Z(n14833) );
  AND U23117 ( .A(n14839), .B(n14840), .Z(n14727) );
  XOR U23118 ( .A(n14807), .B(n14806), .Z(N64076) );
  XNOR U23119 ( .A(n14824), .B(n14825), .Z(n14806) );
  XNOR U23120 ( .A(n14839), .B(n14840), .Z(n14825) );
  XOR U23121 ( .A(n14836), .B(n14835), .Z(n14840) );
  XOR U23122 ( .A(y[6444]), .B(x[6444]), .Z(n14835) );
  XOR U23123 ( .A(n14838), .B(n14837), .Z(n14836) );
  XOR U23124 ( .A(y[6446]), .B(x[6446]), .Z(n14837) );
  XOR U23125 ( .A(y[6445]), .B(x[6445]), .Z(n14838) );
  XOR U23126 ( .A(n14830), .B(n14829), .Z(n14839) );
  XOR U23127 ( .A(n14832), .B(n14831), .Z(n14829) );
  XOR U23128 ( .A(y[6443]), .B(x[6443]), .Z(n14831) );
  XOR U23129 ( .A(y[6442]), .B(x[6442]), .Z(n14832) );
  XOR U23130 ( .A(y[6441]), .B(x[6441]), .Z(n14830) );
  XNOR U23131 ( .A(n14823), .B(n14822), .Z(n14824) );
  XNOR U23132 ( .A(n14819), .B(n14818), .Z(n14822) );
  XOR U23133 ( .A(n14821), .B(n14820), .Z(n14818) );
  XOR U23134 ( .A(y[6440]), .B(x[6440]), .Z(n14820) );
  XOR U23135 ( .A(y[6439]), .B(x[6439]), .Z(n14821) );
  XOR U23136 ( .A(y[6438]), .B(x[6438]), .Z(n14819) );
  XOR U23137 ( .A(n14813), .B(n14812), .Z(n14823) );
  XOR U23138 ( .A(n14815), .B(n14814), .Z(n14812) );
  XOR U23139 ( .A(y[6437]), .B(x[6437]), .Z(n14814) );
  XOR U23140 ( .A(y[6436]), .B(x[6436]), .Z(n14815) );
  XOR U23141 ( .A(y[6435]), .B(x[6435]), .Z(n14813) );
  XNOR U23142 ( .A(n14789), .B(n14790), .Z(n14807) );
  XNOR U23143 ( .A(n14804), .B(n14805), .Z(n14790) );
  XOR U23144 ( .A(n14801), .B(n14800), .Z(n14805) );
  XOR U23145 ( .A(y[6432]), .B(x[6432]), .Z(n14800) );
  XOR U23146 ( .A(n14803), .B(n14802), .Z(n14801) );
  XOR U23147 ( .A(y[6434]), .B(x[6434]), .Z(n14802) );
  XOR U23148 ( .A(y[6433]), .B(x[6433]), .Z(n14803) );
  XOR U23149 ( .A(n14795), .B(n14794), .Z(n14804) );
  XOR U23150 ( .A(n14797), .B(n14796), .Z(n14794) );
  XOR U23151 ( .A(y[6431]), .B(x[6431]), .Z(n14796) );
  XOR U23152 ( .A(y[6430]), .B(x[6430]), .Z(n14797) );
  XOR U23153 ( .A(y[6429]), .B(x[6429]), .Z(n14795) );
  XNOR U23154 ( .A(n14788), .B(n14787), .Z(n14789) );
  XNOR U23155 ( .A(n14784), .B(n14783), .Z(n14787) );
  XOR U23156 ( .A(n14786), .B(n14785), .Z(n14783) );
  XOR U23157 ( .A(y[6428]), .B(x[6428]), .Z(n14785) );
  XOR U23158 ( .A(y[6427]), .B(x[6427]), .Z(n14786) );
  XOR U23159 ( .A(y[6426]), .B(x[6426]), .Z(n14784) );
  XOR U23160 ( .A(n14778), .B(n14777), .Z(n14788) );
  XOR U23161 ( .A(n14780), .B(n14779), .Z(n14777) );
  XOR U23162 ( .A(y[6425]), .B(x[6425]), .Z(n14779) );
  XOR U23163 ( .A(y[6424]), .B(x[6424]), .Z(n14780) );
  XOR U23164 ( .A(y[6423]), .B(x[6423]), .Z(n14778) );
  NAND U23165 ( .A(n14841), .B(n14842), .Z(N64067) );
  NAND U23166 ( .A(n14843), .B(n14844), .Z(n14842) );
  NANDN U23167 ( .A(n14845), .B(n14846), .Z(n14844) );
  NANDN U23168 ( .A(n14846), .B(n14845), .Z(n14841) );
  XOR U23169 ( .A(n14845), .B(n14847), .Z(N64066) );
  XNOR U23170 ( .A(n14843), .B(n14846), .Z(n14847) );
  NAND U23171 ( .A(n14848), .B(n14849), .Z(n14846) );
  NAND U23172 ( .A(n14850), .B(n14851), .Z(n14849) );
  NANDN U23173 ( .A(n14852), .B(n14853), .Z(n14851) );
  NANDN U23174 ( .A(n14853), .B(n14852), .Z(n14848) );
  AND U23175 ( .A(n14854), .B(n14855), .Z(n14843) );
  NAND U23176 ( .A(n14856), .B(n14857), .Z(n14855) );
  NANDN U23177 ( .A(n14858), .B(n14859), .Z(n14857) );
  NANDN U23178 ( .A(n14859), .B(n14858), .Z(n14854) );
  IV U23179 ( .A(n14860), .Z(n14859) );
  AND U23180 ( .A(n14861), .B(n14862), .Z(n14845) );
  NAND U23181 ( .A(n14863), .B(n14864), .Z(n14862) );
  NANDN U23182 ( .A(n14865), .B(n14866), .Z(n14864) );
  NANDN U23183 ( .A(n14866), .B(n14865), .Z(n14861) );
  XOR U23184 ( .A(n14858), .B(n14867), .Z(N64065) );
  XNOR U23185 ( .A(n14856), .B(n14860), .Z(n14867) );
  XOR U23186 ( .A(n14853), .B(n14868), .Z(n14860) );
  XNOR U23187 ( .A(n14850), .B(n14852), .Z(n14868) );
  AND U23188 ( .A(n14869), .B(n14870), .Z(n14852) );
  NANDN U23189 ( .A(n14871), .B(n14872), .Z(n14870) );
  OR U23190 ( .A(n14873), .B(n14874), .Z(n14872) );
  IV U23191 ( .A(n14875), .Z(n14874) );
  NANDN U23192 ( .A(n14875), .B(n14873), .Z(n14869) );
  AND U23193 ( .A(n14876), .B(n14877), .Z(n14850) );
  NAND U23194 ( .A(n14878), .B(n14879), .Z(n14877) );
  NANDN U23195 ( .A(n14880), .B(n14881), .Z(n14879) );
  NANDN U23196 ( .A(n14881), .B(n14880), .Z(n14876) );
  IV U23197 ( .A(n14882), .Z(n14881) );
  NAND U23198 ( .A(n14883), .B(n14884), .Z(n14853) );
  NANDN U23199 ( .A(n14885), .B(n14886), .Z(n14884) );
  NANDN U23200 ( .A(n14887), .B(n14888), .Z(n14886) );
  NANDN U23201 ( .A(n14888), .B(n14887), .Z(n14883) );
  IV U23202 ( .A(n14889), .Z(n14887) );
  AND U23203 ( .A(n14890), .B(n14891), .Z(n14856) );
  NAND U23204 ( .A(n14892), .B(n14893), .Z(n14891) );
  NANDN U23205 ( .A(n14894), .B(n14895), .Z(n14893) );
  NANDN U23206 ( .A(n14895), .B(n14894), .Z(n14890) );
  XOR U23207 ( .A(n14866), .B(n14896), .Z(n14858) );
  XNOR U23208 ( .A(n14863), .B(n14865), .Z(n14896) );
  AND U23209 ( .A(n14897), .B(n14898), .Z(n14865) );
  NANDN U23210 ( .A(n14899), .B(n14900), .Z(n14898) );
  OR U23211 ( .A(n14901), .B(n14902), .Z(n14900) );
  IV U23212 ( .A(n14903), .Z(n14902) );
  NANDN U23213 ( .A(n14903), .B(n14901), .Z(n14897) );
  AND U23214 ( .A(n14904), .B(n14905), .Z(n14863) );
  NAND U23215 ( .A(n14906), .B(n14907), .Z(n14905) );
  NANDN U23216 ( .A(n14908), .B(n14909), .Z(n14907) );
  NANDN U23217 ( .A(n14909), .B(n14908), .Z(n14904) );
  IV U23218 ( .A(n14910), .Z(n14909) );
  NAND U23219 ( .A(n14911), .B(n14912), .Z(n14866) );
  NANDN U23220 ( .A(n14913), .B(n14914), .Z(n14912) );
  NANDN U23221 ( .A(n14915), .B(n14916), .Z(n14914) );
  NANDN U23222 ( .A(n14916), .B(n14915), .Z(n14911) );
  IV U23223 ( .A(n14917), .Z(n14915) );
  XOR U23224 ( .A(n14892), .B(n14918), .Z(N64064) );
  XNOR U23225 ( .A(n14895), .B(n14894), .Z(n14918) );
  XNOR U23226 ( .A(n14906), .B(n14919), .Z(n14894) );
  XNOR U23227 ( .A(n14910), .B(n14908), .Z(n14919) );
  XOR U23228 ( .A(n14916), .B(n14920), .Z(n14908) );
  XNOR U23229 ( .A(n14913), .B(n14917), .Z(n14920) );
  AND U23230 ( .A(n14921), .B(n14922), .Z(n14917) );
  NAND U23231 ( .A(n14923), .B(n14924), .Z(n14922) );
  NAND U23232 ( .A(n14925), .B(n14926), .Z(n14921) );
  AND U23233 ( .A(n14927), .B(n14928), .Z(n14913) );
  NAND U23234 ( .A(n14929), .B(n14930), .Z(n14928) );
  NAND U23235 ( .A(n14931), .B(n14932), .Z(n14927) );
  NANDN U23236 ( .A(n14933), .B(n14934), .Z(n14916) );
  ANDN U23237 ( .B(n14935), .A(n14936), .Z(n14910) );
  XNOR U23238 ( .A(n14901), .B(n14937), .Z(n14906) );
  XNOR U23239 ( .A(n14899), .B(n14903), .Z(n14937) );
  AND U23240 ( .A(n14938), .B(n14939), .Z(n14903) );
  NAND U23241 ( .A(n14940), .B(n14941), .Z(n14939) );
  NAND U23242 ( .A(n14942), .B(n14943), .Z(n14938) );
  AND U23243 ( .A(n14944), .B(n14945), .Z(n14899) );
  NAND U23244 ( .A(n14946), .B(n14947), .Z(n14945) );
  NAND U23245 ( .A(n14948), .B(n14949), .Z(n14944) );
  AND U23246 ( .A(n14950), .B(n14951), .Z(n14901) );
  NAND U23247 ( .A(n14952), .B(n14953), .Z(n14895) );
  XNOR U23248 ( .A(n14878), .B(n14954), .Z(n14892) );
  XNOR U23249 ( .A(n14882), .B(n14880), .Z(n14954) );
  XOR U23250 ( .A(n14888), .B(n14955), .Z(n14880) );
  XNOR U23251 ( .A(n14885), .B(n14889), .Z(n14955) );
  AND U23252 ( .A(n14956), .B(n14957), .Z(n14889) );
  NAND U23253 ( .A(n14958), .B(n14959), .Z(n14957) );
  NAND U23254 ( .A(n14960), .B(n14961), .Z(n14956) );
  AND U23255 ( .A(n14962), .B(n14963), .Z(n14885) );
  NAND U23256 ( .A(n14964), .B(n14965), .Z(n14963) );
  NAND U23257 ( .A(n14966), .B(n14967), .Z(n14962) );
  NANDN U23258 ( .A(n14968), .B(n14969), .Z(n14888) );
  ANDN U23259 ( .B(n14970), .A(n14971), .Z(n14882) );
  XNOR U23260 ( .A(n14873), .B(n14972), .Z(n14878) );
  XNOR U23261 ( .A(n14871), .B(n14875), .Z(n14972) );
  AND U23262 ( .A(n14973), .B(n14974), .Z(n14875) );
  NAND U23263 ( .A(n14975), .B(n14976), .Z(n14974) );
  NAND U23264 ( .A(n14977), .B(n14978), .Z(n14973) );
  AND U23265 ( .A(n14979), .B(n14980), .Z(n14871) );
  NAND U23266 ( .A(n14981), .B(n14982), .Z(n14980) );
  NAND U23267 ( .A(n14983), .B(n14984), .Z(n14979) );
  AND U23268 ( .A(n14985), .B(n14986), .Z(n14873) );
  XOR U23269 ( .A(n14953), .B(n14952), .Z(N64063) );
  XNOR U23270 ( .A(n14970), .B(n14971), .Z(n14952) );
  XNOR U23271 ( .A(n14985), .B(n14986), .Z(n14971) );
  XOR U23272 ( .A(n14982), .B(n14981), .Z(n14986) );
  XOR U23273 ( .A(y[6420]), .B(x[6420]), .Z(n14981) );
  XOR U23274 ( .A(n14984), .B(n14983), .Z(n14982) );
  XOR U23275 ( .A(y[6422]), .B(x[6422]), .Z(n14983) );
  XOR U23276 ( .A(y[6421]), .B(x[6421]), .Z(n14984) );
  XOR U23277 ( .A(n14976), .B(n14975), .Z(n14985) );
  XOR U23278 ( .A(n14978), .B(n14977), .Z(n14975) );
  XOR U23279 ( .A(y[6419]), .B(x[6419]), .Z(n14977) );
  XOR U23280 ( .A(y[6418]), .B(x[6418]), .Z(n14978) );
  XOR U23281 ( .A(y[6417]), .B(x[6417]), .Z(n14976) );
  XNOR U23282 ( .A(n14969), .B(n14968), .Z(n14970) );
  XNOR U23283 ( .A(n14965), .B(n14964), .Z(n14968) );
  XOR U23284 ( .A(n14967), .B(n14966), .Z(n14964) );
  XOR U23285 ( .A(y[6416]), .B(x[6416]), .Z(n14966) );
  XOR U23286 ( .A(y[6415]), .B(x[6415]), .Z(n14967) );
  XOR U23287 ( .A(y[6414]), .B(x[6414]), .Z(n14965) );
  XOR U23288 ( .A(n14959), .B(n14958), .Z(n14969) );
  XOR U23289 ( .A(n14961), .B(n14960), .Z(n14958) );
  XOR U23290 ( .A(y[6413]), .B(x[6413]), .Z(n14960) );
  XOR U23291 ( .A(y[6412]), .B(x[6412]), .Z(n14961) );
  XOR U23292 ( .A(y[6411]), .B(x[6411]), .Z(n14959) );
  XNOR U23293 ( .A(n14935), .B(n14936), .Z(n14953) );
  XNOR U23294 ( .A(n14950), .B(n14951), .Z(n14936) );
  XOR U23295 ( .A(n14947), .B(n14946), .Z(n14951) );
  XOR U23296 ( .A(y[6408]), .B(x[6408]), .Z(n14946) );
  XOR U23297 ( .A(n14949), .B(n14948), .Z(n14947) );
  XOR U23298 ( .A(y[6410]), .B(x[6410]), .Z(n14948) );
  XOR U23299 ( .A(y[6409]), .B(x[6409]), .Z(n14949) );
  XOR U23300 ( .A(n14941), .B(n14940), .Z(n14950) );
  XOR U23301 ( .A(n14943), .B(n14942), .Z(n14940) );
  XOR U23302 ( .A(y[6407]), .B(x[6407]), .Z(n14942) );
  XOR U23303 ( .A(y[6406]), .B(x[6406]), .Z(n14943) );
  XOR U23304 ( .A(y[6405]), .B(x[6405]), .Z(n14941) );
  XNOR U23305 ( .A(n14934), .B(n14933), .Z(n14935) );
  XNOR U23306 ( .A(n14930), .B(n14929), .Z(n14933) );
  XOR U23307 ( .A(n14932), .B(n14931), .Z(n14929) );
  XOR U23308 ( .A(y[6404]), .B(x[6404]), .Z(n14931) );
  XOR U23309 ( .A(y[6403]), .B(x[6403]), .Z(n14932) );
  XOR U23310 ( .A(y[6402]), .B(x[6402]), .Z(n14930) );
  XOR U23311 ( .A(n14924), .B(n14923), .Z(n14934) );
  XOR U23312 ( .A(n14926), .B(n14925), .Z(n14923) );
  XOR U23313 ( .A(y[6401]), .B(x[6401]), .Z(n14925) );
  XOR U23314 ( .A(y[6400]), .B(x[6400]), .Z(n14926) );
  XOR U23315 ( .A(y[6399]), .B(x[6399]), .Z(n14924) );
  NAND U23316 ( .A(n14987), .B(n14988), .Z(N64054) );
  NAND U23317 ( .A(n14989), .B(n14990), .Z(n14988) );
  NANDN U23318 ( .A(n14991), .B(n14992), .Z(n14990) );
  NANDN U23319 ( .A(n14992), .B(n14991), .Z(n14987) );
  XOR U23320 ( .A(n14991), .B(n14993), .Z(N64053) );
  XNOR U23321 ( .A(n14989), .B(n14992), .Z(n14993) );
  NAND U23322 ( .A(n14994), .B(n14995), .Z(n14992) );
  NAND U23323 ( .A(n14996), .B(n14997), .Z(n14995) );
  NANDN U23324 ( .A(n14998), .B(n14999), .Z(n14997) );
  NANDN U23325 ( .A(n14999), .B(n14998), .Z(n14994) );
  AND U23326 ( .A(n15000), .B(n15001), .Z(n14989) );
  NAND U23327 ( .A(n15002), .B(n15003), .Z(n15001) );
  NANDN U23328 ( .A(n15004), .B(n15005), .Z(n15003) );
  NANDN U23329 ( .A(n15005), .B(n15004), .Z(n15000) );
  IV U23330 ( .A(n15006), .Z(n15005) );
  AND U23331 ( .A(n15007), .B(n15008), .Z(n14991) );
  NAND U23332 ( .A(n15009), .B(n15010), .Z(n15008) );
  NANDN U23333 ( .A(n15011), .B(n15012), .Z(n15010) );
  NANDN U23334 ( .A(n15012), .B(n15011), .Z(n15007) );
  XOR U23335 ( .A(n15004), .B(n15013), .Z(N64052) );
  XNOR U23336 ( .A(n15002), .B(n15006), .Z(n15013) );
  XOR U23337 ( .A(n14999), .B(n15014), .Z(n15006) );
  XNOR U23338 ( .A(n14996), .B(n14998), .Z(n15014) );
  AND U23339 ( .A(n15015), .B(n15016), .Z(n14998) );
  NANDN U23340 ( .A(n15017), .B(n15018), .Z(n15016) );
  OR U23341 ( .A(n15019), .B(n15020), .Z(n15018) );
  IV U23342 ( .A(n15021), .Z(n15020) );
  NANDN U23343 ( .A(n15021), .B(n15019), .Z(n15015) );
  AND U23344 ( .A(n15022), .B(n15023), .Z(n14996) );
  NAND U23345 ( .A(n15024), .B(n15025), .Z(n15023) );
  NANDN U23346 ( .A(n15026), .B(n15027), .Z(n15025) );
  NANDN U23347 ( .A(n15027), .B(n15026), .Z(n15022) );
  IV U23348 ( .A(n15028), .Z(n15027) );
  NAND U23349 ( .A(n15029), .B(n15030), .Z(n14999) );
  NANDN U23350 ( .A(n15031), .B(n15032), .Z(n15030) );
  NANDN U23351 ( .A(n15033), .B(n15034), .Z(n15032) );
  NANDN U23352 ( .A(n15034), .B(n15033), .Z(n15029) );
  IV U23353 ( .A(n15035), .Z(n15033) );
  AND U23354 ( .A(n15036), .B(n15037), .Z(n15002) );
  NAND U23355 ( .A(n15038), .B(n15039), .Z(n15037) );
  NANDN U23356 ( .A(n15040), .B(n15041), .Z(n15039) );
  NANDN U23357 ( .A(n15041), .B(n15040), .Z(n15036) );
  XOR U23358 ( .A(n15012), .B(n15042), .Z(n15004) );
  XNOR U23359 ( .A(n15009), .B(n15011), .Z(n15042) );
  AND U23360 ( .A(n15043), .B(n15044), .Z(n15011) );
  NANDN U23361 ( .A(n15045), .B(n15046), .Z(n15044) );
  OR U23362 ( .A(n15047), .B(n15048), .Z(n15046) );
  IV U23363 ( .A(n15049), .Z(n15048) );
  NANDN U23364 ( .A(n15049), .B(n15047), .Z(n15043) );
  AND U23365 ( .A(n15050), .B(n15051), .Z(n15009) );
  NAND U23366 ( .A(n15052), .B(n15053), .Z(n15051) );
  NANDN U23367 ( .A(n15054), .B(n15055), .Z(n15053) );
  NANDN U23368 ( .A(n15055), .B(n15054), .Z(n15050) );
  IV U23369 ( .A(n15056), .Z(n15055) );
  NAND U23370 ( .A(n15057), .B(n15058), .Z(n15012) );
  NANDN U23371 ( .A(n15059), .B(n15060), .Z(n15058) );
  NANDN U23372 ( .A(n15061), .B(n15062), .Z(n15060) );
  NANDN U23373 ( .A(n15062), .B(n15061), .Z(n15057) );
  IV U23374 ( .A(n15063), .Z(n15061) );
  XOR U23375 ( .A(n15038), .B(n15064), .Z(N64051) );
  XNOR U23376 ( .A(n15041), .B(n15040), .Z(n15064) );
  XNOR U23377 ( .A(n15052), .B(n15065), .Z(n15040) );
  XNOR U23378 ( .A(n15056), .B(n15054), .Z(n15065) );
  XOR U23379 ( .A(n15062), .B(n15066), .Z(n15054) );
  XNOR U23380 ( .A(n15059), .B(n15063), .Z(n15066) );
  AND U23381 ( .A(n15067), .B(n15068), .Z(n15063) );
  NAND U23382 ( .A(n15069), .B(n15070), .Z(n15068) );
  NAND U23383 ( .A(n15071), .B(n15072), .Z(n15067) );
  AND U23384 ( .A(n15073), .B(n15074), .Z(n15059) );
  NAND U23385 ( .A(n15075), .B(n15076), .Z(n15074) );
  NAND U23386 ( .A(n15077), .B(n15078), .Z(n15073) );
  NANDN U23387 ( .A(n15079), .B(n15080), .Z(n15062) );
  ANDN U23388 ( .B(n15081), .A(n15082), .Z(n15056) );
  XNOR U23389 ( .A(n15047), .B(n15083), .Z(n15052) );
  XNOR U23390 ( .A(n15045), .B(n15049), .Z(n15083) );
  AND U23391 ( .A(n15084), .B(n15085), .Z(n15049) );
  NAND U23392 ( .A(n15086), .B(n15087), .Z(n15085) );
  NAND U23393 ( .A(n15088), .B(n15089), .Z(n15084) );
  AND U23394 ( .A(n15090), .B(n15091), .Z(n15045) );
  NAND U23395 ( .A(n15092), .B(n15093), .Z(n15091) );
  NAND U23396 ( .A(n15094), .B(n15095), .Z(n15090) );
  AND U23397 ( .A(n15096), .B(n15097), .Z(n15047) );
  NAND U23398 ( .A(n15098), .B(n15099), .Z(n15041) );
  XNOR U23399 ( .A(n15024), .B(n15100), .Z(n15038) );
  XNOR U23400 ( .A(n15028), .B(n15026), .Z(n15100) );
  XOR U23401 ( .A(n15034), .B(n15101), .Z(n15026) );
  XNOR U23402 ( .A(n15031), .B(n15035), .Z(n15101) );
  AND U23403 ( .A(n15102), .B(n15103), .Z(n15035) );
  NAND U23404 ( .A(n15104), .B(n15105), .Z(n15103) );
  NAND U23405 ( .A(n15106), .B(n15107), .Z(n15102) );
  AND U23406 ( .A(n15108), .B(n15109), .Z(n15031) );
  NAND U23407 ( .A(n15110), .B(n15111), .Z(n15109) );
  NAND U23408 ( .A(n15112), .B(n15113), .Z(n15108) );
  NANDN U23409 ( .A(n15114), .B(n15115), .Z(n15034) );
  ANDN U23410 ( .B(n15116), .A(n15117), .Z(n15028) );
  XNOR U23411 ( .A(n15019), .B(n15118), .Z(n15024) );
  XNOR U23412 ( .A(n15017), .B(n15021), .Z(n15118) );
  AND U23413 ( .A(n15119), .B(n15120), .Z(n15021) );
  NAND U23414 ( .A(n15121), .B(n15122), .Z(n15120) );
  NAND U23415 ( .A(n15123), .B(n15124), .Z(n15119) );
  AND U23416 ( .A(n15125), .B(n15126), .Z(n15017) );
  NAND U23417 ( .A(n15127), .B(n15128), .Z(n15126) );
  NAND U23418 ( .A(n15129), .B(n15130), .Z(n15125) );
  AND U23419 ( .A(n15131), .B(n15132), .Z(n15019) );
  XOR U23420 ( .A(n15099), .B(n15098), .Z(N64050) );
  XNOR U23421 ( .A(n15116), .B(n15117), .Z(n15098) );
  XNOR U23422 ( .A(n15131), .B(n15132), .Z(n15117) );
  XOR U23423 ( .A(n15128), .B(n15127), .Z(n15132) );
  XOR U23424 ( .A(y[6396]), .B(x[6396]), .Z(n15127) );
  XOR U23425 ( .A(n15130), .B(n15129), .Z(n15128) );
  XOR U23426 ( .A(y[6398]), .B(x[6398]), .Z(n15129) );
  XOR U23427 ( .A(y[6397]), .B(x[6397]), .Z(n15130) );
  XOR U23428 ( .A(n15122), .B(n15121), .Z(n15131) );
  XOR U23429 ( .A(n15124), .B(n15123), .Z(n15121) );
  XOR U23430 ( .A(y[6395]), .B(x[6395]), .Z(n15123) );
  XOR U23431 ( .A(y[6394]), .B(x[6394]), .Z(n15124) );
  XOR U23432 ( .A(y[6393]), .B(x[6393]), .Z(n15122) );
  XNOR U23433 ( .A(n15115), .B(n15114), .Z(n15116) );
  XNOR U23434 ( .A(n15111), .B(n15110), .Z(n15114) );
  XOR U23435 ( .A(n15113), .B(n15112), .Z(n15110) );
  XOR U23436 ( .A(y[6392]), .B(x[6392]), .Z(n15112) );
  XOR U23437 ( .A(y[6391]), .B(x[6391]), .Z(n15113) );
  XOR U23438 ( .A(y[6390]), .B(x[6390]), .Z(n15111) );
  XOR U23439 ( .A(n15105), .B(n15104), .Z(n15115) );
  XOR U23440 ( .A(n15107), .B(n15106), .Z(n15104) );
  XOR U23441 ( .A(y[6389]), .B(x[6389]), .Z(n15106) );
  XOR U23442 ( .A(y[6388]), .B(x[6388]), .Z(n15107) );
  XOR U23443 ( .A(y[6387]), .B(x[6387]), .Z(n15105) );
  XNOR U23444 ( .A(n15081), .B(n15082), .Z(n15099) );
  XNOR U23445 ( .A(n15096), .B(n15097), .Z(n15082) );
  XOR U23446 ( .A(n15093), .B(n15092), .Z(n15097) );
  XOR U23447 ( .A(y[6384]), .B(x[6384]), .Z(n15092) );
  XOR U23448 ( .A(n15095), .B(n15094), .Z(n15093) );
  XOR U23449 ( .A(y[6386]), .B(x[6386]), .Z(n15094) );
  XOR U23450 ( .A(y[6385]), .B(x[6385]), .Z(n15095) );
  XOR U23451 ( .A(n15087), .B(n15086), .Z(n15096) );
  XOR U23452 ( .A(n15089), .B(n15088), .Z(n15086) );
  XOR U23453 ( .A(y[6383]), .B(x[6383]), .Z(n15088) );
  XOR U23454 ( .A(y[6382]), .B(x[6382]), .Z(n15089) );
  XOR U23455 ( .A(y[6381]), .B(x[6381]), .Z(n15087) );
  XNOR U23456 ( .A(n15080), .B(n15079), .Z(n15081) );
  XNOR U23457 ( .A(n15076), .B(n15075), .Z(n15079) );
  XOR U23458 ( .A(n15078), .B(n15077), .Z(n15075) );
  XOR U23459 ( .A(y[6380]), .B(x[6380]), .Z(n15077) );
  XOR U23460 ( .A(y[6379]), .B(x[6379]), .Z(n15078) );
  XOR U23461 ( .A(y[6378]), .B(x[6378]), .Z(n15076) );
  XOR U23462 ( .A(n15070), .B(n15069), .Z(n15080) );
  XOR U23463 ( .A(n15072), .B(n15071), .Z(n15069) );
  XOR U23464 ( .A(y[6377]), .B(x[6377]), .Z(n15071) );
  XOR U23465 ( .A(y[6376]), .B(x[6376]), .Z(n15072) );
  XOR U23466 ( .A(y[6375]), .B(x[6375]), .Z(n15070) );
  NAND U23467 ( .A(n15133), .B(n15134), .Z(N64041) );
  NAND U23468 ( .A(n15135), .B(n15136), .Z(n15134) );
  NANDN U23469 ( .A(n15137), .B(n15138), .Z(n15136) );
  NANDN U23470 ( .A(n15138), .B(n15137), .Z(n15133) );
  XOR U23471 ( .A(n15137), .B(n15139), .Z(N64040) );
  XNOR U23472 ( .A(n15135), .B(n15138), .Z(n15139) );
  NAND U23473 ( .A(n15140), .B(n15141), .Z(n15138) );
  NAND U23474 ( .A(n15142), .B(n15143), .Z(n15141) );
  NANDN U23475 ( .A(n15144), .B(n15145), .Z(n15143) );
  NANDN U23476 ( .A(n15145), .B(n15144), .Z(n15140) );
  AND U23477 ( .A(n15146), .B(n15147), .Z(n15135) );
  NAND U23478 ( .A(n15148), .B(n15149), .Z(n15147) );
  NANDN U23479 ( .A(n15150), .B(n15151), .Z(n15149) );
  NANDN U23480 ( .A(n15151), .B(n15150), .Z(n15146) );
  IV U23481 ( .A(n15152), .Z(n15151) );
  AND U23482 ( .A(n15153), .B(n15154), .Z(n15137) );
  NAND U23483 ( .A(n15155), .B(n15156), .Z(n15154) );
  NANDN U23484 ( .A(n15157), .B(n15158), .Z(n15156) );
  NANDN U23485 ( .A(n15158), .B(n15157), .Z(n15153) );
  XOR U23486 ( .A(n15150), .B(n15159), .Z(N64039) );
  XNOR U23487 ( .A(n15148), .B(n15152), .Z(n15159) );
  XOR U23488 ( .A(n15145), .B(n15160), .Z(n15152) );
  XNOR U23489 ( .A(n15142), .B(n15144), .Z(n15160) );
  AND U23490 ( .A(n15161), .B(n15162), .Z(n15144) );
  NANDN U23491 ( .A(n15163), .B(n15164), .Z(n15162) );
  OR U23492 ( .A(n15165), .B(n15166), .Z(n15164) );
  IV U23493 ( .A(n15167), .Z(n15166) );
  NANDN U23494 ( .A(n15167), .B(n15165), .Z(n15161) );
  AND U23495 ( .A(n15168), .B(n15169), .Z(n15142) );
  NAND U23496 ( .A(n15170), .B(n15171), .Z(n15169) );
  NANDN U23497 ( .A(n15172), .B(n15173), .Z(n15171) );
  NANDN U23498 ( .A(n15173), .B(n15172), .Z(n15168) );
  IV U23499 ( .A(n15174), .Z(n15173) );
  NAND U23500 ( .A(n15175), .B(n15176), .Z(n15145) );
  NANDN U23501 ( .A(n15177), .B(n15178), .Z(n15176) );
  NANDN U23502 ( .A(n15179), .B(n15180), .Z(n15178) );
  NANDN U23503 ( .A(n15180), .B(n15179), .Z(n15175) );
  IV U23504 ( .A(n15181), .Z(n15179) );
  AND U23505 ( .A(n15182), .B(n15183), .Z(n15148) );
  NAND U23506 ( .A(n15184), .B(n15185), .Z(n15183) );
  NANDN U23507 ( .A(n15186), .B(n15187), .Z(n15185) );
  NANDN U23508 ( .A(n15187), .B(n15186), .Z(n15182) );
  XOR U23509 ( .A(n15158), .B(n15188), .Z(n15150) );
  XNOR U23510 ( .A(n15155), .B(n15157), .Z(n15188) );
  AND U23511 ( .A(n15189), .B(n15190), .Z(n15157) );
  NANDN U23512 ( .A(n15191), .B(n15192), .Z(n15190) );
  OR U23513 ( .A(n15193), .B(n15194), .Z(n15192) );
  IV U23514 ( .A(n15195), .Z(n15194) );
  NANDN U23515 ( .A(n15195), .B(n15193), .Z(n15189) );
  AND U23516 ( .A(n15196), .B(n15197), .Z(n15155) );
  NAND U23517 ( .A(n15198), .B(n15199), .Z(n15197) );
  NANDN U23518 ( .A(n15200), .B(n15201), .Z(n15199) );
  NANDN U23519 ( .A(n15201), .B(n15200), .Z(n15196) );
  IV U23520 ( .A(n15202), .Z(n15201) );
  NAND U23521 ( .A(n15203), .B(n15204), .Z(n15158) );
  NANDN U23522 ( .A(n15205), .B(n15206), .Z(n15204) );
  NANDN U23523 ( .A(n15207), .B(n15208), .Z(n15206) );
  NANDN U23524 ( .A(n15208), .B(n15207), .Z(n15203) );
  IV U23525 ( .A(n15209), .Z(n15207) );
  XOR U23526 ( .A(n15184), .B(n15210), .Z(N64038) );
  XNOR U23527 ( .A(n15187), .B(n15186), .Z(n15210) );
  XNOR U23528 ( .A(n15198), .B(n15211), .Z(n15186) );
  XNOR U23529 ( .A(n15202), .B(n15200), .Z(n15211) );
  XOR U23530 ( .A(n15208), .B(n15212), .Z(n15200) );
  XNOR U23531 ( .A(n15205), .B(n15209), .Z(n15212) );
  AND U23532 ( .A(n15213), .B(n15214), .Z(n15209) );
  NAND U23533 ( .A(n15215), .B(n15216), .Z(n15214) );
  NAND U23534 ( .A(n15217), .B(n15218), .Z(n15213) );
  AND U23535 ( .A(n15219), .B(n15220), .Z(n15205) );
  NAND U23536 ( .A(n15221), .B(n15222), .Z(n15220) );
  NAND U23537 ( .A(n15223), .B(n15224), .Z(n15219) );
  NANDN U23538 ( .A(n15225), .B(n15226), .Z(n15208) );
  ANDN U23539 ( .B(n15227), .A(n15228), .Z(n15202) );
  XNOR U23540 ( .A(n15193), .B(n15229), .Z(n15198) );
  XNOR U23541 ( .A(n15191), .B(n15195), .Z(n15229) );
  AND U23542 ( .A(n15230), .B(n15231), .Z(n15195) );
  NAND U23543 ( .A(n15232), .B(n15233), .Z(n15231) );
  NAND U23544 ( .A(n15234), .B(n15235), .Z(n15230) );
  AND U23545 ( .A(n15236), .B(n15237), .Z(n15191) );
  NAND U23546 ( .A(n15238), .B(n15239), .Z(n15237) );
  NAND U23547 ( .A(n15240), .B(n15241), .Z(n15236) );
  AND U23548 ( .A(n15242), .B(n15243), .Z(n15193) );
  NAND U23549 ( .A(n15244), .B(n15245), .Z(n15187) );
  XNOR U23550 ( .A(n15170), .B(n15246), .Z(n15184) );
  XNOR U23551 ( .A(n15174), .B(n15172), .Z(n15246) );
  XOR U23552 ( .A(n15180), .B(n15247), .Z(n15172) );
  XNOR U23553 ( .A(n15177), .B(n15181), .Z(n15247) );
  AND U23554 ( .A(n15248), .B(n15249), .Z(n15181) );
  NAND U23555 ( .A(n15250), .B(n15251), .Z(n15249) );
  NAND U23556 ( .A(n15252), .B(n15253), .Z(n15248) );
  AND U23557 ( .A(n15254), .B(n15255), .Z(n15177) );
  NAND U23558 ( .A(n15256), .B(n15257), .Z(n15255) );
  NAND U23559 ( .A(n15258), .B(n15259), .Z(n15254) );
  NANDN U23560 ( .A(n15260), .B(n15261), .Z(n15180) );
  ANDN U23561 ( .B(n15262), .A(n15263), .Z(n15174) );
  XNOR U23562 ( .A(n15165), .B(n15264), .Z(n15170) );
  XNOR U23563 ( .A(n15163), .B(n15167), .Z(n15264) );
  AND U23564 ( .A(n15265), .B(n15266), .Z(n15167) );
  NAND U23565 ( .A(n15267), .B(n15268), .Z(n15266) );
  NAND U23566 ( .A(n15269), .B(n15270), .Z(n15265) );
  AND U23567 ( .A(n15271), .B(n15272), .Z(n15163) );
  NAND U23568 ( .A(n15273), .B(n15274), .Z(n15272) );
  NAND U23569 ( .A(n15275), .B(n15276), .Z(n15271) );
  AND U23570 ( .A(n15277), .B(n15278), .Z(n15165) );
  XOR U23571 ( .A(n15245), .B(n15244), .Z(N64037) );
  XNOR U23572 ( .A(n15262), .B(n15263), .Z(n15244) );
  XNOR U23573 ( .A(n15277), .B(n15278), .Z(n15263) );
  XOR U23574 ( .A(n15274), .B(n15273), .Z(n15278) );
  XOR U23575 ( .A(y[6372]), .B(x[6372]), .Z(n15273) );
  XOR U23576 ( .A(n15276), .B(n15275), .Z(n15274) );
  XOR U23577 ( .A(y[6374]), .B(x[6374]), .Z(n15275) );
  XOR U23578 ( .A(y[6373]), .B(x[6373]), .Z(n15276) );
  XOR U23579 ( .A(n15268), .B(n15267), .Z(n15277) );
  XOR U23580 ( .A(n15270), .B(n15269), .Z(n15267) );
  XOR U23581 ( .A(y[6371]), .B(x[6371]), .Z(n15269) );
  XOR U23582 ( .A(y[6370]), .B(x[6370]), .Z(n15270) );
  XOR U23583 ( .A(y[6369]), .B(x[6369]), .Z(n15268) );
  XNOR U23584 ( .A(n15261), .B(n15260), .Z(n15262) );
  XNOR U23585 ( .A(n15257), .B(n15256), .Z(n15260) );
  XOR U23586 ( .A(n15259), .B(n15258), .Z(n15256) );
  XOR U23587 ( .A(y[6368]), .B(x[6368]), .Z(n15258) );
  XOR U23588 ( .A(y[6367]), .B(x[6367]), .Z(n15259) );
  XOR U23589 ( .A(y[6366]), .B(x[6366]), .Z(n15257) );
  XOR U23590 ( .A(n15251), .B(n15250), .Z(n15261) );
  XOR U23591 ( .A(n15253), .B(n15252), .Z(n15250) );
  XOR U23592 ( .A(y[6365]), .B(x[6365]), .Z(n15252) );
  XOR U23593 ( .A(y[6364]), .B(x[6364]), .Z(n15253) );
  XOR U23594 ( .A(y[6363]), .B(x[6363]), .Z(n15251) );
  XNOR U23595 ( .A(n15227), .B(n15228), .Z(n15245) );
  XNOR U23596 ( .A(n15242), .B(n15243), .Z(n15228) );
  XOR U23597 ( .A(n15239), .B(n15238), .Z(n15243) );
  XOR U23598 ( .A(y[6360]), .B(x[6360]), .Z(n15238) );
  XOR U23599 ( .A(n15241), .B(n15240), .Z(n15239) );
  XOR U23600 ( .A(y[6362]), .B(x[6362]), .Z(n15240) );
  XOR U23601 ( .A(y[6361]), .B(x[6361]), .Z(n15241) );
  XOR U23602 ( .A(n15233), .B(n15232), .Z(n15242) );
  XOR U23603 ( .A(n15235), .B(n15234), .Z(n15232) );
  XOR U23604 ( .A(y[6359]), .B(x[6359]), .Z(n15234) );
  XOR U23605 ( .A(y[6358]), .B(x[6358]), .Z(n15235) );
  XOR U23606 ( .A(y[6357]), .B(x[6357]), .Z(n15233) );
  XNOR U23607 ( .A(n15226), .B(n15225), .Z(n15227) );
  XNOR U23608 ( .A(n15222), .B(n15221), .Z(n15225) );
  XOR U23609 ( .A(n15224), .B(n15223), .Z(n15221) );
  XOR U23610 ( .A(y[6356]), .B(x[6356]), .Z(n15223) );
  XOR U23611 ( .A(y[6355]), .B(x[6355]), .Z(n15224) );
  XOR U23612 ( .A(y[6354]), .B(x[6354]), .Z(n15222) );
  XOR U23613 ( .A(n15216), .B(n15215), .Z(n15226) );
  XOR U23614 ( .A(n15218), .B(n15217), .Z(n15215) );
  XOR U23615 ( .A(y[6353]), .B(x[6353]), .Z(n15217) );
  XOR U23616 ( .A(y[6352]), .B(x[6352]), .Z(n15218) );
  XOR U23617 ( .A(y[6351]), .B(x[6351]), .Z(n15216) );
  NAND U23618 ( .A(n15279), .B(n15280), .Z(N64028) );
  NAND U23619 ( .A(n15281), .B(n15282), .Z(n15280) );
  NANDN U23620 ( .A(n15283), .B(n15284), .Z(n15282) );
  NANDN U23621 ( .A(n15284), .B(n15283), .Z(n15279) );
  XOR U23622 ( .A(n15283), .B(n15285), .Z(N64027) );
  XNOR U23623 ( .A(n15281), .B(n15284), .Z(n15285) );
  NAND U23624 ( .A(n15286), .B(n15287), .Z(n15284) );
  NAND U23625 ( .A(n15288), .B(n15289), .Z(n15287) );
  NANDN U23626 ( .A(n15290), .B(n15291), .Z(n15289) );
  NANDN U23627 ( .A(n15291), .B(n15290), .Z(n15286) );
  AND U23628 ( .A(n15292), .B(n15293), .Z(n15281) );
  NAND U23629 ( .A(n15294), .B(n15295), .Z(n15293) );
  NANDN U23630 ( .A(n15296), .B(n15297), .Z(n15295) );
  NANDN U23631 ( .A(n15297), .B(n15296), .Z(n15292) );
  IV U23632 ( .A(n15298), .Z(n15297) );
  AND U23633 ( .A(n15299), .B(n15300), .Z(n15283) );
  NAND U23634 ( .A(n15301), .B(n15302), .Z(n15300) );
  NANDN U23635 ( .A(n15303), .B(n15304), .Z(n15302) );
  NANDN U23636 ( .A(n15304), .B(n15303), .Z(n15299) );
  XOR U23637 ( .A(n15296), .B(n15305), .Z(N64026) );
  XNOR U23638 ( .A(n15294), .B(n15298), .Z(n15305) );
  XOR U23639 ( .A(n15291), .B(n15306), .Z(n15298) );
  XNOR U23640 ( .A(n15288), .B(n15290), .Z(n15306) );
  AND U23641 ( .A(n15307), .B(n15308), .Z(n15290) );
  NANDN U23642 ( .A(n15309), .B(n15310), .Z(n15308) );
  OR U23643 ( .A(n15311), .B(n15312), .Z(n15310) );
  IV U23644 ( .A(n15313), .Z(n15312) );
  NANDN U23645 ( .A(n15313), .B(n15311), .Z(n15307) );
  AND U23646 ( .A(n15314), .B(n15315), .Z(n15288) );
  NAND U23647 ( .A(n15316), .B(n15317), .Z(n15315) );
  NANDN U23648 ( .A(n15318), .B(n15319), .Z(n15317) );
  NANDN U23649 ( .A(n15319), .B(n15318), .Z(n15314) );
  IV U23650 ( .A(n15320), .Z(n15319) );
  NAND U23651 ( .A(n15321), .B(n15322), .Z(n15291) );
  NANDN U23652 ( .A(n15323), .B(n15324), .Z(n15322) );
  NANDN U23653 ( .A(n15325), .B(n15326), .Z(n15324) );
  NANDN U23654 ( .A(n15326), .B(n15325), .Z(n15321) );
  IV U23655 ( .A(n15327), .Z(n15325) );
  AND U23656 ( .A(n15328), .B(n15329), .Z(n15294) );
  NAND U23657 ( .A(n15330), .B(n15331), .Z(n15329) );
  NANDN U23658 ( .A(n15332), .B(n15333), .Z(n15331) );
  NANDN U23659 ( .A(n15333), .B(n15332), .Z(n15328) );
  XOR U23660 ( .A(n15304), .B(n15334), .Z(n15296) );
  XNOR U23661 ( .A(n15301), .B(n15303), .Z(n15334) );
  AND U23662 ( .A(n15335), .B(n15336), .Z(n15303) );
  NANDN U23663 ( .A(n15337), .B(n15338), .Z(n15336) );
  OR U23664 ( .A(n15339), .B(n15340), .Z(n15338) );
  IV U23665 ( .A(n15341), .Z(n15340) );
  NANDN U23666 ( .A(n15341), .B(n15339), .Z(n15335) );
  AND U23667 ( .A(n15342), .B(n15343), .Z(n15301) );
  NAND U23668 ( .A(n15344), .B(n15345), .Z(n15343) );
  NANDN U23669 ( .A(n15346), .B(n15347), .Z(n15345) );
  NANDN U23670 ( .A(n15347), .B(n15346), .Z(n15342) );
  IV U23671 ( .A(n15348), .Z(n15347) );
  NAND U23672 ( .A(n15349), .B(n15350), .Z(n15304) );
  NANDN U23673 ( .A(n15351), .B(n15352), .Z(n15350) );
  NANDN U23674 ( .A(n15353), .B(n15354), .Z(n15352) );
  NANDN U23675 ( .A(n15354), .B(n15353), .Z(n15349) );
  IV U23676 ( .A(n15355), .Z(n15353) );
  XOR U23677 ( .A(n15330), .B(n15356), .Z(N64025) );
  XNOR U23678 ( .A(n15333), .B(n15332), .Z(n15356) );
  XNOR U23679 ( .A(n15344), .B(n15357), .Z(n15332) );
  XNOR U23680 ( .A(n15348), .B(n15346), .Z(n15357) );
  XOR U23681 ( .A(n15354), .B(n15358), .Z(n15346) );
  XNOR U23682 ( .A(n15351), .B(n15355), .Z(n15358) );
  AND U23683 ( .A(n15359), .B(n15360), .Z(n15355) );
  NAND U23684 ( .A(n15361), .B(n15362), .Z(n15360) );
  NAND U23685 ( .A(n15363), .B(n15364), .Z(n15359) );
  AND U23686 ( .A(n15365), .B(n15366), .Z(n15351) );
  NAND U23687 ( .A(n15367), .B(n15368), .Z(n15366) );
  NAND U23688 ( .A(n15369), .B(n15370), .Z(n15365) );
  NANDN U23689 ( .A(n15371), .B(n15372), .Z(n15354) );
  ANDN U23690 ( .B(n15373), .A(n15374), .Z(n15348) );
  XNOR U23691 ( .A(n15339), .B(n15375), .Z(n15344) );
  XNOR U23692 ( .A(n15337), .B(n15341), .Z(n15375) );
  AND U23693 ( .A(n15376), .B(n15377), .Z(n15341) );
  NAND U23694 ( .A(n15378), .B(n15379), .Z(n15377) );
  NAND U23695 ( .A(n15380), .B(n15381), .Z(n15376) );
  AND U23696 ( .A(n15382), .B(n15383), .Z(n15337) );
  NAND U23697 ( .A(n15384), .B(n15385), .Z(n15383) );
  NAND U23698 ( .A(n15386), .B(n15387), .Z(n15382) );
  AND U23699 ( .A(n15388), .B(n15389), .Z(n15339) );
  NAND U23700 ( .A(n15390), .B(n15391), .Z(n15333) );
  XNOR U23701 ( .A(n15316), .B(n15392), .Z(n15330) );
  XNOR U23702 ( .A(n15320), .B(n15318), .Z(n15392) );
  XOR U23703 ( .A(n15326), .B(n15393), .Z(n15318) );
  XNOR U23704 ( .A(n15323), .B(n15327), .Z(n15393) );
  AND U23705 ( .A(n15394), .B(n15395), .Z(n15327) );
  NAND U23706 ( .A(n15396), .B(n15397), .Z(n15395) );
  NAND U23707 ( .A(n15398), .B(n15399), .Z(n15394) );
  AND U23708 ( .A(n15400), .B(n15401), .Z(n15323) );
  NAND U23709 ( .A(n15402), .B(n15403), .Z(n15401) );
  NAND U23710 ( .A(n15404), .B(n15405), .Z(n15400) );
  NANDN U23711 ( .A(n15406), .B(n15407), .Z(n15326) );
  ANDN U23712 ( .B(n15408), .A(n15409), .Z(n15320) );
  XNOR U23713 ( .A(n15311), .B(n15410), .Z(n15316) );
  XNOR U23714 ( .A(n15309), .B(n15313), .Z(n15410) );
  AND U23715 ( .A(n15411), .B(n15412), .Z(n15313) );
  NAND U23716 ( .A(n15413), .B(n15414), .Z(n15412) );
  NAND U23717 ( .A(n15415), .B(n15416), .Z(n15411) );
  AND U23718 ( .A(n15417), .B(n15418), .Z(n15309) );
  NAND U23719 ( .A(n15419), .B(n15420), .Z(n15418) );
  NAND U23720 ( .A(n15421), .B(n15422), .Z(n15417) );
  AND U23721 ( .A(n15423), .B(n15424), .Z(n15311) );
  XOR U23722 ( .A(n15391), .B(n15390), .Z(N64024) );
  XNOR U23723 ( .A(n15408), .B(n15409), .Z(n15390) );
  XNOR U23724 ( .A(n15423), .B(n15424), .Z(n15409) );
  XOR U23725 ( .A(n15420), .B(n15419), .Z(n15424) );
  XOR U23726 ( .A(y[6348]), .B(x[6348]), .Z(n15419) );
  XOR U23727 ( .A(n15422), .B(n15421), .Z(n15420) );
  XOR U23728 ( .A(y[6350]), .B(x[6350]), .Z(n15421) );
  XOR U23729 ( .A(y[6349]), .B(x[6349]), .Z(n15422) );
  XOR U23730 ( .A(n15414), .B(n15413), .Z(n15423) );
  XOR U23731 ( .A(n15416), .B(n15415), .Z(n15413) );
  XOR U23732 ( .A(y[6347]), .B(x[6347]), .Z(n15415) );
  XOR U23733 ( .A(y[6346]), .B(x[6346]), .Z(n15416) );
  XOR U23734 ( .A(y[6345]), .B(x[6345]), .Z(n15414) );
  XNOR U23735 ( .A(n15407), .B(n15406), .Z(n15408) );
  XNOR U23736 ( .A(n15403), .B(n15402), .Z(n15406) );
  XOR U23737 ( .A(n15405), .B(n15404), .Z(n15402) );
  XOR U23738 ( .A(y[6344]), .B(x[6344]), .Z(n15404) );
  XOR U23739 ( .A(y[6343]), .B(x[6343]), .Z(n15405) );
  XOR U23740 ( .A(y[6342]), .B(x[6342]), .Z(n15403) );
  XOR U23741 ( .A(n15397), .B(n15396), .Z(n15407) );
  XOR U23742 ( .A(n15399), .B(n15398), .Z(n15396) );
  XOR U23743 ( .A(y[6341]), .B(x[6341]), .Z(n15398) );
  XOR U23744 ( .A(y[6340]), .B(x[6340]), .Z(n15399) );
  XOR U23745 ( .A(y[6339]), .B(x[6339]), .Z(n15397) );
  XNOR U23746 ( .A(n15373), .B(n15374), .Z(n15391) );
  XNOR U23747 ( .A(n15388), .B(n15389), .Z(n15374) );
  XOR U23748 ( .A(n15385), .B(n15384), .Z(n15389) );
  XOR U23749 ( .A(y[6336]), .B(x[6336]), .Z(n15384) );
  XOR U23750 ( .A(n15387), .B(n15386), .Z(n15385) );
  XOR U23751 ( .A(y[6338]), .B(x[6338]), .Z(n15386) );
  XOR U23752 ( .A(y[6337]), .B(x[6337]), .Z(n15387) );
  XOR U23753 ( .A(n15379), .B(n15378), .Z(n15388) );
  XOR U23754 ( .A(n15381), .B(n15380), .Z(n15378) );
  XOR U23755 ( .A(y[6335]), .B(x[6335]), .Z(n15380) );
  XOR U23756 ( .A(y[6334]), .B(x[6334]), .Z(n15381) );
  XOR U23757 ( .A(y[6333]), .B(x[6333]), .Z(n15379) );
  XNOR U23758 ( .A(n15372), .B(n15371), .Z(n15373) );
  XNOR U23759 ( .A(n15368), .B(n15367), .Z(n15371) );
  XOR U23760 ( .A(n15370), .B(n15369), .Z(n15367) );
  XOR U23761 ( .A(y[6332]), .B(x[6332]), .Z(n15369) );
  XOR U23762 ( .A(y[6331]), .B(x[6331]), .Z(n15370) );
  XOR U23763 ( .A(y[6330]), .B(x[6330]), .Z(n15368) );
  XOR U23764 ( .A(n15362), .B(n15361), .Z(n15372) );
  XOR U23765 ( .A(n15364), .B(n15363), .Z(n15361) );
  XOR U23766 ( .A(y[6329]), .B(x[6329]), .Z(n15363) );
  XOR U23767 ( .A(y[6328]), .B(x[6328]), .Z(n15364) );
  XOR U23768 ( .A(y[6327]), .B(x[6327]), .Z(n15362) );
  NAND U23769 ( .A(n15425), .B(n15426), .Z(N64015) );
  NAND U23770 ( .A(n15427), .B(n15428), .Z(n15426) );
  NANDN U23771 ( .A(n15429), .B(n15430), .Z(n15428) );
  NANDN U23772 ( .A(n15430), .B(n15429), .Z(n15425) );
  XOR U23773 ( .A(n15429), .B(n15431), .Z(N64014) );
  XNOR U23774 ( .A(n15427), .B(n15430), .Z(n15431) );
  NAND U23775 ( .A(n15432), .B(n15433), .Z(n15430) );
  NAND U23776 ( .A(n15434), .B(n15435), .Z(n15433) );
  NANDN U23777 ( .A(n15436), .B(n15437), .Z(n15435) );
  NANDN U23778 ( .A(n15437), .B(n15436), .Z(n15432) );
  AND U23779 ( .A(n15438), .B(n15439), .Z(n15427) );
  NAND U23780 ( .A(n15440), .B(n15441), .Z(n15439) );
  NANDN U23781 ( .A(n15442), .B(n15443), .Z(n15441) );
  NANDN U23782 ( .A(n15443), .B(n15442), .Z(n15438) );
  IV U23783 ( .A(n15444), .Z(n15443) );
  AND U23784 ( .A(n15445), .B(n15446), .Z(n15429) );
  NAND U23785 ( .A(n15447), .B(n15448), .Z(n15446) );
  NANDN U23786 ( .A(n15449), .B(n15450), .Z(n15448) );
  NANDN U23787 ( .A(n15450), .B(n15449), .Z(n15445) );
  XOR U23788 ( .A(n15442), .B(n15451), .Z(N64013) );
  XNOR U23789 ( .A(n15440), .B(n15444), .Z(n15451) );
  XOR U23790 ( .A(n15437), .B(n15452), .Z(n15444) );
  XNOR U23791 ( .A(n15434), .B(n15436), .Z(n15452) );
  AND U23792 ( .A(n15453), .B(n15454), .Z(n15436) );
  NANDN U23793 ( .A(n15455), .B(n15456), .Z(n15454) );
  OR U23794 ( .A(n15457), .B(n15458), .Z(n15456) );
  IV U23795 ( .A(n15459), .Z(n15458) );
  NANDN U23796 ( .A(n15459), .B(n15457), .Z(n15453) );
  AND U23797 ( .A(n15460), .B(n15461), .Z(n15434) );
  NAND U23798 ( .A(n15462), .B(n15463), .Z(n15461) );
  NANDN U23799 ( .A(n15464), .B(n15465), .Z(n15463) );
  NANDN U23800 ( .A(n15465), .B(n15464), .Z(n15460) );
  IV U23801 ( .A(n15466), .Z(n15465) );
  NAND U23802 ( .A(n15467), .B(n15468), .Z(n15437) );
  NANDN U23803 ( .A(n15469), .B(n15470), .Z(n15468) );
  NANDN U23804 ( .A(n15471), .B(n15472), .Z(n15470) );
  NANDN U23805 ( .A(n15472), .B(n15471), .Z(n15467) );
  IV U23806 ( .A(n15473), .Z(n15471) );
  AND U23807 ( .A(n15474), .B(n15475), .Z(n15440) );
  NAND U23808 ( .A(n15476), .B(n15477), .Z(n15475) );
  NANDN U23809 ( .A(n15478), .B(n15479), .Z(n15477) );
  NANDN U23810 ( .A(n15479), .B(n15478), .Z(n15474) );
  XOR U23811 ( .A(n15450), .B(n15480), .Z(n15442) );
  XNOR U23812 ( .A(n15447), .B(n15449), .Z(n15480) );
  AND U23813 ( .A(n15481), .B(n15482), .Z(n15449) );
  NANDN U23814 ( .A(n15483), .B(n15484), .Z(n15482) );
  OR U23815 ( .A(n15485), .B(n15486), .Z(n15484) );
  IV U23816 ( .A(n15487), .Z(n15486) );
  NANDN U23817 ( .A(n15487), .B(n15485), .Z(n15481) );
  AND U23818 ( .A(n15488), .B(n15489), .Z(n15447) );
  NAND U23819 ( .A(n15490), .B(n15491), .Z(n15489) );
  NANDN U23820 ( .A(n15492), .B(n15493), .Z(n15491) );
  NANDN U23821 ( .A(n15493), .B(n15492), .Z(n15488) );
  IV U23822 ( .A(n15494), .Z(n15493) );
  NAND U23823 ( .A(n15495), .B(n15496), .Z(n15450) );
  NANDN U23824 ( .A(n15497), .B(n15498), .Z(n15496) );
  NANDN U23825 ( .A(n15499), .B(n15500), .Z(n15498) );
  NANDN U23826 ( .A(n15500), .B(n15499), .Z(n15495) );
  IV U23827 ( .A(n15501), .Z(n15499) );
  XOR U23828 ( .A(n15476), .B(n15502), .Z(N64012) );
  XNOR U23829 ( .A(n15479), .B(n15478), .Z(n15502) );
  XNOR U23830 ( .A(n15490), .B(n15503), .Z(n15478) );
  XNOR U23831 ( .A(n15494), .B(n15492), .Z(n15503) );
  XOR U23832 ( .A(n15500), .B(n15504), .Z(n15492) );
  XNOR U23833 ( .A(n15497), .B(n15501), .Z(n15504) );
  AND U23834 ( .A(n15505), .B(n15506), .Z(n15501) );
  NAND U23835 ( .A(n15507), .B(n15508), .Z(n15506) );
  NAND U23836 ( .A(n15509), .B(n15510), .Z(n15505) );
  AND U23837 ( .A(n15511), .B(n15512), .Z(n15497) );
  NAND U23838 ( .A(n15513), .B(n15514), .Z(n15512) );
  NAND U23839 ( .A(n15515), .B(n15516), .Z(n15511) );
  NANDN U23840 ( .A(n15517), .B(n15518), .Z(n15500) );
  ANDN U23841 ( .B(n15519), .A(n15520), .Z(n15494) );
  XNOR U23842 ( .A(n15485), .B(n15521), .Z(n15490) );
  XNOR U23843 ( .A(n15483), .B(n15487), .Z(n15521) );
  AND U23844 ( .A(n15522), .B(n15523), .Z(n15487) );
  NAND U23845 ( .A(n15524), .B(n15525), .Z(n15523) );
  NAND U23846 ( .A(n15526), .B(n15527), .Z(n15522) );
  AND U23847 ( .A(n15528), .B(n15529), .Z(n15483) );
  NAND U23848 ( .A(n15530), .B(n15531), .Z(n15529) );
  NAND U23849 ( .A(n15532), .B(n15533), .Z(n15528) );
  AND U23850 ( .A(n15534), .B(n15535), .Z(n15485) );
  NAND U23851 ( .A(n15536), .B(n15537), .Z(n15479) );
  XNOR U23852 ( .A(n15462), .B(n15538), .Z(n15476) );
  XNOR U23853 ( .A(n15466), .B(n15464), .Z(n15538) );
  XOR U23854 ( .A(n15472), .B(n15539), .Z(n15464) );
  XNOR U23855 ( .A(n15469), .B(n15473), .Z(n15539) );
  AND U23856 ( .A(n15540), .B(n15541), .Z(n15473) );
  NAND U23857 ( .A(n15542), .B(n15543), .Z(n15541) );
  NAND U23858 ( .A(n15544), .B(n15545), .Z(n15540) );
  AND U23859 ( .A(n15546), .B(n15547), .Z(n15469) );
  NAND U23860 ( .A(n15548), .B(n15549), .Z(n15547) );
  NAND U23861 ( .A(n15550), .B(n15551), .Z(n15546) );
  NANDN U23862 ( .A(n15552), .B(n15553), .Z(n15472) );
  ANDN U23863 ( .B(n15554), .A(n15555), .Z(n15466) );
  XNOR U23864 ( .A(n15457), .B(n15556), .Z(n15462) );
  XNOR U23865 ( .A(n15455), .B(n15459), .Z(n15556) );
  AND U23866 ( .A(n15557), .B(n15558), .Z(n15459) );
  NAND U23867 ( .A(n15559), .B(n15560), .Z(n15558) );
  NAND U23868 ( .A(n15561), .B(n15562), .Z(n15557) );
  AND U23869 ( .A(n15563), .B(n15564), .Z(n15455) );
  NAND U23870 ( .A(n15565), .B(n15566), .Z(n15564) );
  NAND U23871 ( .A(n15567), .B(n15568), .Z(n15563) );
  AND U23872 ( .A(n15569), .B(n15570), .Z(n15457) );
  XOR U23873 ( .A(n15537), .B(n15536), .Z(N64011) );
  XNOR U23874 ( .A(n15554), .B(n15555), .Z(n15536) );
  XNOR U23875 ( .A(n15569), .B(n15570), .Z(n15555) );
  XOR U23876 ( .A(n15566), .B(n15565), .Z(n15570) );
  XOR U23877 ( .A(y[6324]), .B(x[6324]), .Z(n15565) );
  XOR U23878 ( .A(n15568), .B(n15567), .Z(n15566) );
  XOR U23879 ( .A(y[6326]), .B(x[6326]), .Z(n15567) );
  XOR U23880 ( .A(y[6325]), .B(x[6325]), .Z(n15568) );
  XOR U23881 ( .A(n15560), .B(n15559), .Z(n15569) );
  XOR U23882 ( .A(n15562), .B(n15561), .Z(n15559) );
  XOR U23883 ( .A(y[6323]), .B(x[6323]), .Z(n15561) );
  XOR U23884 ( .A(y[6322]), .B(x[6322]), .Z(n15562) );
  XOR U23885 ( .A(y[6321]), .B(x[6321]), .Z(n15560) );
  XNOR U23886 ( .A(n15553), .B(n15552), .Z(n15554) );
  XNOR U23887 ( .A(n15549), .B(n15548), .Z(n15552) );
  XOR U23888 ( .A(n15551), .B(n15550), .Z(n15548) );
  XOR U23889 ( .A(y[6320]), .B(x[6320]), .Z(n15550) );
  XOR U23890 ( .A(y[6319]), .B(x[6319]), .Z(n15551) );
  XOR U23891 ( .A(y[6318]), .B(x[6318]), .Z(n15549) );
  XOR U23892 ( .A(n15543), .B(n15542), .Z(n15553) );
  XOR U23893 ( .A(n15545), .B(n15544), .Z(n15542) );
  XOR U23894 ( .A(y[6317]), .B(x[6317]), .Z(n15544) );
  XOR U23895 ( .A(y[6316]), .B(x[6316]), .Z(n15545) );
  XOR U23896 ( .A(y[6315]), .B(x[6315]), .Z(n15543) );
  XNOR U23897 ( .A(n15519), .B(n15520), .Z(n15537) );
  XNOR U23898 ( .A(n15534), .B(n15535), .Z(n15520) );
  XOR U23899 ( .A(n15531), .B(n15530), .Z(n15535) );
  XOR U23900 ( .A(y[6312]), .B(x[6312]), .Z(n15530) );
  XOR U23901 ( .A(n15533), .B(n15532), .Z(n15531) );
  XOR U23902 ( .A(y[6314]), .B(x[6314]), .Z(n15532) );
  XOR U23903 ( .A(y[6313]), .B(x[6313]), .Z(n15533) );
  XOR U23904 ( .A(n15525), .B(n15524), .Z(n15534) );
  XOR U23905 ( .A(n15527), .B(n15526), .Z(n15524) );
  XOR U23906 ( .A(y[6311]), .B(x[6311]), .Z(n15526) );
  XOR U23907 ( .A(y[6310]), .B(x[6310]), .Z(n15527) );
  XOR U23908 ( .A(y[6309]), .B(x[6309]), .Z(n15525) );
  XNOR U23909 ( .A(n15518), .B(n15517), .Z(n15519) );
  XNOR U23910 ( .A(n15514), .B(n15513), .Z(n15517) );
  XOR U23911 ( .A(n15516), .B(n15515), .Z(n15513) );
  XOR U23912 ( .A(y[6308]), .B(x[6308]), .Z(n15515) );
  XOR U23913 ( .A(y[6307]), .B(x[6307]), .Z(n15516) );
  XOR U23914 ( .A(y[6306]), .B(x[6306]), .Z(n15514) );
  XOR U23915 ( .A(n15508), .B(n15507), .Z(n15518) );
  XOR U23916 ( .A(n15510), .B(n15509), .Z(n15507) );
  XOR U23917 ( .A(y[6305]), .B(x[6305]), .Z(n15509) );
  XOR U23918 ( .A(y[6304]), .B(x[6304]), .Z(n15510) );
  XOR U23919 ( .A(y[6303]), .B(x[6303]), .Z(n15508) );
  NAND U23920 ( .A(n15571), .B(n15572), .Z(N64002) );
  NAND U23921 ( .A(n15573), .B(n15574), .Z(n15572) );
  NANDN U23922 ( .A(n15575), .B(n15576), .Z(n15574) );
  NANDN U23923 ( .A(n15576), .B(n15575), .Z(n15571) );
  XOR U23924 ( .A(n15575), .B(n15577), .Z(N64001) );
  XNOR U23925 ( .A(n15573), .B(n15576), .Z(n15577) );
  NAND U23926 ( .A(n15578), .B(n15579), .Z(n15576) );
  NAND U23927 ( .A(n15580), .B(n15581), .Z(n15579) );
  NANDN U23928 ( .A(n15582), .B(n15583), .Z(n15581) );
  NANDN U23929 ( .A(n15583), .B(n15582), .Z(n15578) );
  AND U23930 ( .A(n15584), .B(n15585), .Z(n15573) );
  NAND U23931 ( .A(n15586), .B(n15587), .Z(n15585) );
  NANDN U23932 ( .A(n15588), .B(n15589), .Z(n15587) );
  NANDN U23933 ( .A(n15589), .B(n15588), .Z(n15584) );
  IV U23934 ( .A(n15590), .Z(n15589) );
  AND U23935 ( .A(n15591), .B(n15592), .Z(n15575) );
  NAND U23936 ( .A(n15593), .B(n15594), .Z(n15592) );
  NANDN U23937 ( .A(n15595), .B(n15596), .Z(n15594) );
  NANDN U23938 ( .A(n15596), .B(n15595), .Z(n15591) );
  XOR U23939 ( .A(n15588), .B(n15597), .Z(N64000) );
  XNOR U23940 ( .A(n15586), .B(n15590), .Z(n15597) );
  XOR U23941 ( .A(n15583), .B(n15598), .Z(n15590) );
  XNOR U23942 ( .A(n15580), .B(n15582), .Z(n15598) );
  AND U23943 ( .A(n15599), .B(n15600), .Z(n15582) );
  NANDN U23944 ( .A(n15601), .B(n15602), .Z(n15600) );
  OR U23945 ( .A(n15603), .B(n15604), .Z(n15602) );
  IV U23946 ( .A(n15605), .Z(n15604) );
  NANDN U23947 ( .A(n15605), .B(n15603), .Z(n15599) );
  AND U23948 ( .A(n15606), .B(n15607), .Z(n15580) );
  NAND U23949 ( .A(n15608), .B(n15609), .Z(n15607) );
  NANDN U23950 ( .A(n15610), .B(n15611), .Z(n15609) );
  NANDN U23951 ( .A(n15611), .B(n15610), .Z(n15606) );
  IV U23952 ( .A(n15612), .Z(n15611) );
  NAND U23953 ( .A(n15613), .B(n15614), .Z(n15583) );
  NANDN U23954 ( .A(n15615), .B(n15616), .Z(n15614) );
  NANDN U23955 ( .A(n15617), .B(n15618), .Z(n15616) );
  NANDN U23956 ( .A(n15618), .B(n15617), .Z(n15613) );
  IV U23957 ( .A(n15619), .Z(n15617) );
  AND U23958 ( .A(n15620), .B(n15621), .Z(n15586) );
  NAND U23959 ( .A(n15622), .B(n15623), .Z(n15621) );
  NANDN U23960 ( .A(n15624), .B(n15625), .Z(n15623) );
  NANDN U23961 ( .A(n15625), .B(n15624), .Z(n15620) );
  XOR U23962 ( .A(n15596), .B(n15626), .Z(n15588) );
  XNOR U23963 ( .A(n15593), .B(n15595), .Z(n15626) );
  AND U23964 ( .A(n15627), .B(n15628), .Z(n15595) );
  NANDN U23965 ( .A(n15629), .B(n15630), .Z(n15628) );
  OR U23966 ( .A(n15631), .B(n15632), .Z(n15630) );
  IV U23967 ( .A(n15633), .Z(n15632) );
  NANDN U23968 ( .A(n15633), .B(n15631), .Z(n15627) );
  AND U23969 ( .A(n15634), .B(n15635), .Z(n15593) );
  NAND U23970 ( .A(n15636), .B(n15637), .Z(n15635) );
  NANDN U23971 ( .A(n15638), .B(n15639), .Z(n15637) );
  NANDN U23972 ( .A(n15639), .B(n15638), .Z(n15634) );
  IV U23973 ( .A(n15640), .Z(n15639) );
  NAND U23974 ( .A(n15641), .B(n15642), .Z(n15596) );
  NANDN U23975 ( .A(n15643), .B(n15644), .Z(n15642) );
  NANDN U23976 ( .A(n15645), .B(n15646), .Z(n15644) );
  NANDN U23977 ( .A(n15646), .B(n15645), .Z(n15641) );
  IV U23978 ( .A(n15647), .Z(n15645) );
  XOR U23979 ( .A(n15622), .B(n15648), .Z(N63999) );
  XNOR U23980 ( .A(n15625), .B(n15624), .Z(n15648) );
  XNOR U23981 ( .A(n15636), .B(n15649), .Z(n15624) );
  XNOR U23982 ( .A(n15640), .B(n15638), .Z(n15649) );
  XOR U23983 ( .A(n15646), .B(n15650), .Z(n15638) );
  XNOR U23984 ( .A(n15643), .B(n15647), .Z(n15650) );
  AND U23985 ( .A(n15651), .B(n15652), .Z(n15647) );
  NAND U23986 ( .A(n15653), .B(n15654), .Z(n15652) );
  NAND U23987 ( .A(n15655), .B(n15656), .Z(n15651) );
  AND U23988 ( .A(n15657), .B(n15658), .Z(n15643) );
  NAND U23989 ( .A(n15659), .B(n15660), .Z(n15658) );
  NAND U23990 ( .A(n15661), .B(n15662), .Z(n15657) );
  NANDN U23991 ( .A(n15663), .B(n15664), .Z(n15646) );
  ANDN U23992 ( .B(n15665), .A(n15666), .Z(n15640) );
  XNOR U23993 ( .A(n15631), .B(n15667), .Z(n15636) );
  XNOR U23994 ( .A(n15629), .B(n15633), .Z(n15667) );
  AND U23995 ( .A(n15668), .B(n15669), .Z(n15633) );
  NAND U23996 ( .A(n15670), .B(n15671), .Z(n15669) );
  NAND U23997 ( .A(n15672), .B(n15673), .Z(n15668) );
  AND U23998 ( .A(n15674), .B(n15675), .Z(n15629) );
  NAND U23999 ( .A(n15676), .B(n15677), .Z(n15675) );
  NAND U24000 ( .A(n15678), .B(n15679), .Z(n15674) );
  AND U24001 ( .A(n15680), .B(n15681), .Z(n15631) );
  NAND U24002 ( .A(n15682), .B(n15683), .Z(n15625) );
  XNOR U24003 ( .A(n15608), .B(n15684), .Z(n15622) );
  XNOR U24004 ( .A(n15612), .B(n15610), .Z(n15684) );
  XOR U24005 ( .A(n15618), .B(n15685), .Z(n15610) );
  XNOR U24006 ( .A(n15615), .B(n15619), .Z(n15685) );
  AND U24007 ( .A(n15686), .B(n15687), .Z(n15619) );
  NAND U24008 ( .A(n15688), .B(n15689), .Z(n15687) );
  NAND U24009 ( .A(n15690), .B(n15691), .Z(n15686) );
  AND U24010 ( .A(n15692), .B(n15693), .Z(n15615) );
  NAND U24011 ( .A(n15694), .B(n15695), .Z(n15693) );
  NAND U24012 ( .A(n15696), .B(n15697), .Z(n15692) );
  NANDN U24013 ( .A(n15698), .B(n15699), .Z(n15618) );
  ANDN U24014 ( .B(n15700), .A(n15701), .Z(n15612) );
  XNOR U24015 ( .A(n15603), .B(n15702), .Z(n15608) );
  XNOR U24016 ( .A(n15601), .B(n15605), .Z(n15702) );
  AND U24017 ( .A(n15703), .B(n15704), .Z(n15605) );
  NAND U24018 ( .A(n15705), .B(n15706), .Z(n15704) );
  NAND U24019 ( .A(n15707), .B(n15708), .Z(n15703) );
  AND U24020 ( .A(n15709), .B(n15710), .Z(n15601) );
  NAND U24021 ( .A(n15711), .B(n15712), .Z(n15710) );
  NAND U24022 ( .A(n15713), .B(n15714), .Z(n15709) );
  AND U24023 ( .A(n15715), .B(n15716), .Z(n15603) );
  XOR U24024 ( .A(n15683), .B(n15682), .Z(N63998) );
  XNOR U24025 ( .A(n15700), .B(n15701), .Z(n15682) );
  XNOR U24026 ( .A(n15715), .B(n15716), .Z(n15701) );
  XOR U24027 ( .A(n15712), .B(n15711), .Z(n15716) );
  XOR U24028 ( .A(y[6300]), .B(x[6300]), .Z(n15711) );
  XOR U24029 ( .A(n15714), .B(n15713), .Z(n15712) );
  XOR U24030 ( .A(y[6302]), .B(x[6302]), .Z(n15713) );
  XOR U24031 ( .A(y[6301]), .B(x[6301]), .Z(n15714) );
  XOR U24032 ( .A(n15706), .B(n15705), .Z(n15715) );
  XOR U24033 ( .A(n15708), .B(n15707), .Z(n15705) );
  XOR U24034 ( .A(y[6299]), .B(x[6299]), .Z(n15707) );
  XOR U24035 ( .A(y[6298]), .B(x[6298]), .Z(n15708) );
  XOR U24036 ( .A(y[6297]), .B(x[6297]), .Z(n15706) );
  XNOR U24037 ( .A(n15699), .B(n15698), .Z(n15700) );
  XNOR U24038 ( .A(n15695), .B(n15694), .Z(n15698) );
  XOR U24039 ( .A(n15697), .B(n15696), .Z(n15694) );
  XOR U24040 ( .A(y[6296]), .B(x[6296]), .Z(n15696) );
  XOR U24041 ( .A(y[6295]), .B(x[6295]), .Z(n15697) );
  XOR U24042 ( .A(y[6294]), .B(x[6294]), .Z(n15695) );
  XOR U24043 ( .A(n15689), .B(n15688), .Z(n15699) );
  XOR U24044 ( .A(n15691), .B(n15690), .Z(n15688) );
  XOR U24045 ( .A(y[6293]), .B(x[6293]), .Z(n15690) );
  XOR U24046 ( .A(y[6292]), .B(x[6292]), .Z(n15691) );
  XOR U24047 ( .A(y[6291]), .B(x[6291]), .Z(n15689) );
  XNOR U24048 ( .A(n15665), .B(n15666), .Z(n15683) );
  XNOR U24049 ( .A(n15680), .B(n15681), .Z(n15666) );
  XOR U24050 ( .A(n15677), .B(n15676), .Z(n15681) );
  XOR U24051 ( .A(y[6288]), .B(x[6288]), .Z(n15676) );
  XOR U24052 ( .A(n15679), .B(n15678), .Z(n15677) );
  XOR U24053 ( .A(y[6290]), .B(x[6290]), .Z(n15678) );
  XOR U24054 ( .A(y[6289]), .B(x[6289]), .Z(n15679) );
  XOR U24055 ( .A(n15671), .B(n15670), .Z(n15680) );
  XOR U24056 ( .A(n15673), .B(n15672), .Z(n15670) );
  XOR U24057 ( .A(y[6287]), .B(x[6287]), .Z(n15672) );
  XOR U24058 ( .A(y[6286]), .B(x[6286]), .Z(n15673) );
  XOR U24059 ( .A(y[6285]), .B(x[6285]), .Z(n15671) );
  XNOR U24060 ( .A(n15664), .B(n15663), .Z(n15665) );
  XNOR U24061 ( .A(n15660), .B(n15659), .Z(n15663) );
  XOR U24062 ( .A(n15662), .B(n15661), .Z(n15659) );
  XOR U24063 ( .A(y[6284]), .B(x[6284]), .Z(n15661) );
  XOR U24064 ( .A(y[6283]), .B(x[6283]), .Z(n15662) );
  XOR U24065 ( .A(y[6282]), .B(x[6282]), .Z(n15660) );
  XOR U24066 ( .A(n15654), .B(n15653), .Z(n15664) );
  XOR U24067 ( .A(n15656), .B(n15655), .Z(n15653) );
  XOR U24068 ( .A(y[6281]), .B(x[6281]), .Z(n15655) );
  XOR U24069 ( .A(y[6280]), .B(x[6280]), .Z(n15656) );
  XOR U24070 ( .A(y[6279]), .B(x[6279]), .Z(n15654) );
  NAND U24071 ( .A(n15717), .B(n15718), .Z(N63989) );
  NAND U24072 ( .A(n15719), .B(n15720), .Z(n15718) );
  NANDN U24073 ( .A(n15721), .B(n15722), .Z(n15720) );
  NANDN U24074 ( .A(n15722), .B(n15721), .Z(n15717) );
  XOR U24075 ( .A(n15721), .B(n15723), .Z(N63988) );
  XNOR U24076 ( .A(n15719), .B(n15722), .Z(n15723) );
  NAND U24077 ( .A(n15724), .B(n15725), .Z(n15722) );
  NAND U24078 ( .A(n15726), .B(n15727), .Z(n15725) );
  NANDN U24079 ( .A(n15728), .B(n15729), .Z(n15727) );
  NANDN U24080 ( .A(n15729), .B(n15728), .Z(n15724) );
  AND U24081 ( .A(n15730), .B(n15731), .Z(n15719) );
  NAND U24082 ( .A(n15732), .B(n15733), .Z(n15731) );
  NANDN U24083 ( .A(n15734), .B(n15735), .Z(n15733) );
  NANDN U24084 ( .A(n15735), .B(n15734), .Z(n15730) );
  IV U24085 ( .A(n15736), .Z(n15735) );
  AND U24086 ( .A(n15737), .B(n15738), .Z(n15721) );
  NAND U24087 ( .A(n15739), .B(n15740), .Z(n15738) );
  NANDN U24088 ( .A(n15741), .B(n15742), .Z(n15740) );
  NANDN U24089 ( .A(n15742), .B(n15741), .Z(n15737) );
  XOR U24090 ( .A(n15734), .B(n15743), .Z(N63987) );
  XNOR U24091 ( .A(n15732), .B(n15736), .Z(n15743) );
  XOR U24092 ( .A(n15729), .B(n15744), .Z(n15736) );
  XNOR U24093 ( .A(n15726), .B(n15728), .Z(n15744) );
  AND U24094 ( .A(n15745), .B(n15746), .Z(n15728) );
  NANDN U24095 ( .A(n15747), .B(n15748), .Z(n15746) );
  OR U24096 ( .A(n15749), .B(n15750), .Z(n15748) );
  IV U24097 ( .A(n15751), .Z(n15750) );
  NANDN U24098 ( .A(n15751), .B(n15749), .Z(n15745) );
  AND U24099 ( .A(n15752), .B(n15753), .Z(n15726) );
  NAND U24100 ( .A(n15754), .B(n15755), .Z(n15753) );
  NANDN U24101 ( .A(n15756), .B(n15757), .Z(n15755) );
  NANDN U24102 ( .A(n15757), .B(n15756), .Z(n15752) );
  IV U24103 ( .A(n15758), .Z(n15757) );
  NAND U24104 ( .A(n15759), .B(n15760), .Z(n15729) );
  NANDN U24105 ( .A(n15761), .B(n15762), .Z(n15760) );
  NANDN U24106 ( .A(n15763), .B(n15764), .Z(n15762) );
  NANDN U24107 ( .A(n15764), .B(n15763), .Z(n15759) );
  IV U24108 ( .A(n15765), .Z(n15763) );
  AND U24109 ( .A(n15766), .B(n15767), .Z(n15732) );
  NAND U24110 ( .A(n15768), .B(n15769), .Z(n15767) );
  NANDN U24111 ( .A(n15770), .B(n15771), .Z(n15769) );
  NANDN U24112 ( .A(n15771), .B(n15770), .Z(n15766) );
  XOR U24113 ( .A(n15742), .B(n15772), .Z(n15734) );
  XNOR U24114 ( .A(n15739), .B(n15741), .Z(n15772) );
  AND U24115 ( .A(n15773), .B(n15774), .Z(n15741) );
  NANDN U24116 ( .A(n15775), .B(n15776), .Z(n15774) );
  OR U24117 ( .A(n15777), .B(n15778), .Z(n15776) );
  IV U24118 ( .A(n15779), .Z(n15778) );
  NANDN U24119 ( .A(n15779), .B(n15777), .Z(n15773) );
  AND U24120 ( .A(n15780), .B(n15781), .Z(n15739) );
  NAND U24121 ( .A(n15782), .B(n15783), .Z(n15781) );
  NANDN U24122 ( .A(n15784), .B(n15785), .Z(n15783) );
  NANDN U24123 ( .A(n15785), .B(n15784), .Z(n15780) );
  IV U24124 ( .A(n15786), .Z(n15785) );
  NAND U24125 ( .A(n15787), .B(n15788), .Z(n15742) );
  NANDN U24126 ( .A(n15789), .B(n15790), .Z(n15788) );
  NANDN U24127 ( .A(n15791), .B(n15792), .Z(n15790) );
  NANDN U24128 ( .A(n15792), .B(n15791), .Z(n15787) );
  IV U24129 ( .A(n15793), .Z(n15791) );
  XOR U24130 ( .A(n15768), .B(n15794), .Z(N63986) );
  XNOR U24131 ( .A(n15771), .B(n15770), .Z(n15794) );
  XNOR U24132 ( .A(n15782), .B(n15795), .Z(n15770) );
  XNOR U24133 ( .A(n15786), .B(n15784), .Z(n15795) );
  XOR U24134 ( .A(n15792), .B(n15796), .Z(n15784) );
  XNOR U24135 ( .A(n15789), .B(n15793), .Z(n15796) );
  AND U24136 ( .A(n15797), .B(n15798), .Z(n15793) );
  NAND U24137 ( .A(n15799), .B(n15800), .Z(n15798) );
  NAND U24138 ( .A(n15801), .B(n15802), .Z(n15797) );
  AND U24139 ( .A(n15803), .B(n15804), .Z(n15789) );
  NAND U24140 ( .A(n15805), .B(n15806), .Z(n15804) );
  NAND U24141 ( .A(n15807), .B(n15808), .Z(n15803) );
  NANDN U24142 ( .A(n15809), .B(n15810), .Z(n15792) );
  ANDN U24143 ( .B(n15811), .A(n15812), .Z(n15786) );
  XNOR U24144 ( .A(n15777), .B(n15813), .Z(n15782) );
  XNOR U24145 ( .A(n15775), .B(n15779), .Z(n15813) );
  AND U24146 ( .A(n15814), .B(n15815), .Z(n15779) );
  NAND U24147 ( .A(n15816), .B(n15817), .Z(n15815) );
  NAND U24148 ( .A(n15818), .B(n15819), .Z(n15814) );
  AND U24149 ( .A(n15820), .B(n15821), .Z(n15775) );
  NAND U24150 ( .A(n15822), .B(n15823), .Z(n15821) );
  NAND U24151 ( .A(n15824), .B(n15825), .Z(n15820) );
  AND U24152 ( .A(n15826), .B(n15827), .Z(n15777) );
  NAND U24153 ( .A(n15828), .B(n15829), .Z(n15771) );
  XNOR U24154 ( .A(n15754), .B(n15830), .Z(n15768) );
  XNOR U24155 ( .A(n15758), .B(n15756), .Z(n15830) );
  XOR U24156 ( .A(n15764), .B(n15831), .Z(n15756) );
  XNOR U24157 ( .A(n15761), .B(n15765), .Z(n15831) );
  AND U24158 ( .A(n15832), .B(n15833), .Z(n15765) );
  NAND U24159 ( .A(n15834), .B(n15835), .Z(n15833) );
  NAND U24160 ( .A(n15836), .B(n15837), .Z(n15832) );
  AND U24161 ( .A(n15838), .B(n15839), .Z(n15761) );
  NAND U24162 ( .A(n15840), .B(n15841), .Z(n15839) );
  NAND U24163 ( .A(n15842), .B(n15843), .Z(n15838) );
  NANDN U24164 ( .A(n15844), .B(n15845), .Z(n15764) );
  ANDN U24165 ( .B(n15846), .A(n15847), .Z(n15758) );
  XNOR U24166 ( .A(n15749), .B(n15848), .Z(n15754) );
  XNOR U24167 ( .A(n15747), .B(n15751), .Z(n15848) );
  AND U24168 ( .A(n15849), .B(n15850), .Z(n15751) );
  NAND U24169 ( .A(n15851), .B(n15852), .Z(n15850) );
  NAND U24170 ( .A(n15853), .B(n15854), .Z(n15849) );
  AND U24171 ( .A(n15855), .B(n15856), .Z(n15747) );
  NAND U24172 ( .A(n15857), .B(n15858), .Z(n15856) );
  NAND U24173 ( .A(n15859), .B(n15860), .Z(n15855) );
  AND U24174 ( .A(n15861), .B(n15862), .Z(n15749) );
  XOR U24175 ( .A(n15829), .B(n15828), .Z(N63985) );
  XNOR U24176 ( .A(n15846), .B(n15847), .Z(n15828) );
  XNOR U24177 ( .A(n15861), .B(n15862), .Z(n15847) );
  XOR U24178 ( .A(n15858), .B(n15857), .Z(n15862) );
  XOR U24179 ( .A(y[6276]), .B(x[6276]), .Z(n15857) );
  XOR U24180 ( .A(n15860), .B(n15859), .Z(n15858) );
  XOR U24181 ( .A(y[6278]), .B(x[6278]), .Z(n15859) );
  XOR U24182 ( .A(y[6277]), .B(x[6277]), .Z(n15860) );
  XOR U24183 ( .A(n15852), .B(n15851), .Z(n15861) );
  XOR U24184 ( .A(n15854), .B(n15853), .Z(n15851) );
  XOR U24185 ( .A(y[6275]), .B(x[6275]), .Z(n15853) );
  XOR U24186 ( .A(y[6274]), .B(x[6274]), .Z(n15854) );
  XOR U24187 ( .A(y[6273]), .B(x[6273]), .Z(n15852) );
  XNOR U24188 ( .A(n15845), .B(n15844), .Z(n15846) );
  XNOR U24189 ( .A(n15841), .B(n15840), .Z(n15844) );
  XOR U24190 ( .A(n15843), .B(n15842), .Z(n15840) );
  XOR U24191 ( .A(y[6272]), .B(x[6272]), .Z(n15842) );
  XOR U24192 ( .A(y[6271]), .B(x[6271]), .Z(n15843) );
  XOR U24193 ( .A(y[6270]), .B(x[6270]), .Z(n15841) );
  XOR U24194 ( .A(n15835), .B(n15834), .Z(n15845) );
  XOR U24195 ( .A(n15837), .B(n15836), .Z(n15834) );
  XOR U24196 ( .A(y[6269]), .B(x[6269]), .Z(n15836) );
  XOR U24197 ( .A(y[6268]), .B(x[6268]), .Z(n15837) );
  XOR U24198 ( .A(y[6267]), .B(x[6267]), .Z(n15835) );
  XNOR U24199 ( .A(n15811), .B(n15812), .Z(n15829) );
  XNOR U24200 ( .A(n15826), .B(n15827), .Z(n15812) );
  XOR U24201 ( .A(n15823), .B(n15822), .Z(n15827) );
  XOR U24202 ( .A(y[6264]), .B(x[6264]), .Z(n15822) );
  XOR U24203 ( .A(n15825), .B(n15824), .Z(n15823) );
  XOR U24204 ( .A(y[6266]), .B(x[6266]), .Z(n15824) );
  XOR U24205 ( .A(y[6265]), .B(x[6265]), .Z(n15825) );
  XOR U24206 ( .A(n15817), .B(n15816), .Z(n15826) );
  XOR U24207 ( .A(n15819), .B(n15818), .Z(n15816) );
  XOR U24208 ( .A(y[6263]), .B(x[6263]), .Z(n15818) );
  XOR U24209 ( .A(y[6262]), .B(x[6262]), .Z(n15819) );
  XOR U24210 ( .A(y[6261]), .B(x[6261]), .Z(n15817) );
  XNOR U24211 ( .A(n15810), .B(n15809), .Z(n15811) );
  XNOR U24212 ( .A(n15806), .B(n15805), .Z(n15809) );
  XOR U24213 ( .A(n15808), .B(n15807), .Z(n15805) );
  XOR U24214 ( .A(y[6260]), .B(x[6260]), .Z(n15807) );
  XOR U24215 ( .A(y[6259]), .B(x[6259]), .Z(n15808) );
  XOR U24216 ( .A(y[6258]), .B(x[6258]), .Z(n15806) );
  XOR U24217 ( .A(n15800), .B(n15799), .Z(n15810) );
  XOR U24218 ( .A(n15802), .B(n15801), .Z(n15799) );
  XOR U24219 ( .A(y[6257]), .B(x[6257]), .Z(n15801) );
  XOR U24220 ( .A(y[6256]), .B(x[6256]), .Z(n15802) );
  XOR U24221 ( .A(y[6255]), .B(x[6255]), .Z(n15800) );
  NAND U24222 ( .A(n15863), .B(n15864), .Z(N63976) );
  NAND U24223 ( .A(n15865), .B(n15866), .Z(n15864) );
  NANDN U24224 ( .A(n15867), .B(n15868), .Z(n15866) );
  NANDN U24225 ( .A(n15868), .B(n15867), .Z(n15863) );
  XOR U24226 ( .A(n15867), .B(n15869), .Z(N63975) );
  XNOR U24227 ( .A(n15865), .B(n15868), .Z(n15869) );
  NAND U24228 ( .A(n15870), .B(n15871), .Z(n15868) );
  NAND U24229 ( .A(n15872), .B(n15873), .Z(n15871) );
  NANDN U24230 ( .A(n15874), .B(n15875), .Z(n15873) );
  NANDN U24231 ( .A(n15875), .B(n15874), .Z(n15870) );
  AND U24232 ( .A(n15876), .B(n15877), .Z(n15865) );
  NAND U24233 ( .A(n15878), .B(n15879), .Z(n15877) );
  NANDN U24234 ( .A(n15880), .B(n15881), .Z(n15879) );
  NANDN U24235 ( .A(n15881), .B(n15880), .Z(n15876) );
  IV U24236 ( .A(n15882), .Z(n15881) );
  AND U24237 ( .A(n15883), .B(n15884), .Z(n15867) );
  NAND U24238 ( .A(n15885), .B(n15886), .Z(n15884) );
  NANDN U24239 ( .A(n15887), .B(n15888), .Z(n15886) );
  NANDN U24240 ( .A(n15888), .B(n15887), .Z(n15883) );
  XOR U24241 ( .A(n15880), .B(n15889), .Z(N63974) );
  XNOR U24242 ( .A(n15878), .B(n15882), .Z(n15889) );
  XOR U24243 ( .A(n15875), .B(n15890), .Z(n15882) );
  XNOR U24244 ( .A(n15872), .B(n15874), .Z(n15890) );
  AND U24245 ( .A(n15891), .B(n15892), .Z(n15874) );
  NANDN U24246 ( .A(n15893), .B(n15894), .Z(n15892) );
  OR U24247 ( .A(n15895), .B(n15896), .Z(n15894) );
  IV U24248 ( .A(n15897), .Z(n15896) );
  NANDN U24249 ( .A(n15897), .B(n15895), .Z(n15891) );
  AND U24250 ( .A(n15898), .B(n15899), .Z(n15872) );
  NAND U24251 ( .A(n15900), .B(n15901), .Z(n15899) );
  NANDN U24252 ( .A(n15902), .B(n15903), .Z(n15901) );
  NANDN U24253 ( .A(n15903), .B(n15902), .Z(n15898) );
  IV U24254 ( .A(n15904), .Z(n15903) );
  NAND U24255 ( .A(n15905), .B(n15906), .Z(n15875) );
  NANDN U24256 ( .A(n15907), .B(n15908), .Z(n15906) );
  NANDN U24257 ( .A(n15909), .B(n15910), .Z(n15908) );
  NANDN U24258 ( .A(n15910), .B(n15909), .Z(n15905) );
  IV U24259 ( .A(n15911), .Z(n15909) );
  AND U24260 ( .A(n15912), .B(n15913), .Z(n15878) );
  NAND U24261 ( .A(n15914), .B(n15915), .Z(n15913) );
  NANDN U24262 ( .A(n15916), .B(n15917), .Z(n15915) );
  NANDN U24263 ( .A(n15917), .B(n15916), .Z(n15912) );
  XOR U24264 ( .A(n15888), .B(n15918), .Z(n15880) );
  XNOR U24265 ( .A(n15885), .B(n15887), .Z(n15918) );
  AND U24266 ( .A(n15919), .B(n15920), .Z(n15887) );
  NANDN U24267 ( .A(n15921), .B(n15922), .Z(n15920) );
  OR U24268 ( .A(n15923), .B(n15924), .Z(n15922) );
  IV U24269 ( .A(n15925), .Z(n15924) );
  NANDN U24270 ( .A(n15925), .B(n15923), .Z(n15919) );
  AND U24271 ( .A(n15926), .B(n15927), .Z(n15885) );
  NAND U24272 ( .A(n15928), .B(n15929), .Z(n15927) );
  NANDN U24273 ( .A(n15930), .B(n15931), .Z(n15929) );
  NANDN U24274 ( .A(n15931), .B(n15930), .Z(n15926) );
  IV U24275 ( .A(n15932), .Z(n15931) );
  NAND U24276 ( .A(n15933), .B(n15934), .Z(n15888) );
  NANDN U24277 ( .A(n15935), .B(n15936), .Z(n15934) );
  NANDN U24278 ( .A(n15937), .B(n15938), .Z(n15936) );
  NANDN U24279 ( .A(n15938), .B(n15937), .Z(n15933) );
  IV U24280 ( .A(n15939), .Z(n15937) );
  XOR U24281 ( .A(n15914), .B(n15940), .Z(N63973) );
  XNOR U24282 ( .A(n15917), .B(n15916), .Z(n15940) );
  XNOR U24283 ( .A(n15928), .B(n15941), .Z(n15916) );
  XNOR U24284 ( .A(n15932), .B(n15930), .Z(n15941) );
  XOR U24285 ( .A(n15938), .B(n15942), .Z(n15930) );
  XNOR U24286 ( .A(n15935), .B(n15939), .Z(n15942) );
  AND U24287 ( .A(n15943), .B(n15944), .Z(n15939) );
  NAND U24288 ( .A(n15945), .B(n15946), .Z(n15944) );
  NAND U24289 ( .A(n15947), .B(n15948), .Z(n15943) );
  AND U24290 ( .A(n15949), .B(n15950), .Z(n15935) );
  NAND U24291 ( .A(n15951), .B(n15952), .Z(n15950) );
  NAND U24292 ( .A(n15953), .B(n15954), .Z(n15949) );
  NANDN U24293 ( .A(n15955), .B(n15956), .Z(n15938) );
  ANDN U24294 ( .B(n15957), .A(n15958), .Z(n15932) );
  XNOR U24295 ( .A(n15923), .B(n15959), .Z(n15928) );
  XNOR U24296 ( .A(n15921), .B(n15925), .Z(n15959) );
  AND U24297 ( .A(n15960), .B(n15961), .Z(n15925) );
  NAND U24298 ( .A(n15962), .B(n15963), .Z(n15961) );
  NAND U24299 ( .A(n15964), .B(n15965), .Z(n15960) );
  AND U24300 ( .A(n15966), .B(n15967), .Z(n15921) );
  NAND U24301 ( .A(n15968), .B(n15969), .Z(n15967) );
  NAND U24302 ( .A(n15970), .B(n15971), .Z(n15966) );
  AND U24303 ( .A(n15972), .B(n15973), .Z(n15923) );
  NAND U24304 ( .A(n15974), .B(n15975), .Z(n15917) );
  XNOR U24305 ( .A(n15900), .B(n15976), .Z(n15914) );
  XNOR U24306 ( .A(n15904), .B(n15902), .Z(n15976) );
  XOR U24307 ( .A(n15910), .B(n15977), .Z(n15902) );
  XNOR U24308 ( .A(n15907), .B(n15911), .Z(n15977) );
  AND U24309 ( .A(n15978), .B(n15979), .Z(n15911) );
  NAND U24310 ( .A(n15980), .B(n15981), .Z(n15979) );
  NAND U24311 ( .A(n15982), .B(n15983), .Z(n15978) );
  AND U24312 ( .A(n15984), .B(n15985), .Z(n15907) );
  NAND U24313 ( .A(n15986), .B(n15987), .Z(n15985) );
  NAND U24314 ( .A(n15988), .B(n15989), .Z(n15984) );
  NANDN U24315 ( .A(n15990), .B(n15991), .Z(n15910) );
  ANDN U24316 ( .B(n15992), .A(n15993), .Z(n15904) );
  XNOR U24317 ( .A(n15895), .B(n15994), .Z(n15900) );
  XNOR U24318 ( .A(n15893), .B(n15897), .Z(n15994) );
  AND U24319 ( .A(n15995), .B(n15996), .Z(n15897) );
  NAND U24320 ( .A(n15997), .B(n15998), .Z(n15996) );
  NAND U24321 ( .A(n15999), .B(n16000), .Z(n15995) );
  AND U24322 ( .A(n16001), .B(n16002), .Z(n15893) );
  NAND U24323 ( .A(n16003), .B(n16004), .Z(n16002) );
  NAND U24324 ( .A(n16005), .B(n16006), .Z(n16001) );
  AND U24325 ( .A(n16007), .B(n16008), .Z(n15895) );
  XOR U24326 ( .A(n15975), .B(n15974), .Z(N63972) );
  XNOR U24327 ( .A(n15992), .B(n15993), .Z(n15974) );
  XNOR U24328 ( .A(n16007), .B(n16008), .Z(n15993) );
  XOR U24329 ( .A(n16004), .B(n16003), .Z(n16008) );
  XOR U24330 ( .A(y[6252]), .B(x[6252]), .Z(n16003) );
  XOR U24331 ( .A(n16006), .B(n16005), .Z(n16004) );
  XOR U24332 ( .A(y[6254]), .B(x[6254]), .Z(n16005) );
  XOR U24333 ( .A(y[6253]), .B(x[6253]), .Z(n16006) );
  XOR U24334 ( .A(n15998), .B(n15997), .Z(n16007) );
  XOR U24335 ( .A(n16000), .B(n15999), .Z(n15997) );
  XOR U24336 ( .A(y[6251]), .B(x[6251]), .Z(n15999) );
  XOR U24337 ( .A(y[6250]), .B(x[6250]), .Z(n16000) );
  XOR U24338 ( .A(y[6249]), .B(x[6249]), .Z(n15998) );
  XNOR U24339 ( .A(n15991), .B(n15990), .Z(n15992) );
  XNOR U24340 ( .A(n15987), .B(n15986), .Z(n15990) );
  XOR U24341 ( .A(n15989), .B(n15988), .Z(n15986) );
  XOR U24342 ( .A(y[6248]), .B(x[6248]), .Z(n15988) );
  XOR U24343 ( .A(y[6247]), .B(x[6247]), .Z(n15989) );
  XOR U24344 ( .A(y[6246]), .B(x[6246]), .Z(n15987) );
  XOR U24345 ( .A(n15981), .B(n15980), .Z(n15991) );
  XOR U24346 ( .A(n15983), .B(n15982), .Z(n15980) );
  XOR U24347 ( .A(y[6245]), .B(x[6245]), .Z(n15982) );
  XOR U24348 ( .A(y[6244]), .B(x[6244]), .Z(n15983) );
  XOR U24349 ( .A(y[6243]), .B(x[6243]), .Z(n15981) );
  XNOR U24350 ( .A(n15957), .B(n15958), .Z(n15975) );
  XNOR U24351 ( .A(n15972), .B(n15973), .Z(n15958) );
  XOR U24352 ( .A(n15969), .B(n15968), .Z(n15973) );
  XOR U24353 ( .A(y[6240]), .B(x[6240]), .Z(n15968) );
  XOR U24354 ( .A(n15971), .B(n15970), .Z(n15969) );
  XOR U24355 ( .A(y[6242]), .B(x[6242]), .Z(n15970) );
  XOR U24356 ( .A(y[6241]), .B(x[6241]), .Z(n15971) );
  XOR U24357 ( .A(n15963), .B(n15962), .Z(n15972) );
  XOR U24358 ( .A(n15965), .B(n15964), .Z(n15962) );
  XOR U24359 ( .A(y[6239]), .B(x[6239]), .Z(n15964) );
  XOR U24360 ( .A(y[6238]), .B(x[6238]), .Z(n15965) );
  XOR U24361 ( .A(y[6237]), .B(x[6237]), .Z(n15963) );
  XNOR U24362 ( .A(n15956), .B(n15955), .Z(n15957) );
  XNOR U24363 ( .A(n15952), .B(n15951), .Z(n15955) );
  XOR U24364 ( .A(n15954), .B(n15953), .Z(n15951) );
  XOR U24365 ( .A(y[6236]), .B(x[6236]), .Z(n15953) );
  XOR U24366 ( .A(y[6235]), .B(x[6235]), .Z(n15954) );
  XOR U24367 ( .A(y[6234]), .B(x[6234]), .Z(n15952) );
  XOR U24368 ( .A(n15946), .B(n15945), .Z(n15956) );
  XOR U24369 ( .A(n15948), .B(n15947), .Z(n15945) );
  XOR U24370 ( .A(y[6233]), .B(x[6233]), .Z(n15947) );
  XOR U24371 ( .A(y[6232]), .B(x[6232]), .Z(n15948) );
  XOR U24372 ( .A(y[6231]), .B(x[6231]), .Z(n15946) );
  NAND U24373 ( .A(n16009), .B(n16010), .Z(N63963) );
  NAND U24374 ( .A(n16011), .B(n16012), .Z(n16010) );
  NANDN U24375 ( .A(n16013), .B(n16014), .Z(n16012) );
  NANDN U24376 ( .A(n16014), .B(n16013), .Z(n16009) );
  XOR U24377 ( .A(n16013), .B(n16015), .Z(N63962) );
  XNOR U24378 ( .A(n16011), .B(n16014), .Z(n16015) );
  NAND U24379 ( .A(n16016), .B(n16017), .Z(n16014) );
  NAND U24380 ( .A(n16018), .B(n16019), .Z(n16017) );
  NANDN U24381 ( .A(n16020), .B(n16021), .Z(n16019) );
  NANDN U24382 ( .A(n16021), .B(n16020), .Z(n16016) );
  AND U24383 ( .A(n16022), .B(n16023), .Z(n16011) );
  NAND U24384 ( .A(n16024), .B(n16025), .Z(n16023) );
  NANDN U24385 ( .A(n16026), .B(n16027), .Z(n16025) );
  NANDN U24386 ( .A(n16027), .B(n16026), .Z(n16022) );
  IV U24387 ( .A(n16028), .Z(n16027) );
  AND U24388 ( .A(n16029), .B(n16030), .Z(n16013) );
  NAND U24389 ( .A(n16031), .B(n16032), .Z(n16030) );
  NANDN U24390 ( .A(n16033), .B(n16034), .Z(n16032) );
  NANDN U24391 ( .A(n16034), .B(n16033), .Z(n16029) );
  XOR U24392 ( .A(n16026), .B(n16035), .Z(N63961) );
  XNOR U24393 ( .A(n16024), .B(n16028), .Z(n16035) );
  XOR U24394 ( .A(n16021), .B(n16036), .Z(n16028) );
  XNOR U24395 ( .A(n16018), .B(n16020), .Z(n16036) );
  AND U24396 ( .A(n16037), .B(n16038), .Z(n16020) );
  NANDN U24397 ( .A(n16039), .B(n16040), .Z(n16038) );
  OR U24398 ( .A(n16041), .B(n16042), .Z(n16040) );
  IV U24399 ( .A(n16043), .Z(n16042) );
  NANDN U24400 ( .A(n16043), .B(n16041), .Z(n16037) );
  AND U24401 ( .A(n16044), .B(n16045), .Z(n16018) );
  NAND U24402 ( .A(n16046), .B(n16047), .Z(n16045) );
  NANDN U24403 ( .A(n16048), .B(n16049), .Z(n16047) );
  NANDN U24404 ( .A(n16049), .B(n16048), .Z(n16044) );
  IV U24405 ( .A(n16050), .Z(n16049) );
  NAND U24406 ( .A(n16051), .B(n16052), .Z(n16021) );
  NANDN U24407 ( .A(n16053), .B(n16054), .Z(n16052) );
  NANDN U24408 ( .A(n16055), .B(n16056), .Z(n16054) );
  NANDN U24409 ( .A(n16056), .B(n16055), .Z(n16051) );
  IV U24410 ( .A(n16057), .Z(n16055) );
  AND U24411 ( .A(n16058), .B(n16059), .Z(n16024) );
  NAND U24412 ( .A(n16060), .B(n16061), .Z(n16059) );
  NANDN U24413 ( .A(n16062), .B(n16063), .Z(n16061) );
  NANDN U24414 ( .A(n16063), .B(n16062), .Z(n16058) );
  XOR U24415 ( .A(n16034), .B(n16064), .Z(n16026) );
  XNOR U24416 ( .A(n16031), .B(n16033), .Z(n16064) );
  AND U24417 ( .A(n16065), .B(n16066), .Z(n16033) );
  NANDN U24418 ( .A(n16067), .B(n16068), .Z(n16066) );
  OR U24419 ( .A(n16069), .B(n16070), .Z(n16068) );
  IV U24420 ( .A(n16071), .Z(n16070) );
  NANDN U24421 ( .A(n16071), .B(n16069), .Z(n16065) );
  AND U24422 ( .A(n16072), .B(n16073), .Z(n16031) );
  NAND U24423 ( .A(n16074), .B(n16075), .Z(n16073) );
  NANDN U24424 ( .A(n16076), .B(n16077), .Z(n16075) );
  NANDN U24425 ( .A(n16077), .B(n16076), .Z(n16072) );
  IV U24426 ( .A(n16078), .Z(n16077) );
  NAND U24427 ( .A(n16079), .B(n16080), .Z(n16034) );
  NANDN U24428 ( .A(n16081), .B(n16082), .Z(n16080) );
  NANDN U24429 ( .A(n16083), .B(n16084), .Z(n16082) );
  NANDN U24430 ( .A(n16084), .B(n16083), .Z(n16079) );
  IV U24431 ( .A(n16085), .Z(n16083) );
  XOR U24432 ( .A(n16060), .B(n16086), .Z(N63960) );
  XNOR U24433 ( .A(n16063), .B(n16062), .Z(n16086) );
  XNOR U24434 ( .A(n16074), .B(n16087), .Z(n16062) );
  XNOR U24435 ( .A(n16078), .B(n16076), .Z(n16087) );
  XOR U24436 ( .A(n16084), .B(n16088), .Z(n16076) );
  XNOR U24437 ( .A(n16081), .B(n16085), .Z(n16088) );
  AND U24438 ( .A(n16089), .B(n16090), .Z(n16085) );
  NAND U24439 ( .A(n16091), .B(n16092), .Z(n16090) );
  NAND U24440 ( .A(n16093), .B(n16094), .Z(n16089) );
  AND U24441 ( .A(n16095), .B(n16096), .Z(n16081) );
  NAND U24442 ( .A(n16097), .B(n16098), .Z(n16096) );
  NAND U24443 ( .A(n16099), .B(n16100), .Z(n16095) );
  NANDN U24444 ( .A(n16101), .B(n16102), .Z(n16084) );
  ANDN U24445 ( .B(n16103), .A(n16104), .Z(n16078) );
  XNOR U24446 ( .A(n16069), .B(n16105), .Z(n16074) );
  XNOR U24447 ( .A(n16067), .B(n16071), .Z(n16105) );
  AND U24448 ( .A(n16106), .B(n16107), .Z(n16071) );
  NAND U24449 ( .A(n16108), .B(n16109), .Z(n16107) );
  NAND U24450 ( .A(n16110), .B(n16111), .Z(n16106) );
  AND U24451 ( .A(n16112), .B(n16113), .Z(n16067) );
  NAND U24452 ( .A(n16114), .B(n16115), .Z(n16113) );
  NAND U24453 ( .A(n16116), .B(n16117), .Z(n16112) );
  AND U24454 ( .A(n16118), .B(n16119), .Z(n16069) );
  NAND U24455 ( .A(n16120), .B(n16121), .Z(n16063) );
  XNOR U24456 ( .A(n16046), .B(n16122), .Z(n16060) );
  XNOR U24457 ( .A(n16050), .B(n16048), .Z(n16122) );
  XOR U24458 ( .A(n16056), .B(n16123), .Z(n16048) );
  XNOR U24459 ( .A(n16053), .B(n16057), .Z(n16123) );
  AND U24460 ( .A(n16124), .B(n16125), .Z(n16057) );
  NAND U24461 ( .A(n16126), .B(n16127), .Z(n16125) );
  NAND U24462 ( .A(n16128), .B(n16129), .Z(n16124) );
  AND U24463 ( .A(n16130), .B(n16131), .Z(n16053) );
  NAND U24464 ( .A(n16132), .B(n16133), .Z(n16131) );
  NAND U24465 ( .A(n16134), .B(n16135), .Z(n16130) );
  NANDN U24466 ( .A(n16136), .B(n16137), .Z(n16056) );
  ANDN U24467 ( .B(n16138), .A(n16139), .Z(n16050) );
  XNOR U24468 ( .A(n16041), .B(n16140), .Z(n16046) );
  XNOR U24469 ( .A(n16039), .B(n16043), .Z(n16140) );
  AND U24470 ( .A(n16141), .B(n16142), .Z(n16043) );
  NAND U24471 ( .A(n16143), .B(n16144), .Z(n16142) );
  NAND U24472 ( .A(n16145), .B(n16146), .Z(n16141) );
  AND U24473 ( .A(n16147), .B(n16148), .Z(n16039) );
  NAND U24474 ( .A(n16149), .B(n16150), .Z(n16148) );
  NAND U24475 ( .A(n16151), .B(n16152), .Z(n16147) );
  AND U24476 ( .A(n16153), .B(n16154), .Z(n16041) );
  XOR U24477 ( .A(n16121), .B(n16120), .Z(N63959) );
  XNOR U24478 ( .A(n16138), .B(n16139), .Z(n16120) );
  XNOR U24479 ( .A(n16153), .B(n16154), .Z(n16139) );
  XOR U24480 ( .A(n16150), .B(n16149), .Z(n16154) );
  XOR U24481 ( .A(y[6228]), .B(x[6228]), .Z(n16149) );
  XOR U24482 ( .A(n16152), .B(n16151), .Z(n16150) );
  XOR U24483 ( .A(y[6230]), .B(x[6230]), .Z(n16151) );
  XOR U24484 ( .A(y[6229]), .B(x[6229]), .Z(n16152) );
  XOR U24485 ( .A(n16144), .B(n16143), .Z(n16153) );
  XOR U24486 ( .A(n16146), .B(n16145), .Z(n16143) );
  XOR U24487 ( .A(y[6227]), .B(x[6227]), .Z(n16145) );
  XOR U24488 ( .A(y[6226]), .B(x[6226]), .Z(n16146) );
  XOR U24489 ( .A(y[6225]), .B(x[6225]), .Z(n16144) );
  XNOR U24490 ( .A(n16137), .B(n16136), .Z(n16138) );
  XNOR U24491 ( .A(n16133), .B(n16132), .Z(n16136) );
  XOR U24492 ( .A(n16135), .B(n16134), .Z(n16132) );
  XOR U24493 ( .A(y[6224]), .B(x[6224]), .Z(n16134) );
  XOR U24494 ( .A(y[6223]), .B(x[6223]), .Z(n16135) );
  XOR U24495 ( .A(y[6222]), .B(x[6222]), .Z(n16133) );
  XOR U24496 ( .A(n16127), .B(n16126), .Z(n16137) );
  XOR U24497 ( .A(n16129), .B(n16128), .Z(n16126) );
  XOR U24498 ( .A(y[6221]), .B(x[6221]), .Z(n16128) );
  XOR U24499 ( .A(y[6220]), .B(x[6220]), .Z(n16129) );
  XOR U24500 ( .A(y[6219]), .B(x[6219]), .Z(n16127) );
  XNOR U24501 ( .A(n16103), .B(n16104), .Z(n16121) );
  XNOR U24502 ( .A(n16118), .B(n16119), .Z(n16104) );
  XOR U24503 ( .A(n16115), .B(n16114), .Z(n16119) );
  XOR U24504 ( .A(y[6216]), .B(x[6216]), .Z(n16114) );
  XOR U24505 ( .A(n16117), .B(n16116), .Z(n16115) );
  XOR U24506 ( .A(y[6218]), .B(x[6218]), .Z(n16116) );
  XOR U24507 ( .A(y[6217]), .B(x[6217]), .Z(n16117) );
  XOR U24508 ( .A(n16109), .B(n16108), .Z(n16118) );
  XOR U24509 ( .A(n16111), .B(n16110), .Z(n16108) );
  XOR U24510 ( .A(y[6215]), .B(x[6215]), .Z(n16110) );
  XOR U24511 ( .A(y[6214]), .B(x[6214]), .Z(n16111) );
  XOR U24512 ( .A(y[6213]), .B(x[6213]), .Z(n16109) );
  XNOR U24513 ( .A(n16102), .B(n16101), .Z(n16103) );
  XNOR U24514 ( .A(n16098), .B(n16097), .Z(n16101) );
  XOR U24515 ( .A(n16100), .B(n16099), .Z(n16097) );
  XOR U24516 ( .A(y[6212]), .B(x[6212]), .Z(n16099) );
  XOR U24517 ( .A(y[6211]), .B(x[6211]), .Z(n16100) );
  XOR U24518 ( .A(y[6210]), .B(x[6210]), .Z(n16098) );
  XOR U24519 ( .A(n16092), .B(n16091), .Z(n16102) );
  XOR U24520 ( .A(n16094), .B(n16093), .Z(n16091) );
  XOR U24521 ( .A(y[6209]), .B(x[6209]), .Z(n16093) );
  XOR U24522 ( .A(y[6208]), .B(x[6208]), .Z(n16094) );
  XOR U24523 ( .A(y[6207]), .B(x[6207]), .Z(n16092) );
  NAND U24524 ( .A(n16155), .B(n16156), .Z(N63950) );
  NAND U24525 ( .A(n16157), .B(n16158), .Z(n16156) );
  NANDN U24526 ( .A(n16159), .B(n16160), .Z(n16158) );
  NANDN U24527 ( .A(n16160), .B(n16159), .Z(n16155) );
  XOR U24528 ( .A(n16159), .B(n16161), .Z(N63949) );
  XNOR U24529 ( .A(n16157), .B(n16160), .Z(n16161) );
  NAND U24530 ( .A(n16162), .B(n16163), .Z(n16160) );
  NAND U24531 ( .A(n16164), .B(n16165), .Z(n16163) );
  NANDN U24532 ( .A(n16166), .B(n16167), .Z(n16165) );
  NANDN U24533 ( .A(n16167), .B(n16166), .Z(n16162) );
  AND U24534 ( .A(n16168), .B(n16169), .Z(n16157) );
  NAND U24535 ( .A(n16170), .B(n16171), .Z(n16169) );
  NANDN U24536 ( .A(n16172), .B(n16173), .Z(n16171) );
  NANDN U24537 ( .A(n16173), .B(n16172), .Z(n16168) );
  IV U24538 ( .A(n16174), .Z(n16173) );
  AND U24539 ( .A(n16175), .B(n16176), .Z(n16159) );
  NAND U24540 ( .A(n16177), .B(n16178), .Z(n16176) );
  NANDN U24541 ( .A(n16179), .B(n16180), .Z(n16178) );
  NANDN U24542 ( .A(n16180), .B(n16179), .Z(n16175) );
  XOR U24543 ( .A(n16172), .B(n16181), .Z(N63948) );
  XNOR U24544 ( .A(n16170), .B(n16174), .Z(n16181) );
  XOR U24545 ( .A(n16167), .B(n16182), .Z(n16174) );
  XNOR U24546 ( .A(n16164), .B(n16166), .Z(n16182) );
  AND U24547 ( .A(n16183), .B(n16184), .Z(n16166) );
  NANDN U24548 ( .A(n16185), .B(n16186), .Z(n16184) );
  OR U24549 ( .A(n16187), .B(n16188), .Z(n16186) );
  IV U24550 ( .A(n16189), .Z(n16188) );
  NANDN U24551 ( .A(n16189), .B(n16187), .Z(n16183) );
  AND U24552 ( .A(n16190), .B(n16191), .Z(n16164) );
  NAND U24553 ( .A(n16192), .B(n16193), .Z(n16191) );
  NANDN U24554 ( .A(n16194), .B(n16195), .Z(n16193) );
  NANDN U24555 ( .A(n16195), .B(n16194), .Z(n16190) );
  IV U24556 ( .A(n16196), .Z(n16195) );
  NAND U24557 ( .A(n16197), .B(n16198), .Z(n16167) );
  NANDN U24558 ( .A(n16199), .B(n16200), .Z(n16198) );
  NANDN U24559 ( .A(n16201), .B(n16202), .Z(n16200) );
  NANDN U24560 ( .A(n16202), .B(n16201), .Z(n16197) );
  IV U24561 ( .A(n16203), .Z(n16201) );
  AND U24562 ( .A(n16204), .B(n16205), .Z(n16170) );
  NAND U24563 ( .A(n16206), .B(n16207), .Z(n16205) );
  NANDN U24564 ( .A(n16208), .B(n16209), .Z(n16207) );
  NANDN U24565 ( .A(n16209), .B(n16208), .Z(n16204) );
  XOR U24566 ( .A(n16180), .B(n16210), .Z(n16172) );
  XNOR U24567 ( .A(n16177), .B(n16179), .Z(n16210) );
  AND U24568 ( .A(n16211), .B(n16212), .Z(n16179) );
  NANDN U24569 ( .A(n16213), .B(n16214), .Z(n16212) );
  OR U24570 ( .A(n16215), .B(n16216), .Z(n16214) );
  IV U24571 ( .A(n16217), .Z(n16216) );
  NANDN U24572 ( .A(n16217), .B(n16215), .Z(n16211) );
  AND U24573 ( .A(n16218), .B(n16219), .Z(n16177) );
  NAND U24574 ( .A(n16220), .B(n16221), .Z(n16219) );
  NANDN U24575 ( .A(n16222), .B(n16223), .Z(n16221) );
  NANDN U24576 ( .A(n16223), .B(n16222), .Z(n16218) );
  IV U24577 ( .A(n16224), .Z(n16223) );
  NAND U24578 ( .A(n16225), .B(n16226), .Z(n16180) );
  NANDN U24579 ( .A(n16227), .B(n16228), .Z(n16226) );
  NANDN U24580 ( .A(n16229), .B(n16230), .Z(n16228) );
  NANDN U24581 ( .A(n16230), .B(n16229), .Z(n16225) );
  IV U24582 ( .A(n16231), .Z(n16229) );
  XOR U24583 ( .A(n16206), .B(n16232), .Z(N63947) );
  XNOR U24584 ( .A(n16209), .B(n16208), .Z(n16232) );
  XNOR U24585 ( .A(n16220), .B(n16233), .Z(n16208) );
  XNOR U24586 ( .A(n16224), .B(n16222), .Z(n16233) );
  XOR U24587 ( .A(n16230), .B(n16234), .Z(n16222) );
  XNOR U24588 ( .A(n16227), .B(n16231), .Z(n16234) );
  AND U24589 ( .A(n16235), .B(n16236), .Z(n16231) );
  NAND U24590 ( .A(n16237), .B(n16238), .Z(n16236) );
  NAND U24591 ( .A(n16239), .B(n16240), .Z(n16235) );
  AND U24592 ( .A(n16241), .B(n16242), .Z(n16227) );
  NAND U24593 ( .A(n16243), .B(n16244), .Z(n16242) );
  NAND U24594 ( .A(n16245), .B(n16246), .Z(n16241) );
  NANDN U24595 ( .A(n16247), .B(n16248), .Z(n16230) );
  ANDN U24596 ( .B(n16249), .A(n16250), .Z(n16224) );
  XNOR U24597 ( .A(n16215), .B(n16251), .Z(n16220) );
  XNOR U24598 ( .A(n16213), .B(n16217), .Z(n16251) );
  AND U24599 ( .A(n16252), .B(n16253), .Z(n16217) );
  NAND U24600 ( .A(n16254), .B(n16255), .Z(n16253) );
  NAND U24601 ( .A(n16256), .B(n16257), .Z(n16252) );
  AND U24602 ( .A(n16258), .B(n16259), .Z(n16213) );
  NAND U24603 ( .A(n16260), .B(n16261), .Z(n16259) );
  NAND U24604 ( .A(n16262), .B(n16263), .Z(n16258) );
  AND U24605 ( .A(n16264), .B(n16265), .Z(n16215) );
  NAND U24606 ( .A(n16266), .B(n16267), .Z(n16209) );
  XNOR U24607 ( .A(n16192), .B(n16268), .Z(n16206) );
  XNOR U24608 ( .A(n16196), .B(n16194), .Z(n16268) );
  XOR U24609 ( .A(n16202), .B(n16269), .Z(n16194) );
  XNOR U24610 ( .A(n16199), .B(n16203), .Z(n16269) );
  AND U24611 ( .A(n16270), .B(n16271), .Z(n16203) );
  NAND U24612 ( .A(n16272), .B(n16273), .Z(n16271) );
  NAND U24613 ( .A(n16274), .B(n16275), .Z(n16270) );
  AND U24614 ( .A(n16276), .B(n16277), .Z(n16199) );
  NAND U24615 ( .A(n16278), .B(n16279), .Z(n16277) );
  NAND U24616 ( .A(n16280), .B(n16281), .Z(n16276) );
  NANDN U24617 ( .A(n16282), .B(n16283), .Z(n16202) );
  ANDN U24618 ( .B(n16284), .A(n16285), .Z(n16196) );
  XNOR U24619 ( .A(n16187), .B(n16286), .Z(n16192) );
  XNOR U24620 ( .A(n16185), .B(n16189), .Z(n16286) );
  AND U24621 ( .A(n16287), .B(n16288), .Z(n16189) );
  NAND U24622 ( .A(n16289), .B(n16290), .Z(n16288) );
  NAND U24623 ( .A(n16291), .B(n16292), .Z(n16287) );
  AND U24624 ( .A(n16293), .B(n16294), .Z(n16185) );
  NAND U24625 ( .A(n16295), .B(n16296), .Z(n16294) );
  NAND U24626 ( .A(n16297), .B(n16298), .Z(n16293) );
  AND U24627 ( .A(n16299), .B(n16300), .Z(n16187) );
  XOR U24628 ( .A(n16267), .B(n16266), .Z(N63946) );
  XNOR U24629 ( .A(n16284), .B(n16285), .Z(n16266) );
  XNOR U24630 ( .A(n16299), .B(n16300), .Z(n16285) );
  XOR U24631 ( .A(n16296), .B(n16295), .Z(n16300) );
  XOR U24632 ( .A(y[6204]), .B(x[6204]), .Z(n16295) );
  XOR U24633 ( .A(n16298), .B(n16297), .Z(n16296) );
  XOR U24634 ( .A(y[6206]), .B(x[6206]), .Z(n16297) );
  XOR U24635 ( .A(y[6205]), .B(x[6205]), .Z(n16298) );
  XOR U24636 ( .A(n16290), .B(n16289), .Z(n16299) );
  XOR U24637 ( .A(n16292), .B(n16291), .Z(n16289) );
  XOR U24638 ( .A(y[6203]), .B(x[6203]), .Z(n16291) );
  XOR U24639 ( .A(y[6202]), .B(x[6202]), .Z(n16292) );
  XOR U24640 ( .A(y[6201]), .B(x[6201]), .Z(n16290) );
  XNOR U24641 ( .A(n16283), .B(n16282), .Z(n16284) );
  XNOR U24642 ( .A(n16279), .B(n16278), .Z(n16282) );
  XOR U24643 ( .A(n16281), .B(n16280), .Z(n16278) );
  XOR U24644 ( .A(y[6200]), .B(x[6200]), .Z(n16280) );
  XOR U24645 ( .A(y[6199]), .B(x[6199]), .Z(n16281) );
  XOR U24646 ( .A(y[6198]), .B(x[6198]), .Z(n16279) );
  XOR U24647 ( .A(n16273), .B(n16272), .Z(n16283) );
  XOR U24648 ( .A(n16275), .B(n16274), .Z(n16272) );
  XOR U24649 ( .A(y[6197]), .B(x[6197]), .Z(n16274) );
  XOR U24650 ( .A(y[6196]), .B(x[6196]), .Z(n16275) );
  XOR U24651 ( .A(y[6195]), .B(x[6195]), .Z(n16273) );
  XNOR U24652 ( .A(n16249), .B(n16250), .Z(n16267) );
  XNOR U24653 ( .A(n16264), .B(n16265), .Z(n16250) );
  XOR U24654 ( .A(n16261), .B(n16260), .Z(n16265) );
  XOR U24655 ( .A(y[6192]), .B(x[6192]), .Z(n16260) );
  XOR U24656 ( .A(n16263), .B(n16262), .Z(n16261) );
  XOR U24657 ( .A(y[6194]), .B(x[6194]), .Z(n16262) );
  XOR U24658 ( .A(y[6193]), .B(x[6193]), .Z(n16263) );
  XOR U24659 ( .A(n16255), .B(n16254), .Z(n16264) );
  XOR U24660 ( .A(n16257), .B(n16256), .Z(n16254) );
  XOR U24661 ( .A(y[6191]), .B(x[6191]), .Z(n16256) );
  XOR U24662 ( .A(y[6190]), .B(x[6190]), .Z(n16257) );
  XOR U24663 ( .A(y[6189]), .B(x[6189]), .Z(n16255) );
  XNOR U24664 ( .A(n16248), .B(n16247), .Z(n16249) );
  XNOR U24665 ( .A(n16244), .B(n16243), .Z(n16247) );
  XOR U24666 ( .A(n16246), .B(n16245), .Z(n16243) );
  XOR U24667 ( .A(y[6188]), .B(x[6188]), .Z(n16245) );
  XOR U24668 ( .A(y[6187]), .B(x[6187]), .Z(n16246) );
  XOR U24669 ( .A(y[6186]), .B(x[6186]), .Z(n16244) );
  XOR U24670 ( .A(n16238), .B(n16237), .Z(n16248) );
  XOR U24671 ( .A(n16240), .B(n16239), .Z(n16237) );
  XOR U24672 ( .A(y[6185]), .B(x[6185]), .Z(n16239) );
  XOR U24673 ( .A(y[6184]), .B(x[6184]), .Z(n16240) );
  XOR U24674 ( .A(y[6183]), .B(x[6183]), .Z(n16238) );
  NAND U24675 ( .A(n16301), .B(n16302), .Z(N63937) );
  NAND U24676 ( .A(n16303), .B(n16304), .Z(n16302) );
  NANDN U24677 ( .A(n16305), .B(n16306), .Z(n16304) );
  NANDN U24678 ( .A(n16306), .B(n16305), .Z(n16301) );
  XOR U24679 ( .A(n16305), .B(n16307), .Z(N63936) );
  XNOR U24680 ( .A(n16303), .B(n16306), .Z(n16307) );
  NAND U24681 ( .A(n16308), .B(n16309), .Z(n16306) );
  NAND U24682 ( .A(n16310), .B(n16311), .Z(n16309) );
  NANDN U24683 ( .A(n16312), .B(n16313), .Z(n16311) );
  NANDN U24684 ( .A(n16313), .B(n16312), .Z(n16308) );
  AND U24685 ( .A(n16314), .B(n16315), .Z(n16303) );
  NAND U24686 ( .A(n16316), .B(n16317), .Z(n16315) );
  NANDN U24687 ( .A(n16318), .B(n16319), .Z(n16317) );
  NANDN U24688 ( .A(n16319), .B(n16318), .Z(n16314) );
  IV U24689 ( .A(n16320), .Z(n16319) );
  AND U24690 ( .A(n16321), .B(n16322), .Z(n16305) );
  NAND U24691 ( .A(n16323), .B(n16324), .Z(n16322) );
  NANDN U24692 ( .A(n16325), .B(n16326), .Z(n16324) );
  NANDN U24693 ( .A(n16326), .B(n16325), .Z(n16321) );
  XOR U24694 ( .A(n16318), .B(n16327), .Z(N63935) );
  XNOR U24695 ( .A(n16316), .B(n16320), .Z(n16327) );
  XOR U24696 ( .A(n16313), .B(n16328), .Z(n16320) );
  XNOR U24697 ( .A(n16310), .B(n16312), .Z(n16328) );
  AND U24698 ( .A(n16329), .B(n16330), .Z(n16312) );
  NANDN U24699 ( .A(n16331), .B(n16332), .Z(n16330) );
  OR U24700 ( .A(n16333), .B(n16334), .Z(n16332) );
  IV U24701 ( .A(n16335), .Z(n16334) );
  NANDN U24702 ( .A(n16335), .B(n16333), .Z(n16329) );
  AND U24703 ( .A(n16336), .B(n16337), .Z(n16310) );
  NAND U24704 ( .A(n16338), .B(n16339), .Z(n16337) );
  NANDN U24705 ( .A(n16340), .B(n16341), .Z(n16339) );
  NANDN U24706 ( .A(n16341), .B(n16340), .Z(n16336) );
  IV U24707 ( .A(n16342), .Z(n16341) );
  NAND U24708 ( .A(n16343), .B(n16344), .Z(n16313) );
  NANDN U24709 ( .A(n16345), .B(n16346), .Z(n16344) );
  NANDN U24710 ( .A(n16347), .B(n16348), .Z(n16346) );
  NANDN U24711 ( .A(n16348), .B(n16347), .Z(n16343) );
  IV U24712 ( .A(n16349), .Z(n16347) );
  AND U24713 ( .A(n16350), .B(n16351), .Z(n16316) );
  NAND U24714 ( .A(n16352), .B(n16353), .Z(n16351) );
  NANDN U24715 ( .A(n16354), .B(n16355), .Z(n16353) );
  NANDN U24716 ( .A(n16355), .B(n16354), .Z(n16350) );
  XOR U24717 ( .A(n16326), .B(n16356), .Z(n16318) );
  XNOR U24718 ( .A(n16323), .B(n16325), .Z(n16356) );
  AND U24719 ( .A(n16357), .B(n16358), .Z(n16325) );
  NANDN U24720 ( .A(n16359), .B(n16360), .Z(n16358) );
  OR U24721 ( .A(n16361), .B(n16362), .Z(n16360) );
  IV U24722 ( .A(n16363), .Z(n16362) );
  NANDN U24723 ( .A(n16363), .B(n16361), .Z(n16357) );
  AND U24724 ( .A(n16364), .B(n16365), .Z(n16323) );
  NAND U24725 ( .A(n16366), .B(n16367), .Z(n16365) );
  NANDN U24726 ( .A(n16368), .B(n16369), .Z(n16367) );
  NANDN U24727 ( .A(n16369), .B(n16368), .Z(n16364) );
  IV U24728 ( .A(n16370), .Z(n16369) );
  NAND U24729 ( .A(n16371), .B(n16372), .Z(n16326) );
  NANDN U24730 ( .A(n16373), .B(n16374), .Z(n16372) );
  NANDN U24731 ( .A(n16375), .B(n16376), .Z(n16374) );
  NANDN U24732 ( .A(n16376), .B(n16375), .Z(n16371) );
  IV U24733 ( .A(n16377), .Z(n16375) );
  XOR U24734 ( .A(n16352), .B(n16378), .Z(N63934) );
  XNOR U24735 ( .A(n16355), .B(n16354), .Z(n16378) );
  XNOR U24736 ( .A(n16366), .B(n16379), .Z(n16354) );
  XNOR U24737 ( .A(n16370), .B(n16368), .Z(n16379) );
  XOR U24738 ( .A(n16376), .B(n16380), .Z(n16368) );
  XNOR U24739 ( .A(n16373), .B(n16377), .Z(n16380) );
  AND U24740 ( .A(n16381), .B(n16382), .Z(n16377) );
  NAND U24741 ( .A(n16383), .B(n16384), .Z(n16382) );
  NAND U24742 ( .A(n16385), .B(n16386), .Z(n16381) );
  AND U24743 ( .A(n16387), .B(n16388), .Z(n16373) );
  NAND U24744 ( .A(n16389), .B(n16390), .Z(n16388) );
  NAND U24745 ( .A(n16391), .B(n16392), .Z(n16387) );
  NANDN U24746 ( .A(n16393), .B(n16394), .Z(n16376) );
  ANDN U24747 ( .B(n16395), .A(n16396), .Z(n16370) );
  XNOR U24748 ( .A(n16361), .B(n16397), .Z(n16366) );
  XNOR U24749 ( .A(n16359), .B(n16363), .Z(n16397) );
  AND U24750 ( .A(n16398), .B(n16399), .Z(n16363) );
  NAND U24751 ( .A(n16400), .B(n16401), .Z(n16399) );
  NAND U24752 ( .A(n16402), .B(n16403), .Z(n16398) );
  AND U24753 ( .A(n16404), .B(n16405), .Z(n16359) );
  NAND U24754 ( .A(n16406), .B(n16407), .Z(n16405) );
  NAND U24755 ( .A(n16408), .B(n16409), .Z(n16404) );
  AND U24756 ( .A(n16410), .B(n16411), .Z(n16361) );
  NAND U24757 ( .A(n16412), .B(n16413), .Z(n16355) );
  XNOR U24758 ( .A(n16338), .B(n16414), .Z(n16352) );
  XNOR U24759 ( .A(n16342), .B(n16340), .Z(n16414) );
  XOR U24760 ( .A(n16348), .B(n16415), .Z(n16340) );
  XNOR U24761 ( .A(n16345), .B(n16349), .Z(n16415) );
  AND U24762 ( .A(n16416), .B(n16417), .Z(n16349) );
  NAND U24763 ( .A(n16418), .B(n16419), .Z(n16417) );
  NAND U24764 ( .A(n16420), .B(n16421), .Z(n16416) );
  AND U24765 ( .A(n16422), .B(n16423), .Z(n16345) );
  NAND U24766 ( .A(n16424), .B(n16425), .Z(n16423) );
  NAND U24767 ( .A(n16426), .B(n16427), .Z(n16422) );
  NANDN U24768 ( .A(n16428), .B(n16429), .Z(n16348) );
  ANDN U24769 ( .B(n16430), .A(n16431), .Z(n16342) );
  XNOR U24770 ( .A(n16333), .B(n16432), .Z(n16338) );
  XNOR U24771 ( .A(n16331), .B(n16335), .Z(n16432) );
  AND U24772 ( .A(n16433), .B(n16434), .Z(n16335) );
  NAND U24773 ( .A(n16435), .B(n16436), .Z(n16434) );
  NAND U24774 ( .A(n16437), .B(n16438), .Z(n16433) );
  AND U24775 ( .A(n16439), .B(n16440), .Z(n16331) );
  NAND U24776 ( .A(n16441), .B(n16442), .Z(n16440) );
  NAND U24777 ( .A(n16443), .B(n16444), .Z(n16439) );
  AND U24778 ( .A(n16445), .B(n16446), .Z(n16333) );
  XOR U24779 ( .A(n16413), .B(n16412), .Z(N63933) );
  XNOR U24780 ( .A(n16430), .B(n16431), .Z(n16412) );
  XNOR U24781 ( .A(n16445), .B(n16446), .Z(n16431) );
  XOR U24782 ( .A(n16442), .B(n16441), .Z(n16446) );
  XOR U24783 ( .A(y[6180]), .B(x[6180]), .Z(n16441) );
  XOR U24784 ( .A(n16444), .B(n16443), .Z(n16442) );
  XOR U24785 ( .A(y[6182]), .B(x[6182]), .Z(n16443) );
  XOR U24786 ( .A(y[6181]), .B(x[6181]), .Z(n16444) );
  XOR U24787 ( .A(n16436), .B(n16435), .Z(n16445) );
  XOR U24788 ( .A(n16438), .B(n16437), .Z(n16435) );
  XOR U24789 ( .A(y[6179]), .B(x[6179]), .Z(n16437) );
  XOR U24790 ( .A(y[6178]), .B(x[6178]), .Z(n16438) );
  XOR U24791 ( .A(y[6177]), .B(x[6177]), .Z(n16436) );
  XNOR U24792 ( .A(n16429), .B(n16428), .Z(n16430) );
  XNOR U24793 ( .A(n16425), .B(n16424), .Z(n16428) );
  XOR U24794 ( .A(n16427), .B(n16426), .Z(n16424) );
  XOR U24795 ( .A(y[6176]), .B(x[6176]), .Z(n16426) );
  XOR U24796 ( .A(y[6175]), .B(x[6175]), .Z(n16427) );
  XOR U24797 ( .A(y[6174]), .B(x[6174]), .Z(n16425) );
  XOR U24798 ( .A(n16419), .B(n16418), .Z(n16429) );
  XOR U24799 ( .A(n16421), .B(n16420), .Z(n16418) );
  XOR U24800 ( .A(y[6173]), .B(x[6173]), .Z(n16420) );
  XOR U24801 ( .A(y[6172]), .B(x[6172]), .Z(n16421) );
  XOR U24802 ( .A(y[6171]), .B(x[6171]), .Z(n16419) );
  XNOR U24803 ( .A(n16395), .B(n16396), .Z(n16413) );
  XNOR U24804 ( .A(n16410), .B(n16411), .Z(n16396) );
  XOR U24805 ( .A(n16407), .B(n16406), .Z(n16411) );
  XOR U24806 ( .A(y[6168]), .B(x[6168]), .Z(n16406) );
  XOR U24807 ( .A(n16409), .B(n16408), .Z(n16407) );
  XOR U24808 ( .A(y[6170]), .B(x[6170]), .Z(n16408) );
  XOR U24809 ( .A(y[6169]), .B(x[6169]), .Z(n16409) );
  XOR U24810 ( .A(n16401), .B(n16400), .Z(n16410) );
  XOR U24811 ( .A(n16403), .B(n16402), .Z(n16400) );
  XOR U24812 ( .A(y[6167]), .B(x[6167]), .Z(n16402) );
  XOR U24813 ( .A(y[6166]), .B(x[6166]), .Z(n16403) );
  XOR U24814 ( .A(y[6165]), .B(x[6165]), .Z(n16401) );
  XNOR U24815 ( .A(n16394), .B(n16393), .Z(n16395) );
  XNOR U24816 ( .A(n16390), .B(n16389), .Z(n16393) );
  XOR U24817 ( .A(n16392), .B(n16391), .Z(n16389) );
  XOR U24818 ( .A(y[6164]), .B(x[6164]), .Z(n16391) );
  XOR U24819 ( .A(y[6163]), .B(x[6163]), .Z(n16392) );
  XOR U24820 ( .A(y[6162]), .B(x[6162]), .Z(n16390) );
  XOR U24821 ( .A(n16384), .B(n16383), .Z(n16394) );
  XOR U24822 ( .A(n16386), .B(n16385), .Z(n16383) );
  XOR U24823 ( .A(y[6161]), .B(x[6161]), .Z(n16385) );
  XOR U24824 ( .A(y[6160]), .B(x[6160]), .Z(n16386) );
  XOR U24825 ( .A(y[6159]), .B(x[6159]), .Z(n16384) );
  NAND U24826 ( .A(n16447), .B(n16448), .Z(N63924) );
  NAND U24827 ( .A(n16449), .B(n16450), .Z(n16448) );
  NANDN U24828 ( .A(n16451), .B(n16452), .Z(n16450) );
  NANDN U24829 ( .A(n16452), .B(n16451), .Z(n16447) );
  XOR U24830 ( .A(n16451), .B(n16453), .Z(N63923) );
  XNOR U24831 ( .A(n16449), .B(n16452), .Z(n16453) );
  NAND U24832 ( .A(n16454), .B(n16455), .Z(n16452) );
  NAND U24833 ( .A(n16456), .B(n16457), .Z(n16455) );
  NANDN U24834 ( .A(n16458), .B(n16459), .Z(n16457) );
  NANDN U24835 ( .A(n16459), .B(n16458), .Z(n16454) );
  AND U24836 ( .A(n16460), .B(n16461), .Z(n16449) );
  NAND U24837 ( .A(n16462), .B(n16463), .Z(n16461) );
  NANDN U24838 ( .A(n16464), .B(n16465), .Z(n16463) );
  NANDN U24839 ( .A(n16465), .B(n16464), .Z(n16460) );
  IV U24840 ( .A(n16466), .Z(n16465) );
  AND U24841 ( .A(n16467), .B(n16468), .Z(n16451) );
  NAND U24842 ( .A(n16469), .B(n16470), .Z(n16468) );
  NANDN U24843 ( .A(n16471), .B(n16472), .Z(n16470) );
  NANDN U24844 ( .A(n16472), .B(n16471), .Z(n16467) );
  XOR U24845 ( .A(n16464), .B(n16473), .Z(N63922) );
  XNOR U24846 ( .A(n16462), .B(n16466), .Z(n16473) );
  XOR U24847 ( .A(n16459), .B(n16474), .Z(n16466) );
  XNOR U24848 ( .A(n16456), .B(n16458), .Z(n16474) );
  AND U24849 ( .A(n16475), .B(n16476), .Z(n16458) );
  NANDN U24850 ( .A(n16477), .B(n16478), .Z(n16476) );
  OR U24851 ( .A(n16479), .B(n16480), .Z(n16478) );
  IV U24852 ( .A(n16481), .Z(n16480) );
  NANDN U24853 ( .A(n16481), .B(n16479), .Z(n16475) );
  AND U24854 ( .A(n16482), .B(n16483), .Z(n16456) );
  NAND U24855 ( .A(n16484), .B(n16485), .Z(n16483) );
  NANDN U24856 ( .A(n16486), .B(n16487), .Z(n16485) );
  NANDN U24857 ( .A(n16487), .B(n16486), .Z(n16482) );
  IV U24858 ( .A(n16488), .Z(n16487) );
  NAND U24859 ( .A(n16489), .B(n16490), .Z(n16459) );
  NANDN U24860 ( .A(n16491), .B(n16492), .Z(n16490) );
  NANDN U24861 ( .A(n16493), .B(n16494), .Z(n16492) );
  NANDN U24862 ( .A(n16494), .B(n16493), .Z(n16489) );
  IV U24863 ( .A(n16495), .Z(n16493) );
  AND U24864 ( .A(n16496), .B(n16497), .Z(n16462) );
  NAND U24865 ( .A(n16498), .B(n16499), .Z(n16497) );
  NANDN U24866 ( .A(n16500), .B(n16501), .Z(n16499) );
  NANDN U24867 ( .A(n16501), .B(n16500), .Z(n16496) );
  XOR U24868 ( .A(n16472), .B(n16502), .Z(n16464) );
  XNOR U24869 ( .A(n16469), .B(n16471), .Z(n16502) );
  AND U24870 ( .A(n16503), .B(n16504), .Z(n16471) );
  NANDN U24871 ( .A(n16505), .B(n16506), .Z(n16504) );
  OR U24872 ( .A(n16507), .B(n16508), .Z(n16506) );
  IV U24873 ( .A(n16509), .Z(n16508) );
  NANDN U24874 ( .A(n16509), .B(n16507), .Z(n16503) );
  AND U24875 ( .A(n16510), .B(n16511), .Z(n16469) );
  NAND U24876 ( .A(n16512), .B(n16513), .Z(n16511) );
  NANDN U24877 ( .A(n16514), .B(n16515), .Z(n16513) );
  NANDN U24878 ( .A(n16515), .B(n16514), .Z(n16510) );
  IV U24879 ( .A(n16516), .Z(n16515) );
  NAND U24880 ( .A(n16517), .B(n16518), .Z(n16472) );
  NANDN U24881 ( .A(n16519), .B(n16520), .Z(n16518) );
  NANDN U24882 ( .A(n16521), .B(n16522), .Z(n16520) );
  NANDN U24883 ( .A(n16522), .B(n16521), .Z(n16517) );
  IV U24884 ( .A(n16523), .Z(n16521) );
  XOR U24885 ( .A(n16498), .B(n16524), .Z(N63921) );
  XNOR U24886 ( .A(n16501), .B(n16500), .Z(n16524) );
  XNOR U24887 ( .A(n16512), .B(n16525), .Z(n16500) );
  XNOR U24888 ( .A(n16516), .B(n16514), .Z(n16525) );
  XOR U24889 ( .A(n16522), .B(n16526), .Z(n16514) );
  XNOR U24890 ( .A(n16519), .B(n16523), .Z(n16526) );
  AND U24891 ( .A(n16527), .B(n16528), .Z(n16523) );
  NAND U24892 ( .A(n16529), .B(n16530), .Z(n16528) );
  NAND U24893 ( .A(n16531), .B(n16532), .Z(n16527) );
  AND U24894 ( .A(n16533), .B(n16534), .Z(n16519) );
  NAND U24895 ( .A(n16535), .B(n16536), .Z(n16534) );
  NAND U24896 ( .A(n16537), .B(n16538), .Z(n16533) );
  NANDN U24897 ( .A(n16539), .B(n16540), .Z(n16522) );
  ANDN U24898 ( .B(n16541), .A(n16542), .Z(n16516) );
  XNOR U24899 ( .A(n16507), .B(n16543), .Z(n16512) );
  XNOR U24900 ( .A(n16505), .B(n16509), .Z(n16543) );
  AND U24901 ( .A(n16544), .B(n16545), .Z(n16509) );
  NAND U24902 ( .A(n16546), .B(n16547), .Z(n16545) );
  NAND U24903 ( .A(n16548), .B(n16549), .Z(n16544) );
  AND U24904 ( .A(n16550), .B(n16551), .Z(n16505) );
  NAND U24905 ( .A(n16552), .B(n16553), .Z(n16551) );
  NAND U24906 ( .A(n16554), .B(n16555), .Z(n16550) );
  AND U24907 ( .A(n16556), .B(n16557), .Z(n16507) );
  NAND U24908 ( .A(n16558), .B(n16559), .Z(n16501) );
  XNOR U24909 ( .A(n16484), .B(n16560), .Z(n16498) );
  XNOR U24910 ( .A(n16488), .B(n16486), .Z(n16560) );
  XOR U24911 ( .A(n16494), .B(n16561), .Z(n16486) );
  XNOR U24912 ( .A(n16491), .B(n16495), .Z(n16561) );
  AND U24913 ( .A(n16562), .B(n16563), .Z(n16495) );
  NAND U24914 ( .A(n16564), .B(n16565), .Z(n16563) );
  NAND U24915 ( .A(n16566), .B(n16567), .Z(n16562) );
  AND U24916 ( .A(n16568), .B(n16569), .Z(n16491) );
  NAND U24917 ( .A(n16570), .B(n16571), .Z(n16569) );
  NAND U24918 ( .A(n16572), .B(n16573), .Z(n16568) );
  NANDN U24919 ( .A(n16574), .B(n16575), .Z(n16494) );
  ANDN U24920 ( .B(n16576), .A(n16577), .Z(n16488) );
  XNOR U24921 ( .A(n16479), .B(n16578), .Z(n16484) );
  XNOR U24922 ( .A(n16477), .B(n16481), .Z(n16578) );
  AND U24923 ( .A(n16579), .B(n16580), .Z(n16481) );
  NAND U24924 ( .A(n16581), .B(n16582), .Z(n16580) );
  NAND U24925 ( .A(n16583), .B(n16584), .Z(n16579) );
  AND U24926 ( .A(n16585), .B(n16586), .Z(n16477) );
  NAND U24927 ( .A(n16587), .B(n16588), .Z(n16586) );
  NAND U24928 ( .A(n16589), .B(n16590), .Z(n16585) );
  AND U24929 ( .A(n16591), .B(n16592), .Z(n16479) );
  XOR U24930 ( .A(n16559), .B(n16558), .Z(N63920) );
  XNOR U24931 ( .A(n16576), .B(n16577), .Z(n16558) );
  XNOR U24932 ( .A(n16591), .B(n16592), .Z(n16577) );
  XOR U24933 ( .A(n16588), .B(n16587), .Z(n16592) );
  XOR U24934 ( .A(y[6156]), .B(x[6156]), .Z(n16587) );
  XOR U24935 ( .A(n16590), .B(n16589), .Z(n16588) );
  XOR U24936 ( .A(y[6158]), .B(x[6158]), .Z(n16589) );
  XOR U24937 ( .A(y[6157]), .B(x[6157]), .Z(n16590) );
  XOR U24938 ( .A(n16582), .B(n16581), .Z(n16591) );
  XOR U24939 ( .A(n16584), .B(n16583), .Z(n16581) );
  XOR U24940 ( .A(y[6155]), .B(x[6155]), .Z(n16583) );
  XOR U24941 ( .A(y[6154]), .B(x[6154]), .Z(n16584) );
  XOR U24942 ( .A(y[6153]), .B(x[6153]), .Z(n16582) );
  XNOR U24943 ( .A(n16575), .B(n16574), .Z(n16576) );
  XNOR U24944 ( .A(n16571), .B(n16570), .Z(n16574) );
  XOR U24945 ( .A(n16573), .B(n16572), .Z(n16570) );
  XOR U24946 ( .A(y[6152]), .B(x[6152]), .Z(n16572) );
  XOR U24947 ( .A(y[6151]), .B(x[6151]), .Z(n16573) );
  XOR U24948 ( .A(y[6150]), .B(x[6150]), .Z(n16571) );
  XOR U24949 ( .A(n16565), .B(n16564), .Z(n16575) );
  XOR U24950 ( .A(n16567), .B(n16566), .Z(n16564) );
  XOR U24951 ( .A(y[6149]), .B(x[6149]), .Z(n16566) );
  XOR U24952 ( .A(y[6148]), .B(x[6148]), .Z(n16567) );
  XOR U24953 ( .A(y[6147]), .B(x[6147]), .Z(n16565) );
  XNOR U24954 ( .A(n16541), .B(n16542), .Z(n16559) );
  XNOR U24955 ( .A(n16556), .B(n16557), .Z(n16542) );
  XOR U24956 ( .A(n16553), .B(n16552), .Z(n16557) );
  XOR U24957 ( .A(y[6144]), .B(x[6144]), .Z(n16552) );
  XOR U24958 ( .A(n16555), .B(n16554), .Z(n16553) );
  XOR U24959 ( .A(y[6146]), .B(x[6146]), .Z(n16554) );
  XOR U24960 ( .A(y[6145]), .B(x[6145]), .Z(n16555) );
  XOR U24961 ( .A(n16547), .B(n16546), .Z(n16556) );
  XOR U24962 ( .A(n16549), .B(n16548), .Z(n16546) );
  XOR U24963 ( .A(y[6143]), .B(x[6143]), .Z(n16548) );
  XOR U24964 ( .A(y[6142]), .B(x[6142]), .Z(n16549) );
  XOR U24965 ( .A(y[6141]), .B(x[6141]), .Z(n16547) );
  XNOR U24966 ( .A(n16540), .B(n16539), .Z(n16541) );
  XNOR U24967 ( .A(n16536), .B(n16535), .Z(n16539) );
  XOR U24968 ( .A(n16538), .B(n16537), .Z(n16535) );
  XOR U24969 ( .A(y[6140]), .B(x[6140]), .Z(n16537) );
  XOR U24970 ( .A(y[6139]), .B(x[6139]), .Z(n16538) );
  XOR U24971 ( .A(y[6138]), .B(x[6138]), .Z(n16536) );
  XOR U24972 ( .A(n16530), .B(n16529), .Z(n16540) );
  XOR U24973 ( .A(n16532), .B(n16531), .Z(n16529) );
  XOR U24974 ( .A(y[6137]), .B(x[6137]), .Z(n16531) );
  XOR U24975 ( .A(y[6136]), .B(x[6136]), .Z(n16532) );
  XOR U24976 ( .A(y[6135]), .B(x[6135]), .Z(n16530) );
  NAND U24977 ( .A(n16593), .B(n16594), .Z(N63911) );
  NAND U24978 ( .A(n16595), .B(n16596), .Z(n16594) );
  NANDN U24979 ( .A(n16597), .B(n16598), .Z(n16596) );
  NANDN U24980 ( .A(n16598), .B(n16597), .Z(n16593) );
  XOR U24981 ( .A(n16597), .B(n16599), .Z(N63910) );
  XNOR U24982 ( .A(n16595), .B(n16598), .Z(n16599) );
  NAND U24983 ( .A(n16600), .B(n16601), .Z(n16598) );
  NAND U24984 ( .A(n16602), .B(n16603), .Z(n16601) );
  NANDN U24985 ( .A(n16604), .B(n16605), .Z(n16603) );
  NANDN U24986 ( .A(n16605), .B(n16604), .Z(n16600) );
  AND U24987 ( .A(n16606), .B(n16607), .Z(n16595) );
  NAND U24988 ( .A(n16608), .B(n16609), .Z(n16607) );
  NANDN U24989 ( .A(n16610), .B(n16611), .Z(n16609) );
  NANDN U24990 ( .A(n16611), .B(n16610), .Z(n16606) );
  IV U24991 ( .A(n16612), .Z(n16611) );
  AND U24992 ( .A(n16613), .B(n16614), .Z(n16597) );
  NAND U24993 ( .A(n16615), .B(n16616), .Z(n16614) );
  NANDN U24994 ( .A(n16617), .B(n16618), .Z(n16616) );
  NANDN U24995 ( .A(n16618), .B(n16617), .Z(n16613) );
  XOR U24996 ( .A(n16610), .B(n16619), .Z(N63909) );
  XNOR U24997 ( .A(n16608), .B(n16612), .Z(n16619) );
  XOR U24998 ( .A(n16605), .B(n16620), .Z(n16612) );
  XNOR U24999 ( .A(n16602), .B(n16604), .Z(n16620) );
  AND U25000 ( .A(n16621), .B(n16622), .Z(n16604) );
  NANDN U25001 ( .A(n16623), .B(n16624), .Z(n16622) );
  OR U25002 ( .A(n16625), .B(n16626), .Z(n16624) );
  IV U25003 ( .A(n16627), .Z(n16626) );
  NANDN U25004 ( .A(n16627), .B(n16625), .Z(n16621) );
  AND U25005 ( .A(n16628), .B(n16629), .Z(n16602) );
  NAND U25006 ( .A(n16630), .B(n16631), .Z(n16629) );
  NANDN U25007 ( .A(n16632), .B(n16633), .Z(n16631) );
  NANDN U25008 ( .A(n16633), .B(n16632), .Z(n16628) );
  IV U25009 ( .A(n16634), .Z(n16633) );
  NAND U25010 ( .A(n16635), .B(n16636), .Z(n16605) );
  NANDN U25011 ( .A(n16637), .B(n16638), .Z(n16636) );
  NANDN U25012 ( .A(n16639), .B(n16640), .Z(n16638) );
  NANDN U25013 ( .A(n16640), .B(n16639), .Z(n16635) );
  IV U25014 ( .A(n16641), .Z(n16639) );
  AND U25015 ( .A(n16642), .B(n16643), .Z(n16608) );
  NAND U25016 ( .A(n16644), .B(n16645), .Z(n16643) );
  NANDN U25017 ( .A(n16646), .B(n16647), .Z(n16645) );
  NANDN U25018 ( .A(n16647), .B(n16646), .Z(n16642) );
  XOR U25019 ( .A(n16618), .B(n16648), .Z(n16610) );
  XNOR U25020 ( .A(n16615), .B(n16617), .Z(n16648) );
  AND U25021 ( .A(n16649), .B(n16650), .Z(n16617) );
  NANDN U25022 ( .A(n16651), .B(n16652), .Z(n16650) );
  OR U25023 ( .A(n16653), .B(n16654), .Z(n16652) );
  IV U25024 ( .A(n16655), .Z(n16654) );
  NANDN U25025 ( .A(n16655), .B(n16653), .Z(n16649) );
  AND U25026 ( .A(n16656), .B(n16657), .Z(n16615) );
  NAND U25027 ( .A(n16658), .B(n16659), .Z(n16657) );
  NANDN U25028 ( .A(n16660), .B(n16661), .Z(n16659) );
  NANDN U25029 ( .A(n16661), .B(n16660), .Z(n16656) );
  IV U25030 ( .A(n16662), .Z(n16661) );
  NAND U25031 ( .A(n16663), .B(n16664), .Z(n16618) );
  NANDN U25032 ( .A(n16665), .B(n16666), .Z(n16664) );
  NANDN U25033 ( .A(n16667), .B(n16668), .Z(n16666) );
  NANDN U25034 ( .A(n16668), .B(n16667), .Z(n16663) );
  IV U25035 ( .A(n16669), .Z(n16667) );
  XOR U25036 ( .A(n16644), .B(n16670), .Z(N63908) );
  XNOR U25037 ( .A(n16647), .B(n16646), .Z(n16670) );
  XNOR U25038 ( .A(n16658), .B(n16671), .Z(n16646) );
  XNOR U25039 ( .A(n16662), .B(n16660), .Z(n16671) );
  XOR U25040 ( .A(n16668), .B(n16672), .Z(n16660) );
  XNOR U25041 ( .A(n16665), .B(n16669), .Z(n16672) );
  AND U25042 ( .A(n16673), .B(n16674), .Z(n16669) );
  NAND U25043 ( .A(n16675), .B(n16676), .Z(n16674) );
  NAND U25044 ( .A(n16677), .B(n16678), .Z(n16673) );
  AND U25045 ( .A(n16679), .B(n16680), .Z(n16665) );
  NAND U25046 ( .A(n16681), .B(n16682), .Z(n16680) );
  NAND U25047 ( .A(n16683), .B(n16684), .Z(n16679) );
  NANDN U25048 ( .A(n16685), .B(n16686), .Z(n16668) );
  ANDN U25049 ( .B(n16687), .A(n16688), .Z(n16662) );
  XNOR U25050 ( .A(n16653), .B(n16689), .Z(n16658) );
  XNOR U25051 ( .A(n16651), .B(n16655), .Z(n16689) );
  AND U25052 ( .A(n16690), .B(n16691), .Z(n16655) );
  NAND U25053 ( .A(n16692), .B(n16693), .Z(n16691) );
  NAND U25054 ( .A(n16694), .B(n16695), .Z(n16690) );
  AND U25055 ( .A(n16696), .B(n16697), .Z(n16651) );
  NAND U25056 ( .A(n16698), .B(n16699), .Z(n16697) );
  NAND U25057 ( .A(n16700), .B(n16701), .Z(n16696) );
  AND U25058 ( .A(n16702), .B(n16703), .Z(n16653) );
  NAND U25059 ( .A(n16704), .B(n16705), .Z(n16647) );
  XNOR U25060 ( .A(n16630), .B(n16706), .Z(n16644) );
  XNOR U25061 ( .A(n16634), .B(n16632), .Z(n16706) );
  XOR U25062 ( .A(n16640), .B(n16707), .Z(n16632) );
  XNOR U25063 ( .A(n16637), .B(n16641), .Z(n16707) );
  AND U25064 ( .A(n16708), .B(n16709), .Z(n16641) );
  NAND U25065 ( .A(n16710), .B(n16711), .Z(n16709) );
  NAND U25066 ( .A(n16712), .B(n16713), .Z(n16708) );
  AND U25067 ( .A(n16714), .B(n16715), .Z(n16637) );
  NAND U25068 ( .A(n16716), .B(n16717), .Z(n16715) );
  NAND U25069 ( .A(n16718), .B(n16719), .Z(n16714) );
  NANDN U25070 ( .A(n16720), .B(n16721), .Z(n16640) );
  ANDN U25071 ( .B(n16722), .A(n16723), .Z(n16634) );
  XNOR U25072 ( .A(n16625), .B(n16724), .Z(n16630) );
  XNOR U25073 ( .A(n16623), .B(n16627), .Z(n16724) );
  AND U25074 ( .A(n16725), .B(n16726), .Z(n16627) );
  NAND U25075 ( .A(n16727), .B(n16728), .Z(n16726) );
  NAND U25076 ( .A(n16729), .B(n16730), .Z(n16725) );
  AND U25077 ( .A(n16731), .B(n16732), .Z(n16623) );
  NAND U25078 ( .A(n16733), .B(n16734), .Z(n16732) );
  NAND U25079 ( .A(n16735), .B(n16736), .Z(n16731) );
  AND U25080 ( .A(n16737), .B(n16738), .Z(n16625) );
  XOR U25081 ( .A(n16705), .B(n16704), .Z(N63907) );
  XNOR U25082 ( .A(n16722), .B(n16723), .Z(n16704) );
  XNOR U25083 ( .A(n16737), .B(n16738), .Z(n16723) );
  XOR U25084 ( .A(n16734), .B(n16733), .Z(n16738) );
  XOR U25085 ( .A(y[6132]), .B(x[6132]), .Z(n16733) );
  XOR U25086 ( .A(n16736), .B(n16735), .Z(n16734) );
  XOR U25087 ( .A(y[6134]), .B(x[6134]), .Z(n16735) );
  XOR U25088 ( .A(y[6133]), .B(x[6133]), .Z(n16736) );
  XOR U25089 ( .A(n16728), .B(n16727), .Z(n16737) );
  XOR U25090 ( .A(n16730), .B(n16729), .Z(n16727) );
  XOR U25091 ( .A(y[6131]), .B(x[6131]), .Z(n16729) );
  XOR U25092 ( .A(y[6130]), .B(x[6130]), .Z(n16730) );
  XOR U25093 ( .A(y[6129]), .B(x[6129]), .Z(n16728) );
  XNOR U25094 ( .A(n16721), .B(n16720), .Z(n16722) );
  XNOR U25095 ( .A(n16717), .B(n16716), .Z(n16720) );
  XOR U25096 ( .A(n16719), .B(n16718), .Z(n16716) );
  XOR U25097 ( .A(y[6128]), .B(x[6128]), .Z(n16718) );
  XOR U25098 ( .A(y[6127]), .B(x[6127]), .Z(n16719) );
  XOR U25099 ( .A(y[6126]), .B(x[6126]), .Z(n16717) );
  XOR U25100 ( .A(n16711), .B(n16710), .Z(n16721) );
  XOR U25101 ( .A(n16713), .B(n16712), .Z(n16710) );
  XOR U25102 ( .A(y[6125]), .B(x[6125]), .Z(n16712) );
  XOR U25103 ( .A(y[6124]), .B(x[6124]), .Z(n16713) );
  XOR U25104 ( .A(y[6123]), .B(x[6123]), .Z(n16711) );
  XNOR U25105 ( .A(n16687), .B(n16688), .Z(n16705) );
  XNOR U25106 ( .A(n16702), .B(n16703), .Z(n16688) );
  XOR U25107 ( .A(n16699), .B(n16698), .Z(n16703) );
  XOR U25108 ( .A(y[6120]), .B(x[6120]), .Z(n16698) );
  XOR U25109 ( .A(n16701), .B(n16700), .Z(n16699) );
  XOR U25110 ( .A(y[6122]), .B(x[6122]), .Z(n16700) );
  XOR U25111 ( .A(y[6121]), .B(x[6121]), .Z(n16701) );
  XOR U25112 ( .A(n16693), .B(n16692), .Z(n16702) );
  XOR U25113 ( .A(n16695), .B(n16694), .Z(n16692) );
  XOR U25114 ( .A(y[6119]), .B(x[6119]), .Z(n16694) );
  XOR U25115 ( .A(y[6118]), .B(x[6118]), .Z(n16695) );
  XOR U25116 ( .A(y[6117]), .B(x[6117]), .Z(n16693) );
  XNOR U25117 ( .A(n16686), .B(n16685), .Z(n16687) );
  XNOR U25118 ( .A(n16682), .B(n16681), .Z(n16685) );
  XOR U25119 ( .A(n16684), .B(n16683), .Z(n16681) );
  XOR U25120 ( .A(y[6116]), .B(x[6116]), .Z(n16683) );
  XOR U25121 ( .A(y[6115]), .B(x[6115]), .Z(n16684) );
  XOR U25122 ( .A(y[6114]), .B(x[6114]), .Z(n16682) );
  XOR U25123 ( .A(n16676), .B(n16675), .Z(n16686) );
  XOR U25124 ( .A(n16678), .B(n16677), .Z(n16675) );
  XOR U25125 ( .A(y[6113]), .B(x[6113]), .Z(n16677) );
  XOR U25126 ( .A(y[6112]), .B(x[6112]), .Z(n16678) );
  XOR U25127 ( .A(y[6111]), .B(x[6111]), .Z(n16676) );
  NAND U25128 ( .A(n16739), .B(n16740), .Z(N63898) );
  NAND U25129 ( .A(n16741), .B(n16742), .Z(n16740) );
  NANDN U25130 ( .A(n16743), .B(n16744), .Z(n16742) );
  NANDN U25131 ( .A(n16744), .B(n16743), .Z(n16739) );
  XOR U25132 ( .A(n16743), .B(n16745), .Z(N63897) );
  XNOR U25133 ( .A(n16741), .B(n16744), .Z(n16745) );
  NAND U25134 ( .A(n16746), .B(n16747), .Z(n16744) );
  NAND U25135 ( .A(n16748), .B(n16749), .Z(n16747) );
  NANDN U25136 ( .A(n16750), .B(n16751), .Z(n16749) );
  NANDN U25137 ( .A(n16751), .B(n16750), .Z(n16746) );
  AND U25138 ( .A(n16752), .B(n16753), .Z(n16741) );
  NAND U25139 ( .A(n16754), .B(n16755), .Z(n16753) );
  NANDN U25140 ( .A(n16756), .B(n16757), .Z(n16755) );
  NANDN U25141 ( .A(n16757), .B(n16756), .Z(n16752) );
  IV U25142 ( .A(n16758), .Z(n16757) );
  AND U25143 ( .A(n16759), .B(n16760), .Z(n16743) );
  NAND U25144 ( .A(n16761), .B(n16762), .Z(n16760) );
  NANDN U25145 ( .A(n16763), .B(n16764), .Z(n16762) );
  NANDN U25146 ( .A(n16764), .B(n16763), .Z(n16759) );
  XOR U25147 ( .A(n16756), .B(n16765), .Z(N63896) );
  XNOR U25148 ( .A(n16754), .B(n16758), .Z(n16765) );
  XOR U25149 ( .A(n16751), .B(n16766), .Z(n16758) );
  XNOR U25150 ( .A(n16748), .B(n16750), .Z(n16766) );
  AND U25151 ( .A(n16767), .B(n16768), .Z(n16750) );
  NANDN U25152 ( .A(n16769), .B(n16770), .Z(n16768) );
  OR U25153 ( .A(n16771), .B(n16772), .Z(n16770) );
  IV U25154 ( .A(n16773), .Z(n16772) );
  NANDN U25155 ( .A(n16773), .B(n16771), .Z(n16767) );
  AND U25156 ( .A(n16774), .B(n16775), .Z(n16748) );
  NAND U25157 ( .A(n16776), .B(n16777), .Z(n16775) );
  NANDN U25158 ( .A(n16778), .B(n16779), .Z(n16777) );
  NANDN U25159 ( .A(n16779), .B(n16778), .Z(n16774) );
  IV U25160 ( .A(n16780), .Z(n16779) );
  NAND U25161 ( .A(n16781), .B(n16782), .Z(n16751) );
  NANDN U25162 ( .A(n16783), .B(n16784), .Z(n16782) );
  NANDN U25163 ( .A(n16785), .B(n16786), .Z(n16784) );
  NANDN U25164 ( .A(n16786), .B(n16785), .Z(n16781) );
  IV U25165 ( .A(n16787), .Z(n16785) );
  AND U25166 ( .A(n16788), .B(n16789), .Z(n16754) );
  NAND U25167 ( .A(n16790), .B(n16791), .Z(n16789) );
  NANDN U25168 ( .A(n16792), .B(n16793), .Z(n16791) );
  NANDN U25169 ( .A(n16793), .B(n16792), .Z(n16788) );
  XOR U25170 ( .A(n16764), .B(n16794), .Z(n16756) );
  XNOR U25171 ( .A(n16761), .B(n16763), .Z(n16794) );
  AND U25172 ( .A(n16795), .B(n16796), .Z(n16763) );
  NANDN U25173 ( .A(n16797), .B(n16798), .Z(n16796) );
  OR U25174 ( .A(n16799), .B(n16800), .Z(n16798) );
  IV U25175 ( .A(n16801), .Z(n16800) );
  NANDN U25176 ( .A(n16801), .B(n16799), .Z(n16795) );
  AND U25177 ( .A(n16802), .B(n16803), .Z(n16761) );
  NAND U25178 ( .A(n16804), .B(n16805), .Z(n16803) );
  NANDN U25179 ( .A(n16806), .B(n16807), .Z(n16805) );
  NANDN U25180 ( .A(n16807), .B(n16806), .Z(n16802) );
  IV U25181 ( .A(n16808), .Z(n16807) );
  NAND U25182 ( .A(n16809), .B(n16810), .Z(n16764) );
  NANDN U25183 ( .A(n16811), .B(n16812), .Z(n16810) );
  NANDN U25184 ( .A(n16813), .B(n16814), .Z(n16812) );
  NANDN U25185 ( .A(n16814), .B(n16813), .Z(n16809) );
  IV U25186 ( .A(n16815), .Z(n16813) );
  XOR U25187 ( .A(n16790), .B(n16816), .Z(N63895) );
  XNOR U25188 ( .A(n16793), .B(n16792), .Z(n16816) );
  XNOR U25189 ( .A(n16804), .B(n16817), .Z(n16792) );
  XNOR U25190 ( .A(n16808), .B(n16806), .Z(n16817) );
  XOR U25191 ( .A(n16814), .B(n16818), .Z(n16806) );
  XNOR U25192 ( .A(n16811), .B(n16815), .Z(n16818) );
  AND U25193 ( .A(n16819), .B(n16820), .Z(n16815) );
  NAND U25194 ( .A(n16821), .B(n16822), .Z(n16820) );
  NAND U25195 ( .A(n16823), .B(n16824), .Z(n16819) );
  AND U25196 ( .A(n16825), .B(n16826), .Z(n16811) );
  NAND U25197 ( .A(n16827), .B(n16828), .Z(n16826) );
  NAND U25198 ( .A(n16829), .B(n16830), .Z(n16825) );
  NANDN U25199 ( .A(n16831), .B(n16832), .Z(n16814) );
  ANDN U25200 ( .B(n16833), .A(n16834), .Z(n16808) );
  XNOR U25201 ( .A(n16799), .B(n16835), .Z(n16804) );
  XNOR U25202 ( .A(n16797), .B(n16801), .Z(n16835) );
  AND U25203 ( .A(n16836), .B(n16837), .Z(n16801) );
  NAND U25204 ( .A(n16838), .B(n16839), .Z(n16837) );
  NAND U25205 ( .A(n16840), .B(n16841), .Z(n16836) );
  AND U25206 ( .A(n16842), .B(n16843), .Z(n16797) );
  NAND U25207 ( .A(n16844), .B(n16845), .Z(n16843) );
  NAND U25208 ( .A(n16846), .B(n16847), .Z(n16842) );
  AND U25209 ( .A(n16848), .B(n16849), .Z(n16799) );
  NAND U25210 ( .A(n16850), .B(n16851), .Z(n16793) );
  XNOR U25211 ( .A(n16776), .B(n16852), .Z(n16790) );
  XNOR U25212 ( .A(n16780), .B(n16778), .Z(n16852) );
  XOR U25213 ( .A(n16786), .B(n16853), .Z(n16778) );
  XNOR U25214 ( .A(n16783), .B(n16787), .Z(n16853) );
  AND U25215 ( .A(n16854), .B(n16855), .Z(n16787) );
  NAND U25216 ( .A(n16856), .B(n16857), .Z(n16855) );
  NAND U25217 ( .A(n16858), .B(n16859), .Z(n16854) );
  AND U25218 ( .A(n16860), .B(n16861), .Z(n16783) );
  NAND U25219 ( .A(n16862), .B(n16863), .Z(n16861) );
  NAND U25220 ( .A(n16864), .B(n16865), .Z(n16860) );
  NANDN U25221 ( .A(n16866), .B(n16867), .Z(n16786) );
  ANDN U25222 ( .B(n16868), .A(n16869), .Z(n16780) );
  XNOR U25223 ( .A(n16771), .B(n16870), .Z(n16776) );
  XNOR U25224 ( .A(n16769), .B(n16773), .Z(n16870) );
  AND U25225 ( .A(n16871), .B(n16872), .Z(n16773) );
  NAND U25226 ( .A(n16873), .B(n16874), .Z(n16872) );
  NAND U25227 ( .A(n16875), .B(n16876), .Z(n16871) );
  AND U25228 ( .A(n16877), .B(n16878), .Z(n16769) );
  NAND U25229 ( .A(n16879), .B(n16880), .Z(n16878) );
  NAND U25230 ( .A(n16881), .B(n16882), .Z(n16877) );
  AND U25231 ( .A(n16883), .B(n16884), .Z(n16771) );
  XOR U25232 ( .A(n16851), .B(n16850), .Z(N63894) );
  XNOR U25233 ( .A(n16868), .B(n16869), .Z(n16850) );
  XNOR U25234 ( .A(n16883), .B(n16884), .Z(n16869) );
  XOR U25235 ( .A(n16880), .B(n16879), .Z(n16884) );
  XOR U25236 ( .A(y[6108]), .B(x[6108]), .Z(n16879) );
  XOR U25237 ( .A(n16882), .B(n16881), .Z(n16880) );
  XOR U25238 ( .A(y[6110]), .B(x[6110]), .Z(n16881) );
  XOR U25239 ( .A(y[6109]), .B(x[6109]), .Z(n16882) );
  XOR U25240 ( .A(n16874), .B(n16873), .Z(n16883) );
  XOR U25241 ( .A(n16876), .B(n16875), .Z(n16873) );
  XOR U25242 ( .A(y[6107]), .B(x[6107]), .Z(n16875) );
  XOR U25243 ( .A(y[6106]), .B(x[6106]), .Z(n16876) );
  XOR U25244 ( .A(y[6105]), .B(x[6105]), .Z(n16874) );
  XNOR U25245 ( .A(n16867), .B(n16866), .Z(n16868) );
  XNOR U25246 ( .A(n16863), .B(n16862), .Z(n16866) );
  XOR U25247 ( .A(n16865), .B(n16864), .Z(n16862) );
  XOR U25248 ( .A(y[6104]), .B(x[6104]), .Z(n16864) );
  XOR U25249 ( .A(y[6103]), .B(x[6103]), .Z(n16865) );
  XOR U25250 ( .A(y[6102]), .B(x[6102]), .Z(n16863) );
  XOR U25251 ( .A(n16857), .B(n16856), .Z(n16867) );
  XOR U25252 ( .A(n16859), .B(n16858), .Z(n16856) );
  XOR U25253 ( .A(y[6101]), .B(x[6101]), .Z(n16858) );
  XOR U25254 ( .A(y[6100]), .B(x[6100]), .Z(n16859) );
  XOR U25255 ( .A(y[6099]), .B(x[6099]), .Z(n16857) );
  XNOR U25256 ( .A(n16833), .B(n16834), .Z(n16851) );
  XNOR U25257 ( .A(n16848), .B(n16849), .Z(n16834) );
  XOR U25258 ( .A(n16845), .B(n16844), .Z(n16849) );
  XOR U25259 ( .A(y[6096]), .B(x[6096]), .Z(n16844) );
  XOR U25260 ( .A(n16847), .B(n16846), .Z(n16845) );
  XOR U25261 ( .A(y[6098]), .B(x[6098]), .Z(n16846) );
  XOR U25262 ( .A(y[6097]), .B(x[6097]), .Z(n16847) );
  XOR U25263 ( .A(n16839), .B(n16838), .Z(n16848) );
  XOR U25264 ( .A(n16841), .B(n16840), .Z(n16838) );
  XOR U25265 ( .A(y[6095]), .B(x[6095]), .Z(n16840) );
  XOR U25266 ( .A(y[6094]), .B(x[6094]), .Z(n16841) );
  XOR U25267 ( .A(y[6093]), .B(x[6093]), .Z(n16839) );
  XNOR U25268 ( .A(n16832), .B(n16831), .Z(n16833) );
  XNOR U25269 ( .A(n16828), .B(n16827), .Z(n16831) );
  XOR U25270 ( .A(n16830), .B(n16829), .Z(n16827) );
  XOR U25271 ( .A(y[6092]), .B(x[6092]), .Z(n16829) );
  XOR U25272 ( .A(y[6091]), .B(x[6091]), .Z(n16830) );
  XOR U25273 ( .A(y[6090]), .B(x[6090]), .Z(n16828) );
  XOR U25274 ( .A(n16822), .B(n16821), .Z(n16832) );
  XOR U25275 ( .A(n16824), .B(n16823), .Z(n16821) );
  XOR U25276 ( .A(y[6089]), .B(x[6089]), .Z(n16823) );
  XOR U25277 ( .A(y[6088]), .B(x[6088]), .Z(n16824) );
  XOR U25278 ( .A(y[6087]), .B(x[6087]), .Z(n16822) );
  NAND U25279 ( .A(n16885), .B(n16886), .Z(N63885) );
  NAND U25280 ( .A(n16887), .B(n16888), .Z(n16886) );
  NANDN U25281 ( .A(n16889), .B(n16890), .Z(n16888) );
  NANDN U25282 ( .A(n16890), .B(n16889), .Z(n16885) );
  XOR U25283 ( .A(n16889), .B(n16891), .Z(N63884) );
  XNOR U25284 ( .A(n16887), .B(n16890), .Z(n16891) );
  NAND U25285 ( .A(n16892), .B(n16893), .Z(n16890) );
  NAND U25286 ( .A(n16894), .B(n16895), .Z(n16893) );
  NANDN U25287 ( .A(n16896), .B(n16897), .Z(n16895) );
  NANDN U25288 ( .A(n16897), .B(n16896), .Z(n16892) );
  AND U25289 ( .A(n16898), .B(n16899), .Z(n16887) );
  NAND U25290 ( .A(n16900), .B(n16901), .Z(n16899) );
  NANDN U25291 ( .A(n16902), .B(n16903), .Z(n16901) );
  NANDN U25292 ( .A(n16903), .B(n16902), .Z(n16898) );
  IV U25293 ( .A(n16904), .Z(n16903) );
  AND U25294 ( .A(n16905), .B(n16906), .Z(n16889) );
  NAND U25295 ( .A(n16907), .B(n16908), .Z(n16906) );
  NANDN U25296 ( .A(n16909), .B(n16910), .Z(n16908) );
  NANDN U25297 ( .A(n16910), .B(n16909), .Z(n16905) );
  XOR U25298 ( .A(n16902), .B(n16911), .Z(N63883) );
  XNOR U25299 ( .A(n16900), .B(n16904), .Z(n16911) );
  XOR U25300 ( .A(n16897), .B(n16912), .Z(n16904) );
  XNOR U25301 ( .A(n16894), .B(n16896), .Z(n16912) );
  AND U25302 ( .A(n16913), .B(n16914), .Z(n16896) );
  NANDN U25303 ( .A(n16915), .B(n16916), .Z(n16914) );
  OR U25304 ( .A(n16917), .B(n16918), .Z(n16916) );
  IV U25305 ( .A(n16919), .Z(n16918) );
  NANDN U25306 ( .A(n16919), .B(n16917), .Z(n16913) );
  AND U25307 ( .A(n16920), .B(n16921), .Z(n16894) );
  NAND U25308 ( .A(n16922), .B(n16923), .Z(n16921) );
  NANDN U25309 ( .A(n16924), .B(n16925), .Z(n16923) );
  NANDN U25310 ( .A(n16925), .B(n16924), .Z(n16920) );
  IV U25311 ( .A(n16926), .Z(n16925) );
  NAND U25312 ( .A(n16927), .B(n16928), .Z(n16897) );
  NANDN U25313 ( .A(n16929), .B(n16930), .Z(n16928) );
  NANDN U25314 ( .A(n16931), .B(n16932), .Z(n16930) );
  NANDN U25315 ( .A(n16932), .B(n16931), .Z(n16927) );
  IV U25316 ( .A(n16933), .Z(n16931) );
  AND U25317 ( .A(n16934), .B(n16935), .Z(n16900) );
  NAND U25318 ( .A(n16936), .B(n16937), .Z(n16935) );
  NANDN U25319 ( .A(n16938), .B(n16939), .Z(n16937) );
  NANDN U25320 ( .A(n16939), .B(n16938), .Z(n16934) );
  XOR U25321 ( .A(n16910), .B(n16940), .Z(n16902) );
  XNOR U25322 ( .A(n16907), .B(n16909), .Z(n16940) );
  AND U25323 ( .A(n16941), .B(n16942), .Z(n16909) );
  NANDN U25324 ( .A(n16943), .B(n16944), .Z(n16942) );
  OR U25325 ( .A(n16945), .B(n16946), .Z(n16944) );
  IV U25326 ( .A(n16947), .Z(n16946) );
  NANDN U25327 ( .A(n16947), .B(n16945), .Z(n16941) );
  AND U25328 ( .A(n16948), .B(n16949), .Z(n16907) );
  NAND U25329 ( .A(n16950), .B(n16951), .Z(n16949) );
  NANDN U25330 ( .A(n16952), .B(n16953), .Z(n16951) );
  NANDN U25331 ( .A(n16953), .B(n16952), .Z(n16948) );
  IV U25332 ( .A(n16954), .Z(n16953) );
  NAND U25333 ( .A(n16955), .B(n16956), .Z(n16910) );
  NANDN U25334 ( .A(n16957), .B(n16958), .Z(n16956) );
  NANDN U25335 ( .A(n16959), .B(n16960), .Z(n16958) );
  NANDN U25336 ( .A(n16960), .B(n16959), .Z(n16955) );
  IV U25337 ( .A(n16961), .Z(n16959) );
  XOR U25338 ( .A(n16936), .B(n16962), .Z(N63882) );
  XNOR U25339 ( .A(n16939), .B(n16938), .Z(n16962) );
  XNOR U25340 ( .A(n16950), .B(n16963), .Z(n16938) );
  XNOR U25341 ( .A(n16954), .B(n16952), .Z(n16963) );
  XOR U25342 ( .A(n16960), .B(n16964), .Z(n16952) );
  XNOR U25343 ( .A(n16957), .B(n16961), .Z(n16964) );
  AND U25344 ( .A(n16965), .B(n16966), .Z(n16961) );
  NAND U25345 ( .A(n16967), .B(n16968), .Z(n16966) );
  NAND U25346 ( .A(n16969), .B(n16970), .Z(n16965) );
  AND U25347 ( .A(n16971), .B(n16972), .Z(n16957) );
  NAND U25348 ( .A(n16973), .B(n16974), .Z(n16972) );
  NAND U25349 ( .A(n16975), .B(n16976), .Z(n16971) );
  NANDN U25350 ( .A(n16977), .B(n16978), .Z(n16960) );
  ANDN U25351 ( .B(n16979), .A(n16980), .Z(n16954) );
  XNOR U25352 ( .A(n16945), .B(n16981), .Z(n16950) );
  XNOR U25353 ( .A(n16943), .B(n16947), .Z(n16981) );
  AND U25354 ( .A(n16982), .B(n16983), .Z(n16947) );
  NAND U25355 ( .A(n16984), .B(n16985), .Z(n16983) );
  NAND U25356 ( .A(n16986), .B(n16987), .Z(n16982) );
  AND U25357 ( .A(n16988), .B(n16989), .Z(n16943) );
  NAND U25358 ( .A(n16990), .B(n16991), .Z(n16989) );
  NAND U25359 ( .A(n16992), .B(n16993), .Z(n16988) );
  AND U25360 ( .A(n16994), .B(n16995), .Z(n16945) );
  NAND U25361 ( .A(n16996), .B(n16997), .Z(n16939) );
  XNOR U25362 ( .A(n16922), .B(n16998), .Z(n16936) );
  XNOR U25363 ( .A(n16926), .B(n16924), .Z(n16998) );
  XOR U25364 ( .A(n16932), .B(n16999), .Z(n16924) );
  XNOR U25365 ( .A(n16929), .B(n16933), .Z(n16999) );
  AND U25366 ( .A(n17000), .B(n17001), .Z(n16933) );
  NAND U25367 ( .A(n17002), .B(n17003), .Z(n17001) );
  NAND U25368 ( .A(n17004), .B(n17005), .Z(n17000) );
  AND U25369 ( .A(n17006), .B(n17007), .Z(n16929) );
  NAND U25370 ( .A(n17008), .B(n17009), .Z(n17007) );
  NAND U25371 ( .A(n17010), .B(n17011), .Z(n17006) );
  NANDN U25372 ( .A(n17012), .B(n17013), .Z(n16932) );
  ANDN U25373 ( .B(n17014), .A(n17015), .Z(n16926) );
  XNOR U25374 ( .A(n16917), .B(n17016), .Z(n16922) );
  XNOR U25375 ( .A(n16915), .B(n16919), .Z(n17016) );
  AND U25376 ( .A(n17017), .B(n17018), .Z(n16919) );
  NAND U25377 ( .A(n17019), .B(n17020), .Z(n17018) );
  NAND U25378 ( .A(n17021), .B(n17022), .Z(n17017) );
  AND U25379 ( .A(n17023), .B(n17024), .Z(n16915) );
  NAND U25380 ( .A(n17025), .B(n17026), .Z(n17024) );
  NAND U25381 ( .A(n17027), .B(n17028), .Z(n17023) );
  AND U25382 ( .A(n17029), .B(n17030), .Z(n16917) );
  XOR U25383 ( .A(n16997), .B(n16996), .Z(N63881) );
  XNOR U25384 ( .A(n17014), .B(n17015), .Z(n16996) );
  XNOR U25385 ( .A(n17029), .B(n17030), .Z(n17015) );
  XOR U25386 ( .A(n17026), .B(n17025), .Z(n17030) );
  XOR U25387 ( .A(y[6084]), .B(x[6084]), .Z(n17025) );
  XOR U25388 ( .A(n17028), .B(n17027), .Z(n17026) );
  XOR U25389 ( .A(y[6086]), .B(x[6086]), .Z(n17027) );
  XOR U25390 ( .A(y[6085]), .B(x[6085]), .Z(n17028) );
  XOR U25391 ( .A(n17020), .B(n17019), .Z(n17029) );
  XOR U25392 ( .A(n17022), .B(n17021), .Z(n17019) );
  XOR U25393 ( .A(y[6083]), .B(x[6083]), .Z(n17021) );
  XOR U25394 ( .A(y[6082]), .B(x[6082]), .Z(n17022) );
  XOR U25395 ( .A(y[6081]), .B(x[6081]), .Z(n17020) );
  XNOR U25396 ( .A(n17013), .B(n17012), .Z(n17014) );
  XNOR U25397 ( .A(n17009), .B(n17008), .Z(n17012) );
  XOR U25398 ( .A(n17011), .B(n17010), .Z(n17008) );
  XOR U25399 ( .A(y[6080]), .B(x[6080]), .Z(n17010) );
  XOR U25400 ( .A(y[6079]), .B(x[6079]), .Z(n17011) );
  XOR U25401 ( .A(y[6078]), .B(x[6078]), .Z(n17009) );
  XOR U25402 ( .A(n17003), .B(n17002), .Z(n17013) );
  XOR U25403 ( .A(n17005), .B(n17004), .Z(n17002) );
  XOR U25404 ( .A(y[6077]), .B(x[6077]), .Z(n17004) );
  XOR U25405 ( .A(y[6076]), .B(x[6076]), .Z(n17005) );
  XOR U25406 ( .A(y[6075]), .B(x[6075]), .Z(n17003) );
  XNOR U25407 ( .A(n16979), .B(n16980), .Z(n16997) );
  XNOR U25408 ( .A(n16994), .B(n16995), .Z(n16980) );
  XOR U25409 ( .A(n16991), .B(n16990), .Z(n16995) );
  XOR U25410 ( .A(y[6072]), .B(x[6072]), .Z(n16990) );
  XOR U25411 ( .A(n16993), .B(n16992), .Z(n16991) );
  XOR U25412 ( .A(y[6074]), .B(x[6074]), .Z(n16992) );
  XOR U25413 ( .A(y[6073]), .B(x[6073]), .Z(n16993) );
  XOR U25414 ( .A(n16985), .B(n16984), .Z(n16994) );
  XOR U25415 ( .A(n16987), .B(n16986), .Z(n16984) );
  XOR U25416 ( .A(y[6071]), .B(x[6071]), .Z(n16986) );
  XOR U25417 ( .A(y[6070]), .B(x[6070]), .Z(n16987) );
  XOR U25418 ( .A(y[6069]), .B(x[6069]), .Z(n16985) );
  XNOR U25419 ( .A(n16978), .B(n16977), .Z(n16979) );
  XNOR U25420 ( .A(n16974), .B(n16973), .Z(n16977) );
  XOR U25421 ( .A(n16976), .B(n16975), .Z(n16973) );
  XOR U25422 ( .A(y[6068]), .B(x[6068]), .Z(n16975) );
  XOR U25423 ( .A(y[6067]), .B(x[6067]), .Z(n16976) );
  XOR U25424 ( .A(y[6066]), .B(x[6066]), .Z(n16974) );
  XOR U25425 ( .A(n16968), .B(n16967), .Z(n16978) );
  XOR U25426 ( .A(n16970), .B(n16969), .Z(n16967) );
  XOR U25427 ( .A(y[6065]), .B(x[6065]), .Z(n16969) );
  XOR U25428 ( .A(y[6064]), .B(x[6064]), .Z(n16970) );
  XOR U25429 ( .A(y[6063]), .B(x[6063]), .Z(n16968) );
  NAND U25430 ( .A(n17031), .B(n17032), .Z(N63872) );
  NAND U25431 ( .A(n17033), .B(n17034), .Z(n17032) );
  NANDN U25432 ( .A(n17035), .B(n17036), .Z(n17034) );
  NANDN U25433 ( .A(n17036), .B(n17035), .Z(n17031) );
  XOR U25434 ( .A(n17035), .B(n17037), .Z(N63871) );
  XNOR U25435 ( .A(n17033), .B(n17036), .Z(n17037) );
  NAND U25436 ( .A(n17038), .B(n17039), .Z(n17036) );
  NAND U25437 ( .A(n17040), .B(n17041), .Z(n17039) );
  NANDN U25438 ( .A(n17042), .B(n17043), .Z(n17041) );
  NANDN U25439 ( .A(n17043), .B(n17042), .Z(n17038) );
  AND U25440 ( .A(n17044), .B(n17045), .Z(n17033) );
  NAND U25441 ( .A(n17046), .B(n17047), .Z(n17045) );
  NANDN U25442 ( .A(n17048), .B(n17049), .Z(n17047) );
  NANDN U25443 ( .A(n17049), .B(n17048), .Z(n17044) );
  IV U25444 ( .A(n17050), .Z(n17049) );
  AND U25445 ( .A(n17051), .B(n17052), .Z(n17035) );
  NAND U25446 ( .A(n17053), .B(n17054), .Z(n17052) );
  NANDN U25447 ( .A(n17055), .B(n17056), .Z(n17054) );
  NANDN U25448 ( .A(n17056), .B(n17055), .Z(n17051) );
  XOR U25449 ( .A(n17048), .B(n17057), .Z(N63870) );
  XNOR U25450 ( .A(n17046), .B(n17050), .Z(n17057) );
  XOR U25451 ( .A(n17043), .B(n17058), .Z(n17050) );
  XNOR U25452 ( .A(n17040), .B(n17042), .Z(n17058) );
  AND U25453 ( .A(n17059), .B(n17060), .Z(n17042) );
  NANDN U25454 ( .A(n17061), .B(n17062), .Z(n17060) );
  OR U25455 ( .A(n17063), .B(n17064), .Z(n17062) );
  IV U25456 ( .A(n17065), .Z(n17064) );
  NANDN U25457 ( .A(n17065), .B(n17063), .Z(n17059) );
  AND U25458 ( .A(n17066), .B(n17067), .Z(n17040) );
  NAND U25459 ( .A(n17068), .B(n17069), .Z(n17067) );
  NANDN U25460 ( .A(n17070), .B(n17071), .Z(n17069) );
  NANDN U25461 ( .A(n17071), .B(n17070), .Z(n17066) );
  IV U25462 ( .A(n17072), .Z(n17071) );
  NAND U25463 ( .A(n17073), .B(n17074), .Z(n17043) );
  NANDN U25464 ( .A(n17075), .B(n17076), .Z(n17074) );
  NANDN U25465 ( .A(n17077), .B(n17078), .Z(n17076) );
  NANDN U25466 ( .A(n17078), .B(n17077), .Z(n17073) );
  IV U25467 ( .A(n17079), .Z(n17077) );
  AND U25468 ( .A(n17080), .B(n17081), .Z(n17046) );
  NAND U25469 ( .A(n17082), .B(n17083), .Z(n17081) );
  NANDN U25470 ( .A(n17084), .B(n17085), .Z(n17083) );
  NANDN U25471 ( .A(n17085), .B(n17084), .Z(n17080) );
  XOR U25472 ( .A(n17056), .B(n17086), .Z(n17048) );
  XNOR U25473 ( .A(n17053), .B(n17055), .Z(n17086) );
  AND U25474 ( .A(n17087), .B(n17088), .Z(n17055) );
  NANDN U25475 ( .A(n17089), .B(n17090), .Z(n17088) );
  OR U25476 ( .A(n17091), .B(n17092), .Z(n17090) );
  IV U25477 ( .A(n17093), .Z(n17092) );
  NANDN U25478 ( .A(n17093), .B(n17091), .Z(n17087) );
  AND U25479 ( .A(n17094), .B(n17095), .Z(n17053) );
  NAND U25480 ( .A(n17096), .B(n17097), .Z(n17095) );
  NANDN U25481 ( .A(n17098), .B(n17099), .Z(n17097) );
  NANDN U25482 ( .A(n17099), .B(n17098), .Z(n17094) );
  IV U25483 ( .A(n17100), .Z(n17099) );
  NAND U25484 ( .A(n17101), .B(n17102), .Z(n17056) );
  NANDN U25485 ( .A(n17103), .B(n17104), .Z(n17102) );
  NANDN U25486 ( .A(n17105), .B(n17106), .Z(n17104) );
  NANDN U25487 ( .A(n17106), .B(n17105), .Z(n17101) );
  IV U25488 ( .A(n17107), .Z(n17105) );
  XOR U25489 ( .A(n17082), .B(n17108), .Z(N63869) );
  XNOR U25490 ( .A(n17085), .B(n17084), .Z(n17108) );
  XNOR U25491 ( .A(n17096), .B(n17109), .Z(n17084) );
  XNOR U25492 ( .A(n17100), .B(n17098), .Z(n17109) );
  XOR U25493 ( .A(n17106), .B(n17110), .Z(n17098) );
  XNOR U25494 ( .A(n17103), .B(n17107), .Z(n17110) );
  AND U25495 ( .A(n17111), .B(n17112), .Z(n17107) );
  NAND U25496 ( .A(n17113), .B(n17114), .Z(n17112) );
  NAND U25497 ( .A(n17115), .B(n17116), .Z(n17111) );
  AND U25498 ( .A(n17117), .B(n17118), .Z(n17103) );
  NAND U25499 ( .A(n17119), .B(n17120), .Z(n17118) );
  NAND U25500 ( .A(n17121), .B(n17122), .Z(n17117) );
  NANDN U25501 ( .A(n17123), .B(n17124), .Z(n17106) );
  ANDN U25502 ( .B(n17125), .A(n17126), .Z(n17100) );
  XNOR U25503 ( .A(n17091), .B(n17127), .Z(n17096) );
  XNOR U25504 ( .A(n17089), .B(n17093), .Z(n17127) );
  AND U25505 ( .A(n17128), .B(n17129), .Z(n17093) );
  NAND U25506 ( .A(n17130), .B(n17131), .Z(n17129) );
  NAND U25507 ( .A(n17132), .B(n17133), .Z(n17128) );
  AND U25508 ( .A(n17134), .B(n17135), .Z(n17089) );
  NAND U25509 ( .A(n17136), .B(n17137), .Z(n17135) );
  NAND U25510 ( .A(n17138), .B(n17139), .Z(n17134) );
  AND U25511 ( .A(n17140), .B(n17141), .Z(n17091) );
  NAND U25512 ( .A(n17142), .B(n17143), .Z(n17085) );
  XNOR U25513 ( .A(n17068), .B(n17144), .Z(n17082) );
  XNOR U25514 ( .A(n17072), .B(n17070), .Z(n17144) );
  XOR U25515 ( .A(n17078), .B(n17145), .Z(n17070) );
  XNOR U25516 ( .A(n17075), .B(n17079), .Z(n17145) );
  AND U25517 ( .A(n17146), .B(n17147), .Z(n17079) );
  NAND U25518 ( .A(n17148), .B(n17149), .Z(n17147) );
  NAND U25519 ( .A(n17150), .B(n17151), .Z(n17146) );
  AND U25520 ( .A(n17152), .B(n17153), .Z(n17075) );
  NAND U25521 ( .A(n17154), .B(n17155), .Z(n17153) );
  NAND U25522 ( .A(n17156), .B(n17157), .Z(n17152) );
  NANDN U25523 ( .A(n17158), .B(n17159), .Z(n17078) );
  ANDN U25524 ( .B(n17160), .A(n17161), .Z(n17072) );
  XNOR U25525 ( .A(n17063), .B(n17162), .Z(n17068) );
  XNOR U25526 ( .A(n17061), .B(n17065), .Z(n17162) );
  AND U25527 ( .A(n17163), .B(n17164), .Z(n17065) );
  NAND U25528 ( .A(n17165), .B(n17166), .Z(n17164) );
  NAND U25529 ( .A(n17167), .B(n17168), .Z(n17163) );
  AND U25530 ( .A(n17169), .B(n17170), .Z(n17061) );
  NAND U25531 ( .A(n17171), .B(n17172), .Z(n17170) );
  NAND U25532 ( .A(n17173), .B(n17174), .Z(n17169) );
  AND U25533 ( .A(n17175), .B(n17176), .Z(n17063) );
  XOR U25534 ( .A(n17143), .B(n17142), .Z(N63868) );
  XNOR U25535 ( .A(n17160), .B(n17161), .Z(n17142) );
  XNOR U25536 ( .A(n17175), .B(n17176), .Z(n17161) );
  XOR U25537 ( .A(n17172), .B(n17171), .Z(n17176) );
  XOR U25538 ( .A(y[6060]), .B(x[6060]), .Z(n17171) );
  XOR U25539 ( .A(n17174), .B(n17173), .Z(n17172) );
  XOR U25540 ( .A(y[6062]), .B(x[6062]), .Z(n17173) );
  XOR U25541 ( .A(y[6061]), .B(x[6061]), .Z(n17174) );
  XOR U25542 ( .A(n17166), .B(n17165), .Z(n17175) );
  XOR U25543 ( .A(n17168), .B(n17167), .Z(n17165) );
  XOR U25544 ( .A(y[6059]), .B(x[6059]), .Z(n17167) );
  XOR U25545 ( .A(y[6058]), .B(x[6058]), .Z(n17168) );
  XOR U25546 ( .A(y[6057]), .B(x[6057]), .Z(n17166) );
  XNOR U25547 ( .A(n17159), .B(n17158), .Z(n17160) );
  XNOR U25548 ( .A(n17155), .B(n17154), .Z(n17158) );
  XOR U25549 ( .A(n17157), .B(n17156), .Z(n17154) );
  XOR U25550 ( .A(y[6056]), .B(x[6056]), .Z(n17156) );
  XOR U25551 ( .A(y[6055]), .B(x[6055]), .Z(n17157) );
  XOR U25552 ( .A(y[6054]), .B(x[6054]), .Z(n17155) );
  XOR U25553 ( .A(n17149), .B(n17148), .Z(n17159) );
  XOR U25554 ( .A(n17151), .B(n17150), .Z(n17148) );
  XOR U25555 ( .A(y[6053]), .B(x[6053]), .Z(n17150) );
  XOR U25556 ( .A(y[6052]), .B(x[6052]), .Z(n17151) );
  XOR U25557 ( .A(y[6051]), .B(x[6051]), .Z(n17149) );
  XNOR U25558 ( .A(n17125), .B(n17126), .Z(n17143) );
  XNOR U25559 ( .A(n17140), .B(n17141), .Z(n17126) );
  XOR U25560 ( .A(n17137), .B(n17136), .Z(n17141) );
  XOR U25561 ( .A(y[6048]), .B(x[6048]), .Z(n17136) );
  XOR U25562 ( .A(n17139), .B(n17138), .Z(n17137) );
  XOR U25563 ( .A(y[6050]), .B(x[6050]), .Z(n17138) );
  XOR U25564 ( .A(y[6049]), .B(x[6049]), .Z(n17139) );
  XOR U25565 ( .A(n17131), .B(n17130), .Z(n17140) );
  XOR U25566 ( .A(n17133), .B(n17132), .Z(n17130) );
  XOR U25567 ( .A(y[6047]), .B(x[6047]), .Z(n17132) );
  XOR U25568 ( .A(y[6046]), .B(x[6046]), .Z(n17133) );
  XOR U25569 ( .A(y[6045]), .B(x[6045]), .Z(n17131) );
  XNOR U25570 ( .A(n17124), .B(n17123), .Z(n17125) );
  XNOR U25571 ( .A(n17120), .B(n17119), .Z(n17123) );
  XOR U25572 ( .A(n17122), .B(n17121), .Z(n17119) );
  XOR U25573 ( .A(y[6044]), .B(x[6044]), .Z(n17121) );
  XOR U25574 ( .A(y[6043]), .B(x[6043]), .Z(n17122) );
  XOR U25575 ( .A(y[6042]), .B(x[6042]), .Z(n17120) );
  XOR U25576 ( .A(n17114), .B(n17113), .Z(n17124) );
  XOR U25577 ( .A(n17116), .B(n17115), .Z(n17113) );
  XOR U25578 ( .A(y[6041]), .B(x[6041]), .Z(n17115) );
  XOR U25579 ( .A(y[6040]), .B(x[6040]), .Z(n17116) );
  XOR U25580 ( .A(y[6039]), .B(x[6039]), .Z(n17114) );
  NAND U25581 ( .A(n17177), .B(n17178), .Z(N63859) );
  NAND U25582 ( .A(n17179), .B(n17180), .Z(n17178) );
  NANDN U25583 ( .A(n17181), .B(n17182), .Z(n17180) );
  NANDN U25584 ( .A(n17182), .B(n17181), .Z(n17177) );
  XOR U25585 ( .A(n17181), .B(n17183), .Z(N63858) );
  XNOR U25586 ( .A(n17179), .B(n17182), .Z(n17183) );
  NAND U25587 ( .A(n17184), .B(n17185), .Z(n17182) );
  NAND U25588 ( .A(n17186), .B(n17187), .Z(n17185) );
  NANDN U25589 ( .A(n17188), .B(n17189), .Z(n17187) );
  NANDN U25590 ( .A(n17189), .B(n17188), .Z(n17184) );
  AND U25591 ( .A(n17190), .B(n17191), .Z(n17179) );
  NAND U25592 ( .A(n17192), .B(n17193), .Z(n17191) );
  NANDN U25593 ( .A(n17194), .B(n17195), .Z(n17193) );
  NANDN U25594 ( .A(n17195), .B(n17194), .Z(n17190) );
  IV U25595 ( .A(n17196), .Z(n17195) );
  AND U25596 ( .A(n17197), .B(n17198), .Z(n17181) );
  NAND U25597 ( .A(n17199), .B(n17200), .Z(n17198) );
  NANDN U25598 ( .A(n17201), .B(n17202), .Z(n17200) );
  NANDN U25599 ( .A(n17202), .B(n17201), .Z(n17197) );
  XOR U25600 ( .A(n17194), .B(n17203), .Z(N63857) );
  XNOR U25601 ( .A(n17192), .B(n17196), .Z(n17203) );
  XOR U25602 ( .A(n17189), .B(n17204), .Z(n17196) );
  XNOR U25603 ( .A(n17186), .B(n17188), .Z(n17204) );
  AND U25604 ( .A(n17205), .B(n17206), .Z(n17188) );
  NANDN U25605 ( .A(n17207), .B(n17208), .Z(n17206) );
  OR U25606 ( .A(n17209), .B(n17210), .Z(n17208) );
  IV U25607 ( .A(n17211), .Z(n17210) );
  NANDN U25608 ( .A(n17211), .B(n17209), .Z(n17205) );
  AND U25609 ( .A(n17212), .B(n17213), .Z(n17186) );
  NAND U25610 ( .A(n17214), .B(n17215), .Z(n17213) );
  NANDN U25611 ( .A(n17216), .B(n17217), .Z(n17215) );
  NANDN U25612 ( .A(n17217), .B(n17216), .Z(n17212) );
  IV U25613 ( .A(n17218), .Z(n17217) );
  NAND U25614 ( .A(n17219), .B(n17220), .Z(n17189) );
  NANDN U25615 ( .A(n17221), .B(n17222), .Z(n17220) );
  NANDN U25616 ( .A(n17223), .B(n17224), .Z(n17222) );
  NANDN U25617 ( .A(n17224), .B(n17223), .Z(n17219) );
  IV U25618 ( .A(n17225), .Z(n17223) );
  AND U25619 ( .A(n17226), .B(n17227), .Z(n17192) );
  NAND U25620 ( .A(n17228), .B(n17229), .Z(n17227) );
  NANDN U25621 ( .A(n17230), .B(n17231), .Z(n17229) );
  NANDN U25622 ( .A(n17231), .B(n17230), .Z(n17226) );
  XOR U25623 ( .A(n17202), .B(n17232), .Z(n17194) );
  XNOR U25624 ( .A(n17199), .B(n17201), .Z(n17232) );
  AND U25625 ( .A(n17233), .B(n17234), .Z(n17201) );
  NANDN U25626 ( .A(n17235), .B(n17236), .Z(n17234) );
  OR U25627 ( .A(n17237), .B(n17238), .Z(n17236) );
  IV U25628 ( .A(n17239), .Z(n17238) );
  NANDN U25629 ( .A(n17239), .B(n17237), .Z(n17233) );
  AND U25630 ( .A(n17240), .B(n17241), .Z(n17199) );
  NAND U25631 ( .A(n17242), .B(n17243), .Z(n17241) );
  NANDN U25632 ( .A(n17244), .B(n17245), .Z(n17243) );
  NANDN U25633 ( .A(n17245), .B(n17244), .Z(n17240) );
  IV U25634 ( .A(n17246), .Z(n17245) );
  NAND U25635 ( .A(n17247), .B(n17248), .Z(n17202) );
  NANDN U25636 ( .A(n17249), .B(n17250), .Z(n17248) );
  NANDN U25637 ( .A(n17251), .B(n17252), .Z(n17250) );
  NANDN U25638 ( .A(n17252), .B(n17251), .Z(n17247) );
  IV U25639 ( .A(n17253), .Z(n17251) );
  XOR U25640 ( .A(n17228), .B(n17254), .Z(N63856) );
  XNOR U25641 ( .A(n17231), .B(n17230), .Z(n17254) );
  XNOR U25642 ( .A(n17242), .B(n17255), .Z(n17230) );
  XNOR U25643 ( .A(n17246), .B(n17244), .Z(n17255) );
  XOR U25644 ( .A(n17252), .B(n17256), .Z(n17244) );
  XNOR U25645 ( .A(n17249), .B(n17253), .Z(n17256) );
  AND U25646 ( .A(n17257), .B(n17258), .Z(n17253) );
  NAND U25647 ( .A(n17259), .B(n17260), .Z(n17258) );
  NAND U25648 ( .A(n17261), .B(n17262), .Z(n17257) );
  AND U25649 ( .A(n17263), .B(n17264), .Z(n17249) );
  NAND U25650 ( .A(n17265), .B(n17266), .Z(n17264) );
  NAND U25651 ( .A(n17267), .B(n17268), .Z(n17263) );
  NANDN U25652 ( .A(n17269), .B(n17270), .Z(n17252) );
  ANDN U25653 ( .B(n17271), .A(n17272), .Z(n17246) );
  XNOR U25654 ( .A(n17237), .B(n17273), .Z(n17242) );
  XNOR U25655 ( .A(n17235), .B(n17239), .Z(n17273) );
  AND U25656 ( .A(n17274), .B(n17275), .Z(n17239) );
  NAND U25657 ( .A(n17276), .B(n17277), .Z(n17275) );
  NAND U25658 ( .A(n17278), .B(n17279), .Z(n17274) );
  AND U25659 ( .A(n17280), .B(n17281), .Z(n17235) );
  NAND U25660 ( .A(n17282), .B(n17283), .Z(n17281) );
  NAND U25661 ( .A(n17284), .B(n17285), .Z(n17280) );
  AND U25662 ( .A(n17286), .B(n17287), .Z(n17237) );
  NAND U25663 ( .A(n17288), .B(n17289), .Z(n17231) );
  XNOR U25664 ( .A(n17214), .B(n17290), .Z(n17228) );
  XNOR U25665 ( .A(n17218), .B(n17216), .Z(n17290) );
  XOR U25666 ( .A(n17224), .B(n17291), .Z(n17216) );
  XNOR U25667 ( .A(n17221), .B(n17225), .Z(n17291) );
  AND U25668 ( .A(n17292), .B(n17293), .Z(n17225) );
  NAND U25669 ( .A(n17294), .B(n17295), .Z(n17293) );
  NAND U25670 ( .A(n17296), .B(n17297), .Z(n17292) );
  AND U25671 ( .A(n17298), .B(n17299), .Z(n17221) );
  NAND U25672 ( .A(n17300), .B(n17301), .Z(n17299) );
  NAND U25673 ( .A(n17302), .B(n17303), .Z(n17298) );
  NANDN U25674 ( .A(n17304), .B(n17305), .Z(n17224) );
  ANDN U25675 ( .B(n17306), .A(n17307), .Z(n17218) );
  XNOR U25676 ( .A(n17209), .B(n17308), .Z(n17214) );
  XNOR U25677 ( .A(n17207), .B(n17211), .Z(n17308) );
  AND U25678 ( .A(n17309), .B(n17310), .Z(n17211) );
  NAND U25679 ( .A(n17311), .B(n17312), .Z(n17310) );
  NAND U25680 ( .A(n17313), .B(n17314), .Z(n17309) );
  AND U25681 ( .A(n17315), .B(n17316), .Z(n17207) );
  NAND U25682 ( .A(n17317), .B(n17318), .Z(n17316) );
  NAND U25683 ( .A(n17319), .B(n17320), .Z(n17315) );
  AND U25684 ( .A(n17321), .B(n17322), .Z(n17209) );
  XOR U25685 ( .A(n17289), .B(n17288), .Z(N63855) );
  XNOR U25686 ( .A(n17306), .B(n17307), .Z(n17288) );
  XNOR U25687 ( .A(n17321), .B(n17322), .Z(n17307) );
  XOR U25688 ( .A(n17318), .B(n17317), .Z(n17322) );
  XOR U25689 ( .A(y[6036]), .B(x[6036]), .Z(n17317) );
  XOR U25690 ( .A(n17320), .B(n17319), .Z(n17318) );
  XOR U25691 ( .A(y[6038]), .B(x[6038]), .Z(n17319) );
  XOR U25692 ( .A(y[6037]), .B(x[6037]), .Z(n17320) );
  XOR U25693 ( .A(n17312), .B(n17311), .Z(n17321) );
  XOR U25694 ( .A(n17314), .B(n17313), .Z(n17311) );
  XOR U25695 ( .A(y[6035]), .B(x[6035]), .Z(n17313) );
  XOR U25696 ( .A(y[6034]), .B(x[6034]), .Z(n17314) );
  XOR U25697 ( .A(y[6033]), .B(x[6033]), .Z(n17312) );
  XNOR U25698 ( .A(n17305), .B(n17304), .Z(n17306) );
  XNOR U25699 ( .A(n17301), .B(n17300), .Z(n17304) );
  XOR U25700 ( .A(n17303), .B(n17302), .Z(n17300) );
  XOR U25701 ( .A(y[6032]), .B(x[6032]), .Z(n17302) );
  XOR U25702 ( .A(y[6031]), .B(x[6031]), .Z(n17303) );
  XOR U25703 ( .A(y[6030]), .B(x[6030]), .Z(n17301) );
  XOR U25704 ( .A(n17295), .B(n17294), .Z(n17305) );
  XOR U25705 ( .A(n17297), .B(n17296), .Z(n17294) );
  XOR U25706 ( .A(y[6029]), .B(x[6029]), .Z(n17296) );
  XOR U25707 ( .A(y[6028]), .B(x[6028]), .Z(n17297) );
  XOR U25708 ( .A(y[6027]), .B(x[6027]), .Z(n17295) );
  XNOR U25709 ( .A(n17271), .B(n17272), .Z(n17289) );
  XNOR U25710 ( .A(n17286), .B(n17287), .Z(n17272) );
  XOR U25711 ( .A(n17283), .B(n17282), .Z(n17287) );
  XOR U25712 ( .A(y[6024]), .B(x[6024]), .Z(n17282) );
  XOR U25713 ( .A(n17285), .B(n17284), .Z(n17283) );
  XOR U25714 ( .A(y[6026]), .B(x[6026]), .Z(n17284) );
  XOR U25715 ( .A(y[6025]), .B(x[6025]), .Z(n17285) );
  XOR U25716 ( .A(n17277), .B(n17276), .Z(n17286) );
  XOR U25717 ( .A(n17279), .B(n17278), .Z(n17276) );
  XOR U25718 ( .A(y[6023]), .B(x[6023]), .Z(n17278) );
  XOR U25719 ( .A(y[6022]), .B(x[6022]), .Z(n17279) );
  XOR U25720 ( .A(y[6021]), .B(x[6021]), .Z(n17277) );
  XNOR U25721 ( .A(n17270), .B(n17269), .Z(n17271) );
  XNOR U25722 ( .A(n17266), .B(n17265), .Z(n17269) );
  XOR U25723 ( .A(n17268), .B(n17267), .Z(n17265) );
  XOR U25724 ( .A(y[6020]), .B(x[6020]), .Z(n17267) );
  XOR U25725 ( .A(y[6019]), .B(x[6019]), .Z(n17268) );
  XOR U25726 ( .A(y[6018]), .B(x[6018]), .Z(n17266) );
  XOR U25727 ( .A(n17260), .B(n17259), .Z(n17270) );
  XOR U25728 ( .A(n17262), .B(n17261), .Z(n17259) );
  XOR U25729 ( .A(y[6017]), .B(x[6017]), .Z(n17261) );
  XOR U25730 ( .A(y[6016]), .B(x[6016]), .Z(n17262) );
  XOR U25731 ( .A(y[6015]), .B(x[6015]), .Z(n17260) );
  NAND U25732 ( .A(n17323), .B(n17324), .Z(N63846) );
  NAND U25733 ( .A(n17325), .B(n17326), .Z(n17324) );
  NANDN U25734 ( .A(n17327), .B(n17328), .Z(n17326) );
  NANDN U25735 ( .A(n17328), .B(n17327), .Z(n17323) );
  XOR U25736 ( .A(n17327), .B(n17329), .Z(N63845) );
  XNOR U25737 ( .A(n17325), .B(n17328), .Z(n17329) );
  NAND U25738 ( .A(n17330), .B(n17331), .Z(n17328) );
  NAND U25739 ( .A(n17332), .B(n17333), .Z(n17331) );
  NANDN U25740 ( .A(n17334), .B(n17335), .Z(n17333) );
  NANDN U25741 ( .A(n17335), .B(n17334), .Z(n17330) );
  AND U25742 ( .A(n17336), .B(n17337), .Z(n17325) );
  NAND U25743 ( .A(n17338), .B(n17339), .Z(n17337) );
  NANDN U25744 ( .A(n17340), .B(n17341), .Z(n17339) );
  NANDN U25745 ( .A(n17341), .B(n17340), .Z(n17336) );
  IV U25746 ( .A(n17342), .Z(n17341) );
  AND U25747 ( .A(n17343), .B(n17344), .Z(n17327) );
  NAND U25748 ( .A(n17345), .B(n17346), .Z(n17344) );
  NANDN U25749 ( .A(n17347), .B(n17348), .Z(n17346) );
  NANDN U25750 ( .A(n17348), .B(n17347), .Z(n17343) );
  XOR U25751 ( .A(n17340), .B(n17349), .Z(N63844) );
  XNOR U25752 ( .A(n17338), .B(n17342), .Z(n17349) );
  XOR U25753 ( .A(n17335), .B(n17350), .Z(n17342) );
  XNOR U25754 ( .A(n17332), .B(n17334), .Z(n17350) );
  AND U25755 ( .A(n17351), .B(n17352), .Z(n17334) );
  NANDN U25756 ( .A(n17353), .B(n17354), .Z(n17352) );
  OR U25757 ( .A(n17355), .B(n17356), .Z(n17354) );
  IV U25758 ( .A(n17357), .Z(n17356) );
  NANDN U25759 ( .A(n17357), .B(n17355), .Z(n17351) );
  AND U25760 ( .A(n17358), .B(n17359), .Z(n17332) );
  NAND U25761 ( .A(n17360), .B(n17361), .Z(n17359) );
  NANDN U25762 ( .A(n17362), .B(n17363), .Z(n17361) );
  NANDN U25763 ( .A(n17363), .B(n17362), .Z(n17358) );
  IV U25764 ( .A(n17364), .Z(n17363) );
  NAND U25765 ( .A(n17365), .B(n17366), .Z(n17335) );
  NANDN U25766 ( .A(n17367), .B(n17368), .Z(n17366) );
  NANDN U25767 ( .A(n17369), .B(n17370), .Z(n17368) );
  NANDN U25768 ( .A(n17370), .B(n17369), .Z(n17365) );
  IV U25769 ( .A(n17371), .Z(n17369) );
  AND U25770 ( .A(n17372), .B(n17373), .Z(n17338) );
  NAND U25771 ( .A(n17374), .B(n17375), .Z(n17373) );
  NANDN U25772 ( .A(n17376), .B(n17377), .Z(n17375) );
  NANDN U25773 ( .A(n17377), .B(n17376), .Z(n17372) );
  XOR U25774 ( .A(n17348), .B(n17378), .Z(n17340) );
  XNOR U25775 ( .A(n17345), .B(n17347), .Z(n17378) );
  AND U25776 ( .A(n17379), .B(n17380), .Z(n17347) );
  NANDN U25777 ( .A(n17381), .B(n17382), .Z(n17380) );
  OR U25778 ( .A(n17383), .B(n17384), .Z(n17382) );
  IV U25779 ( .A(n17385), .Z(n17384) );
  NANDN U25780 ( .A(n17385), .B(n17383), .Z(n17379) );
  AND U25781 ( .A(n17386), .B(n17387), .Z(n17345) );
  NAND U25782 ( .A(n17388), .B(n17389), .Z(n17387) );
  NANDN U25783 ( .A(n17390), .B(n17391), .Z(n17389) );
  NANDN U25784 ( .A(n17391), .B(n17390), .Z(n17386) );
  IV U25785 ( .A(n17392), .Z(n17391) );
  NAND U25786 ( .A(n17393), .B(n17394), .Z(n17348) );
  NANDN U25787 ( .A(n17395), .B(n17396), .Z(n17394) );
  NANDN U25788 ( .A(n17397), .B(n17398), .Z(n17396) );
  NANDN U25789 ( .A(n17398), .B(n17397), .Z(n17393) );
  IV U25790 ( .A(n17399), .Z(n17397) );
  XOR U25791 ( .A(n17374), .B(n17400), .Z(N63843) );
  XNOR U25792 ( .A(n17377), .B(n17376), .Z(n17400) );
  XNOR U25793 ( .A(n17388), .B(n17401), .Z(n17376) );
  XNOR U25794 ( .A(n17392), .B(n17390), .Z(n17401) );
  XOR U25795 ( .A(n17398), .B(n17402), .Z(n17390) );
  XNOR U25796 ( .A(n17395), .B(n17399), .Z(n17402) );
  AND U25797 ( .A(n17403), .B(n17404), .Z(n17399) );
  NAND U25798 ( .A(n17405), .B(n17406), .Z(n17404) );
  NAND U25799 ( .A(n17407), .B(n17408), .Z(n17403) );
  AND U25800 ( .A(n17409), .B(n17410), .Z(n17395) );
  NAND U25801 ( .A(n17411), .B(n17412), .Z(n17410) );
  NAND U25802 ( .A(n17413), .B(n17414), .Z(n17409) );
  NANDN U25803 ( .A(n17415), .B(n17416), .Z(n17398) );
  ANDN U25804 ( .B(n17417), .A(n17418), .Z(n17392) );
  XNOR U25805 ( .A(n17383), .B(n17419), .Z(n17388) );
  XNOR U25806 ( .A(n17381), .B(n17385), .Z(n17419) );
  AND U25807 ( .A(n17420), .B(n17421), .Z(n17385) );
  NAND U25808 ( .A(n17422), .B(n17423), .Z(n17421) );
  NAND U25809 ( .A(n17424), .B(n17425), .Z(n17420) );
  AND U25810 ( .A(n17426), .B(n17427), .Z(n17381) );
  NAND U25811 ( .A(n17428), .B(n17429), .Z(n17427) );
  NAND U25812 ( .A(n17430), .B(n17431), .Z(n17426) );
  AND U25813 ( .A(n17432), .B(n17433), .Z(n17383) );
  NAND U25814 ( .A(n17434), .B(n17435), .Z(n17377) );
  XNOR U25815 ( .A(n17360), .B(n17436), .Z(n17374) );
  XNOR U25816 ( .A(n17364), .B(n17362), .Z(n17436) );
  XOR U25817 ( .A(n17370), .B(n17437), .Z(n17362) );
  XNOR U25818 ( .A(n17367), .B(n17371), .Z(n17437) );
  AND U25819 ( .A(n17438), .B(n17439), .Z(n17371) );
  NAND U25820 ( .A(n17440), .B(n17441), .Z(n17439) );
  NAND U25821 ( .A(n17442), .B(n17443), .Z(n17438) );
  AND U25822 ( .A(n17444), .B(n17445), .Z(n17367) );
  NAND U25823 ( .A(n17446), .B(n17447), .Z(n17445) );
  NAND U25824 ( .A(n17448), .B(n17449), .Z(n17444) );
  NANDN U25825 ( .A(n17450), .B(n17451), .Z(n17370) );
  ANDN U25826 ( .B(n17452), .A(n17453), .Z(n17364) );
  XNOR U25827 ( .A(n17355), .B(n17454), .Z(n17360) );
  XNOR U25828 ( .A(n17353), .B(n17357), .Z(n17454) );
  AND U25829 ( .A(n17455), .B(n17456), .Z(n17357) );
  NAND U25830 ( .A(n17457), .B(n17458), .Z(n17456) );
  NAND U25831 ( .A(n17459), .B(n17460), .Z(n17455) );
  AND U25832 ( .A(n17461), .B(n17462), .Z(n17353) );
  NAND U25833 ( .A(n17463), .B(n17464), .Z(n17462) );
  NAND U25834 ( .A(n17465), .B(n17466), .Z(n17461) );
  AND U25835 ( .A(n17467), .B(n17468), .Z(n17355) );
  XOR U25836 ( .A(n17435), .B(n17434), .Z(N63842) );
  XNOR U25837 ( .A(n17452), .B(n17453), .Z(n17434) );
  XNOR U25838 ( .A(n17467), .B(n17468), .Z(n17453) );
  XOR U25839 ( .A(n17464), .B(n17463), .Z(n17468) );
  XOR U25840 ( .A(y[6012]), .B(x[6012]), .Z(n17463) );
  XOR U25841 ( .A(n17466), .B(n17465), .Z(n17464) );
  XOR U25842 ( .A(y[6014]), .B(x[6014]), .Z(n17465) );
  XOR U25843 ( .A(y[6013]), .B(x[6013]), .Z(n17466) );
  XOR U25844 ( .A(n17458), .B(n17457), .Z(n17467) );
  XOR U25845 ( .A(n17460), .B(n17459), .Z(n17457) );
  XOR U25846 ( .A(y[6011]), .B(x[6011]), .Z(n17459) );
  XOR U25847 ( .A(y[6010]), .B(x[6010]), .Z(n17460) );
  XOR U25848 ( .A(y[6009]), .B(x[6009]), .Z(n17458) );
  XNOR U25849 ( .A(n17451), .B(n17450), .Z(n17452) );
  XNOR U25850 ( .A(n17447), .B(n17446), .Z(n17450) );
  XOR U25851 ( .A(n17449), .B(n17448), .Z(n17446) );
  XOR U25852 ( .A(y[6008]), .B(x[6008]), .Z(n17448) );
  XOR U25853 ( .A(y[6007]), .B(x[6007]), .Z(n17449) );
  XOR U25854 ( .A(y[6006]), .B(x[6006]), .Z(n17447) );
  XOR U25855 ( .A(n17441), .B(n17440), .Z(n17451) );
  XOR U25856 ( .A(n17443), .B(n17442), .Z(n17440) );
  XOR U25857 ( .A(y[6005]), .B(x[6005]), .Z(n17442) );
  XOR U25858 ( .A(y[6004]), .B(x[6004]), .Z(n17443) );
  XOR U25859 ( .A(y[6003]), .B(x[6003]), .Z(n17441) );
  XNOR U25860 ( .A(n17417), .B(n17418), .Z(n17435) );
  XNOR U25861 ( .A(n17432), .B(n17433), .Z(n17418) );
  XOR U25862 ( .A(n17429), .B(n17428), .Z(n17433) );
  XOR U25863 ( .A(y[6000]), .B(x[6000]), .Z(n17428) );
  XOR U25864 ( .A(n17431), .B(n17430), .Z(n17429) );
  XOR U25865 ( .A(y[6002]), .B(x[6002]), .Z(n17430) );
  XOR U25866 ( .A(y[6001]), .B(x[6001]), .Z(n17431) );
  XOR U25867 ( .A(n17423), .B(n17422), .Z(n17432) );
  XOR U25868 ( .A(n17425), .B(n17424), .Z(n17422) );
  XOR U25869 ( .A(y[5999]), .B(x[5999]), .Z(n17424) );
  XOR U25870 ( .A(y[5998]), .B(x[5998]), .Z(n17425) );
  XOR U25871 ( .A(y[5997]), .B(x[5997]), .Z(n17423) );
  XNOR U25872 ( .A(n17416), .B(n17415), .Z(n17417) );
  XNOR U25873 ( .A(n17412), .B(n17411), .Z(n17415) );
  XOR U25874 ( .A(n17414), .B(n17413), .Z(n17411) );
  XOR U25875 ( .A(y[5996]), .B(x[5996]), .Z(n17413) );
  XOR U25876 ( .A(y[5995]), .B(x[5995]), .Z(n17414) );
  XOR U25877 ( .A(y[5994]), .B(x[5994]), .Z(n17412) );
  XOR U25878 ( .A(n17406), .B(n17405), .Z(n17416) );
  XOR U25879 ( .A(n17408), .B(n17407), .Z(n17405) );
  XOR U25880 ( .A(y[5993]), .B(x[5993]), .Z(n17407) );
  XOR U25881 ( .A(y[5992]), .B(x[5992]), .Z(n17408) );
  XOR U25882 ( .A(y[5991]), .B(x[5991]), .Z(n17406) );
  NAND U25883 ( .A(n17469), .B(n17470), .Z(N63833) );
  NAND U25884 ( .A(n17471), .B(n17472), .Z(n17470) );
  NANDN U25885 ( .A(n17473), .B(n17474), .Z(n17472) );
  NANDN U25886 ( .A(n17474), .B(n17473), .Z(n17469) );
  XOR U25887 ( .A(n17473), .B(n17475), .Z(N63832) );
  XNOR U25888 ( .A(n17471), .B(n17474), .Z(n17475) );
  NAND U25889 ( .A(n17476), .B(n17477), .Z(n17474) );
  NAND U25890 ( .A(n17478), .B(n17479), .Z(n17477) );
  NANDN U25891 ( .A(n17480), .B(n17481), .Z(n17479) );
  NANDN U25892 ( .A(n17481), .B(n17480), .Z(n17476) );
  AND U25893 ( .A(n17482), .B(n17483), .Z(n17471) );
  NAND U25894 ( .A(n17484), .B(n17485), .Z(n17483) );
  NANDN U25895 ( .A(n17486), .B(n17487), .Z(n17485) );
  NANDN U25896 ( .A(n17487), .B(n17486), .Z(n17482) );
  IV U25897 ( .A(n17488), .Z(n17487) );
  AND U25898 ( .A(n17489), .B(n17490), .Z(n17473) );
  NAND U25899 ( .A(n17491), .B(n17492), .Z(n17490) );
  NANDN U25900 ( .A(n17493), .B(n17494), .Z(n17492) );
  NANDN U25901 ( .A(n17494), .B(n17493), .Z(n17489) );
  XOR U25902 ( .A(n17486), .B(n17495), .Z(N63831) );
  XNOR U25903 ( .A(n17484), .B(n17488), .Z(n17495) );
  XOR U25904 ( .A(n17481), .B(n17496), .Z(n17488) );
  XNOR U25905 ( .A(n17478), .B(n17480), .Z(n17496) );
  AND U25906 ( .A(n17497), .B(n17498), .Z(n17480) );
  NANDN U25907 ( .A(n17499), .B(n17500), .Z(n17498) );
  OR U25908 ( .A(n17501), .B(n17502), .Z(n17500) );
  IV U25909 ( .A(n17503), .Z(n17502) );
  NANDN U25910 ( .A(n17503), .B(n17501), .Z(n17497) );
  AND U25911 ( .A(n17504), .B(n17505), .Z(n17478) );
  NAND U25912 ( .A(n17506), .B(n17507), .Z(n17505) );
  NANDN U25913 ( .A(n17508), .B(n17509), .Z(n17507) );
  NANDN U25914 ( .A(n17509), .B(n17508), .Z(n17504) );
  IV U25915 ( .A(n17510), .Z(n17509) );
  NAND U25916 ( .A(n17511), .B(n17512), .Z(n17481) );
  NANDN U25917 ( .A(n17513), .B(n17514), .Z(n17512) );
  NANDN U25918 ( .A(n17515), .B(n17516), .Z(n17514) );
  NANDN U25919 ( .A(n17516), .B(n17515), .Z(n17511) );
  IV U25920 ( .A(n17517), .Z(n17515) );
  AND U25921 ( .A(n17518), .B(n17519), .Z(n17484) );
  NAND U25922 ( .A(n17520), .B(n17521), .Z(n17519) );
  NANDN U25923 ( .A(n17522), .B(n17523), .Z(n17521) );
  NANDN U25924 ( .A(n17523), .B(n17522), .Z(n17518) );
  XOR U25925 ( .A(n17494), .B(n17524), .Z(n17486) );
  XNOR U25926 ( .A(n17491), .B(n17493), .Z(n17524) );
  AND U25927 ( .A(n17525), .B(n17526), .Z(n17493) );
  NANDN U25928 ( .A(n17527), .B(n17528), .Z(n17526) );
  OR U25929 ( .A(n17529), .B(n17530), .Z(n17528) );
  IV U25930 ( .A(n17531), .Z(n17530) );
  NANDN U25931 ( .A(n17531), .B(n17529), .Z(n17525) );
  AND U25932 ( .A(n17532), .B(n17533), .Z(n17491) );
  NAND U25933 ( .A(n17534), .B(n17535), .Z(n17533) );
  NANDN U25934 ( .A(n17536), .B(n17537), .Z(n17535) );
  NANDN U25935 ( .A(n17537), .B(n17536), .Z(n17532) );
  IV U25936 ( .A(n17538), .Z(n17537) );
  NAND U25937 ( .A(n17539), .B(n17540), .Z(n17494) );
  NANDN U25938 ( .A(n17541), .B(n17542), .Z(n17540) );
  NANDN U25939 ( .A(n17543), .B(n17544), .Z(n17542) );
  NANDN U25940 ( .A(n17544), .B(n17543), .Z(n17539) );
  IV U25941 ( .A(n17545), .Z(n17543) );
  XOR U25942 ( .A(n17520), .B(n17546), .Z(N63830) );
  XNOR U25943 ( .A(n17523), .B(n17522), .Z(n17546) );
  XNOR U25944 ( .A(n17534), .B(n17547), .Z(n17522) );
  XNOR U25945 ( .A(n17538), .B(n17536), .Z(n17547) );
  XOR U25946 ( .A(n17544), .B(n17548), .Z(n17536) );
  XNOR U25947 ( .A(n17541), .B(n17545), .Z(n17548) );
  AND U25948 ( .A(n17549), .B(n17550), .Z(n17545) );
  NAND U25949 ( .A(n17551), .B(n17552), .Z(n17550) );
  NAND U25950 ( .A(n17553), .B(n17554), .Z(n17549) );
  AND U25951 ( .A(n17555), .B(n17556), .Z(n17541) );
  NAND U25952 ( .A(n17557), .B(n17558), .Z(n17556) );
  NAND U25953 ( .A(n17559), .B(n17560), .Z(n17555) );
  NANDN U25954 ( .A(n17561), .B(n17562), .Z(n17544) );
  ANDN U25955 ( .B(n17563), .A(n17564), .Z(n17538) );
  XNOR U25956 ( .A(n17529), .B(n17565), .Z(n17534) );
  XNOR U25957 ( .A(n17527), .B(n17531), .Z(n17565) );
  AND U25958 ( .A(n17566), .B(n17567), .Z(n17531) );
  NAND U25959 ( .A(n17568), .B(n17569), .Z(n17567) );
  NAND U25960 ( .A(n17570), .B(n17571), .Z(n17566) );
  AND U25961 ( .A(n17572), .B(n17573), .Z(n17527) );
  NAND U25962 ( .A(n17574), .B(n17575), .Z(n17573) );
  NAND U25963 ( .A(n17576), .B(n17577), .Z(n17572) );
  AND U25964 ( .A(n17578), .B(n17579), .Z(n17529) );
  NAND U25965 ( .A(n17580), .B(n17581), .Z(n17523) );
  XNOR U25966 ( .A(n17506), .B(n17582), .Z(n17520) );
  XNOR U25967 ( .A(n17510), .B(n17508), .Z(n17582) );
  XOR U25968 ( .A(n17516), .B(n17583), .Z(n17508) );
  XNOR U25969 ( .A(n17513), .B(n17517), .Z(n17583) );
  AND U25970 ( .A(n17584), .B(n17585), .Z(n17517) );
  NAND U25971 ( .A(n17586), .B(n17587), .Z(n17585) );
  NAND U25972 ( .A(n17588), .B(n17589), .Z(n17584) );
  AND U25973 ( .A(n17590), .B(n17591), .Z(n17513) );
  NAND U25974 ( .A(n17592), .B(n17593), .Z(n17591) );
  NAND U25975 ( .A(n17594), .B(n17595), .Z(n17590) );
  NANDN U25976 ( .A(n17596), .B(n17597), .Z(n17516) );
  ANDN U25977 ( .B(n17598), .A(n17599), .Z(n17510) );
  XNOR U25978 ( .A(n17501), .B(n17600), .Z(n17506) );
  XNOR U25979 ( .A(n17499), .B(n17503), .Z(n17600) );
  AND U25980 ( .A(n17601), .B(n17602), .Z(n17503) );
  NAND U25981 ( .A(n17603), .B(n17604), .Z(n17602) );
  NAND U25982 ( .A(n17605), .B(n17606), .Z(n17601) );
  AND U25983 ( .A(n17607), .B(n17608), .Z(n17499) );
  NAND U25984 ( .A(n17609), .B(n17610), .Z(n17608) );
  NAND U25985 ( .A(n17611), .B(n17612), .Z(n17607) );
  AND U25986 ( .A(n17613), .B(n17614), .Z(n17501) );
  XOR U25987 ( .A(n17581), .B(n17580), .Z(N63829) );
  XNOR U25988 ( .A(n17598), .B(n17599), .Z(n17580) );
  XNOR U25989 ( .A(n17613), .B(n17614), .Z(n17599) );
  XOR U25990 ( .A(n17610), .B(n17609), .Z(n17614) );
  XOR U25991 ( .A(y[5988]), .B(x[5988]), .Z(n17609) );
  XOR U25992 ( .A(n17612), .B(n17611), .Z(n17610) );
  XOR U25993 ( .A(y[5990]), .B(x[5990]), .Z(n17611) );
  XOR U25994 ( .A(y[5989]), .B(x[5989]), .Z(n17612) );
  XOR U25995 ( .A(n17604), .B(n17603), .Z(n17613) );
  XOR U25996 ( .A(n17606), .B(n17605), .Z(n17603) );
  XOR U25997 ( .A(y[5987]), .B(x[5987]), .Z(n17605) );
  XOR U25998 ( .A(y[5986]), .B(x[5986]), .Z(n17606) );
  XOR U25999 ( .A(y[5985]), .B(x[5985]), .Z(n17604) );
  XNOR U26000 ( .A(n17597), .B(n17596), .Z(n17598) );
  XNOR U26001 ( .A(n17593), .B(n17592), .Z(n17596) );
  XOR U26002 ( .A(n17595), .B(n17594), .Z(n17592) );
  XOR U26003 ( .A(y[5984]), .B(x[5984]), .Z(n17594) );
  XOR U26004 ( .A(y[5983]), .B(x[5983]), .Z(n17595) );
  XOR U26005 ( .A(y[5982]), .B(x[5982]), .Z(n17593) );
  XOR U26006 ( .A(n17587), .B(n17586), .Z(n17597) );
  XOR U26007 ( .A(n17589), .B(n17588), .Z(n17586) );
  XOR U26008 ( .A(y[5981]), .B(x[5981]), .Z(n17588) );
  XOR U26009 ( .A(y[5980]), .B(x[5980]), .Z(n17589) );
  XOR U26010 ( .A(y[5979]), .B(x[5979]), .Z(n17587) );
  XNOR U26011 ( .A(n17563), .B(n17564), .Z(n17581) );
  XNOR U26012 ( .A(n17578), .B(n17579), .Z(n17564) );
  XOR U26013 ( .A(n17575), .B(n17574), .Z(n17579) );
  XOR U26014 ( .A(y[5976]), .B(x[5976]), .Z(n17574) );
  XOR U26015 ( .A(n17577), .B(n17576), .Z(n17575) );
  XOR U26016 ( .A(y[5978]), .B(x[5978]), .Z(n17576) );
  XOR U26017 ( .A(y[5977]), .B(x[5977]), .Z(n17577) );
  XOR U26018 ( .A(n17569), .B(n17568), .Z(n17578) );
  XOR U26019 ( .A(n17571), .B(n17570), .Z(n17568) );
  XOR U26020 ( .A(y[5975]), .B(x[5975]), .Z(n17570) );
  XOR U26021 ( .A(y[5974]), .B(x[5974]), .Z(n17571) );
  XOR U26022 ( .A(y[5973]), .B(x[5973]), .Z(n17569) );
  XNOR U26023 ( .A(n17562), .B(n17561), .Z(n17563) );
  XNOR U26024 ( .A(n17558), .B(n17557), .Z(n17561) );
  XOR U26025 ( .A(n17560), .B(n17559), .Z(n17557) );
  XOR U26026 ( .A(y[5972]), .B(x[5972]), .Z(n17559) );
  XOR U26027 ( .A(y[5971]), .B(x[5971]), .Z(n17560) );
  XOR U26028 ( .A(y[5970]), .B(x[5970]), .Z(n17558) );
  XOR U26029 ( .A(n17552), .B(n17551), .Z(n17562) );
  XOR U26030 ( .A(n17554), .B(n17553), .Z(n17551) );
  XOR U26031 ( .A(y[5969]), .B(x[5969]), .Z(n17553) );
  XOR U26032 ( .A(y[5968]), .B(x[5968]), .Z(n17554) );
  XOR U26033 ( .A(y[5967]), .B(x[5967]), .Z(n17552) );
  NAND U26034 ( .A(n17615), .B(n17616), .Z(N63820) );
  NAND U26035 ( .A(n17617), .B(n17618), .Z(n17616) );
  NANDN U26036 ( .A(n17619), .B(n17620), .Z(n17618) );
  NANDN U26037 ( .A(n17620), .B(n17619), .Z(n17615) );
  XOR U26038 ( .A(n17619), .B(n17621), .Z(N63819) );
  XNOR U26039 ( .A(n17617), .B(n17620), .Z(n17621) );
  NAND U26040 ( .A(n17622), .B(n17623), .Z(n17620) );
  NAND U26041 ( .A(n17624), .B(n17625), .Z(n17623) );
  NANDN U26042 ( .A(n17626), .B(n17627), .Z(n17625) );
  NANDN U26043 ( .A(n17627), .B(n17626), .Z(n17622) );
  AND U26044 ( .A(n17628), .B(n17629), .Z(n17617) );
  NAND U26045 ( .A(n17630), .B(n17631), .Z(n17629) );
  NANDN U26046 ( .A(n17632), .B(n17633), .Z(n17631) );
  NANDN U26047 ( .A(n17633), .B(n17632), .Z(n17628) );
  IV U26048 ( .A(n17634), .Z(n17633) );
  AND U26049 ( .A(n17635), .B(n17636), .Z(n17619) );
  NAND U26050 ( .A(n17637), .B(n17638), .Z(n17636) );
  NANDN U26051 ( .A(n17639), .B(n17640), .Z(n17638) );
  NANDN U26052 ( .A(n17640), .B(n17639), .Z(n17635) );
  XOR U26053 ( .A(n17632), .B(n17641), .Z(N63818) );
  XNOR U26054 ( .A(n17630), .B(n17634), .Z(n17641) );
  XOR U26055 ( .A(n17627), .B(n17642), .Z(n17634) );
  XNOR U26056 ( .A(n17624), .B(n17626), .Z(n17642) );
  AND U26057 ( .A(n17643), .B(n17644), .Z(n17626) );
  NANDN U26058 ( .A(n17645), .B(n17646), .Z(n17644) );
  OR U26059 ( .A(n17647), .B(n17648), .Z(n17646) );
  IV U26060 ( .A(n17649), .Z(n17648) );
  NANDN U26061 ( .A(n17649), .B(n17647), .Z(n17643) );
  AND U26062 ( .A(n17650), .B(n17651), .Z(n17624) );
  NAND U26063 ( .A(n17652), .B(n17653), .Z(n17651) );
  NANDN U26064 ( .A(n17654), .B(n17655), .Z(n17653) );
  NANDN U26065 ( .A(n17655), .B(n17654), .Z(n17650) );
  IV U26066 ( .A(n17656), .Z(n17655) );
  NAND U26067 ( .A(n17657), .B(n17658), .Z(n17627) );
  NANDN U26068 ( .A(n17659), .B(n17660), .Z(n17658) );
  NANDN U26069 ( .A(n17661), .B(n17662), .Z(n17660) );
  NANDN U26070 ( .A(n17662), .B(n17661), .Z(n17657) );
  IV U26071 ( .A(n17663), .Z(n17661) );
  AND U26072 ( .A(n17664), .B(n17665), .Z(n17630) );
  NAND U26073 ( .A(n17666), .B(n17667), .Z(n17665) );
  NANDN U26074 ( .A(n17668), .B(n17669), .Z(n17667) );
  NANDN U26075 ( .A(n17669), .B(n17668), .Z(n17664) );
  XOR U26076 ( .A(n17640), .B(n17670), .Z(n17632) );
  XNOR U26077 ( .A(n17637), .B(n17639), .Z(n17670) );
  AND U26078 ( .A(n17671), .B(n17672), .Z(n17639) );
  NANDN U26079 ( .A(n17673), .B(n17674), .Z(n17672) );
  OR U26080 ( .A(n17675), .B(n17676), .Z(n17674) );
  IV U26081 ( .A(n17677), .Z(n17676) );
  NANDN U26082 ( .A(n17677), .B(n17675), .Z(n17671) );
  AND U26083 ( .A(n17678), .B(n17679), .Z(n17637) );
  NAND U26084 ( .A(n17680), .B(n17681), .Z(n17679) );
  NANDN U26085 ( .A(n17682), .B(n17683), .Z(n17681) );
  NANDN U26086 ( .A(n17683), .B(n17682), .Z(n17678) );
  IV U26087 ( .A(n17684), .Z(n17683) );
  NAND U26088 ( .A(n17685), .B(n17686), .Z(n17640) );
  NANDN U26089 ( .A(n17687), .B(n17688), .Z(n17686) );
  NANDN U26090 ( .A(n17689), .B(n17690), .Z(n17688) );
  NANDN U26091 ( .A(n17690), .B(n17689), .Z(n17685) );
  IV U26092 ( .A(n17691), .Z(n17689) );
  XOR U26093 ( .A(n17666), .B(n17692), .Z(N63817) );
  XNOR U26094 ( .A(n17669), .B(n17668), .Z(n17692) );
  XNOR U26095 ( .A(n17680), .B(n17693), .Z(n17668) );
  XNOR U26096 ( .A(n17684), .B(n17682), .Z(n17693) );
  XOR U26097 ( .A(n17690), .B(n17694), .Z(n17682) );
  XNOR U26098 ( .A(n17687), .B(n17691), .Z(n17694) );
  AND U26099 ( .A(n17695), .B(n17696), .Z(n17691) );
  NAND U26100 ( .A(n17697), .B(n17698), .Z(n17696) );
  NAND U26101 ( .A(n17699), .B(n17700), .Z(n17695) );
  AND U26102 ( .A(n17701), .B(n17702), .Z(n17687) );
  NAND U26103 ( .A(n17703), .B(n17704), .Z(n17702) );
  NAND U26104 ( .A(n17705), .B(n17706), .Z(n17701) );
  NANDN U26105 ( .A(n17707), .B(n17708), .Z(n17690) );
  ANDN U26106 ( .B(n17709), .A(n17710), .Z(n17684) );
  XNOR U26107 ( .A(n17675), .B(n17711), .Z(n17680) );
  XNOR U26108 ( .A(n17673), .B(n17677), .Z(n17711) );
  AND U26109 ( .A(n17712), .B(n17713), .Z(n17677) );
  NAND U26110 ( .A(n17714), .B(n17715), .Z(n17713) );
  NAND U26111 ( .A(n17716), .B(n17717), .Z(n17712) );
  AND U26112 ( .A(n17718), .B(n17719), .Z(n17673) );
  NAND U26113 ( .A(n17720), .B(n17721), .Z(n17719) );
  NAND U26114 ( .A(n17722), .B(n17723), .Z(n17718) );
  AND U26115 ( .A(n17724), .B(n17725), .Z(n17675) );
  NAND U26116 ( .A(n17726), .B(n17727), .Z(n17669) );
  XNOR U26117 ( .A(n17652), .B(n17728), .Z(n17666) );
  XNOR U26118 ( .A(n17656), .B(n17654), .Z(n17728) );
  XOR U26119 ( .A(n17662), .B(n17729), .Z(n17654) );
  XNOR U26120 ( .A(n17659), .B(n17663), .Z(n17729) );
  AND U26121 ( .A(n17730), .B(n17731), .Z(n17663) );
  NAND U26122 ( .A(n17732), .B(n17733), .Z(n17731) );
  NAND U26123 ( .A(n17734), .B(n17735), .Z(n17730) );
  AND U26124 ( .A(n17736), .B(n17737), .Z(n17659) );
  NAND U26125 ( .A(n17738), .B(n17739), .Z(n17737) );
  NAND U26126 ( .A(n17740), .B(n17741), .Z(n17736) );
  NANDN U26127 ( .A(n17742), .B(n17743), .Z(n17662) );
  ANDN U26128 ( .B(n17744), .A(n17745), .Z(n17656) );
  XNOR U26129 ( .A(n17647), .B(n17746), .Z(n17652) );
  XNOR U26130 ( .A(n17645), .B(n17649), .Z(n17746) );
  AND U26131 ( .A(n17747), .B(n17748), .Z(n17649) );
  NAND U26132 ( .A(n17749), .B(n17750), .Z(n17748) );
  NAND U26133 ( .A(n17751), .B(n17752), .Z(n17747) );
  AND U26134 ( .A(n17753), .B(n17754), .Z(n17645) );
  NAND U26135 ( .A(n17755), .B(n17756), .Z(n17754) );
  NAND U26136 ( .A(n17757), .B(n17758), .Z(n17753) );
  AND U26137 ( .A(n17759), .B(n17760), .Z(n17647) );
  XOR U26138 ( .A(n17727), .B(n17726), .Z(N63816) );
  XNOR U26139 ( .A(n17744), .B(n17745), .Z(n17726) );
  XNOR U26140 ( .A(n17759), .B(n17760), .Z(n17745) );
  XOR U26141 ( .A(n17756), .B(n17755), .Z(n17760) );
  XOR U26142 ( .A(y[5964]), .B(x[5964]), .Z(n17755) );
  XOR U26143 ( .A(n17758), .B(n17757), .Z(n17756) );
  XOR U26144 ( .A(y[5966]), .B(x[5966]), .Z(n17757) );
  XOR U26145 ( .A(y[5965]), .B(x[5965]), .Z(n17758) );
  XOR U26146 ( .A(n17750), .B(n17749), .Z(n17759) );
  XOR U26147 ( .A(n17752), .B(n17751), .Z(n17749) );
  XOR U26148 ( .A(y[5963]), .B(x[5963]), .Z(n17751) );
  XOR U26149 ( .A(y[5962]), .B(x[5962]), .Z(n17752) );
  XOR U26150 ( .A(y[5961]), .B(x[5961]), .Z(n17750) );
  XNOR U26151 ( .A(n17743), .B(n17742), .Z(n17744) );
  XNOR U26152 ( .A(n17739), .B(n17738), .Z(n17742) );
  XOR U26153 ( .A(n17741), .B(n17740), .Z(n17738) );
  XOR U26154 ( .A(y[5960]), .B(x[5960]), .Z(n17740) );
  XOR U26155 ( .A(y[5959]), .B(x[5959]), .Z(n17741) );
  XOR U26156 ( .A(y[5958]), .B(x[5958]), .Z(n17739) );
  XOR U26157 ( .A(n17733), .B(n17732), .Z(n17743) );
  XOR U26158 ( .A(n17735), .B(n17734), .Z(n17732) );
  XOR U26159 ( .A(y[5957]), .B(x[5957]), .Z(n17734) );
  XOR U26160 ( .A(y[5956]), .B(x[5956]), .Z(n17735) );
  XOR U26161 ( .A(y[5955]), .B(x[5955]), .Z(n17733) );
  XNOR U26162 ( .A(n17709), .B(n17710), .Z(n17727) );
  XNOR U26163 ( .A(n17724), .B(n17725), .Z(n17710) );
  XOR U26164 ( .A(n17721), .B(n17720), .Z(n17725) );
  XOR U26165 ( .A(y[5952]), .B(x[5952]), .Z(n17720) );
  XOR U26166 ( .A(n17723), .B(n17722), .Z(n17721) );
  XOR U26167 ( .A(y[5954]), .B(x[5954]), .Z(n17722) );
  XOR U26168 ( .A(y[5953]), .B(x[5953]), .Z(n17723) );
  XOR U26169 ( .A(n17715), .B(n17714), .Z(n17724) );
  XOR U26170 ( .A(n17717), .B(n17716), .Z(n17714) );
  XOR U26171 ( .A(y[5951]), .B(x[5951]), .Z(n17716) );
  XOR U26172 ( .A(y[5950]), .B(x[5950]), .Z(n17717) );
  XOR U26173 ( .A(y[5949]), .B(x[5949]), .Z(n17715) );
  XNOR U26174 ( .A(n17708), .B(n17707), .Z(n17709) );
  XNOR U26175 ( .A(n17704), .B(n17703), .Z(n17707) );
  XOR U26176 ( .A(n17706), .B(n17705), .Z(n17703) );
  XOR U26177 ( .A(y[5948]), .B(x[5948]), .Z(n17705) );
  XOR U26178 ( .A(y[5947]), .B(x[5947]), .Z(n17706) );
  XOR U26179 ( .A(y[5946]), .B(x[5946]), .Z(n17704) );
  XOR U26180 ( .A(n17698), .B(n17697), .Z(n17708) );
  XOR U26181 ( .A(n17700), .B(n17699), .Z(n17697) );
  XOR U26182 ( .A(y[5945]), .B(x[5945]), .Z(n17699) );
  XOR U26183 ( .A(y[5944]), .B(x[5944]), .Z(n17700) );
  XOR U26184 ( .A(y[5943]), .B(x[5943]), .Z(n17698) );
  NAND U26185 ( .A(n17761), .B(n17762), .Z(N63807) );
  NAND U26186 ( .A(n17763), .B(n17764), .Z(n17762) );
  NANDN U26187 ( .A(n17765), .B(n17766), .Z(n17764) );
  NANDN U26188 ( .A(n17766), .B(n17765), .Z(n17761) );
  XOR U26189 ( .A(n17765), .B(n17767), .Z(N63806) );
  XNOR U26190 ( .A(n17763), .B(n17766), .Z(n17767) );
  NAND U26191 ( .A(n17768), .B(n17769), .Z(n17766) );
  NAND U26192 ( .A(n17770), .B(n17771), .Z(n17769) );
  NANDN U26193 ( .A(n17772), .B(n17773), .Z(n17771) );
  NANDN U26194 ( .A(n17773), .B(n17772), .Z(n17768) );
  AND U26195 ( .A(n17774), .B(n17775), .Z(n17763) );
  NAND U26196 ( .A(n17776), .B(n17777), .Z(n17775) );
  NANDN U26197 ( .A(n17778), .B(n17779), .Z(n17777) );
  NANDN U26198 ( .A(n17779), .B(n17778), .Z(n17774) );
  IV U26199 ( .A(n17780), .Z(n17779) );
  AND U26200 ( .A(n17781), .B(n17782), .Z(n17765) );
  NAND U26201 ( .A(n17783), .B(n17784), .Z(n17782) );
  NANDN U26202 ( .A(n17785), .B(n17786), .Z(n17784) );
  NANDN U26203 ( .A(n17786), .B(n17785), .Z(n17781) );
  XOR U26204 ( .A(n17778), .B(n17787), .Z(N63805) );
  XNOR U26205 ( .A(n17776), .B(n17780), .Z(n17787) );
  XOR U26206 ( .A(n17773), .B(n17788), .Z(n17780) );
  XNOR U26207 ( .A(n17770), .B(n17772), .Z(n17788) );
  AND U26208 ( .A(n17789), .B(n17790), .Z(n17772) );
  NANDN U26209 ( .A(n17791), .B(n17792), .Z(n17790) );
  OR U26210 ( .A(n17793), .B(n17794), .Z(n17792) );
  IV U26211 ( .A(n17795), .Z(n17794) );
  NANDN U26212 ( .A(n17795), .B(n17793), .Z(n17789) );
  AND U26213 ( .A(n17796), .B(n17797), .Z(n17770) );
  NAND U26214 ( .A(n17798), .B(n17799), .Z(n17797) );
  NANDN U26215 ( .A(n17800), .B(n17801), .Z(n17799) );
  NANDN U26216 ( .A(n17801), .B(n17800), .Z(n17796) );
  IV U26217 ( .A(n17802), .Z(n17801) );
  NAND U26218 ( .A(n17803), .B(n17804), .Z(n17773) );
  NANDN U26219 ( .A(n17805), .B(n17806), .Z(n17804) );
  NANDN U26220 ( .A(n17807), .B(n17808), .Z(n17806) );
  NANDN U26221 ( .A(n17808), .B(n17807), .Z(n17803) );
  IV U26222 ( .A(n17809), .Z(n17807) );
  AND U26223 ( .A(n17810), .B(n17811), .Z(n17776) );
  NAND U26224 ( .A(n17812), .B(n17813), .Z(n17811) );
  NANDN U26225 ( .A(n17814), .B(n17815), .Z(n17813) );
  NANDN U26226 ( .A(n17815), .B(n17814), .Z(n17810) );
  XOR U26227 ( .A(n17786), .B(n17816), .Z(n17778) );
  XNOR U26228 ( .A(n17783), .B(n17785), .Z(n17816) );
  AND U26229 ( .A(n17817), .B(n17818), .Z(n17785) );
  NANDN U26230 ( .A(n17819), .B(n17820), .Z(n17818) );
  OR U26231 ( .A(n17821), .B(n17822), .Z(n17820) );
  IV U26232 ( .A(n17823), .Z(n17822) );
  NANDN U26233 ( .A(n17823), .B(n17821), .Z(n17817) );
  AND U26234 ( .A(n17824), .B(n17825), .Z(n17783) );
  NAND U26235 ( .A(n17826), .B(n17827), .Z(n17825) );
  NANDN U26236 ( .A(n17828), .B(n17829), .Z(n17827) );
  NANDN U26237 ( .A(n17829), .B(n17828), .Z(n17824) );
  IV U26238 ( .A(n17830), .Z(n17829) );
  NAND U26239 ( .A(n17831), .B(n17832), .Z(n17786) );
  NANDN U26240 ( .A(n17833), .B(n17834), .Z(n17832) );
  NANDN U26241 ( .A(n17835), .B(n17836), .Z(n17834) );
  NANDN U26242 ( .A(n17836), .B(n17835), .Z(n17831) );
  IV U26243 ( .A(n17837), .Z(n17835) );
  XOR U26244 ( .A(n17812), .B(n17838), .Z(N63804) );
  XNOR U26245 ( .A(n17815), .B(n17814), .Z(n17838) );
  XNOR U26246 ( .A(n17826), .B(n17839), .Z(n17814) );
  XNOR U26247 ( .A(n17830), .B(n17828), .Z(n17839) );
  XOR U26248 ( .A(n17836), .B(n17840), .Z(n17828) );
  XNOR U26249 ( .A(n17833), .B(n17837), .Z(n17840) );
  AND U26250 ( .A(n17841), .B(n17842), .Z(n17837) );
  NAND U26251 ( .A(n17843), .B(n17844), .Z(n17842) );
  NAND U26252 ( .A(n17845), .B(n17846), .Z(n17841) );
  AND U26253 ( .A(n17847), .B(n17848), .Z(n17833) );
  NAND U26254 ( .A(n17849), .B(n17850), .Z(n17848) );
  NAND U26255 ( .A(n17851), .B(n17852), .Z(n17847) );
  NANDN U26256 ( .A(n17853), .B(n17854), .Z(n17836) );
  ANDN U26257 ( .B(n17855), .A(n17856), .Z(n17830) );
  XNOR U26258 ( .A(n17821), .B(n17857), .Z(n17826) );
  XNOR U26259 ( .A(n17819), .B(n17823), .Z(n17857) );
  AND U26260 ( .A(n17858), .B(n17859), .Z(n17823) );
  NAND U26261 ( .A(n17860), .B(n17861), .Z(n17859) );
  NAND U26262 ( .A(n17862), .B(n17863), .Z(n17858) );
  AND U26263 ( .A(n17864), .B(n17865), .Z(n17819) );
  NAND U26264 ( .A(n17866), .B(n17867), .Z(n17865) );
  NAND U26265 ( .A(n17868), .B(n17869), .Z(n17864) );
  AND U26266 ( .A(n17870), .B(n17871), .Z(n17821) );
  NAND U26267 ( .A(n17872), .B(n17873), .Z(n17815) );
  XNOR U26268 ( .A(n17798), .B(n17874), .Z(n17812) );
  XNOR U26269 ( .A(n17802), .B(n17800), .Z(n17874) );
  XOR U26270 ( .A(n17808), .B(n17875), .Z(n17800) );
  XNOR U26271 ( .A(n17805), .B(n17809), .Z(n17875) );
  AND U26272 ( .A(n17876), .B(n17877), .Z(n17809) );
  NAND U26273 ( .A(n17878), .B(n17879), .Z(n17877) );
  NAND U26274 ( .A(n17880), .B(n17881), .Z(n17876) );
  AND U26275 ( .A(n17882), .B(n17883), .Z(n17805) );
  NAND U26276 ( .A(n17884), .B(n17885), .Z(n17883) );
  NAND U26277 ( .A(n17886), .B(n17887), .Z(n17882) );
  NANDN U26278 ( .A(n17888), .B(n17889), .Z(n17808) );
  ANDN U26279 ( .B(n17890), .A(n17891), .Z(n17802) );
  XNOR U26280 ( .A(n17793), .B(n17892), .Z(n17798) );
  XNOR U26281 ( .A(n17791), .B(n17795), .Z(n17892) );
  AND U26282 ( .A(n17893), .B(n17894), .Z(n17795) );
  NAND U26283 ( .A(n17895), .B(n17896), .Z(n17894) );
  NAND U26284 ( .A(n17897), .B(n17898), .Z(n17893) );
  AND U26285 ( .A(n17899), .B(n17900), .Z(n17791) );
  NAND U26286 ( .A(n17901), .B(n17902), .Z(n17900) );
  NAND U26287 ( .A(n17903), .B(n17904), .Z(n17899) );
  AND U26288 ( .A(n17905), .B(n17906), .Z(n17793) );
  XOR U26289 ( .A(n17873), .B(n17872), .Z(N63803) );
  XNOR U26290 ( .A(n17890), .B(n17891), .Z(n17872) );
  XNOR U26291 ( .A(n17905), .B(n17906), .Z(n17891) );
  XOR U26292 ( .A(n17902), .B(n17901), .Z(n17906) );
  XOR U26293 ( .A(y[5940]), .B(x[5940]), .Z(n17901) );
  XOR U26294 ( .A(n17904), .B(n17903), .Z(n17902) );
  XOR U26295 ( .A(y[5942]), .B(x[5942]), .Z(n17903) );
  XOR U26296 ( .A(y[5941]), .B(x[5941]), .Z(n17904) );
  XOR U26297 ( .A(n17896), .B(n17895), .Z(n17905) );
  XOR U26298 ( .A(n17898), .B(n17897), .Z(n17895) );
  XOR U26299 ( .A(y[5939]), .B(x[5939]), .Z(n17897) );
  XOR U26300 ( .A(y[5938]), .B(x[5938]), .Z(n17898) );
  XOR U26301 ( .A(y[5937]), .B(x[5937]), .Z(n17896) );
  XNOR U26302 ( .A(n17889), .B(n17888), .Z(n17890) );
  XNOR U26303 ( .A(n17885), .B(n17884), .Z(n17888) );
  XOR U26304 ( .A(n17887), .B(n17886), .Z(n17884) );
  XOR U26305 ( .A(y[5936]), .B(x[5936]), .Z(n17886) );
  XOR U26306 ( .A(y[5935]), .B(x[5935]), .Z(n17887) );
  XOR U26307 ( .A(y[5934]), .B(x[5934]), .Z(n17885) );
  XOR U26308 ( .A(n17879), .B(n17878), .Z(n17889) );
  XOR U26309 ( .A(n17881), .B(n17880), .Z(n17878) );
  XOR U26310 ( .A(y[5933]), .B(x[5933]), .Z(n17880) );
  XOR U26311 ( .A(y[5932]), .B(x[5932]), .Z(n17881) );
  XOR U26312 ( .A(y[5931]), .B(x[5931]), .Z(n17879) );
  XNOR U26313 ( .A(n17855), .B(n17856), .Z(n17873) );
  XNOR U26314 ( .A(n17870), .B(n17871), .Z(n17856) );
  XOR U26315 ( .A(n17867), .B(n17866), .Z(n17871) );
  XOR U26316 ( .A(y[5928]), .B(x[5928]), .Z(n17866) );
  XOR U26317 ( .A(n17869), .B(n17868), .Z(n17867) );
  XOR U26318 ( .A(y[5930]), .B(x[5930]), .Z(n17868) );
  XOR U26319 ( .A(y[5929]), .B(x[5929]), .Z(n17869) );
  XOR U26320 ( .A(n17861), .B(n17860), .Z(n17870) );
  XOR U26321 ( .A(n17863), .B(n17862), .Z(n17860) );
  XOR U26322 ( .A(y[5927]), .B(x[5927]), .Z(n17862) );
  XOR U26323 ( .A(y[5926]), .B(x[5926]), .Z(n17863) );
  XOR U26324 ( .A(y[5925]), .B(x[5925]), .Z(n17861) );
  XNOR U26325 ( .A(n17854), .B(n17853), .Z(n17855) );
  XNOR U26326 ( .A(n17850), .B(n17849), .Z(n17853) );
  XOR U26327 ( .A(n17852), .B(n17851), .Z(n17849) );
  XOR U26328 ( .A(y[5924]), .B(x[5924]), .Z(n17851) );
  XOR U26329 ( .A(y[5923]), .B(x[5923]), .Z(n17852) );
  XOR U26330 ( .A(y[5922]), .B(x[5922]), .Z(n17850) );
  XOR U26331 ( .A(n17844), .B(n17843), .Z(n17854) );
  XOR U26332 ( .A(n17846), .B(n17845), .Z(n17843) );
  XOR U26333 ( .A(y[5921]), .B(x[5921]), .Z(n17845) );
  XOR U26334 ( .A(y[5920]), .B(x[5920]), .Z(n17846) );
  XOR U26335 ( .A(y[5919]), .B(x[5919]), .Z(n17844) );
  NAND U26336 ( .A(n17907), .B(n17908), .Z(N63794) );
  NAND U26337 ( .A(n17909), .B(n17910), .Z(n17908) );
  NANDN U26338 ( .A(n17911), .B(n17912), .Z(n17910) );
  NANDN U26339 ( .A(n17912), .B(n17911), .Z(n17907) );
  XOR U26340 ( .A(n17911), .B(n17913), .Z(N63793) );
  XNOR U26341 ( .A(n17909), .B(n17912), .Z(n17913) );
  NAND U26342 ( .A(n17914), .B(n17915), .Z(n17912) );
  NAND U26343 ( .A(n17916), .B(n17917), .Z(n17915) );
  NANDN U26344 ( .A(n17918), .B(n17919), .Z(n17917) );
  NANDN U26345 ( .A(n17919), .B(n17918), .Z(n17914) );
  AND U26346 ( .A(n17920), .B(n17921), .Z(n17909) );
  NAND U26347 ( .A(n17922), .B(n17923), .Z(n17921) );
  NANDN U26348 ( .A(n17924), .B(n17925), .Z(n17923) );
  NANDN U26349 ( .A(n17925), .B(n17924), .Z(n17920) );
  IV U26350 ( .A(n17926), .Z(n17925) );
  AND U26351 ( .A(n17927), .B(n17928), .Z(n17911) );
  NAND U26352 ( .A(n17929), .B(n17930), .Z(n17928) );
  NANDN U26353 ( .A(n17931), .B(n17932), .Z(n17930) );
  NANDN U26354 ( .A(n17932), .B(n17931), .Z(n17927) );
  XOR U26355 ( .A(n17924), .B(n17933), .Z(N63792) );
  XNOR U26356 ( .A(n17922), .B(n17926), .Z(n17933) );
  XOR U26357 ( .A(n17919), .B(n17934), .Z(n17926) );
  XNOR U26358 ( .A(n17916), .B(n17918), .Z(n17934) );
  AND U26359 ( .A(n17935), .B(n17936), .Z(n17918) );
  NANDN U26360 ( .A(n17937), .B(n17938), .Z(n17936) );
  OR U26361 ( .A(n17939), .B(n17940), .Z(n17938) );
  IV U26362 ( .A(n17941), .Z(n17940) );
  NANDN U26363 ( .A(n17941), .B(n17939), .Z(n17935) );
  AND U26364 ( .A(n17942), .B(n17943), .Z(n17916) );
  NAND U26365 ( .A(n17944), .B(n17945), .Z(n17943) );
  NANDN U26366 ( .A(n17946), .B(n17947), .Z(n17945) );
  NANDN U26367 ( .A(n17947), .B(n17946), .Z(n17942) );
  IV U26368 ( .A(n17948), .Z(n17947) );
  NAND U26369 ( .A(n17949), .B(n17950), .Z(n17919) );
  NANDN U26370 ( .A(n17951), .B(n17952), .Z(n17950) );
  NANDN U26371 ( .A(n17953), .B(n17954), .Z(n17952) );
  NANDN U26372 ( .A(n17954), .B(n17953), .Z(n17949) );
  IV U26373 ( .A(n17955), .Z(n17953) );
  AND U26374 ( .A(n17956), .B(n17957), .Z(n17922) );
  NAND U26375 ( .A(n17958), .B(n17959), .Z(n17957) );
  NANDN U26376 ( .A(n17960), .B(n17961), .Z(n17959) );
  NANDN U26377 ( .A(n17961), .B(n17960), .Z(n17956) );
  XOR U26378 ( .A(n17932), .B(n17962), .Z(n17924) );
  XNOR U26379 ( .A(n17929), .B(n17931), .Z(n17962) );
  AND U26380 ( .A(n17963), .B(n17964), .Z(n17931) );
  NANDN U26381 ( .A(n17965), .B(n17966), .Z(n17964) );
  OR U26382 ( .A(n17967), .B(n17968), .Z(n17966) );
  IV U26383 ( .A(n17969), .Z(n17968) );
  NANDN U26384 ( .A(n17969), .B(n17967), .Z(n17963) );
  AND U26385 ( .A(n17970), .B(n17971), .Z(n17929) );
  NAND U26386 ( .A(n17972), .B(n17973), .Z(n17971) );
  NANDN U26387 ( .A(n17974), .B(n17975), .Z(n17973) );
  NANDN U26388 ( .A(n17975), .B(n17974), .Z(n17970) );
  IV U26389 ( .A(n17976), .Z(n17975) );
  NAND U26390 ( .A(n17977), .B(n17978), .Z(n17932) );
  NANDN U26391 ( .A(n17979), .B(n17980), .Z(n17978) );
  NANDN U26392 ( .A(n17981), .B(n17982), .Z(n17980) );
  NANDN U26393 ( .A(n17982), .B(n17981), .Z(n17977) );
  IV U26394 ( .A(n17983), .Z(n17981) );
  XOR U26395 ( .A(n17958), .B(n17984), .Z(N63791) );
  XNOR U26396 ( .A(n17961), .B(n17960), .Z(n17984) );
  XNOR U26397 ( .A(n17972), .B(n17985), .Z(n17960) );
  XNOR U26398 ( .A(n17976), .B(n17974), .Z(n17985) );
  XOR U26399 ( .A(n17982), .B(n17986), .Z(n17974) );
  XNOR U26400 ( .A(n17979), .B(n17983), .Z(n17986) );
  AND U26401 ( .A(n17987), .B(n17988), .Z(n17983) );
  NAND U26402 ( .A(n17989), .B(n17990), .Z(n17988) );
  NAND U26403 ( .A(n17991), .B(n17992), .Z(n17987) );
  AND U26404 ( .A(n17993), .B(n17994), .Z(n17979) );
  NAND U26405 ( .A(n17995), .B(n17996), .Z(n17994) );
  NAND U26406 ( .A(n17997), .B(n17998), .Z(n17993) );
  NANDN U26407 ( .A(n17999), .B(n18000), .Z(n17982) );
  ANDN U26408 ( .B(n18001), .A(n18002), .Z(n17976) );
  XNOR U26409 ( .A(n17967), .B(n18003), .Z(n17972) );
  XNOR U26410 ( .A(n17965), .B(n17969), .Z(n18003) );
  AND U26411 ( .A(n18004), .B(n18005), .Z(n17969) );
  NAND U26412 ( .A(n18006), .B(n18007), .Z(n18005) );
  NAND U26413 ( .A(n18008), .B(n18009), .Z(n18004) );
  AND U26414 ( .A(n18010), .B(n18011), .Z(n17965) );
  NAND U26415 ( .A(n18012), .B(n18013), .Z(n18011) );
  NAND U26416 ( .A(n18014), .B(n18015), .Z(n18010) );
  AND U26417 ( .A(n18016), .B(n18017), .Z(n17967) );
  NAND U26418 ( .A(n18018), .B(n18019), .Z(n17961) );
  XNOR U26419 ( .A(n17944), .B(n18020), .Z(n17958) );
  XNOR U26420 ( .A(n17948), .B(n17946), .Z(n18020) );
  XOR U26421 ( .A(n17954), .B(n18021), .Z(n17946) );
  XNOR U26422 ( .A(n17951), .B(n17955), .Z(n18021) );
  AND U26423 ( .A(n18022), .B(n18023), .Z(n17955) );
  NAND U26424 ( .A(n18024), .B(n18025), .Z(n18023) );
  NAND U26425 ( .A(n18026), .B(n18027), .Z(n18022) );
  AND U26426 ( .A(n18028), .B(n18029), .Z(n17951) );
  NAND U26427 ( .A(n18030), .B(n18031), .Z(n18029) );
  NAND U26428 ( .A(n18032), .B(n18033), .Z(n18028) );
  NANDN U26429 ( .A(n18034), .B(n18035), .Z(n17954) );
  ANDN U26430 ( .B(n18036), .A(n18037), .Z(n17948) );
  XNOR U26431 ( .A(n17939), .B(n18038), .Z(n17944) );
  XNOR U26432 ( .A(n17937), .B(n17941), .Z(n18038) );
  AND U26433 ( .A(n18039), .B(n18040), .Z(n17941) );
  NAND U26434 ( .A(n18041), .B(n18042), .Z(n18040) );
  NAND U26435 ( .A(n18043), .B(n18044), .Z(n18039) );
  AND U26436 ( .A(n18045), .B(n18046), .Z(n17937) );
  NAND U26437 ( .A(n18047), .B(n18048), .Z(n18046) );
  NAND U26438 ( .A(n18049), .B(n18050), .Z(n18045) );
  AND U26439 ( .A(n18051), .B(n18052), .Z(n17939) );
  XOR U26440 ( .A(n18019), .B(n18018), .Z(N63790) );
  XNOR U26441 ( .A(n18036), .B(n18037), .Z(n18018) );
  XNOR U26442 ( .A(n18051), .B(n18052), .Z(n18037) );
  XOR U26443 ( .A(n18048), .B(n18047), .Z(n18052) );
  XOR U26444 ( .A(y[5916]), .B(x[5916]), .Z(n18047) );
  XOR U26445 ( .A(n18050), .B(n18049), .Z(n18048) );
  XOR U26446 ( .A(y[5918]), .B(x[5918]), .Z(n18049) );
  XOR U26447 ( .A(y[5917]), .B(x[5917]), .Z(n18050) );
  XOR U26448 ( .A(n18042), .B(n18041), .Z(n18051) );
  XOR U26449 ( .A(n18044), .B(n18043), .Z(n18041) );
  XOR U26450 ( .A(y[5915]), .B(x[5915]), .Z(n18043) );
  XOR U26451 ( .A(y[5914]), .B(x[5914]), .Z(n18044) );
  XOR U26452 ( .A(y[5913]), .B(x[5913]), .Z(n18042) );
  XNOR U26453 ( .A(n18035), .B(n18034), .Z(n18036) );
  XNOR U26454 ( .A(n18031), .B(n18030), .Z(n18034) );
  XOR U26455 ( .A(n18033), .B(n18032), .Z(n18030) );
  XOR U26456 ( .A(y[5912]), .B(x[5912]), .Z(n18032) );
  XOR U26457 ( .A(y[5911]), .B(x[5911]), .Z(n18033) );
  XOR U26458 ( .A(y[5910]), .B(x[5910]), .Z(n18031) );
  XOR U26459 ( .A(n18025), .B(n18024), .Z(n18035) );
  XOR U26460 ( .A(n18027), .B(n18026), .Z(n18024) );
  XOR U26461 ( .A(y[5909]), .B(x[5909]), .Z(n18026) );
  XOR U26462 ( .A(y[5908]), .B(x[5908]), .Z(n18027) );
  XOR U26463 ( .A(y[5907]), .B(x[5907]), .Z(n18025) );
  XNOR U26464 ( .A(n18001), .B(n18002), .Z(n18019) );
  XNOR U26465 ( .A(n18016), .B(n18017), .Z(n18002) );
  XOR U26466 ( .A(n18013), .B(n18012), .Z(n18017) );
  XOR U26467 ( .A(y[5904]), .B(x[5904]), .Z(n18012) );
  XOR U26468 ( .A(n18015), .B(n18014), .Z(n18013) );
  XOR U26469 ( .A(y[5906]), .B(x[5906]), .Z(n18014) );
  XOR U26470 ( .A(y[5905]), .B(x[5905]), .Z(n18015) );
  XOR U26471 ( .A(n18007), .B(n18006), .Z(n18016) );
  XOR U26472 ( .A(n18009), .B(n18008), .Z(n18006) );
  XOR U26473 ( .A(y[5903]), .B(x[5903]), .Z(n18008) );
  XOR U26474 ( .A(y[5902]), .B(x[5902]), .Z(n18009) );
  XOR U26475 ( .A(y[5901]), .B(x[5901]), .Z(n18007) );
  XNOR U26476 ( .A(n18000), .B(n17999), .Z(n18001) );
  XNOR U26477 ( .A(n17996), .B(n17995), .Z(n17999) );
  XOR U26478 ( .A(n17998), .B(n17997), .Z(n17995) );
  XOR U26479 ( .A(y[5900]), .B(x[5900]), .Z(n17997) );
  XOR U26480 ( .A(y[5899]), .B(x[5899]), .Z(n17998) );
  XOR U26481 ( .A(y[5898]), .B(x[5898]), .Z(n17996) );
  XOR U26482 ( .A(n17990), .B(n17989), .Z(n18000) );
  XOR U26483 ( .A(n17992), .B(n17991), .Z(n17989) );
  XOR U26484 ( .A(y[5897]), .B(x[5897]), .Z(n17991) );
  XOR U26485 ( .A(y[5896]), .B(x[5896]), .Z(n17992) );
  XOR U26486 ( .A(y[5895]), .B(x[5895]), .Z(n17990) );
  NAND U26487 ( .A(n18053), .B(n18054), .Z(N63781) );
  NAND U26488 ( .A(n18055), .B(n18056), .Z(n18054) );
  NANDN U26489 ( .A(n18057), .B(n18058), .Z(n18056) );
  NANDN U26490 ( .A(n18058), .B(n18057), .Z(n18053) );
  XOR U26491 ( .A(n18057), .B(n18059), .Z(N63780) );
  XNOR U26492 ( .A(n18055), .B(n18058), .Z(n18059) );
  NAND U26493 ( .A(n18060), .B(n18061), .Z(n18058) );
  NAND U26494 ( .A(n18062), .B(n18063), .Z(n18061) );
  NANDN U26495 ( .A(n18064), .B(n18065), .Z(n18063) );
  NANDN U26496 ( .A(n18065), .B(n18064), .Z(n18060) );
  AND U26497 ( .A(n18066), .B(n18067), .Z(n18055) );
  NAND U26498 ( .A(n18068), .B(n18069), .Z(n18067) );
  NANDN U26499 ( .A(n18070), .B(n18071), .Z(n18069) );
  NANDN U26500 ( .A(n18071), .B(n18070), .Z(n18066) );
  IV U26501 ( .A(n18072), .Z(n18071) );
  AND U26502 ( .A(n18073), .B(n18074), .Z(n18057) );
  NAND U26503 ( .A(n18075), .B(n18076), .Z(n18074) );
  NANDN U26504 ( .A(n18077), .B(n18078), .Z(n18076) );
  NANDN U26505 ( .A(n18078), .B(n18077), .Z(n18073) );
  XOR U26506 ( .A(n18070), .B(n18079), .Z(N63779) );
  XNOR U26507 ( .A(n18068), .B(n18072), .Z(n18079) );
  XOR U26508 ( .A(n18065), .B(n18080), .Z(n18072) );
  XNOR U26509 ( .A(n18062), .B(n18064), .Z(n18080) );
  AND U26510 ( .A(n18081), .B(n18082), .Z(n18064) );
  NANDN U26511 ( .A(n18083), .B(n18084), .Z(n18082) );
  OR U26512 ( .A(n18085), .B(n18086), .Z(n18084) );
  IV U26513 ( .A(n18087), .Z(n18086) );
  NANDN U26514 ( .A(n18087), .B(n18085), .Z(n18081) );
  AND U26515 ( .A(n18088), .B(n18089), .Z(n18062) );
  NAND U26516 ( .A(n18090), .B(n18091), .Z(n18089) );
  NANDN U26517 ( .A(n18092), .B(n18093), .Z(n18091) );
  NANDN U26518 ( .A(n18093), .B(n18092), .Z(n18088) );
  IV U26519 ( .A(n18094), .Z(n18093) );
  NAND U26520 ( .A(n18095), .B(n18096), .Z(n18065) );
  NANDN U26521 ( .A(n18097), .B(n18098), .Z(n18096) );
  NANDN U26522 ( .A(n18099), .B(n18100), .Z(n18098) );
  NANDN U26523 ( .A(n18100), .B(n18099), .Z(n18095) );
  IV U26524 ( .A(n18101), .Z(n18099) );
  AND U26525 ( .A(n18102), .B(n18103), .Z(n18068) );
  NAND U26526 ( .A(n18104), .B(n18105), .Z(n18103) );
  NANDN U26527 ( .A(n18106), .B(n18107), .Z(n18105) );
  NANDN U26528 ( .A(n18107), .B(n18106), .Z(n18102) );
  XOR U26529 ( .A(n18078), .B(n18108), .Z(n18070) );
  XNOR U26530 ( .A(n18075), .B(n18077), .Z(n18108) );
  AND U26531 ( .A(n18109), .B(n18110), .Z(n18077) );
  NANDN U26532 ( .A(n18111), .B(n18112), .Z(n18110) );
  OR U26533 ( .A(n18113), .B(n18114), .Z(n18112) );
  IV U26534 ( .A(n18115), .Z(n18114) );
  NANDN U26535 ( .A(n18115), .B(n18113), .Z(n18109) );
  AND U26536 ( .A(n18116), .B(n18117), .Z(n18075) );
  NAND U26537 ( .A(n18118), .B(n18119), .Z(n18117) );
  NANDN U26538 ( .A(n18120), .B(n18121), .Z(n18119) );
  NANDN U26539 ( .A(n18121), .B(n18120), .Z(n18116) );
  IV U26540 ( .A(n18122), .Z(n18121) );
  NAND U26541 ( .A(n18123), .B(n18124), .Z(n18078) );
  NANDN U26542 ( .A(n18125), .B(n18126), .Z(n18124) );
  NANDN U26543 ( .A(n18127), .B(n18128), .Z(n18126) );
  NANDN U26544 ( .A(n18128), .B(n18127), .Z(n18123) );
  IV U26545 ( .A(n18129), .Z(n18127) );
  XOR U26546 ( .A(n18104), .B(n18130), .Z(N63778) );
  XNOR U26547 ( .A(n18107), .B(n18106), .Z(n18130) );
  XNOR U26548 ( .A(n18118), .B(n18131), .Z(n18106) );
  XNOR U26549 ( .A(n18122), .B(n18120), .Z(n18131) );
  XOR U26550 ( .A(n18128), .B(n18132), .Z(n18120) );
  XNOR U26551 ( .A(n18125), .B(n18129), .Z(n18132) );
  AND U26552 ( .A(n18133), .B(n18134), .Z(n18129) );
  NAND U26553 ( .A(n18135), .B(n18136), .Z(n18134) );
  NAND U26554 ( .A(n18137), .B(n18138), .Z(n18133) );
  AND U26555 ( .A(n18139), .B(n18140), .Z(n18125) );
  NAND U26556 ( .A(n18141), .B(n18142), .Z(n18140) );
  NAND U26557 ( .A(n18143), .B(n18144), .Z(n18139) );
  NANDN U26558 ( .A(n18145), .B(n18146), .Z(n18128) );
  ANDN U26559 ( .B(n18147), .A(n18148), .Z(n18122) );
  XNOR U26560 ( .A(n18113), .B(n18149), .Z(n18118) );
  XNOR U26561 ( .A(n18111), .B(n18115), .Z(n18149) );
  AND U26562 ( .A(n18150), .B(n18151), .Z(n18115) );
  NAND U26563 ( .A(n18152), .B(n18153), .Z(n18151) );
  NAND U26564 ( .A(n18154), .B(n18155), .Z(n18150) );
  AND U26565 ( .A(n18156), .B(n18157), .Z(n18111) );
  NAND U26566 ( .A(n18158), .B(n18159), .Z(n18157) );
  NAND U26567 ( .A(n18160), .B(n18161), .Z(n18156) );
  AND U26568 ( .A(n18162), .B(n18163), .Z(n18113) );
  NAND U26569 ( .A(n18164), .B(n18165), .Z(n18107) );
  XNOR U26570 ( .A(n18090), .B(n18166), .Z(n18104) );
  XNOR U26571 ( .A(n18094), .B(n18092), .Z(n18166) );
  XOR U26572 ( .A(n18100), .B(n18167), .Z(n18092) );
  XNOR U26573 ( .A(n18097), .B(n18101), .Z(n18167) );
  AND U26574 ( .A(n18168), .B(n18169), .Z(n18101) );
  NAND U26575 ( .A(n18170), .B(n18171), .Z(n18169) );
  NAND U26576 ( .A(n18172), .B(n18173), .Z(n18168) );
  AND U26577 ( .A(n18174), .B(n18175), .Z(n18097) );
  NAND U26578 ( .A(n18176), .B(n18177), .Z(n18175) );
  NAND U26579 ( .A(n18178), .B(n18179), .Z(n18174) );
  NANDN U26580 ( .A(n18180), .B(n18181), .Z(n18100) );
  ANDN U26581 ( .B(n18182), .A(n18183), .Z(n18094) );
  XNOR U26582 ( .A(n18085), .B(n18184), .Z(n18090) );
  XNOR U26583 ( .A(n18083), .B(n18087), .Z(n18184) );
  AND U26584 ( .A(n18185), .B(n18186), .Z(n18087) );
  NAND U26585 ( .A(n18187), .B(n18188), .Z(n18186) );
  NAND U26586 ( .A(n18189), .B(n18190), .Z(n18185) );
  AND U26587 ( .A(n18191), .B(n18192), .Z(n18083) );
  NAND U26588 ( .A(n18193), .B(n18194), .Z(n18192) );
  NAND U26589 ( .A(n18195), .B(n18196), .Z(n18191) );
  AND U26590 ( .A(n18197), .B(n18198), .Z(n18085) );
  XOR U26591 ( .A(n18165), .B(n18164), .Z(N63777) );
  XNOR U26592 ( .A(n18182), .B(n18183), .Z(n18164) );
  XNOR U26593 ( .A(n18197), .B(n18198), .Z(n18183) );
  XOR U26594 ( .A(n18194), .B(n18193), .Z(n18198) );
  XOR U26595 ( .A(y[5892]), .B(x[5892]), .Z(n18193) );
  XOR U26596 ( .A(n18196), .B(n18195), .Z(n18194) );
  XOR U26597 ( .A(y[5894]), .B(x[5894]), .Z(n18195) );
  XOR U26598 ( .A(y[5893]), .B(x[5893]), .Z(n18196) );
  XOR U26599 ( .A(n18188), .B(n18187), .Z(n18197) );
  XOR U26600 ( .A(n18190), .B(n18189), .Z(n18187) );
  XOR U26601 ( .A(y[5891]), .B(x[5891]), .Z(n18189) );
  XOR U26602 ( .A(y[5890]), .B(x[5890]), .Z(n18190) );
  XOR U26603 ( .A(y[5889]), .B(x[5889]), .Z(n18188) );
  XNOR U26604 ( .A(n18181), .B(n18180), .Z(n18182) );
  XNOR U26605 ( .A(n18177), .B(n18176), .Z(n18180) );
  XOR U26606 ( .A(n18179), .B(n18178), .Z(n18176) );
  XOR U26607 ( .A(y[5888]), .B(x[5888]), .Z(n18178) );
  XOR U26608 ( .A(y[5887]), .B(x[5887]), .Z(n18179) );
  XOR U26609 ( .A(y[5886]), .B(x[5886]), .Z(n18177) );
  XOR U26610 ( .A(n18171), .B(n18170), .Z(n18181) );
  XOR U26611 ( .A(n18173), .B(n18172), .Z(n18170) );
  XOR U26612 ( .A(y[5885]), .B(x[5885]), .Z(n18172) );
  XOR U26613 ( .A(y[5884]), .B(x[5884]), .Z(n18173) );
  XOR U26614 ( .A(y[5883]), .B(x[5883]), .Z(n18171) );
  XNOR U26615 ( .A(n18147), .B(n18148), .Z(n18165) );
  XNOR U26616 ( .A(n18162), .B(n18163), .Z(n18148) );
  XOR U26617 ( .A(n18159), .B(n18158), .Z(n18163) );
  XOR U26618 ( .A(y[5880]), .B(x[5880]), .Z(n18158) );
  XOR U26619 ( .A(n18161), .B(n18160), .Z(n18159) );
  XOR U26620 ( .A(y[5882]), .B(x[5882]), .Z(n18160) );
  XOR U26621 ( .A(y[5881]), .B(x[5881]), .Z(n18161) );
  XOR U26622 ( .A(n18153), .B(n18152), .Z(n18162) );
  XOR U26623 ( .A(n18155), .B(n18154), .Z(n18152) );
  XOR U26624 ( .A(y[5879]), .B(x[5879]), .Z(n18154) );
  XOR U26625 ( .A(y[5878]), .B(x[5878]), .Z(n18155) );
  XOR U26626 ( .A(y[5877]), .B(x[5877]), .Z(n18153) );
  XNOR U26627 ( .A(n18146), .B(n18145), .Z(n18147) );
  XNOR U26628 ( .A(n18142), .B(n18141), .Z(n18145) );
  XOR U26629 ( .A(n18144), .B(n18143), .Z(n18141) );
  XOR U26630 ( .A(y[5876]), .B(x[5876]), .Z(n18143) );
  XOR U26631 ( .A(y[5875]), .B(x[5875]), .Z(n18144) );
  XOR U26632 ( .A(y[5874]), .B(x[5874]), .Z(n18142) );
  XOR U26633 ( .A(n18136), .B(n18135), .Z(n18146) );
  XOR U26634 ( .A(n18138), .B(n18137), .Z(n18135) );
  XOR U26635 ( .A(y[5873]), .B(x[5873]), .Z(n18137) );
  XOR U26636 ( .A(y[5872]), .B(x[5872]), .Z(n18138) );
  XOR U26637 ( .A(y[5871]), .B(x[5871]), .Z(n18136) );
  NAND U26638 ( .A(n18199), .B(n18200), .Z(N63768) );
  NAND U26639 ( .A(n18201), .B(n18202), .Z(n18200) );
  NANDN U26640 ( .A(n18203), .B(n18204), .Z(n18202) );
  NANDN U26641 ( .A(n18204), .B(n18203), .Z(n18199) );
  XOR U26642 ( .A(n18203), .B(n18205), .Z(N63767) );
  XNOR U26643 ( .A(n18201), .B(n18204), .Z(n18205) );
  NAND U26644 ( .A(n18206), .B(n18207), .Z(n18204) );
  NAND U26645 ( .A(n18208), .B(n18209), .Z(n18207) );
  NANDN U26646 ( .A(n18210), .B(n18211), .Z(n18209) );
  NANDN U26647 ( .A(n18211), .B(n18210), .Z(n18206) );
  AND U26648 ( .A(n18212), .B(n18213), .Z(n18201) );
  NAND U26649 ( .A(n18214), .B(n18215), .Z(n18213) );
  NANDN U26650 ( .A(n18216), .B(n18217), .Z(n18215) );
  NANDN U26651 ( .A(n18217), .B(n18216), .Z(n18212) );
  IV U26652 ( .A(n18218), .Z(n18217) );
  AND U26653 ( .A(n18219), .B(n18220), .Z(n18203) );
  NAND U26654 ( .A(n18221), .B(n18222), .Z(n18220) );
  NANDN U26655 ( .A(n18223), .B(n18224), .Z(n18222) );
  NANDN U26656 ( .A(n18224), .B(n18223), .Z(n18219) );
  XOR U26657 ( .A(n18216), .B(n18225), .Z(N63766) );
  XNOR U26658 ( .A(n18214), .B(n18218), .Z(n18225) );
  XOR U26659 ( .A(n18211), .B(n18226), .Z(n18218) );
  XNOR U26660 ( .A(n18208), .B(n18210), .Z(n18226) );
  AND U26661 ( .A(n18227), .B(n18228), .Z(n18210) );
  NANDN U26662 ( .A(n18229), .B(n18230), .Z(n18228) );
  OR U26663 ( .A(n18231), .B(n18232), .Z(n18230) );
  IV U26664 ( .A(n18233), .Z(n18232) );
  NANDN U26665 ( .A(n18233), .B(n18231), .Z(n18227) );
  AND U26666 ( .A(n18234), .B(n18235), .Z(n18208) );
  NAND U26667 ( .A(n18236), .B(n18237), .Z(n18235) );
  NANDN U26668 ( .A(n18238), .B(n18239), .Z(n18237) );
  NANDN U26669 ( .A(n18239), .B(n18238), .Z(n18234) );
  IV U26670 ( .A(n18240), .Z(n18239) );
  NAND U26671 ( .A(n18241), .B(n18242), .Z(n18211) );
  NANDN U26672 ( .A(n18243), .B(n18244), .Z(n18242) );
  NANDN U26673 ( .A(n18245), .B(n18246), .Z(n18244) );
  NANDN U26674 ( .A(n18246), .B(n18245), .Z(n18241) );
  IV U26675 ( .A(n18247), .Z(n18245) );
  AND U26676 ( .A(n18248), .B(n18249), .Z(n18214) );
  NAND U26677 ( .A(n18250), .B(n18251), .Z(n18249) );
  NANDN U26678 ( .A(n18252), .B(n18253), .Z(n18251) );
  NANDN U26679 ( .A(n18253), .B(n18252), .Z(n18248) );
  XOR U26680 ( .A(n18224), .B(n18254), .Z(n18216) );
  XNOR U26681 ( .A(n18221), .B(n18223), .Z(n18254) );
  AND U26682 ( .A(n18255), .B(n18256), .Z(n18223) );
  NANDN U26683 ( .A(n18257), .B(n18258), .Z(n18256) );
  OR U26684 ( .A(n18259), .B(n18260), .Z(n18258) );
  IV U26685 ( .A(n18261), .Z(n18260) );
  NANDN U26686 ( .A(n18261), .B(n18259), .Z(n18255) );
  AND U26687 ( .A(n18262), .B(n18263), .Z(n18221) );
  NAND U26688 ( .A(n18264), .B(n18265), .Z(n18263) );
  NANDN U26689 ( .A(n18266), .B(n18267), .Z(n18265) );
  NANDN U26690 ( .A(n18267), .B(n18266), .Z(n18262) );
  IV U26691 ( .A(n18268), .Z(n18267) );
  NAND U26692 ( .A(n18269), .B(n18270), .Z(n18224) );
  NANDN U26693 ( .A(n18271), .B(n18272), .Z(n18270) );
  NANDN U26694 ( .A(n18273), .B(n18274), .Z(n18272) );
  NANDN U26695 ( .A(n18274), .B(n18273), .Z(n18269) );
  IV U26696 ( .A(n18275), .Z(n18273) );
  XOR U26697 ( .A(n18250), .B(n18276), .Z(N63765) );
  XNOR U26698 ( .A(n18253), .B(n18252), .Z(n18276) );
  XNOR U26699 ( .A(n18264), .B(n18277), .Z(n18252) );
  XNOR U26700 ( .A(n18268), .B(n18266), .Z(n18277) );
  XOR U26701 ( .A(n18274), .B(n18278), .Z(n18266) );
  XNOR U26702 ( .A(n18271), .B(n18275), .Z(n18278) );
  AND U26703 ( .A(n18279), .B(n18280), .Z(n18275) );
  NAND U26704 ( .A(n18281), .B(n18282), .Z(n18280) );
  NAND U26705 ( .A(n18283), .B(n18284), .Z(n18279) );
  AND U26706 ( .A(n18285), .B(n18286), .Z(n18271) );
  NAND U26707 ( .A(n18287), .B(n18288), .Z(n18286) );
  NAND U26708 ( .A(n18289), .B(n18290), .Z(n18285) );
  NANDN U26709 ( .A(n18291), .B(n18292), .Z(n18274) );
  ANDN U26710 ( .B(n18293), .A(n18294), .Z(n18268) );
  XNOR U26711 ( .A(n18259), .B(n18295), .Z(n18264) );
  XNOR U26712 ( .A(n18257), .B(n18261), .Z(n18295) );
  AND U26713 ( .A(n18296), .B(n18297), .Z(n18261) );
  NAND U26714 ( .A(n18298), .B(n18299), .Z(n18297) );
  NAND U26715 ( .A(n18300), .B(n18301), .Z(n18296) );
  AND U26716 ( .A(n18302), .B(n18303), .Z(n18257) );
  NAND U26717 ( .A(n18304), .B(n18305), .Z(n18303) );
  NAND U26718 ( .A(n18306), .B(n18307), .Z(n18302) );
  AND U26719 ( .A(n18308), .B(n18309), .Z(n18259) );
  NAND U26720 ( .A(n18310), .B(n18311), .Z(n18253) );
  XNOR U26721 ( .A(n18236), .B(n18312), .Z(n18250) );
  XNOR U26722 ( .A(n18240), .B(n18238), .Z(n18312) );
  XOR U26723 ( .A(n18246), .B(n18313), .Z(n18238) );
  XNOR U26724 ( .A(n18243), .B(n18247), .Z(n18313) );
  AND U26725 ( .A(n18314), .B(n18315), .Z(n18247) );
  NAND U26726 ( .A(n18316), .B(n18317), .Z(n18315) );
  NAND U26727 ( .A(n18318), .B(n18319), .Z(n18314) );
  AND U26728 ( .A(n18320), .B(n18321), .Z(n18243) );
  NAND U26729 ( .A(n18322), .B(n18323), .Z(n18321) );
  NAND U26730 ( .A(n18324), .B(n18325), .Z(n18320) );
  NANDN U26731 ( .A(n18326), .B(n18327), .Z(n18246) );
  ANDN U26732 ( .B(n18328), .A(n18329), .Z(n18240) );
  XNOR U26733 ( .A(n18231), .B(n18330), .Z(n18236) );
  XNOR U26734 ( .A(n18229), .B(n18233), .Z(n18330) );
  AND U26735 ( .A(n18331), .B(n18332), .Z(n18233) );
  NAND U26736 ( .A(n18333), .B(n18334), .Z(n18332) );
  NAND U26737 ( .A(n18335), .B(n18336), .Z(n18331) );
  AND U26738 ( .A(n18337), .B(n18338), .Z(n18229) );
  NAND U26739 ( .A(n18339), .B(n18340), .Z(n18338) );
  NAND U26740 ( .A(n18341), .B(n18342), .Z(n18337) );
  AND U26741 ( .A(n18343), .B(n18344), .Z(n18231) );
  XOR U26742 ( .A(n18311), .B(n18310), .Z(N63764) );
  XNOR U26743 ( .A(n18328), .B(n18329), .Z(n18310) );
  XNOR U26744 ( .A(n18343), .B(n18344), .Z(n18329) );
  XOR U26745 ( .A(n18340), .B(n18339), .Z(n18344) );
  XOR U26746 ( .A(y[5868]), .B(x[5868]), .Z(n18339) );
  XOR U26747 ( .A(n18342), .B(n18341), .Z(n18340) );
  XOR U26748 ( .A(y[5870]), .B(x[5870]), .Z(n18341) );
  XOR U26749 ( .A(y[5869]), .B(x[5869]), .Z(n18342) );
  XOR U26750 ( .A(n18334), .B(n18333), .Z(n18343) );
  XOR U26751 ( .A(n18336), .B(n18335), .Z(n18333) );
  XOR U26752 ( .A(y[5867]), .B(x[5867]), .Z(n18335) );
  XOR U26753 ( .A(y[5866]), .B(x[5866]), .Z(n18336) );
  XOR U26754 ( .A(y[5865]), .B(x[5865]), .Z(n18334) );
  XNOR U26755 ( .A(n18327), .B(n18326), .Z(n18328) );
  XNOR U26756 ( .A(n18323), .B(n18322), .Z(n18326) );
  XOR U26757 ( .A(n18325), .B(n18324), .Z(n18322) );
  XOR U26758 ( .A(y[5864]), .B(x[5864]), .Z(n18324) );
  XOR U26759 ( .A(y[5863]), .B(x[5863]), .Z(n18325) );
  XOR U26760 ( .A(y[5862]), .B(x[5862]), .Z(n18323) );
  XOR U26761 ( .A(n18317), .B(n18316), .Z(n18327) );
  XOR U26762 ( .A(n18319), .B(n18318), .Z(n18316) );
  XOR U26763 ( .A(y[5861]), .B(x[5861]), .Z(n18318) );
  XOR U26764 ( .A(y[5860]), .B(x[5860]), .Z(n18319) );
  XOR U26765 ( .A(y[5859]), .B(x[5859]), .Z(n18317) );
  XNOR U26766 ( .A(n18293), .B(n18294), .Z(n18311) );
  XNOR U26767 ( .A(n18308), .B(n18309), .Z(n18294) );
  XOR U26768 ( .A(n18305), .B(n18304), .Z(n18309) );
  XOR U26769 ( .A(y[5856]), .B(x[5856]), .Z(n18304) );
  XOR U26770 ( .A(n18307), .B(n18306), .Z(n18305) );
  XOR U26771 ( .A(y[5858]), .B(x[5858]), .Z(n18306) );
  XOR U26772 ( .A(y[5857]), .B(x[5857]), .Z(n18307) );
  XOR U26773 ( .A(n18299), .B(n18298), .Z(n18308) );
  XOR U26774 ( .A(n18301), .B(n18300), .Z(n18298) );
  XOR U26775 ( .A(y[5855]), .B(x[5855]), .Z(n18300) );
  XOR U26776 ( .A(y[5854]), .B(x[5854]), .Z(n18301) );
  XOR U26777 ( .A(y[5853]), .B(x[5853]), .Z(n18299) );
  XNOR U26778 ( .A(n18292), .B(n18291), .Z(n18293) );
  XNOR U26779 ( .A(n18288), .B(n18287), .Z(n18291) );
  XOR U26780 ( .A(n18290), .B(n18289), .Z(n18287) );
  XOR U26781 ( .A(y[5852]), .B(x[5852]), .Z(n18289) );
  XOR U26782 ( .A(y[5851]), .B(x[5851]), .Z(n18290) );
  XOR U26783 ( .A(y[5850]), .B(x[5850]), .Z(n18288) );
  XOR U26784 ( .A(n18282), .B(n18281), .Z(n18292) );
  XOR U26785 ( .A(n18284), .B(n18283), .Z(n18281) );
  XOR U26786 ( .A(y[5849]), .B(x[5849]), .Z(n18283) );
  XOR U26787 ( .A(y[5848]), .B(x[5848]), .Z(n18284) );
  XOR U26788 ( .A(y[5847]), .B(x[5847]), .Z(n18282) );
  NAND U26789 ( .A(n18345), .B(n18346), .Z(N63755) );
  NAND U26790 ( .A(n18347), .B(n18348), .Z(n18346) );
  NANDN U26791 ( .A(n18349), .B(n18350), .Z(n18348) );
  NANDN U26792 ( .A(n18350), .B(n18349), .Z(n18345) );
  XOR U26793 ( .A(n18349), .B(n18351), .Z(N63754) );
  XNOR U26794 ( .A(n18347), .B(n18350), .Z(n18351) );
  NAND U26795 ( .A(n18352), .B(n18353), .Z(n18350) );
  NAND U26796 ( .A(n18354), .B(n18355), .Z(n18353) );
  NANDN U26797 ( .A(n18356), .B(n18357), .Z(n18355) );
  NANDN U26798 ( .A(n18357), .B(n18356), .Z(n18352) );
  AND U26799 ( .A(n18358), .B(n18359), .Z(n18347) );
  NAND U26800 ( .A(n18360), .B(n18361), .Z(n18359) );
  NANDN U26801 ( .A(n18362), .B(n18363), .Z(n18361) );
  NANDN U26802 ( .A(n18363), .B(n18362), .Z(n18358) );
  IV U26803 ( .A(n18364), .Z(n18363) );
  AND U26804 ( .A(n18365), .B(n18366), .Z(n18349) );
  NAND U26805 ( .A(n18367), .B(n18368), .Z(n18366) );
  NANDN U26806 ( .A(n18369), .B(n18370), .Z(n18368) );
  NANDN U26807 ( .A(n18370), .B(n18369), .Z(n18365) );
  XOR U26808 ( .A(n18362), .B(n18371), .Z(N63753) );
  XNOR U26809 ( .A(n18360), .B(n18364), .Z(n18371) );
  XOR U26810 ( .A(n18357), .B(n18372), .Z(n18364) );
  XNOR U26811 ( .A(n18354), .B(n18356), .Z(n18372) );
  AND U26812 ( .A(n18373), .B(n18374), .Z(n18356) );
  NANDN U26813 ( .A(n18375), .B(n18376), .Z(n18374) );
  OR U26814 ( .A(n18377), .B(n18378), .Z(n18376) );
  IV U26815 ( .A(n18379), .Z(n18378) );
  NANDN U26816 ( .A(n18379), .B(n18377), .Z(n18373) );
  AND U26817 ( .A(n18380), .B(n18381), .Z(n18354) );
  NAND U26818 ( .A(n18382), .B(n18383), .Z(n18381) );
  NANDN U26819 ( .A(n18384), .B(n18385), .Z(n18383) );
  NANDN U26820 ( .A(n18385), .B(n18384), .Z(n18380) );
  IV U26821 ( .A(n18386), .Z(n18385) );
  NAND U26822 ( .A(n18387), .B(n18388), .Z(n18357) );
  NANDN U26823 ( .A(n18389), .B(n18390), .Z(n18388) );
  NANDN U26824 ( .A(n18391), .B(n18392), .Z(n18390) );
  NANDN U26825 ( .A(n18392), .B(n18391), .Z(n18387) );
  IV U26826 ( .A(n18393), .Z(n18391) );
  AND U26827 ( .A(n18394), .B(n18395), .Z(n18360) );
  NAND U26828 ( .A(n18396), .B(n18397), .Z(n18395) );
  NANDN U26829 ( .A(n18398), .B(n18399), .Z(n18397) );
  NANDN U26830 ( .A(n18399), .B(n18398), .Z(n18394) );
  XOR U26831 ( .A(n18370), .B(n18400), .Z(n18362) );
  XNOR U26832 ( .A(n18367), .B(n18369), .Z(n18400) );
  AND U26833 ( .A(n18401), .B(n18402), .Z(n18369) );
  NANDN U26834 ( .A(n18403), .B(n18404), .Z(n18402) );
  OR U26835 ( .A(n18405), .B(n18406), .Z(n18404) );
  IV U26836 ( .A(n18407), .Z(n18406) );
  NANDN U26837 ( .A(n18407), .B(n18405), .Z(n18401) );
  AND U26838 ( .A(n18408), .B(n18409), .Z(n18367) );
  NAND U26839 ( .A(n18410), .B(n18411), .Z(n18409) );
  NANDN U26840 ( .A(n18412), .B(n18413), .Z(n18411) );
  NANDN U26841 ( .A(n18413), .B(n18412), .Z(n18408) );
  IV U26842 ( .A(n18414), .Z(n18413) );
  NAND U26843 ( .A(n18415), .B(n18416), .Z(n18370) );
  NANDN U26844 ( .A(n18417), .B(n18418), .Z(n18416) );
  NANDN U26845 ( .A(n18419), .B(n18420), .Z(n18418) );
  NANDN U26846 ( .A(n18420), .B(n18419), .Z(n18415) );
  IV U26847 ( .A(n18421), .Z(n18419) );
  XOR U26848 ( .A(n18396), .B(n18422), .Z(N63752) );
  XNOR U26849 ( .A(n18399), .B(n18398), .Z(n18422) );
  XNOR U26850 ( .A(n18410), .B(n18423), .Z(n18398) );
  XNOR U26851 ( .A(n18414), .B(n18412), .Z(n18423) );
  XOR U26852 ( .A(n18420), .B(n18424), .Z(n18412) );
  XNOR U26853 ( .A(n18417), .B(n18421), .Z(n18424) );
  AND U26854 ( .A(n18425), .B(n18426), .Z(n18421) );
  NAND U26855 ( .A(n18427), .B(n18428), .Z(n18426) );
  NAND U26856 ( .A(n18429), .B(n18430), .Z(n18425) );
  AND U26857 ( .A(n18431), .B(n18432), .Z(n18417) );
  NAND U26858 ( .A(n18433), .B(n18434), .Z(n18432) );
  NAND U26859 ( .A(n18435), .B(n18436), .Z(n18431) );
  NANDN U26860 ( .A(n18437), .B(n18438), .Z(n18420) );
  ANDN U26861 ( .B(n18439), .A(n18440), .Z(n18414) );
  XNOR U26862 ( .A(n18405), .B(n18441), .Z(n18410) );
  XNOR U26863 ( .A(n18403), .B(n18407), .Z(n18441) );
  AND U26864 ( .A(n18442), .B(n18443), .Z(n18407) );
  NAND U26865 ( .A(n18444), .B(n18445), .Z(n18443) );
  NAND U26866 ( .A(n18446), .B(n18447), .Z(n18442) );
  AND U26867 ( .A(n18448), .B(n18449), .Z(n18403) );
  NAND U26868 ( .A(n18450), .B(n18451), .Z(n18449) );
  NAND U26869 ( .A(n18452), .B(n18453), .Z(n18448) );
  AND U26870 ( .A(n18454), .B(n18455), .Z(n18405) );
  NAND U26871 ( .A(n18456), .B(n18457), .Z(n18399) );
  XNOR U26872 ( .A(n18382), .B(n18458), .Z(n18396) );
  XNOR U26873 ( .A(n18386), .B(n18384), .Z(n18458) );
  XOR U26874 ( .A(n18392), .B(n18459), .Z(n18384) );
  XNOR U26875 ( .A(n18389), .B(n18393), .Z(n18459) );
  AND U26876 ( .A(n18460), .B(n18461), .Z(n18393) );
  NAND U26877 ( .A(n18462), .B(n18463), .Z(n18461) );
  NAND U26878 ( .A(n18464), .B(n18465), .Z(n18460) );
  AND U26879 ( .A(n18466), .B(n18467), .Z(n18389) );
  NAND U26880 ( .A(n18468), .B(n18469), .Z(n18467) );
  NAND U26881 ( .A(n18470), .B(n18471), .Z(n18466) );
  NANDN U26882 ( .A(n18472), .B(n18473), .Z(n18392) );
  ANDN U26883 ( .B(n18474), .A(n18475), .Z(n18386) );
  XNOR U26884 ( .A(n18377), .B(n18476), .Z(n18382) );
  XNOR U26885 ( .A(n18375), .B(n18379), .Z(n18476) );
  AND U26886 ( .A(n18477), .B(n18478), .Z(n18379) );
  NAND U26887 ( .A(n18479), .B(n18480), .Z(n18478) );
  NAND U26888 ( .A(n18481), .B(n18482), .Z(n18477) );
  AND U26889 ( .A(n18483), .B(n18484), .Z(n18375) );
  NAND U26890 ( .A(n18485), .B(n18486), .Z(n18484) );
  NAND U26891 ( .A(n18487), .B(n18488), .Z(n18483) );
  AND U26892 ( .A(n18489), .B(n18490), .Z(n18377) );
  XOR U26893 ( .A(n18457), .B(n18456), .Z(N63751) );
  XNOR U26894 ( .A(n18474), .B(n18475), .Z(n18456) );
  XNOR U26895 ( .A(n18489), .B(n18490), .Z(n18475) );
  XOR U26896 ( .A(n18486), .B(n18485), .Z(n18490) );
  XOR U26897 ( .A(y[5844]), .B(x[5844]), .Z(n18485) );
  XOR U26898 ( .A(n18488), .B(n18487), .Z(n18486) );
  XOR U26899 ( .A(y[5846]), .B(x[5846]), .Z(n18487) );
  XOR U26900 ( .A(y[5845]), .B(x[5845]), .Z(n18488) );
  XOR U26901 ( .A(n18480), .B(n18479), .Z(n18489) );
  XOR U26902 ( .A(n18482), .B(n18481), .Z(n18479) );
  XOR U26903 ( .A(y[5843]), .B(x[5843]), .Z(n18481) );
  XOR U26904 ( .A(y[5842]), .B(x[5842]), .Z(n18482) );
  XOR U26905 ( .A(y[5841]), .B(x[5841]), .Z(n18480) );
  XNOR U26906 ( .A(n18473), .B(n18472), .Z(n18474) );
  XNOR U26907 ( .A(n18469), .B(n18468), .Z(n18472) );
  XOR U26908 ( .A(n18471), .B(n18470), .Z(n18468) );
  XOR U26909 ( .A(y[5840]), .B(x[5840]), .Z(n18470) );
  XOR U26910 ( .A(y[5839]), .B(x[5839]), .Z(n18471) );
  XOR U26911 ( .A(y[5838]), .B(x[5838]), .Z(n18469) );
  XOR U26912 ( .A(n18463), .B(n18462), .Z(n18473) );
  XOR U26913 ( .A(n18465), .B(n18464), .Z(n18462) );
  XOR U26914 ( .A(y[5837]), .B(x[5837]), .Z(n18464) );
  XOR U26915 ( .A(y[5836]), .B(x[5836]), .Z(n18465) );
  XOR U26916 ( .A(y[5835]), .B(x[5835]), .Z(n18463) );
  XNOR U26917 ( .A(n18439), .B(n18440), .Z(n18457) );
  XNOR U26918 ( .A(n18454), .B(n18455), .Z(n18440) );
  XOR U26919 ( .A(n18451), .B(n18450), .Z(n18455) );
  XOR U26920 ( .A(y[5832]), .B(x[5832]), .Z(n18450) );
  XOR U26921 ( .A(n18453), .B(n18452), .Z(n18451) );
  XOR U26922 ( .A(y[5834]), .B(x[5834]), .Z(n18452) );
  XOR U26923 ( .A(y[5833]), .B(x[5833]), .Z(n18453) );
  XOR U26924 ( .A(n18445), .B(n18444), .Z(n18454) );
  XOR U26925 ( .A(n18447), .B(n18446), .Z(n18444) );
  XOR U26926 ( .A(y[5831]), .B(x[5831]), .Z(n18446) );
  XOR U26927 ( .A(y[5830]), .B(x[5830]), .Z(n18447) );
  XOR U26928 ( .A(y[5829]), .B(x[5829]), .Z(n18445) );
  XNOR U26929 ( .A(n18438), .B(n18437), .Z(n18439) );
  XNOR U26930 ( .A(n18434), .B(n18433), .Z(n18437) );
  XOR U26931 ( .A(n18436), .B(n18435), .Z(n18433) );
  XOR U26932 ( .A(y[5828]), .B(x[5828]), .Z(n18435) );
  XOR U26933 ( .A(y[5827]), .B(x[5827]), .Z(n18436) );
  XOR U26934 ( .A(y[5826]), .B(x[5826]), .Z(n18434) );
  XOR U26935 ( .A(n18428), .B(n18427), .Z(n18438) );
  XOR U26936 ( .A(n18430), .B(n18429), .Z(n18427) );
  XOR U26937 ( .A(y[5825]), .B(x[5825]), .Z(n18429) );
  XOR U26938 ( .A(y[5824]), .B(x[5824]), .Z(n18430) );
  XOR U26939 ( .A(y[5823]), .B(x[5823]), .Z(n18428) );
  NAND U26940 ( .A(n18491), .B(n18492), .Z(N63742) );
  NAND U26941 ( .A(n18493), .B(n18494), .Z(n18492) );
  NANDN U26942 ( .A(n18495), .B(n18496), .Z(n18494) );
  NANDN U26943 ( .A(n18496), .B(n18495), .Z(n18491) );
  XOR U26944 ( .A(n18495), .B(n18497), .Z(N63741) );
  XNOR U26945 ( .A(n18493), .B(n18496), .Z(n18497) );
  NAND U26946 ( .A(n18498), .B(n18499), .Z(n18496) );
  NAND U26947 ( .A(n18500), .B(n18501), .Z(n18499) );
  NANDN U26948 ( .A(n18502), .B(n18503), .Z(n18501) );
  NANDN U26949 ( .A(n18503), .B(n18502), .Z(n18498) );
  AND U26950 ( .A(n18504), .B(n18505), .Z(n18493) );
  NAND U26951 ( .A(n18506), .B(n18507), .Z(n18505) );
  NANDN U26952 ( .A(n18508), .B(n18509), .Z(n18507) );
  NANDN U26953 ( .A(n18509), .B(n18508), .Z(n18504) );
  IV U26954 ( .A(n18510), .Z(n18509) );
  AND U26955 ( .A(n18511), .B(n18512), .Z(n18495) );
  NAND U26956 ( .A(n18513), .B(n18514), .Z(n18512) );
  NANDN U26957 ( .A(n18515), .B(n18516), .Z(n18514) );
  NANDN U26958 ( .A(n18516), .B(n18515), .Z(n18511) );
  XOR U26959 ( .A(n18508), .B(n18517), .Z(N63740) );
  XNOR U26960 ( .A(n18506), .B(n18510), .Z(n18517) );
  XOR U26961 ( .A(n18503), .B(n18518), .Z(n18510) );
  XNOR U26962 ( .A(n18500), .B(n18502), .Z(n18518) );
  AND U26963 ( .A(n18519), .B(n18520), .Z(n18502) );
  NANDN U26964 ( .A(n18521), .B(n18522), .Z(n18520) );
  OR U26965 ( .A(n18523), .B(n18524), .Z(n18522) );
  IV U26966 ( .A(n18525), .Z(n18524) );
  NANDN U26967 ( .A(n18525), .B(n18523), .Z(n18519) );
  AND U26968 ( .A(n18526), .B(n18527), .Z(n18500) );
  NAND U26969 ( .A(n18528), .B(n18529), .Z(n18527) );
  NANDN U26970 ( .A(n18530), .B(n18531), .Z(n18529) );
  NANDN U26971 ( .A(n18531), .B(n18530), .Z(n18526) );
  IV U26972 ( .A(n18532), .Z(n18531) );
  NAND U26973 ( .A(n18533), .B(n18534), .Z(n18503) );
  NANDN U26974 ( .A(n18535), .B(n18536), .Z(n18534) );
  NANDN U26975 ( .A(n18537), .B(n18538), .Z(n18536) );
  NANDN U26976 ( .A(n18538), .B(n18537), .Z(n18533) );
  IV U26977 ( .A(n18539), .Z(n18537) );
  AND U26978 ( .A(n18540), .B(n18541), .Z(n18506) );
  NAND U26979 ( .A(n18542), .B(n18543), .Z(n18541) );
  NANDN U26980 ( .A(n18544), .B(n18545), .Z(n18543) );
  NANDN U26981 ( .A(n18545), .B(n18544), .Z(n18540) );
  XOR U26982 ( .A(n18516), .B(n18546), .Z(n18508) );
  XNOR U26983 ( .A(n18513), .B(n18515), .Z(n18546) );
  AND U26984 ( .A(n18547), .B(n18548), .Z(n18515) );
  NANDN U26985 ( .A(n18549), .B(n18550), .Z(n18548) );
  OR U26986 ( .A(n18551), .B(n18552), .Z(n18550) );
  IV U26987 ( .A(n18553), .Z(n18552) );
  NANDN U26988 ( .A(n18553), .B(n18551), .Z(n18547) );
  AND U26989 ( .A(n18554), .B(n18555), .Z(n18513) );
  NAND U26990 ( .A(n18556), .B(n18557), .Z(n18555) );
  NANDN U26991 ( .A(n18558), .B(n18559), .Z(n18557) );
  NANDN U26992 ( .A(n18559), .B(n18558), .Z(n18554) );
  IV U26993 ( .A(n18560), .Z(n18559) );
  NAND U26994 ( .A(n18561), .B(n18562), .Z(n18516) );
  NANDN U26995 ( .A(n18563), .B(n18564), .Z(n18562) );
  NANDN U26996 ( .A(n18565), .B(n18566), .Z(n18564) );
  NANDN U26997 ( .A(n18566), .B(n18565), .Z(n18561) );
  IV U26998 ( .A(n18567), .Z(n18565) );
  XOR U26999 ( .A(n18542), .B(n18568), .Z(N63739) );
  XNOR U27000 ( .A(n18545), .B(n18544), .Z(n18568) );
  XNOR U27001 ( .A(n18556), .B(n18569), .Z(n18544) );
  XNOR U27002 ( .A(n18560), .B(n18558), .Z(n18569) );
  XOR U27003 ( .A(n18566), .B(n18570), .Z(n18558) );
  XNOR U27004 ( .A(n18563), .B(n18567), .Z(n18570) );
  AND U27005 ( .A(n18571), .B(n18572), .Z(n18567) );
  NAND U27006 ( .A(n18573), .B(n18574), .Z(n18572) );
  NAND U27007 ( .A(n18575), .B(n18576), .Z(n18571) );
  AND U27008 ( .A(n18577), .B(n18578), .Z(n18563) );
  NAND U27009 ( .A(n18579), .B(n18580), .Z(n18578) );
  NAND U27010 ( .A(n18581), .B(n18582), .Z(n18577) );
  NANDN U27011 ( .A(n18583), .B(n18584), .Z(n18566) );
  ANDN U27012 ( .B(n18585), .A(n18586), .Z(n18560) );
  XNOR U27013 ( .A(n18551), .B(n18587), .Z(n18556) );
  XNOR U27014 ( .A(n18549), .B(n18553), .Z(n18587) );
  AND U27015 ( .A(n18588), .B(n18589), .Z(n18553) );
  NAND U27016 ( .A(n18590), .B(n18591), .Z(n18589) );
  NAND U27017 ( .A(n18592), .B(n18593), .Z(n18588) );
  AND U27018 ( .A(n18594), .B(n18595), .Z(n18549) );
  NAND U27019 ( .A(n18596), .B(n18597), .Z(n18595) );
  NAND U27020 ( .A(n18598), .B(n18599), .Z(n18594) );
  AND U27021 ( .A(n18600), .B(n18601), .Z(n18551) );
  NAND U27022 ( .A(n18602), .B(n18603), .Z(n18545) );
  XNOR U27023 ( .A(n18528), .B(n18604), .Z(n18542) );
  XNOR U27024 ( .A(n18532), .B(n18530), .Z(n18604) );
  XOR U27025 ( .A(n18538), .B(n18605), .Z(n18530) );
  XNOR U27026 ( .A(n18535), .B(n18539), .Z(n18605) );
  AND U27027 ( .A(n18606), .B(n18607), .Z(n18539) );
  NAND U27028 ( .A(n18608), .B(n18609), .Z(n18607) );
  NAND U27029 ( .A(n18610), .B(n18611), .Z(n18606) );
  AND U27030 ( .A(n18612), .B(n18613), .Z(n18535) );
  NAND U27031 ( .A(n18614), .B(n18615), .Z(n18613) );
  NAND U27032 ( .A(n18616), .B(n18617), .Z(n18612) );
  NANDN U27033 ( .A(n18618), .B(n18619), .Z(n18538) );
  ANDN U27034 ( .B(n18620), .A(n18621), .Z(n18532) );
  XNOR U27035 ( .A(n18523), .B(n18622), .Z(n18528) );
  XNOR U27036 ( .A(n18521), .B(n18525), .Z(n18622) );
  AND U27037 ( .A(n18623), .B(n18624), .Z(n18525) );
  NAND U27038 ( .A(n18625), .B(n18626), .Z(n18624) );
  NAND U27039 ( .A(n18627), .B(n18628), .Z(n18623) );
  AND U27040 ( .A(n18629), .B(n18630), .Z(n18521) );
  NAND U27041 ( .A(n18631), .B(n18632), .Z(n18630) );
  NAND U27042 ( .A(n18633), .B(n18634), .Z(n18629) );
  AND U27043 ( .A(n18635), .B(n18636), .Z(n18523) );
  XOR U27044 ( .A(n18603), .B(n18602), .Z(N63738) );
  XNOR U27045 ( .A(n18620), .B(n18621), .Z(n18602) );
  XNOR U27046 ( .A(n18635), .B(n18636), .Z(n18621) );
  XOR U27047 ( .A(n18632), .B(n18631), .Z(n18636) );
  XOR U27048 ( .A(y[5820]), .B(x[5820]), .Z(n18631) );
  XOR U27049 ( .A(n18634), .B(n18633), .Z(n18632) );
  XOR U27050 ( .A(y[5822]), .B(x[5822]), .Z(n18633) );
  XOR U27051 ( .A(y[5821]), .B(x[5821]), .Z(n18634) );
  XOR U27052 ( .A(n18626), .B(n18625), .Z(n18635) );
  XOR U27053 ( .A(n18628), .B(n18627), .Z(n18625) );
  XOR U27054 ( .A(y[5819]), .B(x[5819]), .Z(n18627) );
  XOR U27055 ( .A(y[5818]), .B(x[5818]), .Z(n18628) );
  XOR U27056 ( .A(y[5817]), .B(x[5817]), .Z(n18626) );
  XNOR U27057 ( .A(n18619), .B(n18618), .Z(n18620) );
  XNOR U27058 ( .A(n18615), .B(n18614), .Z(n18618) );
  XOR U27059 ( .A(n18617), .B(n18616), .Z(n18614) );
  XOR U27060 ( .A(y[5816]), .B(x[5816]), .Z(n18616) );
  XOR U27061 ( .A(y[5815]), .B(x[5815]), .Z(n18617) );
  XOR U27062 ( .A(y[5814]), .B(x[5814]), .Z(n18615) );
  XOR U27063 ( .A(n18609), .B(n18608), .Z(n18619) );
  XOR U27064 ( .A(n18611), .B(n18610), .Z(n18608) );
  XOR U27065 ( .A(y[5813]), .B(x[5813]), .Z(n18610) );
  XOR U27066 ( .A(y[5812]), .B(x[5812]), .Z(n18611) );
  XOR U27067 ( .A(y[5811]), .B(x[5811]), .Z(n18609) );
  XNOR U27068 ( .A(n18585), .B(n18586), .Z(n18603) );
  XNOR U27069 ( .A(n18600), .B(n18601), .Z(n18586) );
  XOR U27070 ( .A(n18597), .B(n18596), .Z(n18601) );
  XOR U27071 ( .A(y[5808]), .B(x[5808]), .Z(n18596) );
  XOR U27072 ( .A(n18599), .B(n18598), .Z(n18597) );
  XOR U27073 ( .A(y[5810]), .B(x[5810]), .Z(n18598) );
  XOR U27074 ( .A(y[5809]), .B(x[5809]), .Z(n18599) );
  XOR U27075 ( .A(n18591), .B(n18590), .Z(n18600) );
  XOR U27076 ( .A(n18593), .B(n18592), .Z(n18590) );
  XOR U27077 ( .A(y[5807]), .B(x[5807]), .Z(n18592) );
  XOR U27078 ( .A(y[5806]), .B(x[5806]), .Z(n18593) );
  XOR U27079 ( .A(y[5805]), .B(x[5805]), .Z(n18591) );
  XNOR U27080 ( .A(n18584), .B(n18583), .Z(n18585) );
  XNOR U27081 ( .A(n18580), .B(n18579), .Z(n18583) );
  XOR U27082 ( .A(n18582), .B(n18581), .Z(n18579) );
  XOR U27083 ( .A(y[5804]), .B(x[5804]), .Z(n18581) );
  XOR U27084 ( .A(y[5803]), .B(x[5803]), .Z(n18582) );
  XOR U27085 ( .A(y[5802]), .B(x[5802]), .Z(n18580) );
  XOR U27086 ( .A(n18574), .B(n18573), .Z(n18584) );
  XOR U27087 ( .A(n18576), .B(n18575), .Z(n18573) );
  XOR U27088 ( .A(y[5801]), .B(x[5801]), .Z(n18575) );
  XOR U27089 ( .A(y[5800]), .B(x[5800]), .Z(n18576) );
  XOR U27090 ( .A(y[5799]), .B(x[5799]), .Z(n18574) );
  NAND U27091 ( .A(n18637), .B(n18638), .Z(N63729) );
  NAND U27092 ( .A(n18639), .B(n18640), .Z(n18638) );
  NANDN U27093 ( .A(n18641), .B(n18642), .Z(n18640) );
  NANDN U27094 ( .A(n18642), .B(n18641), .Z(n18637) );
  XOR U27095 ( .A(n18641), .B(n18643), .Z(N63728) );
  XNOR U27096 ( .A(n18639), .B(n18642), .Z(n18643) );
  NAND U27097 ( .A(n18644), .B(n18645), .Z(n18642) );
  NAND U27098 ( .A(n18646), .B(n18647), .Z(n18645) );
  NANDN U27099 ( .A(n18648), .B(n18649), .Z(n18647) );
  NANDN U27100 ( .A(n18649), .B(n18648), .Z(n18644) );
  AND U27101 ( .A(n18650), .B(n18651), .Z(n18639) );
  NAND U27102 ( .A(n18652), .B(n18653), .Z(n18651) );
  NANDN U27103 ( .A(n18654), .B(n18655), .Z(n18653) );
  NANDN U27104 ( .A(n18655), .B(n18654), .Z(n18650) );
  IV U27105 ( .A(n18656), .Z(n18655) );
  AND U27106 ( .A(n18657), .B(n18658), .Z(n18641) );
  NAND U27107 ( .A(n18659), .B(n18660), .Z(n18658) );
  NANDN U27108 ( .A(n18661), .B(n18662), .Z(n18660) );
  NANDN U27109 ( .A(n18662), .B(n18661), .Z(n18657) );
  XOR U27110 ( .A(n18654), .B(n18663), .Z(N63727) );
  XNOR U27111 ( .A(n18652), .B(n18656), .Z(n18663) );
  XOR U27112 ( .A(n18649), .B(n18664), .Z(n18656) );
  XNOR U27113 ( .A(n18646), .B(n18648), .Z(n18664) );
  AND U27114 ( .A(n18665), .B(n18666), .Z(n18648) );
  NANDN U27115 ( .A(n18667), .B(n18668), .Z(n18666) );
  OR U27116 ( .A(n18669), .B(n18670), .Z(n18668) );
  IV U27117 ( .A(n18671), .Z(n18670) );
  NANDN U27118 ( .A(n18671), .B(n18669), .Z(n18665) );
  AND U27119 ( .A(n18672), .B(n18673), .Z(n18646) );
  NAND U27120 ( .A(n18674), .B(n18675), .Z(n18673) );
  NANDN U27121 ( .A(n18676), .B(n18677), .Z(n18675) );
  NANDN U27122 ( .A(n18677), .B(n18676), .Z(n18672) );
  IV U27123 ( .A(n18678), .Z(n18677) );
  NAND U27124 ( .A(n18679), .B(n18680), .Z(n18649) );
  NANDN U27125 ( .A(n18681), .B(n18682), .Z(n18680) );
  NANDN U27126 ( .A(n18683), .B(n18684), .Z(n18682) );
  NANDN U27127 ( .A(n18684), .B(n18683), .Z(n18679) );
  IV U27128 ( .A(n18685), .Z(n18683) );
  AND U27129 ( .A(n18686), .B(n18687), .Z(n18652) );
  NAND U27130 ( .A(n18688), .B(n18689), .Z(n18687) );
  NANDN U27131 ( .A(n18690), .B(n18691), .Z(n18689) );
  NANDN U27132 ( .A(n18691), .B(n18690), .Z(n18686) );
  XOR U27133 ( .A(n18662), .B(n18692), .Z(n18654) );
  XNOR U27134 ( .A(n18659), .B(n18661), .Z(n18692) );
  AND U27135 ( .A(n18693), .B(n18694), .Z(n18661) );
  NANDN U27136 ( .A(n18695), .B(n18696), .Z(n18694) );
  OR U27137 ( .A(n18697), .B(n18698), .Z(n18696) );
  IV U27138 ( .A(n18699), .Z(n18698) );
  NANDN U27139 ( .A(n18699), .B(n18697), .Z(n18693) );
  AND U27140 ( .A(n18700), .B(n18701), .Z(n18659) );
  NAND U27141 ( .A(n18702), .B(n18703), .Z(n18701) );
  NANDN U27142 ( .A(n18704), .B(n18705), .Z(n18703) );
  NANDN U27143 ( .A(n18705), .B(n18704), .Z(n18700) );
  IV U27144 ( .A(n18706), .Z(n18705) );
  NAND U27145 ( .A(n18707), .B(n18708), .Z(n18662) );
  NANDN U27146 ( .A(n18709), .B(n18710), .Z(n18708) );
  NANDN U27147 ( .A(n18711), .B(n18712), .Z(n18710) );
  NANDN U27148 ( .A(n18712), .B(n18711), .Z(n18707) );
  IV U27149 ( .A(n18713), .Z(n18711) );
  XOR U27150 ( .A(n18688), .B(n18714), .Z(N63726) );
  XNOR U27151 ( .A(n18691), .B(n18690), .Z(n18714) );
  XNOR U27152 ( .A(n18702), .B(n18715), .Z(n18690) );
  XNOR U27153 ( .A(n18706), .B(n18704), .Z(n18715) );
  XOR U27154 ( .A(n18712), .B(n18716), .Z(n18704) );
  XNOR U27155 ( .A(n18709), .B(n18713), .Z(n18716) );
  AND U27156 ( .A(n18717), .B(n18718), .Z(n18713) );
  NAND U27157 ( .A(n18719), .B(n18720), .Z(n18718) );
  NAND U27158 ( .A(n18721), .B(n18722), .Z(n18717) );
  AND U27159 ( .A(n18723), .B(n18724), .Z(n18709) );
  NAND U27160 ( .A(n18725), .B(n18726), .Z(n18724) );
  NAND U27161 ( .A(n18727), .B(n18728), .Z(n18723) );
  NANDN U27162 ( .A(n18729), .B(n18730), .Z(n18712) );
  ANDN U27163 ( .B(n18731), .A(n18732), .Z(n18706) );
  XNOR U27164 ( .A(n18697), .B(n18733), .Z(n18702) );
  XNOR U27165 ( .A(n18695), .B(n18699), .Z(n18733) );
  AND U27166 ( .A(n18734), .B(n18735), .Z(n18699) );
  NAND U27167 ( .A(n18736), .B(n18737), .Z(n18735) );
  NAND U27168 ( .A(n18738), .B(n18739), .Z(n18734) );
  AND U27169 ( .A(n18740), .B(n18741), .Z(n18695) );
  NAND U27170 ( .A(n18742), .B(n18743), .Z(n18741) );
  NAND U27171 ( .A(n18744), .B(n18745), .Z(n18740) );
  AND U27172 ( .A(n18746), .B(n18747), .Z(n18697) );
  NAND U27173 ( .A(n18748), .B(n18749), .Z(n18691) );
  XNOR U27174 ( .A(n18674), .B(n18750), .Z(n18688) );
  XNOR U27175 ( .A(n18678), .B(n18676), .Z(n18750) );
  XOR U27176 ( .A(n18684), .B(n18751), .Z(n18676) );
  XNOR U27177 ( .A(n18681), .B(n18685), .Z(n18751) );
  AND U27178 ( .A(n18752), .B(n18753), .Z(n18685) );
  NAND U27179 ( .A(n18754), .B(n18755), .Z(n18753) );
  NAND U27180 ( .A(n18756), .B(n18757), .Z(n18752) );
  AND U27181 ( .A(n18758), .B(n18759), .Z(n18681) );
  NAND U27182 ( .A(n18760), .B(n18761), .Z(n18759) );
  NAND U27183 ( .A(n18762), .B(n18763), .Z(n18758) );
  NANDN U27184 ( .A(n18764), .B(n18765), .Z(n18684) );
  ANDN U27185 ( .B(n18766), .A(n18767), .Z(n18678) );
  XNOR U27186 ( .A(n18669), .B(n18768), .Z(n18674) );
  XNOR U27187 ( .A(n18667), .B(n18671), .Z(n18768) );
  AND U27188 ( .A(n18769), .B(n18770), .Z(n18671) );
  NAND U27189 ( .A(n18771), .B(n18772), .Z(n18770) );
  NAND U27190 ( .A(n18773), .B(n18774), .Z(n18769) );
  AND U27191 ( .A(n18775), .B(n18776), .Z(n18667) );
  NAND U27192 ( .A(n18777), .B(n18778), .Z(n18776) );
  NAND U27193 ( .A(n18779), .B(n18780), .Z(n18775) );
  AND U27194 ( .A(n18781), .B(n18782), .Z(n18669) );
  XOR U27195 ( .A(n18749), .B(n18748), .Z(N63725) );
  XNOR U27196 ( .A(n18766), .B(n18767), .Z(n18748) );
  XNOR U27197 ( .A(n18781), .B(n18782), .Z(n18767) );
  XOR U27198 ( .A(n18778), .B(n18777), .Z(n18782) );
  XOR U27199 ( .A(y[5796]), .B(x[5796]), .Z(n18777) );
  XOR U27200 ( .A(n18780), .B(n18779), .Z(n18778) );
  XOR U27201 ( .A(y[5798]), .B(x[5798]), .Z(n18779) );
  XOR U27202 ( .A(y[5797]), .B(x[5797]), .Z(n18780) );
  XOR U27203 ( .A(n18772), .B(n18771), .Z(n18781) );
  XOR U27204 ( .A(n18774), .B(n18773), .Z(n18771) );
  XOR U27205 ( .A(y[5795]), .B(x[5795]), .Z(n18773) );
  XOR U27206 ( .A(y[5794]), .B(x[5794]), .Z(n18774) );
  XOR U27207 ( .A(y[5793]), .B(x[5793]), .Z(n18772) );
  XNOR U27208 ( .A(n18765), .B(n18764), .Z(n18766) );
  XNOR U27209 ( .A(n18761), .B(n18760), .Z(n18764) );
  XOR U27210 ( .A(n18763), .B(n18762), .Z(n18760) );
  XOR U27211 ( .A(y[5792]), .B(x[5792]), .Z(n18762) );
  XOR U27212 ( .A(y[5791]), .B(x[5791]), .Z(n18763) );
  XOR U27213 ( .A(y[5790]), .B(x[5790]), .Z(n18761) );
  XOR U27214 ( .A(n18755), .B(n18754), .Z(n18765) );
  XOR U27215 ( .A(n18757), .B(n18756), .Z(n18754) );
  XOR U27216 ( .A(y[5789]), .B(x[5789]), .Z(n18756) );
  XOR U27217 ( .A(y[5788]), .B(x[5788]), .Z(n18757) );
  XOR U27218 ( .A(y[5787]), .B(x[5787]), .Z(n18755) );
  XNOR U27219 ( .A(n18731), .B(n18732), .Z(n18749) );
  XNOR U27220 ( .A(n18746), .B(n18747), .Z(n18732) );
  XOR U27221 ( .A(n18743), .B(n18742), .Z(n18747) );
  XOR U27222 ( .A(y[5784]), .B(x[5784]), .Z(n18742) );
  XOR U27223 ( .A(n18745), .B(n18744), .Z(n18743) );
  XOR U27224 ( .A(y[5786]), .B(x[5786]), .Z(n18744) );
  XOR U27225 ( .A(y[5785]), .B(x[5785]), .Z(n18745) );
  XOR U27226 ( .A(n18737), .B(n18736), .Z(n18746) );
  XOR U27227 ( .A(n18739), .B(n18738), .Z(n18736) );
  XOR U27228 ( .A(y[5783]), .B(x[5783]), .Z(n18738) );
  XOR U27229 ( .A(y[5782]), .B(x[5782]), .Z(n18739) );
  XOR U27230 ( .A(y[5781]), .B(x[5781]), .Z(n18737) );
  XNOR U27231 ( .A(n18730), .B(n18729), .Z(n18731) );
  XNOR U27232 ( .A(n18726), .B(n18725), .Z(n18729) );
  XOR U27233 ( .A(n18728), .B(n18727), .Z(n18725) );
  XOR U27234 ( .A(y[5780]), .B(x[5780]), .Z(n18727) );
  XOR U27235 ( .A(y[5779]), .B(x[5779]), .Z(n18728) );
  XOR U27236 ( .A(y[5778]), .B(x[5778]), .Z(n18726) );
  XOR U27237 ( .A(n18720), .B(n18719), .Z(n18730) );
  XOR U27238 ( .A(n18722), .B(n18721), .Z(n18719) );
  XOR U27239 ( .A(y[5777]), .B(x[5777]), .Z(n18721) );
  XOR U27240 ( .A(y[5776]), .B(x[5776]), .Z(n18722) );
  XOR U27241 ( .A(y[5775]), .B(x[5775]), .Z(n18720) );
  NAND U27242 ( .A(n18783), .B(n18784), .Z(N63716) );
  NAND U27243 ( .A(n18785), .B(n18786), .Z(n18784) );
  NANDN U27244 ( .A(n18787), .B(n18788), .Z(n18786) );
  NANDN U27245 ( .A(n18788), .B(n18787), .Z(n18783) );
  XOR U27246 ( .A(n18787), .B(n18789), .Z(N63715) );
  XNOR U27247 ( .A(n18785), .B(n18788), .Z(n18789) );
  NAND U27248 ( .A(n18790), .B(n18791), .Z(n18788) );
  NAND U27249 ( .A(n18792), .B(n18793), .Z(n18791) );
  NANDN U27250 ( .A(n18794), .B(n18795), .Z(n18793) );
  NANDN U27251 ( .A(n18795), .B(n18794), .Z(n18790) );
  AND U27252 ( .A(n18796), .B(n18797), .Z(n18785) );
  NAND U27253 ( .A(n18798), .B(n18799), .Z(n18797) );
  NANDN U27254 ( .A(n18800), .B(n18801), .Z(n18799) );
  NANDN U27255 ( .A(n18801), .B(n18800), .Z(n18796) );
  IV U27256 ( .A(n18802), .Z(n18801) );
  AND U27257 ( .A(n18803), .B(n18804), .Z(n18787) );
  NAND U27258 ( .A(n18805), .B(n18806), .Z(n18804) );
  NANDN U27259 ( .A(n18807), .B(n18808), .Z(n18806) );
  NANDN U27260 ( .A(n18808), .B(n18807), .Z(n18803) );
  XOR U27261 ( .A(n18800), .B(n18809), .Z(N63714) );
  XNOR U27262 ( .A(n18798), .B(n18802), .Z(n18809) );
  XOR U27263 ( .A(n18795), .B(n18810), .Z(n18802) );
  XNOR U27264 ( .A(n18792), .B(n18794), .Z(n18810) );
  AND U27265 ( .A(n18811), .B(n18812), .Z(n18794) );
  NANDN U27266 ( .A(n18813), .B(n18814), .Z(n18812) );
  OR U27267 ( .A(n18815), .B(n18816), .Z(n18814) );
  IV U27268 ( .A(n18817), .Z(n18816) );
  NANDN U27269 ( .A(n18817), .B(n18815), .Z(n18811) );
  AND U27270 ( .A(n18818), .B(n18819), .Z(n18792) );
  NAND U27271 ( .A(n18820), .B(n18821), .Z(n18819) );
  NANDN U27272 ( .A(n18822), .B(n18823), .Z(n18821) );
  NANDN U27273 ( .A(n18823), .B(n18822), .Z(n18818) );
  IV U27274 ( .A(n18824), .Z(n18823) );
  NAND U27275 ( .A(n18825), .B(n18826), .Z(n18795) );
  NANDN U27276 ( .A(n18827), .B(n18828), .Z(n18826) );
  NANDN U27277 ( .A(n18829), .B(n18830), .Z(n18828) );
  NANDN U27278 ( .A(n18830), .B(n18829), .Z(n18825) );
  IV U27279 ( .A(n18831), .Z(n18829) );
  AND U27280 ( .A(n18832), .B(n18833), .Z(n18798) );
  NAND U27281 ( .A(n18834), .B(n18835), .Z(n18833) );
  NANDN U27282 ( .A(n18836), .B(n18837), .Z(n18835) );
  NANDN U27283 ( .A(n18837), .B(n18836), .Z(n18832) );
  XOR U27284 ( .A(n18808), .B(n18838), .Z(n18800) );
  XNOR U27285 ( .A(n18805), .B(n18807), .Z(n18838) );
  AND U27286 ( .A(n18839), .B(n18840), .Z(n18807) );
  NANDN U27287 ( .A(n18841), .B(n18842), .Z(n18840) );
  OR U27288 ( .A(n18843), .B(n18844), .Z(n18842) );
  IV U27289 ( .A(n18845), .Z(n18844) );
  NANDN U27290 ( .A(n18845), .B(n18843), .Z(n18839) );
  AND U27291 ( .A(n18846), .B(n18847), .Z(n18805) );
  NAND U27292 ( .A(n18848), .B(n18849), .Z(n18847) );
  NANDN U27293 ( .A(n18850), .B(n18851), .Z(n18849) );
  NANDN U27294 ( .A(n18851), .B(n18850), .Z(n18846) );
  IV U27295 ( .A(n18852), .Z(n18851) );
  NAND U27296 ( .A(n18853), .B(n18854), .Z(n18808) );
  NANDN U27297 ( .A(n18855), .B(n18856), .Z(n18854) );
  NANDN U27298 ( .A(n18857), .B(n18858), .Z(n18856) );
  NANDN U27299 ( .A(n18858), .B(n18857), .Z(n18853) );
  IV U27300 ( .A(n18859), .Z(n18857) );
  XOR U27301 ( .A(n18834), .B(n18860), .Z(N63713) );
  XNOR U27302 ( .A(n18837), .B(n18836), .Z(n18860) );
  XNOR U27303 ( .A(n18848), .B(n18861), .Z(n18836) );
  XNOR U27304 ( .A(n18852), .B(n18850), .Z(n18861) );
  XOR U27305 ( .A(n18858), .B(n18862), .Z(n18850) );
  XNOR U27306 ( .A(n18855), .B(n18859), .Z(n18862) );
  AND U27307 ( .A(n18863), .B(n18864), .Z(n18859) );
  NAND U27308 ( .A(n18865), .B(n18866), .Z(n18864) );
  NAND U27309 ( .A(n18867), .B(n18868), .Z(n18863) );
  AND U27310 ( .A(n18869), .B(n18870), .Z(n18855) );
  NAND U27311 ( .A(n18871), .B(n18872), .Z(n18870) );
  NAND U27312 ( .A(n18873), .B(n18874), .Z(n18869) );
  NANDN U27313 ( .A(n18875), .B(n18876), .Z(n18858) );
  ANDN U27314 ( .B(n18877), .A(n18878), .Z(n18852) );
  XNOR U27315 ( .A(n18843), .B(n18879), .Z(n18848) );
  XNOR U27316 ( .A(n18841), .B(n18845), .Z(n18879) );
  AND U27317 ( .A(n18880), .B(n18881), .Z(n18845) );
  NAND U27318 ( .A(n18882), .B(n18883), .Z(n18881) );
  NAND U27319 ( .A(n18884), .B(n18885), .Z(n18880) );
  AND U27320 ( .A(n18886), .B(n18887), .Z(n18841) );
  NAND U27321 ( .A(n18888), .B(n18889), .Z(n18887) );
  NAND U27322 ( .A(n18890), .B(n18891), .Z(n18886) );
  AND U27323 ( .A(n18892), .B(n18893), .Z(n18843) );
  NAND U27324 ( .A(n18894), .B(n18895), .Z(n18837) );
  XNOR U27325 ( .A(n18820), .B(n18896), .Z(n18834) );
  XNOR U27326 ( .A(n18824), .B(n18822), .Z(n18896) );
  XOR U27327 ( .A(n18830), .B(n18897), .Z(n18822) );
  XNOR U27328 ( .A(n18827), .B(n18831), .Z(n18897) );
  AND U27329 ( .A(n18898), .B(n18899), .Z(n18831) );
  NAND U27330 ( .A(n18900), .B(n18901), .Z(n18899) );
  NAND U27331 ( .A(n18902), .B(n18903), .Z(n18898) );
  AND U27332 ( .A(n18904), .B(n18905), .Z(n18827) );
  NAND U27333 ( .A(n18906), .B(n18907), .Z(n18905) );
  NAND U27334 ( .A(n18908), .B(n18909), .Z(n18904) );
  NANDN U27335 ( .A(n18910), .B(n18911), .Z(n18830) );
  ANDN U27336 ( .B(n18912), .A(n18913), .Z(n18824) );
  XNOR U27337 ( .A(n18815), .B(n18914), .Z(n18820) );
  XNOR U27338 ( .A(n18813), .B(n18817), .Z(n18914) );
  AND U27339 ( .A(n18915), .B(n18916), .Z(n18817) );
  NAND U27340 ( .A(n18917), .B(n18918), .Z(n18916) );
  NAND U27341 ( .A(n18919), .B(n18920), .Z(n18915) );
  AND U27342 ( .A(n18921), .B(n18922), .Z(n18813) );
  NAND U27343 ( .A(n18923), .B(n18924), .Z(n18922) );
  NAND U27344 ( .A(n18925), .B(n18926), .Z(n18921) );
  AND U27345 ( .A(n18927), .B(n18928), .Z(n18815) );
  XOR U27346 ( .A(n18895), .B(n18894), .Z(N63712) );
  XNOR U27347 ( .A(n18912), .B(n18913), .Z(n18894) );
  XNOR U27348 ( .A(n18927), .B(n18928), .Z(n18913) );
  XOR U27349 ( .A(n18924), .B(n18923), .Z(n18928) );
  XOR U27350 ( .A(y[5772]), .B(x[5772]), .Z(n18923) );
  XOR U27351 ( .A(n18926), .B(n18925), .Z(n18924) );
  XOR U27352 ( .A(y[5774]), .B(x[5774]), .Z(n18925) );
  XOR U27353 ( .A(y[5773]), .B(x[5773]), .Z(n18926) );
  XOR U27354 ( .A(n18918), .B(n18917), .Z(n18927) );
  XOR U27355 ( .A(n18920), .B(n18919), .Z(n18917) );
  XOR U27356 ( .A(y[5771]), .B(x[5771]), .Z(n18919) );
  XOR U27357 ( .A(y[5770]), .B(x[5770]), .Z(n18920) );
  XOR U27358 ( .A(y[5769]), .B(x[5769]), .Z(n18918) );
  XNOR U27359 ( .A(n18911), .B(n18910), .Z(n18912) );
  XNOR U27360 ( .A(n18907), .B(n18906), .Z(n18910) );
  XOR U27361 ( .A(n18909), .B(n18908), .Z(n18906) );
  XOR U27362 ( .A(y[5768]), .B(x[5768]), .Z(n18908) );
  XOR U27363 ( .A(y[5767]), .B(x[5767]), .Z(n18909) );
  XOR U27364 ( .A(y[5766]), .B(x[5766]), .Z(n18907) );
  XOR U27365 ( .A(n18901), .B(n18900), .Z(n18911) );
  XOR U27366 ( .A(n18903), .B(n18902), .Z(n18900) );
  XOR U27367 ( .A(y[5765]), .B(x[5765]), .Z(n18902) );
  XOR U27368 ( .A(y[5764]), .B(x[5764]), .Z(n18903) );
  XOR U27369 ( .A(y[5763]), .B(x[5763]), .Z(n18901) );
  XNOR U27370 ( .A(n18877), .B(n18878), .Z(n18895) );
  XNOR U27371 ( .A(n18892), .B(n18893), .Z(n18878) );
  XOR U27372 ( .A(n18889), .B(n18888), .Z(n18893) );
  XOR U27373 ( .A(y[5760]), .B(x[5760]), .Z(n18888) );
  XOR U27374 ( .A(n18891), .B(n18890), .Z(n18889) );
  XOR U27375 ( .A(y[5762]), .B(x[5762]), .Z(n18890) );
  XOR U27376 ( .A(y[5761]), .B(x[5761]), .Z(n18891) );
  XOR U27377 ( .A(n18883), .B(n18882), .Z(n18892) );
  XOR U27378 ( .A(n18885), .B(n18884), .Z(n18882) );
  XOR U27379 ( .A(y[5759]), .B(x[5759]), .Z(n18884) );
  XOR U27380 ( .A(y[5758]), .B(x[5758]), .Z(n18885) );
  XOR U27381 ( .A(y[5757]), .B(x[5757]), .Z(n18883) );
  XNOR U27382 ( .A(n18876), .B(n18875), .Z(n18877) );
  XNOR U27383 ( .A(n18872), .B(n18871), .Z(n18875) );
  XOR U27384 ( .A(n18874), .B(n18873), .Z(n18871) );
  XOR U27385 ( .A(y[5756]), .B(x[5756]), .Z(n18873) );
  XOR U27386 ( .A(y[5755]), .B(x[5755]), .Z(n18874) );
  XOR U27387 ( .A(y[5754]), .B(x[5754]), .Z(n18872) );
  XOR U27388 ( .A(n18866), .B(n18865), .Z(n18876) );
  XOR U27389 ( .A(n18868), .B(n18867), .Z(n18865) );
  XOR U27390 ( .A(y[5753]), .B(x[5753]), .Z(n18867) );
  XOR U27391 ( .A(y[5752]), .B(x[5752]), .Z(n18868) );
  XOR U27392 ( .A(y[5751]), .B(x[5751]), .Z(n18866) );
  NAND U27393 ( .A(n18929), .B(n18930), .Z(N63703) );
  NAND U27394 ( .A(n18931), .B(n18932), .Z(n18930) );
  NANDN U27395 ( .A(n18933), .B(n18934), .Z(n18932) );
  NANDN U27396 ( .A(n18934), .B(n18933), .Z(n18929) );
  XOR U27397 ( .A(n18933), .B(n18935), .Z(N63702) );
  XNOR U27398 ( .A(n18931), .B(n18934), .Z(n18935) );
  NAND U27399 ( .A(n18936), .B(n18937), .Z(n18934) );
  NAND U27400 ( .A(n18938), .B(n18939), .Z(n18937) );
  NANDN U27401 ( .A(n18940), .B(n18941), .Z(n18939) );
  NANDN U27402 ( .A(n18941), .B(n18940), .Z(n18936) );
  AND U27403 ( .A(n18942), .B(n18943), .Z(n18931) );
  NAND U27404 ( .A(n18944), .B(n18945), .Z(n18943) );
  NANDN U27405 ( .A(n18946), .B(n18947), .Z(n18945) );
  NANDN U27406 ( .A(n18947), .B(n18946), .Z(n18942) );
  IV U27407 ( .A(n18948), .Z(n18947) );
  AND U27408 ( .A(n18949), .B(n18950), .Z(n18933) );
  NAND U27409 ( .A(n18951), .B(n18952), .Z(n18950) );
  NANDN U27410 ( .A(n18953), .B(n18954), .Z(n18952) );
  NANDN U27411 ( .A(n18954), .B(n18953), .Z(n18949) );
  XOR U27412 ( .A(n18946), .B(n18955), .Z(N63701) );
  XNOR U27413 ( .A(n18944), .B(n18948), .Z(n18955) );
  XOR U27414 ( .A(n18941), .B(n18956), .Z(n18948) );
  XNOR U27415 ( .A(n18938), .B(n18940), .Z(n18956) );
  AND U27416 ( .A(n18957), .B(n18958), .Z(n18940) );
  NANDN U27417 ( .A(n18959), .B(n18960), .Z(n18958) );
  OR U27418 ( .A(n18961), .B(n18962), .Z(n18960) );
  IV U27419 ( .A(n18963), .Z(n18962) );
  NANDN U27420 ( .A(n18963), .B(n18961), .Z(n18957) );
  AND U27421 ( .A(n18964), .B(n18965), .Z(n18938) );
  NAND U27422 ( .A(n18966), .B(n18967), .Z(n18965) );
  NANDN U27423 ( .A(n18968), .B(n18969), .Z(n18967) );
  NANDN U27424 ( .A(n18969), .B(n18968), .Z(n18964) );
  IV U27425 ( .A(n18970), .Z(n18969) );
  NAND U27426 ( .A(n18971), .B(n18972), .Z(n18941) );
  NANDN U27427 ( .A(n18973), .B(n18974), .Z(n18972) );
  NANDN U27428 ( .A(n18975), .B(n18976), .Z(n18974) );
  NANDN U27429 ( .A(n18976), .B(n18975), .Z(n18971) );
  IV U27430 ( .A(n18977), .Z(n18975) );
  AND U27431 ( .A(n18978), .B(n18979), .Z(n18944) );
  NAND U27432 ( .A(n18980), .B(n18981), .Z(n18979) );
  NANDN U27433 ( .A(n18982), .B(n18983), .Z(n18981) );
  NANDN U27434 ( .A(n18983), .B(n18982), .Z(n18978) );
  XOR U27435 ( .A(n18954), .B(n18984), .Z(n18946) );
  XNOR U27436 ( .A(n18951), .B(n18953), .Z(n18984) );
  AND U27437 ( .A(n18985), .B(n18986), .Z(n18953) );
  NANDN U27438 ( .A(n18987), .B(n18988), .Z(n18986) );
  OR U27439 ( .A(n18989), .B(n18990), .Z(n18988) );
  IV U27440 ( .A(n18991), .Z(n18990) );
  NANDN U27441 ( .A(n18991), .B(n18989), .Z(n18985) );
  AND U27442 ( .A(n18992), .B(n18993), .Z(n18951) );
  NAND U27443 ( .A(n18994), .B(n18995), .Z(n18993) );
  NANDN U27444 ( .A(n18996), .B(n18997), .Z(n18995) );
  NANDN U27445 ( .A(n18997), .B(n18996), .Z(n18992) );
  IV U27446 ( .A(n18998), .Z(n18997) );
  NAND U27447 ( .A(n18999), .B(n19000), .Z(n18954) );
  NANDN U27448 ( .A(n19001), .B(n19002), .Z(n19000) );
  NANDN U27449 ( .A(n19003), .B(n19004), .Z(n19002) );
  NANDN U27450 ( .A(n19004), .B(n19003), .Z(n18999) );
  IV U27451 ( .A(n19005), .Z(n19003) );
  XOR U27452 ( .A(n18980), .B(n19006), .Z(N63700) );
  XNOR U27453 ( .A(n18983), .B(n18982), .Z(n19006) );
  XNOR U27454 ( .A(n18994), .B(n19007), .Z(n18982) );
  XNOR U27455 ( .A(n18998), .B(n18996), .Z(n19007) );
  XOR U27456 ( .A(n19004), .B(n19008), .Z(n18996) );
  XNOR U27457 ( .A(n19001), .B(n19005), .Z(n19008) );
  AND U27458 ( .A(n19009), .B(n19010), .Z(n19005) );
  NAND U27459 ( .A(n19011), .B(n19012), .Z(n19010) );
  NAND U27460 ( .A(n19013), .B(n19014), .Z(n19009) );
  AND U27461 ( .A(n19015), .B(n19016), .Z(n19001) );
  NAND U27462 ( .A(n19017), .B(n19018), .Z(n19016) );
  NAND U27463 ( .A(n19019), .B(n19020), .Z(n19015) );
  NANDN U27464 ( .A(n19021), .B(n19022), .Z(n19004) );
  ANDN U27465 ( .B(n19023), .A(n19024), .Z(n18998) );
  XNOR U27466 ( .A(n18989), .B(n19025), .Z(n18994) );
  XNOR U27467 ( .A(n18987), .B(n18991), .Z(n19025) );
  AND U27468 ( .A(n19026), .B(n19027), .Z(n18991) );
  NAND U27469 ( .A(n19028), .B(n19029), .Z(n19027) );
  NAND U27470 ( .A(n19030), .B(n19031), .Z(n19026) );
  AND U27471 ( .A(n19032), .B(n19033), .Z(n18987) );
  NAND U27472 ( .A(n19034), .B(n19035), .Z(n19033) );
  NAND U27473 ( .A(n19036), .B(n19037), .Z(n19032) );
  AND U27474 ( .A(n19038), .B(n19039), .Z(n18989) );
  NAND U27475 ( .A(n19040), .B(n19041), .Z(n18983) );
  XNOR U27476 ( .A(n18966), .B(n19042), .Z(n18980) );
  XNOR U27477 ( .A(n18970), .B(n18968), .Z(n19042) );
  XOR U27478 ( .A(n18976), .B(n19043), .Z(n18968) );
  XNOR U27479 ( .A(n18973), .B(n18977), .Z(n19043) );
  AND U27480 ( .A(n19044), .B(n19045), .Z(n18977) );
  NAND U27481 ( .A(n19046), .B(n19047), .Z(n19045) );
  NAND U27482 ( .A(n19048), .B(n19049), .Z(n19044) );
  AND U27483 ( .A(n19050), .B(n19051), .Z(n18973) );
  NAND U27484 ( .A(n19052), .B(n19053), .Z(n19051) );
  NAND U27485 ( .A(n19054), .B(n19055), .Z(n19050) );
  NANDN U27486 ( .A(n19056), .B(n19057), .Z(n18976) );
  ANDN U27487 ( .B(n19058), .A(n19059), .Z(n18970) );
  XNOR U27488 ( .A(n18961), .B(n19060), .Z(n18966) );
  XNOR U27489 ( .A(n18959), .B(n18963), .Z(n19060) );
  AND U27490 ( .A(n19061), .B(n19062), .Z(n18963) );
  NAND U27491 ( .A(n19063), .B(n19064), .Z(n19062) );
  NAND U27492 ( .A(n19065), .B(n19066), .Z(n19061) );
  AND U27493 ( .A(n19067), .B(n19068), .Z(n18959) );
  NAND U27494 ( .A(n19069), .B(n19070), .Z(n19068) );
  NAND U27495 ( .A(n19071), .B(n19072), .Z(n19067) );
  AND U27496 ( .A(n19073), .B(n19074), .Z(n18961) );
  XOR U27497 ( .A(n19041), .B(n19040), .Z(N63699) );
  XNOR U27498 ( .A(n19058), .B(n19059), .Z(n19040) );
  XNOR U27499 ( .A(n19073), .B(n19074), .Z(n19059) );
  XOR U27500 ( .A(n19070), .B(n19069), .Z(n19074) );
  XOR U27501 ( .A(y[5748]), .B(x[5748]), .Z(n19069) );
  XOR U27502 ( .A(n19072), .B(n19071), .Z(n19070) );
  XOR U27503 ( .A(y[5750]), .B(x[5750]), .Z(n19071) );
  XOR U27504 ( .A(y[5749]), .B(x[5749]), .Z(n19072) );
  XOR U27505 ( .A(n19064), .B(n19063), .Z(n19073) );
  XOR U27506 ( .A(n19066), .B(n19065), .Z(n19063) );
  XOR U27507 ( .A(y[5747]), .B(x[5747]), .Z(n19065) );
  XOR U27508 ( .A(y[5746]), .B(x[5746]), .Z(n19066) );
  XOR U27509 ( .A(y[5745]), .B(x[5745]), .Z(n19064) );
  XNOR U27510 ( .A(n19057), .B(n19056), .Z(n19058) );
  XNOR U27511 ( .A(n19053), .B(n19052), .Z(n19056) );
  XOR U27512 ( .A(n19055), .B(n19054), .Z(n19052) );
  XOR U27513 ( .A(y[5744]), .B(x[5744]), .Z(n19054) );
  XOR U27514 ( .A(y[5743]), .B(x[5743]), .Z(n19055) );
  XOR U27515 ( .A(y[5742]), .B(x[5742]), .Z(n19053) );
  XOR U27516 ( .A(n19047), .B(n19046), .Z(n19057) );
  XOR U27517 ( .A(n19049), .B(n19048), .Z(n19046) );
  XOR U27518 ( .A(y[5741]), .B(x[5741]), .Z(n19048) );
  XOR U27519 ( .A(y[5740]), .B(x[5740]), .Z(n19049) );
  XOR U27520 ( .A(y[5739]), .B(x[5739]), .Z(n19047) );
  XNOR U27521 ( .A(n19023), .B(n19024), .Z(n19041) );
  XNOR U27522 ( .A(n19038), .B(n19039), .Z(n19024) );
  XOR U27523 ( .A(n19035), .B(n19034), .Z(n19039) );
  XOR U27524 ( .A(y[5736]), .B(x[5736]), .Z(n19034) );
  XOR U27525 ( .A(n19037), .B(n19036), .Z(n19035) );
  XOR U27526 ( .A(y[5738]), .B(x[5738]), .Z(n19036) );
  XOR U27527 ( .A(y[5737]), .B(x[5737]), .Z(n19037) );
  XOR U27528 ( .A(n19029), .B(n19028), .Z(n19038) );
  XOR U27529 ( .A(n19031), .B(n19030), .Z(n19028) );
  XOR U27530 ( .A(y[5735]), .B(x[5735]), .Z(n19030) );
  XOR U27531 ( .A(y[5734]), .B(x[5734]), .Z(n19031) );
  XOR U27532 ( .A(y[5733]), .B(x[5733]), .Z(n19029) );
  XNOR U27533 ( .A(n19022), .B(n19021), .Z(n19023) );
  XNOR U27534 ( .A(n19018), .B(n19017), .Z(n19021) );
  XOR U27535 ( .A(n19020), .B(n19019), .Z(n19017) );
  XOR U27536 ( .A(y[5732]), .B(x[5732]), .Z(n19019) );
  XOR U27537 ( .A(y[5731]), .B(x[5731]), .Z(n19020) );
  XOR U27538 ( .A(y[5730]), .B(x[5730]), .Z(n19018) );
  XOR U27539 ( .A(n19012), .B(n19011), .Z(n19022) );
  XOR U27540 ( .A(n19014), .B(n19013), .Z(n19011) );
  XOR U27541 ( .A(y[5729]), .B(x[5729]), .Z(n19013) );
  XOR U27542 ( .A(y[5728]), .B(x[5728]), .Z(n19014) );
  XOR U27543 ( .A(y[5727]), .B(x[5727]), .Z(n19012) );
  NAND U27544 ( .A(n19075), .B(n19076), .Z(N63690) );
  NAND U27545 ( .A(n19077), .B(n19078), .Z(n19076) );
  NANDN U27546 ( .A(n19079), .B(n19080), .Z(n19078) );
  NANDN U27547 ( .A(n19080), .B(n19079), .Z(n19075) );
  XOR U27548 ( .A(n19079), .B(n19081), .Z(N63689) );
  XNOR U27549 ( .A(n19077), .B(n19080), .Z(n19081) );
  NAND U27550 ( .A(n19082), .B(n19083), .Z(n19080) );
  NAND U27551 ( .A(n19084), .B(n19085), .Z(n19083) );
  NANDN U27552 ( .A(n19086), .B(n19087), .Z(n19085) );
  NANDN U27553 ( .A(n19087), .B(n19086), .Z(n19082) );
  AND U27554 ( .A(n19088), .B(n19089), .Z(n19077) );
  NAND U27555 ( .A(n19090), .B(n19091), .Z(n19089) );
  NANDN U27556 ( .A(n19092), .B(n19093), .Z(n19091) );
  NANDN U27557 ( .A(n19093), .B(n19092), .Z(n19088) );
  IV U27558 ( .A(n19094), .Z(n19093) );
  AND U27559 ( .A(n19095), .B(n19096), .Z(n19079) );
  NAND U27560 ( .A(n19097), .B(n19098), .Z(n19096) );
  NANDN U27561 ( .A(n19099), .B(n19100), .Z(n19098) );
  NANDN U27562 ( .A(n19100), .B(n19099), .Z(n19095) );
  XOR U27563 ( .A(n19092), .B(n19101), .Z(N63688) );
  XNOR U27564 ( .A(n19090), .B(n19094), .Z(n19101) );
  XOR U27565 ( .A(n19087), .B(n19102), .Z(n19094) );
  XNOR U27566 ( .A(n19084), .B(n19086), .Z(n19102) );
  AND U27567 ( .A(n19103), .B(n19104), .Z(n19086) );
  NANDN U27568 ( .A(n19105), .B(n19106), .Z(n19104) );
  OR U27569 ( .A(n19107), .B(n19108), .Z(n19106) );
  IV U27570 ( .A(n19109), .Z(n19108) );
  NANDN U27571 ( .A(n19109), .B(n19107), .Z(n19103) );
  AND U27572 ( .A(n19110), .B(n19111), .Z(n19084) );
  NAND U27573 ( .A(n19112), .B(n19113), .Z(n19111) );
  NANDN U27574 ( .A(n19114), .B(n19115), .Z(n19113) );
  NANDN U27575 ( .A(n19115), .B(n19114), .Z(n19110) );
  IV U27576 ( .A(n19116), .Z(n19115) );
  NAND U27577 ( .A(n19117), .B(n19118), .Z(n19087) );
  NANDN U27578 ( .A(n19119), .B(n19120), .Z(n19118) );
  NANDN U27579 ( .A(n19121), .B(n19122), .Z(n19120) );
  NANDN U27580 ( .A(n19122), .B(n19121), .Z(n19117) );
  IV U27581 ( .A(n19123), .Z(n19121) );
  AND U27582 ( .A(n19124), .B(n19125), .Z(n19090) );
  NAND U27583 ( .A(n19126), .B(n19127), .Z(n19125) );
  NANDN U27584 ( .A(n19128), .B(n19129), .Z(n19127) );
  NANDN U27585 ( .A(n19129), .B(n19128), .Z(n19124) );
  XOR U27586 ( .A(n19100), .B(n19130), .Z(n19092) );
  XNOR U27587 ( .A(n19097), .B(n19099), .Z(n19130) );
  AND U27588 ( .A(n19131), .B(n19132), .Z(n19099) );
  NANDN U27589 ( .A(n19133), .B(n19134), .Z(n19132) );
  OR U27590 ( .A(n19135), .B(n19136), .Z(n19134) );
  IV U27591 ( .A(n19137), .Z(n19136) );
  NANDN U27592 ( .A(n19137), .B(n19135), .Z(n19131) );
  AND U27593 ( .A(n19138), .B(n19139), .Z(n19097) );
  NAND U27594 ( .A(n19140), .B(n19141), .Z(n19139) );
  NANDN U27595 ( .A(n19142), .B(n19143), .Z(n19141) );
  NANDN U27596 ( .A(n19143), .B(n19142), .Z(n19138) );
  IV U27597 ( .A(n19144), .Z(n19143) );
  NAND U27598 ( .A(n19145), .B(n19146), .Z(n19100) );
  NANDN U27599 ( .A(n19147), .B(n19148), .Z(n19146) );
  NANDN U27600 ( .A(n19149), .B(n19150), .Z(n19148) );
  NANDN U27601 ( .A(n19150), .B(n19149), .Z(n19145) );
  IV U27602 ( .A(n19151), .Z(n19149) );
  XOR U27603 ( .A(n19126), .B(n19152), .Z(N63687) );
  XNOR U27604 ( .A(n19129), .B(n19128), .Z(n19152) );
  XNOR U27605 ( .A(n19140), .B(n19153), .Z(n19128) );
  XNOR U27606 ( .A(n19144), .B(n19142), .Z(n19153) );
  XOR U27607 ( .A(n19150), .B(n19154), .Z(n19142) );
  XNOR U27608 ( .A(n19147), .B(n19151), .Z(n19154) );
  AND U27609 ( .A(n19155), .B(n19156), .Z(n19151) );
  NAND U27610 ( .A(n19157), .B(n19158), .Z(n19156) );
  NAND U27611 ( .A(n19159), .B(n19160), .Z(n19155) );
  AND U27612 ( .A(n19161), .B(n19162), .Z(n19147) );
  NAND U27613 ( .A(n19163), .B(n19164), .Z(n19162) );
  NAND U27614 ( .A(n19165), .B(n19166), .Z(n19161) );
  NANDN U27615 ( .A(n19167), .B(n19168), .Z(n19150) );
  ANDN U27616 ( .B(n19169), .A(n19170), .Z(n19144) );
  XNOR U27617 ( .A(n19135), .B(n19171), .Z(n19140) );
  XNOR U27618 ( .A(n19133), .B(n19137), .Z(n19171) );
  AND U27619 ( .A(n19172), .B(n19173), .Z(n19137) );
  NAND U27620 ( .A(n19174), .B(n19175), .Z(n19173) );
  NAND U27621 ( .A(n19176), .B(n19177), .Z(n19172) );
  AND U27622 ( .A(n19178), .B(n19179), .Z(n19133) );
  NAND U27623 ( .A(n19180), .B(n19181), .Z(n19179) );
  NAND U27624 ( .A(n19182), .B(n19183), .Z(n19178) );
  AND U27625 ( .A(n19184), .B(n19185), .Z(n19135) );
  NAND U27626 ( .A(n19186), .B(n19187), .Z(n19129) );
  XNOR U27627 ( .A(n19112), .B(n19188), .Z(n19126) );
  XNOR U27628 ( .A(n19116), .B(n19114), .Z(n19188) );
  XOR U27629 ( .A(n19122), .B(n19189), .Z(n19114) );
  XNOR U27630 ( .A(n19119), .B(n19123), .Z(n19189) );
  AND U27631 ( .A(n19190), .B(n19191), .Z(n19123) );
  NAND U27632 ( .A(n19192), .B(n19193), .Z(n19191) );
  NAND U27633 ( .A(n19194), .B(n19195), .Z(n19190) );
  AND U27634 ( .A(n19196), .B(n19197), .Z(n19119) );
  NAND U27635 ( .A(n19198), .B(n19199), .Z(n19197) );
  NAND U27636 ( .A(n19200), .B(n19201), .Z(n19196) );
  NANDN U27637 ( .A(n19202), .B(n19203), .Z(n19122) );
  ANDN U27638 ( .B(n19204), .A(n19205), .Z(n19116) );
  XNOR U27639 ( .A(n19107), .B(n19206), .Z(n19112) );
  XNOR U27640 ( .A(n19105), .B(n19109), .Z(n19206) );
  AND U27641 ( .A(n19207), .B(n19208), .Z(n19109) );
  NAND U27642 ( .A(n19209), .B(n19210), .Z(n19208) );
  NAND U27643 ( .A(n19211), .B(n19212), .Z(n19207) );
  AND U27644 ( .A(n19213), .B(n19214), .Z(n19105) );
  NAND U27645 ( .A(n19215), .B(n19216), .Z(n19214) );
  NAND U27646 ( .A(n19217), .B(n19218), .Z(n19213) );
  AND U27647 ( .A(n19219), .B(n19220), .Z(n19107) );
  XOR U27648 ( .A(n19187), .B(n19186), .Z(N63686) );
  XNOR U27649 ( .A(n19204), .B(n19205), .Z(n19186) );
  XNOR U27650 ( .A(n19219), .B(n19220), .Z(n19205) );
  XOR U27651 ( .A(n19216), .B(n19215), .Z(n19220) );
  XOR U27652 ( .A(y[5724]), .B(x[5724]), .Z(n19215) );
  XOR U27653 ( .A(n19218), .B(n19217), .Z(n19216) );
  XOR U27654 ( .A(y[5726]), .B(x[5726]), .Z(n19217) );
  XOR U27655 ( .A(y[5725]), .B(x[5725]), .Z(n19218) );
  XOR U27656 ( .A(n19210), .B(n19209), .Z(n19219) );
  XOR U27657 ( .A(n19212), .B(n19211), .Z(n19209) );
  XOR U27658 ( .A(y[5723]), .B(x[5723]), .Z(n19211) );
  XOR U27659 ( .A(y[5722]), .B(x[5722]), .Z(n19212) );
  XOR U27660 ( .A(y[5721]), .B(x[5721]), .Z(n19210) );
  XNOR U27661 ( .A(n19203), .B(n19202), .Z(n19204) );
  XNOR U27662 ( .A(n19199), .B(n19198), .Z(n19202) );
  XOR U27663 ( .A(n19201), .B(n19200), .Z(n19198) );
  XOR U27664 ( .A(y[5720]), .B(x[5720]), .Z(n19200) );
  XOR U27665 ( .A(y[5719]), .B(x[5719]), .Z(n19201) );
  XOR U27666 ( .A(y[5718]), .B(x[5718]), .Z(n19199) );
  XOR U27667 ( .A(n19193), .B(n19192), .Z(n19203) );
  XOR U27668 ( .A(n19195), .B(n19194), .Z(n19192) );
  XOR U27669 ( .A(y[5717]), .B(x[5717]), .Z(n19194) );
  XOR U27670 ( .A(y[5716]), .B(x[5716]), .Z(n19195) );
  XOR U27671 ( .A(y[5715]), .B(x[5715]), .Z(n19193) );
  XNOR U27672 ( .A(n19169), .B(n19170), .Z(n19187) );
  XNOR U27673 ( .A(n19184), .B(n19185), .Z(n19170) );
  XOR U27674 ( .A(n19181), .B(n19180), .Z(n19185) );
  XOR U27675 ( .A(y[5712]), .B(x[5712]), .Z(n19180) );
  XOR U27676 ( .A(n19183), .B(n19182), .Z(n19181) );
  XOR U27677 ( .A(y[5714]), .B(x[5714]), .Z(n19182) );
  XOR U27678 ( .A(y[5713]), .B(x[5713]), .Z(n19183) );
  XOR U27679 ( .A(n19175), .B(n19174), .Z(n19184) );
  XOR U27680 ( .A(n19177), .B(n19176), .Z(n19174) );
  XOR U27681 ( .A(y[5711]), .B(x[5711]), .Z(n19176) );
  XOR U27682 ( .A(y[5710]), .B(x[5710]), .Z(n19177) );
  XOR U27683 ( .A(y[5709]), .B(x[5709]), .Z(n19175) );
  XNOR U27684 ( .A(n19168), .B(n19167), .Z(n19169) );
  XNOR U27685 ( .A(n19164), .B(n19163), .Z(n19167) );
  XOR U27686 ( .A(n19166), .B(n19165), .Z(n19163) );
  XOR U27687 ( .A(y[5708]), .B(x[5708]), .Z(n19165) );
  XOR U27688 ( .A(y[5707]), .B(x[5707]), .Z(n19166) );
  XOR U27689 ( .A(y[5706]), .B(x[5706]), .Z(n19164) );
  XOR U27690 ( .A(n19158), .B(n19157), .Z(n19168) );
  XOR U27691 ( .A(n19160), .B(n19159), .Z(n19157) );
  XOR U27692 ( .A(y[5705]), .B(x[5705]), .Z(n19159) );
  XOR U27693 ( .A(y[5704]), .B(x[5704]), .Z(n19160) );
  XOR U27694 ( .A(y[5703]), .B(x[5703]), .Z(n19158) );
  NAND U27695 ( .A(n19221), .B(n19222), .Z(N63677) );
  NAND U27696 ( .A(n19223), .B(n19224), .Z(n19222) );
  NANDN U27697 ( .A(n19225), .B(n19226), .Z(n19224) );
  NANDN U27698 ( .A(n19226), .B(n19225), .Z(n19221) );
  XOR U27699 ( .A(n19225), .B(n19227), .Z(N63676) );
  XNOR U27700 ( .A(n19223), .B(n19226), .Z(n19227) );
  NAND U27701 ( .A(n19228), .B(n19229), .Z(n19226) );
  NAND U27702 ( .A(n19230), .B(n19231), .Z(n19229) );
  NANDN U27703 ( .A(n19232), .B(n19233), .Z(n19231) );
  NANDN U27704 ( .A(n19233), .B(n19232), .Z(n19228) );
  AND U27705 ( .A(n19234), .B(n19235), .Z(n19223) );
  NAND U27706 ( .A(n19236), .B(n19237), .Z(n19235) );
  NANDN U27707 ( .A(n19238), .B(n19239), .Z(n19237) );
  NANDN U27708 ( .A(n19239), .B(n19238), .Z(n19234) );
  IV U27709 ( .A(n19240), .Z(n19239) );
  AND U27710 ( .A(n19241), .B(n19242), .Z(n19225) );
  NAND U27711 ( .A(n19243), .B(n19244), .Z(n19242) );
  NANDN U27712 ( .A(n19245), .B(n19246), .Z(n19244) );
  NANDN U27713 ( .A(n19246), .B(n19245), .Z(n19241) );
  XOR U27714 ( .A(n19238), .B(n19247), .Z(N63675) );
  XNOR U27715 ( .A(n19236), .B(n19240), .Z(n19247) );
  XOR U27716 ( .A(n19233), .B(n19248), .Z(n19240) );
  XNOR U27717 ( .A(n19230), .B(n19232), .Z(n19248) );
  AND U27718 ( .A(n19249), .B(n19250), .Z(n19232) );
  NANDN U27719 ( .A(n19251), .B(n19252), .Z(n19250) );
  OR U27720 ( .A(n19253), .B(n19254), .Z(n19252) );
  IV U27721 ( .A(n19255), .Z(n19254) );
  NANDN U27722 ( .A(n19255), .B(n19253), .Z(n19249) );
  AND U27723 ( .A(n19256), .B(n19257), .Z(n19230) );
  NAND U27724 ( .A(n19258), .B(n19259), .Z(n19257) );
  NANDN U27725 ( .A(n19260), .B(n19261), .Z(n19259) );
  NANDN U27726 ( .A(n19261), .B(n19260), .Z(n19256) );
  IV U27727 ( .A(n19262), .Z(n19261) );
  NAND U27728 ( .A(n19263), .B(n19264), .Z(n19233) );
  NANDN U27729 ( .A(n19265), .B(n19266), .Z(n19264) );
  NANDN U27730 ( .A(n19267), .B(n19268), .Z(n19266) );
  NANDN U27731 ( .A(n19268), .B(n19267), .Z(n19263) );
  IV U27732 ( .A(n19269), .Z(n19267) );
  AND U27733 ( .A(n19270), .B(n19271), .Z(n19236) );
  NAND U27734 ( .A(n19272), .B(n19273), .Z(n19271) );
  NANDN U27735 ( .A(n19274), .B(n19275), .Z(n19273) );
  NANDN U27736 ( .A(n19275), .B(n19274), .Z(n19270) );
  XOR U27737 ( .A(n19246), .B(n19276), .Z(n19238) );
  XNOR U27738 ( .A(n19243), .B(n19245), .Z(n19276) );
  AND U27739 ( .A(n19277), .B(n19278), .Z(n19245) );
  NANDN U27740 ( .A(n19279), .B(n19280), .Z(n19278) );
  OR U27741 ( .A(n19281), .B(n19282), .Z(n19280) );
  IV U27742 ( .A(n19283), .Z(n19282) );
  NANDN U27743 ( .A(n19283), .B(n19281), .Z(n19277) );
  AND U27744 ( .A(n19284), .B(n19285), .Z(n19243) );
  NAND U27745 ( .A(n19286), .B(n19287), .Z(n19285) );
  NANDN U27746 ( .A(n19288), .B(n19289), .Z(n19287) );
  NANDN U27747 ( .A(n19289), .B(n19288), .Z(n19284) );
  IV U27748 ( .A(n19290), .Z(n19289) );
  NAND U27749 ( .A(n19291), .B(n19292), .Z(n19246) );
  NANDN U27750 ( .A(n19293), .B(n19294), .Z(n19292) );
  NANDN U27751 ( .A(n19295), .B(n19296), .Z(n19294) );
  NANDN U27752 ( .A(n19296), .B(n19295), .Z(n19291) );
  IV U27753 ( .A(n19297), .Z(n19295) );
  XOR U27754 ( .A(n19272), .B(n19298), .Z(N63674) );
  XNOR U27755 ( .A(n19275), .B(n19274), .Z(n19298) );
  XNOR U27756 ( .A(n19286), .B(n19299), .Z(n19274) );
  XNOR U27757 ( .A(n19290), .B(n19288), .Z(n19299) );
  XOR U27758 ( .A(n19296), .B(n19300), .Z(n19288) );
  XNOR U27759 ( .A(n19293), .B(n19297), .Z(n19300) );
  AND U27760 ( .A(n19301), .B(n19302), .Z(n19297) );
  NAND U27761 ( .A(n19303), .B(n19304), .Z(n19302) );
  NAND U27762 ( .A(n19305), .B(n19306), .Z(n19301) );
  AND U27763 ( .A(n19307), .B(n19308), .Z(n19293) );
  NAND U27764 ( .A(n19309), .B(n19310), .Z(n19308) );
  NAND U27765 ( .A(n19311), .B(n19312), .Z(n19307) );
  NANDN U27766 ( .A(n19313), .B(n19314), .Z(n19296) );
  ANDN U27767 ( .B(n19315), .A(n19316), .Z(n19290) );
  XNOR U27768 ( .A(n19281), .B(n19317), .Z(n19286) );
  XNOR U27769 ( .A(n19279), .B(n19283), .Z(n19317) );
  AND U27770 ( .A(n19318), .B(n19319), .Z(n19283) );
  NAND U27771 ( .A(n19320), .B(n19321), .Z(n19319) );
  NAND U27772 ( .A(n19322), .B(n19323), .Z(n19318) );
  AND U27773 ( .A(n19324), .B(n19325), .Z(n19279) );
  NAND U27774 ( .A(n19326), .B(n19327), .Z(n19325) );
  NAND U27775 ( .A(n19328), .B(n19329), .Z(n19324) );
  AND U27776 ( .A(n19330), .B(n19331), .Z(n19281) );
  NAND U27777 ( .A(n19332), .B(n19333), .Z(n19275) );
  XNOR U27778 ( .A(n19258), .B(n19334), .Z(n19272) );
  XNOR U27779 ( .A(n19262), .B(n19260), .Z(n19334) );
  XOR U27780 ( .A(n19268), .B(n19335), .Z(n19260) );
  XNOR U27781 ( .A(n19265), .B(n19269), .Z(n19335) );
  AND U27782 ( .A(n19336), .B(n19337), .Z(n19269) );
  NAND U27783 ( .A(n19338), .B(n19339), .Z(n19337) );
  NAND U27784 ( .A(n19340), .B(n19341), .Z(n19336) );
  AND U27785 ( .A(n19342), .B(n19343), .Z(n19265) );
  NAND U27786 ( .A(n19344), .B(n19345), .Z(n19343) );
  NAND U27787 ( .A(n19346), .B(n19347), .Z(n19342) );
  NANDN U27788 ( .A(n19348), .B(n19349), .Z(n19268) );
  ANDN U27789 ( .B(n19350), .A(n19351), .Z(n19262) );
  XNOR U27790 ( .A(n19253), .B(n19352), .Z(n19258) );
  XNOR U27791 ( .A(n19251), .B(n19255), .Z(n19352) );
  AND U27792 ( .A(n19353), .B(n19354), .Z(n19255) );
  NAND U27793 ( .A(n19355), .B(n19356), .Z(n19354) );
  NAND U27794 ( .A(n19357), .B(n19358), .Z(n19353) );
  AND U27795 ( .A(n19359), .B(n19360), .Z(n19251) );
  NAND U27796 ( .A(n19361), .B(n19362), .Z(n19360) );
  NAND U27797 ( .A(n19363), .B(n19364), .Z(n19359) );
  AND U27798 ( .A(n19365), .B(n19366), .Z(n19253) );
  XOR U27799 ( .A(n19333), .B(n19332), .Z(N63673) );
  XNOR U27800 ( .A(n19350), .B(n19351), .Z(n19332) );
  XNOR U27801 ( .A(n19365), .B(n19366), .Z(n19351) );
  XOR U27802 ( .A(n19362), .B(n19361), .Z(n19366) );
  XOR U27803 ( .A(y[5700]), .B(x[5700]), .Z(n19361) );
  XOR U27804 ( .A(n19364), .B(n19363), .Z(n19362) );
  XOR U27805 ( .A(y[5702]), .B(x[5702]), .Z(n19363) );
  XOR U27806 ( .A(y[5701]), .B(x[5701]), .Z(n19364) );
  XOR U27807 ( .A(n19356), .B(n19355), .Z(n19365) );
  XOR U27808 ( .A(n19358), .B(n19357), .Z(n19355) );
  XOR U27809 ( .A(y[5699]), .B(x[5699]), .Z(n19357) );
  XOR U27810 ( .A(y[5698]), .B(x[5698]), .Z(n19358) );
  XOR U27811 ( .A(y[5697]), .B(x[5697]), .Z(n19356) );
  XNOR U27812 ( .A(n19349), .B(n19348), .Z(n19350) );
  XNOR U27813 ( .A(n19345), .B(n19344), .Z(n19348) );
  XOR U27814 ( .A(n19347), .B(n19346), .Z(n19344) );
  XOR U27815 ( .A(y[5696]), .B(x[5696]), .Z(n19346) );
  XOR U27816 ( .A(y[5695]), .B(x[5695]), .Z(n19347) );
  XOR U27817 ( .A(y[5694]), .B(x[5694]), .Z(n19345) );
  XOR U27818 ( .A(n19339), .B(n19338), .Z(n19349) );
  XOR U27819 ( .A(n19341), .B(n19340), .Z(n19338) );
  XOR U27820 ( .A(y[5693]), .B(x[5693]), .Z(n19340) );
  XOR U27821 ( .A(y[5692]), .B(x[5692]), .Z(n19341) );
  XOR U27822 ( .A(y[5691]), .B(x[5691]), .Z(n19339) );
  XNOR U27823 ( .A(n19315), .B(n19316), .Z(n19333) );
  XNOR U27824 ( .A(n19330), .B(n19331), .Z(n19316) );
  XOR U27825 ( .A(n19327), .B(n19326), .Z(n19331) );
  XOR U27826 ( .A(y[5688]), .B(x[5688]), .Z(n19326) );
  XOR U27827 ( .A(n19329), .B(n19328), .Z(n19327) );
  XOR U27828 ( .A(y[5690]), .B(x[5690]), .Z(n19328) );
  XOR U27829 ( .A(y[5689]), .B(x[5689]), .Z(n19329) );
  XOR U27830 ( .A(n19321), .B(n19320), .Z(n19330) );
  XOR U27831 ( .A(n19323), .B(n19322), .Z(n19320) );
  XOR U27832 ( .A(y[5687]), .B(x[5687]), .Z(n19322) );
  XOR U27833 ( .A(y[5686]), .B(x[5686]), .Z(n19323) );
  XOR U27834 ( .A(y[5685]), .B(x[5685]), .Z(n19321) );
  XNOR U27835 ( .A(n19314), .B(n19313), .Z(n19315) );
  XNOR U27836 ( .A(n19310), .B(n19309), .Z(n19313) );
  XOR U27837 ( .A(n19312), .B(n19311), .Z(n19309) );
  XOR U27838 ( .A(y[5684]), .B(x[5684]), .Z(n19311) );
  XOR U27839 ( .A(y[5683]), .B(x[5683]), .Z(n19312) );
  XOR U27840 ( .A(y[5682]), .B(x[5682]), .Z(n19310) );
  XOR U27841 ( .A(n19304), .B(n19303), .Z(n19314) );
  XOR U27842 ( .A(n19306), .B(n19305), .Z(n19303) );
  XOR U27843 ( .A(y[5681]), .B(x[5681]), .Z(n19305) );
  XOR U27844 ( .A(y[5680]), .B(x[5680]), .Z(n19306) );
  XOR U27845 ( .A(y[5679]), .B(x[5679]), .Z(n19304) );
  NAND U27846 ( .A(n19367), .B(n19368), .Z(N63664) );
  NAND U27847 ( .A(n19369), .B(n19370), .Z(n19368) );
  NANDN U27848 ( .A(n19371), .B(n19372), .Z(n19370) );
  NANDN U27849 ( .A(n19372), .B(n19371), .Z(n19367) );
  XOR U27850 ( .A(n19371), .B(n19373), .Z(N63663) );
  XNOR U27851 ( .A(n19369), .B(n19372), .Z(n19373) );
  NAND U27852 ( .A(n19374), .B(n19375), .Z(n19372) );
  NAND U27853 ( .A(n19376), .B(n19377), .Z(n19375) );
  NANDN U27854 ( .A(n19378), .B(n19379), .Z(n19377) );
  NANDN U27855 ( .A(n19379), .B(n19378), .Z(n19374) );
  AND U27856 ( .A(n19380), .B(n19381), .Z(n19369) );
  NAND U27857 ( .A(n19382), .B(n19383), .Z(n19381) );
  NANDN U27858 ( .A(n19384), .B(n19385), .Z(n19383) );
  NANDN U27859 ( .A(n19385), .B(n19384), .Z(n19380) );
  IV U27860 ( .A(n19386), .Z(n19385) );
  AND U27861 ( .A(n19387), .B(n19388), .Z(n19371) );
  NAND U27862 ( .A(n19389), .B(n19390), .Z(n19388) );
  NANDN U27863 ( .A(n19391), .B(n19392), .Z(n19390) );
  NANDN U27864 ( .A(n19392), .B(n19391), .Z(n19387) );
  XOR U27865 ( .A(n19384), .B(n19393), .Z(N63662) );
  XNOR U27866 ( .A(n19382), .B(n19386), .Z(n19393) );
  XOR U27867 ( .A(n19379), .B(n19394), .Z(n19386) );
  XNOR U27868 ( .A(n19376), .B(n19378), .Z(n19394) );
  AND U27869 ( .A(n19395), .B(n19396), .Z(n19378) );
  NANDN U27870 ( .A(n19397), .B(n19398), .Z(n19396) );
  OR U27871 ( .A(n19399), .B(n19400), .Z(n19398) );
  IV U27872 ( .A(n19401), .Z(n19400) );
  NANDN U27873 ( .A(n19401), .B(n19399), .Z(n19395) );
  AND U27874 ( .A(n19402), .B(n19403), .Z(n19376) );
  NAND U27875 ( .A(n19404), .B(n19405), .Z(n19403) );
  NANDN U27876 ( .A(n19406), .B(n19407), .Z(n19405) );
  NANDN U27877 ( .A(n19407), .B(n19406), .Z(n19402) );
  IV U27878 ( .A(n19408), .Z(n19407) );
  NAND U27879 ( .A(n19409), .B(n19410), .Z(n19379) );
  NANDN U27880 ( .A(n19411), .B(n19412), .Z(n19410) );
  NANDN U27881 ( .A(n19413), .B(n19414), .Z(n19412) );
  NANDN U27882 ( .A(n19414), .B(n19413), .Z(n19409) );
  IV U27883 ( .A(n19415), .Z(n19413) );
  AND U27884 ( .A(n19416), .B(n19417), .Z(n19382) );
  NAND U27885 ( .A(n19418), .B(n19419), .Z(n19417) );
  NANDN U27886 ( .A(n19420), .B(n19421), .Z(n19419) );
  NANDN U27887 ( .A(n19421), .B(n19420), .Z(n19416) );
  XOR U27888 ( .A(n19392), .B(n19422), .Z(n19384) );
  XNOR U27889 ( .A(n19389), .B(n19391), .Z(n19422) );
  AND U27890 ( .A(n19423), .B(n19424), .Z(n19391) );
  NANDN U27891 ( .A(n19425), .B(n19426), .Z(n19424) );
  OR U27892 ( .A(n19427), .B(n19428), .Z(n19426) );
  IV U27893 ( .A(n19429), .Z(n19428) );
  NANDN U27894 ( .A(n19429), .B(n19427), .Z(n19423) );
  AND U27895 ( .A(n19430), .B(n19431), .Z(n19389) );
  NAND U27896 ( .A(n19432), .B(n19433), .Z(n19431) );
  NANDN U27897 ( .A(n19434), .B(n19435), .Z(n19433) );
  NANDN U27898 ( .A(n19435), .B(n19434), .Z(n19430) );
  IV U27899 ( .A(n19436), .Z(n19435) );
  NAND U27900 ( .A(n19437), .B(n19438), .Z(n19392) );
  NANDN U27901 ( .A(n19439), .B(n19440), .Z(n19438) );
  NANDN U27902 ( .A(n19441), .B(n19442), .Z(n19440) );
  NANDN U27903 ( .A(n19442), .B(n19441), .Z(n19437) );
  IV U27904 ( .A(n19443), .Z(n19441) );
  XOR U27905 ( .A(n19418), .B(n19444), .Z(N63661) );
  XNOR U27906 ( .A(n19421), .B(n19420), .Z(n19444) );
  XNOR U27907 ( .A(n19432), .B(n19445), .Z(n19420) );
  XNOR U27908 ( .A(n19436), .B(n19434), .Z(n19445) );
  XOR U27909 ( .A(n19442), .B(n19446), .Z(n19434) );
  XNOR U27910 ( .A(n19439), .B(n19443), .Z(n19446) );
  AND U27911 ( .A(n19447), .B(n19448), .Z(n19443) );
  NAND U27912 ( .A(n19449), .B(n19450), .Z(n19448) );
  NAND U27913 ( .A(n19451), .B(n19452), .Z(n19447) );
  AND U27914 ( .A(n19453), .B(n19454), .Z(n19439) );
  NAND U27915 ( .A(n19455), .B(n19456), .Z(n19454) );
  NAND U27916 ( .A(n19457), .B(n19458), .Z(n19453) );
  NANDN U27917 ( .A(n19459), .B(n19460), .Z(n19442) );
  ANDN U27918 ( .B(n19461), .A(n19462), .Z(n19436) );
  XNOR U27919 ( .A(n19427), .B(n19463), .Z(n19432) );
  XNOR U27920 ( .A(n19425), .B(n19429), .Z(n19463) );
  AND U27921 ( .A(n19464), .B(n19465), .Z(n19429) );
  NAND U27922 ( .A(n19466), .B(n19467), .Z(n19465) );
  NAND U27923 ( .A(n19468), .B(n19469), .Z(n19464) );
  AND U27924 ( .A(n19470), .B(n19471), .Z(n19425) );
  NAND U27925 ( .A(n19472), .B(n19473), .Z(n19471) );
  NAND U27926 ( .A(n19474), .B(n19475), .Z(n19470) );
  AND U27927 ( .A(n19476), .B(n19477), .Z(n19427) );
  NAND U27928 ( .A(n19478), .B(n19479), .Z(n19421) );
  XNOR U27929 ( .A(n19404), .B(n19480), .Z(n19418) );
  XNOR U27930 ( .A(n19408), .B(n19406), .Z(n19480) );
  XOR U27931 ( .A(n19414), .B(n19481), .Z(n19406) );
  XNOR U27932 ( .A(n19411), .B(n19415), .Z(n19481) );
  AND U27933 ( .A(n19482), .B(n19483), .Z(n19415) );
  NAND U27934 ( .A(n19484), .B(n19485), .Z(n19483) );
  NAND U27935 ( .A(n19486), .B(n19487), .Z(n19482) );
  AND U27936 ( .A(n19488), .B(n19489), .Z(n19411) );
  NAND U27937 ( .A(n19490), .B(n19491), .Z(n19489) );
  NAND U27938 ( .A(n19492), .B(n19493), .Z(n19488) );
  NANDN U27939 ( .A(n19494), .B(n19495), .Z(n19414) );
  ANDN U27940 ( .B(n19496), .A(n19497), .Z(n19408) );
  XNOR U27941 ( .A(n19399), .B(n19498), .Z(n19404) );
  XNOR U27942 ( .A(n19397), .B(n19401), .Z(n19498) );
  AND U27943 ( .A(n19499), .B(n19500), .Z(n19401) );
  NAND U27944 ( .A(n19501), .B(n19502), .Z(n19500) );
  NAND U27945 ( .A(n19503), .B(n19504), .Z(n19499) );
  AND U27946 ( .A(n19505), .B(n19506), .Z(n19397) );
  NAND U27947 ( .A(n19507), .B(n19508), .Z(n19506) );
  NAND U27948 ( .A(n19509), .B(n19510), .Z(n19505) );
  AND U27949 ( .A(n19511), .B(n19512), .Z(n19399) );
  XOR U27950 ( .A(n19479), .B(n19478), .Z(N63660) );
  XNOR U27951 ( .A(n19496), .B(n19497), .Z(n19478) );
  XNOR U27952 ( .A(n19511), .B(n19512), .Z(n19497) );
  XOR U27953 ( .A(n19508), .B(n19507), .Z(n19512) );
  XOR U27954 ( .A(y[5676]), .B(x[5676]), .Z(n19507) );
  XOR U27955 ( .A(n19510), .B(n19509), .Z(n19508) );
  XOR U27956 ( .A(y[5678]), .B(x[5678]), .Z(n19509) );
  XOR U27957 ( .A(y[5677]), .B(x[5677]), .Z(n19510) );
  XOR U27958 ( .A(n19502), .B(n19501), .Z(n19511) );
  XOR U27959 ( .A(n19504), .B(n19503), .Z(n19501) );
  XOR U27960 ( .A(y[5675]), .B(x[5675]), .Z(n19503) );
  XOR U27961 ( .A(y[5674]), .B(x[5674]), .Z(n19504) );
  XOR U27962 ( .A(y[5673]), .B(x[5673]), .Z(n19502) );
  XNOR U27963 ( .A(n19495), .B(n19494), .Z(n19496) );
  XNOR U27964 ( .A(n19491), .B(n19490), .Z(n19494) );
  XOR U27965 ( .A(n19493), .B(n19492), .Z(n19490) );
  XOR U27966 ( .A(y[5672]), .B(x[5672]), .Z(n19492) );
  XOR U27967 ( .A(y[5671]), .B(x[5671]), .Z(n19493) );
  XOR U27968 ( .A(y[5670]), .B(x[5670]), .Z(n19491) );
  XOR U27969 ( .A(n19485), .B(n19484), .Z(n19495) );
  XOR U27970 ( .A(n19487), .B(n19486), .Z(n19484) );
  XOR U27971 ( .A(y[5669]), .B(x[5669]), .Z(n19486) );
  XOR U27972 ( .A(y[5668]), .B(x[5668]), .Z(n19487) );
  XOR U27973 ( .A(y[5667]), .B(x[5667]), .Z(n19485) );
  XNOR U27974 ( .A(n19461), .B(n19462), .Z(n19479) );
  XNOR U27975 ( .A(n19476), .B(n19477), .Z(n19462) );
  XOR U27976 ( .A(n19473), .B(n19472), .Z(n19477) );
  XOR U27977 ( .A(y[5664]), .B(x[5664]), .Z(n19472) );
  XOR U27978 ( .A(n19475), .B(n19474), .Z(n19473) );
  XOR U27979 ( .A(y[5666]), .B(x[5666]), .Z(n19474) );
  XOR U27980 ( .A(y[5665]), .B(x[5665]), .Z(n19475) );
  XOR U27981 ( .A(n19467), .B(n19466), .Z(n19476) );
  XOR U27982 ( .A(n19469), .B(n19468), .Z(n19466) );
  XOR U27983 ( .A(y[5663]), .B(x[5663]), .Z(n19468) );
  XOR U27984 ( .A(y[5662]), .B(x[5662]), .Z(n19469) );
  XOR U27985 ( .A(y[5661]), .B(x[5661]), .Z(n19467) );
  XNOR U27986 ( .A(n19460), .B(n19459), .Z(n19461) );
  XNOR U27987 ( .A(n19456), .B(n19455), .Z(n19459) );
  XOR U27988 ( .A(n19458), .B(n19457), .Z(n19455) );
  XOR U27989 ( .A(y[5660]), .B(x[5660]), .Z(n19457) );
  XOR U27990 ( .A(y[5659]), .B(x[5659]), .Z(n19458) );
  XOR U27991 ( .A(y[5658]), .B(x[5658]), .Z(n19456) );
  XOR U27992 ( .A(n19450), .B(n19449), .Z(n19460) );
  XOR U27993 ( .A(n19452), .B(n19451), .Z(n19449) );
  XOR U27994 ( .A(y[5657]), .B(x[5657]), .Z(n19451) );
  XOR U27995 ( .A(y[5656]), .B(x[5656]), .Z(n19452) );
  XOR U27996 ( .A(y[5655]), .B(x[5655]), .Z(n19450) );
  NAND U27997 ( .A(n19513), .B(n19514), .Z(N63651) );
  NAND U27998 ( .A(n19515), .B(n19516), .Z(n19514) );
  NANDN U27999 ( .A(n19517), .B(n19518), .Z(n19516) );
  NANDN U28000 ( .A(n19518), .B(n19517), .Z(n19513) );
  XOR U28001 ( .A(n19517), .B(n19519), .Z(N63650) );
  XNOR U28002 ( .A(n19515), .B(n19518), .Z(n19519) );
  NAND U28003 ( .A(n19520), .B(n19521), .Z(n19518) );
  NAND U28004 ( .A(n19522), .B(n19523), .Z(n19521) );
  NANDN U28005 ( .A(n19524), .B(n19525), .Z(n19523) );
  NANDN U28006 ( .A(n19525), .B(n19524), .Z(n19520) );
  AND U28007 ( .A(n19526), .B(n19527), .Z(n19515) );
  NAND U28008 ( .A(n19528), .B(n19529), .Z(n19527) );
  NANDN U28009 ( .A(n19530), .B(n19531), .Z(n19529) );
  NANDN U28010 ( .A(n19531), .B(n19530), .Z(n19526) );
  IV U28011 ( .A(n19532), .Z(n19531) );
  AND U28012 ( .A(n19533), .B(n19534), .Z(n19517) );
  NAND U28013 ( .A(n19535), .B(n19536), .Z(n19534) );
  NANDN U28014 ( .A(n19537), .B(n19538), .Z(n19536) );
  NANDN U28015 ( .A(n19538), .B(n19537), .Z(n19533) );
  XOR U28016 ( .A(n19530), .B(n19539), .Z(N63649) );
  XNOR U28017 ( .A(n19528), .B(n19532), .Z(n19539) );
  XOR U28018 ( .A(n19525), .B(n19540), .Z(n19532) );
  XNOR U28019 ( .A(n19522), .B(n19524), .Z(n19540) );
  AND U28020 ( .A(n19541), .B(n19542), .Z(n19524) );
  NANDN U28021 ( .A(n19543), .B(n19544), .Z(n19542) );
  OR U28022 ( .A(n19545), .B(n19546), .Z(n19544) );
  IV U28023 ( .A(n19547), .Z(n19546) );
  NANDN U28024 ( .A(n19547), .B(n19545), .Z(n19541) );
  AND U28025 ( .A(n19548), .B(n19549), .Z(n19522) );
  NAND U28026 ( .A(n19550), .B(n19551), .Z(n19549) );
  NANDN U28027 ( .A(n19552), .B(n19553), .Z(n19551) );
  NANDN U28028 ( .A(n19553), .B(n19552), .Z(n19548) );
  IV U28029 ( .A(n19554), .Z(n19553) );
  NAND U28030 ( .A(n19555), .B(n19556), .Z(n19525) );
  NANDN U28031 ( .A(n19557), .B(n19558), .Z(n19556) );
  NANDN U28032 ( .A(n19559), .B(n19560), .Z(n19558) );
  NANDN U28033 ( .A(n19560), .B(n19559), .Z(n19555) );
  IV U28034 ( .A(n19561), .Z(n19559) );
  AND U28035 ( .A(n19562), .B(n19563), .Z(n19528) );
  NAND U28036 ( .A(n19564), .B(n19565), .Z(n19563) );
  NANDN U28037 ( .A(n19566), .B(n19567), .Z(n19565) );
  NANDN U28038 ( .A(n19567), .B(n19566), .Z(n19562) );
  XOR U28039 ( .A(n19538), .B(n19568), .Z(n19530) );
  XNOR U28040 ( .A(n19535), .B(n19537), .Z(n19568) );
  AND U28041 ( .A(n19569), .B(n19570), .Z(n19537) );
  NANDN U28042 ( .A(n19571), .B(n19572), .Z(n19570) );
  OR U28043 ( .A(n19573), .B(n19574), .Z(n19572) );
  IV U28044 ( .A(n19575), .Z(n19574) );
  NANDN U28045 ( .A(n19575), .B(n19573), .Z(n19569) );
  AND U28046 ( .A(n19576), .B(n19577), .Z(n19535) );
  NAND U28047 ( .A(n19578), .B(n19579), .Z(n19577) );
  NANDN U28048 ( .A(n19580), .B(n19581), .Z(n19579) );
  NANDN U28049 ( .A(n19581), .B(n19580), .Z(n19576) );
  IV U28050 ( .A(n19582), .Z(n19581) );
  NAND U28051 ( .A(n19583), .B(n19584), .Z(n19538) );
  NANDN U28052 ( .A(n19585), .B(n19586), .Z(n19584) );
  NANDN U28053 ( .A(n19587), .B(n19588), .Z(n19586) );
  NANDN U28054 ( .A(n19588), .B(n19587), .Z(n19583) );
  IV U28055 ( .A(n19589), .Z(n19587) );
  XOR U28056 ( .A(n19564), .B(n19590), .Z(N63648) );
  XNOR U28057 ( .A(n19567), .B(n19566), .Z(n19590) );
  XNOR U28058 ( .A(n19578), .B(n19591), .Z(n19566) );
  XNOR U28059 ( .A(n19582), .B(n19580), .Z(n19591) );
  XOR U28060 ( .A(n19588), .B(n19592), .Z(n19580) );
  XNOR U28061 ( .A(n19585), .B(n19589), .Z(n19592) );
  AND U28062 ( .A(n19593), .B(n19594), .Z(n19589) );
  NAND U28063 ( .A(n19595), .B(n19596), .Z(n19594) );
  NAND U28064 ( .A(n19597), .B(n19598), .Z(n19593) );
  AND U28065 ( .A(n19599), .B(n19600), .Z(n19585) );
  NAND U28066 ( .A(n19601), .B(n19602), .Z(n19600) );
  NAND U28067 ( .A(n19603), .B(n19604), .Z(n19599) );
  NANDN U28068 ( .A(n19605), .B(n19606), .Z(n19588) );
  ANDN U28069 ( .B(n19607), .A(n19608), .Z(n19582) );
  XNOR U28070 ( .A(n19573), .B(n19609), .Z(n19578) );
  XNOR U28071 ( .A(n19571), .B(n19575), .Z(n19609) );
  AND U28072 ( .A(n19610), .B(n19611), .Z(n19575) );
  NAND U28073 ( .A(n19612), .B(n19613), .Z(n19611) );
  NAND U28074 ( .A(n19614), .B(n19615), .Z(n19610) );
  AND U28075 ( .A(n19616), .B(n19617), .Z(n19571) );
  NAND U28076 ( .A(n19618), .B(n19619), .Z(n19617) );
  NAND U28077 ( .A(n19620), .B(n19621), .Z(n19616) );
  AND U28078 ( .A(n19622), .B(n19623), .Z(n19573) );
  NAND U28079 ( .A(n19624), .B(n19625), .Z(n19567) );
  XNOR U28080 ( .A(n19550), .B(n19626), .Z(n19564) );
  XNOR U28081 ( .A(n19554), .B(n19552), .Z(n19626) );
  XOR U28082 ( .A(n19560), .B(n19627), .Z(n19552) );
  XNOR U28083 ( .A(n19557), .B(n19561), .Z(n19627) );
  AND U28084 ( .A(n19628), .B(n19629), .Z(n19561) );
  NAND U28085 ( .A(n19630), .B(n19631), .Z(n19629) );
  NAND U28086 ( .A(n19632), .B(n19633), .Z(n19628) );
  AND U28087 ( .A(n19634), .B(n19635), .Z(n19557) );
  NAND U28088 ( .A(n19636), .B(n19637), .Z(n19635) );
  NAND U28089 ( .A(n19638), .B(n19639), .Z(n19634) );
  NANDN U28090 ( .A(n19640), .B(n19641), .Z(n19560) );
  ANDN U28091 ( .B(n19642), .A(n19643), .Z(n19554) );
  XNOR U28092 ( .A(n19545), .B(n19644), .Z(n19550) );
  XNOR U28093 ( .A(n19543), .B(n19547), .Z(n19644) );
  AND U28094 ( .A(n19645), .B(n19646), .Z(n19547) );
  NAND U28095 ( .A(n19647), .B(n19648), .Z(n19646) );
  NAND U28096 ( .A(n19649), .B(n19650), .Z(n19645) );
  AND U28097 ( .A(n19651), .B(n19652), .Z(n19543) );
  NAND U28098 ( .A(n19653), .B(n19654), .Z(n19652) );
  NAND U28099 ( .A(n19655), .B(n19656), .Z(n19651) );
  AND U28100 ( .A(n19657), .B(n19658), .Z(n19545) );
  XOR U28101 ( .A(n19625), .B(n19624), .Z(N63647) );
  XNOR U28102 ( .A(n19642), .B(n19643), .Z(n19624) );
  XNOR U28103 ( .A(n19657), .B(n19658), .Z(n19643) );
  XOR U28104 ( .A(n19654), .B(n19653), .Z(n19658) );
  XOR U28105 ( .A(y[5652]), .B(x[5652]), .Z(n19653) );
  XOR U28106 ( .A(n19656), .B(n19655), .Z(n19654) );
  XOR U28107 ( .A(y[5654]), .B(x[5654]), .Z(n19655) );
  XOR U28108 ( .A(y[5653]), .B(x[5653]), .Z(n19656) );
  XOR U28109 ( .A(n19648), .B(n19647), .Z(n19657) );
  XOR U28110 ( .A(n19650), .B(n19649), .Z(n19647) );
  XOR U28111 ( .A(y[5651]), .B(x[5651]), .Z(n19649) );
  XOR U28112 ( .A(y[5650]), .B(x[5650]), .Z(n19650) );
  XOR U28113 ( .A(y[5649]), .B(x[5649]), .Z(n19648) );
  XNOR U28114 ( .A(n19641), .B(n19640), .Z(n19642) );
  XNOR U28115 ( .A(n19637), .B(n19636), .Z(n19640) );
  XOR U28116 ( .A(n19639), .B(n19638), .Z(n19636) );
  XOR U28117 ( .A(y[5648]), .B(x[5648]), .Z(n19638) );
  XOR U28118 ( .A(y[5647]), .B(x[5647]), .Z(n19639) );
  XOR U28119 ( .A(y[5646]), .B(x[5646]), .Z(n19637) );
  XOR U28120 ( .A(n19631), .B(n19630), .Z(n19641) );
  XOR U28121 ( .A(n19633), .B(n19632), .Z(n19630) );
  XOR U28122 ( .A(y[5645]), .B(x[5645]), .Z(n19632) );
  XOR U28123 ( .A(y[5644]), .B(x[5644]), .Z(n19633) );
  XOR U28124 ( .A(y[5643]), .B(x[5643]), .Z(n19631) );
  XNOR U28125 ( .A(n19607), .B(n19608), .Z(n19625) );
  XNOR U28126 ( .A(n19622), .B(n19623), .Z(n19608) );
  XOR U28127 ( .A(n19619), .B(n19618), .Z(n19623) );
  XOR U28128 ( .A(y[5640]), .B(x[5640]), .Z(n19618) );
  XOR U28129 ( .A(n19621), .B(n19620), .Z(n19619) );
  XOR U28130 ( .A(y[5642]), .B(x[5642]), .Z(n19620) );
  XOR U28131 ( .A(y[5641]), .B(x[5641]), .Z(n19621) );
  XOR U28132 ( .A(n19613), .B(n19612), .Z(n19622) );
  XOR U28133 ( .A(n19615), .B(n19614), .Z(n19612) );
  XOR U28134 ( .A(y[5639]), .B(x[5639]), .Z(n19614) );
  XOR U28135 ( .A(y[5638]), .B(x[5638]), .Z(n19615) );
  XOR U28136 ( .A(y[5637]), .B(x[5637]), .Z(n19613) );
  XNOR U28137 ( .A(n19606), .B(n19605), .Z(n19607) );
  XNOR U28138 ( .A(n19602), .B(n19601), .Z(n19605) );
  XOR U28139 ( .A(n19604), .B(n19603), .Z(n19601) );
  XOR U28140 ( .A(y[5636]), .B(x[5636]), .Z(n19603) );
  XOR U28141 ( .A(y[5635]), .B(x[5635]), .Z(n19604) );
  XOR U28142 ( .A(y[5634]), .B(x[5634]), .Z(n19602) );
  XOR U28143 ( .A(n19596), .B(n19595), .Z(n19606) );
  XOR U28144 ( .A(n19598), .B(n19597), .Z(n19595) );
  XOR U28145 ( .A(y[5633]), .B(x[5633]), .Z(n19597) );
  XOR U28146 ( .A(y[5632]), .B(x[5632]), .Z(n19598) );
  XOR U28147 ( .A(y[5631]), .B(x[5631]), .Z(n19596) );
  NAND U28148 ( .A(n19659), .B(n19660), .Z(N63638) );
  NAND U28149 ( .A(n19661), .B(n19662), .Z(n19660) );
  NANDN U28150 ( .A(n19663), .B(n19664), .Z(n19662) );
  NANDN U28151 ( .A(n19664), .B(n19663), .Z(n19659) );
  XOR U28152 ( .A(n19663), .B(n19665), .Z(N63637) );
  XNOR U28153 ( .A(n19661), .B(n19664), .Z(n19665) );
  NAND U28154 ( .A(n19666), .B(n19667), .Z(n19664) );
  NAND U28155 ( .A(n19668), .B(n19669), .Z(n19667) );
  NANDN U28156 ( .A(n19670), .B(n19671), .Z(n19669) );
  NANDN U28157 ( .A(n19671), .B(n19670), .Z(n19666) );
  AND U28158 ( .A(n19672), .B(n19673), .Z(n19661) );
  NAND U28159 ( .A(n19674), .B(n19675), .Z(n19673) );
  NANDN U28160 ( .A(n19676), .B(n19677), .Z(n19675) );
  NANDN U28161 ( .A(n19677), .B(n19676), .Z(n19672) );
  IV U28162 ( .A(n19678), .Z(n19677) );
  AND U28163 ( .A(n19679), .B(n19680), .Z(n19663) );
  NAND U28164 ( .A(n19681), .B(n19682), .Z(n19680) );
  NANDN U28165 ( .A(n19683), .B(n19684), .Z(n19682) );
  NANDN U28166 ( .A(n19684), .B(n19683), .Z(n19679) );
  XOR U28167 ( .A(n19676), .B(n19685), .Z(N63636) );
  XNOR U28168 ( .A(n19674), .B(n19678), .Z(n19685) );
  XOR U28169 ( .A(n19671), .B(n19686), .Z(n19678) );
  XNOR U28170 ( .A(n19668), .B(n19670), .Z(n19686) );
  AND U28171 ( .A(n19687), .B(n19688), .Z(n19670) );
  NANDN U28172 ( .A(n19689), .B(n19690), .Z(n19688) );
  OR U28173 ( .A(n19691), .B(n19692), .Z(n19690) );
  IV U28174 ( .A(n19693), .Z(n19692) );
  NANDN U28175 ( .A(n19693), .B(n19691), .Z(n19687) );
  AND U28176 ( .A(n19694), .B(n19695), .Z(n19668) );
  NAND U28177 ( .A(n19696), .B(n19697), .Z(n19695) );
  NANDN U28178 ( .A(n19698), .B(n19699), .Z(n19697) );
  NANDN U28179 ( .A(n19699), .B(n19698), .Z(n19694) );
  IV U28180 ( .A(n19700), .Z(n19699) );
  NAND U28181 ( .A(n19701), .B(n19702), .Z(n19671) );
  NANDN U28182 ( .A(n19703), .B(n19704), .Z(n19702) );
  NANDN U28183 ( .A(n19705), .B(n19706), .Z(n19704) );
  NANDN U28184 ( .A(n19706), .B(n19705), .Z(n19701) );
  IV U28185 ( .A(n19707), .Z(n19705) );
  AND U28186 ( .A(n19708), .B(n19709), .Z(n19674) );
  NAND U28187 ( .A(n19710), .B(n19711), .Z(n19709) );
  NANDN U28188 ( .A(n19712), .B(n19713), .Z(n19711) );
  NANDN U28189 ( .A(n19713), .B(n19712), .Z(n19708) );
  XOR U28190 ( .A(n19684), .B(n19714), .Z(n19676) );
  XNOR U28191 ( .A(n19681), .B(n19683), .Z(n19714) );
  AND U28192 ( .A(n19715), .B(n19716), .Z(n19683) );
  NANDN U28193 ( .A(n19717), .B(n19718), .Z(n19716) );
  OR U28194 ( .A(n19719), .B(n19720), .Z(n19718) );
  IV U28195 ( .A(n19721), .Z(n19720) );
  NANDN U28196 ( .A(n19721), .B(n19719), .Z(n19715) );
  AND U28197 ( .A(n19722), .B(n19723), .Z(n19681) );
  NAND U28198 ( .A(n19724), .B(n19725), .Z(n19723) );
  NANDN U28199 ( .A(n19726), .B(n19727), .Z(n19725) );
  NANDN U28200 ( .A(n19727), .B(n19726), .Z(n19722) );
  IV U28201 ( .A(n19728), .Z(n19727) );
  NAND U28202 ( .A(n19729), .B(n19730), .Z(n19684) );
  NANDN U28203 ( .A(n19731), .B(n19732), .Z(n19730) );
  NANDN U28204 ( .A(n19733), .B(n19734), .Z(n19732) );
  NANDN U28205 ( .A(n19734), .B(n19733), .Z(n19729) );
  IV U28206 ( .A(n19735), .Z(n19733) );
  XOR U28207 ( .A(n19710), .B(n19736), .Z(N63635) );
  XNOR U28208 ( .A(n19713), .B(n19712), .Z(n19736) );
  XNOR U28209 ( .A(n19724), .B(n19737), .Z(n19712) );
  XNOR U28210 ( .A(n19728), .B(n19726), .Z(n19737) );
  XOR U28211 ( .A(n19734), .B(n19738), .Z(n19726) );
  XNOR U28212 ( .A(n19731), .B(n19735), .Z(n19738) );
  AND U28213 ( .A(n19739), .B(n19740), .Z(n19735) );
  NAND U28214 ( .A(n19741), .B(n19742), .Z(n19740) );
  NAND U28215 ( .A(n19743), .B(n19744), .Z(n19739) );
  AND U28216 ( .A(n19745), .B(n19746), .Z(n19731) );
  NAND U28217 ( .A(n19747), .B(n19748), .Z(n19746) );
  NAND U28218 ( .A(n19749), .B(n19750), .Z(n19745) );
  NANDN U28219 ( .A(n19751), .B(n19752), .Z(n19734) );
  ANDN U28220 ( .B(n19753), .A(n19754), .Z(n19728) );
  XNOR U28221 ( .A(n19719), .B(n19755), .Z(n19724) );
  XNOR U28222 ( .A(n19717), .B(n19721), .Z(n19755) );
  AND U28223 ( .A(n19756), .B(n19757), .Z(n19721) );
  NAND U28224 ( .A(n19758), .B(n19759), .Z(n19757) );
  NAND U28225 ( .A(n19760), .B(n19761), .Z(n19756) );
  AND U28226 ( .A(n19762), .B(n19763), .Z(n19717) );
  NAND U28227 ( .A(n19764), .B(n19765), .Z(n19763) );
  NAND U28228 ( .A(n19766), .B(n19767), .Z(n19762) );
  AND U28229 ( .A(n19768), .B(n19769), .Z(n19719) );
  NAND U28230 ( .A(n19770), .B(n19771), .Z(n19713) );
  XNOR U28231 ( .A(n19696), .B(n19772), .Z(n19710) );
  XNOR U28232 ( .A(n19700), .B(n19698), .Z(n19772) );
  XOR U28233 ( .A(n19706), .B(n19773), .Z(n19698) );
  XNOR U28234 ( .A(n19703), .B(n19707), .Z(n19773) );
  AND U28235 ( .A(n19774), .B(n19775), .Z(n19707) );
  NAND U28236 ( .A(n19776), .B(n19777), .Z(n19775) );
  NAND U28237 ( .A(n19778), .B(n19779), .Z(n19774) );
  AND U28238 ( .A(n19780), .B(n19781), .Z(n19703) );
  NAND U28239 ( .A(n19782), .B(n19783), .Z(n19781) );
  NAND U28240 ( .A(n19784), .B(n19785), .Z(n19780) );
  NANDN U28241 ( .A(n19786), .B(n19787), .Z(n19706) );
  ANDN U28242 ( .B(n19788), .A(n19789), .Z(n19700) );
  XNOR U28243 ( .A(n19691), .B(n19790), .Z(n19696) );
  XNOR U28244 ( .A(n19689), .B(n19693), .Z(n19790) );
  AND U28245 ( .A(n19791), .B(n19792), .Z(n19693) );
  NAND U28246 ( .A(n19793), .B(n19794), .Z(n19792) );
  NAND U28247 ( .A(n19795), .B(n19796), .Z(n19791) );
  AND U28248 ( .A(n19797), .B(n19798), .Z(n19689) );
  NAND U28249 ( .A(n19799), .B(n19800), .Z(n19798) );
  NAND U28250 ( .A(n19801), .B(n19802), .Z(n19797) );
  AND U28251 ( .A(n19803), .B(n19804), .Z(n19691) );
  XOR U28252 ( .A(n19771), .B(n19770), .Z(N63634) );
  XNOR U28253 ( .A(n19788), .B(n19789), .Z(n19770) );
  XNOR U28254 ( .A(n19803), .B(n19804), .Z(n19789) );
  XOR U28255 ( .A(n19800), .B(n19799), .Z(n19804) );
  XOR U28256 ( .A(y[5628]), .B(x[5628]), .Z(n19799) );
  XOR U28257 ( .A(n19802), .B(n19801), .Z(n19800) );
  XOR U28258 ( .A(y[5630]), .B(x[5630]), .Z(n19801) );
  XOR U28259 ( .A(y[5629]), .B(x[5629]), .Z(n19802) );
  XOR U28260 ( .A(n19794), .B(n19793), .Z(n19803) );
  XOR U28261 ( .A(n19796), .B(n19795), .Z(n19793) );
  XOR U28262 ( .A(y[5627]), .B(x[5627]), .Z(n19795) );
  XOR U28263 ( .A(y[5626]), .B(x[5626]), .Z(n19796) );
  XOR U28264 ( .A(y[5625]), .B(x[5625]), .Z(n19794) );
  XNOR U28265 ( .A(n19787), .B(n19786), .Z(n19788) );
  XNOR U28266 ( .A(n19783), .B(n19782), .Z(n19786) );
  XOR U28267 ( .A(n19785), .B(n19784), .Z(n19782) );
  XOR U28268 ( .A(y[5624]), .B(x[5624]), .Z(n19784) );
  XOR U28269 ( .A(y[5623]), .B(x[5623]), .Z(n19785) );
  XOR U28270 ( .A(y[5622]), .B(x[5622]), .Z(n19783) );
  XOR U28271 ( .A(n19777), .B(n19776), .Z(n19787) );
  XOR U28272 ( .A(n19779), .B(n19778), .Z(n19776) );
  XOR U28273 ( .A(y[5621]), .B(x[5621]), .Z(n19778) );
  XOR U28274 ( .A(y[5620]), .B(x[5620]), .Z(n19779) );
  XOR U28275 ( .A(y[5619]), .B(x[5619]), .Z(n19777) );
  XNOR U28276 ( .A(n19753), .B(n19754), .Z(n19771) );
  XNOR U28277 ( .A(n19768), .B(n19769), .Z(n19754) );
  XOR U28278 ( .A(n19765), .B(n19764), .Z(n19769) );
  XOR U28279 ( .A(y[5616]), .B(x[5616]), .Z(n19764) );
  XOR U28280 ( .A(n19767), .B(n19766), .Z(n19765) );
  XOR U28281 ( .A(y[5618]), .B(x[5618]), .Z(n19766) );
  XOR U28282 ( .A(y[5617]), .B(x[5617]), .Z(n19767) );
  XOR U28283 ( .A(n19759), .B(n19758), .Z(n19768) );
  XOR U28284 ( .A(n19761), .B(n19760), .Z(n19758) );
  XOR U28285 ( .A(y[5615]), .B(x[5615]), .Z(n19760) );
  XOR U28286 ( .A(y[5614]), .B(x[5614]), .Z(n19761) );
  XOR U28287 ( .A(y[5613]), .B(x[5613]), .Z(n19759) );
  XNOR U28288 ( .A(n19752), .B(n19751), .Z(n19753) );
  XNOR U28289 ( .A(n19748), .B(n19747), .Z(n19751) );
  XOR U28290 ( .A(n19750), .B(n19749), .Z(n19747) );
  XOR U28291 ( .A(y[5612]), .B(x[5612]), .Z(n19749) );
  XOR U28292 ( .A(y[5611]), .B(x[5611]), .Z(n19750) );
  XOR U28293 ( .A(y[5610]), .B(x[5610]), .Z(n19748) );
  XOR U28294 ( .A(n19742), .B(n19741), .Z(n19752) );
  XOR U28295 ( .A(n19744), .B(n19743), .Z(n19741) );
  XOR U28296 ( .A(y[5609]), .B(x[5609]), .Z(n19743) );
  XOR U28297 ( .A(y[5608]), .B(x[5608]), .Z(n19744) );
  XOR U28298 ( .A(y[5607]), .B(x[5607]), .Z(n19742) );
  NAND U28299 ( .A(n19805), .B(n19806), .Z(N63625) );
  NAND U28300 ( .A(n19807), .B(n19808), .Z(n19806) );
  NANDN U28301 ( .A(n19809), .B(n19810), .Z(n19808) );
  NANDN U28302 ( .A(n19810), .B(n19809), .Z(n19805) );
  XOR U28303 ( .A(n19809), .B(n19811), .Z(N63624) );
  XNOR U28304 ( .A(n19807), .B(n19810), .Z(n19811) );
  NAND U28305 ( .A(n19812), .B(n19813), .Z(n19810) );
  NAND U28306 ( .A(n19814), .B(n19815), .Z(n19813) );
  NANDN U28307 ( .A(n19816), .B(n19817), .Z(n19815) );
  NANDN U28308 ( .A(n19817), .B(n19816), .Z(n19812) );
  AND U28309 ( .A(n19818), .B(n19819), .Z(n19807) );
  NAND U28310 ( .A(n19820), .B(n19821), .Z(n19819) );
  NANDN U28311 ( .A(n19822), .B(n19823), .Z(n19821) );
  NANDN U28312 ( .A(n19823), .B(n19822), .Z(n19818) );
  IV U28313 ( .A(n19824), .Z(n19823) );
  AND U28314 ( .A(n19825), .B(n19826), .Z(n19809) );
  NAND U28315 ( .A(n19827), .B(n19828), .Z(n19826) );
  NANDN U28316 ( .A(n19829), .B(n19830), .Z(n19828) );
  NANDN U28317 ( .A(n19830), .B(n19829), .Z(n19825) );
  XOR U28318 ( .A(n19822), .B(n19831), .Z(N63623) );
  XNOR U28319 ( .A(n19820), .B(n19824), .Z(n19831) );
  XOR U28320 ( .A(n19817), .B(n19832), .Z(n19824) );
  XNOR U28321 ( .A(n19814), .B(n19816), .Z(n19832) );
  AND U28322 ( .A(n19833), .B(n19834), .Z(n19816) );
  NANDN U28323 ( .A(n19835), .B(n19836), .Z(n19834) );
  OR U28324 ( .A(n19837), .B(n19838), .Z(n19836) );
  IV U28325 ( .A(n19839), .Z(n19838) );
  NANDN U28326 ( .A(n19839), .B(n19837), .Z(n19833) );
  AND U28327 ( .A(n19840), .B(n19841), .Z(n19814) );
  NAND U28328 ( .A(n19842), .B(n19843), .Z(n19841) );
  NANDN U28329 ( .A(n19844), .B(n19845), .Z(n19843) );
  NANDN U28330 ( .A(n19845), .B(n19844), .Z(n19840) );
  IV U28331 ( .A(n19846), .Z(n19845) );
  NAND U28332 ( .A(n19847), .B(n19848), .Z(n19817) );
  NANDN U28333 ( .A(n19849), .B(n19850), .Z(n19848) );
  NANDN U28334 ( .A(n19851), .B(n19852), .Z(n19850) );
  NANDN U28335 ( .A(n19852), .B(n19851), .Z(n19847) );
  IV U28336 ( .A(n19853), .Z(n19851) );
  AND U28337 ( .A(n19854), .B(n19855), .Z(n19820) );
  NAND U28338 ( .A(n19856), .B(n19857), .Z(n19855) );
  NANDN U28339 ( .A(n19858), .B(n19859), .Z(n19857) );
  NANDN U28340 ( .A(n19859), .B(n19858), .Z(n19854) );
  XOR U28341 ( .A(n19830), .B(n19860), .Z(n19822) );
  XNOR U28342 ( .A(n19827), .B(n19829), .Z(n19860) );
  AND U28343 ( .A(n19861), .B(n19862), .Z(n19829) );
  NANDN U28344 ( .A(n19863), .B(n19864), .Z(n19862) );
  OR U28345 ( .A(n19865), .B(n19866), .Z(n19864) );
  IV U28346 ( .A(n19867), .Z(n19866) );
  NANDN U28347 ( .A(n19867), .B(n19865), .Z(n19861) );
  AND U28348 ( .A(n19868), .B(n19869), .Z(n19827) );
  NAND U28349 ( .A(n19870), .B(n19871), .Z(n19869) );
  NANDN U28350 ( .A(n19872), .B(n19873), .Z(n19871) );
  NANDN U28351 ( .A(n19873), .B(n19872), .Z(n19868) );
  IV U28352 ( .A(n19874), .Z(n19873) );
  NAND U28353 ( .A(n19875), .B(n19876), .Z(n19830) );
  NANDN U28354 ( .A(n19877), .B(n19878), .Z(n19876) );
  NANDN U28355 ( .A(n19879), .B(n19880), .Z(n19878) );
  NANDN U28356 ( .A(n19880), .B(n19879), .Z(n19875) );
  IV U28357 ( .A(n19881), .Z(n19879) );
  XOR U28358 ( .A(n19856), .B(n19882), .Z(N63622) );
  XNOR U28359 ( .A(n19859), .B(n19858), .Z(n19882) );
  XNOR U28360 ( .A(n19870), .B(n19883), .Z(n19858) );
  XNOR U28361 ( .A(n19874), .B(n19872), .Z(n19883) );
  XOR U28362 ( .A(n19880), .B(n19884), .Z(n19872) );
  XNOR U28363 ( .A(n19877), .B(n19881), .Z(n19884) );
  AND U28364 ( .A(n19885), .B(n19886), .Z(n19881) );
  NAND U28365 ( .A(n19887), .B(n19888), .Z(n19886) );
  NAND U28366 ( .A(n19889), .B(n19890), .Z(n19885) );
  AND U28367 ( .A(n19891), .B(n19892), .Z(n19877) );
  NAND U28368 ( .A(n19893), .B(n19894), .Z(n19892) );
  NAND U28369 ( .A(n19895), .B(n19896), .Z(n19891) );
  NANDN U28370 ( .A(n19897), .B(n19898), .Z(n19880) );
  ANDN U28371 ( .B(n19899), .A(n19900), .Z(n19874) );
  XNOR U28372 ( .A(n19865), .B(n19901), .Z(n19870) );
  XNOR U28373 ( .A(n19863), .B(n19867), .Z(n19901) );
  AND U28374 ( .A(n19902), .B(n19903), .Z(n19867) );
  NAND U28375 ( .A(n19904), .B(n19905), .Z(n19903) );
  NAND U28376 ( .A(n19906), .B(n19907), .Z(n19902) );
  AND U28377 ( .A(n19908), .B(n19909), .Z(n19863) );
  NAND U28378 ( .A(n19910), .B(n19911), .Z(n19909) );
  NAND U28379 ( .A(n19912), .B(n19913), .Z(n19908) );
  AND U28380 ( .A(n19914), .B(n19915), .Z(n19865) );
  NAND U28381 ( .A(n19916), .B(n19917), .Z(n19859) );
  XNOR U28382 ( .A(n19842), .B(n19918), .Z(n19856) );
  XNOR U28383 ( .A(n19846), .B(n19844), .Z(n19918) );
  XOR U28384 ( .A(n19852), .B(n19919), .Z(n19844) );
  XNOR U28385 ( .A(n19849), .B(n19853), .Z(n19919) );
  AND U28386 ( .A(n19920), .B(n19921), .Z(n19853) );
  NAND U28387 ( .A(n19922), .B(n19923), .Z(n19921) );
  NAND U28388 ( .A(n19924), .B(n19925), .Z(n19920) );
  AND U28389 ( .A(n19926), .B(n19927), .Z(n19849) );
  NAND U28390 ( .A(n19928), .B(n19929), .Z(n19927) );
  NAND U28391 ( .A(n19930), .B(n19931), .Z(n19926) );
  NANDN U28392 ( .A(n19932), .B(n19933), .Z(n19852) );
  ANDN U28393 ( .B(n19934), .A(n19935), .Z(n19846) );
  XNOR U28394 ( .A(n19837), .B(n19936), .Z(n19842) );
  XNOR U28395 ( .A(n19835), .B(n19839), .Z(n19936) );
  AND U28396 ( .A(n19937), .B(n19938), .Z(n19839) );
  NAND U28397 ( .A(n19939), .B(n19940), .Z(n19938) );
  NAND U28398 ( .A(n19941), .B(n19942), .Z(n19937) );
  AND U28399 ( .A(n19943), .B(n19944), .Z(n19835) );
  NAND U28400 ( .A(n19945), .B(n19946), .Z(n19944) );
  NAND U28401 ( .A(n19947), .B(n19948), .Z(n19943) );
  AND U28402 ( .A(n19949), .B(n19950), .Z(n19837) );
  XOR U28403 ( .A(n19917), .B(n19916), .Z(N63621) );
  XNOR U28404 ( .A(n19934), .B(n19935), .Z(n19916) );
  XNOR U28405 ( .A(n19949), .B(n19950), .Z(n19935) );
  XOR U28406 ( .A(n19946), .B(n19945), .Z(n19950) );
  XOR U28407 ( .A(y[5604]), .B(x[5604]), .Z(n19945) );
  XOR U28408 ( .A(n19948), .B(n19947), .Z(n19946) );
  XOR U28409 ( .A(y[5606]), .B(x[5606]), .Z(n19947) );
  XOR U28410 ( .A(y[5605]), .B(x[5605]), .Z(n19948) );
  XOR U28411 ( .A(n19940), .B(n19939), .Z(n19949) );
  XOR U28412 ( .A(n19942), .B(n19941), .Z(n19939) );
  XOR U28413 ( .A(y[5603]), .B(x[5603]), .Z(n19941) );
  XOR U28414 ( .A(y[5602]), .B(x[5602]), .Z(n19942) );
  XOR U28415 ( .A(y[5601]), .B(x[5601]), .Z(n19940) );
  XNOR U28416 ( .A(n19933), .B(n19932), .Z(n19934) );
  XNOR U28417 ( .A(n19929), .B(n19928), .Z(n19932) );
  XOR U28418 ( .A(n19931), .B(n19930), .Z(n19928) );
  XOR U28419 ( .A(y[5600]), .B(x[5600]), .Z(n19930) );
  XOR U28420 ( .A(y[5599]), .B(x[5599]), .Z(n19931) );
  XOR U28421 ( .A(y[5598]), .B(x[5598]), .Z(n19929) );
  XOR U28422 ( .A(n19923), .B(n19922), .Z(n19933) );
  XOR U28423 ( .A(n19925), .B(n19924), .Z(n19922) );
  XOR U28424 ( .A(y[5597]), .B(x[5597]), .Z(n19924) );
  XOR U28425 ( .A(y[5596]), .B(x[5596]), .Z(n19925) );
  XOR U28426 ( .A(y[5595]), .B(x[5595]), .Z(n19923) );
  XNOR U28427 ( .A(n19899), .B(n19900), .Z(n19917) );
  XNOR U28428 ( .A(n19914), .B(n19915), .Z(n19900) );
  XOR U28429 ( .A(n19911), .B(n19910), .Z(n19915) );
  XOR U28430 ( .A(y[5592]), .B(x[5592]), .Z(n19910) );
  XOR U28431 ( .A(n19913), .B(n19912), .Z(n19911) );
  XOR U28432 ( .A(y[5594]), .B(x[5594]), .Z(n19912) );
  XOR U28433 ( .A(y[5593]), .B(x[5593]), .Z(n19913) );
  XOR U28434 ( .A(n19905), .B(n19904), .Z(n19914) );
  XOR U28435 ( .A(n19907), .B(n19906), .Z(n19904) );
  XOR U28436 ( .A(y[5591]), .B(x[5591]), .Z(n19906) );
  XOR U28437 ( .A(y[5590]), .B(x[5590]), .Z(n19907) );
  XOR U28438 ( .A(y[5589]), .B(x[5589]), .Z(n19905) );
  XNOR U28439 ( .A(n19898), .B(n19897), .Z(n19899) );
  XNOR U28440 ( .A(n19894), .B(n19893), .Z(n19897) );
  XOR U28441 ( .A(n19896), .B(n19895), .Z(n19893) );
  XOR U28442 ( .A(y[5588]), .B(x[5588]), .Z(n19895) );
  XOR U28443 ( .A(y[5587]), .B(x[5587]), .Z(n19896) );
  XOR U28444 ( .A(y[5586]), .B(x[5586]), .Z(n19894) );
  XOR U28445 ( .A(n19888), .B(n19887), .Z(n19898) );
  XOR U28446 ( .A(n19890), .B(n19889), .Z(n19887) );
  XOR U28447 ( .A(y[5585]), .B(x[5585]), .Z(n19889) );
  XOR U28448 ( .A(y[5584]), .B(x[5584]), .Z(n19890) );
  XOR U28449 ( .A(y[5583]), .B(x[5583]), .Z(n19888) );
  NAND U28450 ( .A(n19951), .B(n19952), .Z(N63612) );
  NAND U28451 ( .A(n19953), .B(n19954), .Z(n19952) );
  NANDN U28452 ( .A(n19955), .B(n19956), .Z(n19954) );
  NANDN U28453 ( .A(n19956), .B(n19955), .Z(n19951) );
  XOR U28454 ( .A(n19955), .B(n19957), .Z(N63611) );
  XNOR U28455 ( .A(n19953), .B(n19956), .Z(n19957) );
  NAND U28456 ( .A(n19958), .B(n19959), .Z(n19956) );
  NAND U28457 ( .A(n19960), .B(n19961), .Z(n19959) );
  NANDN U28458 ( .A(n19962), .B(n19963), .Z(n19961) );
  NANDN U28459 ( .A(n19963), .B(n19962), .Z(n19958) );
  AND U28460 ( .A(n19964), .B(n19965), .Z(n19953) );
  NAND U28461 ( .A(n19966), .B(n19967), .Z(n19965) );
  NANDN U28462 ( .A(n19968), .B(n19969), .Z(n19967) );
  NANDN U28463 ( .A(n19969), .B(n19968), .Z(n19964) );
  IV U28464 ( .A(n19970), .Z(n19969) );
  AND U28465 ( .A(n19971), .B(n19972), .Z(n19955) );
  NAND U28466 ( .A(n19973), .B(n19974), .Z(n19972) );
  NANDN U28467 ( .A(n19975), .B(n19976), .Z(n19974) );
  NANDN U28468 ( .A(n19976), .B(n19975), .Z(n19971) );
  XOR U28469 ( .A(n19968), .B(n19977), .Z(N63610) );
  XNOR U28470 ( .A(n19966), .B(n19970), .Z(n19977) );
  XOR U28471 ( .A(n19963), .B(n19978), .Z(n19970) );
  XNOR U28472 ( .A(n19960), .B(n19962), .Z(n19978) );
  AND U28473 ( .A(n19979), .B(n19980), .Z(n19962) );
  NANDN U28474 ( .A(n19981), .B(n19982), .Z(n19980) );
  OR U28475 ( .A(n19983), .B(n19984), .Z(n19982) );
  IV U28476 ( .A(n19985), .Z(n19984) );
  NANDN U28477 ( .A(n19985), .B(n19983), .Z(n19979) );
  AND U28478 ( .A(n19986), .B(n19987), .Z(n19960) );
  NAND U28479 ( .A(n19988), .B(n19989), .Z(n19987) );
  NANDN U28480 ( .A(n19990), .B(n19991), .Z(n19989) );
  NANDN U28481 ( .A(n19991), .B(n19990), .Z(n19986) );
  IV U28482 ( .A(n19992), .Z(n19991) );
  NAND U28483 ( .A(n19993), .B(n19994), .Z(n19963) );
  NANDN U28484 ( .A(n19995), .B(n19996), .Z(n19994) );
  NANDN U28485 ( .A(n19997), .B(n19998), .Z(n19996) );
  NANDN U28486 ( .A(n19998), .B(n19997), .Z(n19993) );
  IV U28487 ( .A(n19999), .Z(n19997) );
  AND U28488 ( .A(n20000), .B(n20001), .Z(n19966) );
  NAND U28489 ( .A(n20002), .B(n20003), .Z(n20001) );
  NANDN U28490 ( .A(n20004), .B(n20005), .Z(n20003) );
  NANDN U28491 ( .A(n20005), .B(n20004), .Z(n20000) );
  XOR U28492 ( .A(n19976), .B(n20006), .Z(n19968) );
  XNOR U28493 ( .A(n19973), .B(n19975), .Z(n20006) );
  AND U28494 ( .A(n20007), .B(n20008), .Z(n19975) );
  NANDN U28495 ( .A(n20009), .B(n20010), .Z(n20008) );
  OR U28496 ( .A(n20011), .B(n20012), .Z(n20010) );
  IV U28497 ( .A(n20013), .Z(n20012) );
  NANDN U28498 ( .A(n20013), .B(n20011), .Z(n20007) );
  AND U28499 ( .A(n20014), .B(n20015), .Z(n19973) );
  NAND U28500 ( .A(n20016), .B(n20017), .Z(n20015) );
  NANDN U28501 ( .A(n20018), .B(n20019), .Z(n20017) );
  NANDN U28502 ( .A(n20019), .B(n20018), .Z(n20014) );
  IV U28503 ( .A(n20020), .Z(n20019) );
  NAND U28504 ( .A(n20021), .B(n20022), .Z(n19976) );
  NANDN U28505 ( .A(n20023), .B(n20024), .Z(n20022) );
  NANDN U28506 ( .A(n20025), .B(n20026), .Z(n20024) );
  NANDN U28507 ( .A(n20026), .B(n20025), .Z(n20021) );
  IV U28508 ( .A(n20027), .Z(n20025) );
  XOR U28509 ( .A(n20002), .B(n20028), .Z(N63609) );
  XNOR U28510 ( .A(n20005), .B(n20004), .Z(n20028) );
  XNOR U28511 ( .A(n20016), .B(n20029), .Z(n20004) );
  XNOR U28512 ( .A(n20020), .B(n20018), .Z(n20029) );
  XOR U28513 ( .A(n20026), .B(n20030), .Z(n20018) );
  XNOR U28514 ( .A(n20023), .B(n20027), .Z(n20030) );
  AND U28515 ( .A(n20031), .B(n20032), .Z(n20027) );
  NAND U28516 ( .A(n20033), .B(n20034), .Z(n20032) );
  NAND U28517 ( .A(n20035), .B(n20036), .Z(n20031) );
  AND U28518 ( .A(n20037), .B(n20038), .Z(n20023) );
  NAND U28519 ( .A(n20039), .B(n20040), .Z(n20038) );
  NAND U28520 ( .A(n20041), .B(n20042), .Z(n20037) );
  NANDN U28521 ( .A(n20043), .B(n20044), .Z(n20026) );
  ANDN U28522 ( .B(n20045), .A(n20046), .Z(n20020) );
  XNOR U28523 ( .A(n20011), .B(n20047), .Z(n20016) );
  XNOR U28524 ( .A(n20009), .B(n20013), .Z(n20047) );
  AND U28525 ( .A(n20048), .B(n20049), .Z(n20013) );
  NAND U28526 ( .A(n20050), .B(n20051), .Z(n20049) );
  NAND U28527 ( .A(n20052), .B(n20053), .Z(n20048) );
  AND U28528 ( .A(n20054), .B(n20055), .Z(n20009) );
  NAND U28529 ( .A(n20056), .B(n20057), .Z(n20055) );
  NAND U28530 ( .A(n20058), .B(n20059), .Z(n20054) );
  AND U28531 ( .A(n20060), .B(n20061), .Z(n20011) );
  NAND U28532 ( .A(n20062), .B(n20063), .Z(n20005) );
  XNOR U28533 ( .A(n19988), .B(n20064), .Z(n20002) );
  XNOR U28534 ( .A(n19992), .B(n19990), .Z(n20064) );
  XOR U28535 ( .A(n19998), .B(n20065), .Z(n19990) );
  XNOR U28536 ( .A(n19995), .B(n19999), .Z(n20065) );
  AND U28537 ( .A(n20066), .B(n20067), .Z(n19999) );
  NAND U28538 ( .A(n20068), .B(n20069), .Z(n20067) );
  NAND U28539 ( .A(n20070), .B(n20071), .Z(n20066) );
  AND U28540 ( .A(n20072), .B(n20073), .Z(n19995) );
  NAND U28541 ( .A(n20074), .B(n20075), .Z(n20073) );
  NAND U28542 ( .A(n20076), .B(n20077), .Z(n20072) );
  NANDN U28543 ( .A(n20078), .B(n20079), .Z(n19998) );
  ANDN U28544 ( .B(n20080), .A(n20081), .Z(n19992) );
  XNOR U28545 ( .A(n19983), .B(n20082), .Z(n19988) );
  XNOR U28546 ( .A(n19981), .B(n19985), .Z(n20082) );
  AND U28547 ( .A(n20083), .B(n20084), .Z(n19985) );
  NAND U28548 ( .A(n20085), .B(n20086), .Z(n20084) );
  NAND U28549 ( .A(n20087), .B(n20088), .Z(n20083) );
  AND U28550 ( .A(n20089), .B(n20090), .Z(n19981) );
  NAND U28551 ( .A(n20091), .B(n20092), .Z(n20090) );
  NAND U28552 ( .A(n20093), .B(n20094), .Z(n20089) );
  AND U28553 ( .A(n20095), .B(n20096), .Z(n19983) );
  XOR U28554 ( .A(n20063), .B(n20062), .Z(N63608) );
  XNOR U28555 ( .A(n20080), .B(n20081), .Z(n20062) );
  XNOR U28556 ( .A(n20095), .B(n20096), .Z(n20081) );
  XOR U28557 ( .A(n20092), .B(n20091), .Z(n20096) );
  XOR U28558 ( .A(y[5580]), .B(x[5580]), .Z(n20091) );
  XOR U28559 ( .A(n20094), .B(n20093), .Z(n20092) );
  XOR U28560 ( .A(y[5582]), .B(x[5582]), .Z(n20093) );
  XOR U28561 ( .A(y[5581]), .B(x[5581]), .Z(n20094) );
  XOR U28562 ( .A(n20086), .B(n20085), .Z(n20095) );
  XOR U28563 ( .A(n20088), .B(n20087), .Z(n20085) );
  XOR U28564 ( .A(y[5579]), .B(x[5579]), .Z(n20087) );
  XOR U28565 ( .A(y[5578]), .B(x[5578]), .Z(n20088) );
  XOR U28566 ( .A(y[5577]), .B(x[5577]), .Z(n20086) );
  XNOR U28567 ( .A(n20079), .B(n20078), .Z(n20080) );
  XNOR U28568 ( .A(n20075), .B(n20074), .Z(n20078) );
  XOR U28569 ( .A(n20077), .B(n20076), .Z(n20074) );
  XOR U28570 ( .A(y[5576]), .B(x[5576]), .Z(n20076) );
  XOR U28571 ( .A(y[5575]), .B(x[5575]), .Z(n20077) );
  XOR U28572 ( .A(y[5574]), .B(x[5574]), .Z(n20075) );
  XOR U28573 ( .A(n20069), .B(n20068), .Z(n20079) );
  XOR U28574 ( .A(n20071), .B(n20070), .Z(n20068) );
  XOR U28575 ( .A(y[5573]), .B(x[5573]), .Z(n20070) );
  XOR U28576 ( .A(y[5572]), .B(x[5572]), .Z(n20071) );
  XOR U28577 ( .A(y[5571]), .B(x[5571]), .Z(n20069) );
  XNOR U28578 ( .A(n20045), .B(n20046), .Z(n20063) );
  XNOR U28579 ( .A(n20060), .B(n20061), .Z(n20046) );
  XOR U28580 ( .A(n20057), .B(n20056), .Z(n20061) );
  XOR U28581 ( .A(y[5568]), .B(x[5568]), .Z(n20056) );
  XOR U28582 ( .A(n20059), .B(n20058), .Z(n20057) );
  XOR U28583 ( .A(y[5570]), .B(x[5570]), .Z(n20058) );
  XOR U28584 ( .A(y[5569]), .B(x[5569]), .Z(n20059) );
  XOR U28585 ( .A(n20051), .B(n20050), .Z(n20060) );
  XOR U28586 ( .A(n20053), .B(n20052), .Z(n20050) );
  XOR U28587 ( .A(y[5567]), .B(x[5567]), .Z(n20052) );
  XOR U28588 ( .A(y[5566]), .B(x[5566]), .Z(n20053) );
  XOR U28589 ( .A(y[5565]), .B(x[5565]), .Z(n20051) );
  XNOR U28590 ( .A(n20044), .B(n20043), .Z(n20045) );
  XNOR U28591 ( .A(n20040), .B(n20039), .Z(n20043) );
  XOR U28592 ( .A(n20042), .B(n20041), .Z(n20039) );
  XOR U28593 ( .A(y[5564]), .B(x[5564]), .Z(n20041) );
  XOR U28594 ( .A(y[5563]), .B(x[5563]), .Z(n20042) );
  XOR U28595 ( .A(y[5562]), .B(x[5562]), .Z(n20040) );
  XOR U28596 ( .A(n20034), .B(n20033), .Z(n20044) );
  XOR U28597 ( .A(n20036), .B(n20035), .Z(n20033) );
  XOR U28598 ( .A(y[5561]), .B(x[5561]), .Z(n20035) );
  XOR U28599 ( .A(y[5560]), .B(x[5560]), .Z(n20036) );
  XOR U28600 ( .A(y[5559]), .B(x[5559]), .Z(n20034) );
  NAND U28601 ( .A(n20097), .B(n20098), .Z(N63599) );
  NAND U28602 ( .A(n20099), .B(n20100), .Z(n20098) );
  NANDN U28603 ( .A(n20101), .B(n20102), .Z(n20100) );
  NANDN U28604 ( .A(n20102), .B(n20101), .Z(n20097) );
  XOR U28605 ( .A(n20101), .B(n20103), .Z(N63598) );
  XNOR U28606 ( .A(n20099), .B(n20102), .Z(n20103) );
  NAND U28607 ( .A(n20104), .B(n20105), .Z(n20102) );
  NAND U28608 ( .A(n20106), .B(n20107), .Z(n20105) );
  NANDN U28609 ( .A(n20108), .B(n20109), .Z(n20107) );
  NANDN U28610 ( .A(n20109), .B(n20108), .Z(n20104) );
  AND U28611 ( .A(n20110), .B(n20111), .Z(n20099) );
  NAND U28612 ( .A(n20112), .B(n20113), .Z(n20111) );
  NANDN U28613 ( .A(n20114), .B(n20115), .Z(n20113) );
  NANDN U28614 ( .A(n20115), .B(n20114), .Z(n20110) );
  IV U28615 ( .A(n20116), .Z(n20115) );
  AND U28616 ( .A(n20117), .B(n20118), .Z(n20101) );
  NAND U28617 ( .A(n20119), .B(n20120), .Z(n20118) );
  NANDN U28618 ( .A(n20121), .B(n20122), .Z(n20120) );
  NANDN U28619 ( .A(n20122), .B(n20121), .Z(n20117) );
  XOR U28620 ( .A(n20114), .B(n20123), .Z(N63597) );
  XNOR U28621 ( .A(n20112), .B(n20116), .Z(n20123) );
  XOR U28622 ( .A(n20109), .B(n20124), .Z(n20116) );
  XNOR U28623 ( .A(n20106), .B(n20108), .Z(n20124) );
  AND U28624 ( .A(n20125), .B(n20126), .Z(n20108) );
  NANDN U28625 ( .A(n20127), .B(n20128), .Z(n20126) );
  OR U28626 ( .A(n20129), .B(n20130), .Z(n20128) );
  IV U28627 ( .A(n20131), .Z(n20130) );
  NANDN U28628 ( .A(n20131), .B(n20129), .Z(n20125) );
  AND U28629 ( .A(n20132), .B(n20133), .Z(n20106) );
  NAND U28630 ( .A(n20134), .B(n20135), .Z(n20133) );
  NANDN U28631 ( .A(n20136), .B(n20137), .Z(n20135) );
  NANDN U28632 ( .A(n20137), .B(n20136), .Z(n20132) );
  IV U28633 ( .A(n20138), .Z(n20137) );
  NAND U28634 ( .A(n20139), .B(n20140), .Z(n20109) );
  NANDN U28635 ( .A(n20141), .B(n20142), .Z(n20140) );
  NANDN U28636 ( .A(n20143), .B(n20144), .Z(n20142) );
  NANDN U28637 ( .A(n20144), .B(n20143), .Z(n20139) );
  IV U28638 ( .A(n20145), .Z(n20143) );
  AND U28639 ( .A(n20146), .B(n20147), .Z(n20112) );
  NAND U28640 ( .A(n20148), .B(n20149), .Z(n20147) );
  NANDN U28641 ( .A(n20150), .B(n20151), .Z(n20149) );
  NANDN U28642 ( .A(n20151), .B(n20150), .Z(n20146) );
  XOR U28643 ( .A(n20122), .B(n20152), .Z(n20114) );
  XNOR U28644 ( .A(n20119), .B(n20121), .Z(n20152) );
  AND U28645 ( .A(n20153), .B(n20154), .Z(n20121) );
  NANDN U28646 ( .A(n20155), .B(n20156), .Z(n20154) );
  OR U28647 ( .A(n20157), .B(n20158), .Z(n20156) );
  IV U28648 ( .A(n20159), .Z(n20158) );
  NANDN U28649 ( .A(n20159), .B(n20157), .Z(n20153) );
  AND U28650 ( .A(n20160), .B(n20161), .Z(n20119) );
  NAND U28651 ( .A(n20162), .B(n20163), .Z(n20161) );
  NANDN U28652 ( .A(n20164), .B(n20165), .Z(n20163) );
  NANDN U28653 ( .A(n20165), .B(n20164), .Z(n20160) );
  IV U28654 ( .A(n20166), .Z(n20165) );
  NAND U28655 ( .A(n20167), .B(n20168), .Z(n20122) );
  NANDN U28656 ( .A(n20169), .B(n20170), .Z(n20168) );
  NANDN U28657 ( .A(n20171), .B(n20172), .Z(n20170) );
  NANDN U28658 ( .A(n20172), .B(n20171), .Z(n20167) );
  IV U28659 ( .A(n20173), .Z(n20171) );
  XOR U28660 ( .A(n20148), .B(n20174), .Z(N63596) );
  XNOR U28661 ( .A(n20151), .B(n20150), .Z(n20174) );
  XNOR U28662 ( .A(n20162), .B(n20175), .Z(n20150) );
  XNOR U28663 ( .A(n20166), .B(n20164), .Z(n20175) );
  XOR U28664 ( .A(n20172), .B(n20176), .Z(n20164) );
  XNOR U28665 ( .A(n20169), .B(n20173), .Z(n20176) );
  AND U28666 ( .A(n20177), .B(n20178), .Z(n20173) );
  NAND U28667 ( .A(n20179), .B(n20180), .Z(n20178) );
  NAND U28668 ( .A(n20181), .B(n20182), .Z(n20177) );
  AND U28669 ( .A(n20183), .B(n20184), .Z(n20169) );
  NAND U28670 ( .A(n20185), .B(n20186), .Z(n20184) );
  NAND U28671 ( .A(n20187), .B(n20188), .Z(n20183) );
  NANDN U28672 ( .A(n20189), .B(n20190), .Z(n20172) );
  ANDN U28673 ( .B(n20191), .A(n20192), .Z(n20166) );
  XNOR U28674 ( .A(n20157), .B(n20193), .Z(n20162) );
  XNOR U28675 ( .A(n20155), .B(n20159), .Z(n20193) );
  AND U28676 ( .A(n20194), .B(n20195), .Z(n20159) );
  NAND U28677 ( .A(n20196), .B(n20197), .Z(n20195) );
  NAND U28678 ( .A(n20198), .B(n20199), .Z(n20194) );
  AND U28679 ( .A(n20200), .B(n20201), .Z(n20155) );
  NAND U28680 ( .A(n20202), .B(n20203), .Z(n20201) );
  NAND U28681 ( .A(n20204), .B(n20205), .Z(n20200) );
  AND U28682 ( .A(n20206), .B(n20207), .Z(n20157) );
  NAND U28683 ( .A(n20208), .B(n20209), .Z(n20151) );
  XNOR U28684 ( .A(n20134), .B(n20210), .Z(n20148) );
  XNOR U28685 ( .A(n20138), .B(n20136), .Z(n20210) );
  XOR U28686 ( .A(n20144), .B(n20211), .Z(n20136) );
  XNOR U28687 ( .A(n20141), .B(n20145), .Z(n20211) );
  AND U28688 ( .A(n20212), .B(n20213), .Z(n20145) );
  NAND U28689 ( .A(n20214), .B(n20215), .Z(n20213) );
  NAND U28690 ( .A(n20216), .B(n20217), .Z(n20212) );
  AND U28691 ( .A(n20218), .B(n20219), .Z(n20141) );
  NAND U28692 ( .A(n20220), .B(n20221), .Z(n20219) );
  NAND U28693 ( .A(n20222), .B(n20223), .Z(n20218) );
  NANDN U28694 ( .A(n20224), .B(n20225), .Z(n20144) );
  ANDN U28695 ( .B(n20226), .A(n20227), .Z(n20138) );
  XNOR U28696 ( .A(n20129), .B(n20228), .Z(n20134) );
  XNOR U28697 ( .A(n20127), .B(n20131), .Z(n20228) );
  AND U28698 ( .A(n20229), .B(n20230), .Z(n20131) );
  NAND U28699 ( .A(n20231), .B(n20232), .Z(n20230) );
  NAND U28700 ( .A(n20233), .B(n20234), .Z(n20229) );
  AND U28701 ( .A(n20235), .B(n20236), .Z(n20127) );
  NAND U28702 ( .A(n20237), .B(n20238), .Z(n20236) );
  NAND U28703 ( .A(n20239), .B(n20240), .Z(n20235) );
  AND U28704 ( .A(n20241), .B(n20242), .Z(n20129) );
  XOR U28705 ( .A(n20209), .B(n20208), .Z(N63595) );
  XNOR U28706 ( .A(n20226), .B(n20227), .Z(n20208) );
  XNOR U28707 ( .A(n20241), .B(n20242), .Z(n20227) );
  XOR U28708 ( .A(n20238), .B(n20237), .Z(n20242) );
  XOR U28709 ( .A(y[5556]), .B(x[5556]), .Z(n20237) );
  XOR U28710 ( .A(n20240), .B(n20239), .Z(n20238) );
  XOR U28711 ( .A(y[5558]), .B(x[5558]), .Z(n20239) );
  XOR U28712 ( .A(y[5557]), .B(x[5557]), .Z(n20240) );
  XOR U28713 ( .A(n20232), .B(n20231), .Z(n20241) );
  XOR U28714 ( .A(n20234), .B(n20233), .Z(n20231) );
  XOR U28715 ( .A(y[5555]), .B(x[5555]), .Z(n20233) );
  XOR U28716 ( .A(y[5554]), .B(x[5554]), .Z(n20234) );
  XOR U28717 ( .A(y[5553]), .B(x[5553]), .Z(n20232) );
  XNOR U28718 ( .A(n20225), .B(n20224), .Z(n20226) );
  XNOR U28719 ( .A(n20221), .B(n20220), .Z(n20224) );
  XOR U28720 ( .A(n20223), .B(n20222), .Z(n20220) );
  XOR U28721 ( .A(y[5552]), .B(x[5552]), .Z(n20222) );
  XOR U28722 ( .A(y[5551]), .B(x[5551]), .Z(n20223) );
  XOR U28723 ( .A(y[5550]), .B(x[5550]), .Z(n20221) );
  XOR U28724 ( .A(n20215), .B(n20214), .Z(n20225) );
  XOR U28725 ( .A(n20217), .B(n20216), .Z(n20214) );
  XOR U28726 ( .A(y[5549]), .B(x[5549]), .Z(n20216) );
  XOR U28727 ( .A(y[5548]), .B(x[5548]), .Z(n20217) );
  XOR U28728 ( .A(y[5547]), .B(x[5547]), .Z(n20215) );
  XNOR U28729 ( .A(n20191), .B(n20192), .Z(n20209) );
  XNOR U28730 ( .A(n20206), .B(n20207), .Z(n20192) );
  XOR U28731 ( .A(n20203), .B(n20202), .Z(n20207) );
  XOR U28732 ( .A(y[5544]), .B(x[5544]), .Z(n20202) );
  XOR U28733 ( .A(n20205), .B(n20204), .Z(n20203) );
  XOR U28734 ( .A(y[5546]), .B(x[5546]), .Z(n20204) );
  XOR U28735 ( .A(y[5545]), .B(x[5545]), .Z(n20205) );
  XOR U28736 ( .A(n20197), .B(n20196), .Z(n20206) );
  XOR U28737 ( .A(n20199), .B(n20198), .Z(n20196) );
  XOR U28738 ( .A(y[5543]), .B(x[5543]), .Z(n20198) );
  XOR U28739 ( .A(y[5542]), .B(x[5542]), .Z(n20199) );
  XOR U28740 ( .A(y[5541]), .B(x[5541]), .Z(n20197) );
  XNOR U28741 ( .A(n20190), .B(n20189), .Z(n20191) );
  XNOR U28742 ( .A(n20186), .B(n20185), .Z(n20189) );
  XOR U28743 ( .A(n20188), .B(n20187), .Z(n20185) );
  XOR U28744 ( .A(y[5540]), .B(x[5540]), .Z(n20187) );
  XOR U28745 ( .A(y[5539]), .B(x[5539]), .Z(n20188) );
  XOR U28746 ( .A(y[5538]), .B(x[5538]), .Z(n20186) );
  XOR U28747 ( .A(n20180), .B(n20179), .Z(n20190) );
  XOR U28748 ( .A(n20182), .B(n20181), .Z(n20179) );
  XOR U28749 ( .A(y[5537]), .B(x[5537]), .Z(n20181) );
  XOR U28750 ( .A(y[5536]), .B(x[5536]), .Z(n20182) );
  XOR U28751 ( .A(y[5535]), .B(x[5535]), .Z(n20180) );
  NAND U28752 ( .A(n20243), .B(n20244), .Z(N63586) );
  NAND U28753 ( .A(n20245), .B(n20246), .Z(n20244) );
  NANDN U28754 ( .A(n20247), .B(n20248), .Z(n20246) );
  NANDN U28755 ( .A(n20248), .B(n20247), .Z(n20243) );
  XOR U28756 ( .A(n20247), .B(n20249), .Z(N63585) );
  XNOR U28757 ( .A(n20245), .B(n20248), .Z(n20249) );
  NAND U28758 ( .A(n20250), .B(n20251), .Z(n20248) );
  NAND U28759 ( .A(n20252), .B(n20253), .Z(n20251) );
  NANDN U28760 ( .A(n20254), .B(n20255), .Z(n20253) );
  NANDN U28761 ( .A(n20255), .B(n20254), .Z(n20250) );
  AND U28762 ( .A(n20256), .B(n20257), .Z(n20245) );
  NAND U28763 ( .A(n20258), .B(n20259), .Z(n20257) );
  NANDN U28764 ( .A(n20260), .B(n20261), .Z(n20259) );
  NANDN U28765 ( .A(n20261), .B(n20260), .Z(n20256) );
  IV U28766 ( .A(n20262), .Z(n20261) );
  AND U28767 ( .A(n20263), .B(n20264), .Z(n20247) );
  NAND U28768 ( .A(n20265), .B(n20266), .Z(n20264) );
  NANDN U28769 ( .A(n20267), .B(n20268), .Z(n20266) );
  NANDN U28770 ( .A(n20268), .B(n20267), .Z(n20263) );
  XOR U28771 ( .A(n20260), .B(n20269), .Z(N63584) );
  XNOR U28772 ( .A(n20258), .B(n20262), .Z(n20269) );
  XOR U28773 ( .A(n20255), .B(n20270), .Z(n20262) );
  XNOR U28774 ( .A(n20252), .B(n20254), .Z(n20270) );
  AND U28775 ( .A(n20271), .B(n20272), .Z(n20254) );
  NANDN U28776 ( .A(n20273), .B(n20274), .Z(n20272) );
  OR U28777 ( .A(n20275), .B(n20276), .Z(n20274) );
  IV U28778 ( .A(n20277), .Z(n20276) );
  NANDN U28779 ( .A(n20277), .B(n20275), .Z(n20271) );
  AND U28780 ( .A(n20278), .B(n20279), .Z(n20252) );
  NAND U28781 ( .A(n20280), .B(n20281), .Z(n20279) );
  NANDN U28782 ( .A(n20282), .B(n20283), .Z(n20281) );
  NANDN U28783 ( .A(n20283), .B(n20282), .Z(n20278) );
  IV U28784 ( .A(n20284), .Z(n20283) );
  NAND U28785 ( .A(n20285), .B(n20286), .Z(n20255) );
  NANDN U28786 ( .A(n20287), .B(n20288), .Z(n20286) );
  NANDN U28787 ( .A(n20289), .B(n20290), .Z(n20288) );
  NANDN U28788 ( .A(n20290), .B(n20289), .Z(n20285) );
  IV U28789 ( .A(n20291), .Z(n20289) );
  AND U28790 ( .A(n20292), .B(n20293), .Z(n20258) );
  NAND U28791 ( .A(n20294), .B(n20295), .Z(n20293) );
  NANDN U28792 ( .A(n20296), .B(n20297), .Z(n20295) );
  NANDN U28793 ( .A(n20297), .B(n20296), .Z(n20292) );
  XOR U28794 ( .A(n20268), .B(n20298), .Z(n20260) );
  XNOR U28795 ( .A(n20265), .B(n20267), .Z(n20298) );
  AND U28796 ( .A(n20299), .B(n20300), .Z(n20267) );
  NANDN U28797 ( .A(n20301), .B(n20302), .Z(n20300) );
  OR U28798 ( .A(n20303), .B(n20304), .Z(n20302) );
  IV U28799 ( .A(n20305), .Z(n20304) );
  NANDN U28800 ( .A(n20305), .B(n20303), .Z(n20299) );
  AND U28801 ( .A(n20306), .B(n20307), .Z(n20265) );
  NAND U28802 ( .A(n20308), .B(n20309), .Z(n20307) );
  NANDN U28803 ( .A(n20310), .B(n20311), .Z(n20309) );
  NANDN U28804 ( .A(n20311), .B(n20310), .Z(n20306) );
  IV U28805 ( .A(n20312), .Z(n20311) );
  NAND U28806 ( .A(n20313), .B(n20314), .Z(n20268) );
  NANDN U28807 ( .A(n20315), .B(n20316), .Z(n20314) );
  NANDN U28808 ( .A(n20317), .B(n20318), .Z(n20316) );
  NANDN U28809 ( .A(n20318), .B(n20317), .Z(n20313) );
  IV U28810 ( .A(n20319), .Z(n20317) );
  XOR U28811 ( .A(n20294), .B(n20320), .Z(N63583) );
  XNOR U28812 ( .A(n20297), .B(n20296), .Z(n20320) );
  XNOR U28813 ( .A(n20308), .B(n20321), .Z(n20296) );
  XNOR U28814 ( .A(n20312), .B(n20310), .Z(n20321) );
  XOR U28815 ( .A(n20318), .B(n20322), .Z(n20310) );
  XNOR U28816 ( .A(n20315), .B(n20319), .Z(n20322) );
  AND U28817 ( .A(n20323), .B(n20324), .Z(n20319) );
  NAND U28818 ( .A(n20325), .B(n20326), .Z(n20324) );
  NAND U28819 ( .A(n20327), .B(n20328), .Z(n20323) );
  AND U28820 ( .A(n20329), .B(n20330), .Z(n20315) );
  NAND U28821 ( .A(n20331), .B(n20332), .Z(n20330) );
  NAND U28822 ( .A(n20333), .B(n20334), .Z(n20329) );
  NANDN U28823 ( .A(n20335), .B(n20336), .Z(n20318) );
  ANDN U28824 ( .B(n20337), .A(n20338), .Z(n20312) );
  XNOR U28825 ( .A(n20303), .B(n20339), .Z(n20308) );
  XNOR U28826 ( .A(n20301), .B(n20305), .Z(n20339) );
  AND U28827 ( .A(n20340), .B(n20341), .Z(n20305) );
  NAND U28828 ( .A(n20342), .B(n20343), .Z(n20341) );
  NAND U28829 ( .A(n20344), .B(n20345), .Z(n20340) );
  AND U28830 ( .A(n20346), .B(n20347), .Z(n20301) );
  NAND U28831 ( .A(n20348), .B(n20349), .Z(n20347) );
  NAND U28832 ( .A(n20350), .B(n20351), .Z(n20346) );
  AND U28833 ( .A(n20352), .B(n20353), .Z(n20303) );
  NAND U28834 ( .A(n20354), .B(n20355), .Z(n20297) );
  XNOR U28835 ( .A(n20280), .B(n20356), .Z(n20294) );
  XNOR U28836 ( .A(n20284), .B(n20282), .Z(n20356) );
  XOR U28837 ( .A(n20290), .B(n20357), .Z(n20282) );
  XNOR U28838 ( .A(n20287), .B(n20291), .Z(n20357) );
  AND U28839 ( .A(n20358), .B(n20359), .Z(n20291) );
  NAND U28840 ( .A(n20360), .B(n20361), .Z(n20359) );
  NAND U28841 ( .A(n20362), .B(n20363), .Z(n20358) );
  AND U28842 ( .A(n20364), .B(n20365), .Z(n20287) );
  NAND U28843 ( .A(n20366), .B(n20367), .Z(n20365) );
  NAND U28844 ( .A(n20368), .B(n20369), .Z(n20364) );
  NANDN U28845 ( .A(n20370), .B(n20371), .Z(n20290) );
  ANDN U28846 ( .B(n20372), .A(n20373), .Z(n20284) );
  XNOR U28847 ( .A(n20275), .B(n20374), .Z(n20280) );
  XNOR U28848 ( .A(n20273), .B(n20277), .Z(n20374) );
  AND U28849 ( .A(n20375), .B(n20376), .Z(n20277) );
  NAND U28850 ( .A(n20377), .B(n20378), .Z(n20376) );
  NAND U28851 ( .A(n20379), .B(n20380), .Z(n20375) );
  AND U28852 ( .A(n20381), .B(n20382), .Z(n20273) );
  NAND U28853 ( .A(n20383), .B(n20384), .Z(n20382) );
  NAND U28854 ( .A(n20385), .B(n20386), .Z(n20381) );
  AND U28855 ( .A(n20387), .B(n20388), .Z(n20275) );
  XOR U28856 ( .A(n20355), .B(n20354), .Z(N63582) );
  XNOR U28857 ( .A(n20372), .B(n20373), .Z(n20354) );
  XNOR U28858 ( .A(n20387), .B(n20388), .Z(n20373) );
  XOR U28859 ( .A(n20384), .B(n20383), .Z(n20388) );
  XOR U28860 ( .A(y[5532]), .B(x[5532]), .Z(n20383) );
  XOR U28861 ( .A(n20386), .B(n20385), .Z(n20384) );
  XOR U28862 ( .A(y[5534]), .B(x[5534]), .Z(n20385) );
  XOR U28863 ( .A(y[5533]), .B(x[5533]), .Z(n20386) );
  XOR U28864 ( .A(n20378), .B(n20377), .Z(n20387) );
  XOR U28865 ( .A(n20380), .B(n20379), .Z(n20377) );
  XOR U28866 ( .A(y[5531]), .B(x[5531]), .Z(n20379) );
  XOR U28867 ( .A(y[5530]), .B(x[5530]), .Z(n20380) );
  XOR U28868 ( .A(y[5529]), .B(x[5529]), .Z(n20378) );
  XNOR U28869 ( .A(n20371), .B(n20370), .Z(n20372) );
  XNOR U28870 ( .A(n20367), .B(n20366), .Z(n20370) );
  XOR U28871 ( .A(n20369), .B(n20368), .Z(n20366) );
  XOR U28872 ( .A(y[5528]), .B(x[5528]), .Z(n20368) );
  XOR U28873 ( .A(y[5527]), .B(x[5527]), .Z(n20369) );
  XOR U28874 ( .A(y[5526]), .B(x[5526]), .Z(n20367) );
  XOR U28875 ( .A(n20361), .B(n20360), .Z(n20371) );
  XOR U28876 ( .A(n20363), .B(n20362), .Z(n20360) );
  XOR U28877 ( .A(y[5525]), .B(x[5525]), .Z(n20362) );
  XOR U28878 ( .A(y[5524]), .B(x[5524]), .Z(n20363) );
  XOR U28879 ( .A(y[5523]), .B(x[5523]), .Z(n20361) );
  XNOR U28880 ( .A(n20337), .B(n20338), .Z(n20355) );
  XNOR U28881 ( .A(n20352), .B(n20353), .Z(n20338) );
  XOR U28882 ( .A(n20349), .B(n20348), .Z(n20353) );
  XOR U28883 ( .A(y[5520]), .B(x[5520]), .Z(n20348) );
  XOR U28884 ( .A(n20351), .B(n20350), .Z(n20349) );
  XOR U28885 ( .A(y[5522]), .B(x[5522]), .Z(n20350) );
  XOR U28886 ( .A(y[5521]), .B(x[5521]), .Z(n20351) );
  XOR U28887 ( .A(n20343), .B(n20342), .Z(n20352) );
  XOR U28888 ( .A(n20345), .B(n20344), .Z(n20342) );
  XOR U28889 ( .A(y[5519]), .B(x[5519]), .Z(n20344) );
  XOR U28890 ( .A(y[5518]), .B(x[5518]), .Z(n20345) );
  XOR U28891 ( .A(y[5517]), .B(x[5517]), .Z(n20343) );
  XNOR U28892 ( .A(n20336), .B(n20335), .Z(n20337) );
  XNOR U28893 ( .A(n20332), .B(n20331), .Z(n20335) );
  XOR U28894 ( .A(n20334), .B(n20333), .Z(n20331) );
  XOR U28895 ( .A(y[5516]), .B(x[5516]), .Z(n20333) );
  XOR U28896 ( .A(y[5515]), .B(x[5515]), .Z(n20334) );
  XOR U28897 ( .A(y[5514]), .B(x[5514]), .Z(n20332) );
  XOR U28898 ( .A(n20326), .B(n20325), .Z(n20336) );
  XOR U28899 ( .A(n20328), .B(n20327), .Z(n20325) );
  XOR U28900 ( .A(y[5513]), .B(x[5513]), .Z(n20327) );
  XOR U28901 ( .A(y[5512]), .B(x[5512]), .Z(n20328) );
  XOR U28902 ( .A(y[5511]), .B(x[5511]), .Z(n20326) );
  NAND U28903 ( .A(n20389), .B(n20390), .Z(N63573) );
  NAND U28904 ( .A(n20391), .B(n20392), .Z(n20390) );
  NANDN U28905 ( .A(n20393), .B(n20394), .Z(n20392) );
  NANDN U28906 ( .A(n20394), .B(n20393), .Z(n20389) );
  XOR U28907 ( .A(n20393), .B(n20395), .Z(N63572) );
  XNOR U28908 ( .A(n20391), .B(n20394), .Z(n20395) );
  NAND U28909 ( .A(n20396), .B(n20397), .Z(n20394) );
  NAND U28910 ( .A(n20398), .B(n20399), .Z(n20397) );
  NANDN U28911 ( .A(n20400), .B(n20401), .Z(n20399) );
  NANDN U28912 ( .A(n20401), .B(n20400), .Z(n20396) );
  AND U28913 ( .A(n20402), .B(n20403), .Z(n20391) );
  NAND U28914 ( .A(n20404), .B(n20405), .Z(n20403) );
  NANDN U28915 ( .A(n20406), .B(n20407), .Z(n20405) );
  NANDN U28916 ( .A(n20407), .B(n20406), .Z(n20402) );
  IV U28917 ( .A(n20408), .Z(n20407) );
  AND U28918 ( .A(n20409), .B(n20410), .Z(n20393) );
  NAND U28919 ( .A(n20411), .B(n20412), .Z(n20410) );
  NANDN U28920 ( .A(n20413), .B(n20414), .Z(n20412) );
  NANDN U28921 ( .A(n20414), .B(n20413), .Z(n20409) );
  XOR U28922 ( .A(n20406), .B(n20415), .Z(N63571) );
  XNOR U28923 ( .A(n20404), .B(n20408), .Z(n20415) );
  XOR U28924 ( .A(n20401), .B(n20416), .Z(n20408) );
  XNOR U28925 ( .A(n20398), .B(n20400), .Z(n20416) );
  AND U28926 ( .A(n20417), .B(n20418), .Z(n20400) );
  NANDN U28927 ( .A(n20419), .B(n20420), .Z(n20418) );
  OR U28928 ( .A(n20421), .B(n20422), .Z(n20420) );
  IV U28929 ( .A(n20423), .Z(n20422) );
  NANDN U28930 ( .A(n20423), .B(n20421), .Z(n20417) );
  AND U28931 ( .A(n20424), .B(n20425), .Z(n20398) );
  NAND U28932 ( .A(n20426), .B(n20427), .Z(n20425) );
  NANDN U28933 ( .A(n20428), .B(n20429), .Z(n20427) );
  NANDN U28934 ( .A(n20429), .B(n20428), .Z(n20424) );
  IV U28935 ( .A(n20430), .Z(n20429) );
  NAND U28936 ( .A(n20431), .B(n20432), .Z(n20401) );
  NANDN U28937 ( .A(n20433), .B(n20434), .Z(n20432) );
  NANDN U28938 ( .A(n20435), .B(n20436), .Z(n20434) );
  NANDN U28939 ( .A(n20436), .B(n20435), .Z(n20431) );
  IV U28940 ( .A(n20437), .Z(n20435) );
  AND U28941 ( .A(n20438), .B(n20439), .Z(n20404) );
  NAND U28942 ( .A(n20440), .B(n20441), .Z(n20439) );
  NANDN U28943 ( .A(n20442), .B(n20443), .Z(n20441) );
  NANDN U28944 ( .A(n20443), .B(n20442), .Z(n20438) );
  XOR U28945 ( .A(n20414), .B(n20444), .Z(n20406) );
  XNOR U28946 ( .A(n20411), .B(n20413), .Z(n20444) );
  AND U28947 ( .A(n20445), .B(n20446), .Z(n20413) );
  NANDN U28948 ( .A(n20447), .B(n20448), .Z(n20446) );
  OR U28949 ( .A(n20449), .B(n20450), .Z(n20448) );
  IV U28950 ( .A(n20451), .Z(n20450) );
  NANDN U28951 ( .A(n20451), .B(n20449), .Z(n20445) );
  AND U28952 ( .A(n20452), .B(n20453), .Z(n20411) );
  NAND U28953 ( .A(n20454), .B(n20455), .Z(n20453) );
  NANDN U28954 ( .A(n20456), .B(n20457), .Z(n20455) );
  NANDN U28955 ( .A(n20457), .B(n20456), .Z(n20452) );
  IV U28956 ( .A(n20458), .Z(n20457) );
  NAND U28957 ( .A(n20459), .B(n20460), .Z(n20414) );
  NANDN U28958 ( .A(n20461), .B(n20462), .Z(n20460) );
  NANDN U28959 ( .A(n20463), .B(n20464), .Z(n20462) );
  NANDN U28960 ( .A(n20464), .B(n20463), .Z(n20459) );
  IV U28961 ( .A(n20465), .Z(n20463) );
  XOR U28962 ( .A(n20440), .B(n20466), .Z(N63570) );
  XNOR U28963 ( .A(n20443), .B(n20442), .Z(n20466) );
  XNOR U28964 ( .A(n20454), .B(n20467), .Z(n20442) );
  XNOR U28965 ( .A(n20458), .B(n20456), .Z(n20467) );
  XOR U28966 ( .A(n20464), .B(n20468), .Z(n20456) );
  XNOR U28967 ( .A(n20461), .B(n20465), .Z(n20468) );
  AND U28968 ( .A(n20469), .B(n20470), .Z(n20465) );
  NAND U28969 ( .A(n20471), .B(n20472), .Z(n20470) );
  NAND U28970 ( .A(n20473), .B(n20474), .Z(n20469) );
  AND U28971 ( .A(n20475), .B(n20476), .Z(n20461) );
  NAND U28972 ( .A(n20477), .B(n20478), .Z(n20476) );
  NAND U28973 ( .A(n20479), .B(n20480), .Z(n20475) );
  NANDN U28974 ( .A(n20481), .B(n20482), .Z(n20464) );
  ANDN U28975 ( .B(n20483), .A(n20484), .Z(n20458) );
  XNOR U28976 ( .A(n20449), .B(n20485), .Z(n20454) );
  XNOR U28977 ( .A(n20447), .B(n20451), .Z(n20485) );
  AND U28978 ( .A(n20486), .B(n20487), .Z(n20451) );
  NAND U28979 ( .A(n20488), .B(n20489), .Z(n20487) );
  NAND U28980 ( .A(n20490), .B(n20491), .Z(n20486) );
  AND U28981 ( .A(n20492), .B(n20493), .Z(n20447) );
  NAND U28982 ( .A(n20494), .B(n20495), .Z(n20493) );
  NAND U28983 ( .A(n20496), .B(n20497), .Z(n20492) );
  AND U28984 ( .A(n20498), .B(n20499), .Z(n20449) );
  NAND U28985 ( .A(n20500), .B(n20501), .Z(n20443) );
  XNOR U28986 ( .A(n20426), .B(n20502), .Z(n20440) );
  XNOR U28987 ( .A(n20430), .B(n20428), .Z(n20502) );
  XOR U28988 ( .A(n20436), .B(n20503), .Z(n20428) );
  XNOR U28989 ( .A(n20433), .B(n20437), .Z(n20503) );
  AND U28990 ( .A(n20504), .B(n20505), .Z(n20437) );
  NAND U28991 ( .A(n20506), .B(n20507), .Z(n20505) );
  NAND U28992 ( .A(n20508), .B(n20509), .Z(n20504) );
  AND U28993 ( .A(n20510), .B(n20511), .Z(n20433) );
  NAND U28994 ( .A(n20512), .B(n20513), .Z(n20511) );
  NAND U28995 ( .A(n20514), .B(n20515), .Z(n20510) );
  NANDN U28996 ( .A(n20516), .B(n20517), .Z(n20436) );
  ANDN U28997 ( .B(n20518), .A(n20519), .Z(n20430) );
  XNOR U28998 ( .A(n20421), .B(n20520), .Z(n20426) );
  XNOR U28999 ( .A(n20419), .B(n20423), .Z(n20520) );
  AND U29000 ( .A(n20521), .B(n20522), .Z(n20423) );
  NAND U29001 ( .A(n20523), .B(n20524), .Z(n20522) );
  NAND U29002 ( .A(n20525), .B(n20526), .Z(n20521) );
  AND U29003 ( .A(n20527), .B(n20528), .Z(n20419) );
  NAND U29004 ( .A(n20529), .B(n20530), .Z(n20528) );
  NAND U29005 ( .A(n20531), .B(n20532), .Z(n20527) );
  AND U29006 ( .A(n20533), .B(n20534), .Z(n20421) );
  XOR U29007 ( .A(n20501), .B(n20500), .Z(N63569) );
  XNOR U29008 ( .A(n20518), .B(n20519), .Z(n20500) );
  XNOR U29009 ( .A(n20533), .B(n20534), .Z(n20519) );
  XOR U29010 ( .A(n20530), .B(n20529), .Z(n20534) );
  XOR U29011 ( .A(y[5508]), .B(x[5508]), .Z(n20529) );
  XOR U29012 ( .A(n20532), .B(n20531), .Z(n20530) );
  XOR U29013 ( .A(y[5510]), .B(x[5510]), .Z(n20531) );
  XOR U29014 ( .A(y[5509]), .B(x[5509]), .Z(n20532) );
  XOR U29015 ( .A(n20524), .B(n20523), .Z(n20533) );
  XOR U29016 ( .A(n20526), .B(n20525), .Z(n20523) );
  XOR U29017 ( .A(y[5507]), .B(x[5507]), .Z(n20525) );
  XOR U29018 ( .A(y[5506]), .B(x[5506]), .Z(n20526) );
  XOR U29019 ( .A(y[5505]), .B(x[5505]), .Z(n20524) );
  XNOR U29020 ( .A(n20517), .B(n20516), .Z(n20518) );
  XNOR U29021 ( .A(n20513), .B(n20512), .Z(n20516) );
  XOR U29022 ( .A(n20515), .B(n20514), .Z(n20512) );
  XOR U29023 ( .A(y[5504]), .B(x[5504]), .Z(n20514) );
  XOR U29024 ( .A(y[5503]), .B(x[5503]), .Z(n20515) );
  XOR U29025 ( .A(y[5502]), .B(x[5502]), .Z(n20513) );
  XOR U29026 ( .A(n20507), .B(n20506), .Z(n20517) );
  XOR U29027 ( .A(n20509), .B(n20508), .Z(n20506) );
  XOR U29028 ( .A(y[5501]), .B(x[5501]), .Z(n20508) );
  XOR U29029 ( .A(y[5500]), .B(x[5500]), .Z(n20509) );
  XOR U29030 ( .A(y[5499]), .B(x[5499]), .Z(n20507) );
  XNOR U29031 ( .A(n20483), .B(n20484), .Z(n20501) );
  XNOR U29032 ( .A(n20498), .B(n20499), .Z(n20484) );
  XOR U29033 ( .A(n20495), .B(n20494), .Z(n20499) );
  XOR U29034 ( .A(y[5496]), .B(x[5496]), .Z(n20494) );
  XOR U29035 ( .A(n20497), .B(n20496), .Z(n20495) );
  XOR U29036 ( .A(y[5498]), .B(x[5498]), .Z(n20496) );
  XOR U29037 ( .A(y[5497]), .B(x[5497]), .Z(n20497) );
  XOR U29038 ( .A(n20489), .B(n20488), .Z(n20498) );
  XOR U29039 ( .A(n20491), .B(n20490), .Z(n20488) );
  XOR U29040 ( .A(y[5495]), .B(x[5495]), .Z(n20490) );
  XOR U29041 ( .A(y[5494]), .B(x[5494]), .Z(n20491) );
  XOR U29042 ( .A(y[5493]), .B(x[5493]), .Z(n20489) );
  XNOR U29043 ( .A(n20482), .B(n20481), .Z(n20483) );
  XNOR U29044 ( .A(n20478), .B(n20477), .Z(n20481) );
  XOR U29045 ( .A(n20480), .B(n20479), .Z(n20477) );
  XOR U29046 ( .A(y[5492]), .B(x[5492]), .Z(n20479) );
  XOR U29047 ( .A(y[5491]), .B(x[5491]), .Z(n20480) );
  XOR U29048 ( .A(y[5490]), .B(x[5490]), .Z(n20478) );
  XOR U29049 ( .A(n20472), .B(n20471), .Z(n20482) );
  XOR U29050 ( .A(n20474), .B(n20473), .Z(n20471) );
  XOR U29051 ( .A(y[5489]), .B(x[5489]), .Z(n20473) );
  XOR U29052 ( .A(y[5488]), .B(x[5488]), .Z(n20474) );
  XOR U29053 ( .A(y[5487]), .B(x[5487]), .Z(n20472) );
  NAND U29054 ( .A(n20535), .B(n20536), .Z(N63560) );
  NAND U29055 ( .A(n20537), .B(n20538), .Z(n20536) );
  NANDN U29056 ( .A(n20539), .B(n20540), .Z(n20538) );
  NANDN U29057 ( .A(n20540), .B(n20539), .Z(n20535) );
  XOR U29058 ( .A(n20539), .B(n20541), .Z(N63559) );
  XNOR U29059 ( .A(n20537), .B(n20540), .Z(n20541) );
  NAND U29060 ( .A(n20542), .B(n20543), .Z(n20540) );
  NAND U29061 ( .A(n20544), .B(n20545), .Z(n20543) );
  NANDN U29062 ( .A(n20546), .B(n20547), .Z(n20545) );
  NANDN U29063 ( .A(n20547), .B(n20546), .Z(n20542) );
  AND U29064 ( .A(n20548), .B(n20549), .Z(n20537) );
  NAND U29065 ( .A(n20550), .B(n20551), .Z(n20549) );
  NANDN U29066 ( .A(n20552), .B(n20553), .Z(n20551) );
  NANDN U29067 ( .A(n20553), .B(n20552), .Z(n20548) );
  IV U29068 ( .A(n20554), .Z(n20553) );
  AND U29069 ( .A(n20555), .B(n20556), .Z(n20539) );
  NAND U29070 ( .A(n20557), .B(n20558), .Z(n20556) );
  NANDN U29071 ( .A(n20559), .B(n20560), .Z(n20558) );
  NANDN U29072 ( .A(n20560), .B(n20559), .Z(n20555) );
  XOR U29073 ( .A(n20552), .B(n20561), .Z(N63558) );
  XNOR U29074 ( .A(n20550), .B(n20554), .Z(n20561) );
  XOR U29075 ( .A(n20547), .B(n20562), .Z(n20554) );
  XNOR U29076 ( .A(n20544), .B(n20546), .Z(n20562) );
  AND U29077 ( .A(n20563), .B(n20564), .Z(n20546) );
  NANDN U29078 ( .A(n20565), .B(n20566), .Z(n20564) );
  OR U29079 ( .A(n20567), .B(n20568), .Z(n20566) );
  IV U29080 ( .A(n20569), .Z(n20568) );
  NANDN U29081 ( .A(n20569), .B(n20567), .Z(n20563) );
  AND U29082 ( .A(n20570), .B(n20571), .Z(n20544) );
  NAND U29083 ( .A(n20572), .B(n20573), .Z(n20571) );
  NANDN U29084 ( .A(n20574), .B(n20575), .Z(n20573) );
  NANDN U29085 ( .A(n20575), .B(n20574), .Z(n20570) );
  IV U29086 ( .A(n20576), .Z(n20575) );
  NAND U29087 ( .A(n20577), .B(n20578), .Z(n20547) );
  NANDN U29088 ( .A(n20579), .B(n20580), .Z(n20578) );
  NANDN U29089 ( .A(n20581), .B(n20582), .Z(n20580) );
  NANDN U29090 ( .A(n20582), .B(n20581), .Z(n20577) );
  IV U29091 ( .A(n20583), .Z(n20581) );
  AND U29092 ( .A(n20584), .B(n20585), .Z(n20550) );
  NAND U29093 ( .A(n20586), .B(n20587), .Z(n20585) );
  NANDN U29094 ( .A(n20588), .B(n20589), .Z(n20587) );
  NANDN U29095 ( .A(n20589), .B(n20588), .Z(n20584) );
  XOR U29096 ( .A(n20560), .B(n20590), .Z(n20552) );
  XNOR U29097 ( .A(n20557), .B(n20559), .Z(n20590) );
  AND U29098 ( .A(n20591), .B(n20592), .Z(n20559) );
  NANDN U29099 ( .A(n20593), .B(n20594), .Z(n20592) );
  OR U29100 ( .A(n20595), .B(n20596), .Z(n20594) );
  IV U29101 ( .A(n20597), .Z(n20596) );
  NANDN U29102 ( .A(n20597), .B(n20595), .Z(n20591) );
  AND U29103 ( .A(n20598), .B(n20599), .Z(n20557) );
  NAND U29104 ( .A(n20600), .B(n20601), .Z(n20599) );
  NANDN U29105 ( .A(n20602), .B(n20603), .Z(n20601) );
  NANDN U29106 ( .A(n20603), .B(n20602), .Z(n20598) );
  IV U29107 ( .A(n20604), .Z(n20603) );
  NAND U29108 ( .A(n20605), .B(n20606), .Z(n20560) );
  NANDN U29109 ( .A(n20607), .B(n20608), .Z(n20606) );
  NANDN U29110 ( .A(n20609), .B(n20610), .Z(n20608) );
  NANDN U29111 ( .A(n20610), .B(n20609), .Z(n20605) );
  IV U29112 ( .A(n20611), .Z(n20609) );
  XOR U29113 ( .A(n20586), .B(n20612), .Z(N63557) );
  XNOR U29114 ( .A(n20589), .B(n20588), .Z(n20612) );
  XNOR U29115 ( .A(n20600), .B(n20613), .Z(n20588) );
  XNOR U29116 ( .A(n20604), .B(n20602), .Z(n20613) );
  XOR U29117 ( .A(n20610), .B(n20614), .Z(n20602) );
  XNOR U29118 ( .A(n20607), .B(n20611), .Z(n20614) );
  AND U29119 ( .A(n20615), .B(n20616), .Z(n20611) );
  NAND U29120 ( .A(n20617), .B(n20618), .Z(n20616) );
  NAND U29121 ( .A(n20619), .B(n20620), .Z(n20615) );
  AND U29122 ( .A(n20621), .B(n20622), .Z(n20607) );
  NAND U29123 ( .A(n20623), .B(n20624), .Z(n20622) );
  NAND U29124 ( .A(n20625), .B(n20626), .Z(n20621) );
  NANDN U29125 ( .A(n20627), .B(n20628), .Z(n20610) );
  ANDN U29126 ( .B(n20629), .A(n20630), .Z(n20604) );
  XNOR U29127 ( .A(n20595), .B(n20631), .Z(n20600) );
  XNOR U29128 ( .A(n20593), .B(n20597), .Z(n20631) );
  AND U29129 ( .A(n20632), .B(n20633), .Z(n20597) );
  NAND U29130 ( .A(n20634), .B(n20635), .Z(n20633) );
  NAND U29131 ( .A(n20636), .B(n20637), .Z(n20632) );
  AND U29132 ( .A(n20638), .B(n20639), .Z(n20593) );
  NAND U29133 ( .A(n20640), .B(n20641), .Z(n20639) );
  NAND U29134 ( .A(n20642), .B(n20643), .Z(n20638) );
  AND U29135 ( .A(n20644), .B(n20645), .Z(n20595) );
  NAND U29136 ( .A(n20646), .B(n20647), .Z(n20589) );
  XNOR U29137 ( .A(n20572), .B(n20648), .Z(n20586) );
  XNOR U29138 ( .A(n20576), .B(n20574), .Z(n20648) );
  XOR U29139 ( .A(n20582), .B(n20649), .Z(n20574) );
  XNOR U29140 ( .A(n20579), .B(n20583), .Z(n20649) );
  AND U29141 ( .A(n20650), .B(n20651), .Z(n20583) );
  NAND U29142 ( .A(n20652), .B(n20653), .Z(n20651) );
  NAND U29143 ( .A(n20654), .B(n20655), .Z(n20650) );
  AND U29144 ( .A(n20656), .B(n20657), .Z(n20579) );
  NAND U29145 ( .A(n20658), .B(n20659), .Z(n20657) );
  NAND U29146 ( .A(n20660), .B(n20661), .Z(n20656) );
  NANDN U29147 ( .A(n20662), .B(n20663), .Z(n20582) );
  ANDN U29148 ( .B(n20664), .A(n20665), .Z(n20576) );
  XNOR U29149 ( .A(n20567), .B(n20666), .Z(n20572) );
  XNOR U29150 ( .A(n20565), .B(n20569), .Z(n20666) );
  AND U29151 ( .A(n20667), .B(n20668), .Z(n20569) );
  NAND U29152 ( .A(n20669), .B(n20670), .Z(n20668) );
  NAND U29153 ( .A(n20671), .B(n20672), .Z(n20667) );
  AND U29154 ( .A(n20673), .B(n20674), .Z(n20565) );
  NAND U29155 ( .A(n20675), .B(n20676), .Z(n20674) );
  NAND U29156 ( .A(n20677), .B(n20678), .Z(n20673) );
  AND U29157 ( .A(n20679), .B(n20680), .Z(n20567) );
  XOR U29158 ( .A(n20647), .B(n20646), .Z(N63556) );
  XNOR U29159 ( .A(n20664), .B(n20665), .Z(n20646) );
  XNOR U29160 ( .A(n20679), .B(n20680), .Z(n20665) );
  XOR U29161 ( .A(n20676), .B(n20675), .Z(n20680) );
  XOR U29162 ( .A(y[5484]), .B(x[5484]), .Z(n20675) );
  XOR U29163 ( .A(n20678), .B(n20677), .Z(n20676) );
  XOR U29164 ( .A(y[5486]), .B(x[5486]), .Z(n20677) );
  XOR U29165 ( .A(y[5485]), .B(x[5485]), .Z(n20678) );
  XOR U29166 ( .A(n20670), .B(n20669), .Z(n20679) );
  XOR U29167 ( .A(n20672), .B(n20671), .Z(n20669) );
  XOR U29168 ( .A(y[5483]), .B(x[5483]), .Z(n20671) );
  XOR U29169 ( .A(y[5482]), .B(x[5482]), .Z(n20672) );
  XOR U29170 ( .A(y[5481]), .B(x[5481]), .Z(n20670) );
  XNOR U29171 ( .A(n20663), .B(n20662), .Z(n20664) );
  XNOR U29172 ( .A(n20659), .B(n20658), .Z(n20662) );
  XOR U29173 ( .A(n20661), .B(n20660), .Z(n20658) );
  XOR U29174 ( .A(y[5480]), .B(x[5480]), .Z(n20660) );
  XOR U29175 ( .A(y[5479]), .B(x[5479]), .Z(n20661) );
  XOR U29176 ( .A(y[5478]), .B(x[5478]), .Z(n20659) );
  XOR U29177 ( .A(n20653), .B(n20652), .Z(n20663) );
  XOR U29178 ( .A(n20655), .B(n20654), .Z(n20652) );
  XOR U29179 ( .A(y[5477]), .B(x[5477]), .Z(n20654) );
  XOR U29180 ( .A(y[5476]), .B(x[5476]), .Z(n20655) );
  XOR U29181 ( .A(y[5475]), .B(x[5475]), .Z(n20653) );
  XNOR U29182 ( .A(n20629), .B(n20630), .Z(n20647) );
  XNOR U29183 ( .A(n20644), .B(n20645), .Z(n20630) );
  XOR U29184 ( .A(n20641), .B(n20640), .Z(n20645) );
  XOR U29185 ( .A(y[5472]), .B(x[5472]), .Z(n20640) );
  XOR U29186 ( .A(n20643), .B(n20642), .Z(n20641) );
  XOR U29187 ( .A(y[5474]), .B(x[5474]), .Z(n20642) );
  XOR U29188 ( .A(y[5473]), .B(x[5473]), .Z(n20643) );
  XOR U29189 ( .A(n20635), .B(n20634), .Z(n20644) );
  XOR U29190 ( .A(n20637), .B(n20636), .Z(n20634) );
  XOR U29191 ( .A(y[5471]), .B(x[5471]), .Z(n20636) );
  XOR U29192 ( .A(y[5470]), .B(x[5470]), .Z(n20637) );
  XOR U29193 ( .A(y[5469]), .B(x[5469]), .Z(n20635) );
  XNOR U29194 ( .A(n20628), .B(n20627), .Z(n20629) );
  XNOR U29195 ( .A(n20624), .B(n20623), .Z(n20627) );
  XOR U29196 ( .A(n20626), .B(n20625), .Z(n20623) );
  XOR U29197 ( .A(y[5468]), .B(x[5468]), .Z(n20625) );
  XOR U29198 ( .A(y[5467]), .B(x[5467]), .Z(n20626) );
  XOR U29199 ( .A(y[5466]), .B(x[5466]), .Z(n20624) );
  XOR U29200 ( .A(n20618), .B(n20617), .Z(n20628) );
  XOR U29201 ( .A(n20620), .B(n20619), .Z(n20617) );
  XOR U29202 ( .A(y[5465]), .B(x[5465]), .Z(n20619) );
  XOR U29203 ( .A(y[5464]), .B(x[5464]), .Z(n20620) );
  XOR U29204 ( .A(y[5463]), .B(x[5463]), .Z(n20618) );
  NAND U29205 ( .A(n20681), .B(n20682), .Z(N63547) );
  NAND U29206 ( .A(n20683), .B(n20684), .Z(n20682) );
  NANDN U29207 ( .A(n20685), .B(n20686), .Z(n20684) );
  NANDN U29208 ( .A(n20686), .B(n20685), .Z(n20681) );
  XOR U29209 ( .A(n20685), .B(n20687), .Z(N63546) );
  XNOR U29210 ( .A(n20683), .B(n20686), .Z(n20687) );
  NAND U29211 ( .A(n20688), .B(n20689), .Z(n20686) );
  NAND U29212 ( .A(n20690), .B(n20691), .Z(n20689) );
  NANDN U29213 ( .A(n20692), .B(n20693), .Z(n20691) );
  NANDN U29214 ( .A(n20693), .B(n20692), .Z(n20688) );
  AND U29215 ( .A(n20694), .B(n20695), .Z(n20683) );
  NAND U29216 ( .A(n20696), .B(n20697), .Z(n20695) );
  NANDN U29217 ( .A(n20698), .B(n20699), .Z(n20697) );
  NANDN U29218 ( .A(n20699), .B(n20698), .Z(n20694) );
  IV U29219 ( .A(n20700), .Z(n20699) );
  AND U29220 ( .A(n20701), .B(n20702), .Z(n20685) );
  NAND U29221 ( .A(n20703), .B(n20704), .Z(n20702) );
  NANDN U29222 ( .A(n20705), .B(n20706), .Z(n20704) );
  NANDN U29223 ( .A(n20706), .B(n20705), .Z(n20701) );
  XOR U29224 ( .A(n20698), .B(n20707), .Z(N63545) );
  XNOR U29225 ( .A(n20696), .B(n20700), .Z(n20707) );
  XOR U29226 ( .A(n20693), .B(n20708), .Z(n20700) );
  XNOR U29227 ( .A(n20690), .B(n20692), .Z(n20708) );
  AND U29228 ( .A(n20709), .B(n20710), .Z(n20692) );
  NANDN U29229 ( .A(n20711), .B(n20712), .Z(n20710) );
  OR U29230 ( .A(n20713), .B(n20714), .Z(n20712) );
  IV U29231 ( .A(n20715), .Z(n20714) );
  NANDN U29232 ( .A(n20715), .B(n20713), .Z(n20709) );
  AND U29233 ( .A(n20716), .B(n20717), .Z(n20690) );
  NAND U29234 ( .A(n20718), .B(n20719), .Z(n20717) );
  NANDN U29235 ( .A(n20720), .B(n20721), .Z(n20719) );
  NANDN U29236 ( .A(n20721), .B(n20720), .Z(n20716) );
  IV U29237 ( .A(n20722), .Z(n20721) );
  NAND U29238 ( .A(n20723), .B(n20724), .Z(n20693) );
  NANDN U29239 ( .A(n20725), .B(n20726), .Z(n20724) );
  NANDN U29240 ( .A(n20727), .B(n20728), .Z(n20726) );
  NANDN U29241 ( .A(n20728), .B(n20727), .Z(n20723) );
  IV U29242 ( .A(n20729), .Z(n20727) );
  AND U29243 ( .A(n20730), .B(n20731), .Z(n20696) );
  NAND U29244 ( .A(n20732), .B(n20733), .Z(n20731) );
  NANDN U29245 ( .A(n20734), .B(n20735), .Z(n20733) );
  NANDN U29246 ( .A(n20735), .B(n20734), .Z(n20730) );
  XOR U29247 ( .A(n20706), .B(n20736), .Z(n20698) );
  XNOR U29248 ( .A(n20703), .B(n20705), .Z(n20736) );
  AND U29249 ( .A(n20737), .B(n20738), .Z(n20705) );
  NANDN U29250 ( .A(n20739), .B(n20740), .Z(n20738) );
  OR U29251 ( .A(n20741), .B(n20742), .Z(n20740) );
  IV U29252 ( .A(n20743), .Z(n20742) );
  NANDN U29253 ( .A(n20743), .B(n20741), .Z(n20737) );
  AND U29254 ( .A(n20744), .B(n20745), .Z(n20703) );
  NAND U29255 ( .A(n20746), .B(n20747), .Z(n20745) );
  NANDN U29256 ( .A(n20748), .B(n20749), .Z(n20747) );
  NANDN U29257 ( .A(n20749), .B(n20748), .Z(n20744) );
  IV U29258 ( .A(n20750), .Z(n20749) );
  NAND U29259 ( .A(n20751), .B(n20752), .Z(n20706) );
  NANDN U29260 ( .A(n20753), .B(n20754), .Z(n20752) );
  NANDN U29261 ( .A(n20755), .B(n20756), .Z(n20754) );
  NANDN U29262 ( .A(n20756), .B(n20755), .Z(n20751) );
  IV U29263 ( .A(n20757), .Z(n20755) );
  XOR U29264 ( .A(n20732), .B(n20758), .Z(N63544) );
  XNOR U29265 ( .A(n20735), .B(n20734), .Z(n20758) );
  XNOR U29266 ( .A(n20746), .B(n20759), .Z(n20734) );
  XNOR U29267 ( .A(n20750), .B(n20748), .Z(n20759) );
  XOR U29268 ( .A(n20756), .B(n20760), .Z(n20748) );
  XNOR U29269 ( .A(n20753), .B(n20757), .Z(n20760) );
  AND U29270 ( .A(n20761), .B(n20762), .Z(n20757) );
  NAND U29271 ( .A(n20763), .B(n20764), .Z(n20762) );
  NAND U29272 ( .A(n20765), .B(n20766), .Z(n20761) );
  AND U29273 ( .A(n20767), .B(n20768), .Z(n20753) );
  NAND U29274 ( .A(n20769), .B(n20770), .Z(n20768) );
  NAND U29275 ( .A(n20771), .B(n20772), .Z(n20767) );
  NANDN U29276 ( .A(n20773), .B(n20774), .Z(n20756) );
  ANDN U29277 ( .B(n20775), .A(n20776), .Z(n20750) );
  XNOR U29278 ( .A(n20741), .B(n20777), .Z(n20746) );
  XNOR U29279 ( .A(n20739), .B(n20743), .Z(n20777) );
  AND U29280 ( .A(n20778), .B(n20779), .Z(n20743) );
  NAND U29281 ( .A(n20780), .B(n20781), .Z(n20779) );
  NAND U29282 ( .A(n20782), .B(n20783), .Z(n20778) );
  AND U29283 ( .A(n20784), .B(n20785), .Z(n20739) );
  NAND U29284 ( .A(n20786), .B(n20787), .Z(n20785) );
  NAND U29285 ( .A(n20788), .B(n20789), .Z(n20784) );
  AND U29286 ( .A(n20790), .B(n20791), .Z(n20741) );
  NAND U29287 ( .A(n20792), .B(n20793), .Z(n20735) );
  XNOR U29288 ( .A(n20718), .B(n20794), .Z(n20732) );
  XNOR U29289 ( .A(n20722), .B(n20720), .Z(n20794) );
  XOR U29290 ( .A(n20728), .B(n20795), .Z(n20720) );
  XNOR U29291 ( .A(n20725), .B(n20729), .Z(n20795) );
  AND U29292 ( .A(n20796), .B(n20797), .Z(n20729) );
  NAND U29293 ( .A(n20798), .B(n20799), .Z(n20797) );
  NAND U29294 ( .A(n20800), .B(n20801), .Z(n20796) );
  AND U29295 ( .A(n20802), .B(n20803), .Z(n20725) );
  NAND U29296 ( .A(n20804), .B(n20805), .Z(n20803) );
  NAND U29297 ( .A(n20806), .B(n20807), .Z(n20802) );
  NANDN U29298 ( .A(n20808), .B(n20809), .Z(n20728) );
  ANDN U29299 ( .B(n20810), .A(n20811), .Z(n20722) );
  XNOR U29300 ( .A(n20713), .B(n20812), .Z(n20718) );
  XNOR U29301 ( .A(n20711), .B(n20715), .Z(n20812) );
  AND U29302 ( .A(n20813), .B(n20814), .Z(n20715) );
  NAND U29303 ( .A(n20815), .B(n20816), .Z(n20814) );
  NAND U29304 ( .A(n20817), .B(n20818), .Z(n20813) );
  AND U29305 ( .A(n20819), .B(n20820), .Z(n20711) );
  NAND U29306 ( .A(n20821), .B(n20822), .Z(n20820) );
  NAND U29307 ( .A(n20823), .B(n20824), .Z(n20819) );
  AND U29308 ( .A(n20825), .B(n20826), .Z(n20713) );
  XOR U29309 ( .A(n20793), .B(n20792), .Z(N63543) );
  XNOR U29310 ( .A(n20810), .B(n20811), .Z(n20792) );
  XNOR U29311 ( .A(n20825), .B(n20826), .Z(n20811) );
  XOR U29312 ( .A(n20822), .B(n20821), .Z(n20826) );
  XOR U29313 ( .A(y[5460]), .B(x[5460]), .Z(n20821) );
  XOR U29314 ( .A(n20824), .B(n20823), .Z(n20822) );
  XOR U29315 ( .A(y[5462]), .B(x[5462]), .Z(n20823) );
  XOR U29316 ( .A(y[5461]), .B(x[5461]), .Z(n20824) );
  XOR U29317 ( .A(n20816), .B(n20815), .Z(n20825) );
  XOR U29318 ( .A(n20818), .B(n20817), .Z(n20815) );
  XOR U29319 ( .A(y[5459]), .B(x[5459]), .Z(n20817) );
  XOR U29320 ( .A(y[5458]), .B(x[5458]), .Z(n20818) );
  XOR U29321 ( .A(y[5457]), .B(x[5457]), .Z(n20816) );
  XNOR U29322 ( .A(n20809), .B(n20808), .Z(n20810) );
  XNOR U29323 ( .A(n20805), .B(n20804), .Z(n20808) );
  XOR U29324 ( .A(n20807), .B(n20806), .Z(n20804) );
  XOR U29325 ( .A(y[5456]), .B(x[5456]), .Z(n20806) );
  XOR U29326 ( .A(y[5455]), .B(x[5455]), .Z(n20807) );
  XOR U29327 ( .A(y[5454]), .B(x[5454]), .Z(n20805) );
  XOR U29328 ( .A(n20799), .B(n20798), .Z(n20809) );
  XOR U29329 ( .A(n20801), .B(n20800), .Z(n20798) );
  XOR U29330 ( .A(y[5453]), .B(x[5453]), .Z(n20800) );
  XOR U29331 ( .A(y[5452]), .B(x[5452]), .Z(n20801) );
  XOR U29332 ( .A(y[5451]), .B(x[5451]), .Z(n20799) );
  XNOR U29333 ( .A(n20775), .B(n20776), .Z(n20793) );
  XNOR U29334 ( .A(n20790), .B(n20791), .Z(n20776) );
  XOR U29335 ( .A(n20787), .B(n20786), .Z(n20791) );
  XOR U29336 ( .A(y[5448]), .B(x[5448]), .Z(n20786) );
  XOR U29337 ( .A(n20789), .B(n20788), .Z(n20787) );
  XOR U29338 ( .A(y[5450]), .B(x[5450]), .Z(n20788) );
  XOR U29339 ( .A(y[5449]), .B(x[5449]), .Z(n20789) );
  XOR U29340 ( .A(n20781), .B(n20780), .Z(n20790) );
  XOR U29341 ( .A(n20783), .B(n20782), .Z(n20780) );
  XOR U29342 ( .A(y[5447]), .B(x[5447]), .Z(n20782) );
  XOR U29343 ( .A(y[5446]), .B(x[5446]), .Z(n20783) );
  XOR U29344 ( .A(y[5445]), .B(x[5445]), .Z(n20781) );
  XNOR U29345 ( .A(n20774), .B(n20773), .Z(n20775) );
  XNOR U29346 ( .A(n20770), .B(n20769), .Z(n20773) );
  XOR U29347 ( .A(n20772), .B(n20771), .Z(n20769) );
  XOR U29348 ( .A(y[5444]), .B(x[5444]), .Z(n20771) );
  XOR U29349 ( .A(y[5443]), .B(x[5443]), .Z(n20772) );
  XOR U29350 ( .A(y[5442]), .B(x[5442]), .Z(n20770) );
  XOR U29351 ( .A(n20764), .B(n20763), .Z(n20774) );
  XOR U29352 ( .A(n20766), .B(n20765), .Z(n20763) );
  XOR U29353 ( .A(y[5441]), .B(x[5441]), .Z(n20765) );
  XOR U29354 ( .A(y[5440]), .B(x[5440]), .Z(n20766) );
  XOR U29355 ( .A(y[5439]), .B(x[5439]), .Z(n20764) );
  NAND U29356 ( .A(n20827), .B(n20828), .Z(N63534) );
  NAND U29357 ( .A(n20829), .B(n20830), .Z(n20828) );
  NANDN U29358 ( .A(n20831), .B(n20832), .Z(n20830) );
  NANDN U29359 ( .A(n20832), .B(n20831), .Z(n20827) );
  XOR U29360 ( .A(n20831), .B(n20833), .Z(N63533) );
  XNOR U29361 ( .A(n20829), .B(n20832), .Z(n20833) );
  NAND U29362 ( .A(n20834), .B(n20835), .Z(n20832) );
  NAND U29363 ( .A(n20836), .B(n20837), .Z(n20835) );
  NANDN U29364 ( .A(n20838), .B(n20839), .Z(n20837) );
  NANDN U29365 ( .A(n20839), .B(n20838), .Z(n20834) );
  AND U29366 ( .A(n20840), .B(n20841), .Z(n20829) );
  NAND U29367 ( .A(n20842), .B(n20843), .Z(n20841) );
  NANDN U29368 ( .A(n20844), .B(n20845), .Z(n20843) );
  NANDN U29369 ( .A(n20845), .B(n20844), .Z(n20840) );
  IV U29370 ( .A(n20846), .Z(n20845) );
  AND U29371 ( .A(n20847), .B(n20848), .Z(n20831) );
  NAND U29372 ( .A(n20849), .B(n20850), .Z(n20848) );
  NANDN U29373 ( .A(n20851), .B(n20852), .Z(n20850) );
  NANDN U29374 ( .A(n20852), .B(n20851), .Z(n20847) );
  XOR U29375 ( .A(n20844), .B(n20853), .Z(N63532) );
  XNOR U29376 ( .A(n20842), .B(n20846), .Z(n20853) );
  XOR U29377 ( .A(n20839), .B(n20854), .Z(n20846) );
  XNOR U29378 ( .A(n20836), .B(n20838), .Z(n20854) );
  AND U29379 ( .A(n20855), .B(n20856), .Z(n20838) );
  NANDN U29380 ( .A(n20857), .B(n20858), .Z(n20856) );
  OR U29381 ( .A(n20859), .B(n20860), .Z(n20858) );
  IV U29382 ( .A(n20861), .Z(n20860) );
  NANDN U29383 ( .A(n20861), .B(n20859), .Z(n20855) );
  AND U29384 ( .A(n20862), .B(n20863), .Z(n20836) );
  NAND U29385 ( .A(n20864), .B(n20865), .Z(n20863) );
  NANDN U29386 ( .A(n20866), .B(n20867), .Z(n20865) );
  NANDN U29387 ( .A(n20867), .B(n20866), .Z(n20862) );
  IV U29388 ( .A(n20868), .Z(n20867) );
  NAND U29389 ( .A(n20869), .B(n20870), .Z(n20839) );
  NANDN U29390 ( .A(n20871), .B(n20872), .Z(n20870) );
  NANDN U29391 ( .A(n20873), .B(n20874), .Z(n20872) );
  NANDN U29392 ( .A(n20874), .B(n20873), .Z(n20869) );
  IV U29393 ( .A(n20875), .Z(n20873) );
  AND U29394 ( .A(n20876), .B(n20877), .Z(n20842) );
  NAND U29395 ( .A(n20878), .B(n20879), .Z(n20877) );
  NANDN U29396 ( .A(n20880), .B(n20881), .Z(n20879) );
  NANDN U29397 ( .A(n20881), .B(n20880), .Z(n20876) );
  XOR U29398 ( .A(n20852), .B(n20882), .Z(n20844) );
  XNOR U29399 ( .A(n20849), .B(n20851), .Z(n20882) );
  AND U29400 ( .A(n20883), .B(n20884), .Z(n20851) );
  NANDN U29401 ( .A(n20885), .B(n20886), .Z(n20884) );
  OR U29402 ( .A(n20887), .B(n20888), .Z(n20886) );
  IV U29403 ( .A(n20889), .Z(n20888) );
  NANDN U29404 ( .A(n20889), .B(n20887), .Z(n20883) );
  AND U29405 ( .A(n20890), .B(n20891), .Z(n20849) );
  NAND U29406 ( .A(n20892), .B(n20893), .Z(n20891) );
  NANDN U29407 ( .A(n20894), .B(n20895), .Z(n20893) );
  NANDN U29408 ( .A(n20895), .B(n20894), .Z(n20890) );
  IV U29409 ( .A(n20896), .Z(n20895) );
  NAND U29410 ( .A(n20897), .B(n20898), .Z(n20852) );
  NANDN U29411 ( .A(n20899), .B(n20900), .Z(n20898) );
  NANDN U29412 ( .A(n20901), .B(n20902), .Z(n20900) );
  NANDN U29413 ( .A(n20902), .B(n20901), .Z(n20897) );
  IV U29414 ( .A(n20903), .Z(n20901) );
  XOR U29415 ( .A(n20878), .B(n20904), .Z(N63531) );
  XNOR U29416 ( .A(n20881), .B(n20880), .Z(n20904) );
  XNOR U29417 ( .A(n20892), .B(n20905), .Z(n20880) );
  XNOR U29418 ( .A(n20896), .B(n20894), .Z(n20905) );
  XOR U29419 ( .A(n20902), .B(n20906), .Z(n20894) );
  XNOR U29420 ( .A(n20899), .B(n20903), .Z(n20906) );
  AND U29421 ( .A(n20907), .B(n20908), .Z(n20903) );
  NAND U29422 ( .A(n20909), .B(n20910), .Z(n20908) );
  NAND U29423 ( .A(n20911), .B(n20912), .Z(n20907) );
  AND U29424 ( .A(n20913), .B(n20914), .Z(n20899) );
  NAND U29425 ( .A(n20915), .B(n20916), .Z(n20914) );
  NAND U29426 ( .A(n20917), .B(n20918), .Z(n20913) );
  NANDN U29427 ( .A(n20919), .B(n20920), .Z(n20902) );
  ANDN U29428 ( .B(n20921), .A(n20922), .Z(n20896) );
  XNOR U29429 ( .A(n20887), .B(n20923), .Z(n20892) );
  XNOR U29430 ( .A(n20885), .B(n20889), .Z(n20923) );
  AND U29431 ( .A(n20924), .B(n20925), .Z(n20889) );
  NAND U29432 ( .A(n20926), .B(n20927), .Z(n20925) );
  NAND U29433 ( .A(n20928), .B(n20929), .Z(n20924) );
  AND U29434 ( .A(n20930), .B(n20931), .Z(n20885) );
  NAND U29435 ( .A(n20932), .B(n20933), .Z(n20931) );
  NAND U29436 ( .A(n20934), .B(n20935), .Z(n20930) );
  AND U29437 ( .A(n20936), .B(n20937), .Z(n20887) );
  NAND U29438 ( .A(n20938), .B(n20939), .Z(n20881) );
  XNOR U29439 ( .A(n20864), .B(n20940), .Z(n20878) );
  XNOR U29440 ( .A(n20868), .B(n20866), .Z(n20940) );
  XOR U29441 ( .A(n20874), .B(n20941), .Z(n20866) );
  XNOR U29442 ( .A(n20871), .B(n20875), .Z(n20941) );
  AND U29443 ( .A(n20942), .B(n20943), .Z(n20875) );
  NAND U29444 ( .A(n20944), .B(n20945), .Z(n20943) );
  NAND U29445 ( .A(n20946), .B(n20947), .Z(n20942) );
  AND U29446 ( .A(n20948), .B(n20949), .Z(n20871) );
  NAND U29447 ( .A(n20950), .B(n20951), .Z(n20949) );
  NAND U29448 ( .A(n20952), .B(n20953), .Z(n20948) );
  NANDN U29449 ( .A(n20954), .B(n20955), .Z(n20874) );
  ANDN U29450 ( .B(n20956), .A(n20957), .Z(n20868) );
  XNOR U29451 ( .A(n20859), .B(n20958), .Z(n20864) );
  XNOR U29452 ( .A(n20857), .B(n20861), .Z(n20958) );
  AND U29453 ( .A(n20959), .B(n20960), .Z(n20861) );
  NAND U29454 ( .A(n20961), .B(n20962), .Z(n20960) );
  NAND U29455 ( .A(n20963), .B(n20964), .Z(n20959) );
  AND U29456 ( .A(n20965), .B(n20966), .Z(n20857) );
  NAND U29457 ( .A(n20967), .B(n20968), .Z(n20966) );
  NAND U29458 ( .A(n20969), .B(n20970), .Z(n20965) );
  AND U29459 ( .A(n20971), .B(n20972), .Z(n20859) );
  XOR U29460 ( .A(n20939), .B(n20938), .Z(N63530) );
  XNOR U29461 ( .A(n20956), .B(n20957), .Z(n20938) );
  XNOR U29462 ( .A(n20971), .B(n20972), .Z(n20957) );
  XOR U29463 ( .A(n20968), .B(n20967), .Z(n20972) );
  XOR U29464 ( .A(y[5436]), .B(x[5436]), .Z(n20967) );
  XOR U29465 ( .A(n20970), .B(n20969), .Z(n20968) );
  XOR U29466 ( .A(y[5438]), .B(x[5438]), .Z(n20969) );
  XOR U29467 ( .A(y[5437]), .B(x[5437]), .Z(n20970) );
  XOR U29468 ( .A(n20962), .B(n20961), .Z(n20971) );
  XOR U29469 ( .A(n20964), .B(n20963), .Z(n20961) );
  XOR U29470 ( .A(y[5435]), .B(x[5435]), .Z(n20963) );
  XOR U29471 ( .A(y[5434]), .B(x[5434]), .Z(n20964) );
  XOR U29472 ( .A(y[5433]), .B(x[5433]), .Z(n20962) );
  XNOR U29473 ( .A(n20955), .B(n20954), .Z(n20956) );
  XNOR U29474 ( .A(n20951), .B(n20950), .Z(n20954) );
  XOR U29475 ( .A(n20953), .B(n20952), .Z(n20950) );
  XOR U29476 ( .A(y[5432]), .B(x[5432]), .Z(n20952) );
  XOR U29477 ( .A(y[5431]), .B(x[5431]), .Z(n20953) );
  XOR U29478 ( .A(y[5430]), .B(x[5430]), .Z(n20951) );
  XOR U29479 ( .A(n20945), .B(n20944), .Z(n20955) );
  XOR U29480 ( .A(n20947), .B(n20946), .Z(n20944) );
  XOR U29481 ( .A(y[5429]), .B(x[5429]), .Z(n20946) );
  XOR U29482 ( .A(y[5428]), .B(x[5428]), .Z(n20947) );
  XOR U29483 ( .A(y[5427]), .B(x[5427]), .Z(n20945) );
  XNOR U29484 ( .A(n20921), .B(n20922), .Z(n20939) );
  XNOR U29485 ( .A(n20936), .B(n20937), .Z(n20922) );
  XOR U29486 ( .A(n20933), .B(n20932), .Z(n20937) );
  XOR U29487 ( .A(y[5424]), .B(x[5424]), .Z(n20932) );
  XOR U29488 ( .A(n20935), .B(n20934), .Z(n20933) );
  XOR U29489 ( .A(y[5426]), .B(x[5426]), .Z(n20934) );
  XOR U29490 ( .A(y[5425]), .B(x[5425]), .Z(n20935) );
  XOR U29491 ( .A(n20927), .B(n20926), .Z(n20936) );
  XOR U29492 ( .A(n20929), .B(n20928), .Z(n20926) );
  XOR U29493 ( .A(y[5423]), .B(x[5423]), .Z(n20928) );
  XOR U29494 ( .A(y[5422]), .B(x[5422]), .Z(n20929) );
  XOR U29495 ( .A(y[5421]), .B(x[5421]), .Z(n20927) );
  XNOR U29496 ( .A(n20920), .B(n20919), .Z(n20921) );
  XNOR U29497 ( .A(n20916), .B(n20915), .Z(n20919) );
  XOR U29498 ( .A(n20918), .B(n20917), .Z(n20915) );
  XOR U29499 ( .A(y[5420]), .B(x[5420]), .Z(n20917) );
  XOR U29500 ( .A(y[5419]), .B(x[5419]), .Z(n20918) );
  XOR U29501 ( .A(y[5418]), .B(x[5418]), .Z(n20916) );
  XOR U29502 ( .A(n20910), .B(n20909), .Z(n20920) );
  XOR U29503 ( .A(n20912), .B(n20911), .Z(n20909) );
  XOR U29504 ( .A(y[5417]), .B(x[5417]), .Z(n20911) );
  XOR U29505 ( .A(y[5416]), .B(x[5416]), .Z(n20912) );
  XOR U29506 ( .A(y[5415]), .B(x[5415]), .Z(n20910) );
  NAND U29507 ( .A(n20973), .B(n20974), .Z(N63521) );
  NAND U29508 ( .A(n20975), .B(n20976), .Z(n20974) );
  NANDN U29509 ( .A(n20977), .B(n20978), .Z(n20976) );
  NANDN U29510 ( .A(n20978), .B(n20977), .Z(n20973) );
  XOR U29511 ( .A(n20977), .B(n20979), .Z(N63520) );
  XNOR U29512 ( .A(n20975), .B(n20978), .Z(n20979) );
  NAND U29513 ( .A(n20980), .B(n20981), .Z(n20978) );
  NAND U29514 ( .A(n20982), .B(n20983), .Z(n20981) );
  NANDN U29515 ( .A(n20984), .B(n20985), .Z(n20983) );
  NANDN U29516 ( .A(n20985), .B(n20984), .Z(n20980) );
  AND U29517 ( .A(n20986), .B(n20987), .Z(n20975) );
  NAND U29518 ( .A(n20988), .B(n20989), .Z(n20987) );
  NANDN U29519 ( .A(n20990), .B(n20991), .Z(n20989) );
  NANDN U29520 ( .A(n20991), .B(n20990), .Z(n20986) );
  IV U29521 ( .A(n20992), .Z(n20991) );
  AND U29522 ( .A(n20993), .B(n20994), .Z(n20977) );
  NAND U29523 ( .A(n20995), .B(n20996), .Z(n20994) );
  NANDN U29524 ( .A(n20997), .B(n20998), .Z(n20996) );
  NANDN U29525 ( .A(n20998), .B(n20997), .Z(n20993) );
  XOR U29526 ( .A(n20990), .B(n20999), .Z(N63519) );
  XNOR U29527 ( .A(n20988), .B(n20992), .Z(n20999) );
  XOR U29528 ( .A(n20985), .B(n21000), .Z(n20992) );
  XNOR U29529 ( .A(n20982), .B(n20984), .Z(n21000) );
  AND U29530 ( .A(n21001), .B(n21002), .Z(n20984) );
  NANDN U29531 ( .A(n21003), .B(n21004), .Z(n21002) );
  OR U29532 ( .A(n21005), .B(n21006), .Z(n21004) );
  IV U29533 ( .A(n21007), .Z(n21006) );
  NANDN U29534 ( .A(n21007), .B(n21005), .Z(n21001) );
  AND U29535 ( .A(n21008), .B(n21009), .Z(n20982) );
  NAND U29536 ( .A(n21010), .B(n21011), .Z(n21009) );
  NANDN U29537 ( .A(n21012), .B(n21013), .Z(n21011) );
  NANDN U29538 ( .A(n21013), .B(n21012), .Z(n21008) );
  IV U29539 ( .A(n21014), .Z(n21013) );
  NAND U29540 ( .A(n21015), .B(n21016), .Z(n20985) );
  NANDN U29541 ( .A(n21017), .B(n21018), .Z(n21016) );
  NANDN U29542 ( .A(n21019), .B(n21020), .Z(n21018) );
  NANDN U29543 ( .A(n21020), .B(n21019), .Z(n21015) );
  IV U29544 ( .A(n21021), .Z(n21019) );
  AND U29545 ( .A(n21022), .B(n21023), .Z(n20988) );
  NAND U29546 ( .A(n21024), .B(n21025), .Z(n21023) );
  NANDN U29547 ( .A(n21026), .B(n21027), .Z(n21025) );
  NANDN U29548 ( .A(n21027), .B(n21026), .Z(n21022) );
  XOR U29549 ( .A(n20998), .B(n21028), .Z(n20990) );
  XNOR U29550 ( .A(n20995), .B(n20997), .Z(n21028) );
  AND U29551 ( .A(n21029), .B(n21030), .Z(n20997) );
  NANDN U29552 ( .A(n21031), .B(n21032), .Z(n21030) );
  OR U29553 ( .A(n21033), .B(n21034), .Z(n21032) );
  IV U29554 ( .A(n21035), .Z(n21034) );
  NANDN U29555 ( .A(n21035), .B(n21033), .Z(n21029) );
  AND U29556 ( .A(n21036), .B(n21037), .Z(n20995) );
  NAND U29557 ( .A(n21038), .B(n21039), .Z(n21037) );
  NANDN U29558 ( .A(n21040), .B(n21041), .Z(n21039) );
  NANDN U29559 ( .A(n21041), .B(n21040), .Z(n21036) );
  IV U29560 ( .A(n21042), .Z(n21041) );
  NAND U29561 ( .A(n21043), .B(n21044), .Z(n20998) );
  NANDN U29562 ( .A(n21045), .B(n21046), .Z(n21044) );
  NANDN U29563 ( .A(n21047), .B(n21048), .Z(n21046) );
  NANDN U29564 ( .A(n21048), .B(n21047), .Z(n21043) );
  IV U29565 ( .A(n21049), .Z(n21047) );
  XOR U29566 ( .A(n21024), .B(n21050), .Z(N63518) );
  XNOR U29567 ( .A(n21027), .B(n21026), .Z(n21050) );
  XNOR U29568 ( .A(n21038), .B(n21051), .Z(n21026) );
  XNOR U29569 ( .A(n21042), .B(n21040), .Z(n21051) );
  XOR U29570 ( .A(n21048), .B(n21052), .Z(n21040) );
  XNOR U29571 ( .A(n21045), .B(n21049), .Z(n21052) );
  AND U29572 ( .A(n21053), .B(n21054), .Z(n21049) );
  NAND U29573 ( .A(n21055), .B(n21056), .Z(n21054) );
  NAND U29574 ( .A(n21057), .B(n21058), .Z(n21053) );
  AND U29575 ( .A(n21059), .B(n21060), .Z(n21045) );
  NAND U29576 ( .A(n21061), .B(n21062), .Z(n21060) );
  NAND U29577 ( .A(n21063), .B(n21064), .Z(n21059) );
  NANDN U29578 ( .A(n21065), .B(n21066), .Z(n21048) );
  ANDN U29579 ( .B(n21067), .A(n21068), .Z(n21042) );
  XNOR U29580 ( .A(n21033), .B(n21069), .Z(n21038) );
  XNOR U29581 ( .A(n21031), .B(n21035), .Z(n21069) );
  AND U29582 ( .A(n21070), .B(n21071), .Z(n21035) );
  NAND U29583 ( .A(n21072), .B(n21073), .Z(n21071) );
  NAND U29584 ( .A(n21074), .B(n21075), .Z(n21070) );
  AND U29585 ( .A(n21076), .B(n21077), .Z(n21031) );
  NAND U29586 ( .A(n21078), .B(n21079), .Z(n21077) );
  NAND U29587 ( .A(n21080), .B(n21081), .Z(n21076) );
  AND U29588 ( .A(n21082), .B(n21083), .Z(n21033) );
  NAND U29589 ( .A(n21084), .B(n21085), .Z(n21027) );
  XNOR U29590 ( .A(n21010), .B(n21086), .Z(n21024) );
  XNOR U29591 ( .A(n21014), .B(n21012), .Z(n21086) );
  XOR U29592 ( .A(n21020), .B(n21087), .Z(n21012) );
  XNOR U29593 ( .A(n21017), .B(n21021), .Z(n21087) );
  AND U29594 ( .A(n21088), .B(n21089), .Z(n21021) );
  NAND U29595 ( .A(n21090), .B(n21091), .Z(n21089) );
  NAND U29596 ( .A(n21092), .B(n21093), .Z(n21088) );
  AND U29597 ( .A(n21094), .B(n21095), .Z(n21017) );
  NAND U29598 ( .A(n21096), .B(n21097), .Z(n21095) );
  NAND U29599 ( .A(n21098), .B(n21099), .Z(n21094) );
  NANDN U29600 ( .A(n21100), .B(n21101), .Z(n21020) );
  ANDN U29601 ( .B(n21102), .A(n21103), .Z(n21014) );
  XNOR U29602 ( .A(n21005), .B(n21104), .Z(n21010) );
  XNOR U29603 ( .A(n21003), .B(n21007), .Z(n21104) );
  AND U29604 ( .A(n21105), .B(n21106), .Z(n21007) );
  NAND U29605 ( .A(n21107), .B(n21108), .Z(n21106) );
  NAND U29606 ( .A(n21109), .B(n21110), .Z(n21105) );
  AND U29607 ( .A(n21111), .B(n21112), .Z(n21003) );
  NAND U29608 ( .A(n21113), .B(n21114), .Z(n21112) );
  NAND U29609 ( .A(n21115), .B(n21116), .Z(n21111) );
  AND U29610 ( .A(n21117), .B(n21118), .Z(n21005) );
  XOR U29611 ( .A(n21085), .B(n21084), .Z(N63517) );
  XNOR U29612 ( .A(n21102), .B(n21103), .Z(n21084) );
  XNOR U29613 ( .A(n21117), .B(n21118), .Z(n21103) );
  XOR U29614 ( .A(n21114), .B(n21113), .Z(n21118) );
  XOR U29615 ( .A(y[5412]), .B(x[5412]), .Z(n21113) );
  XOR U29616 ( .A(n21116), .B(n21115), .Z(n21114) );
  XOR U29617 ( .A(y[5414]), .B(x[5414]), .Z(n21115) );
  XOR U29618 ( .A(y[5413]), .B(x[5413]), .Z(n21116) );
  XOR U29619 ( .A(n21108), .B(n21107), .Z(n21117) );
  XOR U29620 ( .A(n21110), .B(n21109), .Z(n21107) );
  XOR U29621 ( .A(y[5411]), .B(x[5411]), .Z(n21109) );
  XOR U29622 ( .A(y[5410]), .B(x[5410]), .Z(n21110) );
  XOR U29623 ( .A(y[5409]), .B(x[5409]), .Z(n21108) );
  XNOR U29624 ( .A(n21101), .B(n21100), .Z(n21102) );
  XNOR U29625 ( .A(n21097), .B(n21096), .Z(n21100) );
  XOR U29626 ( .A(n21099), .B(n21098), .Z(n21096) );
  XOR U29627 ( .A(y[5408]), .B(x[5408]), .Z(n21098) );
  XOR U29628 ( .A(y[5407]), .B(x[5407]), .Z(n21099) );
  XOR U29629 ( .A(y[5406]), .B(x[5406]), .Z(n21097) );
  XOR U29630 ( .A(n21091), .B(n21090), .Z(n21101) );
  XOR U29631 ( .A(n21093), .B(n21092), .Z(n21090) );
  XOR U29632 ( .A(y[5405]), .B(x[5405]), .Z(n21092) );
  XOR U29633 ( .A(y[5404]), .B(x[5404]), .Z(n21093) );
  XOR U29634 ( .A(y[5403]), .B(x[5403]), .Z(n21091) );
  XNOR U29635 ( .A(n21067), .B(n21068), .Z(n21085) );
  XNOR U29636 ( .A(n21082), .B(n21083), .Z(n21068) );
  XOR U29637 ( .A(n21079), .B(n21078), .Z(n21083) );
  XOR U29638 ( .A(y[5400]), .B(x[5400]), .Z(n21078) );
  XOR U29639 ( .A(n21081), .B(n21080), .Z(n21079) );
  XOR U29640 ( .A(y[5402]), .B(x[5402]), .Z(n21080) );
  XOR U29641 ( .A(y[5401]), .B(x[5401]), .Z(n21081) );
  XOR U29642 ( .A(n21073), .B(n21072), .Z(n21082) );
  XOR U29643 ( .A(n21075), .B(n21074), .Z(n21072) );
  XOR U29644 ( .A(y[5399]), .B(x[5399]), .Z(n21074) );
  XOR U29645 ( .A(y[5398]), .B(x[5398]), .Z(n21075) );
  XOR U29646 ( .A(y[5397]), .B(x[5397]), .Z(n21073) );
  XNOR U29647 ( .A(n21066), .B(n21065), .Z(n21067) );
  XNOR U29648 ( .A(n21062), .B(n21061), .Z(n21065) );
  XOR U29649 ( .A(n21064), .B(n21063), .Z(n21061) );
  XOR U29650 ( .A(y[5396]), .B(x[5396]), .Z(n21063) );
  XOR U29651 ( .A(y[5395]), .B(x[5395]), .Z(n21064) );
  XOR U29652 ( .A(y[5394]), .B(x[5394]), .Z(n21062) );
  XOR U29653 ( .A(n21056), .B(n21055), .Z(n21066) );
  XOR U29654 ( .A(n21058), .B(n21057), .Z(n21055) );
  XOR U29655 ( .A(y[5393]), .B(x[5393]), .Z(n21057) );
  XOR U29656 ( .A(y[5392]), .B(x[5392]), .Z(n21058) );
  XOR U29657 ( .A(y[5391]), .B(x[5391]), .Z(n21056) );
  NAND U29658 ( .A(n21119), .B(n21120), .Z(N63508) );
  NAND U29659 ( .A(n21121), .B(n21122), .Z(n21120) );
  NANDN U29660 ( .A(n21123), .B(n21124), .Z(n21122) );
  NANDN U29661 ( .A(n21124), .B(n21123), .Z(n21119) );
  XOR U29662 ( .A(n21123), .B(n21125), .Z(N63507) );
  XNOR U29663 ( .A(n21121), .B(n21124), .Z(n21125) );
  NAND U29664 ( .A(n21126), .B(n21127), .Z(n21124) );
  NAND U29665 ( .A(n21128), .B(n21129), .Z(n21127) );
  NANDN U29666 ( .A(n21130), .B(n21131), .Z(n21129) );
  NANDN U29667 ( .A(n21131), .B(n21130), .Z(n21126) );
  AND U29668 ( .A(n21132), .B(n21133), .Z(n21121) );
  NAND U29669 ( .A(n21134), .B(n21135), .Z(n21133) );
  NANDN U29670 ( .A(n21136), .B(n21137), .Z(n21135) );
  NANDN U29671 ( .A(n21137), .B(n21136), .Z(n21132) );
  IV U29672 ( .A(n21138), .Z(n21137) );
  AND U29673 ( .A(n21139), .B(n21140), .Z(n21123) );
  NAND U29674 ( .A(n21141), .B(n21142), .Z(n21140) );
  NANDN U29675 ( .A(n21143), .B(n21144), .Z(n21142) );
  NANDN U29676 ( .A(n21144), .B(n21143), .Z(n21139) );
  XOR U29677 ( .A(n21136), .B(n21145), .Z(N63506) );
  XNOR U29678 ( .A(n21134), .B(n21138), .Z(n21145) );
  XOR U29679 ( .A(n21131), .B(n21146), .Z(n21138) );
  XNOR U29680 ( .A(n21128), .B(n21130), .Z(n21146) );
  AND U29681 ( .A(n21147), .B(n21148), .Z(n21130) );
  NANDN U29682 ( .A(n21149), .B(n21150), .Z(n21148) );
  OR U29683 ( .A(n21151), .B(n21152), .Z(n21150) );
  IV U29684 ( .A(n21153), .Z(n21152) );
  NANDN U29685 ( .A(n21153), .B(n21151), .Z(n21147) );
  AND U29686 ( .A(n21154), .B(n21155), .Z(n21128) );
  NAND U29687 ( .A(n21156), .B(n21157), .Z(n21155) );
  NANDN U29688 ( .A(n21158), .B(n21159), .Z(n21157) );
  NANDN U29689 ( .A(n21159), .B(n21158), .Z(n21154) );
  IV U29690 ( .A(n21160), .Z(n21159) );
  NAND U29691 ( .A(n21161), .B(n21162), .Z(n21131) );
  NANDN U29692 ( .A(n21163), .B(n21164), .Z(n21162) );
  NANDN U29693 ( .A(n21165), .B(n21166), .Z(n21164) );
  NANDN U29694 ( .A(n21166), .B(n21165), .Z(n21161) );
  IV U29695 ( .A(n21167), .Z(n21165) );
  AND U29696 ( .A(n21168), .B(n21169), .Z(n21134) );
  NAND U29697 ( .A(n21170), .B(n21171), .Z(n21169) );
  NANDN U29698 ( .A(n21172), .B(n21173), .Z(n21171) );
  NANDN U29699 ( .A(n21173), .B(n21172), .Z(n21168) );
  XOR U29700 ( .A(n21144), .B(n21174), .Z(n21136) );
  XNOR U29701 ( .A(n21141), .B(n21143), .Z(n21174) );
  AND U29702 ( .A(n21175), .B(n21176), .Z(n21143) );
  NANDN U29703 ( .A(n21177), .B(n21178), .Z(n21176) );
  OR U29704 ( .A(n21179), .B(n21180), .Z(n21178) );
  IV U29705 ( .A(n21181), .Z(n21180) );
  NANDN U29706 ( .A(n21181), .B(n21179), .Z(n21175) );
  AND U29707 ( .A(n21182), .B(n21183), .Z(n21141) );
  NAND U29708 ( .A(n21184), .B(n21185), .Z(n21183) );
  NANDN U29709 ( .A(n21186), .B(n21187), .Z(n21185) );
  NANDN U29710 ( .A(n21187), .B(n21186), .Z(n21182) );
  IV U29711 ( .A(n21188), .Z(n21187) );
  NAND U29712 ( .A(n21189), .B(n21190), .Z(n21144) );
  NANDN U29713 ( .A(n21191), .B(n21192), .Z(n21190) );
  NANDN U29714 ( .A(n21193), .B(n21194), .Z(n21192) );
  NANDN U29715 ( .A(n21194), .B(n21193), .Z(n21189) );
  IV U29716 ( .A(n21195), .Z(n21193) );
  XOR U29717 ( .A(n21170), .B(n21196), .Z(N63505) );
  XNOR U29718 ( .A(n21173), .B(n21172), .Z(n21196) );
  XNOR U29719 ( .A(n21184), .B(n21197), .Z(n21172) );
  XNOR U29720 ( .A(n21188), .B(n21186), .Z(n21197) );
  XOR U29721 ( .A(n21194), .B(n21198), .Z(n21186) );
  XNOR U29722 ( .A(n21191), .B(n21195), .Z(n21198) );
  AND U29723 ( .A(n21199), .B(n21200), .Z(n21195) );
  NAND U29724 ( .A(n21201), .B(n21202), .Z(n21200) );
  NAND U29725 ( .A(n21203), .B(n21204), .Z(n21199) );
  AND U29726 ( .A(n21205), .B(n21206), .Z(n21191) );
  NAND U29727 ( .A(n21207), .B(n21208), .Z(n21206) );
  NAND U29728 ( .A(n21209), .B(n21210), .Z(n21205) );
  NANDN U29729 ( .A(n21211), .B(n21212), .Z(n21194) );
  ANDN U29730 ( .B(n21213), .A(n21214), .Z(n21188) );
  XNOR U29731 ( .A(n21179), .B(n21215), .Z(n21184) );
  XNOR U29732 ( .A(n21177), .B(n21181), .Z(n21215) );
  AND U29733 ( .A(n21216), .B(n21217), .Z(n21181) );
  NAND U29734 ( .A(n21218), .B(n21219), .Z(n21217) );
  NAND U29735 ( .A(n21220), .B(n21221), .Z(n21216) );
  AND U29736 ( .A(n21222), .B(n21223), .Z(n21177) );
  NAND U29737 ( .A(n21224), .B(n21225), .Z(n21223) );
  NAND U29738 ( .A(n21226), .B(n21227), .Z(n21222) );
  AND U29739 ( .A(n21228), .B(n21229), .Z(n21179) );
  NAND U29740 ( .A(n21230), .B(n21231), .Z(n21173) );
  XNOR U29741 ( .A(n21156), .B(n21232), .Z(n21170) );
  XNOR U29742 ( .A(n21160), .B(n21158), .Z(n21232) );
  XOR U29743 ( .A(n21166), .B(n21233), .Z(n21158) );
  XNOR U29744 ( .A(n21163), .B(n21167), .Z(n21233) );
  AND U29745 ( .A(n21234), .B(n21235), .Z(n21167) );
  NAND U29746 ( .A(n21236), .B(n21237), .Z(n21235) );
  NAND U29747 ( .A(n21238), .B(n21239), .Z(n21234) );
  AND U29748 ( .A(n21240), .B(n21241), .Z(n21163) );
  NAND U29749 ( .A(n21242), .B(n21243), .Z(n21241) );
  NAND U29750 ( .A(n21244), .B(n21245), .Z(n21240) );
  NANDN U29751 ( .A(n21246), .B(n21247), .Z(n21166) );
  ANDN U29752 ( .B(n21248), .A(n21249), .Z(n21160) );
  XNOR U29753 ( .A(n21151), .B(n21250), .Z(n21156) );
  XNOR U29754 ( .A(n21149), .B(n21153), .Z(n21250) );
  AND U29755 ( .A(n21251), .B(n21252), .Z(n21153) );
  NAND U29756 ( .A(n21253), .B(n21254), .Z(n21252) );
  NAND U29757 ( .A(n21255), .B(n21256), .Z(n21251) );
  AND U29758 ( .A(n21257), .B(n21258), .Z(n21149) );
  NAND U29759 ( .A(n21259), .B(n21260), .Z(n21258) );
  NAND U29760 ( .A(n21261), .B(n21262), .Z(n21257) );
  AND U29761 ( .A(n21263), .B(n21264), .Z(n21151) );
  XOR U29762 ( .A(n21231), .B(n21230), .Z(N63504) );
  XNOR U29763 ( .A(n21248), .B(n21249), .Z(n21230) );
  XNOR U29764 ( .A(n21263), .B(n21264), .Z(n21249) );
  XOR U29765 ( .A(n21260), .B(n21259), .Z(n21264) );
  XOR U29766 ( .A(y[5388]), .B(x[5388]), .Z(n21259) );
  XOR U29767 ( .A(n21262), .B(n21261), .Z(n21260) );
  XOR U29768 ( .A(y[5390]), .B(x[5390]), .Z(n21261) );
  XOR U29769 ( .A(y[5389]), .B(x[5389]), .Z(n21262) );
  XOR U29770 ( .A(n21254), .B(n21253), .Z(n21263) );
  XOR U29771 ( .A(n21256), .B(n21255), .Z(n21253) );
  XOR U29772 ( .A(y[5387]), .B(x[5387]), .Z(n21255) );
  XOR U29773 ( .A(y[5386]), .B(x[5386]), .Z(n21256) );
  XOR U29774 ( .A(y[5385]), .B(x[5385]), .Z(n21254) );
  XNOR U29775 ( .A(n21247), .B(n21246), .Z(n21248) );
  XNOR U29776 ( .A(n21243), .B(n21242), .Z(n21246) );
  XOR U29777 ( .A(n21245), .B(n21244), .Z(n21242) );
  XOR U29778 ( .A(y[5384]), .B(x[5384]), .Z(n21244) );
  XOR U29779 ( .A(y[5383]), .B(x[5383]), .Z(n21245) );
  XOR U29780 ( .A(y[5382]), .B(x[5382]), .Z(n21243) );
  XOR U29781 ( .A(n21237), .B(n21236), .Z(n21247) );
  XOR U29782 ( .A(n21239), .B(n21238), .Z(n21236) );
  XOR U29783 ( .A(y[5381]), .B(x[5381]), .Z(n21238) );
  XOR U29784 ( .A(y[5380]), .B(x[5380]), .Z(n21239) );
  XOR U29785 ( .A(y[5379]), .B(x[5379]), .Z(n21237) );
  XNOR U29786 ( .A(n21213), .B(n21214), .Z(n21231) );
  XNOR U29787 ( .A(n21228), .B(n21229), .Z(n21214) );
  XOR U29788 ( .A(n21225), .B(n21224), .Z(n21229) );
  XOR U29789 ( .A(y[5376]), .B(x[5376]), .Z(n21224) );
  XOR U29790 ( .A(n21227), .B(n21226), .Z(n21225) );
  XOR U29791 ( .A(y[5378]), .B(x[5378]), .Z(n21226) );
  XOR U29792 ( .A(y[5377]), .B(x[5377]), .Z(n21227) );
  XOR U29793 ( .A(n21219), .B(n21218), .Z(n21228) );
  XOR U29794 ( .A(n21221), .B(n21220), .Z(n21218) );
  XOR U29795 ( .A(y[5375]), .B(x[5375]), .Z(n21220) );
  XOR U29796 ( .A(y[5374]), .B(x[5374]), .Z(n21221) );
  XOR U29797 ( .A(y[5373]), .B(x[5373]), .Z(n21219) );
  XNOR U29798 ( .A(n21212), .B(n21211), .Z(n21213) );
  XNOR U29799 ( .A(n21208), .B(n21207), .Z(n21211) );
  XOR U29800 ( .A(n21210), .B(n21209), .Z(n21207) );
  XOR U29801 ( .A(y[5372]), .B(x[5372]), .Z(n21209) );
  XOR U29802 ( .A(y[5371]), .B(x[5371]), .Z(n21210) );
  XOR U29803 ( .A(y[5370]), .B(x[5370]), .Z(n21208) );
  XOR U29804 ( .A(n21202), .B(n21201), .Z(n21212) );
  XOR U29805 ( .A(n21204), .B(n21203), .Z(n21201) );
  XOR U29806 ( .A(y[5369]), .B(x[5369]), .Z(n21203) );
  XOR U29807 ( .A(y[5368]), .B(x[5368]), .Z(n21204) );
  XOR U29808 ( .A(y[5367]), .B(x[5367]), .Z(n21202) );
  NAND U29809 ( .A(n21265), .B(n21266), .Z(N63495) );
  NAND U29810 ( .A(n21267), .B(n21268), .Z(n21266) );
  NANDN U29811 ( .A(n21269), .B(n21270), .Z(n21268) );
  NANDN U29812 ( .A(n21270), .B(n21269), .Z(n21265) );
  XOR U29813 ( .A(n21269), .B(n21271), .Z(N63494) );
  XNOR U29814 ( .A(n21267), .B(n21270), .Z(n21271) );
  NAND U29815 ( .A(n21272), .B(n21273), .Z(n21270) );
  NAND U29816 ( .A(n21274), .B(n21275), .Z(n21273) );
  NANDN U29817 ( .A(n21276), .B(n21277), .Z(n21275) );
  NANDN U29818 ( .A(n21277), .B(n21276), .Z(n21272) );
  AND U29819 ( .A(n21278), .B(n21279), .Z(n21267) );
  NAND U29820 ( .A(n21280), .B(n21281), .Z(n21279) );
  NANDN U29821 ( .A(n21282), .B(n21283), .Z(n21281) );
  NANDN U29822 ( .A(n21283), .B(n21282), .Z(n21278) );
  IV U29823 ( .A(n21284), .Z(n21283) );
  AND U29824 ( .A(n21285), .B(n21286), .Z(n21269) );
  NAND U29825 ( .A(n21287), .B(n21288), .Z(n21286) );
  NANDN U29826 ( .A(n21289), .B(n21290), .Z(n21288) );
  NANDN U29827 ( .A(n21290), .B(n21289), .Z(n21285) );
  XOR U29828 ( .A(n21282), .B(n21291), .Z(N63493) );
  XNOR U29829 ( .A(n21280), .B(n21284), .Z(n21291) );
  XOR U29830 ( .A(n21277), .B(n21292), .Z(n21284) );
  XNOR U29831 ( .A(n21274), .B(n21276), .Z(n21292) );
  AND U29832 ( .A(n21293), .B(n21294), .Z(n21276) );
  NANDN U29833 ( .A(n21295), .B(n21296), .Z(n21294) );
  OR U29834 ( .A(n21297), .B(n21298), .Z(n21296) );
  IV U29835 ( .A(n21299), .Z(n21298) );
  NANDN U29836 ( .A(n21299), .B(n21297), .Z(n21293) );
  AND U29837 ( .A(n21300), .B(n21301), .Z(n21274) );
  NAND U29838 ( .A(n21302), .B(n21303), .Z(n21301) );
  NANDN U29839 ( .A(n21304), .B(n21305), .Z(n21303) );
  NANDN U29840 ( .A(n21305), .B(n21304), .Z(n21300) );
  IV U29841 ( .A(n21306), .Z(n21305) );
  NAND U29842 ( .A(n21307), .B(n21308), .Z(n21277) );
  NANDN U29843 ( .A(n21309), .B(n21310), .Z(n21308) );
  NANDN U29844 ( .A(n21311), .B(n21312), .Z(n21310) );
  NANDN U29845 ( .A(n21312), .B(n21311), .Z(n21307) );
  IV U29846 ( .A(n21313), .Z(n21311) );
  AND U29847 ( .A(n21314), .B(n21315), .Z(n21280) );
  NAND U29848 ( .A(n21316), .B(n21317), .Z(n21315) );
  NANDN U29849 ( .A(n21318), .B(n21319), .Z(n21317) );
  NANDN U29850 ( .A(n21319), .B(n21318), .Z(n21314) );
  XOR U29851 ( .A(n21290), .B(n21320), .Z(n21282) );
  XNOR U29852 ( .A(n21287), .B(n21289), .Z(n21320) );
  AND U29853 ( .A(n21321), .B(n21322), .Z(n21289) );
  NANDN U29854 ( .A(n21323), .B(n21324), .Z(n21322) );
  OR U29855 ( .A(n21325), .B(n21326), .Z(n21324) );
  IV U29856 ( .A(n21327), .Z(n21326) );
  NANDN U29857 ( .A(n21327), .B(n21325), .Z(n21321) );
  AND U29858 ( .A(n21328), .B(n21329), .Z(n21287) );
  NAND U29859 ( .A(n21330), .B(n21331), .Z(n21329) );
  NANDN U29860 ( .A(n21332), .B(n21333), .Z(n21331) );
  NANDN U29861 ( .A(n21333), .B(n21332), .Z(n21328) );
  IV U29862 ( .A(n21334), .Z(n21333) );
  NAND U29863 ( .A(n21335), .B(n21336), .Z(n21290) );
  NANDN U29864 ( .A(n21337), .B(n21338), .Z(n21336) );
  NANDN U29865 ( .A(n21339), .B(n21340), .Z(n21338) );
  NANDN U29866 ( .A(n21340), .B(n21339), .Z(n21335) );
  IV U29867 ( .A(n21341), .Z(n21339) );
  XOR U29868 ( .A(n21316), .B(n21342), .Z(N63492) );
  XNOR U29869 ( .A(n21319), .B(n21318), .Z(n21342) );
  XNOR U29870 ( .A(n21330), .B(n21343), .Z(n21318) );
  XNOR U29871 ( .A(n21334), .B(n21332), .Z(n21343) );
  XOR U29872 ( .A(n21340), .B(n21344), .Z(n21332) );
  XNOR U29873 ( .A(n21337), .B(n21341), .Z(n21344) );
  AND U29874 ( .A(n21345), .B(n21346), .Z(n21341) );
  NAND U29875 ( .A(n21347), .B(n21348), .Z(n21346) );
  NAND U29876 ( .A(n21349), .B(n21350), .Z(n21345) );
  AND U29877 ( .A(n21351), .B(n21352), .Z(n21337) );
  NAND U29878 ( .A(n21353), .B(n21354), .Z(n21352) );
  NAND U29879 ( .A(n21355), .B(n21356), .Z(n21351) );
  NANDN U29880 ( .A(n21357), .B(n21358), .Z(n21340) );
  ANDN U29881 ( .B(n21359), .A(n21360), .Z(n21334) );
  XNOR U29882 ( .A(n21325), .B(n21361), .Z(n21330) );
  XNOR U29883 ( .A(n21323), .B(n21327), .Z(n21361) );
  AND U29884 ( .A(n21362), .B(n21363), .Z(n21327) );
  NAND U29885 ( .A(n21364), .B(n21365), .Z(n21363) );
  NAND U29886 ( .A(n21366), .B(n21367), .Z(n21362) );
  AND U29887 ( .A(n21368), .B(n21369), .Z(n21323) );
  NAND U29888 ( .A(n21370), .B(n21371), .Z(n21369) );
  NAND U29889 ( .A(n21372), .B(n21373), .Z(n21368) );
  AND U29890 ( .A(n21374), .B(n21375), .Z(n21325) );
  NAND U29891 ( .A(n21376), .B(n21377), .Z(n21319) );
  XNOR U29892 ( .A(n21302), .B(n21378), .Z(n21316) );
  XNOR U29893 ( .A(n21306), .B(n21304), .Z(n21378) );
  XOR U29894 ( .A(n21312), .B(n21379), .Z(n21304) );
  XNOR U29895 ( .A(n21309), .B(n21313), .Z(n21379) );
  AND U29896 ( .A(n21380), .B(n21381), .Z(n21313) );
  NAND U29897 ( .A(n21382), .B(n21383), .Z(n21381) );
  NAND U29898 ( .A(n21384), .B(n21385), .Z(n21380) );
  AND U29899 ( .A(n21386), .B(n21387), .Z(n21309) );
  NAND U29900 ( .A(n21388), .B(n21389), .Z(n21387) );
  NAND U29901 ( .A(n21390), .B(n21391), .Z(n21386) );
  NANDN U29902 ( .A(n21392), .B(n21393), .Z(n21312) );
  ANDN U29903 ( .B(n21394), .A(n21395), .Z(n21306) );
  XNOR U29904 ( .A(n21297), .B(n21396), .Z(n21302) );
  XNOR U29905 ( .A(n21295), .B(n21299), .Z(n21396) );
  AND U29906 ( .A(n21397), .B(n21398), .Z(n21299) );
  NAND U29907 ( .A(n21399), .B(n21400), .Z(n21398) );
  NAND U29908 ( .A(n21401), .B(n21402), .Z(n21397) );
  AND U29909 ( .A(n21403), .B(n21404), .Z(n21295) );
  NAND U29910 ( .A(n21405), .B(n21406), .Z(n21404) );
  NAND U29911 ( .A(n21407), .B(n21408), .Z(n21403) );
  AND U29912 ( .A(n21409), .B(n21410), .Z(n21297) );
  XOR U29913 ( .A(n21377), .B(n21376), .Z(N63491) );
  XNOR U29914 ( .A(n21394), .B(n21395), .Z(n21376) );
  XNOR U29915 ( .A(n21409), .B(n21410), .Z(n21395) );
  XOR U29916 ( .A(n21406), .B(n21405), .Z(n21410) );
  XOR U29917 ( .A(y[5364]), .B(x[5364]), .Z(n21405) );
  XOR U29918 ( .A(n21408), .B(n21407), .Z(n21406) );
  XOR U29919 ( .A(y[5366]), .B(x[5366]), .Z(n21407) );
  XOR U29920 ( .A(y[5365]), .B(x[5365]), .Z(n21408) );
  XOR U29921 ( .A(n21400), .B(n21399), .Z(n21409) );
  XOR U29922 ( .A(n21402), .B(n21401), .Z(n21399) );
  XOR U29923 ( .A(y[5363]), .B(x[5363]), .Z(n21401) );
  XOR U29924 ( .A(y[5362]), .B(x[5362]), .Z(n21402) );
  XOR U29925 ( .A(y[5361]), .B(x[5361]), .Z(n21400) );
  XNOR U29926 ( .A(n21393), .B(n21392), .Z(n21394) );
  XNOR U29927 ( .A(n21389), .B(n21388), .Z(n21392) );
  XOR U29928 ( .A(n21391), .B(n21390), .Z(n21388) );
  XOR U29929 ( .A(y[5360]), .B(x[5360]), .Z(n21390) );
  XOR U29930 ( .A(y[5359]), .B(x[5359]), .Z(n21391) );
  XOR U29931 ( .A(y[5358]), .B(x[5358]), .Z(n21389) );
  XOR U29932 ( .A(n21383), .B(n21382), .Z(n21393) );
  XOR U29933 ( .A(n21385), .B(n21384), .Z(n21382) );
  XOR U29934 ( .A(y[5357]), .B(x[5357]), .Z(n21384) );
  XOR U29935 ( .A(y[5356]), .B(x[5356]), .Z(n21385) );
  XOR U29936 ( .A(y[5355]), .B(x[5355]), .Z(n21383) );
  XNOR U29937 ( .A(n21359), .B(n21360), .Z(n21377) );
  XNOR U29938 ( .A(n21374), .B(n21375), .Z(n21360) );
  XOR U29939 ( .A(n21371), .B(n21370), .Z(n21375) );
  XOR U29940 ( .A(y[5352]), .B(x[5352]), .Z(n21370) );
  XOR U29941 ( .A(n21373), .B(n21372), .Z(n21371) );
  XOR U29942 ( .A(y[5354]), .B(x[5354]), .Z(n21372) );
  XOR U29943 ( .A(y[5353]), .B(x[5353]), .Z(n21373) );
  XOR U29944 ( .A(n21365), .B(n21364), .Z(n21374) );
  XOR U29945 ( .A(n21367), .B(n21366), .Z(n21364) );
  XOR U29946 ( .A(y[5351]), .B(x[5351]), .Z(n21366) );
  XOR U29947 ( .A(y[5350]), .B(x[5350]), .Z(n21367) );
  XOR U29948 ( .A(y[5349]), .B(x[5349]), .Z(n21365) );
  XNOR U29949 ( .A(n21358), .B(n21357), .Z(n21359) );
  XNOR U29950 ( .A(n21354), .B(n21353), .Z(n21357) );
  XOR U29951 ( .A(n21356), .B(n21355), .Z(n21353) );
  XOR U29952 ( .A(y[5348]), .B(x[5348]), .Z(n21355) );
  XOR U29953 ( .A(y[5347]), .B(x[5347]), .Z(n21356) );
  XOR U29954 ( .A(y[5346]), .B(x[5346]), .Z(n21354) );
  XOR U29955 ( .A(n21348), .B(n21347), .Z(n21358) );
  XOR U29956 ( .A(n21350), .B(n21349), .Z(n21347) );
  XOR U29957 ( .A(y[5345]), .B(x[5345]), .Z(n21349) );
  XOR U29958 ( .A(y[5344]), .B(x[5344]), .Z(n21350) );
  XOR U29959 ( .A(y[5343]), .B(x[5343]), .Z(n21348) );
  NAND U29960 ( .A(n21411), .B(n21412), .Z(N63482) );
  NAND U29961 ( .A(n21413), .B(n21414), .Z(n21412) );
  NANDN U29962 ( .A(n21415), .B(n21416), .Z(n21414) );
  NANDN U29963 ( .A(n21416), .B(n21415), .Z(n21411) );
  XOR U29964 ( .A(n21415), .B(n21417), .Z(N63481) );
  XNOR U29965 ( .A(n21413), .B(n21416), .Z(n21417) );
  NAND U29966 ( .A(n21418), .B(n21419), .Z(n21416) );
  NAND U29967 ( .A(n21420), .B(n21421), .Z(n21419) );
  NANDN U29968 ( .A(n21422), .B(n21423), .Z(n21421) );
  NANDN U29969 ( .A(n21423), .B(n21422), .Z(n21418) );
  AND U29970 ( .A(n21424), .B(n21425), .Z(n21413) );
  NAND U29971 ( .A(n21426), .B(n21427), .Z(n21425) );
  NANDN U29972 ( .A(n21428), .B(n21429), .Z(n21427) );
  NANDN U29973 ( .A(n21429), .B(n21428), .Z(n21424) );
  IV U29974 ( .A(n21430), .Z(n21429) );
  AND U29975 ( .A(n21431), .B(n21432), .Z(n21415) );
  NAND U29976 ( .A(n21433), .B(n21434), .Z(n21432) );
  NANDN U29977 ( .A(n21435), .B(n21436), .Z(n21434) );
  NANDN U29978 ( .A(n21436), .B(n21435), .Z(n21431) );
  XOR U29979 ( .A(n21428), .B(n21437), .Z(N63480) );
  XNOR U29980 ( .A(n21426), .B(n21430), .Z(n21437) );
  XOR U29981 ( .A(n21423), .B(n21438), .Z(n21430) );
  XNOR U29982 ( .A(n21420), .B(n21422), .Z(n21438) );
  AND U29983 ( .A(n21439), .B(n21440), .Z(n21422) );
  NANDN U29984 ( .A(n21441), .B(n21442), .Z(n21440) );
  OR U29985 ( .A(n21443), .B(n21444), .Z(n21442) );
  IV U29986 ( .A(n21445), .Z(n21444) );
  NANDN U29987 ( .A(n21445), .B(n21443), .Z(n21439) );
  AND U29988 ( .A(n21446), .B(n21447), .Z(n21420) );
  NAND U29989 ( .A(n21448), .B(n21449), .Z(n21447) );
  NANDN U29990 ( .A(n21450), .B(n21451), .Z(n21449) );
  NANDN U29991 ( .A(n21451), .B(n21450), .Z(n21446) );
  IV U29992 ( .A(n21452), .Z(n21451) );
  NAND U29993 ( .A(n21453), .B(n21454), .Z(n21423) );
  NANDN U29994 ( .A(n21455), .B(n21456), .Z(n21454) );
  NANDN U29995 ( .A(n21457), .B(n21458), .Z(n21456) );
  NANDN U29996 ( .A(n21458), .B(n21457), .Z(n21453) );
  IV U29997 ( .A(n21459), .Z(n21457) );
  AND U29998 ( .A(n21460), .B(n21461), .Z(n21426) );
  NAND U29999 ( .A(n21462), .B(n21463), .Z(n21461) );
  NANDN U30000 ( .A(n21464), .B(n21465), .Z(n21463) );
  NANDN U30001 ( .A(n21465), .B(n21464), .Z(n21460) );
  XOR U30002 ( .A(n21436), .B(n21466), .Z(n21428) );
  XNOR U30003 ( .A(n21433), .B(n21435), .Z(n21466) );
  AND U30004 ( .A(n21467), .B(n21468), .Z(n21435) );
  NANDN U30005 ( .A(n21469), .B(n21470), .Z(n21468) );
  OR U30006 ( .A(n21471), .B(n21472), .Z(n21470) );
  IV U30007 ( .A(n21473), .Z(n21472) );
  NANDN U30008 ( .A(n21473), .B(n21471), .Z(n21467) );
  AND U30009 ( .A(n21474), .B(n21475), .Z(n21433) );
  NAND U30010 ( .A(n21476), .B(n21477), .Z(n21475) );
  NANDN U30011 ( .A(n21478), .B(n21479), .Z(n21477) );
  NANDN U30012 ( .A(n21479), .B(n21478), .Z(n21474) );
  IV U30013 ( .A(n21480), .Z(n21479) );
  NAND U30014 ( .A(n21481), .B(n21482), .Z(n21436) );
  NANDN U30015 ( .A(n21483), .B(n21484), .Z(n21482) );
  NANDN U30016 ( .A(n21485), .B(n21486), .Z(n21484) );
  NANDN U30017 ( .A(n21486), .B(n21485), .Z(n21481) );
  IV U30018 ( .A(n21487), .Z(n21485) );
  XOR U30019 ( .A(n21462), .B(n21488), .Z(N63479) );
  XNOR U30020 ( .A(n21465), .B(n21464), .Z(n21488) );
  XNOR U30021 ( .A(n21476), .B(n21489), .Z(n21464) );
  XNOR U30022 ( .A(n21480), .B(n21478), .Z(n21489) );
  XOR U30023 ( .A(n21486), .B(n21490), .Z(n21478) );
  XNOR U30024 ( .A(n21483), .B(n21487), .Z(n21490) );
  AND U30025 ( .A(n21491), .B(n21492), .Z(n21487) );
  NAND U30026 ( .A(n21493), .B(n21494), .Z(n21492) );
  NAND U30027 ( .A(n21495), .B(n21496), .Z(n21491) );
  AND U30028 ( .A(n21497), .B(n21498), .Z(n21483) );
  NAND U30029 ( .A(n21499), .B(n21500), .Z(n21498) );
  NAND U30030 ( .A(n21501), .B(n21502), .Z(n21497) );
  NANDN U30031 ( .A(n21503), .B(n21504), .Z(n21486) );
  ANDN U30032 ( .B(n21505), .A(n21506), .Z(n21480) );
  XNOR U30033 ( .A(n21471), .B(n21507), .Z(n21476) );
  XNOR U30034 ( .A(n21469), .B(n21473), .Z(n21507) );
  AND U30035 ( .A(n21508), .B(n21509), .Z(n21473) );
  NAND U30036 ( .A(n21510), .B(n21511), .Z(n21509) );
  NAND U30037 ( .A(n21512), .B(n21513), .Z(n21508) );
  AND U30038 ( .A(n21514), .B(n21515), .Z(n21469) );
  NAND U30039 ( .A(n21516), .B(n21517), .Z(n21515) );
  NAND U30040 ( .A(n21518), .B(n21519), .Z(n21514) );
  AND U30041 ( .A(n21520), .B(n21521), .Z(n21471) );
  NAND U30042 ( .A(n21522), .B(n21523), .Z(n21465) );
  XNOR U30043 ( .A(n21448), .B(n21524), .Z(n21462) );
  XNOR U30044 ( .A(n21452), .B(n21450), .Z(n21524) );
  XOR U30045 ( .A(n21458), .B(n21525), .Z(n21450) );
  XNOR U30046 ( .A(n21455), .B(n21459), .Z(n21525) );
  AND U30047 ( .A(n21526), .B(n21527), .Z(n21459) );
  NAND U30048 ( .A(n21528), .B(n21529), .Z(n21527) );
  NAND U30049 ( .A(n21530), .B(n21531), .Z(n21526) );
  AND U30050 ( .A(n21532), .B(n21533), .Z(n21455) );
  NAND U30051 ( .A(n21534), .B(n21535), .Z(n21533) );
  NAND U30052 ( .A(n21536), .B(n21537), .Z(n21532) );
  NANDN U30053 ( .A(n21538), .B(n21539), .Z(n21458) );
  ANDN U30054 ( .B(n21540), .A(n21541), .Z(n21452) );
  XNOR U30055 ( .A(n21443), .B(n21542), .Z(n21448) );
  XNOR U30056 ( .A(n21441), .B(n21445), .Z(n21542) );
  AND U30057 ( .A(n21543), .B(n21544), .Z(n21445) );
  NAND U30058 ( .A(n21545), .B(n21546), .Z(n21544) );
  NAND U30059 ( .A(n21547), .B(n21548), .Z(n21543) );
  AND U30060 ( .A(n21549), .B(n21550), .Z(n21441) );
  NAND U30061 ( .A(n21551), .B(n21552), .Z(n21550) );
  NAND U30062 ( .A(n21553), .B(n21554), .Z(n21549) );
  AND U30063 ( .A(n21555), .B(n21556), .Z(n21443) );
  XOR U30064 ( .A(n21523), .B(n21522), .Z(N63478) );
  XNOR U30065 ( .A(n21540), .B(n21541), .Z(n21522) );
  XNOR U30066 ( .A(n21555), .B(n21556), .Z(n21541) );
  XOR U30067 ( .A(n21552), .B(n21551), .Z(n21556) );
  XOR U30068 ( .A(y[5340]), .B(x[5340]), .Z(n21551) );
  XOR U30069 ( .A(n21554), .B(n21553), .Z(n21552) );
  XOR U30070 ( .A(y[5342]), .B(x[5342]), .Z(n21553) );
  XOR U30071 ( .A(y[5341]), .B(x[5341]), .Z(n21554) );
  XOR U30072 ( .A(n21546), .B(n21545), .Z(n21555) );
  XOR U30073 ( .A(n21548), .B(n21547), .Z(n21545) );
  XOR U30074 ( .A(y[5339]), .B(x[5339]), .Z(n21547) );
  XOR U30075 ( .A(y[5338]), .B(x[5338]), .Z(n21548) );
  XOR U30076 ( .A(y[5337]), .B(x[5337]), .Z(n21546) );
  XNOR U30077 ( .A(n21539), .B(n21538), .Z(n21540) );
  XNOR U30078 ( .A(n21535), .B(n21534), .Z(n21538) );
  XOR U30079 ( .A(n21537), .B(n21536), .Z(n21534) );
  XOR U30080 ( .A(y[5336]), .B(x[5336]), .Z(n21536) );
  XOR U30081 ( .A(y[5335]), .B(x[5335]), .Z(n21537) );
  XOR U30082 ( .A(y[5334]), .B(x[5334]), .Z(n21535) );
  XOR U30083 ( .A(n21529), .B(n21528), .Z(n21539) );
  XOR U30084 ( .A(n21531), .B(n21530), .Z(n21528) );
  XOR U30085 ( .A(y[5333]), .B(x[5333]), .Z(n21530) );
  XOR U30086 ( .A(y[5332]), .B(x[5332]), .Z(n21531) );
  XOR U30087 ( .A(y[5331]), .B(x[5331]), .Z(n21529) );
  XNOR U30088 ( .A(n21505), .B(n21506), .Z(n21523) );
  XNOR U30089 ( .A(n21520), .B(n21521), .Z(n21506) );
  XOR U30090 ( .A(n21517), .B(n21516), .Z(n21521) );
  XOR U30091 ( .A(y[5328]), .B(x[5328]), .Z(n21516) );
  XOR U30092 ( .A(n21519), .B(n21518), .Z(n21517) );
  XOR U30093 ( .A(y[5330]), .B(x[5330]), .Z(n21518) );
  XOR U30094 ( .A(y[5329]), .B(x[5329]), .Z(n21519) );
  XOR U30095 ( .A(n21511), .B(n21510), .Z(n21520) );
  XOR U30096 ( .A(n21513), .B(n21512), .Z(n21510) );
  XOR U30097 ( .A(y[5327]), .B(x[5327]), .Z(n21512) );
  XOR U30098 ( .A(y[5326]), .B(x[5326]), .Z(n21513) );
  XOR U30099 ( .A(y[5325]), .B(x[5325]), .Z(n21511) );
  XNOR U30100 ( .A(n21504), .B(n21503), .Z(n21505) );
  XNOR U30101 ( .A(n21500), .B(n21499), .Z(n21503) );
  XOR U30102 ( .A(n21502), .B(n21501), .Z(n21499) );
  XOR U30103 ( .A(y[5324]), .B(x[5324]), .Z(n21501) );
  XOR U30104 ( .A(y[5323]), .B(x[5323]), .Z(n21502) );
  XOR U30105 ( .A(y[5322]), .B(x[5322]), .Z(n21500) );
  XOR U30106 ( .A(n21494), .B(n21493), .Z(n21504) );
  XOR U30107 ( .A(n21496), .B(n21495), .Z(n21493) );
  XOR U30108 ( .A(y[5321]), .B(x[5321]), .Z(n21495) );
  XOR U30109 ( .A(y[5320]), .B(x[5320]), .Z(n21496) );
  XOR U30110 ( .A(y[5319]), .B(x[5319]), .Z(n21494) );
  NAND U30111 ( .A(n21557), .B(n21558), .Z(N63469) );
  NAND U30112 ( .A(n21559), .B(n21560), .Z(n21558) );
  NANDN U30113 ( .A(n21561), .B(n21562), .Z(n21560) );
  NANDN U30114 ( .A(n21562), .B(n21561), .Z(n21557) );
  XOR U30115 ( .A(n21561), .B(n21563), .Z(N63468) );
  XNOR U30116 ( .A(n21559), .B(n21562), .Z(n21563) );
  NAND U30117 ( .A(n21564), .B(n21565), .Z(n21562) );
  NAND U30118 ( .A(n21566), .B(n21567), .Z(n21565) );
  NANDN U30119 ( .A(n21568), .B(n21569), .Z(n21567) );
  NANDN U30120 ( .A(n21569), .B(n21568), .Z(n21564) );
  AND U30121 ( .A(n21570), .B(n21571), .Z(n21559) );
  NAND U30122 ( .A(n21572), .B(n21573), .Z(n21571) );
  NANDN U30123 ( .A(n21574), .B(n21575), .Z(n21573) );
  NANDN U30124 ( .A(n21575), .B(n21574), .Z(n21570) );
  IV U30125 ( .A(n21576), .Z(n21575) );
  AND U30126 ( .A(n21577), .B(n21578), .Z(n21561) );
  NAND U30127 ( .A(n21579), .B(n21580), .Z(n21578) );
  NANDN U30128 ( .A(n21581), .B(n21582), .Z(n21580) );
  NANDN U30129 ( .A(n21582), .B(n21581), .Z(n21577) );
  XOR U30130 ( .A(n21574), .B(n21583), .Z(N63467) );
  XNOR U30131 ( .A(n21572), .B(n21576), .Z(n21583) );
  XOR U30132 ( .A(n21569), .B(n21584), .Z(n21576) );
  XNOR U30133 ( .A(n21566), .B(n21568), .Z(n21584) );
  AND U30134 ( .A(n21585), .B(n21586), .Z(n21568) );
  NANDN U30135 ( .A(n21587), .B(n21588), .Z(n21586) );
  OR U30136 ( .A(n21589), .B(n21590), .Z(n21588) );
  IV U30137 ( .A(n21591), .Z(n21590) );
  NANDN U30138 ( .A(n21591), .B(n21589), .Z(n21585) );
  AND U30139 ( .A(n21592), .B(n21593), .Z(n21566) );
  NAND U30140 ( .A(n21594), .B(n21595), .Z(n21593) );
  NANDN U30141 ( .A(n21596), .B(n21597), .Z(n21595) );
  NANDN U30142 ( .A(n21597), .B(n21596), .Z(n21592) );
  IV U30143 ( .A(n21598), .Z(n21597) );
  NAND U30144 ( .A(n21599), .B(n21600), .Z(n21569) );
  NANDN U30145 ( .A(n21601), .B(n21602), .Z(n21600) );
  NANDN U30146 ( .A(n21603), .B(n21604), .Z(n21602) );
  NANDN U30147 ( .A(n21604), .B(n21603), .Z(n21599) );
  IV U30148 ( .A(n21605), .Z(n21603) );
  AND U30149 ( .A(n21606), .B(n21607), .Z(n21572) );
  NAND U30150 ( .A(n21608), .B(n21609), .Z(n21607) );
  NANDN U30151 ( .A(n21610), .B(n21611), .Z(n21609) );
  NANDN U30152 ( .A(n21611), .B(n21610), .Z(n21606) );
  XOR U30153 ( .A(n21582), .B(n21612), .Z(n21574) );
  XNOR U30154 ( .A(n21579), .B(n21581), .Z(n21612) );
  AND U30155 ( .A(n21613), .B(n21614), .Z(n21581) );
  NANDN U30156 ( .A(n21615), .B(n21616), .Z(n21614) );
  OR U30157 ( .A(n21617), .B(n21618), .Z(n21616) );
  IV U30158 ( .A(n21619), .Z(n21618) );
  NANDN U30159 ( .A(n21619), .B(n21617), .Z(n21613) );
  AND U30160 ( .A(n21620), .B(n21621), .Z(n21579) );
  NAND U30161 ( .A(n21622), .B(n21623), .Z(n21621) );
  NANDN U30162 ( .A(n21624), .B(n21625), .Z(n21623) );
  NANDN U30163 ( .A(n21625), .B(n21624), .Z(n21620) );
  IV U30164 ( .A(n21626), .Z(n21625) );
  NAND U30165 ( .A(n21627), .B(n21628), .Z(n21582) );
  NANDN U30166 ( .A(n21629), .B(n21630), .Z(n21628) );
  NANDN U30167 ( .A(n21631), .B(n21632), .Z(n21630) );
  NANDN U30168 ( .A(n21632), .B(n21631), .Z(n21627) );
  IV U30169 ( .A(n21633), .Z(n21631) );
  XOR U30170 ( .A(n21608), .B(n21634), .Z(N63466) );
  XNOR U30171 ( .A(n21611), .B(n21610), .Z(n21634) );
  XNOR U30172 ( .A(n21622), .B(n21635), .Z(n21610) );
  XNOR U30173 ( .A(n21626), .B(n21624), .Z(n21635) );
  XOR U30174 ( .A(n21632), .B(n21636), .Z(n21624) );
  XNOR U30175 ( .A(n21629), .B(n21633), .Z(n21636) );
  AND U30176 ( .A(n21637), .B(n21638), .Z(n21633) );
  NAND U30177 ( .A(n21639), .B(n21640), .Z(n21638) );
  NAND U30178 ( .A(n21641), .B(n21642), .Z(n21637) );
  AND U30179 ( .A(n21643), .B(n21644), .Z(n21629) );
  NAND U30180 ( .A(n21645), .B(n21646), .Z(n21644) );
  NAND U30181 ( .A(n21647), .B(n21648), .Z(n21643) );
  NANDN U30182 ( .A(n21649), .B(n21650), .Z(n21632) );
  ANDN U30183 ( .B(n21651), .A(n21652), .Z(n21626) );
  XNOR U30184 ( .A(n21617), .B(n21653), .Z(n21622) );
  XNOR U30185 ( .A(n21615), .B(n21619), .Z(n21653) );
  AND U30186 ( .A(n21654), .B(n21655), .Z(n21619) );
  NAND U30187 ( .A(n21656), .B(n21657), .Z(n21655) );
  NAND U30188 ( .A(n21658), .B(n21659), .Z(n21654) );
  AND U30189 ( .A(n21660), .B(n21661), .Z(n21615) );
  NAND U30190 ( .A(n21662), .B(n21663), .Z(n21661) );
  NAND U30191 ( .A(n21664), .B(n21665), .Z(n21660) );
  AND U30192 ( .A(n21666), .B(n21667), .Z(n21617) );
  NAND U30193 ( .A(n21668), .B(n21669), .Z(n21611) );
  XNOR U30194 ( .A(n21594), .B(n21670), .Z(n21608) );
  XNOR U30195 ( .A(n21598), .B(n21596), .Z(n21670) );
  XOR U30196 ( .A(n21604), .B(n21671), .Z(n21596) );
  XNOR U30197 ( .A(n21601), .B(n21605), .Z(n21671) );
  AND U30198 ( .A(n21672), .B(n21673), .Z(n21605) );
  NAND U30199 ( .A(n21674), .B(n21675), .Z(n21673) );
  NAND U30200 ( .A(n21676), .B(n21677), .Z(n21672) );
  AND U30201 ( .A(n21678), .B(n21679), .Z(n21601) );
  NAND U30202 ( .A(n21680), .B(n21681), .Z(n21679) );
  NAND U30203 ( .A(n21682), .B(n21683), .Z(n21678) );
  NANDN U30204 ( .A(n21684), .B(n21685), .Z(n21604) );
  ANDN U30205 ( .B(n21686), .A(n21687), .Z(n21598) );
  XNOR U30206 ( .A(n21589), .B(n21688), .Z(n21594) );
  XNOR U30207 ( .A(n21587), .B(n21591), .Z(n21688) );
  AND U30208 ( .A(n21689), .B(n21690), .Z(n21591) );
  NAND U30209 ( .A(n21691), .B(n21692), .Z(n21690) );
  NAND U30210 ( .A(n21693), .B(n21694), .Z(n21689) );
  AND U30211 ( .A(n21695), .B(n21696), .Z(n21587) );
  NAND U30212 ( .A(n21697), .B(n21698), .Z(n21696) );
  NAND U30213 ( .A(n21699), .B(n21700), .Z(n21695) );
  AND U30214 ( .A(n21701), .B(n21702), .Z(n21589) );
  XOR U30215 ( .A(n21669), .B(n21668), .Z(N63465) );
  XNOR U30216 ( .A(n21686), .B(n21687), .Z(n21668) );
  XNOR U30217 ( .A(n21701), .B(n21702), .Z(n21687) );
  XOR U30218 ( .A(n21698), .B(n21697), .Z(n21702) );
  XOR U30219 ( .A(y[5316]), .B(x[5316]), .Z(n21697) );
  XOR U30220 ( .A(n21700), .B(n21699), .Z(n21698) );
  XOR U30221 ( .A(y[5318]), .B(x[5318]), .Z(n21699) );
  XOR U30222 ( .A(y[5317]), .B(x[5317]), .Z(n21700) );
  XOR U30223 ( .A(n21692), .B(n21691), .Z(n21701) );
  XOR U30224 ( .A(n21694), .B(n21693), .Z(n21691) );
  XOR U30225 ( .A(y[5315]), .B(x[5315]), .Z(n21693) );
  XOR U30226 ( .A(y[5314]), .B(x[5314]), .Z(n21694) );
  XOR U30227 ( .A(y[5313]), .B(x[5313]), .Z(n21692) );
  XNOR U30228 ( .A(n21685), .B(n21684), .Z(n21686) );
  XNOR U30229 ( .A(n21681), .B(n21680), .Z(n21684) );
  XOR U30230 ( .A(n21683), .B(n21682), .Z(n21680) );
  XOR U30231 ( .A(y[5312]), .B(x[5312]), .Z(n21682) );
  XOR U30232 ( .A(y[5311]), .B(x[5311]), .Z(n21683) );
  XOR U30233 ( .A(y[5310]), .B(x[5310]), .Z(n21681) );
  XOR U30234 ( .A(n21675), .B(n21674), .Z(n21685) );
  XOR U30235 ( .A(n21677), .B(n21676), .Z(n21674) );
  XOR U30236 ( .A(y[5309]), .B(x[5309]), .Z(n21676) );
  XOR U30237 ( .A(y[5308]), .B(x[5308]), .Z(n21677) );
  XOR U30238 ( .A(y[5307]), .B(x[5307]), .Z(n21675) );
  XNOR U30239 ( .A(n21651), .B(n21652), .Z(n21669) );
  XNOR U30240 ( .A(n21666), .B(n21667), .Z(n21652) );
  XOR U30241 ( .A(n21663), .B(n21662), .Z(n21667) );
  XOR U30242 ( .A(y[5304]), .B(x[5304]), .Z(n21662) );
  XOR U30243 ( .A(n21665), .B(n21664), .Z(n21663) );
  XOR U30244 ( .A(y[5306]), .B(x[5306]), .Z(n21664) );
  XOR U30245 ( .A(y[5305]), .B(x[5305]), .Z(n21665) );
  XOR U30246 ( .A(n21657), .B(n21656), .Z(n21666) );
  XOR U30247 ( .A(n21659), .B(n21658), .Z(n21656) );
  XOR U30248 ( .A(y[5303]), .B(x[5303]), .Z(n21658) );
  XOR U30249 ( .A(y[5302]), .B(x[5302]), .Z(n21659) );
  XOR U30250 ( .A(y[5301]), .B(x[5301]), .Z(n21657) );
  XNOR U30251 ( .A(n21650), .B(n21649), .Z(n21651) );
  XNOR U30252 ( .A(n21646), .B(n21645), .Z(n21649) );
  XOR U30253 ( .A(n21648), .B(n21647), .Z(n21645) );
  XOR U30254 ( .A(y[5300]), .B(x[5300]), .Z(n21647) );
  XOR U30255 ( .A(y[5299]), .B(x[5299]), .Z(n21648) );
  XOR U30256 ( .A(y[5298]), .B(x[5298]), .Z(n21646) );
  XOR U30257 ( .A(n21640), .B(n21639), .Z(n21650) );
  XOR U30258 ( .A(n21642), .B(n21641), .Z(n21639) );
  XOR U30259 ( .A(y[5297]), .B(x[5297]), .Z(n21641) );
  XOR U30260 ( .A(y[5296]), .B(x[5296]), .Z(n21642) );
  XOR U30261 ( .A(y[5295]), .B(x[5295]), .Z(n21640) );
  NAND U30262 ( .A(n21703), .B(n21704), .Z(N63456) );
  NAND U30263 ( .A(n21705), .B(n21706), .Z(n21704) );
  NANDN U30264 ( .A(n21707), .B(n21708), .Z(n21706) );
  NANDN U30265 ( .A(n21708), .B(n21707), .Z(n21703) );
  XOR U30266 ( .A(n21707), .B(n21709), .Z(N63455) );
  XNOR U30267 ( .A(n21705), .B(n21708), .Z(n21709) );
  NAND U30268 ( .A(n21710), .B(n21711), .Z(n21708) );
  NAND U30269 ( .A(n21712), .B(n21713), .Z(n21711) );
  NANDN U30270 ( .A(n21714), .B(n21715), .Z(n21713) );
  NANDN U30271 ( .A(n21715), .B(n21714), .Z(n21710) );
  AND U30272 ( .A(n21716), .B(n21717), .Z(n21705) );
  NAND U30273 ( .A(n21718), .B(n21719), .Z(n21717) );
  NANDN U30274 ( .A(n21720), .B(n21721), .Z(n21719) );
  NANDN U30275 ( .A(n21721), .B(n21720), .Z(n21716) );
  IV U30276 ( .A(n21722), .Z(n21721) );
  AND U30277 ( .A(n21723), .B(n21724), .Z(n21707) );
  NAND U30278 ( .A(n21725), .B(n21726), .Z(n21724) );
  NANDN U30279 ( .A(n21727), .B(n21728), .Z(n21726) );
  NANDN U30280 ( .A(n21728), .B(n21727), .Z(n21723) );
  XOR U30281 ( .A(n21720), .B(n21729), .Z(N63454) );
  XNOR U30282 ( .A(n21718), .B(n21722), .Z(n21729) );
  XOR U30283 ( .A(n21715), .B(n21730), .Z(n21722) );
  XNOR U30284 ( .A(n21712), .B(n21714), .Z(n21730) );
  AND U30285 ( .A(n21731), .B(n21732), .Z(n21714) );
  NANDN U30286 ( .A(n21733), .B(n21734), .Z(n21732) );
  OR U30287 ( .A(n21735), .B(n21736), .Z(n21734) );
  IV U30288 ( .A(n21737), .Z(n21736) );
  NANDN U30289 ( .A(n21737), .B(n21735), .Z(n21731) );
  AND U30290 ( .A(n21738), .B(n21739), .Z(n21712) );
  NAND U30291 ( .A(n21740), .B(n21741), .Z(n21739) );
  NANDN U30292 ( .A(n21742), .B(n21743), .Z(n21741) );
  NANDN U30293 ( .A(n21743), .B(n21742), .Z(n21738) );
  IV U30294 ( .A(n21744), .Z(n21743) );
  NAND U30295 ( .A(n21745), .B(n21746), .Z(n21715) );
  NANDN U30296 ( .A(n21747), .B(n21748), .Z(n21746) );
  NANDN U30297 ( .A(n21749), .B(n21750), .Z(n21748) );
  NANDN U30298 ( .A(n21750), .B(n21749), .Z(n21745) );
  IV U30299 ( .A(n21751), .Z(n21749) );
  AND U30300 ( .A(n21752), .B(n21753), .Z(n21718) );
  NAND U30301 ( .A(n21754), .B(n21755), .Z(n21753) );
  NANDN U30302 ( .A(n21756), .B(n21757), .Z(n21755) );
  NANDN U30303 ( .A(n21757), .B(n21756), .Z(n21752) );
  XOR U30304 ( .A(n21728), .B(n21758), .Z(n21720) );
  XNOR U30305 ( .A(n21725), .B(n21727), .Z(n21758) );
  AND U30306 ( .A(n21759), .B(n21760), .Z(n21727) );
  NANDN U30307 ( .A(n21761), .B(n21762), .Z(n21760) );
  OR U30308 ( .A(n21763), .B(n21764), .Z(n21762) );
  IV U30309 ( .A(n21765), .Z(n21764) );
  NANDN U30310 ( .A(n21765), .B(n21763), .Z(n21759) );
  AND U30311 ( .A(n21766), .B(n21767), .Z(n21725) );
  NAND U30312 ( .A(n21768), .B(n21769), .Z(n21767) );
  NANDN U30313 ( .A(n21770), .B(n21771), .Z(n21769) );
  NANDN U30314 ( .A(n21771), .B(n21770), .Z(n21766) );
  IV U30315 ( .A(n21772), .Z(n21771) );
  NAND U30316 ( .A(n21773), .B(n21774), .Z(n21728) );
  NANDN U30317 ( .A(n21775), .B(n21776), .Z(n21774) );
  NANDN U30318 ( .A(n21777), .B(n21778), .Z(n21776) );
  NANDN U30319 ( .A(n21778), .B(n21777), .Z(n21773) );
  IV U30320 ( .A(n21779), .Z(n21777) );
  XOR U30321 ( .A(n21754), .B(n21780), .Z(N63453) );
  XNOR U30322 ( .A(n21757), .B(n21756), .Z(n21780) );
  XNOR U30323 ( .A(n21768), .B(n21781), .Z(n21756) );
  XNOR U30324 ( .A(n21772), .B(n21770), .Z(n21781) );
  XOR U30325 ( .A(n21778), .B(n21782), .Z(n21770) );
  XNOR U30326 ( .A(n21775), .B(n21779), .Z(n21782) );
  AND U30327 ( .A(n21783), .B(n21784), .Z(n21779) );
  NAND U30328 ( .A(n21785), .B(n21786), .Z(n21784) );
  NAND U30329 ( .A(n21787), .B(n21788), .Z(n21783) );
  AND U30330 ( .A(n21789), .B(n21790), .Z(n21775) );
  NAND U30331 ( .A(n21791), .B(n21792), .Z(n21790) );
  NAND U30332 ( .A(n21793), .B(n21794), .Z(n21789) );
  NANDN U30333 ( .A(n21795), .B(n21796), .Z(n21778) );
  ANDN U30334 ( .B(n21797), .A(n21798), .Z(n21772) );
  XNOR U30335 ( .A(n21763), .B(n21799), .Z(n21768) );
  XNOR U30336 ( .A(n21761), .B(n21765), .Z(n21799) );
  AND U30337 ( .A(n21800), .B(n21801), .Z(n21765) );
  NAND U30338 ( .A(n21802), .B(n21803), .Z(n21801) );
  NAND U30339 ( .A(n21804), .B(n21805), .Z(n21800) );
  AND U30340 ( .A(n21806), .B(n21807), .Z(n21761) );
  NAND U30341 ( .A(n21808), .B(n21809), .Z(n21807) );
  NAND U30342 ( .A(n21810), .B(n21811), .Z(n21806) );
  AND U30343 ( .A(n21812), .B(n21813), .Z(n21763) );
  NAND U30344 ( .A(n21814), .B(n21815), .Z(n21757) );
  XNOR U30345 ( .A(n21740), .B(n21816), .Z(n21754) );
  XNOR U30346 ( .A(n21744), .B(n21742), .Z(n21816) );
  XOR U30347 ( .A(n21750), .B(n21817), .Z(n21742) );
  XNOR U30348 ( .A(n21747), .B(n21751), .Z(n21817) );
  AND U30349 ( .A(n21818), .B(n21819), .Z(n21751) );
  NAND U30350 ( .A(n21820), .B(n21821), .Z(n21819) );
  NAND U30351 ( .A(n21822), .B(n21823), .Z(n21818) );
  AND U30352 ( .A(n21824), .B(n21825), .Z(n21747) );
  NAND U30353 ( .A(n21826), .B(n21827), .Z(n21825) );
  NAND U30354 ( .A(n21828), .B(n21829), .Z(n21824) );
  NANDN U30355 ( .A(n21830), .B(n21831), .Z(n21750) );
  ANDN U30356 ( .B(n21832), .A(n21833), .Z(n21744) );
  XNOR U30357 ( .A(n21735), .B(n21834), .Z(n21740) );
  XNOR U30358 ( .A(n21733), .B(n21737), .Z(n21834) );
  AND U30359 ( .A(n21835), .B(n21836), .Z(n21737) );
  NAND U30360 ( .A(n21837), .B(n21838), .Z(n21836) );
  NAND U30361 ( .A(n21839), .B(n21840), .Z(n21835) );
  AND U30362 ( .A(n21841), .B(n21842), .Z(n21733) );
  NAND U30363 ( .A(n21843), .B(n21844), .Z(n21842) );
  NAND U30364 ( .A(n21845), .B(n21846), .Z(n21841) );
  AND U30365 ( .A(n21847), .B(n21848), .Z(n21735) );
  XOR U30366 ( .A(n21815), .B(n21814), .Z(N63452) );
  XNOR U30367 ( .A(n21832), .B(n21833), .Z(n21814) );
  XNOR U30368 ( .A(n21847), .B(n21848), .Z(n21833) );
  XOR U30369 ( .A(n21844), .B(n21843), .Z(n21848) );
  XOR U30370 ( .A(y[5292]), .B(x[5292]), .Z(n21843) );
  XOR U30371 ( .A(n21846), .B(n21845), .Z(n21844) );
  XOR U30372 ( .A(y[5294]), .B(x[5294]), .Z(n21845) );
  XOR U30373 ( .A(y[5293]), .B(x[5293]), .Z(n21846) );
  XOR U30374 ( .A(n21838), .B(n21837), .Z(n21847) );
  XOR U30375 ( .A(n21840), .B(n21839), .Z(n21837) );
  XOR U30376 ( .A(y[5291]), .B(x[5291]), .Z(n21839) );
  XOR U30377 ( .A(y[5290]), .B(x[5290]), .Z(n21840) );
  XOR U30378 ( .A(y[5289]), .B(x[5289]), .Z(n21838) );
  XNOR U30379 ( .A(n21831), .B(n21830), .Z(n21832) );
  XNOR U30380 ( .A(n21827), .B(n21826), .Z(n21830) );
  XOR U30381 ( .A(n21829), .B(n21828), .Z(n21826) );
  XOR U30382 ( .A(y[5288]), .B(x[5288]), .Z(n21828) );
  XOR U30383 ( .A(y[5287]), .B(x[5287]), .Z(n21829) );
  XOR U30384 ( .A(y[5286]), .B(x[5286]), .Z(n21827) );
  XOR U30385 ( .A(n21821), .B(n21820), .Z(n21831) );
  XOR U30386 ( .A(n21823), .B(n21822), .Z(n21820) );
  XOR U30387 ( .A(y[5285]), .B(x[5285]), .Z(n21822) );
  XOR U30388 ( .A(y[5284]), .B(x[5284]), .Z(n21823) );
  XOR U30389 ( .A(y[5283]), .B(x[5283]), .Z(n21821) );
  XNOR U30390 ( .A(n21797), .B(n21798), .Z(n21815) );
  XNOR U30391 ( .A(n21812), .B(n21813), .Z(n21798) );
  XOR U30392 ( .A(n21809), .B(n21808), .Z(n21813) );
  XOR U30393 ( .A(y[5280]), .B(x[5280]), .Z(n21808) );
  XOR U30394 ( .A(n21811), .B(n21810), .Z(n21809) );
  XOR U30395 ( .A(y[5282]), .B(x[5282]), .Z(n21810) );
  XOR U30396 ( .A(y[5281]), .B(x[5281]), .Z(n21811) );
  XOR U30397 ( .A(n21803), .B(n21802), .Z(n21812) );
  XOR U30398 ( .A(n21805), .B(n21804), .Z(n21802) );
  XOR U30399 ( .A(y[5279]), .B(x[5279]), .Z(n21804) );
  XOR U30400 ( .A(y[5278]), .B(x[5278]), .Z(n21805) );
  XOR U30401 ( .A(y[5277]), .B(x[5277]), .Z(n21803) );
  XNOR U30402 ( .A(n21796), .B(n21795), .Z(n21797) );
  XNOR U30403 ( .A(n21792), .B(n21791), .Z(n21795) );
  XOR U30404 ( .A(n21794), .B(n21793), .Z(n21791) );
  XOR U30405 ( .A(y[5276]), .B(x[5276]), .Z(n21793) );
  XOR U30406 ( .A(y[5275]), .B(x[5275]), .Z(n21794) );
  XOR U30407 ( .A(y[5274]), .B(x[5274]), .Z(n21792) );
  XOR U30408 ( .A(n21786), .B(n21785), .Z(n21796) );
  XOR U30409 ( .A(n21788), .B(n21787), .Z(n21785) );
  XOR U30410 ( .A(y[5273]), .B(x[5273]), .Z(n21787) );
  XOR U30411 ( .A(y[5272]), .B(x[5272]), .Z(n21788) );
  XOR U30412 ( .A(y[5271]), .B(x[5271]), .Z(n21786) );
  NAND U30413 ( .A(n21849), .B(n21850), .Z(N63443) );
  NAND U30414 ( .A(n21851), .B(n21852), .Z(n21850) );
  NANDN U30415 ( .A(n21853), .B(n21854), .Z(n21852) );
  NANDN U30416 ( .A(n21854), .B(n21853), .Z(n21849) );
  XOR U30417 ( .A(n21853), .B(n21855), .Z(N63442) );
  XNOR U30418 ( .A(n21851), .B(n21854), .Z(n21855) );
  NAND U30419 ( .A(n21856), .B(n21857), .Z(n21854) );
  NAND U30420 ( .A(n21858), .B(n21859), .Z(n21857) );
  NANDN U30421 ( .A(n21860), .B(n21861), .Z(n21859) );
  NANDN U30422 ( .A(n21861), .B(n21860), .Z(n21856) );
  AND U30423 ( .A(n21862), .B(n21863), .Z(n21851) );
  NAND U30424 ( .A(n21864), .B(n21865), .Z(n21863) );
  NANDN U30425 ( .A(n21866), .B(n21867), .Z(n21865) );
  NANDN U30426 ( .A(n21867), .B(n21866), .Z(n21862) );
  IV U30427 ( .A(n21868), .Z(n21867) );
  AND U30428 ( .A(n21869), .B(n21870), .Z(n21853) );
  NAND U30429 ( .A(n21871), .B(n21872), .Z(n21870) );
  NANDN U30430 ( .A(n21873), .B(n21874), .Z(n21872) );
  NANDN U30431 ( .A(n21874), .B(n21873), .Z(n21869) );
  XOR U30432 ( .A(n21866), .B(n21875), .Z(N63441) );
  XNOR U30433 ( .A(n21864), .B(n21868), .Z(n21875) );
  XOR U30434 ( .A(n21861), .B(n21876), .Z(n21868) );
  XNOR U30435 ( .A(n21858), .B(n21860), .Z(n21876) );
  AND U30436 ( .A(n21877), .B(n21878), .Z(n21860) );
  NANDN U30437 ( .A(n21879), .B(n21880), .Z(n21878) );
  OR U30438 ( .A(n21881), .B(n21882), .Z(n21880) );
  IV U30439 ( .A(n21883), .Z(n21882) );
  NANDN U30440 ( .A(n21883), .B(n21881), .Z(n21877) );
  AND U30441 ( .A(n21884), .B(n21885), .Z(n21858) );
  NAND U30442 ( .A(n21886), .B(n21887), .Z(n21885) );
  NANDN U30443 ( .A(n21888), .B(n21889), .Z(n21887) );
  NANDN U30444 ( .A(n21889), .B(n21888), .Z(n21884) );
  IV U30445 ( .A(n21890), .Z(n21889) );
  NAND U30446 ( .A(n21891), .B(n21892), .Z(n21861) );
  NANDN U30447 ( .A(n21893), .B(n21894), .Z(n21892) );
  NANDN U30448 ( .A(n21895), .B(n21896), .Z(n21894) );
  NANDN U30449 ( .A(n21896), .B(n21895), .Z(n21891) );
  IV U30450 ( .A(n21897), .Z(n21895) );
  AND U30451 ( .A(n21898), .B(n21899), .Z(n21864) );
  NAND U30452 ( .A(n21900), .B(n21901), .Z(n21899) );
  NANDN U30453 ( .A(n21902), .B(n21903), .Z(n21901) );
  NANDN U30454 ( .A(n21903), .B(n21902), .Z(n21898) );
  XOR U30455 ( .A(n21874), .B(n21904), .Z(n21866) );
  XNOR U30456 ( .A(n21871), .B(n21873), .Z(n21904) );
  AND U30457 ( .A(n21905), .B(n21906), .Z(n21873) );
  NANDN U30458 ( .A(n21907), .B(n21908), .Z(n21906) );
  OR U30459 ( .A(n21909), .B(n21910), .Z(n21908) );
  IV U30460 ( .A(n21911), .Z(n21910) );
  NANDN U30461 ( .A(n21911), .B(n21909), .Z(n21905) );
  AND U30462 ( .A(n21912), .B(n21913), .Z(n21871) );
  NAND U30463 ( .A(n21914), .B(n21915), .Z(n21913) );
  NANDN U30464 ( .A(n21916), .B(n21917), .Z(n21915) );
  NANDN U30465 ( .A(n21917), .B(n21916), .Z(n21912) );
  IV U30466 ( .A(n21918), .Z(n21917) );
  NAND U30467 ( .A(n21919), .B(n21920), .Z(n21874) );
  NANDN U30468 ( .A(n21921), .B(n21922), .Z(n21920) );
  NANDN U30469 ( .A(n21923), .B(n21924), .Z(n21922) );
  NANDN U30470 ( .A(n21924), .B(n21923), .Z(n21919) );
  IV U30471 ( .A(n21925), .Z(n21923) );
  XOR U30472 ( .A(n21900), .B(n21926), .Z(N63440) );
  XNOR U30473 ( .A(n21903), .B(n21902), .Z(n21926) );
  XNOR U30474 ( .A(n21914), .B(n21927), .Z(n21902) );
  XNOR U30475 ( .A(n21918), .B(n21916), .Z(n21927) );
  XOR U30476 ( .A(n21924), .B(n21928), .Z(n21916) );
  XNOR U30477 ( .A(n21921), .B(n21925), .Z(n21928) );
  AND U30478 ( .A(n21929), .B(n21930), .Z(n21925) );
  NAND U30479 ( .A(n21931), .B(n21932), .Z(n21930) );
  NAND U30480 ( .A(n21933), .B(n21934), .Z(n21929) );
  AND U30481 ( .A(n21935), .B(n21936), .Z(n21921) );
  NAND U30482 ( .A(n21937), .B(n21938), .Z(n21936) );
  NAND U30483 ( .A(n21939), .B(n21940), .Z(n21935) );
  NANDN U30484 ( .A(n21941), .B(n21942), .Z(n21924) );
  ANDN U30485 ( .B(n21943), .A(n21944), .Z(n21918) );
  XNOR U30486 ( .A(n21909), .B(n21945), .Z(n21914) );
  XNOR U30487 ( .A(n21907), .B(n21911), .Z(n21945) );
  AND U30488 ( .A(n21946), .B(n21947), .Z(n21911) );
  NAND U30489 ( .A(n21948), .B(n21949), .Z(n21947) );
  NAND U30490 ( .A(n21950), .B(n21951), .Z(n21946) );
  AND U30491 ( .A(n21952), .B(n21953), .Z(n21907) );
  NAND U30492 ( .A(n21954), .B(n21955), .Z(n21953) );
  NAND U30493 ( .A(n21956), .B(n21957), .Z(n21952) );
  AND U30494 ( .A(n21958), .B(n21959), .Z(n21909) );
  NAND U30495 ( .A(n21960), .B(n21961), .Z(n21903) );
  XNOR U30496 ( .A(n21886), .B(n21962), .Z(n21900) );
  XNOR U30497 ( .A(n21890), .B(n21888), .Z(n21962) );
  XOR U30498 ( .A(n21896), .B(n21963), .Z(n21888) );
  XNOR U30499 ( .A(n21893), .B(n21897), .Z(n21963) );
  AND U30500 ( .A(n21964), .B(n21965), .Z(n21897) );
  NAND U30501 ( .A(n21966), .B(n21967), .Z(n21965) );
  NAND U30502 ( .A(n21968), .B(n21969), .Z(n21964) );
  AND U30503 ( .A(n21970), .B(n21971), .Z(n21893) );
  NAND U30504 ( .A(n21972), .B(n21973), .Z(n21971) );
  NAND U30505 ( .A(n21974), .B(n21975), .Z(n21970) );
  NANDN U30506 ( .A(n21976), .B(n21977), .Z(n21896) );
  ANDN U30507 ( .B(n21978), .A(n21979), .Z(n21890) );
  XNOR U30508 ( .A(n21881), .B(n21980), .Z(n21886) );
  XNOR U30509 ( .A(n21879), .B(n21883), .Z(n21980) );
  AND U30510 ( .A(n21981), .B(n21982), .Z(n21883) );
  NAND U30511 ( .A(n21983), .B(n21984), .Z(n21982) );
  NAND U30512 ( .A(n21985), .B(n21986), .Z(n21981) );
  AND U30513 ( .A(n21987), .B(n21988), .Z(n21879) );
  NAND U30514 ( .A(n21989), .B(n21990), .Z(n21988) );
  NAND U30515 ( .A(n21991), .B(n21992), .Z(n21987) );
  AND U30516 ( .A(n21993), .B(n21994), .Z(n21881) );
  XOR U30517 ( .A(n21961), .B(n21960), .Z(N63439) );
  XNOR U30518 ( .A(n21978), .B(n21979), .Z(n21960) );
  XNOR U30519 ( .A(n21993), .B(n21994), .Z(n21979) );
  XOR U30520 ( .A(n21990), .B(n21989), .Z(n21994) );
  XOR U30521 ( .A(y[5268]), .B(x[5268]), .Z(n21989) );
  XOR U30522 ( .A(n21992), .B(n21991), .Z(n21990) );
  XOR U30523 ( .A(y[5270]), .B(x[5270]), .Z(n21991) );
  XOR U30524 ( .A(y[5269]), .B(x[5269]), .Z(n21992) );
  XOR U30525 ( .A(n21984), .B(n21983), .Z(n21993) );
  XOR U30526 ( .A(n21986), .B(n21985), .Z(n21983) );
  XOR U30527 ( .A(y[5267]), .B(x[5267]), .Z(n21985) );
  XOR U30528 ( .A(y[5266]), .B(x[5266]), .Z(n21986) );
  XOR U30529 ( .A(y[5265]), .B(x[5265]), .Z(n21984) );
  XNOR U30530 ( .A(n21977), .B(n21976), .Z(n21978) );
  XNOR U30531 ( .A(n21973), .B(n21972), .Z(n21976) );
  XOR U30532 ( .A(n21975), .B(n21974), .Z(n21972) );
  XOR U30533 ( .A(y[5264]), .B(x[5264]), .Z(n21974) );
  XOR U30534 ( .A(y[5263]), .B(x[5263]), .Z(n21975) );
  XOR U30535 ( .A(y[5262]), .B(x[5262]), .Z(n21973) );
  XOR U30536 ( .A(n21967), .B(n21966), .Z(n21977) );
  XOR U30537 ( .A(n21969), .B(n21968), .Z(n21966) );
  XOR U30538 ( .A(y[5261]), .B(x[5261]), .Z(n21968) );
  XOR U30539 ( .A(y[5260]), .B(x[5260]), .Z(n21969) );
  XOR U30540 ( .A(y[5259]), .B(x[5259]), .Z(n21967) );
  XNOR U30541 ( .A(n21943), .B(n21944), .Z(n21961) );
  XNOR U30542 ( .A(n21958), .B(n21959), .Z(n21944) );
  XOR U30543 ( .A(n21955), .B(n21954), .Z(n21959) );
  XOR U30544 ( .A(y[5256]), .B(x[5256]), .Z(n21954) );
  XOR U30545 ( .A(n21957), .B(n21956), .Z(n21955) );
  XOR U30546 ( .A(y[5258]), .B(x[5258]), .Z(n21956) );
  XOR U30547 ( .A(y[5257]), .B(x[5257]), .Z(n21957) );
  XOR U30548 ( .A(n21949), .B(n21948), .Z(n21958) );
  XOR U30549 ( .A(n21951), .B(n21950), .Z(n21948) );
  XOR U30550 ( .A(y[5255]), .B(x[5255]), .Z(n21950) );
  XOR U30551 ( .A(y[5254]), .B(x[5254]), .Z(n21951) );
  XOR U30552 ( .A(y[5253]), .B(x[5253]), .Z(n21949) );
  XNOR U30553 ( .A(n21942), .B(n21941), .Z(n21943) );
  XNOR U30554 ( .A(n21938), .B(n21937), .Z(n21941) );
  XOR U30555 ( .A(n21940), .B(n21939), .Z(n21937) );
  XOR U30556 ( .A(y[5252]), .B(x[5252]), .Z(n21939) );
  XOR U30557 ( .A(y[5251]), .B(x[5251]), .Z(n21940) );
  XOR U30558 ( .A(y[5250]), .B(x[5250]), .Z(n21938) );
  XOR U30559 ( .A(n21932), .B(n21931), .Z(n21942) );
  XOR U30560 ( .A(n21934), .B(n21933), .Z(n21931) );
  XOR U30561 ( .A(y[5249]), .B(x[5249]), .Z(n21933) );
  XOR U30562 ( .A(y[5248]), .B(x[5248]), .Z(n21934) );
  XOR U30563 ( .A(y[5247]), .B(x[5247]), .Z(n21932) );
  NAND U30564 ( .A(n21995), .B(n21996), .Z(N63430) );
  NAND U30565 ( .A(n21997), .B(n21998), .Z(n21996) );
  NANDN U30566 ( .A(n21999), .B(n22000), .Z(n21998) );
  NANDN U30567 ( .A(n22000), .B(n21999), .Z(n21995) );
  XOR U30568 ( .A(n21999), .B(n22001), .Z(N63429) );
  XNOR U30569 ( .A(n21997), .B(n22000), .Z(n22001) );
  NAND U30570 ( .A(n22002), .B(n22003), .Z(n22000) );
  NAND U30571 ( .A(n22004), .B(n22005), .Z(n22003) );
  NANDN U30572 ( .A(n22006), .B(n22007), .Z(n22005) );
  NANDN U30573 ( .A(n22007), .B(n22006), .Z(n22002) );
  AND U30574 ( .A(n22008), .B(n22009), .Z(n21997) );
  NAND U30575 ( .A(n22010), .B(n22011), .Z(n22009) );
  NANDN U30576 ( .A(n22012), .B(n22013), .Z(n22011) );
  NANDN U30577 ( .A(n22013), .B(n22012), .Z(n22008) );
  IV U30578 ( .A(n22014), .Z(n22013) );
  AND U30579 ( .A(n22015), .B(n22016), .Z(n21999) );
  NAND U30580 ( .A(n22017), .B(n22018), .Z(n22016) );
  NANDN U30581 ( .A(n22019), .B(n22020), .Z(n22018) );
  NANDN U30582 ( .A(n22020), .B(n22019), .Z(n22015) );
  XOR U30583 ( .A(n22012), .B(n22021), .Z(N63428) );
  XNOR U30584 ( .A(n22010), .B(n22014), .Z(n22021) );
  XOR U30585 ( .A(n22007), .B(n22022), .Z(n22014) );
  XNOR U30586 ( .A(n22004), .B(n22006), .Z(n22022) );
  AND U30587 ( .A(n22023), .B(n22024), .Z(n22006) );
  NANDN U30588 ( .A(n22025), .B(n22026), .Z(n22024) );
  OR U30589 ( .A(n22027), .B(n22028), .Z(n22026) );
  IV U30590 ( .A(n22029), .Z(n22028) );
  NANDN U30591 ( .A(n22029), .B(n22027), .Z(n22023) );
  AND U30592 ( .A(n22030), .B(n22031), .Z(n22004) );
  NAND U30593 ( .A(n22032), .B(n22033), .Z(n22031) );
  NANDN U30594 ( .A(n22034), .B(n22035), .Z(n22033) );
  NANDN U30595 ( .A(n22035), .B(n22034), .Z(n22030) );
  IV U30596 ( .A(n22036), .Z(n22035) );
  NAND U30597 ( .A(n22037), .B(n22038), .Z(n22007) );
  NANDN U30598 ( .A(n22039), .B(n22040), .Z(n22038) );
  NANDN U30599 ( .A(n22041), .B(n22042), .Z(n22040) );
  NANDN U30600 ( .A(n22042), .B(n22041), .Z(n22037) );
  IV U30601 ( .A(n22043), .Z(n22041) );
  AND U30602 ( .A(n22044), .B(n22045), .Z(n22010) );
  NAND U30603 ( .A(n22046), .B(n22047), .Z(n22045) );
  NANDN U30604 ( .A(n22048), .B(n22049), .Z(n22047) );
  NANDN U30605 ( .A(n22049), .B(n22048), .Z(n22044) );
  XOR U30606 ( .A(n22020), .B(n22050), .Z(n22012) );
  XNOR U30607 ( .A(n22017), .B(n22019), .Z(n22050) );
  AND U30608 ( .A(n22051), .B(n22052), .Z(n22019) );
  NANDN U30609 ( .A(n22053), .B(n22054), .Z(n22052) );
  OR U30610 ( .A(n22055), .B(n22056), .Z(n22054) );
  IV U30611 ( .A(n22057), .Z(n22056) );
  NANDN U30612 ( .A(n22057), .B(n22055), .Z(n22051) );
  AND U30613 ( .A(n22058), .B(n22059), .Z(n22017) );
  NAND U30614 ( .A(n22060), .B(n22061), .Z(n22059) );
  NANDN U30615 ( .A(n22062), .B(n22063), .Z(n22061) );
  NANDN U30616 ( .A(n22063), .B(n22062), .Z(n22058) );
  IV U30617 ( .A(n22064), .Z(n22063) );
  NAND U30618 ( .A(n22065), .B(n22066), .Z(n22020) );
  NANDN U30619 ( .A(n22067), .B(n22068), .Z(n22066) );
  NANDN U30620 ( .A(n22069), .B(n22070), .Z(n22068) );
  NANDN U30621 ( .A(n22070), .B(n22069), .Z(n22065) );
  IV U30622 ( .A(n22071), .Z(n22069) );
  XOR U30623 ( .A(n22046), .B(n22072), .Z(N63427) );
  XNOR U30624 ( .A(n22049), .B(n22048), .Z(n22072) );
  XNOR U30625 ( .A(n22060), .B(n22073), .Z(n22048) );
  XNOR U30626 ( .A(n22064), .B(n22062), .Z(n22073) );
  XOR U30627 ( .A(n22070), .B(n22074), .Z(n22062) );
  XNOR U30628 ( .A(n22067), .B(n22071), .Z(n22074) );
  AND U30629 ( .A(n22075), .B(n22076), .Z(n22071) );
  NAND U30630 ( .A(n22077), .B(n22078), .Z(n22076) );
  NAND U30631 ( .A(n22079), .B(n22080), .Z(n22075) );
  AND U30632 ( .A(n22081), .B(n22082), .Z(n22067) );
  NAND U30633 ( .A(n22083), .B(n22084), .Z(n22082) );
  NAND U30634 ( .A(n22085), .B(n22086), .Z(n22081) );
  NANDN U30635 ( .A(n22087), .B(n22088), .Z(n22070) );
  ANDN U30636 ( .B(n22089), .A(n22090), .Z(n22064) );
  XNOR U30637 ( .A(n22055), .B(n22091), .Z(n22060) );
  XNOR U30638 ( .A(n22053), .B(n22057), .Z(n22091) );
  AND U30639 ( .A(n22092), .B(n22093), .Z(n22057) );
  NAND U30640 ( .A(n22094), .B(n22095), .Z(n22093) );
  NAND U30641 ( .A(n22096), .B(n22097), .Z(n22092) );
  AND U30642 ( .A(n22098), .B(n22099), .Z(n22053) );
  NAND U30643 ( .A(n22100), .B(n22101), .Z(n22099) );
  NAND U30644 ( .A(n22102), .B(n22103), .Z(n22098) );
  AND U30645 ( .A(n22104), .B(n22105), .Z(n22055) );
  NAND U30646 ( .A(n22106), .B(n22107), .Z(n22049) );
  XNOR U30647 ( .A(n22032), .B(n22108), .Z(n22046) );
  XNOR U30648 ( .A(n22036), .B(n22034), .Z(n22108) );
  XOR U30649 ( .A(n22042), .B(n22109), .Z(n22034) );
  XNOR U30650 ( .A(n22039), .B(n22043), .Z(n22109) );
  AND U30651 ( .A(n22110), .B(n22111), .Z(n22043) );
  NAND U30652 ( .A(n22112), .B(n22113), .Z(n22111) );
  NAND U30653 ( .A(n22114), .B(n22115), .Z(n22110) );
  AND U30654 ( .A(n22116), .B(n22117), .Z(n22039) );
  NAND U30655 ( .A(n22118), .B(n22119), .Z(n22117) );
  NAND U30656 ( .A(n22120), .B(n22121), .Z(n22116) );
  NANDN U30657 ( .A(n22122), .B(n22123), .Z(n22042) );
  ANDN U30658 ( .B(n22124), .A(n22125), .Z(n22036) );
  XNOR U30659 ( .A(n22027), .B(n22126), .Z(n22032) );
  XNOR U30660 ( .A(n22025), .B(n22029), .Z(n22126) );
  AND U30661 ( .A(n22127), .B(n22128), .Z(n22029) );
  NAND U30662 ( .A(n22129), .B(n22130), .Z(n22128) );
  NAND U30663 ( .A(n22131), .B(n22132), .Z(n22127) );
  AND U30664 ( .A(n22133), .B(n22134), .Z(n22025) );
  NAND U30665 ( .A(n22135), .B(n22136), .Z(n22134) );
  NAND U30666 ( .A(n22137), .B(n22138), .Z(n22133) );
  AND U30667 ( .A(n22139), .B(n22140), .Z(n22027) );
  XOR U30668 ( .A(n22107), .B(n22106), .Z(N63426) );
  XNOR U30669 ( .A(n22124), .B(n22125), .Z(n22106) );
  XNOR U30670 ( .A(n22139), .B(n22140), .Z(n22125) );
  XOR U30671 ( .A(n22136), .B(n22135), .Z(n22140) );
  XOR U30672 ( .A(y[5244]), .B(x[5244]), .Z(n22135) );
  XOR U30673 ( .A(n22138), .B(n22137), .Z(n22136) );
  XOR U30674 ( .A(y[5246]), .B(x[5246]), .Z(n22137) );
  XOR U30675 ( .A(y[5245]), .B(x[5245]), .Z(n22138) );
  XOR U30676 ( .A(n22130), .B(n22129), .Z(n22139) );
  XOR U30677 ( .A(n22132), .B(n22131), .Z(n22129) );
  XOR U30678 ( .A(y[5243]), .B(x[5243]), .Z(n22131) );
  XOR U30679 ( .A(y[5242]), .B(x[5242]), .Z(n22132) );
  XOR U30680 ( .A(y[5241]), .B(x[5241]), .Z(n22130) );
  XNOR U30681 ( .A(n22123), .B(n22122), .Z(n22124) );
  XNOR U30682 ( .A(n22119), .B(n22118), .Z(n22122) );
  XOR U30683 ( .A(n22121), .B(n22120), .Z(n22118) );
  XOR U30684 ( .A(y[5240]), .B(x[5240]), .Z(n22120) );
  XOR U30685 ( .A(y[5239]), .B(x[5239]), .Z(n22121) );
  XOR U30686 ( .A(y[5238]), .B(x[5238]), .Z(n22119) );
  XOR U30687 ( .A(n22113), .B(n22112), .Z(n22123) );
  XOR U30688 ( .A(n22115), .B(n22114), .Z(n22112) );
  XOR U30689 ( .A(y[5237]), .B(x[5237]), .Z(n22114) );
  XOR U30690 ( .A(y[5236]), .B(x[5236]), .Z(n22115) );
  XOR U30691 ( .A(y[5235]), .B(x[5235]), .Z(n22113) );
  XNOR U30692 ( .A(n22089), .B(n22090), .Z(n22107) );
  XNOR U30693 ( .A(n22104), .B(n22105), .Z(n22090) );
  XOR U30694 ( .A(n22101), .B(n22100), .Z(n22105) );
  XOR U30695 ( .A(y[5232]), .B(x[5232]), .Z(n22100) );
  XOR U30696 ( .A(n22103), .B(n22102), .Z(n22101) );
  XOR U30697 ( .A(y[5234]), .B(x[5234]), .Z(n22102) );
  XOR U30698 ( .A(y[5233]), .B(x[5233]), .Z(n22103) );
  XOR U30699 ( .A(n22095), .B(n22094), .Z(n22104) );
  XOR U30700 ( .A(n22097), .B(n22096), .Z(n22094) );
  XOR U30701 ( .A(y[5231]), .B(x[5231]), .Z(n22096) );
  XOR U30702 ( .A(y[5230]), .B(x[5230]), .Z(n22097) );
  XOR U30703 ( .A(y[5229]), .B(x[5229]), .Z(n22095) );
  XNOR U30704 ( .A(n22088), .B(n22087), .Z(n22089) );
  XNOR U30705 ( .A(n22084), .B(n22083), .Z(n22087) );
  XOR U30706 ( .A(n22086), .B(n22085), .Z(n22083) );
  XOR U30707 ( .A(y[5228]), .B(x[5228]), .Z(n22085) );
  XOR U30708 ( .A(y[5227]), .B(x[5227]), .Z(n22086) );
  XOR U30709 ( .A(y[5226]), .B(x[5226]), .Z(n22084) );
  XOR U30710 ( .A(n22078), .B(n22077), .Z(n22088) );
  XOR U30711 ( .A(n22080), .B(n22079), .Z(n22077) );
  XOR U30712 ( .A(y[5225]), .B(x[5225]), .Z(n22079) );
  XOR U30713 ( .A(y[5224]), .B(x[5224]), .Z(n22080) );
  XOR U30714 ( .A(y[5223]), .B(x[5223]), .Z(n22078) );
  NAND U30715 ( .A(n22141), .B(n22142), .Z(N63417) );
  NAND U30716 ( .A(n22143), .B(n22144), .Z(n22142) );
  NANDN U30717 ( .A(n22145), .B(n22146), .Z(n22144) );
  NANDN U30718 ( .A(n22146), .B(n22145), .Z(n22141) );
  XOR U30719 ( .A(n22145), .B(n22147), .Z(N63416) );
  XNOR U30720 ( .A(n22143), .B(n22146), .Z(n22147) );
  NAND U30721 ( .A(n22148), .B(n22149), .Z(n22146) );
  NAND U30722 ( .A(n22150), .B(n22151), .Z(n22149) );
  NANDN U30723 ( .A(n22152), .B(n22153), .Z(n22151) );
  NANDN U30724 ( .A(n22153), .B(n22152), .Z(n22148) );
  AND U30725 ( .A(n22154), .B(n22155), .Z(n22143) );
  NAND U30726 ( .A(n22156), .B(n22157), .Z(n22155) );
  NANDN U30727 ( .A(n22158), .B(n22159), .Z(n22157) );
  NANDN U30728 ( .A(n22159), .B(n22158), .Z(n22154) );
  IV U30729 ( .A(n22160), .Z(n22159) );
  AND U30730 ( .A(n22161), .B(n22162), .Z(n22145) );
  NAND U30731 ( .A(n22163), .B(n22164), .Z(n22162) );
  NANDN U30732 ( .A(n22165), .B(n22166), .Z(n22164) );
  NANDN U30733 ( .A(n22166), .B(n22165), .Z(n22161) );
  XOR U30734 ( .A(n22158), .B(n22167), .Z(N63415) );
  XNOR U30735 ( .A(n22156), .B(n22160), .Z(n22167) );
  XOR U30736 ( .A(n22153), .B(n22168), .Z(n22160) );
  XNOR U30737 ( .A(n22150), .B(n22152), .Z(n22168) );
  AND U30738 ( .A(n22169), .B(n22170), .Z(n22152) );
  NANDN U30739 ( .A(n22171), .B(n22172), .Z(n22170) );
  OR U30740 ( .A(n22173), .B(n22174), .Z(n22172) );
  IV U30741 ( .A(n22175), .Z(n22174) );
  NANDN U30742 ( .A(n22175), .B(n22173), .Z(n22169) );
  AND U30743 ( .A(n22176), .B(n22177), .Z(n22150) );
  NAND U30744 ( .A(n22178), .B(n22179), .Z(n22177) );
  NANDN U30745 ( .A(n22180), .B(n22181), .Z(n22179) );
  NANDN U30746 ( .A(n22181), .B(n22180), .Z(n22176) );
  IV U30747 ( .A(n22182), .Z(n22181) );
  NAND U30748 ( .A(n22183), .B(n22184), .Z(n22153) );
  NANDN U30749 ( .A(n22185), .B(n22186), .Z(n22184) );
  NANDN U30750 ( .A(n22187), .B(n22188), .Z(n22186) );
  NANDN U30751 ( .A(n22188), .B(n22187), .Z(n22183) );
  IV U30752 ( .A(n22189), .Z(n22187) );
  AND U30753 ( .A(n22190), .B(n22191), .Z(n22156) );
  NAND U30754 ( .A(n22192), .B(n22193), .Z(n22191) );
  NANDN U30755 ( .A(n22194), .B(n22195), .Z(n22193) );
  NANDN U30756 ( .A(n22195), .B(n22194), .Z(n22190) );
  XOR U30757 ( .A(n22166), .B(n22196), .Z(n22158) );
  XNOR U30758 ( .A(n22163), .B(n22165), .Z(n22196) );
  AND U30759 ( .A(n22197), .B(n22198), .Z(n22165) );
  NANDN U30760 ( .A(n22199), .B(n22200), .Z(n22198) );
  OR U30761 ( .A(n22201), .B(n22202), .Z(n22200) );
  IV U30762 ( .A(n22203), .Z(n22202) );
  NANDN U30763 ( .A(n22203), .B(n22201), .Z(n22197) );
  AND U30764 ( .A(n22204), .B(n22205), .Z(n22163) );
  NAND U30765 ( .A(n22206), .B(n22207), .Z(n22205) );
  NANDN U30766 ( .A(n22208), .B(n22209), .Z(n22207) );
  NANDN U30767 ( .A(n22209), .B(n22208), .Z(n22204) );
  IV U30768 ( .A(n22210), .Z(n22209) );
  NAND U30769 ( .A(n22211), .B(n22212), .Z(n22166) );
  NANDN U30770 ( .A(n22213), .B(n22214), .Z(n22212) );
  NANDN U30771 ( .A(n22215), .B(n22216), .Z(n22214) );
  NANDN U30772 ( .A(n22216), .B(n22215), .Z(n22211) );
  IV U30773 ( .A(n22217), .Z(n22215) );
  XOR U30774 ( .A(n22192), .B(n22218), .Z(N63414) );
  XNOR U30775 ( .A(n22195), .B(n22194), .Z(n22218) );
  XNOR U30776 ( .A(n22206), .B(n22219), .Z(n22194) );
  XNOR U30777 ( .A(n22210), .B(n22208), .Z(n22219) );
  XOR U30778 ( .A(n22216), .B(n22220), .Z(n22208) );
  XNOR U30779 ( .A(n22213), .B(n22217), .Z(n22220) );
  AND U30780 ( .A(n22221), .B(n22222), .Z(n22217) );
  NAND U30781 ( .A(n22223), .B(n22224), .Z(n22222) );
  NAND U30782 ( .A(n22225), .B(n22226), .Z(n22221) );
  AND U30783 ( .A(n22227), .B(n22228), .Z(n22213) );
  NAND U30784 ( .A(n22229), .B(n22230), .Z(n22228) );
  NAND U30785 ( .A(n22231), .B(n22232), .Z(n22227) );
  NANDN U30786 ( .A(n22233), .B(n22234), .Z(n22216) );
  ANDN U30787 ( .B(n22235), .A(n22236), .Z(n22210) );
  XNOR U30788 ( .A(n22201), .B(n22237), .Z(n22206) );
  XNOR U30789 ( .A(n22199), .B(n22203), .Z(n22237) );
  AND U30790 ( .A(n22238), .B(n22239), .Z(n22203) );
  NAND U30791 ( .A(n22240), .B(n22241), .Z(n22239) );
  NAND U30792 ( .A(n22242), .B(n22243), .Z(n22238) );
  AND U30793 ( .A(n22244), .B(n22245), .Z(n22199) );
  NAND U30794 ( .A(n22246), .B(n22247), .Z(n22245) );
  NAND U30795 ( .A(n22248), .B(n22249), .Z(n22244) );
  AND U30796 ( .A(n22250), .B(n22251), .Z(n22201) );
  NAND U30797 ( .A(n22252), .B(n22253), .Z(n22195) );
  XNOR U30798 ( .A(n22178), .B(n22254), .Z(n22192) );
  XNOR U30799 ( .A(n22182), .B(n22180), .Z(n22254) );
  XOR U30800 ( .A(n22188), .B(n22255), .Z(n22180) );
  XNOR U30801 ( .A(n22185), .B(n22189), .Z(n22255) );
  AND U30802 ( .A(n22256), .B(n22257), .Z(n22189) );
  NAND U30803 ( .A(n22258), .B(n22259), .Z(n22257) );
  NAND U30804 ( .A(n22260), .B(n22261), .Z(n22256) );
  AND U30805 ( .A(n22262), .B(n22263), .Z(n22185) );
  NAND U30806 ( .A(n22264), .B(n22265), .Z(n22263) );
  NAND U30807 ( .A(n22266), .B(n22267), .Z(n22262) );
  NANDN U30808 ( .A(n22268), .B(n22269), .Z(n22188) );
  ANDN U30809 ( .B(n22270), .A(n22271), .Z(n22182) );
  XNOR U30810 ( .A(n22173), .B(n22272), .Z(n22178) );
  XNOR U30811 ( .A(n22171), .B(n22175), .Z(n22272) );
  AND U30812 ( .A(n22273), .B(n22274), .Z(n22175) );
  NAND U30813 ( .A(n22275), .B(n22276), .Z(n22274) );
  NAND U30814 ( .A(n22277), .B(n22278), .Z(n22273) );
  AND U30815 ( .A(n22279), .B(n22280), .Z(n22171) );
  NAND U30816 ( .A(n22281), .B(n22282), .Z(n22280) );
  NAND U30817 ( .A(n22283), .B(n22284), .Z(n22279) );
  AND U30818 ( .A(n22285), .B(n22286), .Z(n22173) );
  XOR U30819 ( .A(n22253), .B(n22252), .Z(N63413) );
  XNOR U30820 ( .A(n22270), .B(n22271), .Z(n22252) );
  XNOR U30821 ( .A(n22285), .B(n22286), .Z(n22271) );
  XOR U30822 ( .A(n22282), .B(n22281), .Z(n22286) );
  XOR U30823 ( .A(y[5220]), .B(x[5220]), .Z(n22281) );
  XOR U30824 ( .A(n22284), .B(n22283), .Z(n22282) );
  XOR U30825 ( .A(y[5222]), .B(x[5222]), .Z(n22283) );
  XOR U30826 ( .A(y[5221]), .B(x[5221]), .Z(n22284) );
  XOR U30827 ( .A(n22276), .B(n22275), .Z(n22285) );
  XOR U30828 ( .A(n22278), .B(n22277), .Z(n22275) );
  XOR U30829 ( .A(y[5219]), .B(x[5219]), .Z(n22277) );
  XOR U30830 ( .A(y[5218]), .B(x[5218]), .Z(n22278) );
  XOR U30831 ( .A(y[5217]), .B(x[5217]), .Z(n22276) );
  XNOR U30832 ( .A(n22269), .B(n22268), .Z(n22270) );
  XNOR U30833 ( .A(n22265), .B(n22264), .Z(n22268) );
  XOR U30834 ( .A(n22267), .B(n22266), .Z(n22264) );
  XOR U30835 ( .A(y[5216]), .B(x[5216]), .Z(n22266) );
  XOR U30836 ( .A(y[5215]), .B(x[5215]), .Z(n22267) );
  XOR U30837 ( .A(y[5214]), .B(x[5214]), .Z(n22265) );
  XOR U30838 ( .A(n22259), .B(n22258), .Z(n22269) );
  XOR U30839 ( .A(n22261), .B(n22260), .Z(n22258) );
  XOR U30840 ( .A(y[5213]), .B(x[5213]), .Z(n22260) );
  XOR U30841 ( .A(y[5212]), .B(x[5212]), .Z(n22261) );
  XOR U30842 ( .A(y[5211]), .B(x[5211]), .Z(n22259) );
  XNOR U30843 ( .A(n22235), .B(n22236), .Z(n22253) );
  XNOR U30844 ( .A(n22250), .B(n22251), .Z(n22236) );
  XOR U30845 ( .A(n22247), .B(n22246), .Z(n22251) );
  XOR U30846 ( .A(y[5208]), .B(x[5208]), .Z(n22246) );
  XOR U30847 ( .A(n22249), .B(n22248), .Z(n22247) );
  XOR U30848 ( .A(y[5210]), .B(x[5210]), .Z(n22248) );
  XOR U30849 ( .A(y[5209]), .B(x[5209]), .Z(n22249) );
  XOR U30850 ( .A(n22241), .B(n22240), .Z(n22250) );
  XOR U30851 ( .A(n22243), .B(n22242), .Z(n22240) );
  XOR U30852 ( .A(y[5207]), .B(x[5207]), .Z(n22242) );
  XOR U30853 ( .A(y[5206]), .B(x[5206]), .Z(n22243) );
  XOR U30854 ( .A(y[5205]), .B(x[5205]), .Z(n22241) );
  XNOR U30855 ( .A(n22234), .B(n22233), .Z(n22235) );
  XNOR U30856 ( .A(n22230), .B(n22229), .Z(n22233) );
  XOR U30857 ( .A(n22232), .B(n22231), .Z(n22229) );
  XOR U30858 ( .A(y[5204]), .B(x[5204]), .Z(n22231) );
  XOR U30859 ( .A(y[5203]), .B(x[5203]), .Z(n22232) );
  XOR U30860 ( .A(y[5202]), .B(x[5202]), .Z(n22230) );
  XOR U30861 ( .A(n22224), .B(n22223), .Z(n22234) );
  XOR U30862 ( .A(n22226), .B(n22225), .Z(n22223) );
  XOR U30863 ( .A(y[5201]), .B(x[5201]), .Z(n22225) );
  XOR U30864 ( .A(y[5200]), .B(x[5200]), .Z(n22226) );
  XOR U30865 ( .A(y[5199]), .B(x[5199]), .Z(n22224) );
  NAND U30866 ( .A(n22287), .B(n22288), .Z(N63404) );
  NAND U30867 ( .A(n22289), .B(n22290), .Z(n22288) );
  NANDN U30868 ( .A(n22291), .B(n22292), .Z(n22290) );
  NANDN U30869 ( .A(n22292), .B(n22291), .Z(n22287) );
  XOR U30870 ( .A(n22291), .B(n22293), .Z(N63403) );
  XNOR U30871 ( .A(n22289), .B(n22292), .Z(n22293) );
  NAND U30872 ( .A(n22294), .B(n22295), .Z(n22292) );
  NAND U30873 ( .A(n22296), .B(n22297), .Z(n22295) );
  NANDN U30874 ( .A(n22298), .B(n22299), .Z(n22297) );
  NANDN U30875 ( .A(n22299), .B(n22298), .Z(n22294) );
  AND U30876 ( .A(n22300), .B(n22301), .Z(n22289) );
  NAND U30877 ( .A(n22302), .B(n22303), .Z(n22301) );
  NANDN U30878 ( .A(n22304), .B(n22305), .Z(n22303) );
  NANDN U30879 ( .A(n22305), .B(n22304), .Z(n22300) );
  IV U30880 ( .A(n22306), .Z(n22305) );
  AND U30881 ( .A(n22307), .B(n22308), .Z(n22291) );
  NAND U30882 ( .A(n22309), .B(n22310), .Z(n22308) );
  NANDN U30883 ( .A(n22311), .B(n22312), .Z(n22310) );
  NANDN U30884 ( .A(n22312), .B(n22311), .Z(n22307) );
  XOR U30885 ( .A(n22304), .B(n22313), .Z(N63402) );
  XNOR U30886 ( .A(n22302), .B(n22306), .Z(n22313) );
  XOR U30887 ( .A(n22299), .B(n22314), .Z(n22306) );
  XNOR U30888 ( .A(n22296), .B(n22298), .Z(n22314) );
  AND U30889 ( .A(n22315), .B(n22316), .Z(n22298) );
  NANDN U30890 ( .A(n22317), .B(n22318), .Z(n22316) );
  OR U30891 ( .A(n22319), .B(n22320), .Z(n22318) );
  IV U30892 ( .A(n22321), .Z(n22320) );
  NANDN U30893 ( .A(n22321), .B(n22319), .Z(n22315) );
  AND U30894 ( .A(n22322), .B(n22323), .Z(n22296) );
  NAND U30895 ( .A(n22324), .B(n22325), .Z(n22323) );
  NANDN U30896 ( .A(n22326), .B(n22327), .Z(n22325) );
  NANDN U30897 ( .A(n22327), .B(n22326), .Z(n22322) );
  IV U30898 ( .A(n22328), .Z(n22327) );
  NAND U30899 ( .A(n22329), .B(n22330), .Z(n22299) );
  NANDN U30900 ( .A(n22331), .B(n22332), .Z(n22330) );
  NANDN U30901 ( .A(n22333), .B(n22334), .Z(n22332) );
  NANDN U30902 ( .A(n22334), .B(n22333), .Z(n22329) );
  IV U30903 ( .A(n22335), .Z(n22333) );
  AND U30904 ( .A(n22336), .B(n22337), .Z(n22302) );
  NAND U30905 ( .A(n22338), .B(n22339), .Z(n22337) );
  NANDN U30906 ( .A(n22340), .B(n22341), .Z(n22339) );
  NANDN U30907 ( .A(n22341), .B(n22340), .Z(n22336) );
  XOR U30908 ( .A(n22312), .B(n22342), .Z(n22304) );
  XNOR U30909 ( .A(n22309), .B(n22311), .Z(n22342) );
  AND U30910 ( .A(n22343), .B(n22344), .Z(n22311) );
  NANDN U30911 ( .A(n22345), .B(n22346), .Z(n22344) );
  OR U30912 ( .A(n22347), .B(n22348), .Z(n22346) );
  IV U30913 ( .A(n22349), .Z(n22348) );
  NANDN U30914 ( .A(n22349), .B(n22347), .Z(n22343) );
  AND U30915 ( .A(n22350), .B(n22351), .Z(n22309) );
  NAND U30916 ( .A(n22352), .B(n22353), .Z(n22351) );
  NANDN U30917 ( .A(n22354), .B(n22355), .Z(n22353) );
  NANDN U30918 ( .A(n22355), .B(n22354), .Z(n22350) );
  IV U30919 ( .A(n22356), .Z(n22355) );
  NAND U30920 ( .A(n22357), .B(n22358), .Z(n22312) );
  NANDN U30921 ( .A(n22359), .B(n22360), .Z(n22358) );
  NANDN U30922 ( .A(n22361), .B(n22362), .Z(n22360) );
  NANDN U30923 ( .A(n22362), .B(n22361), .Z(n22357) );
  IV U30924 ( .A(n22363), .Z(n22361) );
  XOR U30925 ( .A(n22338), .B(n22364), .Z(N63401) );
  XNOR U30926 ( .A(n22341), .B(n22340), .Z(n22364) );
  XNOR U30927 ( .A(n22352), .B(n22365), .Z(n22340) );
  XNOR U30928 ( .A(n22356), .B(n22354), .Z(n22365) );
  XOR U30929 ( .A(n22362), .B(n22366), .Z(n22354) );
  XNOR U30930 ( .A(n22359), .B(n22363), .Z(n22366) );
  AND U30931 ( .A(n22367), .B(n22368), .Z(n22363) );
  NAND U30932 ( .A(n22369), .B(n22370), .Z(n22368) );
  NAND U30933 ( .A(n22371), .B(n22372), .Z(n22367) );
  AND U30934 ( .A(n22373), .B(n22374), .Z(n22359) );
  NAND U30935 ( .A(n22375), .B(n22376), .Z(n22374) );
  NAND U30936 ( .A(n22377), .B(n22378), .Z(n22373) );
  NANDN U30937 ( .A(n22379), .B(n22380), .Z(n22362) );
  ANDN U30938 ( .B(n22381), .A(n22382), .Z(n22356) );
  XNOR U30939 ( .A(n22347), .B(n22383), .Z(n22352) );
  XNOR U30940 ( .A(n22345), .B(n22349), .Z(n22383) );
  AND U30941 ( .A(n22384), .B(n22385), .Z(n22349) );
  NAND U30942 ( .A(n22386), .B(n22387), .Z(n22385) );
  NAND U30943 ( .A(n22388), .B(n22389), .Z(n22384) );
  AND U30944 ( .A(n22390), .B(n22391), .Z(n22345) );
  NAND U30945 ( .A(n22392), .B(n22393), .Z(n22391) );
  NAND U30946 ( .A(n22394), .B(n22395), .Z(n22390) );
  AND U30947 ( .A(n22396), .B(n22397), .Z(n22347) );
  NAND U30948 ( .A(n22398), .B(n22399), .Z(n22341) );
  XNOR U30949 ( .A(n22324), .B(n22400), .Z(n22338) );
  XNOR U30950 ( .A(n22328), .B(n22326), .Z(n22400) );
  XOR U30951 ( .A(n22334), .B(n22401), .Z(n22326) );
  XNOR U30952 ( .A(n22331), .B(n22335), .Z(n22401) );
  AND U30953 ( .A(n22402), .B(n22403), .Z(n22335) );
  NAND U30954 ( .A(n22404), .B(n22405), .Z(n22403) );
  NAND U30955 ( .A(n22406), .B(n22407), .Z(n22402) );
  AND U30956 ( .A(n22408), .B(n22409), .Z(n22331) );
  NAND U30957 ( .A(n22410), .B(n22411), .Z(n22409) );
  NAND U30958 ( .A(n22412), .B(n22413), .Z(n22408) );
  NANDN U30959 ( .A(n22414), .B(n22415), .Z(n22334) );
  ANDN U30960 ( .B(n22416), .A(n22417), .Z(n22328) );
  XNOR U30961 ( .A(n22319), .B(n22418), .Z(n22324) );
  XNOR U30962 ( .A(n22317), .B(n22321), .Z(n22418) );
  AND U30963 ( .A(n22419), .B(n22420), .Z(n22321) );
  NAND U30964 ( .A(n22421), .B(n22422), .Z(n22420) );
  NAND U30965 ( .A(n22423), .B(n22424), .Z(n22419) );
  AND U30966 ( .A(n22425), .B(n22426), .Z(n22317) );
  NAND U30967 ( .A(n22427), .B(n22428), .Z(n22426) );
  NAND U30968 ( .A(n22429), .B(n22430), .Z(n22425) );
  AND U30969 ( .A(n22431), .B(n22432), .Z(n22319) );
  XOR U30970 ( .A(n22399), .B(n22398), .Z(N63400) );
  XNOR U30971 ( .A(n22416), .B(n22417), .Z(n22398) );
  XNOR U30972 ( .A(n22431), .B(n22432), .Z(n22417) );
  XOR U30973 ( .A(n22428), .B(n22427), .Z(n22432) );
  XOR U30974 ( .A(y[5196]), .B(x[5196]), .Z(n22427) );
  XOR U30975 ( .A(n22430), .B(n22429), .Z(n22428) );
  XOR U30976 ( .A(y[5198]), .B(x[5198]), .Z(n22429) );
  XOR U30977 ( .A(y[5197]), .B(x[5197]), .Z(n22430) );
  XOR U30978 ( .A(n22422), .B(n22421), .Z(n22431) );
  XOR U30979 ( .A(n22424), .B(n22423), .Z(n22421) );
  XOR U30980 ( .A(y[5195]), .B(x[5195]), .Z(n22423) );
  XOR U30981 ( .A(y[5194]), .B(x[5194]), .Z(n22424) );
  XOR U30982 ( .A(y[5193]), .B(x[5193]), .Z(n22422) );
  XNOR U30983 ( .A(n22415), .B(n22414), .Z(n22416) );
  XNOR U30984 ( .A(n22411), .B(n22410), .Z(n22414) );
  XOR U30985 ( .A(n22413), .B(n22412), .Z(n22410) );
  XOR U30986 ( .A(y[5192]), .B(x[5192]), .Z(n22412) );
  XOR U30987 ( .A(y[5191]), .B(x[5191]), .Z(n22413) );
  XOR U30988 ( .A(y[5190]), .B(x[5190]), .Z(n22411) );
  XOR U30989 ( .A(n22405), .B(n22404), .Z(n22415) );
  XOR U30990 ( .A(n22407), .B(n22406), .Z(n22404) );
  XOR U30991 ( .A(y[5189]), .B(x[5189]), .Z(n22406) );
  XOR U30992 ( .A(y[5188]), .B(x[5188]), .Z(n22407) );
  XOR U30993 ( .A(y[5187]), .B(x[5187]), .Z(n22405) );
  XNOR U30994 ( .A(n22381), .B(n22382), .Z(n22399) );
  XNOR U30995 ( .A(n22396), .B(n22397), .Z(n22382) );
  XOR U30996 ( .A(n22393), .B(n22392), .Z(n22397) );
  XOR U30997 ( .A(y[5184]), .B(x[5184]), .Z(n22392) );
  XOR U30998 ( .A(n22395), .B(n22394), .Z(n22393) );
  XOR U30999 ( .A(y[5186]), .B(x[5186]), .Z(n22394) );
  XOR U31000 ( .A(y[5185]), .B(x[5185]), .Z(n22395) );
  XOR U31001 ( .A(n22387), .B(n22386), .Z(n22396) );
  XOR U31002 ( .A(n22389), .B(n22388), .Z(n22386) );
  XOR U31003 ( .A(y[5183]), .B(x[5183]), .Z(n22388) );
  XOR U31004 ( .A(y[5182]), .B(x[5182]), .Z(n22389) );
  XOR U31005 ( .A(y[5181]), .B(x[5181]), .Z(n22387) );
  XNOR U31006 ( .A(n22380), .B(n22379), .Z(n22381) );
  XNOR U31007 ( .A(n22376), .B(n22375), .Z(n22379) );
  XOR U31008 ( .A(n22378), .B(n22377), .Z(n22375) );
  XOR U31009 ( .A(y[5180]), .B(x[5180]), .Z(n22377) );
  XOR U31010 ( .A(y[5179]), .B(x[5179]), .Z(n22378) );
  XOR U31011 ( .A(y[5178]), .B(x[5178]), .Z(n22376) );
  XOR U31012 ( .A(n22370), .B(n22369), .Z(n22380) );
  XOR U31013 ( .A(n22372), .B(n22371), .Z(n22369) );
  XOR U31014 ( .A(y[5177]), .B(x[5177]), .Z(n22371) );
  XOR U31015 ( .A(y[5176]), .B(x[5176]), .Z(n22372) );
  XOR U31016 ( .A(y[5175]), .B(x[5175]), .Z(n22370) );
  NAND U31017 ( .A(n22433), .B(n22434), .Z(N63391) );
  NAND U31018 ( .A(n22435), .B(n22436), .Z(n22434) );
  NANDN U31019 ( .A(n22437), .B(n22438), .Z(n22436) );
  NANDN U31020 ( .A(n22438), .B(n22437), .Z(n22433) );
  XOR U31021 ( .A(n22437), .B(n22439), .Z(N63390) );
  XNOR U31022 ( .A(n22435), .B(n22438), .Z(n22439) );
  NAND U31023 ( .A(n22440), .B(n22441), .Z(n22438) );
  NAND U31024 ( .A(n22442), .B(n22443), .Z(n22441) );
  NANDN U31025 ( .A(n22444), .B(n22445), .Z(n22443) );
  NANDN U31026 ( .A(n22445), .B(n22444), .Z(n22440) );
  AND U31027 ( .A(n22446), .B(n22447), .Z(n22435) );
  NAND U31028 ( .A(n22448), .B(n22449), .Z(n22447) );
  NANDN U31029 ( .A(n22450), .B(n22451), .Z(n22449) );
  NANDN U31030 ( .A(n22451), .B(n22450), .Z(n22446) );
  IV U31031 ( .A(n22452), .Z(n22451) );
  AND U31032 ( .A(n22453), .B(n22454), .Z(n22437) );
  NAND U31033 ( .A(n22455), .B(n22456), .Z(n22454) );
  NANDN U31034 ( .A(n22457), .B(n22458), .Z(n22456) );
  NANDN U31035 ( .A(n22458), .B(n22457), .Z(n22453) );
  XOR U31036 ( .A(n22450), .B(n22459), .Z(N63389) );
  XNOR U31037 ( .A(n22448), .B(n22452), .Z(n22459) );
  XOR U31038 ( .A(n22445), .B(n22460), .Z(n22452) );
  XNOR U31039 ( .A(n22442), .B(n22444), .Z(n22460) );
  AND U31040 ( .A(n22461), .B(n22462), .Z(n22444) );
  NANDN U31041 ( .A(n22463), .B(n22464), .Z(n22462) );
  OR U31042 ( .A(n22465), .B(n22466), .Z(n22464) );
  IV U31043 ( .A(n22467), .Z(n22466) );
  NANDN U31044 ( .A(n22467), .B(n22465), .Z(n22461) );
  AND U31045 ( .A(n22468), .B(n22469), .Z(n22442) );
  NAND U31046 ( .A(n22470), .B(n22471), .Z(n22469) );
  NANDN U31047 ( .A(n22472), .B(n22473), .Z(n22471) );
  NANDN U31048 ( .A(n22473), .B(n22472), .Z(n22468) );
  IV U31049 ( .A(n22474), .Z(n22473) );
  NAND U31050 ( .A(n22475), .B(n22476), .Z(n22445) );
  NANDN U31051 ( .A(n22477), .B(n22478), .Z(n22476) );
  NANDN U31052 ( .A(n22479), .B(n22480), .Z(n22478) );
  NANDN U31053 ( .A(n22480), .B(n22479), .Z(n22475) );
  IV U31054 ( .A(n22481), .Z(n22479) );
  AND U31055 ( .A(n22482), .B(n22483), .Z(n22448) );
  NAND U31056 ( .A(n22484), .B(n22485), .Z(n22483) );
  NANDN U31057 ( .A(n22486), .B(n22487), .Z(n22485) );
  NANDN U31058 ( .A(n22487), .B(n22486), .Z(n22482) );
  XOR U31059 ( .A(n22458), .B(n22488), .Z(n22450) );
  XNOR U31060 ( .A(n22455), .B(n22457), .Z(n22488) );
  AND U31061 ( .A(n22489), .B(n22490), .Z(n22457) );
  NANDN U31062 ( .A(n22491), .B(n22492), .Z(n22490) );
  OR U31063 ( .A(n22493), .B(n22494), .Z(n22492) );
  IV U31064 ( .A(n22495), .Z(n22494) );
  NANDN U31065 ( .A(n22495), .B(n22493), .Z(n22489) );
  AND U31066 ( .A(n22496), .B(n22497), .Z(n22455) );
  NAND U31067 ( .A(n22498), .B(n22499), .Z(n22497) );
  NANDN U31068 ( .A(n22500), .B(n22501), .Z(n22499) );
  NANDN U31069 ( .A(n22501), .B(n22500), .Z(n22496) );
  IV U31070 ( .A(n22502), .Z(n22501) );
  NAND U31071 ( .A(n22503), .B(n22504), .Z(n22458) );
  NANDN U31072 ( .A(n22505), .B(n22506), .Z(n22504) );
  NANDN U31073 ( .A(n22507), .B(n22508), .Z(n22506) );
  NANDN U31074 ( .A(n22508), .B(n22507), .Z(n22503) );
  IV U31075 ( .A(n22509), .Z(n22507) );
  XOR U31076 ( .A(n22484), .B(n22510), .Z(N63388) );
  XNOR U31077 ( .A(n22487), .B(n22486), .Z(n22510) );
  XNOR U31078 ( .A(n22498), .B(n22511), .Z(n22486) );
  XNOR U31079 ( .A(n22502), .B(n22500), .Z(n22511) );
  XOR U31080 ( .A(n22508), .B(n22512), .Z(n22500) );
  XNOR U31081 ( .A(n22505), .B(n22509), .Z(n22512) );
  AND U31082 ( .A(n22513), .B(n22514), .Z(n22509) );
  NAND U31083 ( .A(n22515), .B(n22516), .Z(n22514) );
  NAND U31084 ( .A(n22517), .B(n22518), .Z(n22513) );
  AND U31085 ( .A(n22519), .B(n22520), .Z(n22505) );
  NAND U31086 ( .A(n22521), .B(n22522), .Z(n22520) );
  NAND U31087 ( .A(n22523), .B(n22524), .Z(n22519) );
  NANDN U31088 ( .A(n22525), .B(n22526), .Z(n22508) );
  ANDN U31089 ( .B(n22527), .A(n22528), .Z(n22502) );
  XNOR U31090 ( .A(n22493), .B(n22529), .Z(n22498) );
  XNOR U31091 ( .A(n22491), .B(n22495), .Z(n22529) );
  AND U31092 ( .A(n22530), .B(n22531), .Z(n22495) );
  NAND U31093 ( .A(n22532), .B(n22533), .Z(n22531) );
  NAND U31094 ( .A(n22534), .B(n22535), .Z(n22530) );
  AND U31095 ( .A(n22536), .B(n22537), .Z(n22491) );
  NAND U31096 ( .A(n22538), .B(n22539), .Z(n22537) );
  NAND U31097 ( .A(n22540), .B(n22541), .Z(n22536) );
  AND U31098 ( .A(n22542), .B(n22543), .Z(n22493) );
  NAND U31099 ( .A(n22544), .B(n22545), .Z(n22487) );
  XNOR U31100 ( .A(n22470), .B(n22546), .Z(n22484) );
  XNOR U31101 ( .A(n22474), .B(n22472), .Z(n22546) );
  XOR U31102 ( .A(n22480), .B(n22547), .Z(n22472) );
  XNOR U31103 ( .A(n22477), .B(n22481), .Z(n22547) );
  AND U31104 ( .A(n22548), .B(n22549), .Z(n22481) );
  NAND U31105 ( .A(n22550), .B(n22551), .Z(n22549) );
  NAND U31106 ( .A(n22552), .B(n22553), .Z(n22548) );
  AND U31107 ( .A(n22554), .B(n22555), .Z(n22477) );
  NAND U31108 ( .A(n22556), .B(n22557), .Z(n22555) );
  NAND U31109 ( .A(n22558), .B(n22559), .Z(n22554) );
  NANDN U31110 ( .A(n22560), .B(n22561), .Z(n22480) );
  ANDN U31111 ( .B(n22562), .A(n22563), .Z(n22474) );
  XNOR U31112 ( .A(n22465), .B(n22564), .Z(n22470) );
  XNOR U31113 ( .A(n22463), .B(n22467), .Z(n22564) );
  AND U31114 ( .A(n22565), .B(n22566), .Z(n22467) );
  NAND U31115 ( .A(n22567), .B(n22568), .Z(n22566) );
  NAND U31116 ( .A(n22569), .B(n22570), .Z(n22565) );
  AND U31117 ( .A(n22571), .B(n22572), .Z(n22463) );
  NAND U31118 ( .A(n22573), .B(n22574), .Z(n22572) );
  NAND U31119 ( .A(n22575), .B(n22576), .Z(n22571) );
  AND U31120 ( .A(n22577), .B(n22578), .Z(n22465) );
  XOR U31121 ( .A(n22545), .B(n22544), .Z(N63387) );
  XNOR U31122 ( .A(n22562), .B(n22563), .Z(n22544) );
  XNOR U31123 ( .A(n22577), .B(n22578), .Z(n22563) );
  XOR U31124 ( .A(n22574), .B(n22573), .Z(n22578) );
  XOR U31125 ( .A(y[5172]), .B(x[5172]), .Z(n22573) );
  XOR U31126 ( .A(n22576), .B(n22575), .Z(n22574) );
  XOR U31127 ( .A(y[5174]), .B(x[5174]), .Z(n22575) );
  XOR U31128 ( .A(y[5173]), .B(x[5173]), .Z(n22576) );
  XOR U31129 ( .A(n22568), .B(n22567), .Z(n22577) );
  XOR U31130 ( .A(n22570), .B(n22569), .Z(n22567) );
  XOR U31131 ( .A(y[5171]), .B(x[5171]), .Z(n22569) );
  XOR U31132 ( .A(y[5170]), .B(x[5170]), .Z(n22570) );
  XOR U31133 ( .A(y[5169]), .B(x[5169]), .Z(n22568) );
  XNOR U31134 ( .A(n22561), .B(n22560), .Z(n22562) );
  XNOR U31135 ( .A(n22557), .B(n22556), .Z(n22560) );
  XOR U31136 ( .A(n22559), .B(n22558), .Z(n22556) );
  XOR U31137 ( .A(y[5168]), .B(x[5168]), .Z(n22558) );
  XOR U31138 ( .A(y[5167]), .B(x[5167]), .Z(n22559) );
  XOR U31139 ( .A(y[5166]), .B(x[5166]), .Z(n22557) );
  XOR U31140 ( .A(n22551), .B(n22550), .Z(n22561) );
  XOR U31141 ( .A(n22553), .B(n22552), .Z(n22550) );
  XOR U31142 ( .A(y[5165]), .B(x[5165]), .Z(n22552) );
  XOR U31143 ( .A(y[5164]), .B(x[5164]), .Z(n22553) );
  XOR U31144 ( .A(y[5163]), .B(x[5163]), .Z(n22551) );
  XNOR U31145 ( .A(n22527), .B(n22528), .Z(n22545) );
  XNOR U31146 ( .A(n22542), .B(n22543), .Z(n22528) );
  XOR U31147 ( .A(n22539), .B(n22538), .Z(n22543) );
  XOR U31148 ( .A(y[5160]), .B(x[5160]), .Z(n22538) );
  XOR U31149 ( .A(n22541), .B(n22540), .Z(n22539) );
  XOR U31150 ( .A(y[5162]), .B(x[5162]), .Z(n22540) );
  XOR U31151 ( .A(y[5161]), .B(x[5161]), .Z(n22541) );
  XOR U31152 ( .A(n22533), .B(n22532), .Z(n22542) );
  XOR U31153 ( .A(n22535), .B(n22534), .Z(n22532) );
  XOR U31154 ( .A(y[5159]), .B(x[5159]), .Z(n22534) );
  XOR U31155 ( .A(y[5158]), .B(x[5158]), .Z(n22535) );
  XOR U31156 ( .A(y[5157]), .B(x[5157]), .Z(n22533) );
  XNOR U31157 ( .A(n22526), .B(n22525), .Z(n22527) );
  XNOR U31158 ( .A(n22522), .B(n22521), .Z(n22525) );
  XOR U31159 ( .A(n22524), .B(n22523), .Z(n22521) );
  XOR U31160 ( .A(y[5156]), .B(x[5156]), .Z(n22523) );
  XOR U31161 ( .A(y[5155]), .B(x[5155]), .Z(n22524) );
  XOR U31162 ( .A(y[5154]), .B(x[5154]), .Z(n22522) );
  XOR U31163 ( .A(n22516), .B(n22515), .Z(n22526) );
  XOR U31164 ( .A(n22518), .B(n22517), .Z(n22515) );
  XOR U31165 ( .A(y[5153]), .B(x[5153]), .Z(n22517) );
  XOR U31166 ( .A(y[5152]), .B(x[5152]), .Z(n22518) );
  XOR U31167 ( .A(y[5151]), .B(x[5151]), .Z(n22516) );
  NAND U31168 ( .A(n22579), .B(n22580), .Z(N63378) );
  NAND U31169 ( .A(n22581), .B(n22582), .Z(n22580) );
  NANDN U31170 ( .A(n22583), .B(n22584), .Z(n22582) );
  NANDN U31171 ( .A(n22584), .B(n22583), .Z(n22579) );
  XOR U31172 ( .A(n22583), .B(n22585), .Z(N63377) );
  XNOR U31173 ( .A(n22581), .B(n22584), .Z(n22585) );
  NAND U31174 ( .A(n22586), .B(n22587), .Z(n22584) );
  NAND U31175 ( .A(n22588), .B(n22589), .Z(n22587) );
  NANDN U31176 ( .A(n22590), .B(n22591), .Z(n22589) );
  NANDN U31177 ( .A(n22591), .B(n22590), .Z(n22586) );
  AND U31178 ( .A(n22592), .B(n22593), .Z(n22581) );
  NAND U31179 ( .A(n22594), .B(n22595), .Z(n22593) );
  NANDN U31180 ( .A(n22596), .B(n22597), .Z(n22595) );
  NANDN U31181 ( .A(n22597), .B(n22596), .Z(n22592) );
  IV U31182 ( .A(n22598), .Z(n22597) );
  AND U31183 ( .A(n22599), .B(n22600), .Z(n22583) );
  NAND U31184 ( .A(n22601), .B(n22602), .Z(n22600) );
  NANDN U31185 ( .A(n22603), .B(n22604), .Z(n22602) );
  NANDN U31186 ( .A(n22604), .B(n22603), .Z(n22599) );
  XOR U31187 ( .A(n22596), .B(n22605), .Z(N63376) );
  XNOR U31188 ( .A(n22594), .B(n22598), .Z(n22605) );
  XOR U31189 ( .A(n22591), .B(n22606), .Z(n22598) );
  XNOR U31190 ( .A(n22588), .B(n22590), .Z(n22606) );
  AND U31191 ( .A(n22607), .B(n22608), .Z(n22590) );
  NANDN U31192 ( .A(n22609), .B(n22610), .Z(n22608) );
  OR U31193 ( .A(n22611), .B(n22612), .Z(n22610) );
  IV U31194 ( .A(n22613), .Z(n22612) );
  NANDN U31195 ( .A(n22613), .B(n22611), .Z(n22607) );
  AND U31196 ( .A(n22614), .B(n22615), .Z(n22588) );
  NAND U31197 ( .A(n22616), .B(n22617), .Z(n22615) );
  NANDN U31198 ( .A(n22618), .B(n22619), .Z(n22617) );
  NANDN U31199 ( .A(n22619), .B(n22618), .Z(n22614) );
  IV U31200 ( .A(n22620), .Z(n22619) );
  NAND U31201 ( .A(n22621), .B(n22622), .Z(n22591) );
  NANDN U31202 ( .A(n22623), .B(n22624), .Z(n22622) );
  NANDN U31203 ( .A(n22625), .B(n22626), .Z(n22624) );
  NANDN U31204 ( .A(n22626), .B(n22625), .Z(n22621) );
  IV U31205 ( .A(n22627), .Z(n22625) );
  AND U31206 ( .A(n22628), .B(n22629), .Z(n22594) );
  NAND U31207 ( .A(n22630), .B(n22631), .Z(n22629) );
  NANDN U31208 ( .A(n22632), .B(n22633), .Z(n22631) );
  NANDN U31209 ( .A(n22633), .B(n22632), .Z(n22628) );
  XOR U31210 ( .A(n22604), .B(n22634), .Z(n22596) );
  XNOR U31211 ( .A(n22601), .B(n22603), .Z(n22634) );
  AND U31212 ( .A(n22635), .B(n22636), .Z(n22603) );
  NANDN U31213 ( .A(n22637), .B(n22638), .Z(n22636) );
  OR U31214 ( .A(n22639), .B(n22640), .Z(n22638) );
  IV U31215 ( .A(n22641), .Z(n22640) );
  NANDN U31216 ( .A(n22641), .B(n22639), .Z(n22635) );
  AND U31217 ( .A(n22642), .B(n22643), .Z(n22601) );
  NAND U31218 ( .A(n22644), .B(n22645), .Z(n22643) );
  NANDN U31219 ( .A(n22646), .B(n22647), .Z(n22645) );
  NANDN U31220 ( .A(n22647), .B(n22646), .Z(n22642) );
  IV U31221 ( .A(n22648), .Z(n22647) );
  NAND U31222 ( .A(n22649), .B(n22650), .Z(n22604) );
  NANDN U31223 ( .A(n22651), .B(n22652), .Z(n22650) );
  NANDN U31224 ( .A(n22653), .B(n22654), .Z(n22652) );
  NANDN U31225 ( .A(n22654), .B(n22653), .Z(n22649) );
  IV U31226 ( .A(n22655), .Z(n22653) );
  XOR U31227 ( .A(n22630), .B(n22656), .Z(N63375) );
  XNOR U31228 ( .A(n22633), .B(n22632), .Z(n22656) );
  XNOR U31229 ( .A(n22644), .B(n22657), .Z(n22632) );
  XNOR U31230 ( .A(n22648), .B(n22646), .Z(n22657) );
  XOR U31231 ( .A(n22654), .B(n22658), .Z(n22646) );
  XNOR U31232 ( .A(n22651), .B(n22655), .Z(n22658) );
  AND U31233 ( .A(n22659), .B(n22660), .Z(n22655) );
  NAND U31234 ( .A(n22661), .B(n22662), .Z(n22660) );
  NAND U31235 ( .A(n22663), .B(n22664), .Z(n22659) );
  AND U31236 ( .A(n22665), .B(n22666), .Z(n22651) );
  NAND U31237 ( .A(n22667), .B(n22668), .Z(n22666) );
  NAND U31238 ( .A(n22669), .B(n22670), .Z(n22665) );
  NANDN U31239 ( .A(n22671), .B(n22672), .Z(n22654) );
  ANDN U31240 ( .B(n22673), .A(n22674), .Z(n22648) );
  XNOR U31241 ( .A(n22639), .B(n22675), .Z(n22644) );
  XNOR U31242 ( .A(n22637), .B(n22641), .Z(n22675) );
  AND U31243 ( .A(n22676), .B(n22677), .Z(n22641) );
  NAND U31244 ( .A(n22678), .B(n22679), .Z(n22677) );
  NAND U31245 ( .A(n22680), .B(n22681), .Z(n22676) );
  AND U31246 ( .A(n22682), .B(n22683), .Z(n22637) );
  NAND U31247 ( .A(n22684), .B(n22685), .Z(n22683) );
  NAND U31248 ( .A(n22686), .B(n22687), .Z(n22682) );
  AND U31249 ( .A(n22688), .B(n22689), .Z(n22639) );
  NAND U31250 ( .A(n22690), .B(n22691), .Z(n22633) );
  XNOR U31251 ( .A(n22616), .B(n22692), .Z(n22630) );
  XNOR U31252 ( .A(n22620), .B(n22618), .Z(n22692) );
  XOR U31253 ( .A(n22626), .B(n22693), .Z(n22618) );
  XNOR U31254 ( .A(n22623), .B(n22627), .Z(n22693) );
  AND U31255 ( .A(n22694), .B(n22695), .Z(n22627) );
  NAND U31256 ( .A(n22696), .B(n22697), .Z(n22695) );
  NAND U31257 ( .A(n22698), .B(n22699), .Z(n22694) );
  AND U31258 ( .A(n22700), .B(n22701), .Z(n22623) );
  NAND U31259 ( .A(n22702), .B(n22703), .Z(n22701) );
  NAND U31260 ( .A(n22704), .B(n22705), .Z(n22700) );
  NANDN U31261 ( .A(n22706), .B(n22707), .Z(n22626) );
  ANDN U31262 ( .B(n22708), .A(n22709), .Z(n22620) );
  XNOR U31263 ( .A(n22611), .B(n22710), .Z(n22616) );
  XNOR U31264 ( .A(n22609), .B(n22613), .Z(n22710) );
  AND U31265 ( .A(n22711), .B(n22712), .Z(n22613) );
  NAND U31266 ( .A(n22713), .B(n22714), .Z(n22712) );
  NAND U31267 ( .A(n22715), .B(n22716), .Z(n22711) );
  AND U31268 ( .A(n22717), .B(n22718), .Z(n22609) );
  NAND U31269 ( .A(n22719), .B(n22720), .Z(n22718) );
  NAND U31270 ( .A(n22721), .B(n22722), .Z(n22717) );
  AND U31271 ( .A(n22723), .B(n22724), .Z(n22611) );
  XOR U31272 ( .A(n22691), .B(n22690), .Z(N63374) );
  XNOR U31273 ( .A(n22708), .B(n22709), .Z(n22690) );
  XNOR U31274 ( .A(n22723), .B(n22724), .Z(n22709) );
  XOR U31275 ( .A(n22720), .B(n22719), .Z(n22724) );
  XOR U31276 ( .A(y[5148]), .B(x[5148]), .Z(n22719) );
  XOR U31277 ( .A(n22722), .B(n22721), .Z(n22720) );
  XOR U31278 ( .A(y[5150]), .B(x[5150]), .Z(n22721) );
  XOR U31279 ( .A(y[5149]), .B(x[5149]), .Z(n22722) );
  XOR U31280 ( .A(n22714), .B(n22713), .Z(n22723) );
  XOR U31281 ( .A(n22716), .B(n22715), .Z(n22713) );
  XOR U31282 ( .A(y[5147]), .B(x[5147]), .Z(n22715) );
  XOR U31283 ( .A(y[5146]), .B(x[5146]), .Z(n22716) );
  XOR U31284 ( .A(y[5145]), .B(x[5145]), .Z(n22714) );
  XNOR U31285 ( .A(n22707), .B(n22706), .Z(n22708) );
  XNOR U31286 ( .A(n22703), .B(n22702), .Z(n22706) );
  XOR U31287 ( .A(n22705), .B(n22704), .Z(n22702) );
  XOR U31288 ( .A(y[5144]), .B(x[5144]), .Z(n22704) );
  XOR U31289 ( .A(y[5143]), .B(x[5143]), .Z(n22705) );
  XOR U31290 ( .A(y[5142]), .B(x[5142]), .Z(n22703) );
  XOR U31291 ( .A(n22697), .B(n22696), .Z(n22707) );
  XOR U31292 ( .A(n22699), .B(n22698), .Z(n22696) );
  XOR U31293 ( .A(y[5141]), .B(x[5141]), .Z(n22698) );
  XOR U31294 ( .A(y[5140]), .B(x[5140]), .Z(n22699) );
  XOR U31295 ( .A(y[5139]), .B(x[5139]), .Z(n22697) );
  XNOR U31296 ( .A(n22673), .B(n22674), .Z(n22691) );
  XNOR U31297 ( .A(n22688), .B(n22689), .Z(n22674) );
  XOR U31298 ( .A(n22685), .B(n22684), .Z(n22689) );
  XOR U31299 ( .A(y[5136]), .B(x[5136]), .Z(n22684) );
  XOR U31300 ( .A(n22687), .B(n22686), .Z(n22685) );
  XOR U31301 ( .A(y[5138]), .B(x[5138]), .Z(n22686) );
  XOR U31302 ( .A(y[5137]), .B(x[5137]), .Z(n22687) );
  XOR U31303 ( .A(n22679), .B(n22678), .Z(n22688) );
  XOR U31304 ( .A(n22681), .B(n22680), .Z(n22678) );
  XOR U31305 ( .A(y[5135]), .B(x[5135]), .Z(n22680) );
  XOR U31306 ( .A(y[5134]), .B(x[5134]), .Z(n22681) );
  XOR U31307 ( .A(y[5133]), .B(x[5133]), .Z(n22679) );
  XNOR U31308 ( .A(n22672), .B(n22671), .Z(n22673) );
  XNOR U31309 ( .A(n22668), .B(n22667), .Z(n22671) );
  XOR U31310 ( .A(n22670), .B(n22669), .Z(n22667) );
  XOR U31311 ( .A(y[5132]), .B(x[5132]), .Z(n22669) );
  XOR U31312 ( .A(y[5131]), .B(x[5131]), .Z(n22670) );
  XOR U31313 ( .A(y[5130]), .B(x[5130]), .Z(n22668) );
  XOR U31314 ( .A(n22662), .B(n22661), .Z(n22672) );
  XOR U31315 ( .A(n22664), .B(n22663), .Z(n22661) );
  XOR U31316 ( .A(y[5129]), .B(x[5129]), .Z(n22663) );
  XOR U31317 ( .A(y[5128]), .B(x[5128]), .Z(n22664) );
  XOR U31318 ( .A(y[5127]), .B(x[5127]), .Z(n22662) );
  NAND U31319 ( .A(n22725), .B(n22726), .Z(N63365) );
  NAND U31320 ( .A(n22727), .B(n22728), .Z(n22726) );
  NANDN U31321 ( .A(n22729), .B(n22730), .Z(n22728) );
  NANDN U31322 ( .A(n22730), .B(n22729), .Z(n22725) );
  XOR U31323 ( .A(n22729), .B(n22731), .Z(N63364) );
  XNOR U31324 ( .A(n22727), .B(n22730), .Z(n22731) );
  NAND U31325 ( .A(n22732), .B(n22733), .Z(n22730) );
  NAND U31326 ( .A(n22734), .B(n22735), .Z(n22733) );
  NANDN U31327 ( .A(n22736), .B(n22737), .Z(n22735) );
  NANDN U31328 ( .A(n22737), .B(n22736), .Z(n22732) );
  AND U31329 ( .A(n22738), .B(n22739), .Z(n22727) );
  NAND U31330 ( .A(n22740), .B(n22741), .Z(n22739) );
  NANDN U31331 ( .A(n22742), .B(n22743), .Z(n22741) );
  NANDN U31332 ( .A(n22743), .B(n22742), .Z(n22738) );
  IV U31333 ( .A(n22744), .Z(n22743) );
  AND U31334 ( .A(n22745), .B(n22746), .Z(n22729) );
  NAND U31335 ( .A(n22747), .B(n22748), .Z(n22746) );
  NANDN U31336 ( .A(n22749), .B(n22750), .Z(n22748) );
  NANDN U31337 ( .A(n22750), .B(n22749), .Z(n22745) );
  XOR U31338 ( .A(n22742), .B(n22751), .Z(N63363) );
  XNOR U31339 ( .A(n22740), .B(n22744), .Z(n22751) );
  XOR U31340 ( .A(n22737), .B(n22752), .Z(n22744) );
  XNOR U31341 ( .A(n22734), .B(n22736), .Z(n22752) );
  AND U31342 ( .A(n22753), .B(n22754), .Z(n22736) );
  NANDN U31343 ( .A(n22755), .B(n22756), .Z(n22754) );
  OR U31344 ( .A(n22757), .B(n22758), .Z(n22756) );
  IV U31345 ( .A(n22759), .Z(n22758) );
  NANDN U31346 ( .A(n22759), .B(n22757), .Z(n22753) );
  AND U31347 ( .A(n22760), .B(n22761), .Z(n22734) );
  NAND U31348 ( .A(n22762), .B(n22763), .Z(n22761) );
  NANDN U31349 ( .A(n22764), .B(n22765), .Z(n22763) );
  NANDN U31350 ( .A(n22765), .B(n22764), .Z(n22760) );
  IV U31351 ( .A(n22766), .Z(n22765) );
  NAND U31352 ( .A(n22767), .B(n22768), .Z(n22737) );
  NANDN U31353 ( .A(n22769), .B(n22770), .Z(n22768) );
  NANDN U31354 ( .A(n22771), .B(n22772), .Z(n22770) );
  NANDN U31355 ( .A(n22772), .B(n22771), .Z(n22767) );
  IV U31356 ( .A(n22773), .Z(n22771) );
  AND U31357 ( .A(n22774), .B(n22775), .Z(n22740) );
  NAND U31358 ( .A(n22776), .B(n22777), .Z(n22775) );
  NANDN U31359 ( .A(n22778), .B(n22779), .Z(n22777) );
  NANDN U31360 ( .A(n22779), .B(n22778), .Z(n22774) );
  XOR U31361 ( .A(n22750), .B(n22780), .Z(n22742) );
  XNOR U31362 ( .A(n22747), .B(n22749), .Z(n22780) );
  AND U31363 ( .A(n22781), .B(n22782), .Z(n22749) );
  NANDN U31364 ( .A(n22783), .B(n22784), .Z(n22782) );
  OR U31365 ( .A(n22785), .B(n22786), .Z(n22784) );
  IV U31366 ( .A(n22787), .Z(n22786) );
  NANDN U31367 ( .A(n22787), .B(n22785), .Z(n22781) );
  AND U31368 ( .A(n22788), .B(n22789), .Z(n22747) );
  NAND U31369 ( .A(n22790), .B(n22791), .Z(n22789) );
  NANDN U31370 ( .A(n22792), .B(n22793), .Z(n22791) );
  NANDN U31371 ( .A(n22793), .B(n22792), .Z(n22788) );
  IV U31372 ( .A(n22794), .Z(n22793) );
  NAND U31373 ( .A(n22795), .B(n22796), .Z(n22750) );
  NANDN U31374 ( .A(n22797), .B(n22798), .Z(n22796) );
  NANDN U31375 ( .A(n22799), .B(n22800), .Z(n22798) );
  NANDN U31376 ( .A(n22800), .B(n22799), .Z(n22795) );
  IV U31377 ( .A(n22801), .Z(n22799) );
  XOR U31378 ( .A(n22776), .B(n22802), .Z(N63362) );
  XNOR U31379 ( .A(n22779), .B(n22778), .Z(n22802) );
  XNOR U31380 ( .A(n22790), .B(n22803), .Z(n22778) );
  XNOR U31381 ( .A(n22794), .B(n22792), .Z(n22803) );
  XOR U31382 ( .A(n22800), .B(n22804), .Z(n22792) );
  XNOR U31383 ( .A(n22797), .B(n22801), .Z(n22804) );
  AND U31384 ( .A(n22805), .B(n22806), .Z(n22801) );
  NAND U31385 ( .A(n22807), .B(n22808), .Z(n22806) );
  NAND U31386 ( .A(n22809), .B(n22810), .Z(n22805) );
  AND U31387 ( .A(n22811), .B(n22812), .Z(n22797) );
  NAND U31388 ( .A(n22813), .B(n22814), .Z(n22812) );
  NAND U31389 ( .A(n22815), .B(n22816), .Z(n22811) );
  NANDN U31390 ( .A(n22817), .B(n22818), .Z(n22800) );
  ANDN U31391 ( .B(n22819), .A(n22820), .Z(n22794) );
  XNOR U31392 ( .A(n22785), .B(n22821), .Z(n22790) );
  XNOR U31393 ( .A(n22783), .B(n22787), .Z(n22821) );
  AND U31394 ( .A(n22822), .B(n22823), .Z(n22787) );
  NAND U31395 ( .A(n22824), .B(n22825), .Z(n22823) );
  NAND U31396 ( .A(n22826), .B(n22827), .Z(n22822) );
  AND U31397 ( .A(n22828), .B(n22829), .Z(n22783) );
  NAND U31398 ( .A(n22830), .B(n22831), .Z(n22829) );
  NAND U31399 ( .A(n22832), .B(n22833), .Z(n22828) );
  AND U31400 ( .A(n22834), .B(n22835), .Z(n22785) );
  NAND U31401 ( .A(n22836), .B(n22837), .Z(n22779) );
  XNOR U31402 ( .A(n22762), .B(n22838), .Z(n22776) );
  XNOR U31403 ( .A(n22766), .B(n22764), .Z(n22838) );
  XOR U31404 ( .A(n22772), .B(n22839), .Z(n22764) );
  XNOR U31405 ( .A(n22769), .B(n22773), .Z(n22839) );
  AND U31406 ( .A(n22840), .B(n22841), .Z(n22773) );
  NAND U31407 ( .A(n22842), .B(n22843), .Z(n22841) );
  NAND U31408 ( .A(n22844), .B(n22845), .Z(n22840) );
  AND U31409 ( .A(n22846), .B(n22847), .Z(n22769) );
  NAND U31410 ( .A(n22848), .B(n22849), .Z(n22847) );
  NAND U31411 ( .A(n22850), .B(n22851), .Z(n22846) );
  NANDN U31412 ( .A(n22852), .B(n22853), .Z(n22772) );
  ANDN U31413 ( .B(n22854), .A(n22855), .Z(n22766) );
  XNOR U31414 ( .A(n22757), .B(n22856), .Z(n22762) );
  XNOR U31415 ( .A(n22755), .B(n22759), .Z(n22856) );
  AND U31416 ( .A(n22857), .B(n22858), .Z(n22759) );
  NAND U31417 ( .A(n22859), .B(n22860), .Z(n22858) );
  NAND U31418 ( .A(n22861), .B(n22862), .Z(n22857) );
  AND U31419 ( .A(n22863), .B(n22864), .Z(n22755) );
  NAND U31420 ( .A(n22865), .B(n22866), .Z(n22864) );
  NAND U31421 ( .A(n22867), .B(n22868), .Z(n22863) );
  AND U31422 ( .A(n22869), .B(n22870), .Z(n22757) );
  XOR U31423 ( .A(n22837), .B(n22836), .Z(N63361) );
  XNOR U31424 ( .A(n22854), .B(n22855), .Z(n22836) );
  XNOR U31425 ( .A(n22869), .B(n22870), .Z(n22855) );
  XOR U31426 ( .A(n22866), .B(n22865), .Z(n22870) );
  XOR U31427 ( .A(y[5124]), .B(x[5124]), .Z(n22865) );
  XOR U31428 ( .A(n22868), .B(n22867), .Z(n22866) );
  XOR U31429 ( .A(y[5126]), .B(x[5126]), .Z(n22867) );
  XOR U31430 ( .A(y[5125]), .B(x[5125]), .Z(n22868) );
  XOR U31431 ( .A(n22860), .B(n22859), .Z(n22869) );
  XOR U31432 ( .A(n22862), .B(n22861), .Z(n22859) );
  XOR U31433 ( .A(y[5123]), .B(x[5123]), .Z(n22861) );
  XOR U31434 ( .A(y[5122]), .B(x[5122]), .Z(n22862) );
  XOR U31435 ( .A(y[5121]), .B(x[5121]), .Z(n22860) );
  XNOR U31436 ( .A(n22853), .B(n22852), .Z(n22854) );
  XNOR U31437 ( .A(n22849), .B(n22848), .Z(n22852) );
  XOR U31438 ( .A(n22851), .B(n22850), .Z(n22848) );
  XOR U31439 ( .A(y[5120]), .B(x[5120]), .Z(n22850) );
  XOR U31440 ( .A(y[5119]), .B(x[5119]), .Z(n22851) );
  XOR U31441 ( .A(y[5118]), .B(x[5118]), .Z(n22849) );
  XOR U31442 ( .A(n22843), .B(n22842), .Z(n22853) );
  XOR U31443 ( .A(n22845), .B(n22844), .Z(n22842) );
  XOR U31444 ( .A(y[5117]), .B(x[5117]), .Z(n22844) );
  XOR U31445 ( .A(y[5116]), .B(x[5116]), .Z(n22845) );
  XOR U31446 ( .A(y[5115]), .B(x[5115]), .Z(n22843) );
  XNOR U31447 ( .A(n22819), .B(n22820), .Z(n22837) );
  XNOR U31448 ( .A(n22834), .B(n22835), .Z(n22820) );
  XOR U31449 ( .A(n22831), .B(n22830), .Z(n22835) );
  XOR U31450 ( .A(y[5112]), .B(x[5112]), .Z(n22830) );
  XOR U31451 ( .A(n22833), .B(n22832), .Z(n22831) );
  XOR U31452 ( .A(y[5114]), .B(x[5114]), .Z(n22832) );
  XOR U31453 ( .A(y[5113]), .B(x[5113]), .Z(n22833) );
  XOR U31454 ( .A(n22825), .B(n22824), .Z(n22834) );
  XOR U31455 ( .A(n22827), .B(n22826), .Z(n22824) );
  XOR U31456 ( .A(y[5111]), .B(x[5111]), .Z(n22826) );
  XOR U31457 ( .A(y[5110]), .B(x[5110]), .Z(n22827) );
  XOR U31458 ( .A(y[5109]), .B(x[5109]), .Z(n22825) );
  XNOR U31459 ( .A(n22818), .B(n22817), .Z(n22819) );
  XNOR U31460 ( .A(n22814), .B(n22813), .Z(n22817) );
  XOR U31461 ( .A(n22816), .B(n22815), .Z(n22813) );
  XOR U31462 ( .A(y[5108]), .B(x[5108]), .Z(n22815) );
  XOR U31463 ( .A(y[5107]), .B(x[5107]), .Z(n22816) );
  XOR U31464 ( .A(y[5106]), .B(x[5106]), .Z(n22814) );
  XOR U31465 ( .A(n22808), .B(n22807), .Z(n22818) );
  XOR U31466 ( .A(n22810), .B(n22809), .Z(n22807) );
  XOR U31467 ( .A(y[5105]), .B(x[5105]), .Z(n22809) );
  XOR U31468 ( .A(y[5104]), .B(x[5104]), .Z(n22810) );
  XOR U31469 ( .A(y[5103]), .B(x[5103]), .Z(n22808) );
  NAND U31470 ( .A(n22871), .B(n22872), .Z(N63352) );
  NAND U31471 ( .A(n22873), .B(n22874), .Z(n22872) );
  NANDN U31472 ( .A(n22875), .B(n22876), .Z(n22874) );
  NANDN U31473 ( .A(n22876), .B(n22875), .Z(n22871) );
  XOR U31474 ( .A(n22875), .B(n22877), .Z(N63351) );
  XNOR U31475 ( .A(n22873), .B(n22876), .Z(n22877) );
  NAND U31476 ( .A(n22878), .B(n22879), .Z(n22876) );
  NAND U31477 ( .A(n22880), .B(n22881), .Z(n22879) );
  NANDN U31478 ( .A(n22882), .B(n22883), .Z(n22881) );
  NANDN U31479 ( .A(n22883), .B(n22882), .Z(n22878) );
  AND U31480 ( .A(n22884), .B(n22885), .Z(n22873) );
  NAND U31481 ( .A(n22886), .B(n22887), .Z(n22885) );
  NANDN U31482 ( .A(n22888), .B(n22889), .Z(n22887) );
  NANDN U31483 ( .A(n22889), .B(n22888), .Z(n22884) );
  IV U31484 ( .A(n22890), .Z(n22889) );
  AND U31485 ( .A(n22891), .B(n22892), .Z(n22875) );
  NAND U31486 ( .A(n22893), .B(n22894), .Z(n22892) );
  NANDN U31487 ( .A(n22895), .B(n22896), .Z(n22894) );
  NANDN U31488 ( .A(n22896), .B(n22895), .Z(n22891) );
  XOR U31489 ( .A(n22888), .B(n22897), .Z(N63350) );
  XNOR U31490 ( .A(n22886), .B(n22890), .Z(n22897) );
  XOR U31491 ( .A(n22883), .B(n22898), .Z(n22890) );
  XNOR U31492 ( .A(n22880), .B(n22882), .Z(n22898) );
  AND U31493 ( .A(n22899), .B(n22900), .Z(n22882) );
  NANDN U31494 ( .A(n22901), .B(n22902), .Z(n22900) );
  OR U31495 ( .A(n22903), .B(n22904), .Z(n22902) );
  IV U31496 ( .A(n22905), .Z(n22904) );
  NANDN U31497 ( .A(n22905), .B(n22903), .Z(n22899) );
  AND U31498 ( .A(n22906), .B(n22907), .Z(n22880) );
  NAND U31499 ( .A(n22908), .B(n22909), .Z(n22907) );
  NANDN U31500 ( .A(n22910), .B(n22911), .Z(n22909) );
  NANDN U31501 ( .A(n22911), .B(n22910), .Z(n22906) );
  IV U31502 ( .A(n22912), .Z(n22911) );
  NAND U31503 ( .A(n22913), .B(n22914), .Z(n22883) );
  NANDN U31504 ( .A(n22915), .B(n22916), .Z(n22914) );
  NANDN U31505 ( .A(n22917), .B(n22918), .Z(n22916) );
  NANDN U31506 ( .A(n22918), .B(n22917), .Z(n22913) );
  IV U31507 ( .A(n22919), .Z(n22917) );
  AND U31508 ( .A(n22920), .B(n22921), .Z(n22886) );
  NAND U31509 ( .A(n22922), .B(n22923), .Z(n22921) );
  NANDN U31510 ( .A(n22924), .B(n22925), .Z(n22923) );
  NANDN U31511 ( .A(n22925), .B(n22924), .Z(n22920) );
  XOR U31512 ( .A(n22896), .B(n22926), .Z(n22888) );
  XNOR U31513 ( .A(n22893), .B(n22895), .Z(n22926) );
  AND U31514 ( .A(n22927), .B(n22928), .Z(n22895) );
  NANDN U31515 ( .A(n22929), .B(n22930), .Z(n22928) );
  OR U31516 ( .A(n22931), .B(n22932), .Z(n22930) );
  IV U31517 ( .A(n22933), .Z(n22932) );
  NANDN U31518 ( .A(n22933), .B(n22931), .Z(n22927) );
  AND U31519 ( .A(n22934), .B(n22935), .Z(n22893) );
  NAND U31520 ( .A(n22936), .B(n22937), .Z(n22935) );
  NANDN U31521 ( .A(n22938), .B(n22939), .Z(n22937) );
  NANDN U31522 ( .A(n22939), .B(n22938), .Z(n22934) );
  IV U31523 ( .A(n22940), .Z(n22939) );
  NAND U31524 ( .A(n22941), .B(n22942), .Z(n22896) );
  NANDN U31525 ( .A(n22943), .B(n22944), .Z(n22942) );
  NANDN U31526 ( .A(n22945), .B(n22946), .Z(n22944) );
  NANDN U31527 ( .A(n22946), .B(n22945), .Z(n22941) );
  IV U31528 ( .A(n22947), .Z(n22945) );
  XOR U31529 ( .A(n22922), .B(n22948), .Z(N63349) );
  XNOR U31530 ( .A(n22925), .B(n22924), .Z(n22948) );
  XNOR U31531 ( .A(n22936), .B(n22949), .Z(n22924) );
  XNOR U31532 ( .A(n22940), .B(n22938), .Z(n22949) );
  XOR U31533 ( .A(n22946), .B(n22950), .Z(n22938) );
  XNOR U31534 ( .A(n22943), .B(n22947), .Z(n22950) );
  AND U31535 ( .A(n22951), .B(n22952), .Z(n22947) );
  NAND U31536 ( .A(n22953), .B(n22954), .Z(n22952) );
  NAND U31537 ( .A(n22955), .B(n22956), .Z(n22951) );
  AND U31538 ( .A(n22957), .B(n22958), .Z(n22943) );
  NAND U31539 ( .A(n22959), .B(n22960), .Z(n22958) );
  NAND U31540 ( .A(n22961), .B(n22962), .Z(n22957) );
  NANDN U31541 ( .A(n22963), .B(n22964), .Z(n22946) );
  ANDN U31542 ( .B(n22965), .A(n22966), .Z(n22940) );
  XNOR U31543 ( .A(n22931), .B(n22967), .Z(n22936) );
  XNOR U31544 ( .A(n22929), .B(n22933), .Z(n22967) );
  AND U31545 ( .A(n22968), .B(n22969), .Z(n22933) );
  NAND U31546 ( .A(n22970), .B(n22971), .Z(n22969) );
  NAND U31547 ( .A(n22972), .B(n22973), .Z(n22968) );
  AND U31548 ( .A(n22974), .B(n22975), .Z(n22929) );
  NAND U31549 ( .A(n22976), .B(n22977), .Z(n22975) );
  NAND U31550 ( .A(n22978), .B(n22979), .Z(n22974) );
  AND U31551 ( .A(n22980), .B(n22981), .Z(n22931) );
  NAND U31552 ( .A(n22982), .B(n22983), .Z(n22925) );
  XNOR U31553 ( .A(n22908), .B(n22984), .Z(n22922) );
  XNOR U31554 ( .A(n22912), .B(n22910), .Z(n22984) );
  XOR U31555 ( .A(n22918), .B(n22985), .Z(n22910) );
  XNOR U31556 ( .A(n22915), .B(n22919), .Z(n22985) );
  AND U31557 ( .A(n22986), .B(n22987), .Z(n22919) );
  NAND U31558 ( .A(n22988), .B(n22989), .Z(n22987) );
  NAND U31559 ( .A(n22990), .B(n22991), .Z(n22986) );
  AND U31560 ( .A(n22992), .B(n22993), .Z(n22915) );
  NAND U31561 ( .A(n22994), .B(n22995), .Z(n22993) );
  NAND U31562 ( .A(n22996), .B(n22997), .Z(n22992) );
  NANDN U31563 ( .A(n22998), .B(n22999), .Z(n22918) );
  ANDN U31564 ( .B(n23000), .A(n23001), .Z(n22912) );
  XNOR U31565 ( .A(n22903), .B(n23002), .Z(n22908) );
  XNOR U31566 ( .A(n22901), .B(n22905), .Z(n23002) );
  AND U31567 ( .A(n23003), .B(n23004), .Z(n22905) );
  NAND U31568 ( .A(n23005), .B(n23006), .Z(n23004) );
  NAND U31569 ( .A(n23007), .B(n23008), .Z(n23003) );
  AND U31570 ( .A(n23009), .B(n23010), .Z(n22901) );
  NAND U31571 ( .A(n23011), .B(n23012), .Z(n23010) );
  NAND U31572 ( .A(n23013), .B(n23014), .Z(n23009) );
  AND U31573 ( .A(n23015), .B(n23016), .Z(n22903) );
  XOR U31574 ( .A(n22983), .B(n22982), .Z(N63348) );
  XNOR U31575 ( .A(n23000), .B(n23001), .Z(n22982) );
  XNOR U31576 ( .A(n23015), .B(n23016), .Z(n23001) );
  XOR U31577 ( .A(n23012), .B(n23011), .Z(n23016) );
  XOR U31578 ( .A(y[5100]), .B(x[5100]), .Z(n23011) );
  XOR U31579 ( .A(n23014), .B(n23013), .Z(n23012) );
  XOR U31580 ( .A(y[5102]), .B(x[5102]), .Z(n23013) );
  XOR U31581 ( .A(y[5101]), .B(x[5101]), .Z(n23014) );
  XOR U31582 ( .A(n23006), .B(n23005), .Z(n23015) );
  XOR U31583 ( .A(n23008), .B(n23007), .Z(n23005) );
  XOR U31584 ( .A(y[5099]), .B(x[5099]), .Z(n23007) );
  XOR U31585 ( .A(y[5098]), .B(x[5098]), .Z(n23008) );
  XOR U31586 ( .A(y[5097]), .B(x[5097]), .Z(n23006) );
  XNOR U31587 ( .A(n22999), .B(n22998), .Z(n23000) );
  XNOR U31588 ( .A(n22995), .B(n22994), .Z(n22998) );
  XOR U31589 ( .A(n22997), .B(n22996), .Z(n22994) );
  XOR U31590 ( .A(y[5096]), .B(x[5096]), .Z(n22996) );
  XOR U31591 ( .A(y[5095]), .B(x[5095]), .Z(n22997) );
  XOR U31592 ( .A(y[5094]), .B(x[5094]), .Z(n22995) );
  XOR U31593 ( .A(n22989), .B(n22988), .Z(n22999) );
  XOR U31594 ( .A(n22991), .B(n22990), .Z(n22988) );
  XOR U31595 ( .A(y[5093]), .B(x[5093]), .Z(n22990) );
  XOR U31596 ( .A(y[5092]), .B(x[5092]), .Z(n22991) );
  XOR U31597 ( .A(y[5091]), .B(x[5091]), .Z(n22989) );
  XNOR U31598 ( .A(n22965), .B(n22966), .Z(n22983) );
  XNOR U31599 ( .A(n22980), .B(n22981), .Z(n22966) );
  XOR U31600 ( .A(n22977), .B(n22976), .Z(n22981) );
  XOR U31601 ( .A(y[5088]), .B(x[5088]), .Z(n22976) );
  XOR U31602 ( .A(n22979), .B(n22978), .Z(n22977) );
  XOR U31603 ( .A(y[5090]), .B(x[5090]), .Z(n22978) );
  XOR U31604 ( .A(y[5089]), .B(x[5089]), .Z(n22979) );
  XOR U31605 ( .A(n22971), .B(n22970), .Z(n22980) );
  XOR U31606 ( .A(n22973), .B(n22972), .Z(n22970) );
  XOR U31607 ( .A(y[5087]), .B(x[5087]), .Z(n22972) );
  XOR U31608 ( .A(y[5086]), .B(x[5086]), .Z(n22973) );
  XOR U31609 ( .A(y[5085]), .B(x[5085]), .Z(n22971) );
  XNOR U31610 ( .A(n22964), .B(n22963), .Z(n22965) );
  XNOR U31611 ( .A(n22960), .B(n22959), .Z(n22963) );
  XOR U31612 ( .A(n22962), .B(n22961), .Z(n22959) );
  XOR U31613 ( .A(y[5084]), .B(x[5084]), .Z(n22961) );
  XOR U31614 ( .A(y[5083]), .B(x[5083]), .Z(n22962) );
  XOR U31615 ( .A(y[5082]), .B(x[5082]), .Z(n22960) );
  XOR U31616 ( .A(n22954), .B(n22953), .Z(n22964) );
  XOR U31617 ( .A(n22956), .B(n22955), .Z(n22953) );
  XOR U31618 ( .A(y[5081]), .B(x[5081]), .Z(n22955) );
  XOR U31619 ( .A(y[5080]), .B(x[5080]), .Z(n22956) );
  XOR U31620 ( .A(y[5079]), .B(x[5079]), .Z(n22954) );
  NAND U31621 ( .A(n23017), .B(n23018), .Z(N63339) );
  NAND U31622 ( .A(n23019), .B(n23020), .Z(n23018) );
  NANDN U31623 ( .A(n23021), .B(n23022), .Z(n23020) );
  NANDN U31624 ( .A(n23022), .B(n23021), .Z(n23017) );
  XOR U31625 ( .A(n23021), .B(n23023), .Z(N63338) );
  XNOR U31626 ( .A(n23019), .B(n23022), .Z(n23023) );
  NAND U31627 ( .A(n23024), .B(n23025), .Z(n23022) );
  NAND U31628 ( .A(n23026), .B(n23027), .Z(n23025) );
  NANDN U31629 ( .A(n23028), .B(n23029), .Z(n23027) );
  NANDN U31630 ( .A(n23029), .B(n23028), .Z(n23024) );
  AND U31631 ( .A(n23030), .B(n23031), .Z(n23019) );
  NAND U31632 ( .A(n23032), .B(n23033), .Z(n23031) );
  NANDN U31633 ( .A(n23034), .B(n23035), .Z(n23033) );
  NANDN U31634 ( .A(n23035), .B(n23034), .Z(n23030) );
  IV U31635 ( .A(n23036), .Z(n23035) );
  AND U31636 ( .A(n23037), .B(n23038), .Z(n23021) );
  NAND U31637 ( .A(n23039), .B(n23040), .Z(n23038) );
  NANDN U31638 ( .A(n23041), .B(n23042), .Z(n23040) );
  NANDN U31639 ( .A(n23042), .B(n23041), .Z(n23037) );
  XOR U31640 ( .A(n23034), .B(n23043), .Z(N63337) );
  XNOR U31641 ( .A(n23032), .B(n23036), .Z(n23043) );
  XOR U31642 ( .A(n23029), .B(n23044), .Z(n23036) );
  XNOR U31643 ( .A(n23026), .B(n23028), .Z(n23044) );
  AND U31644 ( .A(n23045), .B(n23046), .Z(n23028) );
  NANDN U31645 ( .A(n23047), .B(n23048), .Z(n23046) );
  OR U31646 ( .A(n23049), .B(n23050), .Z(n23048) );
  IV U31647 ( .A(n23051), .Z(n23050) );
  NANDN U31648 ( .A(n23051), .B(n23049), .Z(n23045) );
  AND U31649 ( .A(n23052), .B(n23053), .Z(n23026) );
  NAND U31650 ( .A(n23054), .B(n23055), .Z(n23053) );
  NANDN U31651 ( .A(n23056), .B(n23057), .Z(n23055) );
  NANDN U31652 ( .A(n23057), .B(n23056), .Z(n23052) );
  IV U31653 ( .A(n23058), .Z(n23057) );
  NAND U31654 ( .A(n23059), .B(n23060), .Z(n23029) );
  NANDN U31655 ( .A(n23061), .B(n23062), .Z(n23060) );
  NANDN U31656 ( .A(n23063), .B(n23064), .Z(n23062) );
  NANDN U31657 ( .A(n23064), .B(n23063), .Z(n23059) );
  IV U31658 ( .A(n23065), .Z(n23063) );
  AND U31659 ( .A(n23066), .B(n23067), .Z(n23032) );
  NAND U31660 ( .A(n23068), .B(n23069), .Z(n23067) );
  NANDN U31661 ( .A(n23070), .B(n23071), .Z(n23069) );
  NANDN U31662 ( .A(n23071), .B(n23070), .Z(n23066) );
  XOR U31663 ( .A(n23042), .B(n23072), .Z(n23034) );
  XNOR U31664 ( .A(n23039), .B(n23041), .Z(n23072) );
  AND U31665 ( .A(n23073), .B(n23074), .Z(n23041) );
  NANDN U31666 ( .A(n23075), .B(n23076), .Z(n23074) );
  OR U31667 ( .A(n23077), .B(n23078), .Z(n23076) );
  IV U31668 ( .A(n23079), .Z(n23078) );
  NANDN U31669 ( .A(n23079), .B(n23077), .Z(n23073) );
  AND U31670 ( .A(n23080), .B(n23081), .Z(n23039) );
  NAND U31671 ( .A(n23082), .B(n23083), .Z(n23081) );
  NANDN U31672 ( .A(n23084), .B(n23085), .Z(n23083) );
  NANDN U31673 ( .A(n23085), .B(n23084), .Z(n23080) );
  IV U31674 ( .A(n23086), .Z(n23085) );
  NAND U31675 ( .A(n23087), .B(n23088), .Z(n23042) );
  NANDN U31676 ( .A(n23089), .B(n23090), .Z(n23088) );
  NANDN U31677 ( .A(n23091), .B(n23092), .Z(n23090) );
  NANDN U31678 ( .A(n23092), .B(n23091), .Z(n23087) );
  IV U31679 ( .A(n23093), .Z(n23091) );
  XOR U31680 ( .A(n23068), .B(n23094), .Z(N63336) );
  XNOR U31681 ( .A(n23071), .B(n23070), .Z(n23094) );
  XNOR U31682 ( .A(n23082), .B(n23095), .Z(n23070) );
  XNOR U31683 ( .A(n23086), .B(n23084), .Z(n23095) );
  XOR U31684 ( .A(n23092), .B(n23096), .Z(n23084) );
  XNOR U31685 ( .A(n23089), .B(n23093), .Z(n23096) );
  AND U31686 ( .A(n23097), .B(n23098), .Z(n23093) );
  NAND U31687 ( .A(n23099), .B(n23100), .Z(n23098) );
  NAND U31688 ( .A(n23101), .B(n23102), .Z(n23097) );
  AND U31689 ( .A(n23103), .B(n23104), .Z(n23089) );
  NAND U31690 ( .A(n23105), .B(n23106), .Z(n23104) );
  NAND U31691 ( .A(n23107), .B(n23108), .Z(n23103) );
  NANDN U31692 ( .A(n23109), .B(n23110), .Z(n23092) );
  ANDN U31693 ( .B(n23111), .A(n23112), .Z(n23086) );
  XNOR U31694 ( .A(n23077), .B(n23113), .Z(n23082) );
  XNOR U31695 ( .A(n23075), .B(n23079), .Z(n23113) );
  AND U31696 ( .A(n23114), .B(n23115), .Z(n23079) );
  NAND U31697 ( .A(n23116), .B(n23117), .Z(n23115) );
  NAND U31698 ( .A(n23118), .B(n23119), .Z(n23114) );
  AND U31699 ( .A(n23120), .B(n23121), .Z(n23075) );
  NAND U31700 ( .A(n23122), .B(n23123), .Z(n23121) );
  NAND U31701 ( .A(n23124), .B(n23125), .Z(n23120) );
  AND U31702 ( .A(n23126), .B(n23127), .Z(n23077) );
  NAND U31703 ( .A(n23128), .B(n23129), .Z(n23071) );
  XNOR U31704 ( .A(n23054), .B(n23130), .Z(n23068) );
  XNOR U31705 ( .A(n23058), .B(n23056), .Z(n23130) );
  XOR U31706 ( .A(n23064), .B(n23131), .Z(n23056) );
  XNOR U31707 ( .A(n23061), .B(n23065), .Z(n23131) );
  AND U31708 ( .A(n23132), .B(n23133), .Z(n23065) );
  NAND U31709 ( .A(n23134), .B(n23135), .Z(n23133) );
  NAND U31710 ( .A(n23136), .B(n23137), .Z(n23132) );
  AND U31711 ( .A(n23138), .B(n23139), .Z(n23061) );
  NAND U31712 ( .A(n23140), .B(n23141), .Z(n23139) );
  NAND U31713 ( .A(n23142), .B(n23143), .Z(n23138) );
  NANDN U31714 ( .A(n23144), .B(n23145), .Z(n23064) );
  ANDN U31715 ( .B(n23146), .A(n23147), .Z(n23058) );
  XNOR U31716 ( .A(n23049), .B(n23148), .Z(n23054) );
  XNOR U31717 ( .A(n23047), .B(n23051), .Z(n23148) );
  AND U31718 ( .A(n23149), .B(n23150), .Z(n23051) );
  NAND U31719 ( .A(n23151), .B(n23152), .Z(n23150) );
  NAND U31720 ( .A(n23153), .B(n23154), .Z(n23149) );
  AND U31721 ( .A(n23155), .B(n23156), .Z(n23047) );
  NAND U31722 ( .A(n23157), .B(n23158), .Z(n23156) );
  NAND U31723 ( .A(n23159), .B(n23160), .Z(n23155) );
  AND U31724 ( .A(n23161), .B(n23162), .Z(n23049) );
  XOR U31725 ( .A(n23129), .B(n23128), .Z(N63335) );
  XNOR U31726 ( .A(n23146), .B(n23147), .Z(n23128) );
  XNOR U31727 ( .A(n23161), .B(n23162), .Z(n23147) );
  XOR U31728 ( .A(n23158), .B(n23157), .Z(n23162) );
  XOR U31729 ( .A(y[5076]), .B(x[5076]), .Z(n23157) );
  XOR U31730 ( .A(n23160), .B(n23159), .Z(n23158) );
  XOR U31731 ( .A(y[5078]), .B(x[5078]), .Z(n23159) );
  XOR U31732 ( .A(y[5077]), .B(x[5077]), .Z(n23160) );
  XOR U31733 ( .A(n23152), .B(n23151), .Z(n23161) );
  XOR U31734 ( .A(n23154), .B(n23153), .Z(n23151) );
  XOR U31735 ( .A(y[5075]), .B(x[5075]), .Z(n23153) );
  XOR U31736 ( .A(y[5074]), .B(x[5074]), .Z(n23154) );
  XOR U31737 ( .A(y[5073]), .B(x[5073]), .Z(n23152) );
  XNOR U31738 ( .A(n23145), .B(n23144), .Z(n23146) );
  XNOR U31739 ( .A(n23141), .B(n23140), .Z(n23144) );
  XOR U31740 ( .A(n23143), .B(n23142), .Z(n23140) );
  XOR U31741 ( .A(y[5072]), .B(x[5072]), .Z(n23142) );
  XOR U31742 ( .A(y[5071]), .B(x[5071]), .Z(n23143) );
  XOR U31743 ( .A(y[5070]), .B(x[5070]), .Z(n23141) );
  XOR U31744 ( .A(n23135), .B(n23134), .Z(n23145) );
  XOR U31745 ( .A(n23137), .B(n23136), .Z(n23134) );
  XOR U31746 ( .A(y[5069]), .B(x[5069]), .Z(n23136) );
  XOR U31747 ( .A(y[5068]), .B(x[5068]), .Z(n23137) );
  XOR U31748 ( .A(y[5067]), .B(x[5067]), .Z(n23135) );
  XNOR U31749 ( .A(n23111), .B(n23112), .Z(n23129) );
  XNOR U31750 ( .A(n23126), .B(n23127), .Z(n23112) );
  XOR U31751 ( .A(n23123), .B(n23122), .Z(n23127) );
  XOR U31752 ( .A(y[5064]), .B(x[5064]), .Z(n23122) );
  XOR U31753 ( .A(n23125), .B(n23124), .Z(n23123) );
  XOR U31754 ( .A(y[5066]), .B(x[5066]), .Z(n23124) );
  XOR U31755 ( .A(y[5065]), .B(x[5065]), .Z(n23125) );
  XOR U31756 ( .A(n23117), .B(n23116), .Z(n23126) );
  XOR U31757 ( .A(n23119), .B(n23118), .Z(n23116) );
  XOR U31758 ( .A(y[5063]), .B(x[5063]), .Z(n23118) );
  XOR U31759 ( .A(y[5062]), .B(x[5062]), .Z(n23119) );
  XOR U31760 ( .A(y[5061]), .B(x[5061]), .Z(n23117) );
  XNOR U31761 ( .A(n23110), .B(n23109), .Z(n23111) );
  XNOR U31762 ( .A(n23106), .B(n23105), .Z(n23109) );
  XOR U31763 ( .A(n23108), .B(n23107), .Z(n23105) );
  XOR U31764 ( .A(y[5060]), .B(x[5060]), .Z(n23107) );
  XOR U31765 ( .A(y[5059]), .B(x[5059]), .Z(n23108) );
  XOR U31766 ( .A(y[5058]), .B(x[5058]), .Z(n23106) );
  XOR U31767 ( .A(n23100), .B(n23099), .Z(n23110) );
  XOR U31768 ( .A(n23102), .B(n23101), .Z(n23099) );
  XOR U31769 ( .A(y[5057]), .B(x[5057]), .Z(n23101) );
  XOR U31770 ( .A(y[5056]), .B(x[5056]), .Z(n23102) );
  XOR U31771 ( .A(y[5055]), .B(x[5055]), .Z(n23100) );
  NAND U31772 ( .A(n23163), .B(n23164), .Z(N63326) );
  NAND U31773 ( .A(n23165), .B(n23166), .Z(n23164) );
  NANDN U31774 ( .A(n23167), .B(n23168), .Z(n23166) );
  NANDN U31775 ( .A(n23168), .B(n23167), .Z(n23163) );
  XOR U31776 ( .A(n23167), .B(n23169), .Z(N63325) );
  XNOR U31777 ( .A(n23165), .B(n23168), .Z(n23169) );
  NAND U31778 ( .A(n23170), .B(n23171), .Z(n23168) );
  NAND U31779 ( .A(n23172), .B(n23173), .Z(n23171) );
  NANDN U31780 ( .A(n23174), .B(n23175), .Z(n23173) );
  NANDN U31781 ( .A(n23175), .B(n23174), .Z(n23170) );
  AND U31782 ( .A(n23176), .B(n23177), .Z(n23165) );
  NAND U31783 ( .A(n23178), .B(n23179), .Z(n23177) );
  NANDN U31784 ( .A(n23180), .B(n23181), .Z(n23179) );
  NANDN U31785 ( .A(n23181), .B(n23180), .Z(n23176) );
  IV U31786 ( .A(n23182), .Z(n23181) );
  AND U31787 ( .A(n23183), .B(n23184), .Z(n23167) );
  NAND U31788 ( .A(n23185), .B(n23186), .Z(n23184) );
  NANDN U31789 ( .A(n23187), .B(n23188), .Z(n23186) );
  NANDN U31790 ( .A(n23188), .B(n23187), .Z(n23183) );
  XOR U31791 ( .A(n23180), .B(n23189), .Z(N63324) );
  XNOR U31792 ( .A(n23178), .B(n23182), .Z(n23189) );
  XOR U31793 ( .A(n23175), .B(n23190), .Z(n23182) );
  XNOR U31794 ( .A(n23172), .B(n23174), .Z(n23190) );
  AND U31795 ( .A(n23191), .B(n23192), .Z(n23174) );
  NANDN U31796 ( .A(n23193), .B(n23194), .Z(n23192) );
  OR U31797 ( .A(n23195), .B(n23196), .Z(n23194) );
  IV U31798 ( .A(n23197), .Z(n23196) );
  NANDN U31799 ( .A(n23197), .B(n23195), .Z(n23191) );
  AND U31800 ( .A(n23198), .B(n23199), .Z(n23172) );
  NAND U31801 ( .A(n23200), .B(n23201), .Z(n23199) );
  NANDN U31802 ( .A(n23202), .B(n23203), .Z(n23201) );
  NANDN U31803 ( .A(n23203), .B(n23202), .Z(n23198) );
  IV U31804 ( .A(n23204), .Z(n23203) );
  NAND U31805 ( .A(n23205), .B(n23206), .Z(n23175) );
  NANDN U31806 ( .A(n23207), .B(n23208), .Z(n23206) );
  NANDN U31807 ( .A(n23209), .B(n23210), .Z(n23208) );
  NANDN U31808 ( .A(n23210), .B(n23209), .Z(n23205) );
  IV U31809 ( .A(n23211), .Z(n23209) );
  AND U31810 ( .A(n23212), .B(n23213), .Z(n23178) );
  NAND U31811 ( .A(n23214), .B(n23215), .Z(n23213) );
  NANDN U31812 ( .A(n23216), .B(n23217), .Z(n23215) );
  NANDN U31813 ( .A(n23217), .B(n23216), .Z(n23212) );
  XOR U31814 ( .A(n23188), .B(n23218), .Z(n23180) );
  XNOR U31815 ( .A(n23185), .B(n23187), .Z(n23218) );
  AND U31816 ( .A(n23219), .B(n23220), .Z(n23187) );
  NANDN U31817 ( .A(n23221), .B(n23222), .Z(n23220) );
  OR U31818 ( .A(n23223), .B(n23224), .Z(n23222) );
  IV U31819 ( .A(n23225), .Z(n23224) );
  NANDN U31820 ( .A(n23225), .B(n23223), .Z(n23219) );
  AND U31821 ( .A(n23226), .B(n23227), .Z(n23185) );
  NAND U31822 ( .A(n23228), .B(n23229), .Z(n23227) );
  NANDN U31823 ( .A(n23230), .B(n23231), .Z(n23229) );
  NANDN U31824 ( .A(n23231), .B(n23230), .Z(n23226) );
  IV U31825 ( .A(n23232), .Z(n23231) );
  NAND U31826 ( .A(n23233), .B(n23234), .Z(n23188) );
  NANDN U31827 ( .A(n23235), .B(n23236), .Z(n23234) );
  NANDN U31828 ( .A(n23237), .B(n23238), .Z(n23236) );
  NANDN U31829 ( .A(n23238), .B(n23237), .Z(n23233) );
  IV U31830 ( .A(n23239), .Z(n23237) );
  XOR U31831 ( .A(n23214), .B(n23240), .Z(N63323) );
  XNOR U31832 ( .A(n23217), .B(n23216), .Z(n23240) );
  XNOR U31833 ( .A(n23228), .B(n23241), .Z(n23216) );
  XNOR U31834 ( .A(n23232), .B(n23230), .Z(n23241) );
  XOR U31835 ( .A(n23238), .B(n23242), .Z(n23230) );
  XNOR U31836 ( .A(n23235), .B(n23239), .Z(n23242) );
  AND U31837 ( .A(n23243), .B(n23244), .Z(n23239) );
  NAND U31838 ( .A(n23245), .B(n23246), .Z(n23244) );
  NAND U31839 ( .A(n23247), .B(n23248), .Z(n23243) );
  AND U31840 ( .A(n23249), .B(n23250), .Z(n23235) );
  NAND U31841 ( .A(n23251), .B(n23252), .Z(n23250) );
  NAND U31842 ( .A(n23253), .B(n23254), .Z(n23249) );
  NANDN U31843 ( .A(n23255), .B(n23256), .Z(n23238) );
  ANDN U31844 ( .B(n23257), .A(n23258), .Z(n23232) );
  XNOR U31845 ( .A(n23223), .B(n23259), .Z(n23228) );
  XNOR U31846 ( .A(n23221), .B(n23225), .Z(n23259) );
  AND U31847 ( .A(n23260), .B(n23261), .Z(n23225) );
  NAND U31848 ( .A(n23262), .B(n23263), .Z(n23261) );
  NAND U31849 ( .A(n23264), .B(n23265), .Z(n23260) );
  AND U31850 ( .A(n23266), .B(n23267), .Z(n23221) );
  NAND U31851 ( .A(n23268), .B(n23269), .Z(n23267) );
  NAND U31852 ( .A(n23270), .B(n23271), .Z(n23266) );
  AND U31853 ( .A(n23272), .B(n23273), .Z(n23223) );
  NAND U31854 ( .A(n23274), .B(n23275), .Z(n23217) );
  XNOR U31855 ( .A(n23200), .B(n23276), .Z(n23214) );
  XNOR U31856 ( .A(n23204), .B(n23202), .Z(n23276) );
  XOR U31857 ( .A(n23210), .B(n23277), .Z(n23202) );
  XNOR U31858 ( .A(n23207), .B(n23211), .Z(n23277) );
  AND U31859 ( .A(n23278), .B(n23279), .Z(n23211) );
  NAND U31860 ( .A(n23280), .B(n23281), .Z(n23279) );
  NAND U31861 ( .A(n23282), .B(n23283), .Z(n23278) );
  AND U31862 ( .A(n23284), .B(n23285), .Z(n23207) );
  NAND U31863 ( .A(n23286), .B(n23287), .Z(n23285) );
  NAND U31864 ( .A(n23288), .B(n23289), .Z(n23284) );
  NANDN U31865 ( .A(n23290), .B(n23291), .Z(n23210) );
  ANDN U31866 ( .B(n23292), .A(n23293), .Z(n23204) );
  XNOR U31867 ( .A(n23195), .B(n23294), .Z(n23200) );
  XNOR U31868 ( .A(n23193), .B(n23197), .Z(n23294) );
  AND U31869 ( .A(n23295), .B(n23296), .Z(n23197) );
  NAND U31870 ( .A(n23297), .B(n23298), .Z(n23296) );
  NAND U31871 ( .A(n23299), .B(n23300), .Z(n23295) );
  AND U31872 ( .A(n23301), .B(n23302), .Z(n23193) );
  NAND U31873 ( .A(n23303), .B(n23304), .Z(n23302) );
  NAND U31874 ( .A(n23305), .B(n23306), .Z(n23301) );
  AND U31875 ( .A(n23307), .B(n23308), .Z(n23195) );
  XOR U31876 ( .A(n23275), .B(n23274), .Z(N63322) );
  XNOR U31877 ( .A(n23292), .B(n23293), .Z(n23274) );
  XNOR U31878 ( .A(n23307), .B(n23308), .Z(n23293) );
  XOR U31879 ( .A(n23304), .B(n23303), .Z(n23308) );
  XOR U31880 ( .A(y[5052]), .B(x[5052]), .Z(n23303) );
  XOR U31881 ( .A(n23306), .B(n23305), .Z(n23304) );
  XOR U31882 ( .A(y[5054]), .B(x[5054]), .Z(n23305) );
  XOR U31883 ( .A(y[5053]), .B(x[5053]), .Z(n23306) );
  XOR U31884 ( .A(n23298), .B(n23297), .Z(n23307) );
  XOR U31885 ( .A(n23300), .B(n23299), .Z(n23297) );
  XOR U31886 ( .A(y[5051]), .B(x[5051]), .Z(n23299) );
  XOR U31887 ( .A(y[5050]), .B(x[5050]), .Z(n23300) );
  XOR U31888 ( .A(y[5049]), .B(x[5049]), .Z(n23298) );
  XNOR U31889 ( .A(n23291), .B(n23290), .Z(n23292) );
  XNOR U31890 ( .A(n23287), .B(n23286), .Z(n23290) );
  XOR U31891 ( .A(n23289), .B(n23288), .Z(n23286) );
  XOR U31892 ( .A(y[5048]), .B(x[5048]), .Z(n23288) );
  XOR U31893 ( .A(y[5047]), .B(x[5047]), .Z(n23289) );
  XOR U31894 ( .A(y[5046]), .B(x[5046]), .Z(n23287) );
  XOR U31895 ( .A(n23281), .B(n23280), .Z(n23291) );
  XOR U31896 ( .A(n23283), .B(n23282), .Z(n23280) );
  XOR U31897 ( .A(y[5045]), .B(x[5045]), .Z(n23282) );
  XOR U31898 ( .A(y[5044]), .B(x[5044]), .Z(n23283) );
  XOR U31899 ( .A(y[5043]), .B(x[5043]), .Z(n23281) );
  XNOR U31900 ( .A(n23257), .B(n23258), .Z(n23275) );
  XNOR U31901 ( .A(n23272), .B(n23273), .Z(n23258) );
  XOR U31902 ( .A(n23269), .B(n23268), .Z(n23273) );
  XOR U31903 ( .A(y[5040]), .B(x[5040]), .Z(n23268) );
  XOR U31904 ( .A(n23271), .B(n23270), .Z(n23269) );
  XOR U31905 ( .A(y[5042]), .B(x[5042]), .Z(n23270) );
  XOR U31906 ( .A(y[5041]), .B(x[5041]), .Z(n23271) );
  XOR U31907 ( .A(n23263), .B(n23262), .Z(n23272) );
  XOR U31908 ( .A(n23265), .B(n23264), .Z(n23262) );
  XOR U31909 ( .A(y[5039]), .B(x[5039]), .Z(n23264) );
  XOR U31910 ( .A(y[5038]), .B(x[5038]), .Z(n23265) );
  XOR U31911 ( .A(y[5037]), .B(x[5037]), .Z(n23263) );
  XNOR U31912 ( .A(n23256), .B(n23255), .Z(n23257) );
  XNOR U31913 ( .A(n23252), .B(n23251), .Z(n23255) );
  XOR U31914 ( .A(n23254), .B(n23253), .Z(n23251) );
  XOR U31915 ( .A(y[5036]), .B(x[5036]), .Z(n23253) );
  XOR U31916 ( .A(y[5035]), .B(x[5035]), .Z(n23254) );
  XOR U31917 ( .A(y[5034]), .B(x[5034]), .Z(n23252) );
  XOR U31918 ( .A(n23246), .B(n23245), .Z(n23256) );
  XOR U31919 ( .A(n23248), .B(n23247), .Z(n23245) );
  XOR U31920 ( .A(y[5033]), .B(x[5033]), .Z(n23247) );
  XOR U31921 ( .A(y[5032]), .B(x[5032]), .Z(n23248) );
  XOR U31922 ( .A(y[5031]), .B(x[5031]), .Z(n23246) );
  NAND U31923 ( .A(n23309), .B(n23310), .Z(N63313) );
  NAND U31924 ( .A(n23311), .B(n23312), .Z(n23310) );
  NANDN U31925 ( .A(n23313), .B(n23314), .Z(n23312) );
  NANDN U31926 ( .A(n23314), .B(n23313), .Z(n23309) );
  XOR U31927 ( .A(n23313), .B(n23315), .Z(N63312) );
  XNOR U31928 ( .A(n23311), .B(n23314), .Z(n23315) );
  NAND U31929 ( .A(n23316), .B(n23317), .Z(n23314) );
  NAND U31930 ( .A(n23318), .B(n23319), .Z(n23317) );
  NANDN U31931 ( .A(n23320), .B(n23321), .Z(n23319) );
  NANDN U31932 ( .A(n23321), .B(n23320), .Z(n23316) );
  AND U31933 ( .A(n23322), .B(n23323), .Z(n23311) );
  NAND U31934 ( .A(n23324), .B(n23325), .Z(n23323) );
  NANDN U31935 ( .A(n23326), .B(n23327), .Z(n23325) );
  NANDN U31936 ( .A(n23327), .B(n23326), .Z(n23322) );
  IV U31937 ( .A(n23328), .Z(n23327) );
  AND U31938 ( .A(n23329), .B(n23330), .Z(n23313) );
  NAND U31939 ( .A(n23331), .B(n23332), .Z(n23330) );
  NANDN U31940 ( .A(n23333), .B(n23334), .Z(n23332) );
  NANDN U31941 ( .A(n23334), .B(n23333), .Z(n23329) );
  XOR U31942 ( .A(n23326), .B(n23335), .Z(N63311) );
  XNOR U31943 ( .A(n23324), .B(n23328), .Z(n23335) );
  XOR U31944 ( .A(n23321), .B(n23336), .Z(n23328) );
  XNOR U31945 ( .A(n23318), .B(n23320), .Z(n23336) );
  AND U31946 ( .A(n23337), .B(n23338), .Z(n23320) );
  NANDN U31947 ( .A(n23339), .B(n23340), .Z(n23338) );
  OR U31948 ( .A(n23341), .B(n23342), .Z(n23340) );
  IV U31949 ( .A(n23343), .Z(n23342) );
  NANDN U31950 ( .A(n23343), .B(n23341), .Z(n23337) );
  AND U31951 ( .A(n23344), .B(n23345), .Z(n23318) );
  NAND U31952 ( .A(n23346), .B(n23347), .Z(n23345) );
  NANDN U31953 ( .A(n23348), .B(n23349), .Z(n23347) );
  NANDN U31954 ( .A(n23349), .B(n23348), .Z(n23344) );
  IV U31955 ( .A(n23350), .Z(n23349) );
  NAND U31956 ( .A(n23351), .B(n23352), .Z(n23321) );
  NANDN U31957 ( .A(n23353), .B(n23354), .Z(n23352) );
  NANDN U31958 ( .A(n23355), .B(n23356), .Z(n23354) );
  NANDN U31959 ( .A(n23356), .B(n23355), .Z(n23351) );
  IV U31960 ( .A(n23357), .Z(n23355) );
  AND U31961 ( .A(n23358), .B(n23359), .Z(n23324) );
  NAND U31962 ( .A(n23360), .B(n23361), .Z(n23359) );
  NANDN U31963 ( .A(n23362), .B(n23363), .Z(n23361) );
  NANDN U31964 ( .A(n23363), .B(n23362), .Z(n23358) );
  XOR U31965 ( .A(n23334), .B(n23364), .Z(n23326) );
  XNOR U31966 ( .A(n23331), .B(n23333), .Z(n23364) );
  AND U31967 ( .A(n23365), .B(n23366), .Z(n23333) );
  NANDN U31968 ( .A(n23367), .B(n23368), .Z(n23366) );
  OR U31969 ( .A(n23369), .B(n23370), .Z(n23368) );
  IV U31970 ( .A(n23371), .Z(n23370) );
  NANDN U31971 ( .A(n23371), .B(n23369), .Z(n23365) );
  AND U31972 ( .A(n23372), .B(n23373), .Z(n23331) );
  NAND U31973 ( .A(n23374), .B(n23375), .Z(n23373) );
  NANDN U31974 ( .A(n23376), .B(n23377), .Z(n23375) );
  NANDN U31975 ( .A(n23377), .B(n23376), .Z(n23372) );
  IV U31976 ( .A(n23378), .Z(n23377) );
  NAND U31977 ( .A(n23379), .B(n23380), .Z(n23334) );
  NANDN U31978 ( .A(n23381), .B(n23382), .Z(n23380) );
  NANDN U31979 ( .A(n23383), .B(n23384), .Z(n23382) );
  NANDN U31980 ( .A(n23384), .B(n23383), .Z(n23379) );
  IV U31981 ( .A(n23385), .Z(n23383) );
  XOR U31982 ( .A(n23360), .B(n23386), .Z(N63310) );
  XNOR U31983 ( .A(n23363), .B(n23362), .Z(n23386) );
  XNOR U31984 ( .A(n23374), .B(n23387), .Z(n23362) );
  XNOR U31985 ( .A(n23378), .B(n23376), .Z(n23387) );
  XOR U31986 ( .A(n23384), .B(n23388), .Z(n23376) );
  XNOR U31987 ( .A(n23381), .B(n23385), .Z(n23388) );
  AND U31988 ( .A(n23389), .B(n23390), .Z(n23385) );
  NAND U31989 ( .A(n23391), .B(n23392), .Z(n23390) );
  NAND U31990 ( .A(n23393), .B(n23394), .Z(n23389) );
  AND U31991 ( .A(n23395), .B(n23396), .Z(n23381) );
  NAND U31992 ( .A(n23397), .B(n23398), .Z(n23396) );
  NAND U31993 ( .A(n23399), .B(n23400), .Z(n23395) );
  NANDN U31994 ( .A(n23401), .B(n23402), .Z(n23384) );
  ANDN U31995 ( .B(n23403), .A(n23404), .Z(n23378) );
  XNOR U31996 ( .A(n23369), .B(n23405), .Z(n23374) );
  XNOR U31997 ( .A(n23367), .B(n23371), .Z(n23405) );
  AND U31998 ( .A(n23406), .B(n23407), .Z(n23371) );
  NAND U31999 ( .A(n23408), .B(n23409), .Z(n23407) );
  NAND U32000 ( .A(n23410), .B(n23411), .Z(n23406) );
  AND U32001 ( .A(n23412), .B(n23413), .Z(n23367) );
  NAND U32002 ( .A(n23414), .B(n23415), .Z(n23413) );
  NAND U32003 ( .A(n23416), .B(n23417), .Z(n23412) );
  AND U32004 ( .A(n23418), .B(n23419), .Z(n23369) );
  NAND U32005 ( .A(n23420), .B(n23421), .Z(n23363) );
  XNOR U32006 ( .A(n23346), .B(n23422), .Z(n23360) );
  XNOR U32007 ( .A(n23350), .B(n23348), .Z(n23422) );
  XOR U32008 ( .A(n23356), .B(n23423), .Z(n23348) );
  XNOR U32009 ( .A(n23353), .B(n23357), .Z(n23423) );
  AND U32010 ( .A(n23424), .B(n23425), .Z(n23357) );
  NAND U32011 ( .A(n23426), .B(n23427), .Z(n23425) );
  NAND U32012 ( .A(n23428), .B(n23429), .Z(n23424) );
  AND U32013 ( .A(n23430), .B(n23431), .Z(n23353) );
  NAND U32014 ( .A(n23432), .B(n23433), .Z(n23431) );
  NAND U32015 ( .A(n23434), .B(n23435), .Z(n23430) );
  NANDN U32016 ( .A(n23436), .B(n23437), .Z(n23356) );
  ANDN U32017 ( .B(n23438), .A(n23439), .Z(n23350) );
  XNOR U32018 ( .A(n23341), .B(n23440), .Z(n23346) );
  XNOR U32019 ( .A(n23339), .B(n23343), .Z(n23440) );
  AND U32020 ( .A(n23441), .B(n23442), .Z(n23343) );
  NAND U32021 ( .A(n23443), .B(n23444), .Z(n23442) );
  NAND U32022 ( .A(n23445), .B(n23446), .Z(n23441) );
  AND U32023 ( .A(n23447), .B(n23448), .Z(n23339) );
  NAND U32024 ( .A(n23449), .B(n23450), .Z(n23448) );
  NAND U32025 ( .A(n23451), .B(n23452), .Z(n23447) );
  AND U32026 ( .A(n23453), .B(n23454), .Z(n23341) );
  XOR U32027 ( .A(n23421), .B(n23420), .Z(N63309) );
  XNOR U32028 ( .A(n23438), .B(n23439), .Z(n23420) );
  XNOR U32029 ( .A(n23453), .B(n23454), .Z(n23439) );
  XOR U32030 ( .A(n23450), .B(n23449), .Z(n23454) );
  XOR U32031 ( .A(y[5028]), .B(x[5028]), .Z(n23449) );
  XOR U32032 ( .A(n23452), .B(n23451), .Z(n23450) );
  XOR U32033 ( .A(y[5030]), .B(x[5030]), .Z(n23451) );
  XOR U32034 ( .A(y[5029]), .B(x[5029]), .Z(n23452) );
  XOR U32035 ( .A(n23444), .B(n23443), .Z(n23453) );
  XOR U32036 ( .A(n23446), .B(n23445), .Z(n23443) );
  XOR U32037 ( .A(y[5027]), .B(x[5027]), .Z(n23445) );
  XOR U32038 ( .A(y[5026]), .B(x[5026]), .Z(n23446) );
  XOR U32039 ( .A(y[5025]), .B(x[5025]), .Z(n23444) );
  XNOR U32040 ( .A(n23437), .B(n23436), .Z(n23438) );
  XNOR U32041 ( .A(n23433), .B(n23432), .Z(n23436) );
  XOR U32042 ( .A(n23435), .B(n23434), .Z(n23432) );
  XOR U32043 ( .A(y[5024]), .B(x[5024]), .Z(n23434) );
  XOR U32044 ( .A(y[5023]), .B(x[5023]), .Z(n23435) );
  XOR U32045 ( .A(y[5022]), .B(x[5022]), .Z(n23433) );
  XOR U32046 ( .A(n23427), .B(n23426), .Z(n23437) );
  XOR U32047 ( .A(n23429), .B(n23428), .Z(n23426) );
  XOR U32048 ( .A(y[5021]), .B(x[5021]), .Z(n23428) );
  XOR U32049 ( .A(y[5020]), .B(x[5020]), .Z(n23429) );
  XOR U32050 ( .A(y[5019]), .B(x[5019]), .Z(n23427) );
  XNOR U32051 ( .A(n23403), .B(n23404), .Z(n23421) );
  XNOR U32052 ( .A(n23418), .B(n23419), .Z(n23404) );
  XOR U32053 ( .A(n23415), .B(n23414), .Z(n23419) );
  XOR U32054 ( .A(y[5016]), .B(x[5016]), .Z(n23414) );
  XOR U32055 ( .A(n23417), .B(n23416), .Z(n23415) );
  XOR U32056 ( .A(y[5018]), .B(x[5018]), .Z(n23416) );
  XOR U32057 ( .A(y[5017]), .B(x[5017]), .Z(n23417) );
  XOR U32058 ( .A(n23409), .B(n23408), .Z(n23418) );
  XOR U32059 ( .A(n23411), .B(n23410), .Z(n23408) );
  XOR U32060 ( .A(y[5015]), .B(x[5015]), .Z(n23410) );
  XOR U32061 ( .A(y[5014]), .B(x[5014]), .Z(n23411) );
  XOR U32062 ( .A(y[5013]), .B(x[5013]), .Z(n23409) );
  XNOR U32063 ( .A(n23402), .B(n23401), .Z(n23403) );
  XNOR U32064 ( .A(n23398), .B(n23397), .Z(n23401) );
  XOR U32065 ( .A(n23400), .B(n23399), .Z(n23397) );
  XOR U32066 ( .A(y[5012]), .B(x[5012]), .Z(n23399) );
  XOR U32067 ( .A(y[5011]), .B(x[5011]), .Z(n23400) );
  XOR U32068 ( .A(y[5010]), .B(x[5010]), .Z(n23398) );
  XOR U32069 ( .A(n23392), .B(n23391), .Z(n23402) );
  XOR U32070 ( .A(n23394), .B(n23393), .Z(n23391) );
  XOR U32071 ( .A(y[5009]), .B(x[5009]), .Z(n23393) );
  XOR U32072 ( .A(y[5008]), .B(x[5008]), .Z(n23394) );
  XOR U32073 ( .A(y[5007]), .B(x[5007]), .Z(n23392) );
  NAND U32074 ( .A(n23455), .B(n23456), .Z(N63300) );
  NAND U32075 ( .A(n23457), .B(n23458), .Z(n23456) );
  NANDN U32076 ( .A(n23459), .B(n23460), .Z(n23458) );
  NANDN U32077 ( .A(n23460), .B(n23459), .Z(n23455) );
  XOR U32078 ( .A(n23459), .B(n23461), .Z(N63299) );
  XNOR U32079 ( .A(n23457), .B(n23460), .Z(n23461) );
  NAND U32080 ( .A(n23462), .B(n23463), .Z(n23460) );
  NAND U32081 ( .A(n23464), .B(n23465), .Z(n23463) );
  NANDN U32082 ( .A(n23466), .B(n23467), .Z(n23465) );
  NANDN U32083 ( .A(n23467), .B(n23466), .Z(n23462) );
  AND U32084 ( .A(n23468), .B(n23469), .Z(n23457) );
  NAND U32085 ( .A(n23470), .B(n23471), .Z(n23469) );
  NANDN U32086 ( .A(n23472), .B(n23473), .Z(n23471) );
  NANDN U32087 ( .A(n23473), .B(n23472), .Z(n23468) );
  IV U32088 ( .A(n23474), .Z(n23473) );
  AND U32089 ( .A(n23475), .B(n23476), .Z(n23459) );
  NAND U32090 ( .A(n23477), .B(n23478), .Z(n23476) );
  NANDN U32091 ( .A(n23479), .B(n23480), .Z(n23478) );
  NANDN U32092 ( .A(n23480), .B(n23479), .Z(n23475) );
  XOR U32093 ( .A(n23472), .B(n23481), .Z(N63298) );
  XNOR U32094 ( .A(n23470), .B(n23474), .Z(n23481) );
  XOR U32095 ( .A(n23467), .B(n23482), .Z(n23474) );
  XNOR U32096 ( .A(n23464), .B(n23466), .Z(n23482) );
  AND U32097 ( .A(n23483), .B(n23484), .Z(n23466) );
  NANDN U32098 ( .A(n23485), .B(n23486), .Z(n23484) );
  OR U32099 ( .A(n23487), .B(n23488), .Z(n23486) );
  IV U32100 ( .A(n23489), .Z(n23488) );
  NANDN U32101 ( .A(n23489), .B(n23487), .Z(n23483) );
  AND U32102 ( .A(n23490), .B(n23491), .Z(n23464) );
  NAND U32103 ( .A(n23492), .B(n23493), .Z(n23491) );
  NANDN U32104 ( .A(n23494), .B(n23495), .Z(n23493) );
  NANDN U32105 ( .A(n23495), .B(n23494), .Z(n23490) );
  IV U32106 ( .A(n23496), .Z(n23495) );
  NAND U32107 ( .A(n23497), .B(n23498), .Z(n23467) );
  NANDN U32108 ( .A(n23499), .B(n23500), .Z(n23498) );
  NANDN U32109 ( .A(n23501), .B(n23502), .Z(n23500) );
  NANDN U32110 ( .A(n23502), .B(n23501), .Z(n23497) );
  IV U32111 ( .A(n23503), .Z(n23501) );
  AND U32112 ( .A(n23504), .B(n23505), .Z(n23470) );
  NAND U32113 ( .A(n23506), .B(n23507), .Z(n23505) );
  NANDN U32114 ( .A(n23508), .B(n23509), .Z(n23507) );
  NANDN U32115 ( .A(n23509), .B(n23508), .Z(n23504) );
  XOR U32116 ( .A(n23480), .B(n23510), .Z(n23472) );
  XNOR U32117 ( .A(n23477), .B(n23479), .Z(n23510) );
  AND U32118 ( .A(n23511), .B(n23512), .Z(n23479) );
  NANDN U32119 ( .A(n23513), .B(n23514), .Z(n23512) );
  OR U32120 ( .A(n23515), .B(n23516), .Z(n23514) );
  IV U32121 ( .A(n23517), .Z(n23516) );
  NANDN U32122 ( .A(n23517), .B(n23515), .Z(n23511) );
  AND U32123 ( .A(n23518), .B(n23519), .Z(n23477) );
  NAND U32124 ( .A(n23520), .B(n23521), .Z(n23519) );
  NANDN U32125 ( .A(n23522), .B(n23523), .Z(n23521) );
  NANDN U32126 ( .A(n23523), .B(n23522), .Z(n23518) );
  IV U32127 ( .A(n23524), .Z(n23523) );
  NAND U32128 ( .A(n23525), .B(n23526), .Z(n23480) );
  NANDN U32129 ( .A(n23527), .B(n23528), .Z(n23526) );
  NANDN U32130 ( .A(n23529), .B(n23530), .Z(n23528) );
  NANDN U32131 ( .A(n23530), .B(n23529), .Z(n23525) );
  IV U32132 ( .A(n23531), .Z(n23529) );
  XOR U32133 ( .A(n23506), .B(n23532), .Z(N63297) );
  XNOR U32134 ( .A(n23509), .B(n23508), .Z(n23532) );
  XNOR U32135 ( .A(n23520), .B(n23533), .Z(n23508) );
  XNOR U32136 ( .A(n23524), .B(n23522), .Z(n23533) );
  XOR U32137 ( .A(n23530), .B(n23534), .Z(n23522) );
  XNOR U32138 ( .A(n23527), .B(n23531), .Z(n23534) );
  AND U32139 ( .A(n23535), .B(n23536), .Z(n23531) );
  NAND U32140 ( .A(n23537), .B(n23538), .Z(n23536) );
  NAND U32141 ( .A(n23539), .B(n23540), .Z(n23535) );
  AND U32142 ( .A(n23541), .B(n23542), .Z(n23527) );
  NAND U32143 ( .A(n23543), .B(n23544), .Z(n23542) );
  NAND U32144 ( .A(n23545), .B(n23546), .Z(n23541) );
  NANDN U32145 ( .A(n23547), .B(n23548), .Z(n23530) );
  ANDN U32146 ( .B(n23549), .A(n23550), .Z(n23524) );
  XNOR U32147 ( .A(n23515), .B(n23551), .Z(n23520) );
  XNOR U32148 ( .A(n23513), .B(n23517), .Z(n23551) );
  AND U32149 ( .A(n23552), .B(n23553), .Z(n23517) );
  NAND U32150 ( .A(n23554), .B(n23555), .Z(n23553) );
  NAND U32151 ( .A(n23556), .B(n23557), .Z(n23552) );
  AND U32152 ( .A(n23558), .B(n23559), .Z(n23513) );
  NAND U32153 ( .A(n23560), .B(n23561), .Z(n23559) );
  NAND U32154 ( .A(n23562), .B(n23563), .Z(n23558) );
  AND U32155 ( .A(n23564), .B(n23565), .Z(n23515) );
  NAND U32156 ( .A(n23566), .B(n23567), .Z(n23509) );
  XNOR U32157 ( .A(n23492), .B(n23568), .Z(n23506) );
  XNOR U32158 ( .A(n23496), .B(n23494), .Z(n23568) );
  XOR U32159 ( .A(n23502), .B(n23569), .Z(n23494) );
  XNOR U32160 ( .A(n23499), .B(n23503), .Z(n23569) );
  AND U32161 ( .A(n23570), .B(n23571), .Z(n23503) );
  NAND U32162 ( .A(n23572), .B(n23573), .Z(n23571) );
  NAND U32163 ( .A(n23574), .B(n23575), .Z(n23570) );
  AND U32164 ( .A(n23576), .B(n23577), .Z(n23499) );
  NAND U32165 ( .A(n23578), .B(n23579), .Z(n23577) );
  NAND U32166 ( .A(n23580), .B(n23581), .Z(n23576) );
  NANDN U32167 ( .A(n23582), .B(n23583), .Z(n23502) );
  ANDN U32168 ( .B(n23584), .A(n23585), .Z(n23496) );
  XNOR U32169 ( .A(n23487), .B(n23586), .Z(n23492) );
  XNOR U32170 ( .A(n23485), .B(n23489), .Z(n23586) );
  AND U32171 ( .A(n23587), .B(n23588), .Z(n23489) );
  NAND U32172 ( .A(n23589), .B(n23590), .Z(n23588) );
  NAND U32173 ( .A(n23591), .B(n23592), .Z(n23587) );
  AND U32174 ( .A(n23593), .B(n23594), .Z(n23485) );
  NAND U32175 ( .A(n23595), .B(n23596), .Z(n23594) );
  NAND U32176 ( .A(n23597), .B(n23598), .Z(n23593) );
  AND U32177 ( .A(n23599), .B(n23600), .Z(n23487) );
  XOR U32178 ( .A(n23567), .B(n23566), .Z(N63296) );
  XNOR U32179 ( .A(n23584), .B(n23585), .Z(n23566) );
  XNOR U32180 ( .A(n23599), .B(n23600), .Z(n23585) );
  XOR U32181 ( .A(n23596), .B(n23595), .Z(n23600) );
  XOR U32182 ( .A(y[5004]), .B(x[5004]), .Z(n23595) );
  XOR U32183 ( .A(n23598), .B(n23597), .Z(n23596) );
  XOR U32184 ( .A(y[5006]), .B(x[5006]), .Z(n23597) );
  XOR U32185 ( .A(y[5005]), .B(x[5005]), .Z(n23598) );
  XOR U32186 ( .A(n23590), .B(n23589), .Z(n23599) );
  XOR U32187 ( .A(n23592), .B(n23591), .Z(n23589) );
  XOR U32188 ( .A(y[5003]), .B(x[5003]), .Z(n23591) );
  XOR U32189 ( .A(y[5002]), .B(x[5002]), .Z(n23592) );
  XOR U32190 ( .A(y[5001]), .B(x[5001]), .Z(n23590) );
  XNOR U32191 ( .A(n23583), .B(n23582), .Z(n23584) );
  XNOR U32192 ( .A(n23579), .B(n23578), .Z(n23582) );
  XOR U32193 ( .A(n23581), .B(n23580), .Z(n23578) );
  XOR U32194 ( .A(y[5000]), .B(x[5000]), .Z(n23580) );
  XOR U32195 ( .A(y[4999]), .B(x[4999]), .Z(n23581) );
  XOR U32196 ( .A(y[4998]), .B(x[4998]), .Z(n23579) );
  XOR U32197 ( .A(n23573), .B(n23572), .Z(n23583) );
  XOR U32198 ( .A(n23575), .B(n23574), .Z(n23572) );
  XOR U32199 ( .A(y[4997]), .B(x[4997]), .Z(n23574) );
  XOR U32200 ( .A(y[4996]), .B(x[4996]), .Z(n23575) );
  XOR U32201 ( .A(y[4995]), .B(x[4995]), .Z(n23573) );
  XNOR U32202 ( .A(n23549), .B(n23550), .Z(n23567) );
  XNOR U32203 ( .A(n23564), .B(n23565), .Z(n23550) );
  XOR U32204 ( .A(n23561), .B(n23560), .Z(n23565) );
  XOR U32205 ( .A(y[4992]), .B(x[4992]), .Z(n23560) );
  XOR U32206 ( .A(n23563), .B(n23562), .Z(n23561) );
  XOR U32207 ( .A(y[4994]), .B(x[4994]), .Z(n23562) );
  XOR U32208 ( .A(y[4993]), .B(x[4993]), .Z(n23563) );
  XOR U32209 ( .A(n23555), .B(n23554), .Z(n23564) );
  XOR U32210 ( .A(n23557), .B(n23556), .Z(n23554) );
  XOR U32211 ( .A(y[4991]), .B(x[4991]), .Z(n23556) );
  XOR U32212 ( .A(y[4990]), .B(x[4990]), .Z(n23557) );
  XOR U32213 ( .A(y[4989]), .B(x[4989]), .Z(n23555) );
  XNOR U32214 ( .A(n23548), .B(n23547), .Z(n23549) );
  XNOR U32215 ( .A(n23544), .B(n23543), .Z(n23547) );
  XOR U32216 ( .A(n23546), .B(n23545), .Z(n23543) );
  XOR U32217 ( .A(y[4988]), .B(x[4988]), .Z(n23545) );
  XOR U32218 ( .A(y[4987]), .B(x[4987]), .Z(n23546) );
  XOR U32219 ( .A(y[4986]), .B(x[4986]), .Z(n23544) );
  XOR U32220 ( .A(n23538), .B(n23537), .Z(n23548) );
  XOR U32221 ( .A(n23540), .B(n23539), .Z(n23537) );
  XOR U32222 ( .A(y[4985]), .B(x[4985]), .Z(n23539) );
  XOR U32223 ( .A(y[4984]), .B(x[4984]), .Z(n23540) );
  XOR U32224 ( .A(y[4983]), .B(x[4983]), .Z(n23538) );
  NAND U32225 ( .A(n23601), .B(n23602), .Z(N63287) );
  NAND U32226 ( .A(n23603), .B(n23604), .Z(n23602) );
  NANDN U32227 ( .A(n23605), .B(n23606), .Z(n23604) );
  NANDN U32228 ( .A(n23606), .B(n23605), .Z(n23601) );
  XOR U32229 ( .A(n23605), .B(n23607), .Z(N63286) );
  XNOR U32230 ( .A(n23603), .B(n23606), .Z(n23607) );
  NAND U32231 ( .A(n23608), .B(n23609), .Z(n23606) );
  NAND U32232 ( .A(n23610), .B(n23611), .Z(n23609) );
  NANDN U32233 ( .A(n23612), .B(n23613), .Z(n23611) );
  NANDN U32234 ( .A(n23613), .B(n23612), .Z(n23608) );
  AND U32235 ( .A(n23614), .B(n23615), .Z(n23603) );
  NAND U32236 ( .A(n23616), .B(n23617), .Z(n23615) );
  NANDN U32237 ( .A(n23618), .B(n23619), .Z(n23617) );
  NANDN U32238 ( .A(n23619), .B(n23618), .Z(n23614) );
  IV U32239 ( .A(n23620), .Z(n23619) );
  AND U32240 ( .A(n23621), .B(n23622), .Z(n23605) );
  NAND U32241 ( .A(n23623), .B(n23624), .Z(n23622) );
  NANDN U32242 ( .A(n23625), .B(n23626), .Z(n23624) );
  NANDN U32243 ( .A(n23626), .B(n23625), .Z(n23621) );
  XOR U32244 ( .A(n23618), .B(n23627), .Z(N63285) );
  XNOR U32245 ( .A(n23616), .B(n23620), .Z(n23627) );
  XOR U32246 ( .A(n23613), .B(n23628), .Z(n23620) );
  XNOR U32247 ( .A(n23610), .B(n23612), .Z(n23628) );
  AND U32248 ( .A(n23629), .B(n23630), .Z(n23612) );
  NANDN U32249 ( .A(n23631), .B(n23632), .Z(n23630) );
  OR U32250 ( .A(n23633), .B(n23634), .Z(n23632) );
  IV U32251 ( .A(n23635), .Z(n23634) );
  NANDN U32252 ( .A(n23635), .B(n23633), .Z(n23629) );
  AND U32253 ( .A(n23636), .B(n23637), .Z(n23610) );
  NAND U32254 ( .A(n23638), .B(n23639), .Z(n23637) );
  NANDN U32255 ( .A(n23640), .B(n23641), .Z(n23639) );
  NANDN U32256 ( .A(n23641), .B(n23640), .Z(n23636) );
  IV U32257 ( .A(n23642), .Z(n23641) );
  NAND U32258 ( .A(n23643), .B(n23644), .Z(n23613) );
  NANDN U32259 ( .A(n23645), .B(n23646), .Z(n23644) );
  NANDN U32260 ( .A(n23647), .B(n23648), .Z(n23646) );
  NANDN U32261 ( .A(n23648), .B(n23647), .Z(n23643) );
  IV U32262 ( .A(n23649), .Z(n23647) );
  AND U32263 ( .A(n23650), .B(n23651), .Z(n23616) );
  NAND U32264 ( .A(n23652), .B(n23653), .Z(n23651) );
  NANDN U32265 ( .A(n23654), .B(n23655), .Z(n23653) );
  NANDN U32266 ( .A(n23655), .B(n23654), .Z(n23650) );
  XOR U32267 ( .A(n23626), .B(n23656), .Z(n23618) );
  XNOR U32268 ( .A(n23623), .B(n23625), .Z(n23656) );
  AND U32269 ( .A(n23657), .B(n23658), .Z(n23625) );
  NANDN U32270 ( .A(n23659), .B(n23660), .Z(n23658) );
  OR U32271 ( .A(n23661), .B(n23662), .Z(n23660) );
  IV U32272 ( .A(n23663), .Z(n23662) );
  NANDN U32273 ( .A(n23663), .B(n23661), .Z(n23657) );
  AND U32274 ( .A(n23664), .B(n23665), .Z(n23623) );
  NAND U32275 ( .A(n23666), .B(n23667), .Z(n23665) );
  NANDN U32276 ( .A(n23668), .B(n23669), .Z(n23667) );
  NANDN U32277 ( .A(n23669), .B(n23668), .Z(n23664) );
  IV U32278 ( .A(n23670), .Z(n23669) );
  NAND U32279 ( .A(n23671), .B(n23672), .Z(n23626) );
  NANDN U32280 ( .A(n23673), .B(n23674), .Z(n23672) );
  NANDN U32281 ( .A(n23675), .B(n23676), .Z(n23674) );
  NANDN U32282 ( .A(n23676), .B(n23675), .Z(n23671) );
  IV U32283 ( .A(n23677), .Z(n23675) );
  XOR U32284 ( .A(n23652), .B(n23678), .Z(N63284) );
  XNOR U32285 ( .A(n23655), .B(n23654), .Z(n23678) );
  XNOR U32286 ( .A(n23666), .B(n23679), .Z(n23654) );
  XNOR U32287 ( .A(n23670), .B(n23668), .Z(n23679) );
  XOR U32288 ( .A(n23676), .B(n23680), .Z(n23668) );
  XNOR U32289 ( .A(n23673), .B(n23677), .Z(n23680) );
  AND U32290 ( .A(n23681), .B(n23682), .Z(n23677) );
  NAND U32291 ( .A(n23683), .B(n23684), .Z(n23682) );
  NAND U32292 ( .A(n23685), .B(n23686), .Z(n23681) );
  AND U32293 ( .A(n23687), .B(n23688), .Z(n23673) );
  NAND U32294 ( .A(n23689), .B(n23690), .Z(n23688) );
  NAND U32295 ( .A(n23691), .B(n23692), .Z(n23687) );
  NANDN U32296 ( .A(n23693), .B(n23694), .Z(n23676) );
  ANDN U32297 ( .B(n23695), .A(n23696), .Z(n23670) );
  XNOR U32298 ( .A(n23661), .B(n23697), .Z(n23666) );
  XNOR U32299 ( .A(n23659), .B(n23663), .Z(n23697) );
  AND U32300 ( .A(n23698), .B(n23699), .Z(n23663) );
  NAND U32301 ( .A(n23700), .B(n23701), .Z(n23699) );
  NAND U32302 ( .A(n23702), .B(n23703), .Z(n23698) );
  AND U32303 ( .A(n23704), .B(n23705), .Z(n23659) );
  NAND U32304 ( .A(n23706), .B(n23707), .Z(n23705) );
  NAND U32305 ( .A(n23708), .B(n23709), .Z(n23704) );
  AND U32306 ( .A(n23710), .B(n23711), .Z(n23661) );
  NAND U32307 ( .A(n23712), .B(n23713), .Z(n23655) );
  XNOR U32308 ( .A(n23638), .B(n23714), .Z(n23652) );
  XNOR U32309 ( .A(n23642), .B(n23640), .Z(n23714) );
  XOR U32310 ( .A(n23648), .B(n23715), .Z(n23640) );
  XNOR U32311 ( .A(n23645), .B(n23649), .Z(n23715) );
  AND U32312 ( .A(n23716), .B(n23717), .Z(n23649) );
  NAND U32313 ( .A(n23718), .B(n23719), .Z(n23717) );
  NAND U32314 ( .A(n23720), .B(n23721), .Z(n23716) );
  AND U32315 ( .A(n23722), .B(n23723), .Z(n23645) );
  NAND U32316 ( .A(n23724), .B(n23725), .Z(n23723) );
  NAND U32317 ( .A(n23726), .B(n23727), .Z(n23722) );
  NANDN U32318 ( .A(n23728), .B(n23729), .Z(n23648) );
  ANDN U32319 ( .B(n23730), .A(n23731), .Z(n23642) );
  XNOR U32320 ( .A(n23633), .B(n23732), .Z(n23638) );
  XNOR U32321 ( .A(n23631), .B(n23635), .Z(n23732) );
  AND U32322 ( .A(n23733), .B(n23734), .Z(n23635) );
  NAND U32323 ( .A(n23735), .B(n23736), .Z(n23734) );
  NAND U32324 ( .A(n23737), .B(n23738), .Z(n23733) );
  AND U32325 ( .A(n23739), .B(n23740), .Z(n23631) );
  NAND U32326 ( .A(n23741), .B(n23742), .Z(n23740) );
  NAND U32327 ( .A(n23743), .B(n23744), .Z(n23739) );
  AND U32328 ( .A(n23745), .B(n23746), .Z(n23633) );
  XOR U32329 ( .A(n23713), .B(n23712), .Z(N63283) );
  XNOR U32330 ( .A(n23730), .B(n23731), .Z(n23712) );
  XNOR U32331 ( .A(n23745), .B(n23746), .Z(n23731) );
  XOR U32332 ( .A(n23742), .B(n23741), .Z(n23746) );
  XOR U32333 ( .A(y[4980]), .B(x[4980]), .Z(n23741) );
  XOR U32334 ( .A(n23744), .B(n23743), .Z(n23742) );
  XOR U32335 ( .A(y[4982]), .B(x[4982]), .Z(n23743) );
  XOR U32336 ( .A(y[4981]), .B(x[4981]), .Z(n23744) );
  XOR U32337 ( .A(n23736), .B(n23735), .Z(n23745) );
  XOR U32338 ( .A(n23738), .B(n23737), .Z(n23735) );
  XOR U32339 ( .A(y[4979]), .B(x[4979]), .Z(n23737) );
  XOR U32340 ( .A(y[4978]), .B(x[4978]), .Z(n23738) );
  XOR U32341 ( .A(y[4977]), .B(x[4977]), .Z(n23736) );
  XNOR U32342 ( .A(n23729), .B(n23728), .Z(n23730) );
  XNOR U32343 ( .A(n23725), .B(n23724), .Z(n23728) );
  XOR U32344 ( .A(n23727), .B(n23726), .Z(n23724) );
  XOR U32345 ( .A(y[4976]), .B(x[4976]), .Z(n23726) );
  XOR U32346 ( .A(y[4975]), .B(x[4975]), .Z(n23727) );
  XOR U32347 ( .A(y[4974]), .B(x[4974]), .Z(n23725) );
  XOR U32348 ( .A(n23719), .B(n23718), .Z(n23729) );
  XOR U32349 ( .A(n23721), .B(n23720), .Z(n23718) );
  XOR U32350 ( .A(y[4973]), .B(x[4973]), .Z(n23720) );
  XOR U32351 ( .A(y[4972]), .B(x[4972]), .Z(n23721) );
  XOR U32352 ( .A(y[4971]), .B(x[4971]), .Z(n23719) );
  XNOR U32353 ( .A(n23695), .B(n23696), .Z(n23713) );
  XNOR U32354 ( .A(n23710), .B(n23711), .Z(n23696) );
  XOR U32355 ( .A(n23707), .B(n23706), .Z(n23711) );
  XOR U32356 ( .A(y[4968]), .B(x[4968]), .Z(n23706) );
  XOR U32357 ( .A(n23709), .B(n23708), .Z(n23707) );
  XOR U32358 ( .A(y[4970]), .B(x[4970]), .Z(n23708) );
  XOR U32359 ( .A(y[4969]), .B(x[4969]), .Z(n23709) );
  XOR U32360 ( .A(n23701), .B(n23700), .Z(n23710) );
  XOR U32361 ( .A(n23703), .B(n23702), .Z(n23700) );
  XOR U32362 ( .A(y[4967]), .B(x[4967]), .Z(n23702) );
  XOR U32363 ( .A(y[4966]), .B(x[4966]), .Z(n23703) );
  XOR U32364 ( .A(y[4965]), .B(x[4965]), .Z(n23701) );
  XNOR U32365 ( .A(n23694), .B(n23693), .Z(n23695) );
  XNOR U32366 ( .A(n23690), .B(n23689), .Z(n23693) );
  XOR U32367 ( .A(n23692), .B(n23691), .Z(n23689) );
  XOR U32368 ( .A(y[4964]), .B(x[4964]), .Z(n23691) );
  XOR U32369 ( .A(y[4963]), .B(x[4963]), .Z(n23692) );
  XOR U32370 ( .A(y[4962]), .B(x[4962]), .Z(n23690) );
  XOR U32371 ( .A(n23684), .B(n23683), .Z(n23694) );
  XOR U32372 ( .A(n23686), .B(n23685), .Z(n23683) );
  XOR U32373 ( .A(y[4961]), .B(x[4961]), .Z(n23685) );
  XOR U32374 ( .A(y[4960]), .B(x[4960]), .Z(n23686) );
  XOR U32375 ( .A(y[4959]), .B(x[4959]), .Z(n23684) );
  NAND U32376 ( .A(n23747), .B(n23748), .Z(N63274) );
  NAND U32377 ( .A(n23749), .B(n23750), .Z(n23748) );
  NANDN U32378 ( .A(n23751), .B(n23752), .Z(n23750) );
  NANDN U32379 ( .A(n23752), .B(n23751), .Z(n23747) );
  XOR U32380 ( .A(n23751), .B(n23753), .Z(N63273) );
  XNOR U32381 ( .A(n23749), .B(n23752), .Z(n23753) );
  NAND U32382 ( .A(n23754), .B(n23755), .Z(n23752) );
  NAND U32383 ( .A(n23756), .B(n23757), .Z(n23755) );
  NANDN U32384 ( .A(n23758), .B(n23759), .Z(n23757) );
  NANDN U32385 ( .A(n23759), .B(n23758), .Z(n23754) );
  AND U32386 ( .A(n23760), .B(n23761), .Z(n23749) );
  NAND U32387 ( .A(n23762), .B(n23763), .Z(n23761) );
  NANDN U32388 ( .A(n23764), .B(n23765), .Z(n23763) );
  NANDN U32389 ( .A(n23765), .B(n23764), .Z(n23760) );
  IV U32390 ( .A(n23766), .Z(n23765) );
  AND U32391 ( .A(n23767), .B(n23768), .Z(n23751) );
  NAND U32392 ( .A(n23769), .B(n23770), .Z(n23768) );
  NANDN U32393 ( .A(n23771), .B(n23772), .Z(n23770) );
  NANDN U32394 ( .A(n23772), .B(n23771), .Z(n23767) );
  XOR U32395 ( .A(n23764), .B(n23773), .Z(N63272) );
  XNOR U32396 ( .A(n23762), .B(n23766), .Z(n23773) );
  XOR U32397 ( .A(n23759), .B(n23774), .Z(n23766) );
  XNOR U32398 ( .A(n23756), .B(n23758), .Z(n23774) );
  AND U32399 ( .A(n23775), .B(n23776), .Z(n23758) );
  NANDN U32400 ( .A(n23777), .B(n23778), .Z(n23776) );
  OR U32401 ( .A(n23779), .B(n23780), .Z(n23778) );
  IV U32402 ( .A(n23781), .Z(n23780) );
  NANDN U32403 ( .A(n23781), .B(n23779), .Z(n23775) );
  AND U32404 ( .A(n23782), .B(n23783), .Z(n23756) );
  NAND U32405 ( .A(n23784), .B(n23785), .Z(n23783) );
  NANDN U32406 ( .A(n23786), .B(n23787), .Z(n23785) );
  NANDN U32407 ( .A(n23787), .B(n23786), .Z(n23782) );
  IV U32408 ( .A(n23788), .Z(n23787) );
  NAND U32409 ( .A(n23789), .B(n23790), .Z(n23759) );
  NANDN U32410 ( .A(n23791), .B(n23792), .Z(n23790) );
  NANDN U32411 ( .A(n23793), .B(n23794), .Z(n23792) );
  NANDN U32412 ( .A(n23794), .B(n23793), .Z(n23789) );
  IV U32413 ( .A(n23795), .Z(n23793) );
  AND U32414 ( .A(n23796), .B(n23797), .Z(n23762) );
  NAND U32415 ( .A(n23798), .B(n23799), .Z(n23797) );
  NANDN U32416 ( .A(n23800), .B(n23801), .Z(n23799) );
  NANDN U32417 ( .A(n23801), .B(n23800), .Z(n23796) );
  XOR U32418 ( .A(n23772), .B(n23802), .Z(n23764) );
  XNOR U32419 ( .A(n23769), .B(n23771), .Z(n23802) );
  AND U32420 ( .A(n23803), .B(n23804), .Z(n23771) );
  NANDN U32421 ( .A(n23805), .B(n23806), .Z(n23804) );
  OR U32422 ( .A(n23807), .B(n23808), .Z(n23806) );
  IV U32423 ( .A(n23809), .Z(n23808) );
  NANDN U32424 ( .A(n23809), .B(n23807), .Z(n23803) );
  AND U32425 ( .A(n23810), .B(n23811), .Z(n23769) );
  NAND U32426 ( .A(n23812), .B(n23813), .Z(n23811) );
  NANDN U32427 ( .A(n23814), .B(n23815), .Z(n23813) );
  NANDN U32428 ( .A(n23815), .B(n23814), .Z(n23810) );
  IV U32429 ( .A(n23816), .Z(n23815) );
  NAND U32430 ( .A(n23817), .B(n23818), .Z(n23772) );
  NANDN U32431 ( .A(n23819), .B(n23820), .Z(n23818) );
  NANDN U32432 ( .A(n23821), .B(n23822), .Z(n23820) );
  NANDN U32433 ( .A(n23822), .B(n23821), .Z(n23817) );
  IV U32434 ( .A(n23823), .Z(n23821) );
  XOR U32435 ( .A(n23798), .B(n23824), .Z(N63271) );
  XNOR U32436 ( .A(n23801), .B(n23800), .Z(n23824) );
  XNOR U32437 ( .A(n23812), .B(n23825), .Z(n23800) );
  XNOR U32438 ( .A(n23816), .B(n23814), .Z(n23825) );
  XOR U32439 ( .A(n23822), .B(n23826), .Z(n23814) );
  XNOR U32440 ( .A(n23819), .B(n23823), .Z(n23826) );
  AND U32441 ( .A(n23827), .B(n23828), .Z(n23823) );
  NAND U32442 ( .A(n23829), .B(n23830), .Z(n23828) );
  NAND U32443 ( .A(n23831), .B(n23832), .Z(n23827) );
  AND U32444 ( .A(n23833), .B(n23834), .Z(n23819) );
  NAND U32445 ( .A(n23835), .B(n23836), .Z(n23834) );
  NAND U32446 ( .A(n23837), .B(n23838), .Z(n23833) );
  NANDN U32447 ( .A(n23839), .B(n23840), .Z(n23822) );
  ANDN U32448 ( .B(n23841), .A(n23842), .Z(n23816) );
  XNOR U32449 ( .A(n23807), .B(n23843), .Z(n23812) );
  XNOR U32450 ( .A(n23805), .B(n23809), .Z(n23843) );
  AND U32451 ( .A(n23844), .B(n23845), .Z(n23809) );
  NAND U32452 ( .A(n23846), .B(n23847), .Z(n23845) );
  NAND U32453 ( .A(n23848), .B(n23849), .Z(n23844) );
  AND U32454 ( .A(n23850), .B(n23851), .Z(n23805) );
  NAND U32455 ( .A(n23852), .B(n23853), .Z(n23851) );
  NAND U32456 ( .A(n23854), .B(n23855), .Z(n23850) );
  AND U32457 ( .A(n23856), .B(n23857), .Z(n23807) );
  NAND U32458 ( .A(n23858), .B(n23859), .Z(n23801) );
  XNOR U32459 ( .A(n23784), .B(n23860), .Z(n23798) );
  XNOR U32460 ( .A(n23788), .B(n23786), .Z(n23860) );
  XOR U32461 ( .A(n23794), .B(n23861), .Z(n23786) );
  XNOR U32462 ( .A(n23791), .B(n23795), .Z(n23861) );
  AND U32463 ( .A(n23862), .B(n23863), .Z(n23795) );
  NAND U32464 ( .A(n23864), .B(n23865), .Z(n23863) );
  NAND U32465 ( .A(n23866), .B(n23867), .Z(n23862) );
  AND U32466 ( .A(n23868), .B(n23869), .Z(n23791) );
  NAND U32467 ( .A(n23870), .B(n23871), .Z(n23869) );
  NAND U32468 ( .A(n23872), .B(n23873), .Z(n23868) );
  NANDN U32469 ( .A(n23874), .B(n23875), .Z(n23794) );
  ANDN U32470 ( .B(n23876), .A(n23877), .Z(n23788) );
  XNOR U32471 ( .A(n23779), .B(n23878), .Z(n23784) );
  XNOR U32472 ( .A(n23777), .B(n23781), .Z(n23878) );
  AND U32473 ( .A(n23879), .B(n23880), .Z(n23781) );
  NAND U32474 ( .A(n23881), .B(n23882), .Z(n23880) );
  NAND U32475 ( .A(n23883), .B(n23884), .Z(n23879) );
  AND U32476 ( .A(n23885), .B(n23886), .Z(n23777) );
  NAND U32477 ( .A(n23887), .B(n23888), .Z(n23886) );
  NAND U32478 ( .A(n23889), .B(n23890), .Z(n23885) );
  AND U32479 ( .A(n23891), .B(n23892), .Z(n23779) );
  XOR U32480 ( .A(n23859), .B(n23858), .Z(N63270) );
  XNOR U32481 ( .A(n23876), .B(n23877), .Z(n23858) );
  XNOR U32482 ( .A(n23891), .B(n23892), .Z(n23877) );
  XOR U32483 ( .A(n23888), .B(n23887), .Z(n23892) );
  XOR U32484 ( .A(y[4956]), .B(x[4956]), .Z(n23887) );
  XOR U32485 ( .A(n23890), .B(n23889), .Z(n23888) );
  XOR U32486 ( .A(y[4958]), .B(x[4958]), .Z(n23889) );
  XOR U32487 ( .A(y[4957]), .B(x[4957]), .Z(n23890) );
  XOR U32488 ( .A(n23882), .B(n23881), .Z(n23891) );
  XOR U32489 ( .A(n23884), .B(n23883), .Z(n23881) );
  XOR U32490 ( .A(y[4955]), .B(x[4955]), .Z(n23883) );
  XOR U32491 ( .A(y[4954]), .B(x[4954]), .Z(n23884) );
  XOR U32492 ( .A(y[4953]), .B(x[4953]), .Z(n23882) );
  XNOR U32493 ( .A(n23875), .B(n23874), .Z(n23876) );
  XNOR U32494 ( .A(n23871), .B(n23870), .Z(n23874) );
  XOR U32495 ( .A(n23873), .B(n23872), .Z(n23870) );
  XOR U32496 ( .A(y[4952]), .B(x[4952]), .Z(n23872) );
  XOR U32497 ( .A(y[4951]), .B(x[4951]), .Z(n23873) );
  XOR U32498 ( .A(y[4950]), .B(x[4950]), .Z(n23871) );
  XOR U32499 ( .A(n23865), .B(n23864), .Z(n23875) );
  XOR U32500 ( .A(n23867), .B(n23866), .Z(n23864) );
  XOR U32501 ( .A(y[4949]), .B(x[4949]), .Z(n23866) );
  XOR U32502 ( .A(y[4948]), .B(x[4948]), .Z(n23867) );
  XOR U32503 ( .A(y[4947]), .B(x[4947]), .Z(n23865) );
  XNOR U32504 ( .A(n23841), .B(n23842), .Z(n23859) );
  XNOR U32505 ( .A(n23856), .B(n23857), .Z(n23842) );
  XOR U32506 ( .A(n23853), .B(n23852), .Z(n23857) );
  XOR U32507 ( .A(y[4944]), .B(x[4944]), .Z(n23852) );
  XOR U32508 ( .A(n23855), .B(n23854), .Z(n23853) );
  XOR U32509 ( .A(y[4946]), .B(x[4946]), .Z(n23854) );
  XOR U32510 ( .A(y[4945]), .B(x[4945]), .Z(n23855) );
  XOR U32511 ( .A(n23847), .B(n23846), .Z(n23856) );
  XOR U32512 ( .A(n23849), .B(n23848), .Z(n23846) );
  XOR U32513 ( .A(y[4943]), .B(x[4943]), .Z(n23848) );
  XOR U32514 ( .A(y[4942]), .B(x[4942]), .Z(n23849) );
  XOR U32515 ( .A(y[4941]), .B(x[4941]), .Z(n23847) );
  XNOR U32516 ( .A(n23840), .B(n23839), .Z(n23841) );
  XNOR U32517 ( .A(n23836), .B(n23835), .Z(n23839) );
  XOR U32518 ( .A(n23838), .B(n23837), .Z(n23835) );
  XOR U32519 ( .A(y[4940]), .B(x[4940]), .Z(n23837) );
  XOR U32520 ( .A(y[4939]), .B(x[4939]), .Z(n23838) );
  XOR U32521 ( .A(y[4938]), .B(x[4938]), .Z(n23836) );
  XOR U32522 ( .A(n23830), .B(n23829), .Z(n23840) );
  XOR U32523 ( .A(n23832), .B(n23831), .Z(n23829) );
  XOR U32524 ( .A(y[4937]), .B(x[4937]), .Z(n23831) );
  XOR U32525 ( .A(y[4936]), .B(x[4936]), .Z(n23832) );
  XOR U32526 ( .A(y[4935]), .B(x[4935]), .Z(n23830) );
  NAND U32527 ( .A(n23893), .B(n23894), .Z(N63261) );
  NAND U32528 ( .A(n23895), .B(n23896), .Z(n23894) );
  NANDN U32529 ( .A(n23897), .B(n23898), .Z(n23896) );
  NANDN U32530 ( .A(n23898), .B(n23897), .Z(n23893) );
  XOR U32531 ( .A(n23897), .B(n23899), .Z(N63260) );
  XNOR U32532 ( .A(n23895), .B(n23898), .Z(n23899) );
  NAND U32533 ( .A(n23900), .B(n23901), .Z(n23898) );
  NAND U32534 ( .A(n23902), .B(n23903), .Z(n23901) );
  NANDN U32535 ( .A(n23904), .B(n23905), .Z(n23903) );
  NANDN U32536 ( .A(n23905), .B(n23904), .Z(n23900) );
  AND U32537 ( .A(n23906), .B(n23907), .Z(n23895) );
  NAND U32538 ( .A(n23908), .B(n23909), .Z(n23907) );
  NANDN U32539 ( .A(n23910), .B(n23911), .Z(n23909) );
  NANDN U32540 ( .A(n23911), .B(n23910), .Z(n23906) );
  IV U32541 ( .A(n23912), .Z(n23911) );
  AND U32542 ( .A(n23913), .B(n23914), .Z(n23897) );
  NAND U32543 ( .A(n23915), .B(n23916), .Z(n23914) );
  NANDN U32544 ( .A(n23917), .B(n23918), .Z(n23916) );
  NANDN U32545 ( .A(n23918), .B(n23917), .Z(n23913) );
  XOR U32546 ( .A(n23910), .B(n23919), .Z(N63259) );
  XNOR U32547 ( .A(n23908), .B(n23912), .Z(n23919) );
  XOR U32548 ( .A(n23905), .B(n23920), .Z(n23912) );
  XNOR U32549 ( .A(n23902), .B(n23904), .Z(n23920) );
  AND U32550 ( .A(n23921), .B(n23922), .Z(n23904) );
  NANDN U32551 ( .A(n23923), .B(n23924), .Z(n23922) );
  OR U32552 ( .A(n23925), .B(n23926), .Z(n23924) );
  IV U32553 ( .A(n23927), .Z(n23926) );
  NANDN U32554 ( .A(n23927), .B(n23925), .Z(n23921) );
  AND U32555 ( .A(n23928), .B(n23929), .Z(n23902) );
  NAND U32556 ( .A(n23930), .B(n23931), .Z(n23929) );
  NANDN U32557 ( .A(n23932), .B(n23933), .Z(n23931) );
  NANDN U32558 ( .A(n23933), .B(n23932), .Z(n23928) );
  IV U32559 ( .A(n23934), .Z(n23933) );
  NAND U32560 ( .A(n23935), .B(n23936), .Z(n23905) );
  NANDN U32561 ( .A(n23937), .B(n23938), .Z(n23936) );
  NANDN U32562 ( .A(n23939), .B(n23940), .Z(n23938) );
  NANDN U32563 ( .A(n23940), .B(n23939), .Z(n23935) );
  IV U32564 ( .A(n23941), .Z(n23939) );
  AND U32565 ( .A(n23942), .B(n23943), .Z(n23908) );
  NAND U32566 ( .A(n23944), .B(n23945), .Z(n23943) );
  NANDN U32567 ( .A(n23946), .B(n23947), .Z(n23945) );
  NANDN U32568 ( .A(n23947), .B(n23946), .Z(n23942) );
  XOR U32569 ( .A(n23918), .B(n23948), .Z(n23910) );
  XNOR U32570 ( .A(n23915), .B(n23917), .Z(n23948) );
  AND U32571 ( .A(n23949), .B(n23950), .Z(n23917) );
  NANDN U32572 ( .A(n23951), .B(n23952), .Z(n23950) );
  OR U32573 ( .A(n23953), .B(n23954), .Z(n23952) );
  IV U32574 ( .A(n23955), .Z(n23954) );
  NANDN U32575 ( .A(n23955), .B(n23953), .Z(n23949) );
  AND U32576 ( .A(n23956), .B(n23957), .Z(n23915) );
  NAND U32577 ( .A(n23958), .B(n23959), .Z(n23957) );
  NANDN U32578 ( .A(n23960), .B(n23961), .Z(n23959) );
  NANDN U32579 ( .A(n23961), .B(n23960), .Z(n23956) );
  IV U32580 ( .A(n23962), .Z(n23961) );
  NAND U32581 ( .A(n23963), .B(n23964), .Z(n23918) );
  NANDN U32582 ( .A(n23965), .B(n23966), .Z(n23964) );
  NANDN U32583 ( .A(n23967), .B(n23968), .Z(n23966) );
  NANDN U32584 ( .A(n23968), .B(n23967), .Z(n23963) );
  IV U32585 ( .A(n23969), .Z(n23967) );
  XOR U32586 ( .A(n23944), .B(n23970), .Z(N63258) );
  XNOR U32587 ( .A(n23947), .B(n23946), .Z(n23970) );
  XNOR U32588 ( .A(n23958), .B(n23971), .Z(n23946) );
  XNOR U32589 ( .A(n23962), .B(n23960), .Z(n23971) );
  XOR U32590 ( .A(n23968), .B(n23972), .Z(n23960) );
  XNOR U32591 ( .A(n23965), .B(n23969), .Z(n23972) );
  AND U32592 ( .A(n23973), .B(n23974), .Z(n23969) );
  NAND U32593 ( .A(n23975), .B(n23976), .Z(n23974) );
  NAND U32594 ( .A(n23977), .B(n23978), .Z(n23973) );
  AND U32595 ( .A(n23979), .B(n23980), .Z(n23965) );
  NAND U32596 ( .A(n23981), .B(n23982), .Z(n23980) );
  NAND U32597 ( .A(n23983), .B(n23984), .Z(n23979) );
  NANDN U32598 ( .A(n23985), .B(n23986), .Z(n23968) );
  ANDN U32599 ( .B(n23987), .A(n23988), .Z(n23962) );
  XNOR U32600 ( .A(n23953), .B(n23989), .Z(n23958) );
  XNOR U32601 ( .A(n23951), .B(n23955), .Z(n23989) );
  AND U32602 ( .A(n23990), .B(n23991), .Z(n23955) );
  NAND U32603 ( .A(n23992), .B(n23993), .Z(n23991) );
  NAND U32604 ( .A(n23994), .B(n23995), .Z(n23990) );
  AND U32605 ( .A(n23996), .B(n23997), .Z(n23951) );
  NAND U32606 ( .A(n23998), .B(n23999), .Z(n23997) );
  NAND U32607 ( .A(n24000), .B(n24001), .Z(n23996) );
  AND U32608 ( .A(n24002), .B(n24003), .Z(n23953) );
  NAND U32609 ( .A(n24004), .B(n24005), .Z(n23947) );
  XNOR U32610 ( .A(n23930), .B(n24006), .Z(n23944) );
  XNOR U32611 ( .A(n23934), .B(n23932), .Z(n24006) );
  XOR U32612 ( .A(n23940), .B(n24007), .Z(n23932) );
  XNOR U32613 ( .A(n23937), .B(n23941), .Z(n24007) );
  AND U32614 ( .A(n24008), .B(n24009), .Z(n23941) );
  NAND U32615 ( .A(n24010), .B(n24011), .Z(n24009) );
  NAND U32616 ( .A(n24012), .B(n24013), .Z(n24008) );
  AND U32617 ( .A(n24014), .B(n24015), .Z(n23937) );
  NAND U32618 ( .A(n24016), .B(n24017), .Z(n24015) );
  NAND U32619 ( .A(n24018), .B(n24019), .Z(n24014) );
  NANDN U32620 ( .A(n24020), .B(n24021), .Z(n23940) );
  ANDN U32621 ( .B(n24022), .A(n24023), .Z(n23934) );
  XNOR U32622 ( .A(n23925), .B(n24024), .Z(n23930) );
  XNOR U32623 ( .A(n23923), .B(n23927), .Z(n24024) );
  AND U32624 ( .A(n24025), .B(n24026), .Z(n23927) );
  NAND U32625 ( .A(n24027), .B(n24028), .Z(n24026) );
  NAND U32626 ( .A(n24029), .B(n24030), .Z(n24025) );
  AND U32627 ( .A(n24031), .B(n24032), .Z(n23923) );
  NAND U32628 ( .A(n24033), .B(n24034), .Z(n24032) );
  NAND U32629 ( .A(n24035), .B(n24036), .Z(n24031) );
  AND U32630 ( .A(n24037), .B(n24038), .Z(n23925) );
  XOR U32631 ( .A(n24005), .B(n24004), .Z(N63257) );
  XNOR U32632 ( .A(n24022), .B(n24023), .Z(n24004) );
  XNOR U32633 ( .A(n24037), .B(n24038), .Z(n24023) );
  XOR U32634 ( .A(n24034), .B(n24033), .Z(n24038) );
  XOR U32635 ( .A(y[4932]), .B(x[4932]), .Z(n24033) );
  XOR U32636 ( .A(n24036), .B(n24035), .Z(n24034) );
  XOR U32637 ( .A(y[4934]), .B(x[4934]), .Z(n24035) );
  XOR U32638 ( .A(y[4933]), .B(x[4933]), .Z(n24036) );
  XOR U32639 ( .A(n24028), .B(n24027), .Z(n24037) );
  XOR U32640 ( .A(n24030), .B(n24029), .Z(n24027) );
  XOR U32641 ( .A(y[4931]), .B(x[4931]), .Z(n24029) );
  XOR U32642 ( .A(y[4930]), .B(x[4930]), .Z(n24030) );
  XOR U32643 ( .A(y[4929]), .B(x[4929]), .Z(n24028) );
  XNOR U32644 ( .A(n24021), .B(n24020), .Z(n24022) );
  XNOR U32645 ( .A(n24017), .B(n24016), .Z(n24020) );
  XOR U32646 ( .A(n24019), .B(n24018), .Z(n24016) );
  XOR U32647 ( .A(y[4928]), .B(x[4928]), .Z(n24018) );
  XOR U32648 ( .A(y[4927]), .B(x[4927]), .Z(n24019) );
  XOR U32649 ( .A(y[4926]), .B(x[4926]), .Z(n24017) );
  XOR U32650 ( .A(n24011), .B(n24010), .Z(n24021) );
  XOR U32651 ( .A(n24013), .B(n24012), .Z(n24010) );
  XOR U32652 ( .A(y[4925]), .B(x[4925]), .Z(n24012) );
  XOR U32653 ( .A(y[4924]), .B(x[4924]), .Z(n24013) );
  XOR U32654 ( .A(y[4923]), .B(x[4923]), .Z(n24011) );
  XNOR U32655 ( .A(n23987), .B(n23988), .Z(n24005) );
  XNOR U32656 ( .A(n24002), .B(n24003), .Z(n23988) );
  XOR U32657 ( .A(n23999), .B(n23998), .Z(n24003) );
  XOR U32658 ( .A(y[4920]), .B(x[4920]), .Z(n23998) );
  XOR U32659 ( .A(n24001), .B(n24000), .Z(n23999) );
  XOR U32660 ( .A(y[4922]), .B(x[4922]), .Z(n24000) );
  XOR U32661 ( .A(y[4921]), .B(x[4921]), .Z(n24001) );
  XOR U32662 ( .A(n23993), .B(n23992), .Z(n24002) );
  XOR U32663 ( .A(n23995), .B(n23994), .Z(n23992) );
  XOR U32664 ( .A(y[4919]), .B(x[4919]), .Z(n23994) );
  XOR U32665 ( .A(y[4918]), .B(x[4918]), .Z(n23995) );
  XOR U32666 ( .A(y[4917]), .B(x[4917]), .Z(n23993) );
  XNOR U32667 ( .A(n23986), .B(n23985), .Z(n23987) );
  XNOR U32668 ( .A(n23982), .B(n23981), .Z(n23985) );
  XOR U32669 ( .A(n23984), .B(n23983), .Z(n23981) );
  XOR U32670 ( .A(y[4916]), .B(x[4916]), .Z(n23983) );
  XOR U32671 ( .A(y[4915]), .B(x[4915]), .Z(n23984) );
  XOR U32672 ( .A(y[4914]), .B(x[4914]), .Z(n23982) );
  XOR U32673 ( .A(n23976), .B(n23975), .Z(n23986) );
  XOR U32674 ( .A(n23978), .B(n23977), .Z(n23975) );
  XOR U32675 ( .A(y[4913]), .B(x[4913]), .Z(n23977) );
  XOR U32676 ( .A(y[4912]), .B(x[4912]), .Z(n23978) );
  XOR U32677 ( .A(y[4911]), .B(x[4911]), .Z(n23976) );
  NAND U32678 ( .A(n24039), .B(n24040), .Z(N63248) );
  NAND U32679 ( .A(n24041), .B(n24042), .Z(n24040) );
  NANDN U32680 ( .A(n24043), .B(n24044), .Z(n24042) );
  NANDN U32681 ( .A(n24044), .B(n24043), .Z(n24039) );
  XOR U32682 ( .A(n24043), .B(n24045), .Z(N63247) );
  XNOR U32683 ( .A(n24041), .B(n24044), .Z(n24045) );
  NAND U32684 ( .A(n24046), .B(n24047), .Z(n24044) );
  NAND U32685 ( .A(n24048), .B(n24049), .Z(n24047) );
  NANDN U32686 ( .A(n24050), .B(n24051), .Z(n24049) );
  NANDN U32687 ( .A(n24051), .B(n24050), .Z(n24046) );
  AND U32688 ( .A(n24052), .B(n24053), .Z(n24041) );
  NAND U32689 ( .A(n24054), .B(n24055), .Z(n24053) );
  NANDN U32690 ( .A(n24056), .B(n24057), .Z(n24055) );
  NANDN U32691 ( .A(n24057), .B(n24056), .Z(n24052) );
  IV U32692 ( .A(n24058), .Z(n24057) );
  AND U32693 ( .A(n24059), .B(n24060), .Z(n24043) );
  NAND U32694 ( .A(n24061), .B(n24062), .Z(n24060) );
  NANDN U32695 ( .A(n24063), .B(n24064), .Z(n24062) );
  NANDN U32696 ( .A(n24064), .B(n24063), .Z(n24059) );
  XOR U32697 ( .A(n24056), .B(n24065), .Z(N63246) );
  XNOR U32698 ( .A(n24054), .B(n24058), .Z(n24065) );
  XOR U32699 ( .A(n24051), .B(n24066), .Z(n24058) );
  XNOR U32700 ( .A(n24048), .B(n24050), .Z(n24066) );
  AND U32701 ( .A(n24067), .B(n24068), .Z(n24050) );
  NANDN U32702 ( .A(n24069), .B(n24070), .Z(n24068) );
  OR U32703 ( .A(n24071), .B(n24072), .Z(n24070) );
  IV U32704 ( .A(n24073), .Z(n24072) );
  NANDN U32705 ( .A(n24073), .B(n24071), .Z(n24067) );
  AND U32706 ( .A(n24074), .B(n24075), .Z(n24048) );
  NAND U32707 ( .A(n24076), .B(n24077), .Z(n24075) );
  NANDN U32708 ( .A(n24078), .B(n24079), .Z(n24077) );
  NANDN U32709 ( .A(n24079), .B(n24078), .Z(n24074) );
  IV U32710 ( .A(n24080), .Z(n24079) );
  NAND U32711 ( .A(n24081), .B(n24082), .Z(n24051) );
  NANDN U32712 ( .A(n24083), .B(n24084), .Z(n24082) );
  NANDN U32713 ( .A(n24085), .B(n24086), .Z(n24084) );
  NANDN U32714 ( .A(n24086), .B(n24085), .Z(n24081) );
  IV U32715 ( .A(n24087), .Z(n24085) );
  AND U32716 ( .A(n24088), .B(n24089), .Z(n24054) );
  NAND U32717 ( .A(n24090), .B(n24091), .Z(n24089) );
  NANDN U32718 ( .A(n24092), .B(n24093), .Z(n24091) );
  NANDN U32719 ( .A(n24093), .B(n24092), .Z(n24088) );
  XOR U32720 ( .A(n24064), .B(n24094), .Z(n24056) );
  XNOR U32721 ( .A(n24061), .B(n24063), .Z(n24094) );
  AND U32722 ( .A(n24095), .B(n24096), .Z(n24063) );
  NANDN U32723 ( .A(n24097), .B(n24098), .Z(n24096) );
  OR U32724 ( .A(n24099), .B(n24100), .Z(n24098) );
  IV U32725 ( .A(n24101), .Z(n24100) );
  NANDN U32726 ( .A(n24101), .B(n24099), .Z(n24095) );
  AND U32727 ( .A(n24102), .B(n24103), .Z(n24061) );
  NAND U32728 ( .A(n24104), .B(n24105), .Z(n24103) );
  NANDN U32729 ( .A(n24106), .B(n24107), .Z(n24105) );
  NANDN U32730 ( .A(n24107), .B(n24106), .Z(n24102) );
  IV U32731 ( .A(n24108), .Z(n24107) );
  NAND U32732 ( .A(n24109), .B(n24110), .Z(n24064) );
  NANDN U32733 ( .A(n24111), .B(n24112), .Z(n24110) );
  NANDN U32734 ( .A(n24113), .B(n24114), .Z(n24112) );
  NANDN U32735 ( .A(n24114), .B(n24113), .Z(n24109) );
  IV U32736 ( .A(n24115), .Z(n24113) );
  XOR U32737 ( .A(n24090), .B(n24116), .Z(N63245) );
  XNOR U32738 ( .A(n24093), .B(n24092), .Z(n24116) );
  XNOR U32739 ( .A(n24104), .B(n24117), .Z(n24092) );
  XNOR U32740 ( .A(n24108), .B(n24106), .Z(n24117) );
  XOR U32741 ( .A(n24114), .B(n24118), .Z(n24106) );
  XNOR U32742 ( .A(n24111), .B(n24115), .Z(n24118) );
  AND U32743 ( .A(n24119), .B(n24120), .Z(n24115) );
  NAND U32744 ( .A(n24121), .B(n24122), .Z(n24120) );
  NAND U32745 ( .A(n24123), .B(n24124), .Z(n24119) );
  AND U32746 ( .A(n24125), .B(n24126), .Z(n24111) );
  NAND U32747 ( .A(n24127), .B(n24128), .Z(n24126) );
  NAND U32748 ( .A(n24129), .B(n24130), .Z(n24125) );
  NANDN U32749 ( .A(n24131), .B(n24132), .Z(n24114) );
  ANDN U32750 ( .B(n24133), .A(n24134), .Z(n24108) );
  XNOR U32751 ( .A(n24099), .B(n24135), .Z(n24104) );
  XNOR U32752 ( .A(n24097), .B(n24101), .Z(n24135) );
  AND U32753 ( .A(n24136), .B(n24137), .Z(n24101) );
  NAND U32754 ( .A(n24138), .B(n24139), .Z(n24137) );
  NAND U32755 ( .A(n24140), .B(n24141), .Z(n24136) );
  AND U32756 ( .A(n24142), .B(n24143), .Z(n24097) );
  NAND U32757 ( .A(n24144), .B(n24145), .Z(n24143) );
  NAND U32758 ( .A(n24146), .B(n24147), .Z(n24142) );
  AND U32759 ( .A(n24148), .B(n24149), .Z(n24099) );
  NAND U32760 ( .A(n24150), .B(n24151), .Z(n24093) );
  XNOR U32761 ( .A(n24076), .B(n24152), .Z(n24090) );
  XNOR U32762 ( .A(n24080), .B(n24078), .Z(n24152) );
  XOR U32763 ( .A(n24086), .B(n24153), .Z(n24078) );
  XNOR U32764 ( .A(n24083), .B(n24087), .Z(n24153) );
  AND U32765 ( .A(n24154), .B(n24155), .Z(n24087) );
  NAND U32766 ( .A(n24156), .B(n24157), .Z(n24155) );
  NAND U32767 ( .A(n24158), .B(n24159), .Z(n24154) );
  AND U32768 ( .A(n24160), .B(n24161), .Z(n24083) );
  NAND U32769 ( .A(n24162), .B(n24163), .Z(n24161) );
  NAND U32770 ( .A(n24164), .B(n24165), .Z(n24160) );
  NANDN U32771 ( .A(n24166), .B(n24167), .Z(n24086) );
  ANDN U32772 ( .B(n24168), .A(n24169), .Z(n24080) );
  XNOR U32773 ( .A(n24071), .B(n24170), .Z(n24076) );
  XNOR U32774 ( .A(n24069), .B(n24073), .Z(n24170) );
  AND U32775 ( .A(n24171), .B(n24172), .Z(n24073) );
  NAND U32776 ( .A(n24173), .B(n24174), .Z(n24172) );
  NAND U32777 ( .A(n24175), .B(n24176), .Z(n24171) );
  AND U32778 ( .A(n24177), .B(n24178), .Z(n24069) );
  NAND U32779 ( .A(n24179), .B(n24180), .Z(n24178) );
  NAND U32780 ( .A(n24181), .B(n24182), .Z(n24177) );
  AND U32781 ( .A(n24183), .B(n24184), .Z(n24071) );
  XOR U32782 ( .A(n24151), .B(n24150), .Z(N63244) );
  XNOR U32783 ( .A(n24168), .B(n24169), .Z(n24150) );
  XNOR U32784 ( .A(n24183), .B(n24184), .Z(n24169) );
  XOR U32785 ( .A(n24180), .B(n24179), .Z(n24184) );
  XOR U32786 ( .A(y[4908]), .B(x[4908]), .Z(n24179) );
  XOR U32787 ( .A(n24182), .B(n24181), .Z(n24180) );
  XOR U32788 ( .A(y[4910]), .B(x[4910]), .Z(n24181) );
  XOR U32789 ( .A(y[4909]), .B(x[4909]), .Z(n24182) );
  XOR U32790 ( .A(n24174), .B(n24173), .Z(n24183) );
  XOR U32791 ( .A(n24176), .B(n24175), .Z(n24173) );
  XOR U32792 ( .A(y[4907]), .B(x[4907]), .Z(n24175) );
  XOR U32793 ( .A(y[4906]), .B(x[4906]), .Z(n24176) );
  XOR U32794 ( .A(y[4905]), .B(x[4905]), .Z(n24174) );
  XNOR U32795 ( .A(n24167), .B(n24166), .Z(n24168) );
  XNOR U32796 ( .A(n24163), .B(n24162), .Z(n24166) );
  XOR U32797 ( .A(n24165), .B(n24164), .Z(n24162) );
  XOR U32798 ( .A(y[4904]), .B(x[4904]), .Z(n24164) );
  XOR U32799 ( .A(y[4903]), .B(x[4903]), .Z(n24165) );
  XOR U32800 ( .A(y[4902]), .B(x[4902]), .Z(n24163) );
  XOR U32801 ( .A(n24157), .B(n24156), .Z(n24167) );
  XOR U32802 ( .A(n24159), .B(n24158), .Z(n24156) );
  XOR U32803 ( .A(y[4901]), .B(x[4901]), .Z(n24158) );
  XOR U32804 ( .A(y[4900]), .B(x[4900]), .Z(n24159) );
  XOR U32805 ( .A(y[4899]), .B(x[4899]), .Z(n24157) );
  XNOR U32806 ( .A(n24133), .B(n24134), .Z(n24151) );
  XNOR U32807 ( .A(n24148), .B(n24149), .Z(n24134) );
  XOR U32808 ( .A(n24145), .B(n24144), .Z(n24149) );
  XOR U32809 ( .A(y[4896]), .B(x[4896]), .Z(n24144) );
  XOR U32810 ( .A(n24147), .B(n24146), .Z(n24145) );
  XOR U32811 ( .A(y[4898]), .B(x[4898]), .Z(n24146) );
  XOR U32812 ( .A(y[4897]), .B(x[4897]), .Z(n24147) );
  XOR U32813 ( .A(n24139), .B(n24138), .Z(n24148) );
  XOR U32814 ( .A(n24141), .B(n24140), .Z(n24138) );
  XOR U32815 ( .A(y[4895]), .B(x[4895]), .Z(n24140) );
  XOR U32816 ( .A(y[4894]), .B(x[4894]), .Z(n24141) );
  XOR U32817 ( .A(y[4893]), .B(x[4893]), .Z(n24139) );
  XNOR U32818 ( .A(n24132), .B(n24131), .Z(n24133) );
  XNOR U32819 ( .A(n24128), .B(n24127), .Z(n24131) );
  XOR U32820 ( .A(n24130), .B(n24129), .Z(n24127) );
  XOR U32821 ( .A(y[4892]), .B(x[4892]), .Z(n24129) );
  XOR U32822 ( .A(y[4891]), .B(x[4891]), .Z(n24130) );
  XOR U32823 ( .A(y[4890]), .B(x[4890]), .Z(n24128) );
  XOR U32824 ( .A(n24122), .B(n24121), .Z(n24132) );
  XOR U32825 ( .A(n24124), .B(n24123), .Z(n24121) );
  XOR U32826 ( .A(y[4889]), .B(x[4889]), .Z(n24123) );
  XOR U32827 ( .A(y[4888]), .B(x[4888]), .Z(n24124) );
  XOR U32828 ( .A(y[4887]), .B(x[4887]), .Z(n24122) );
  NAND U32829 ( .A(n24185), .B(n24186), .Z(N63235) );
  NAND U32830 ( .A(n24187), .B(n24188), .Z(n24186) );
  NANDN U32831 ( .A(n24189), .B(n24190), .Z(n24188) );
  NANDN U32832 ( .A(n24190), .B(n24189), .Z(n24185) );
  XOR U32833 ( .A(n24189), .B(n24191), .Z(N63234) );
  XNOR U32834 ( .A(n24187), .B(n24190), .Z(n24191) );
  NAND U32835 ( .A(n24192), .B(n24193), .Z(n24190) );
  NAND U32836 ( .A(n24194), .B(n24195), .Z(n24193) );
  NANDN U32837 ( .A(n24196), .B(n24197), .Z(n24195) );
  NANDN U32838 ( .A(n24197), .B(n24196), .Z(n24192) );
  AND U32839 ( .A(n24198), .B(n24199), .Z(n24187) );
  NAND U32840 ( .A(n24200), .B(n24201), .Z(n24199) );
  NANDN U32841 ( .A(n24202), .B(n24203), .Z(n24201) );
  NANDN U32842 ( .A(n24203), .B(n24202), .Z(n24198) );
  IV U32843 ( .A(n24204), .Z(n24203) );
  AND U32844 ( .A(n24205), .B(n24206), .Z(n24189) );
  NAND U32845 ( .A(n24207), .B(n24208), .Z(n24206) );
  NANDN U32846 ( .A(n24209), .B(n24210), .Z(n24208) );
  NANDN U32847 ( .A(n24210), .B(n24209), .Z(n24205) );
  XOR U32848 ( .A(n24202), .B(n24211), .Z(N63233) );
  XNOR U32849 ( .A(n24200), .B(n24204), .Z(n24211) );
  XOR U32850 ( .A(n24197), .B(n24212), .Z(n24204) );
  XNOR U32851 ( .A(n24194), .B(n24196), .Z(n24212) );
  AND U32852 ( .A(n24213), .B(n24214), .Z(n24196) );
  NANDN U32853 ( .A(n24215), .B(n24216), .Z(n24214) );
  OR U32854 ( .A(n24217), .B(n24218), .Z(n24216) );
  IV U32855 ( .A(n24219), .Z(n24218) );
  NANDN U32856 ( .A(n24219), .B(n24217), .Z(n24213) );
  AND U32857 ( .A(n24220), .B(n24221), .Z(n24194) );
  NAND U32858 ( .A(n24222), .B(n24223), .Z(n24221) );
  NANDN U32859 ( .A(n24224), .B(n24225), .Z(n24223) );
  NANDN U32860 ( .A(n24225), .B(n24224), .Z(n24220) );
  IV U32861 ( .A(n24226), .Z(n24225) );
  NAND U32862 ( .A(n24227), .B(n24228), .Z(n24197) );
  NANDN U32863 ( .A(n24229), .B(n24230), .Z(n24228) );
  NANDN U32864 ( .A(n24231), .B(n24232), .Z(n24230) );
  NANDN U32865 ( .A(n24232), .B(n24231), .Z(n24227) );
  IV U32866 ( .A(n24233), .Z(n24231) );
  AND U32867 ( .A(n24234), .B(n24235), .Z(n24200) );
  NAND U32868 ( .A(n24236), .B(n24237), .Z(n24235) );
  NANDN U32869 ( .A(n24238), .B(n24239), .Z(n24237) );
  NANDN U32870 ( .A(n24239), .B(n24238), .Z(n24234) );
  XOR U32871 ( .A(n24210), .B(n24240), .Z(n24202) );
  XNOR U32872 ( .A(n24207), .B(n24209), .Z(n24240) );
  AND U32873 ( .A(n24241), .B(n24242), .Z(n24209) );
  NANDN U32874 ( .A(n24243), .B(n24244), .Z(n24242) );
  OR U32875 ( .A(n24245), .B(n24246), .Z(n24244) );
  IV U32876 ( .A(n24247), .Z(n24246) );
  NANDN U32877 ( .A(n24247), .B(n24245), .Z(n24241) );
  AND U32878 ( .A(n24248), .B(n24249), .Z(n24207) );
  NAND U32879 ( .A(n24250), .B(n24251), .Z(n24249) );
  NANDN U32880 ( .A(n24252), .B(n24253), .Z(n24251) );
  NANDN U32881 ( .A(n24253), .B(n24252), .Z(n24248) );
  IV U32882 ( .A(n24254), .Z(n24253) );
  NAND U32883 ( .A(n24255), .B(n24256), .Z(n24210) );
  NANDN U32884 ( .A(n24257), .B(n24258), .Z(n24256) );
  NANDN U32885 ( .A(n24259), .B(n24260), .Z(n24258) );
  NANDN U32886 ( .A(n24260), .B(n24259), .Z(n24255) );
  IV U32887 ( .A(n24261), .Z(n24259) );
  XOR U32888 ( .A(n24236), .B(n24262), .Z(N63232) );
  XNOR U32889 ( .A(n24239), .B(n24238), .Z(n24262) );
  XNOR U32890 ( .A(n24250), .B(n24263), .Z(n24238) );
  XNOR U32891 ( .A(n24254), .B(n24252), .Z(n24263) );
  XOR U32892 ( .A(n24260), .B(n24264), .Z(n24252) );
  XNOR U32893 ( .A(n24257), .B(n24261), .Z(n24264) );
  AND U32894 ( .A(n24265), .B(n24266), .Z(n24261) );
  NAND U32895 ( .A(n24267), .B(n24268), .Z(n24266) );
  NAND U32896 ( .A(n24269), .B(n24270), .Z(n24265) );
  AND U32897 ( .A(n24271), .B(n24272), .Z(n24257) );
  NAND U32898 ( .A(n24273), .B(n24274), .Z(n24272) );
  NAND U32899 ( .A(n24275), .B(n24276), .Z(n24271) );
  NANDN U32900 ( .A(n24277), .B(n24278), .Z(n24260) );
  ANDN U32901 ( .B(n24279), .A(n24280), .Z(n24254) );
  XNOR U32902 ( .A(n24245), .B(n24281), .Z(n24250) );
  XNOR U32903 ( .A(n24243), .B(n24247), .Z(n24281) );
  AND U32904 ( .A(n24282), .B(n24283), .Z(n24247) );
  NAND U32905 ( .A(n24284), .B(n24285), .Z(n24283) );
  NAND U32906 ( .A(n24286), .B(n24287), .Z(n24282) );
  AND U32907 ( .A(n24288), .B(n24289), .Z(n24243) );
  NAND U32908 ( .A(n24290), .B(n24291), .Z(n24289) );
  NAND U32909 ( .A(n24292), .B(n24293), .Z(n24288) );
  AND U32910 ( .A(n24294), .B(n24295), .Z(n24245) );
  NAND U32911 ( .A(n24296), .B(n24297), .Z(n24239) );
  XNOR U32912 ( .A(n24222), .B(n24298), .Z(n24236) );
  XNOR U32913 ( .A(n24226), .B(n24224), .Z(n24298) );
  XOR U32914 ( .A(n24232), .B(n24299), .Z(n24224) );
  XNOR U32915 ( .A(n24229), .B(n24233), .Z(n24299) );
  AND U32916 ( .A(n24300), .B(n24301), .Z(n24233) );
  NAND U32917 ( .A(n24302), .B(n24303), .Z(n24301) );
  NAND U32918 ( .A(n24304), .B(n24305), .Z(n24300) );
  AND U32919 ( .A(n24306), .B(n24307), .Z(n24229) );
  NAND U32920 ( .A(n24308), .B(n24309), .Z(n24307) );
  NAND U32921 ( .A(n24310), .B(n24311), .Z(n24306) );
  NANDN U32922 ( .A(n24312), .B(n24313), .Z(n24232) );
  ANDN U32923 ( .B(n24314), .A(n24315), .Z(n24226) );
  XNOR U32924 ( .A(n24217), .B(n24316), .Z(n24222) );
  XNOR U32925 ( .A(n24215), .B(n24219), .Z(n24316) );
  AND U32926 ( .A(n24317), .B(n24318), .Z(n24219) );
  NAND U32927 ( .A(n24319), .B(n24320), .Z(n24318) );
  NAND U32928 ( .A(n24321), .B(n24322), .Z(n24317) );
  AND U32929 ( .A(n24323), .B(n24324), .Z(n24215) );
  NAND U32930 ( .A(n24325), .B(n24326), .Z(n24324) );
  NAND U32931 ( .A(n24327), .B(n24328), .Z(n24323) );
  AND U32932 ( .A(n24329), .B(n24330), .Z(n24217) );
  XOR U32933 ( .A(n24297), .B(n24296), .Z(N63231) );
  XNOR U32934 ( .A(n24314), .B(n24315), .Z(n24296) );
  XNOR U32935 ( .A(n24329), .B(n24330), .Z(n24315) );
  XOR U32936 ( .A(n24326), .B(n24325), .Z(n24330) );
  XOR U32937 ( .A(y[4884]), .B(x[4884]), .Z(n24325) );
  XOR U32938 ( .A(n24328), .B(n24327), .Z(n24326) );
  XOR U32939 ( .A(y[4886]), .B(x[4886]), .Z(n24327) );
  XOR U32940 ( .A(y[4885]), .B(x[4885]), .Z(n24328) );
  XOR U32941 ( .A(n24320), .B(n24319), .Z(n24329) );
  XOR U32942 ( .A(n24322), .B(n24321), .Z(n24319) );
  XOR U32943 ( .A(y[4883]), .B(x[4883]), .Z(n24321) );
  XOR U32944 ( .A(y[4882]), .B(x[4882]), .Z(n24322) );
  XOR U32945 ( .A(y[4881]), .B(x[4881]), .Z(n24320) );
  XNOR U32946 ( .A(n24313), .B(n24312), .Z(n24314) );
  XNOR U32947 ( .A(n24309), .B(n24308), .Z(n24312) );
  XOR U32948 ( .A(n24311), .B(n24310), .Z(n24308) );
  XOR U32949 ( .A(y[4880]), .B(x[4880]), .Z(n24310) );
  XOR U32950 ( .A(y[4879]), .B(x[4879]), .Z(n24311) );
  XOR U32951 ( .A(y[4878]), .B(x[4878]), .Z(n24309) );
  XOR U32952 ( .A(n24303), .B(n24302), .Z(n24313) );
  XOR U32953 ( .A(n24305), .B(n24304), .Z(n24302) );
  XOR U32954 ( .A(y[4877]), .B(x[4877]), .Z(n24304) );
  XOR U32955 ( .A(y[4876]), .B(x[4876]), .Z(n24305) );
  XOR U32956 ( .A(y[4875]), .B(x[4875]), .Z(n24303) );
  XNOR U32957 ( .A(n24279), .B(n24280), .Z(n24297) );
  XNOR U32958 ( .A(n24294), .B(n24295), .Z(n24280) );
  XOR U32959 ( .A(n24291), .B(n24290), .Z(n24295) );
  XOR U32960 ( .A(y[4872]), .B(x[4872]), .Z(n24290) );
  XOR U32961 ( .A(n24293), .B(n24292), .Z(n24291) );
  XOR U32962 ( .A(y[4874]), .B(x[4874]), .Z(n24292) );
  XOR U32963 ( .A(y[4873]), .B(x[4873]), .Z(n24293) );
  XOR U32964 ( .A(n24285), .B(n24284), .Z(n24294) );
  XOR U32965 ( .A(n24287), .B(n24286), .Z(n24284) );
  XOR U32966 ( .A(y[4871]), .B(x[4871]), .Z(n24286) );
  XOR U32967 ( .A(y[4870]), .B(x[4870]), .Z(n24287) );
  XOR U32968 ( .A(y[4869]), .B(x[4869]), .Z(n24285) );
  XNOR U32969 ( .A(n24278), .B(n24277), .Z(n24279) );
  XNOR U32970 ( .A(n24274), .B(n24273), .Z(n24277) );
  XOR U32971 ( .A(n24276), .B(n24275), .Z(n24273) );
  XOR U32972 ( .A(y[4868]), .B(x[4868]), .Z(n24275) );
  XOR U32973 ( .A(y[4867]), .B(x[4867]), .Z(n24276) );
  XOR U32974 ( .A(y[4866]), .B(x[4866]), .Z(n24274) );
  XOR U32975 ( .A(n24268), .B(n24267), .Z(n24278) );
  XOR U32976 ( .A(n24270), .B(n24269), .Z(n24267) );
  XOR U32977 ( .A(y[4865]), .B(x[4865]), .Z(n24269) );
  XOR U32978 ( .A(y[4864]), .B(x[4864]), .Z(n24270) );
  XOR U32979 ( .A(y[4863]), .B(x[4863]), .Z(n24268) );
  NAND U32980 ( .A(n24331), .B(n24332), .Z(N63222) );
  NAND U32981 ( .A(n24333), .B(n24334), .Z(n24332) );
  NANDN U32982 ( .A(n24335), .B(n24336), .Z(n24334) );
  NANDN U32983 ( .A(n24336), .B(n24335), .Z(n24331) );
  XOR U32984 ( .A(n24335), .B(n24337), .Z(N63221) );
  XNOR U32985 ( .A(n24333), .B(n24336), .Z(n24337) );
  NAND U32986 ( .A(n24338), .B(n24339), .Z(n24336) );
  NAND U32987 ( .A(n24340), .B(n24341), .Z(n24339) );
  NANDN U32988 ( .A(n24342), .B(n24343), .Z(n24341) );
  NANDN U32989 ( .A(n24343), .B(n24342), .Z(n24338) );
  AND U32990 ( .A(n24344), .B(n24345), .Z(n24333) );
  NAND U32991 ( .A(n24346), .B(n24347), .Z(n24345) );
  NANDN U32992 ( .A(n24348), .B(n24349), .Z(n24347) );
  NANDN U32993 ( .A(n24349), .B(n24348), .Z(n24344) );
  IV U32994 ( .A(n24350), .Z(n24349) );
  AND U32995 ( .A(n24351), .B(n24352), .Z(n24335) );
  NAND U32996 ( .A(n24353), .B(n24354), .Z(n24352) );
  NANDN U32997 ( .A(n24355), .B(n24356), .Z(n24354) );
  NANDN U32998 ( .A(n24356), .B(n24355), .Z(n24351) );
  XOR U32999 ( .A(n24348), .B(n24357), .Z(N63220) );
  XNOR U33000 ( .A(n24346), .B(n24350), .Z(n24357) );
  XOR U33001 ( .A(n24343), .B(n24358), .Z(n24350) );
  XNOR U33002 ( .A(n24340), .B(n24342), .Z(n24358) );
  AND U33003 ( .A(n24359), .B(n24360), .Z(n24342) );
  NANDN U33004 ( .A(n24361), .B(n24362), .Z(n24360) );
  OR U33005 ( .A(n24363), .B(n24364), .Z(n24362) );
  IV U33006 ( .A(n24365), .Z(n24364) );
  NANDN U33007 ( .A(n24365), .B(n24363), .Z(n24359) );
  AND U33008 ( .A(n24366), .B(n24367), .Z(n24340) );
  NAND U33009 ( .A(n24368), .B(n24369), .Z(n24367) );
  NANDN U33010 ( .A(n24370), .B(n24371), .Z(n24369) );
  NANDN U33011 ( .A(n24371), .B(n24370), .Z(n24366) );
  IV U33012 ( .A(n24372), .Z(n24371) );
  NAND U33013 ( .A(n24373), .B(n24374), .Z(n24343) );
  NANDN U33014 ( .A(n24375), .B(n24376), .Z(n24374) );
  NANDN U33015 ( .A(n24377), .B(n24378), .Z(n24376) );
  NANDN U33016 ( .A(n24378), .B(n24377), .Z(n24373) );
  IV U33017 ( .A(n24379), .Z(n24377) );
  AND U33018 ( .A(n24380), .B(n24381), .Z(n24346) );
  NAND U33019 ( .A(n24382), .B(n24383), .Z(n24381) );
  NANDN U33020 ( .A(n24384), .B(n24385), .Z(n24383) );
  NANDN U33021 ( .A(n24385), .B(n24384), .Z(n24380) );
  XOR U33022 ( .A(n24356), .B(n24386), .Z(n24348) );
  XNOR U33023 ( .A(n24353), .B(n24355), .Z(n24386) );
  AND U33024 ( .A(n24387), .B(n24388), .Z(n24355) );
  NANDN U33025 ( .A(n24389), .B(n24390), .Z(n24388) );
  OR U33026 ( .A(n24391), .B(n24392), .Z(n24390) );
  IV U33027 ( .A(n24393), .Z(n24392) );
  NANDN U33028 ( .A(n24393), .B(n24391), .Z(n24387) );
  AND U33029 ( .A(n24394), .B(n24395), .Z(n24353) );
  NAND U33030 ( .A(n24396), .B(n24397), .Z(n24395) );
  NANDN U33031 ( .A(n24398), .B(n24399), .Z(n24397) );
  NANDN U33032 ( .A(n24399), .B(n24398), .Z(n24394) );
  IV U33033 ( .A(n24400), .Z(n24399) );
  NAND U33034 ( .A(n24401), .B(n24402), .Z(n24356) );
  NANDN U33035 ( .A(n24403), .B(n24404), .Z(n24402) );
  NANDN U33036 ( .A(n24405), .B(n24406), .Z(n24404) );
  NANDN U33037 ( .A(n24406), .B(n24405), .Z(n24401) );
  IV U33038 ( .A(n24407), .Z(n24405) );
  XOR U33039 ( .A(n24382), .B(n24408), .Z(N63219) );
  XNOR U33040 ( .A(n24385), .B(n24384), .Z(n24408) );
  XNOR U33041 ( .A(n24396), .B(n24409), .Z(n24384) );
  XNOR U33042 ( .A(n24400), .B(n24398), .Z(n24409) );
  XOR U33043 ( .A(n24406), .B(n24410), .Z(n24398) );
  XNOR U33044 ( .A(n24403), .B(n24407), .Z(n24410) );
  AND U33045 ( .A(n24411), .B(n24412), .Z(n24407) );
  NAND U33046 ( .A(n24413), .B(n24414), .Z(n24412) );
  NAND U33047 ( .A(n24415), .B(n24416), .Z(n24411) );
  AND U33048 ( .A(n24417), .B(n24418), .Z(n24403) );
  NAND U33049 ( .A(n24419), .B(n24420), .Z(n24418) );
  NAND U33050 ( .A(n24421), .B(n24422), .Z(n24417) );
  NANDN U33051 ( .A(n24423), .B(n24424), .Z(n24406) );
  ANDN U33052 ( .B(n24425), .A(n24426), .Z(n24400) );
  XNOR U33053 ( .A(n24391), .B(n24427), .Z(n24396) );
  XNOR U33054 ( .A(n24389), .B(n24393), .Z(n24427) );
  AND U33055 ( .A(n24428), .B(n24429), .Z(n24393) );
  NAND U33056 ( .A(n24430), .B(n24431), .Z(n24429) );
  NAND U33057 ( .A(n24432), .B(n24433), .Z(n24428) );
  AND U33058 ( .A(n24434), .B(n24435), .Z(n24389) );
  NAND U33059 ( .A(n24436), .B(n24437), .Z(n24435) );
  NAND U33060 ( .A(n24438), .B(n24439), .Z(n24434) );
  AND U33061 ( .A(n24440), .B(n24441), .Z(n24391) );
  NAND U33062 ( .A(n24442), .B(n24443), .Z(n24385) );
  XNOR U33063 ( .A(n24368), .B(n24444), .Z(n24382) );
  XNOR U33064 ( .A(n24372), .B(n24370), .Z(n24444) );
  XOR U33065 ( .A(n24378), .B(n24445), .Z(n24370) );
  XNOR U33066 ( .A(n24375), .B(n24379), .Z(n24445) );
  AND U33067 ( .A(n24446), .B(n24447), .Z(n24379) );
  NAND U33068 ( .A(n24448), .B(n24449), .Z(n24447) );
  NAND U33069 ( .A(n24450), .B(n24451), .Z(n24446) );
  AND U33070 ( .A(n24452), .B(n24453), .Z(n24375) );
  NAND U33071 ( .A(n24454), .B(n24455), .Z(n24453) );
  NAND U33072 ( .A(n24456), .B(n24457), .Z(n24452) );
  NANDN U33073 ( .A(n24458), .B(n24459), .Z(n24378) );
  ANDN U33074 ( .B(n24460), .A(n24461), .Z(n24372) );
  XNOR U33075 ( .A(n24363), .B(n24462), .Z(n24368) );
  XNOR U33076 ( .A(n24361), .B(n24365), .Z(n24462) );
  AND U33077 ( .A(n24463), .B(n24464), .Z(n24365) );
  NAND U33078 ( .A(n24465), .B(n24466), .Z(n24464) );
  NAND U33079 ( .A(n24467), .B(n24468), .Z(n24463) );
  AND U33080 ( .A(n24469), .B(n24470), .Z(n24361) );
  NAND U33081 ( .A(n24471), .B(n24472), .Z(n24470) );
  NAND U33082 ( .A(n24473), .B(n24474), .Z(n24469) );
  AND U33083 ( .A(n24475), .B(n24476), .Z(n24363) );
  XOR U33084 ( .A(n24443), .B(n24442), .Z(N63218) );
  XNOR U33085 ( .A(n24460), .B(n24461), .Z(n24442) );
  XNOR U33086 ( .A(n24475), .B(n24476), .Z(n24461) );
  XOR U33087 ( .A(n24472), .B(n24471), .Z(n24476) );
  XOR U33088 ( .A(y[4860]), .B(x[4860]), .Z(n24471) );
  XOR U33089 ( .A(n24474), .B(n24473), .Z(n24472) );
  XOR U33090 ( .A(y[4862]), .B(x[4862]), .Z(n24473) );
  XOR U33091 ( .A(y[4861]), .B(x[4861]), .Z(n24474) );
  XOR U33092 ( .A(n24466), .B(n24465), .Z(n24475) );
  XOR U33093 ( .A(n24468), .B(n24467), .Z(n24465) );
  XOR U33094 ( .A(y[4859]), .B(x[4859]), .Z(n24467) );
  XOR U33095 ( .A(y[4858]), .B(x[4858]), .Z(n24468) );
  XOR U33096 ( .A(y[4857]), .B(x[4857]), .Z(n24466) );
  XNOR U33097 ( .A(n24459), .B(n24458), .Z(n24460) );
  XNOR U33098 ( .A(n24455), .B(n24454), .Z(n24458) );
  XOR U33099 ( .A(n24457), .B(n24456), .Z(n24454) );
  XOR U33100 ( .A(y[4856]), .B(x[4856]), .Z(n24456) );
  XOR U33101 ( .A(y[4855]), .B(x[4855]), .Z(n24457) );
  XOR U33102 ( .A(y[4854]), .B(x[4854]), .Z(n24455) );
  XOR U33103 ( .A(n24449), .B(n24448), .Z(n24459) );
  XOR U33104 ( .A(n24451), .B(n24450), .Z(n24448) );
  XOR U33105 ( .A(y[4853]), .B(x[4853]), .Z(n24450) );
  XOR U33106 ( .A(y[4852]), .B(x[4852]), .Z(n24451) );
  XOR U33107 ( .A(y[4851]), .B(x[4851]), .Z(n24449) );
  XNOR U33108 ( .A(n24425), .B(n24426), .Z(n24443) );
  XNOR U33109 ( .A(n24440), .B(n24441), .Z(n24426) );
  XOR U33110 ( .A(n24437), .B(n24436), .Z(n24441) );
  XOR U33111 ( .A(y[4848]), .B(x[4848]), .Z(n24436) );
  XOR U33112 ( .A(n24439), .B(n24438), .Z(n24437) );
  XOR U33113 ( .A(y[4850]), .B(x[4850]), .Z(n24438) );
  XOR U33114 ( .A(y[4849]), .B(x[4849]), .Z(n24439) );
  XOR U33115 ( .A(n24431), .B(n24430), .Z(n24440) );
  XOR U33116 ( .A(n24433), .B(n24432), .Z(n24430) );
  XOR U33117 ( .A(y[4847]), .B(x[4847]), .Z(n24432) );
  XOR U33118 ( .A(y[4846]), .B(x[4846]), .Z(n24433) );
  XOR U33119 ( .A(y[4845]), .B(x[4845]), .Z(n24431) );
  XNOR U33120 ( .A(n24424), .B(n24423), .Z(n24425) );
  XNOR U33121 ( .A(n24420), .B(n24419), .Z(n24423) );
  XOR U33122 ( .A(n24422), .B(n24421), .Z(n24419) );
  XOR U33123 ( .A(y[4844]), .B(x[4844]), .Z(n24421) );
  XOR U33124 ( .A(y[4843]), .B(x[4843]), .Z(n24422) );
  XOR U33125 ( .A(y[4842]), .B(x[4842]), .Z(n24420) );
  XOR U33126 ( .A(n24414), .B(n24413), .Z(n24424) );
  XOR U33127 ( .A(n24416), .B(n24415), .Z(n24413) );
  XOR U33128 ( .A(y[4841]), .B(x[4841]), .Z(n24415) );
  XOR U33129 ( .A(y[4840]), .B(x[4840]), .Z(n24416) );
  XOR U33130 ( .A(y[4839]), .B(x[4839]), .Z(n24414) );
  NAND U33131 ( .A(n24477), .B(n24478), .Z(N63209) );
  NAND U33132 ( .A(n24479), .B(n24480), .Z(n24478) );
  NANDN U33133 ( .A(n24481), .B(n24482), .Z(n24480) );
  NANDN U33134 ( .A(n24482), .B(n24481), .Z(n24477) );
  XOR U33135 ( .A(n24481), .B(n24483), .Z(N63208) );
  XNOR U33136 ( .A(n24479), .B(n24482), .Z(n24483) );
  NAND U33137 ( .A(n24484), .B(n24485), .Z(n24482) );
  NAND U33138 ( .A(n24486), .B(n24487), .Z(n24485) );
  NANDN U33139 ( .A(n24488), .B(n24489), .Z(n24487) );
  NANDN U33140 ( .A(n24489), .B(n24488), .Z(n24484) );
  AND U33141 ( .A(n24490), .B(n24491), .Z(n24479) );
  NAND U33142 ( .A(n24492), .B(n24493), .Z(n24491) );
  NANDN U33143 ( .A(n24494), .B(n24495), .Z(n24493) );
  NANDN U33144 ( .A(n24495), .B(n24494), .Z(n24490) );
  IV U33145 ( .A(n24496), .Z(n24495) );
  AND U33146 ( .A(n24497), .B(n24498), .Z(n24481) );
  NAND U33147 ( .A(n24499), .B(n24500), .Z(n24498) );
  NANDN U33148 ( .A(n24501), .B(n24502), .Z(n24500) );
  NANDN U33149 ( .A(n24502), .B(n24501), .Z(n24497) );
  XOR U33150 ( .A(n24494), .B(n24503), .Z(N63207) );
  XNOR U33151 ( .A(n24492), .B(n24496), .Z(n24503) );
  XOR U33152 ( .A(n24489), .B(n24504), .Z(n24496) );
  XNOR U33153 ( .A(n24486), .B(n24488), .Z(n24504) );
  AND U33154 ( .A(n24505), .B(n24506), .Z(n24488) );
  NANDN U33155 ( .A(n24507), .B(n24508), .Z(n24506) );
  OR U33156 ( .A(n24509), .B(n24510), .Z(n24508) );
  IV U33157 ( .A(n24511), .Z(n24510) );
  NANDN U33158 ( .A(n24511), .B(n24509), .Z(n24505) );
  AND U33159 ( .A(n24512), .B(n24513), .Z(n24486) );
  NAND U33160 ( .A(n24514), .B(n24515), .Z(n24513) );
  NANDN U33161 ( .A(n24516), .B(n24517), .Z(n24515) );
  NANDN U33162 ( .A(n24517), .B(n24516), .Z(n24512) );
  IV U33163 ( .A(n24518), .Z(n24517) );
  NAND U33164 ( .A(n24519), .B(n24520), .Z(n24489) );
  NANDN U33165 ( .A(n24521), .B(n24522), .Z(n24520) );
  NANDN U33166 ( .A(n24523), .B(n24524), .Z(n24522) );
  NANDN U33167 ( .A(n24524), .B(n24523), .Z(n24519) );
  IV U33168 ( .A(n24525), .Z(n24523) );
  AND U33169 ( .A(n24526), .B(n24527), .Z(n24492) );
  NAND U33170 ( .A(n24528), .B(n24529), .Z(n24527) );
  NANDN U33171 ( .A(n24530), .B(n24531), .Z(n24529) );
  NANDN U33172 ( .A(n24531), .B(n24530), .Z(n24526) );
  XOR U33173 ( .A(n24502), .B(n24532), .Z(n24494) );
  XNOR U33174 ( .A(n24499), .B(n24501), .Z(n24532) );
  AND U33175 ( .A(n24533), .B(n24534), .Z(n24501) );
  NANDN U33176 ( .A(n24535), .B(n24536), .Z(n24534) );
  OR U33177 ( .A(n24537), .B(n24538), .Z(n24536) );
  IV U33178 ( .A(n24539), .Z(n24538) );
  NANDN U33179 ( .A(n24539), .B(n24537), .Z(n24533) );
  AND U33180 ( .A(n24540), .B(n24541), .Z(n24499) );
  NAND U33181 ( .A(n24542), .B(n24543), .Z(n24541) );
  NANDN U33182 ( .A(n24544), .B(n24545), .Z(n24543) );
  NANDN U33183 ( .A(n24545), .B(n24544), .Z(n24540) );
  IV U33184 ( .A(n24546), .Z(n24545) );
  NAND U33185 ( .A(n24547), .B(n24548), .Z(n24502) );
  NANDN U33186 ( .A(n24549), .B(n24550), .Z(n24548) );
  NANDN U33187 ( .A(n24551), .B(n24552), .Z(n24550) );
  NANDN U33188 ( .A(n24552), .B(n24551), .Z(n24547) );
  IV U33189 ( .A(n24553), .Z(n24551) );
  XOR U33190 ( .A(n24528), .B(n24554), .Z(N63206) );
  XNOR U33191 ( .A(n24531), .B(n24530), .Z(n24554) );
  XNOR U33192 ( .A(n24542), .B(n24555), .Z(n24530) );
  XNOR U33193 ( .A(n24546), .B(n24544), .Z(n24555) );
  XOR U33194 ( .A(n24552), .B(n24556), .Z(n24544) );
  XNOR U33195 ( .A(n24549), .B(n24553), .Z(n24556) );
  AND U33196 ( .A(n24557), .B(n24558), .Z(n24553) );
  NAND U33197 ( .A(n24559), .B(n24560), .Z(n24558) );
  NAND U33198 ( .A(n24561), .B(n24562), .Z(n24557) );
  AND U33199 ( .A(n24563), .B(n24564), .Z(n24549) );
  NAND U33200 ( .A(n24565), .B(n24566), .Z(n24564) );
  NAND U33201 ( .A(n24567), .B(n24568), .Z(n24563) );
  NANDN U33202 ( .A(n24569), .B(n24570), .Z(n24552) );
  ANDN U33203 ( .B(n24571), .A(n24572), .Z(n24546) );
  XNOR U33204 ( .A(n24537), .B(n24573), .Z(n24542) );
  XNOR U33205 ( .A(n24535), .B(n24539), .Z(n24573) );
  AND U33206 ( .A(n24574), .B(n24575), .Z(n24539) );
  NAND U33207 ( .A(n24576), .B(n24577), .Z(n24575) );
  NAND U33208 ( .A(n24578), .B(n24579), .Z(n24574) );
  AND U33209 ( .A(n24580), .B(n24581), .Z(n24535) );
  NAND U33210 ( .A(n24582), .B(n24583), .Z(n24581) );
  NAND U33211 ( .A(n24584), .B(n24585), .Z(n24580) );
  AND U33212 ( .A(n24586), .B(n24587), .Z(n24537) );
  NAND U33213 ( .A(n24588), .B(n24589), .Z(n24531) );
  XNOR U33214 ( .A(n24514), .B(n24590), .Z(n24528) );
  XNOR U33215 ( .A(n24518), .B(n24516), .Z(n24590) );
  XOR U33216 ( .A(n24524), .B(n24591), .Z(n24516) );
  XNOR U33217 ( .A(n24521), .B(n24525), .Z(n24591) );
  AND U33218 ( .A(n24592), .B(n24593), .Z(n24525) );
  NAND U33219 ( .A(n24594), .B(n24595), .Z(n24593) );
  NAND U33220 ( .A(n24596), .B(n24597), .Z(n24592) );
  AND U33221 ( .A(n24598), .B(n24599), .Z(n24521) );
  NAND U33222 ( .A(n24600), .B(n24601), .Z(n24599) );
  NAND U33223 ( .A(n24602), .B(n24603), .Z(n24598) );
  NANDN U33224 ( .A(n24604), .B(n24605), .Z(n24524) );
  ANDN U33225 ( .B(n24606), .A(n24607), .Z(n24518) );
  XNOR U33226 ( .A(n24509), .B(n24608), .Z(n24514) );
  XNOR U33227 ( .A(n24507), .B(n24511), .Z(n24608) );
  AND U33228 ( .A(n24609), .B(n24610), .Z(n24511) );
  NAND U33229 ( .A(n24611), .B(n24612), .Z(n24610) );
  NAND U33230 ( .A(n24613), .B(n24614), .Z(n24609) );
  AND U33231 ( .A(n24615), .B(n24616), .Z(n24507) );
  NAND U33232 ( .A(n24617), .B(n24618), .Z(n24616) );
  NAND U33233 ( .A(n24619), .B(n24620), .Z(n24615) );
  AND U33234 ( .A(n24621), .B(n24622), .Z(n24509) );
  XOR U33235 ( .A(n24589), .B(n24588), .Z(N63205) );
  XNOR U33236 ( .A(n24606), .B(n24607), .Z(n24588) );
  XNOR U33237 ( .A(n24621), .B(n24622), .Z(n24607) );
  XOR U33238 ( .A(n24618), .B(n24617), .Z(n24622) );
  XOR U33239 ( .A(y[4836]), .B(x[4836]), .Z(n24617) );
  XOR U33240 ( .A(n24620), .B(n24619), .Z(n24618) );
  XOR U33241 ( .A(y[4838]), .B(x[4838]), .Z(n24619) );
  XOR U33242 ( .A(y[4837]), .B(x[4837]), .Z(n24620) );
  XOR U33243 ( .A(n24612), .B(n24611), .Z(n24621) );
  XOR U33244 ( .A(n24614), .B(n24613), .Z(n24611) );
  XOR U33245 ( .A(y[4835]), .B(x[4835]), .Z(n24613) );
  XOR U33246 ( .A(y[4834]), .B(x[4834]), .Z(n24614) );
  XOR U33247 ( .A(y[4833]), .B(x[4833]), .Z(n24612) );
  XNOR U33248 ( .A(n24605), .B(n24604), .Z(n24606) );
  XNOR U33249 ( .A(n24601), .B(n24600), .Z(n24604) );
  XOR U33250 ( .A(n24603), .B(n24602), .Z(n24600) );
  XOR U33251 ( .A(y[4832]), .B(x[4832]), .Z(n24602) );
  XOR U33252 ( .A(y[4831]), .B(x[4831]), .Z(n24603) );
  XOR U33253 ( .A(y[4830]), .B(x[4830]), .Z(n24601) );
  XOR U33254 ( .A(n24595), .B(n24594), .Z(n24605) );
  XOR U33255 ( .A(n24597), .B(n24596), .Z(n24594) );
  XOR U33256 ( .A(y[4829]), .B(x[4829]), .Z(n24596) );
  XOR U33257 ( .A(y[4828]), .B(x[4828]), .Z(n24597) );
  XOR U33258 ( .A(y[4827]), .B(x[4827]), .Z(n24595) );
  XNOR U33259 ( .A(n24571), .B(n24572), .Z(n24589) );
  XNOR U33260 ( .A(n24586), .B(n24587), .Z(n24572) );
  XOR U33261 ( .A(n24583), .B(n24582), .Z(n24587) );
  XOR U33262 ( .A(y[4824]), .B(x[4824]), .Z(n24582) );
  XOR U33263 ( .A(n24585), .B(n24584), .Z(n24583) );
  XOR U33264 ( .A(y[4826]), .B(x[4826]), .Z(n24584) );
  XOR U33265 ( .A(y[4825]), .B(x[4825]), .Z(n24585) );
  XOR U33266 ( .A(n24577), .B(n24576), .Z(n24586) );
  XOR U33267 ( .A(n24579), .B(n24578), .Z(n24576) );
  XOR U33268 ( .A(y[4823]), .B(x[4823]), .Z(n24578) );
  XOR U33269 ( .A(y[4822]), .B(x[4822]), .Z(n24579) );
  XOR U33270 ( .A(y[4821]), .B(x[4821]), .Z(n24577) );
  XNOR U33271 ( .A(n24570), .B(n24569), .Z(n24571) );
  XNOR U33272 ( .A(n24566), .B(n24565), .Z(n24569) );
  XOR U33273 ( .A(n24568), .B(n24567), .Z(n24565) );
  XOR U33274 ( .A(y[4820]), .B(x[4820]), .Z(n24567) );
  XOR U33275 ( .A(y[4819]), .B(x[4819]), .Z(n24568) );
  XOR U33276 ( .A(y[4818]), .B(x[4818]), .Z(n24566) );
  XOR U33277 ( .A(n24560), .B(n24559), .Z(n24570) );
  XOR U33278 ( .A(n24562), .B(n24561), .Z(n24559) );
  XOR U33279 ( .A(y[4817]), .B(x[4817]), .Z(n24561) );
  XOR U33280 ( .A(y[4816]), .B(x[4816]), .Z(n24562) );
  XOR U33281 ( .A(y[4815]), .B(x[4815]), .Z(n24560) );
  NAND U33282 ( .A(n24623), .B(n24624), .Z(N63196) );
  NAND U33283 ( .A(n24625), .B(n24626), .Z(n24624) );
  NANDN U33284 ( .A(n24627), .B(n24628), .Z(n24626) );
  NANDN U33285 ( .A(n24628), .B(n24627), .Z(n24623) );
  XOR U33286 ( .A(n24627), .B(n24629), .Z(N63195) );
  XNOR U33287 ( .A(n24625), .B(n24628), .Z(n24629) );
  NAND U33288 ( .A(n24630), .B(n24631), .Z(n24628) );
  NAND U33289 ( .A(n24632), .B(n24633), .Z(n24631) );
  NANDN U33290 ( .A(n24634), .B(n24635), .Z(n24633) );
  NANDN U33291 ( .A(n24635), .B(n24634), .Z(n24630) );
  AND U33292 ( .A(n24636), .B(n24637), .Z(n24625) );
  NAND U33293 ( .A(n24638), .B(n24639), .Z(n24637) );
  NANDN U33294 ( .A(n24640), .B(n24641), .Z(n24639) );
  NANDN U33295 ( .A(n24641), .B(n24640), .Z(n24636) );
  IV U33296 ( .A(n24642), .Z(n24641) );
  AND U33297 ( .A(n24643), .B(n24644), .Z(n24627) );
  NAND U33298 ( .A(n24645), .B(n24646), .Z(n24644) );
  NANDN U33299 ( .A(n24647), .B(n24648), .Z(n24646) );
  NANDN U33300 ( .A(n24648), .B(n24647), .Z(n24643) );
  XOR U33301 ( .A(n24640), .B(n24649), .Z(N63194) );
  XNOR U33302 ( .A(n24638), .B(n24642), .Z(n24649) );
  XOR U33303 ( .A(n24635), .B(n24650), .Z(n24642) );
  XNOR U33304 ( .A(n24632), .B(n24634), .Z(n24650) );
  AND U33305 ( .A(n24651), .B(n24652), .Z(n24634) );
  NANDN U33306 ( .A(n24653), .B(n24654), .Z(n24652) );
  OR U33307 ( .A(n24655), .B(n24656), .Z(n24654) );
  IV U33308 ( .A(n24657), .Z(n24656) );
  NANDN U33309 ( .A(n24657), .B(n24655), .Z(n24651) );
  AND U33310 ( .A(n24658), .B(n24659), .Z(n24632) );
  NAND U33311 ( .A(n24660), .B(n24661), .Z(n24659) );
  NANDN U33312 ( .A(n24662), .B(n24663), .Z(n24661) );
  NANDN U33313 ( .A(n24663), .B(n24662), .Z(n24658) );
  IV U33314 ( .A(n24664), .Z(n24663) );
  NAND U33315 ( .A(n24665), .B(n24666), .Z(n24635) );
  NANDN U33316 ( .A(n24667), .B(n24668), .Z(n24666) );
  NANDN U33317 ( .A(n24669), .B(n24670), .Z(n24668) );
  NANDN U33318 ( .A(n24670), .B(n24669), .Z(n24665) );
  IV U33319 ( .A(n24671), .Z(n24669) );
  AND U33320 ( .A(n24672), .B(n24673), .Z(n24638) );
  NAND U33321 ( .A(n24674), .B(n24675), .Z(n24673) );
  NANDN U33322 ( .A(n24676), .B(n24677), .Z(n24675) );
  NANDN U33323 ( .A(n24677), .B(n24676), .Z(n24672) );
  XOR U33324 ( .A(n24648), .B(n24678), .Z(n24640) );
  XNOR U33325 ( .A(n24645), .B(n24647), .Z(n24678) );
  AND U33326 ( .A(n24679), .B(n24680), .Z(n24647) );
  NANDN U33327 ( .A(n24681), .B(n24682), .Z(n24680) );
  OR U33328 ( .A(n24683), .B(n24684), .Z(n24682) );
  IV U33329 ( .A(n24685), .Z(n24684) );
  NANDN U33330 ( .A(n24685), .B(n24683), .Z(n24679) );
  AND U33331 ( .A(n24686), .B(n24687), .Z(n24645) );
  NAND U33332 ( .A(n24688), .B(n24689), .Z(n24687) );
  NANDN U33333 ( .A(n24690), .B(n24691), .Z(n24689) );
  NANDN U33334 ( .A(n24691), .B(n24690), .Z(n24686) );
  IV U33335 ( .A(n24692), .Z(n24691) );
  NAND U33336 ( .A(n24693), .B(n24694), .Z(n24648) );
  NANDN U33337 ( .A(n24695), .B(n24696), .Z(n24694) );
  NANDN U33338 ( .A(n24697), .B(n24698), .Z(n24696) );
  NANDN U33339 ( .A(n24698), .B(n24697), .Z(n24693) );
  IV U33340 ( .A(n24699), .Z(n24697) );
  XOR U33341 ( .A(n24674), .B(n24700), .Z(N63193) );
  XNOR U33342 ( .A(n24677), .B(n24676), .Z(n24700) );
  XNOR U33343 ( .A(n24688), .B(n24701), .Z(n24676) );
  XNOR U33344 ( .A(n24692), .B(n24690), .Z(n24701) );
  XOR U33345 ( .A(n24698), .B(n24702), .Z(n24690) );
  XNOR U33346 ( .A(n24695), .B(n24699), .Z(n24702) );
  AND U33347 ( .A(n24703), .B(n24704), .Z(n24699) );
  NAND U33348 ( .A(n24705), .B(n24706), .Z(n24704) );
  NAND U33349 ( .A(n24707), .B(n24708), .Z(n24703) );
  AND U33350 ( .A(n24709), .B(n24710), .Z(n24695) );
  NAND U33351 ( .A(n24711), .B(n24712), .Z(n24710) );
  NAND U33352 ( .A(n24713), .B(n24714), .Z(n24709) );
  NANDN U33353 ( .A(n24715), .B(n24716), .Z(n24698) );
  ANDN U33354 ( .B(n24717), .A(n24718), .Z(n24692) );
  XNOR U33355 ( .A(n24683), .B(n24719), .Z(n24688) );
  XNOR U33356 ( .A(n24681), .B(n24685), .Z(n24719) );
  AND U33357 ( .A(n24720), .B(n24721), .Z(n24685) );
  NAND U33358 ( .A(n24722), .B(n24723), .Z(n24721) );
  NAND U33359 ( .A(n24724), .B(n24725), .Z(n24720) );
  AND U33360 ( .A(n24726), .B(n24727), .Z(n24681) );
  NAND U33361 ( .A(n24728), .B(n24729), .Z(n24727) );
  NAND U33362 ( .A(n24730), .B(n24731), .Z(n24726) );
  AND U33363 ( .A(n24732), .B(n24733), .Z(n24683) );
  NAND U33364 ( .A(n24734), .B(n24735), .Z(n24677) );
  XNOR U33365 ( .A(n24660), .B(n24736), .Z(n24674) );
  XNOR U33366 ( .A(n24664), .B(n24662), .Z(n24736) );
  XOR U33367 ( .A(n24670), .B(n24737), .Z(n24662) );
  XNOR U33368 ( .A(n24667), .B(n24671), .Z(n24737) );
  AND U33369 ( .A(n24738), .B(n24739), .Z(n24671) );
  NAND U33370 ( .A(n24740), .B(n24741), .Z(n24739) );
  NAND U33371 ( .A(n24742), .B(n24743), .Z(n24738) );
  AND U33372 ( .A(n24744), .B(n24745), .Z(n24667) );
  NAND U33373 ( .A(n24746), .B(n24747), .Z(n24745) );
  NAND U33374 ( .A(n24748), .B(n24749), .Z(n24744) );
  NANDN U33375 ( .A(n24750), .B(n24751), .Z(n24670) );
  ANDN U33376 ( .B(n24752), .A(n24753), .Z(n24664) );
  XNOR U33377 ( .A(n24655), .B(n24754), .Z(n24660) );
  XNOR U33378 ( .A(n24653), .B(n24657), .Z(n24754) );
  AND U33379 ( .A(n24755), .B(n24756), .Z(n24657) );
  NAND U33380 ( .A(n24757), .B(n24758), .Z(n24756) );
  NAND U33381 ( .A(n24759), .B(n24760), .Z(n24755) );
  AND U33382 ( .A(n24761), .B(n24762), .Z(n24653) );
  NAND U33383 ( .A(n24763), .B(n24764), .Z(n24762) );
  NAND U33384 ( .A(n24765), .B(n24766), .Z(n24761) );
  AND U33385 ( .A(n24767), .B(n24768), .Z(n24655) );
  XOR U33386 ( .A(n24735), .B(n24734), .Z(N63192) );
  XNOR U33387 ( .A(n24752), .B(n24753), .Z(n24734) );
  XNOR U33388 ( .A(n24767), .B(n24768), .Z(n24753) );
  XOR U33389 ( .A(n24764), .B(n24763), .Z(n24768) );
  XOR U33390 ( .A(y[4812]), .B(x[4812]), .Z(n24763) );
  XOR U33391 ( .A(n24766), .B(n24765), .Z(n24764) );
  XOR U33392 ( .A(y[4814]), .B(x[4814]), .Z(n24765) );
  XOR U33393 ( .A(y[4813]), .B(x[4813]), .Z(n24766) );
  XOR U33394 ( .A(n24758), .B(n24757), .Z(n24767) );
  XOR U33395 ( .A(n24760), .B(n24759), .Z(n24757) );
  XOR U33396 ( .A(y[4811]), .B(x[4811]), .Z(n24759) );
  XOR U33397 ( .A(y[4810]), .B(x[4810]), .Z(n24760) );
  XOR U33398 ( .A(y[4809]), .B(x[4809]), .Z(n24758) );
  XNOR U33399 ( .A(n24751), .B(n24750), .Z(n24752) );
  XNOR U33400 ( .A(n24747), .B(n24746), .Z(n24750) );
  XOR U33401 ( .A(n24749), .B(n24748), .Z(n24746) );
  XOR U33402 ( .A(y[4808]), .B(x[4808]), .Z(n24748) );
  XOR U33403 ( .A(y[4807]), .B(x[4807]), .Z(n24749) );
  XOR U33404 ( .A(y[4806]), .B(x[4806]), .Z(n24747) );
  XOR U33405 ( .A(n24741), .B(n24740), .Z(n24751) );
  XOR U33406 ( .A(n24743), .B(n24742), .Z(n24740) );
  XOR U33407 ( .A(y[4805]), .B(x[4805]), .Z(n24742) );
  XOR U33408 ( .A(y[4804]), .B(x[4804]), .Z(n24743) );
  XOR U33409 ( .A(y[4803]), .B(x[4803]), .Z(n24741) );
  XNOR U33410 ( .A(n24717), .B(n24718), .Z(n24735) );
  XNOR U33411 ( .A(n24732), .B(n24733), .Z(n24718) );
  XOR U33412 ( .A(n24729), .B(n24728), .Z(n24733) );
  XOR U33413 ( .A(y[4800]), .B(x[4800]), .Z(n24728) );
  XOR U33414 ( .A(n24731), .B(n24730), .Z(n24729) );
  XOR U33415 ( .A(y[4802]), .B(x[4802]), .Z(n24730) );
  XOR U33416 ( .A(y[4801]), .B(x[4801]), .Z(n24731) );
  XOR U33417 ( .A(n24723), .B(n24722), .Z(n24732) );
  XOR U33418 ( .A(n24725), .B(n24724), .Z(n24722) );
  XOR U33419 ( .A(y[4799]), .B(x[4799]), .Z(n24724) );
  XOR U33420 ( .A(y[4798]), .B(x[4798]), .Z(n24725) );
  XOR U33421 ( .A(y[4797]), .B(x[4797]), .Z(n24723) );
  XNOR U33422 ( .A(n24716), .B(n24715), .Z(n24717) );
  XNOR U33423 ( .A(n24712), .B(n24711), .Z(n24715) );
  XOR U33424 ( .A(n24714), .B(n24713), .Z(n24711) );
  XOR U33425 ( .A(y[4796]), .B(x[4796]), .Z(n24713) );
  XOR U33426 ( .A(y[4795]), .B(x[4795]), .Z(n24714) );
  XOR U33427 ( .A(y[4794]), .B(x[4794]), .Z(n24712) );
  XOR U33428 ( .A(n24706), .B(n24705), .Z(n24716) );
  XOR U33429 ( .A(n24708), .B(n24707), .Z(n24705) );
  XOR U33430 ( .A(y[4793]), .B(x[4793]), .Z(n24707) );
  XOR U33431 ( .A(y[4792]), .B(x[4792]), .Z(n24708) );
  XOR U33432 ( .A(y[4791]), .B(x[4791]), .Z(n24706) );
  NAND U33433 ( .A(n24769), .B(n24770), .Z(N63183) );
  NAND U33434 ( .A(n24771), .B(n24772), .Z(n24770) );
  NANDN U33435 ( .A(n24773), .B(n24774), .Z(n24772) );
  NANDN U33436 ( .A(n24774), .B(n24773), .Z(n24769) );
  XOR U33437 ( .A(n24773), .B(n24775), .Z(N63182) );
  XNOR U33438 ( .A(n24771), .B(n24774), .Z(n24775) );
  NAND U33439 ( .A(n24776), .B(n24777), .Z(n24774) );
  NAND U33440 ( .A(n24778), .B(n24779), .Z(n24777) );
  NANDN U33441 ( .A(n24780), .B(n24781), .Z(n24779) );
  NANDN U33442 ( .A(n24781), .B(n24780), .Z(n24776) );
  AND U33443 ( .A(n24782), .B(n24783), .Z(n24771) );
  NAND U33444 ( .A(n24784), .B(n24785), .Z(n24783) );
  NANDN U33445 ( .A(n24786), .B(n24787), .Z(n24785) );
  NANDN U33446 ( .A(n24787), .B(n24786), .Z(n24782) );
  IV U33447 ( .A(n24788), .Z(n24787) );
  AND U33448 ( .A(n24789), .B(n24790), .Z(n24773) );
  NAND U33449 ( .A(n24791), .B(n24792), .Z(n24790) );
  NANDN U33450 ( .A(n24793), .B(n24794), .Z(n24792) );
  NANDN U33451 ( .A(n24794), .B(n24793), .Z(n24789) );
  XOR U33452 ( .A(n24786), .B(n24795), .Z(N63181) );
  XNOR U33453 ( .A(n24784), .B(n24788), .Z(n24795) );
  XOR U33454 ( .A(n24781), .B(n24796), .Z(n24788) );
  XNOR U33455 ( .A(n24778), .B(n24780), .Z(n24796) );
  AND U33456 ( .A(n24797), .B(n24798), .Z(n24780) );
  NANDN U33457 ( .A(n24799), .B(n24800), .Z(n24798) );
  OR U33458 ( .A(n24801), .B(n24802), .Z(n24800) );
  IV U33459 ( .A(n24803), .Z(n24802) );
  NANDN U33460 ( .A(n24803), .B(n24801), .Z(n24797) );
  AND U33461 ( .A(n24804), .B(n24805), .Z(n24778) );
  NAND U33462 ( .A(n24806), .B(n24807), .Z(n24805) );
  NANDN U33463 ( .A(n24808), .B(n24809), .Z(n24807) );
  NANDN U33464 ( .A(n24809), .B(n24808), .Z(n24804) );
  IV U33465 ( .A(n24810), .Z(n24809) );
  NAND U33466 ( .A(n24811), .B(n24812), .Z(n24781) );
  NANDN U33467 ( .A(n24813), .B(n24814), .Z(n24812) );
  NANDN U33468 ( .A(n24815), .B(n24816), .Z(n24814) );
  NANDN U33469 ( .A(n24816), .B(n24815), .Z(n24811) );
  IV U33470 ( .A(n24817), .Z(n24815) );
  AND U33471 ( .A(n24818), .B(n24819), .Z(n24784) );
  NAND U33472 ( .A(n24820), .B(n24821), .Z(n24819) );
  NANDN U33473 ( .A(n24822), .B(n24823), .Z(n24821) );
  NANDN U33474 ( .A(n24823), .B(n24822), .Z(n24818) );
  XOR U33475 ( .A(n24794), .B(n24824), .Z(n24786) );
  XNOR U33476 ( .A(n24791), .B(n24793), .Z(n24824) );
  AND U33477 ( .A(n24825), .B(n24826), .Z(n24793) );
  NANDN U33478 ( .A(n24827), .B(n24828), .Z(n24826) );
  OR U33479 ( .A(n24829), .B(n24830), .Z(n24828) );
  IV U33480 ( .A(n24831), .Z(n24830) );
  NANDN U33481 ( .A(n24831), .B(n24829), .Z(n24825) );
  AND U33482 ( .A(n24832), .B(n24833), .Z(n24791) );
  NAND U33483 ( .A(n24834), .B(n24835), .Z(n24833) );
  NANDN U33484 ( .A(n24836), .B(n24837), .Z(n24835) );
  NANDN U33485 ( .A(n24837), .B(n24836), .Z(n24832) );
  IV U33486 ( .A(n24838), .Z(n24837) );
  NAND U33487 ( .A(n24839), .B(n24840), .Z(n24794) );
  NANDN U33488 ( .A(n24841), .B(n24842), .Z(n24840) );
  NANDN U33489 ( .A(n24843), .B(n24844), .Z(n24842) );
  NANDN U33490 ( .A(n24844), .B(n24843), .Z(n24839) );
  IV U33491 ( .A(n24845), .Z(n24843) );
  XOR U33492 ( .A(n24820), .B(n24846), .Z(N63180) );
  XNOR U33493 ( .A(n24823), .B(n24822), .Z(n24846) );
  XNOR U33494 ( .A(n24834), .B(n24847), .Z(n24822) );
  XNOR U33495 ( .A(n24838), .B(n24836), .Z(n24847) );
  XOR U33496 ( .A(n24844), .B(n24848), .Z(n24836) );
  XNOR U33497 ( .A(n24841), .B(n24845), .Z(n24848) );
  AND U33498 ( .A(n24849), .B(n24850), .Z(n24845) );
  NAND U33499 ( .A(n24851), .B(n24852), .Z(n24850) );
  NAND U33500 ( .A(n24853), .B(n24854), .Z(n24849) );
  AND U33501 ( .A(n24855), .B(n24856), .Z(n24841) );
  NAND U33502 ( .A(n24857), .B(n24858), .Z(n24856) );
  NAND U33503 ( .A(n24859), .B(n24860), .Z(n24855) );
  NANDN U33504 ( .A(n24861), .B(n24862), .Z(n24844) );
  ANDN U33505 ( .B(n24863), .A(n24864), .Z(n24838) );
  XNOR U33506 ( .A(n24829), .B(n24865), .Z(n24834) );
  XNOR U33507 ( .A(n24827), .B(n24831), .Z(n24865) );
  AND U33508 ( .A(n24866), .B(n24867), .Z(n24831) );
  NAND U33509 ( .A(n24868), .B(n24869), .Z(n24867) );
  NAND U33510 ( .A(n24870), .B(n24871), .Z(n24866) );
  AND U33511 ( .A(n24872), .B(n24873), .Z(n24827) );
  NAND U33512 ( .A(n24874), .B(n24875), .Z(n24873) );
  NAND U33513 ( .A(n24876), .B(n24877), .Z(n24872) );
  AND U33514 ( .A(n24878), .B(n24879), .Z(n24829) );
  NAND U33515 ( .A(n24880), .B(n24881), .Z(n24823) );
  XNOR U33516 ( .A(n24806), .B(n24882), .Z(n24820) );
  XNOR U33517 ( .A(n24810), .B(n24808), .Z(n24882) );
  XOR U33518 ( .A(n24816), .B(n24883), .Z(n24808) );
  XNOR U33519 ( .A(n24813), .B(n24817), .Z(n24883) );
  AND U33520 ( .A(n24884), .B(n24885), .Z(n24817) );
  NAND U33521 ( .A(n24886), .B(n24887), .Z(n24885) );
  NAND U33522 ( .A(n24888), .B(n24889), .Z(n24884) );
  AND U33523 ( .A(n24890), .B(n24891), .Z(n24813) );
  NAND U33524 ( .A(n24892), .B(n24893), .Z(n24891) );
  NAND U33525 ( .A(n24894), .B(n24895), .Z(n24890) );
  NANDN U33526 ( .A(n24896), .B(n24897), .Z(n24816) );
  ANDN U33527 ( .B(n24898), .A(n24899), .Z(n24810) );
  XNOR U33528 ( .A(n24801), .B(n24900), .Z(n24806) );
  XNOR U33529 ( .A(n24799), .B(n24803), .Z(n24900) );
  AND U33530 ( .A(n24901), .B(n24902), .Z(n24803) );
  NAND U33531 ( .A(n24903), .B(n24904), .Z(n24902) );
  NAND U33532 ( .A(n24905), .B(n24906), .Z(n24901) );
  AND U33533 ( .A(n24907), .B(n24908), .Z(n24799) );
  NAND U33534 ( .A(n24909), .B(n24910), .Z(n24908) );
  NAND U33535 ( .A(n24911), .B(n24912), .Z(n24907) );
  AND U33536 ( .A(n24913), .B(n24914), .Z(n24801) );
  XOR U33537 ( .A(n24881), .B(n24880), .Z(N63179) );
  XNOR U33538 ( .A(n24898), .B(n24899), .Z(n24880) );
  XNOR U33539 ( .A(n24913), .B(n24914), .Z(n24899) );
  XOR U33540 ( .A(n24910), .B(n24909), .Z(n24914) );
  XOR U33541 ( .A(y[4788]), .B(x[4788]), .Z(n24909) );
  XOR U33542 ( .A(n24912), .B(n24911), .Z(n24910) );
  XOR U33543 ( .A(y[4790]), .B(x[4790]), .Z(n24911) );
  XOR U33544 ( .A(y[4789]), .B(x[4789]), .Z(n24912) );
  XOR U33545 ( .A(n24904), .B(n24903), .Z(n24913) );
  XOR U33546 ( .A(n24906), .B(n24905), .Z(n24903) );
  XOR U33547 ( .A(y[4787]), .B(x[4787]), .Z(n24905) );
  XOR U33548 ( .A(y[4786]), .B(x[4786]), .Z(n24906) );
  XOR U33549 ( .A(y[4785]), .B(x[4785]), .Z(n24904) );
  XNOR U33550 ( .A(n24897), .B(n24896), .Z(n24898) );
  XNOR U33551 ( .A(n24893), .B(n24892), .Z(n24896) );
  XOR U33552 ( .A(n24895), .B(n24894), .Z(n24892) );
  XOR U33553 ( .A(y[4784]), .B(x[4784]), .Z(n24894) );
  XOR U33554 ( .A(y[4783]), .B(x[4783]), .Z(n24895) );
  XOR U33555 ( .A(y[4782]), .B(x[4782]), .Z(n24893) );
  XOR U33556 ( .A(n24887), .B(n24886), .Z(n24897) );
  XOR U33557 ( .A(n24889), .B(n24888), .Z(n24886) );
  XOR U33558 ( .A(y[4781]), .B(x[4781]), .Z(n24888) );
  XOR U33559 ( .A(y[4780]), .B(x[4780]), .Z(n24889) );
  XOR U33560 ( .A(y[4779]), .B(x[4779]), .Z(n24887) );
  XNOR U33561 ( .A(n24863), .B(n24864), .Z(n24881) );
  XNOR U33562 ( .A(n24878), .B(n24879), .Z(n24864) );
  XOR U33563 ( .A(n24875), .B(n24874), .Z(n24879) );
  XOR U33564 ( .A(y[4776]), .B(x[4776]), .Z(n24874) );
  XOR U33565 ( .A(n24877), .B(n24876), .Z(n24875) );
  XOR U33566 ( .A(y[4778]), .B(x[4778]), .Z(n24876) );
  XOR U33567 ( .A(y[4777]), .B(x[4777]), .Z(n24877) );
  XOR U33568 ( .A(n24869), .B(n24868), .Z(n24878) );
  XOR U33569 ( .A(n24871), .B(n24870), .Z(n24868) );
  XOR U33570 ( .A(y[4775]), .B(x[4775]), .Z(n24870) );
  XOR U33571 ( .A(y[4774]), .B(x[4774]), .Z(n24871) );
  XOR U33572 ( .A(y[4773]), .B(x[4773]), .Z(n24869) );
  XNOR U33573 ( .A(n24862), .B(n24861), .Z(n24863) );
  XNOR U33574 ( .A(n24858), .B(n24857), .Z(n24861) );
  XOR U33575 ( .A(n24860), .B(n24859), .Z(n24857) );
  XOR U33576 ( .A(y[4772]), .B(x[4772]), .Z(n24859) );
  XOR U33577 ( .A(y[4771]), .B(x[4771]), .Z(n24860) );
  XOR U33578 ( .A(y[4770]), .B(x[4770]), .Z(n24858) );
  XOR U33579 ( .A(n24852), .B(n24851), .Z(n24862) );
  XOR U33580 ( .A(n24854), .B(n24853), .Z(n24851) );
  XOR U33581 ( .A(y[4769]), .B(x[4769]), .Z(n24853) );
  XOR U33582 ( .A(y[4768]), .B(x[4768]), .Z(n24854) );
  XOR U33583 ( .A(y[4767]), .B(x[4767]), .Z(n24852) );
  NAND U33584 ( .A(n24915), .B(n24916), .Z(N63170) );
  NAND U33585 ( .A(n24917), .B(n24918), .Z(n24916) );
  NANDN U33586 ( .A(n24919), .B(n24920), .Z(n24918) );
  NANDN U33587 ( .A(n24920), .B(n24919), .Z(n24915) );
  XOR U33588 ( .A(n24919), .B(n24921), .Z(N63169) );
  XNOR U33589 ( .A(n24917), .B(n24920), .Z(n24921) );
  NAND U33590 ( .A(n24922), .B(n24923), .Z(n24920) );
  NAND U33591 ( .A(n24924), .B(n24925), .Z(n24923) );
  NANDN U33592 ( .A(n24926), .B(n24927), .Z(n24925) );
  NANDN U33593 ( .A(n24927), .B(n24926), .Z(n24922) );
  AND U33594 ( .A(n24928), .B(n24929), .Z(n24917) );
  NAND U33595 ( .A(n24930), .B(n24931), .Z(n24929) );
  NANDN U33596 ( .A(n24932), .B(n24933), .Z(n24931) );
  NANDN U33597 ( .A(n24933), .B(n24932), .Z(n24928) );
  IV U33598 ( .A(n24934), .Z(n24933) );
  AND U33599 ( .A(n24935), .B(n24936), .Z(n24919) );
  NAND U33600 ( .A(n24937), .B(n24938), .Z(n24936) );
  NANDN U33601 ( .A(n24939), .B(n24940), .Z(n24938) );
  NANDN U33602 ( .A(n24940), .B(n24939), .Z(n24935) );
  XOR U33603 ( .A(n24932), .B(n24941), .Z(N63168) );
  XNOR U33604 ( .A(n24930), .B(n24934), .Z(n24941) );
  XOR U33605 ( .A(n24927), .B(n24942), .Z(n24934) );
  XNOR U33606 ( .A(n24924), .B(n24926), .Z(n24942) );
  AND U33607 ( .A(n24943), .B(n24944), .Z(n24926) );
  NANDN U33608 ( .A(n24945), .B(n24946), .Z(n24944) );
  OR U33609 ( .A(n24947), .B(n24948), .Z(n24946) );
  IV U33610 ( .A(n24949), .Z(n24948) );
  NANDN U33611 ( .A(n24949), .B(n24947), .Z(n24943) );
  AND U33612 ( .A(n24950), .B(n24951), .Z(n24924) );
  NAND U33613 ( .A(n24952), .B(n24953), .Z(n24951) );
  NANDN U33614 ( .A(n24954), .B(n24955), .Z(n24953) );
  NANDN U33615 ( .A(n24955), .B(n24954), .Z(n24950) );
  IV U33616 ( .A(n24956), .Z(n24955) );
  NAND U33617 ( .A(n24957), .B(n24958), .Z(n24927) );
  NANDN U33618 ( .A(n24959), .B(n24960), .Z(n24958) );
  NANDN U33619 ( .A(n24961), .B(n24962), .Z(n24960) );
  NANDN U33620 ( .A(n24962), .B(n24961), .Z(n24957) );
  IV U33621 ( .A(n24963), .Z(n24961) );
  AND U33622 ( .A(n24964), .B(n24965), .Z(n24930) );
  NAND U33623 ( .A(n24966), .B(n24967), .Z(n24965) );
  NANDN U33624 ( .A(n24968), .B(n24969), .Z(n24967) );
  NANDN U33625 ( .A(n24969), .B(n24968), .Z(n24964) );
  XOR U33626 ( .A(n24940), .B(n24970), .Z(n24932) );
  XNOR U33627 ( .A(n24937), .B(n24939), .Z(n24970) );
  AND U33628 ( .A(n24971), .B(n24972), .Z(n24939) );
  NANDN U33629 ( .A(n24973), .B(n24974), .Z(n24972) );
  OR U33630 ( .A(n24975), .B(n24976), .Z(n24974) );
  IV U33631 ( .A(n24977), .Z(n24976) );
  NANDN U33632 ( .A(n24977), .B(n24975), .Z(n24971) );
  AND U33633 ( .A(n24978), .B(n24979), .Z(n24937) );
  NAND U33634 ( .A(n24980), .B(n24981), .Z(n24979) );
  NANDN U33635 ( .A(n24982), .B(n24983), .Z(n24981) );
  NANDN U33636 ( .A(n24983), .B(n24982), .Z(n24978) );
  IV U33637 ( .A(n24984), .Z(n24983) );
  NAND U33638 ( .A(n24985), .B(n24986), .Z(n24940) );
  NANDN U33639 ( .A(n24987), .B(n24988), .Z(n24986) );
  NANDN U33640 ( .A(n24989), .B(n24990), .Z(n24988) );
  NANDN U33641 ( .A(n24990), .B(n24989), .Z(n24985) );
  IV U33642 ( .A(n24991), .Z(n24989) );
  XOR U33643 ( .A(n24966), .B(n24992), .Z(N63167) );
  XNOR U33644 ( .A(n24969), .B(n24968), .Z(n24992) );
  XNOR U33645 ( .A(n24980), .B(n24993), .Z(n24968) );
  XNOR U33646 ( .A(n24984), .B(n24982), .Z(n24993) );
  XOR U33647 ( .A(n24990), .B(n24994), .Z(n24982) );
  XNOR U33648 ( .A(n24987), .B(n24991), .Z(n24994) );
  AND U33649 ( .A(n24995), .B(n24996), .Z(n24991) );
  NAND U33650 ( .A(n24997), .B(n24998), .Z(n24996) );
  NAND U33651 ( .A(n24999), .B(n25000), .Z(n24995) );
  AND U33652 ( .A(n25001), .B(n25002), .Z(n24987) );
  NAND U33653 ( .A(n25003), .B(n25004), .Z(n25002) );
  NAND U33654 ( .A(n25005), .B(n25006), .Z(n25001) );
  NANDN U33655 ( .A(n25007), .B(n25008), .Z(n24990) );
  ANDN U33656 ( .B(n25009), .A(n25010), .Z(n24984) );
  XNOR U33657 ( .A(n24975), .B(n25011), .Z(n24980) );
  XNOR U33658 ( .A(n24973), .B(n24977), .Z(n25011) );
  AND U33659 ( .A(n25012), .B(n25013), .Z(n24977) );
  NAND U33660 ( .A(n25014), .B(n25015), .Z(n25013) );
  NAND U33661 ( .A(n25016), .B(n25017), .Z(n25012) );
  AND U33662 ( .A(n25018), .B(n25019), .Z(n24973) );
  NAND U33663 ( .A(n25020), .B(n25021), .Z(n25019) );
  NAND U33664 ( .A(n25022), .B(n25023), .Z(n25018) );
  AND U33665 ( .A(n25024), .B(n25025), .Z(n24975) );
  NAND U33666 ( .A(n25026), .B(n25027), .Z(n24969) );
  XNOR U33667 ( .A(n24952), .B(n25028), .Z(n24966) );
  XNOR U33668 ( .A(n24956), .B(n24954), .Z(n25028) );
  XOR U33669 ( .A(n24962), .B(n25029), .Z(n24954) );
  XNOR U33670 ( .A(n24959), .B(n24963), .Z(n25029) );
  AND U33671 ( .A(n25030), .B(n25031), .Z(n24963) );
  NAND U33672 ( .A(n25032), .B(n25033), .Z(n25031) );
  NAND U33673 ( .A(n25034), .B(n25035), .Z(n25030) );
  AND U33674 ( .A(n25036), .B(n25037), .Z(n24959) );
  NAND U33675 ( .A(n25038), .B(n25039), .Z(n25037) );
  NAND U33676 ( .A(n25040), .B(n25041), .Z(n25036) );
  NANDN U33677 ( .A(n25042), .B(n25043), .Z(n24962) );
  ANDN U33678 ( .B(n25044), .A(n25045), .Z(n24956) );
  XNOR U33679 ( .A(n24947), .B(n25046), .Z(n24952) );
  XNOR U33680 ( .A(n24945), .B(n24949), .Z(n25046) );
  AND U33681 ( .A(n25047), .B(n25048), .Z(n24949) );
  NAND U33682 ( .A(n25049), .B(n25050), .Z(n25048) );
  NAND U33683 ( .A(n25051), .B(n25052), .Z(n25047) );
  AND U33684 ( .A(n25053), .B(n25054), .Z(n24945) );
  NAND U33685 ( .A(n25055), .B(n25056), .Z(n25054) );
  NAND U33686 ( .A(n25057), .B(n25058), .Z(n25053) );
  AND U33687 ( .A(n25059), .B(n25060), .Z(n24947) );
  XOR U33688 ( .A(n25027), .B(n25026), .Z(N63166) );
  XNOR U33689 ( .A(n25044), .B(n25045), .Z(n25026) );
  XNOR U33690 ( .A(n25059), .B(n25060), .Z(n25045) );
  XOR U33691 ( .A(n25056), .B(n25055), .Z(n25060) );
  XOR U33692 ( .A(y[4764]), .B(x[4764]), .Z(n25055) );
  XOR U33693 ( .A(n25058), .B(n25057), .Z(n25056) );
  XOR U33694 ( .A(y[4766]), .B(x[4766]), .Z(n25057) );
  XOR U33695 ( .A(y[4765]), .B(x[4765]), .Z(n25058) );
  XOR U33696 ( .A(n25050), .B(n25049), .Z(n25059) );
  XOR U33697 ( .A(n25052), .B(n25051), .Z(n25049) );
  XOR U33698 ( .A(y[4763]), .B(x[4763]), .Z(n25051) );
  XOR U33699 ( .A(y[4762]), .B(x[4762]), .Z(n25052) );
  XOR U33700 ( .A(y[4761]), .B(x[4761]), .Z(n25050) );
  XNOR U33701 ( .A(n25043), .B(n25042), .Z(n25044) );
  XNOR U33702 ( .A(n25039), .B(n25038), .Z(n25042) );
  XOR U33703 ( .A(n25041), .B(n25040), .Z(n25038) );
  XOR U33704 ( .A(y[4760]), .B(x[4760]), .Z(n25040) );
  XOR U33705 ( .A(y[4759]), .B(x[4759]), .Z(n25041) );
  XOR U33706 ( .A(y[4758]), .B(x[4758]), .Z(n25039) );
  XOR U33707 ( .A(n25033), .B(n25032), .Z(n25043) );
  XOR U33708 ( .A(n25035), .B(n25034), .Z(n25032) );
  XOR U33709 ( .A(y[4757]), .B(x[4757]), .Z(n25034) );
  XOR U33710 ( .A(y[4756]), .B(x[4756]), .Z(n25035) );
  XOR U33711 ( .A(y[4755]), .B(x[4755]), .Z(n25033) );
  XNOR U33712 ( .A(n25009), .B(n25010), .Z(n25027) );
  XNOR U33713 ( .A(n25024), .B(n25025), .Z(n25010) );
  XOR U33714 ( .A(n25021), .B(n25020), .Z(n25025) );
  XOR U33715 ( .A(y[4752]), .B(x[4752]), .Z(n25020) );
  XOR U33716 ( .A(n25023), .B(n25022), .Z(n25021) );
  XOR U33717 ( .A(y[4754]), .B(x[4754]), .Z(n25022) );
  XOR U33718 ( .A(y[4753]), .B(x[4753]), .Z(n25023) );
  XOR U33719 ( .A(n25015), .B(n25014), .Z(n25024) );
  XOR U33720 ( .A(n25017), .B(n25016), .Z(n25014) );
  XOR U33721 ( .A(y[4751]), .B(x[4751]), .Z(n25016) );
  XOR U33722 ( .A(y[4750]), .B(x[4750]), .Z(n25017) );
  XOR U33723 ( .A(y[4749]), .B(x[4749]), .Z(n25015) );
  XNOR U33724 ( .A(n25008), .B(n25007), .Z(n25009) );
  XNOR U33725 ( .A(n25004), .B(n25003), .Z(n25007) );
  XOR U33726 ( .A(n25006), .B(n25005), .Z(n25003) );
  XOR U33727 ( .A(y[4748]), .B(x[4748]), .Z(n25005) );
  XOR U33728 ( .A(y[4747]), .B(x[4747]), .Z(n25006) );
  XOR U33729 ( .A(y[4746]), .B(x[4746]), .Z(n25004) );
  XOR U33730 ( .A(n24998), .B(n24997), .Z(n25008) );
  XOR U33731 ( .A(n25000), .B(n24999), .Z(n24997) );
  XOR U33732 ( .A(y[4745]), .B(x[4745]), .Z(n24999) );
  XOR U33733 ( .A(y[4744]), .B(x[4744]), .Z(n25000) );
  XOR U33734 ( .A(y[4743]), .B(x[4743]), .Z(n24998) );
  NAND U33735 ( .A(n25061), .B(n25062), .Z(N63157) );
  NAND U33736 ( .A(n25063), .B(n25064), .Z(n25062) );
  NANDN U33737 ( .A(n25065), .B(n25066), .Z(n25064) );
  NANDN U33738 ( .A(n25066), .B(n25065), .Z(n25061) );
  XOR U33739 ( .A(n25065), .B(n25067), .Z(N63156) );
  XNOR U33740 ( .A(n25063), .B(n25066), .Z(n25067) );
  NAND U33741 ( .A(n25068), .B(n25069), .Z(n25066) );
  NAND U33742 ( .A(n25070), .B(n25071), .Z(n25069) );
  NANDN U33743 ( .A(n25072), .B(n25073), .Z(n25071) );
  NANDN U33744 ( .A(n25073), .B(n25072), .Z(n25068) );
  AND U33745 ( .A(n25074), .B(n25075), .Z(n25063) );
  NAND U33746 ( .A(n25076), .B(n25077), .Z(n25075) );
  NANDN U33747 ( .A(n25078), .B(n25079), .Z(n25077) );
  NANDN U33748 ( .A(n25079), .B(n25078), .Z(n25074) );
  IV U33749 ( .A(n25080), .Z(n25079) );
  AND U33750 ( .A(n25081), .B(n25082), .Z(n25065) );
  NAND U33751 ( .A(n25083), .B(n25084), .Z(n25082) );
  NANDN U33752 ( .A(n25085), .B(n25086), .Z(n25084) );
  NANDN U33753 ( .A(n25086), .B(n25085), .Z(n25081) );
  XOR U33754 ( .A(n25078), .B(n25087), .Z(N63155) );
  XNOR U33755 ( .A(n25076), .B(n25080), .Z(n25087) );
  XOR U33756 ( .A(n25073), .B(n25088), .Z(n25080) );
  XNOR U33757 ( .A(n25070), .B(n25072), .Z(n25088) );
  AND U33758 ( .A(n25089), .B(n25090), .Z(n25072) );
  NANDN U33759 ( .A(n25091), .B(n25092), .Z(n25090) );
  OR U33760 ( .A(n25093), .B(n25094), .Z(n25092) );
  IV U33761 ( .A(n25095), .Z(n25094) );
  NANDN U33762 ( .A(n25095), .B(n25093), .Z(n25089) );
  AND U33763 ( .A(n25096), .B(n25097), .Z(n25070) );
  NAND U33764 ( .A(n25098), .B(n25099), .Z(n25097) );
  NANDN U33765 ( .A(n25100), .B(n25101), .Z(n25099) );
  NANDN U33766 ( .A(n25101), .B(n25100), .Z(n25096) );
  IV U33767 ( .A(n25102), .Z(n25101) );
  NAND U33768 ( .A(n25103), .B(n25104), .Z(n25073) );
  NANDN U33769 ( .A(n25105), .B(n25106), .Z(n25104) );
  NANDN U33770 ( .A(n25107), .B(n25108), .Z(n25106) );
  NANDN U33771 ( .A(n25108), .B(n25107), .Z(n25103) );
  IV U33772 ( .A(n25109), .Z(n25107) );
  AND U33773 ( .A(n25110), .B(n25111), .Z(n25076) );
  NAND U33774 ( .A(n25112), .B(n25113), .Z(n25111) );
  NANDN U33775 ( .A(n25114), .B(n25115), .Z(n25113) );
  NANDN U33776 ( .A(n25115), .B(n25114), .Z(n25110) );
  XOR U33777 ( .A(n25086), .B(n25116), .Z(n25078) );
  XNOR U33778 ( .A(n25083), .B(n25085), .Z(n25116) );
  AND U33779 ( .A(n25117), .B(n25118), .Z(n25085) );
  NANDN U33780 ( .A(n25119), .B(n25120), .Z(n25118) );
  OR U33781 ( .A(n25121), .B(n25122), .Z(n25120) );
  IV U33782 ( .A(n25123), .Z(n25122) );
  NANDN U33783 ( .A(n25123), .B(n25121), .Z(n25117) );
  AND U33784 ( .A(n25124), .B(n25125), .Z(n25083) );
  NAND U33785 ( .A(n25126), .B(n25127), .Z(n25125) );
  NANDN U33786 ( .A(n25128), .B(n25129), .Z(n25127) );
  NANDN U33787 ( .A(n25129), .B(n25128), .Z(n25124) );
  IV U33788 ( .A(n25130), .Z(n25129) );
  NAND U33789 ( .A(n25131), .B(n25132), .Z(n25086) );
  NANDN U33790 ( .A(n25133), .B(n25134), .Z(n25132) );
  NANDN U33791 ( .A(n25135), .B(n25136), .Z(n25134) );
  NANDN U33792 ( .A(n25136), .B(n25135), .Z(n25131) );
  IV U33793 ( .A(n25137), .Z(n25135) );
  XOR U33794 ( .A(n25112), .B(n25138), .Z(N63154) );
  XNOR U33795 ( .A(n25115), .B(n25114), .Z(n25138) );
  XNOR U33796 ( .A(n25126), .B(n25139), .Z(n25114) );
  XNOR U33797 ( .A(n25130), .B(n25128), .Z(n25139) );
  XOR U33798 ( .A(n25136), .B(n25140), .Z(n25128) );
  XNOR U33799 ( .A(n25133), .B(n25137), .Z(n25140) );
  AND U33800 ( .A(n25141), .B(n25142), .Z(n25137) );
  NAND U33801 ( .A(n25143), .B(n25144), .Z(n25142) );
  NAND U33802 ( .A(n25145), .B(n25146), .Z(n25141) );
  AND U33803 ( .A(n25147), .B(n25148), .Z(n25133) );
  NAND U33804 ( .A(n25149), .B(n25150), .Z(n25148) );
  NAND U33805 ( .A(n25151), .B(n25152), .Z(n25147) );
  NANDN U33806 ( .A(n25153), .B(n25154), .Z(n25136) );
  ANDN U33807 ( .B(n25155), .A(n25156), .Z(n25130) );
  XNOR U33808 ( .A(n25121), .B(n25157), .Z(n25126) );
  XNOR U33809 ( .A(n25119), .B(n25123), .Z(n25157) );
  AND U33810 ( .A(n25158), .B(n25159), .Z(n25123) );
  NAND U33811 ( .A(n25160), .B(n25161), .Z(n25159) );
  NAND U33812 ( .A(n25162), .B(n25163), .Z(n25158) );
  AND U33813 ( .A(n25164), .B(n25165), .Z(n25119) );
  NAND U33814 ( .A(n25166), .B(n25167), .Z(n25165) );
  NAND U33815 ( .A(n25168), .B(n25169), .Z(n25164) );
  AND U33816 ( .A(n25170), .B(n25171), .Z(n25121) );
  NAND U33817 ( .A(n25172), .B(n25173), .Z(n25115) );
  XNOR U33818 ( .A(n25098), .B(n25174), .Z(n25112) );
  XNOR U33819 ( .A(n25102), .B(n25100), .Z(n25174) );
  XOR U33820 ( .A(n25108), .B(n25175), .Z(n25100) );
  XNOR U33821 ( .A(n25105), .B(n25109), .Z(n25175) );
  AND U33822 ( .A(n25176), .B(n25177), .Z(n25109) );
  NAND U33823 ( .A(n25178), .B(n25179), .Z(n25177) );
  NAND U33824 ( .A(n25180), .B(n25181), .Z(n25176) );
  AND U33825 ( .A(n25182), .B(n25183), .Z(n25105) );
  NAND U33826 ( .A(n25184), .B(n25185), .Z(n25183) );
  NAND U33827 ( .A(n25186), .B(n25187), .Z(n25182) );
  NANDN U33828 ( .A(n25188), .B(n25189), .Z(n25108) );
  ANDN U33829 ( .B(n25190), .A(n25191), .Z(n25102) );
  XNOR U33830 ( .A(n25093), .B(n25192), .Z(n25098) );
  XNOR U33831 ( .A(n25091), .B(n25095), .Z(n25192) );
  AND U33832 ( .A(n25193), .B(n25194), .Z(n25095) );
  NAND U33833 ( .A(n25195), .B(n25196), .Z(n25194) );
  NAND U33834 ( .A(n25197), .B(n25198), .Z(n25193) );
  AND U33835 ( .A(n25199), .B(n25200), .Z(n25091) );
  NAND U33836 ( .A(n25201), .B(n25202), .Z(n25200) );
  NAND U33837 ( .A(n25203), .B(n25204), .Z(n25199) );
  AND U33838 ( .A(n25205), .B(n25206), .Z(n25093) );
  XOR U33839 ( .A(n25173), .B(n25172), .Z(N63153) );
  XNOR U33840 ( .A(n25190), .B(n25191), .Z(n25172) );
  XNOR U33841 ( .A(n25205), .B(n25206), .Z(n25191) );
  XOR U33842 ( .A(n25202), .B(n25201), .Z(n25206) );
  XOR U33843 ( .A(y[4740]), .B(x[4740]), .Z(n25201) );
  XOR U33844 ( .A(n25204), .B(n25203), .Z(n25202) );
  XOR U33845 ( .A(y[4742]), .B(x[4742]), .Z(n25203) );
  XOR U33846 ( .A(y[4741]), .B(x[4741]), .Z(n25204) );
  XOR U33847 ( .A(n25196), .B(n25195), .Z(n25205) );
  XOR U33848 ( .A(n25198), .B(n25197), .Z(n25195) );
  XOR U33849 ( .A(y[4739]), .B(x[4739]), .Z(n25197) );
  XOR U33850 ( .A(y[4738]), .B(x[4738]), .Z(n25198) );
  XOR U33851 ( .A(y[4737]), .B(x[4737]), .Z(n25196) );
  XNOR U33852 ( .A(n25189), .B(n25188), .Z(n25190) );
  XNOR U33853 ( .A(n25185), .B(n25184), .Z(n25188) );
  XOR U33854 ( .A(n25187), .B(n25186), .Z(n25184) );
  XOR U33855 ( .A(y[4736]), .B(x[4736]), .Z(n25186) );
  XOR U33856 ( .A(y[4735]), .B(x[4735]), .Z(n25187) );
  XOR U33857 ( .A(y[4734]), .B(x[4734]), .Z(n25185) );
  XOR U33858 ( .A(n25179), .B(n25178), .Z(n25189) );
  XOR U33859 ( .A(n25181), .B(n25180), .Z(n25178) );
  XOR U33860 ( .A(y[4733]), .B(x[4733]), .Z(n25180) );
  XOR U33861 ( .A(y[4732]), .B(x[4732]), .Z(n25181) );
  XOR U33862 ( .A(y[4731]), .B(x[4731]), .Z(n25179) );
  XNOR U33863 ( .A(n25155), .B(n25156), .Z(n25173) );
  XNOR U33864 ( .A(n25170), .B(n25171), .Z(n25156) );
  XOR U33865 ( .A(n25167), .B(n25166), .Z(n25171) );
  XOR U33866 ( .A(y[4728]), .B(x[4728]), .Z(n25166) );
  XOR U33867 ( .A(n25169), .B(n25168), .Z(n25167) );
  XOR U33868 ( .A(y[4730]), .B(x[4730]), .Z(n25168) );
  XOR U33869 ( .A(y[4729]), .B(x[4729]), .Z(n25169) );
  XOR U33870 ( .A(n25161), .B(n25160), .Z(n25170) );
  XOR U33871 ( .A(n25163), .B(n25162), .Z(n25160) );
  XOR U33872 ( .A(y[4727]), .B(x[4727]), .Z(n25162) );
  XOR U33873 ( .A(y[4726]), .B(x[4726]), .Z(n25163) );
  XOR U33874 ( .A(y[4725]), .B(x[4725]), .Z(n25161) );
  XNOR U33875 ( .A(n25154), .B(n25153), .Z(n25155) );
  XNOR U33876 ( .A(n25150), .B(n25149), .Z(n25153) );
  XOR U33877 ( .A(n25152), .B(n25151), .Z(n25149) );
  XOR U33878 ( .A(y[4724]), .B(x[4724]), .Z(n25151) );
  XOR U33879 ( .A(y[4723]), .B(x[4723]), .Z(n25152) );
  XOR U33880 ( .A(y[4722]), .B(x[4722]), .Z(n25150) );
  XOR U33881 ( .A(n25144), .B(n25143), .Z(n25154) );
  XOR U33882 ( .A(n25146), .B(n25145), .Z(n25143) );
  XOR U33883 ( .A(y[4721]), .B(x[4721]), .Z(n25145) );
  XOR U33884 ( .A(y[4720]), .B(x[4720]), .Z(n25146) );
  XOR U33885 ( .A(y[4719]), .B(x[4719]), .Z(n25144) );
  NAND U33886 ( .A(n25207), .B(n25208), .Z(N63144) );
  NAND U33887 ( .A(n25209), .B(n25210), .Z(n25208) );
  NANDN U33888 ( .A(n25211), .B(n25212), .Z(n25210) );
  NANDN U33889 ( .A(n25212), .B(n25211), .Z(n25207) );
  XOR U33890 ( .A(n25211), .B(n25213), .Z(N63143) );
  XNOR U33891 ( .A(n25209), .B(n25212), .Z(n25213) );
  NAND U33892 ( .A(n25214), .B(n25215), .Z(n25212) );
  NAND U33893 ( .A(n25216), .B(n25217), .Z(n25215) );
  NANDN U33894 ( .A(n25218), .B(n25219), .Z(n25217) );
  NANDN U33895 ( .A(n25219), .B(n25218), .Z(n25214) );
  AND U33896 ( .A(n25220), .B(n25221), .Z(n25209) );
  NAND U33897 ( .A(n25222), .B(n25223), .Z(n25221) );
  NANDN U33898 ( .A(n25224), .B(n25225), .Z(n25223) );
  NANDN U33899 ( .A(n25225), .B(n25224), .Z(n25220) );
  IV U33900 ( .A(n25226), .Z(n25225) );
  AND U33901 ( .A(n25227), .B(n25228), .Z(n25211) );
  NAND U33902 ( .A(n25229), .B(n25230), .Z(n25228) );
  NANDN U33903 ( .A(n25231), .B(n25232), .Z(n25230) );
  NANDN U33904 ( .A(n25232), .B(n25231), .Z(n25227) );
  XOR U33905 ( .A(n25224), .B(n25233), .Z(N63142) );
  XNOR U33906 ( .A(n25222), .B(n25226), .Z(n25233) );
  XOR U33907 ( .A(n25219), .B(n25234), .Z(n25226) );
  XNOR U33908 ( .A(n25216), .B(n25218), .Z(n25234) );
  AND U33909 ( .A(n25235), .B(n25236), .Z(n25218) );
  NANDN U33910 ( .A(n25237), .B(n25238), .Z(n25236) );
  OR U33911 ( .A(n25239), .B(n25240), .Z(n25238) );
  IV U33912 ( .A(n25241), .Z(n25240) );
  NANDN U33913 ( .A(n25241), .B(n25239), .Z(n25235) );
  AND U33914 ( .A(n25242), .B(n25243), .Z(n25216) );
  NAND U33915 ( .A(n25244), .B(n25245), .Z(n25243) );
  NANDN U33916 ( .A(n25246), .B(n25247), .Z(n25245) );
  NANDN U33917 ( .A(n25247), .B(n25246), .Z(n25242) );
  IV U33918 ( .A(n25248), .Z(n25247) );
  NAND U33919 ( .A(n25249), .B(n25250), .Z(n25219) );
  NANDN U33920 ( .A(n25251), .B(n25252), .Z(n25250) );
  NANDN U33921 ( .A(n25253), .B(n25254), .Z(n25252) );
  NANDN U33922 ( .A(n25254), .B(n25253), .Z(n25249) );
  IV U33923 ( .A(n25255), .Z(n25253) );
  AND U33924 ( .A(n25256), .B(n25257), .Z(n25222) );
  NAND U33925 ( .A(n25258), .B(n25259), .Z(n25257) );
  NANDN U33926 ( .A(n25260), .B(n25261), .Z(n25259) );
  NANDN U33927 ( .A(n25261), .B(n25260), .Z(n25256) );
  XOR U33928 ( .A(n25232), .B(n25262), .Z(n25224) );
  XNOR U33929 ( .A(n25229), .B(n25231), .Z(n25262) );
  AND U33930 ( .A(n25263), .B(n25264), .Z(n25231) );
  NANDN U33931 ( .A(n25265), .B(n25266), .Z(n25264) );
  OR U33932 ( .A(n25267), .B(n25268), .Z(n25266) );
  IV U33933 ( .A(n25269), .Z(n25268) );
  NANDN U33934 ( .A(n25269), .B(n25267), .Z(n25263) );
  AND U33935 ( .A(n25270), .B(n25271), .Z(n25229) );
  NAND U33936 ( .A(n25272), .B(n25273), .Z(n25271) );
  NANDN U33937 ( .A(n25274), .B(n25275), .Z(n25273) );
  NANDN U33938 ( .A(n25275), .B(n25274), .Z(n25270) );
  IV U33939 ( .A(n25276), .Z(n25275) );
  NAND U33940 ( .A(n25277), .B(n25278), .Z(n25232) );
  NANDN U33941 ( .A(n25279), .B(n25280), .Z(n25278) );
  NANDN U33942 ( .A(n25281), .B(n25282), .Z(n25280) );
  NANDN U33943 ( .A(n25282), .B(n25281), .Z(n25277) );
  IV U33944 ( .A(n25283), .Z(n25281) );
  XOR U33945 ( .A(n25258), .B(n25284), .Z(N63141) );
  XNOR U33946 ( .A(n25261), .B(n25260), .Z(n25284) );
  XNOR U33947 ( .A(n25272), .B(n25285), .Z(n25260) );
  XNOR U33948 ( .A(n25276), .B(n25274), .Z(n25285) );
  XOR U33949 ( .A(n25282), .B(n25286), .Z(n25274) );
  XNOR U33950 ( .A(n25279), .B(n25283), .Z(n25286) );
  AND U33951 ( .A(n25287), .B(n25288), .Z(n25283) );
  NAND U33952 ( .A(n25289), .B(n25290), .Z(n25288) );
  NAND U33953 ( .A(n25291), .B(n25292), .Z(n25287) );
  AND U33954 ( .A(n25293), .B(n25294), .Z(n25279) );
  NAND U33955 ( .A(n25295), .B(n25296), .Z(n25294) );
  NAND U33956 ( .A(n25297), .B(n25298), .Z(n25293) );
  NANDN U33957 ( .A(n25299), .B(n25300), .Z(n25282) );
  ANDN U33958 ( .B(n25301), .A(n25302), .Z(n25276) );
  XNOR U33959 ( .A(n25267), .B(n25303), .Z(n25272) );
  XNOR U33960 ( .A(n25265), .B(n25269), .Z(n25303) );
  AND U33961 ( .A(n25304), .B(n25305), .Z(n25269) );
  NAND U33962 ( .A(n25306), .B(n25307), .Z(n25305) );
  NAND U33963 ( .A(n25308), .B(n25309), .Z(n25304) );
  AND U33964 ( .A(n25310), .B(n25311), .Z(n25265) );
  NAND U33965 ( .A(n25312), .B(n25313), .Z(n25311) );
  NAND U33966 ( .A(n25314), .B(n25315), .Z(n25310) );
  AND U33967 ( .A(n25316), .B(n25317), .Z(n25267) );
  NAND U33968 ( .A(n25318), .B(n25319), .Z(n25261) );
  XNOR U33969 ( .A(n25244), .B(n25320), .Z(n25258) );
  XNOR U33970 ( .A(n25248), .B(n25246), .Z(n25320) );
  XOR U33971 ( .A(n25254), .B(n25321), .Z(n25246) );
  XNOR U33972 ( .A(n25251), .B(n25255), .Z(n25321) );
  AND U33973 ( .A(n25322), .B(n25323), .Z(n25255) );
  NAND U33974 ( .A(n25324), .B(n25325), .Z(n25323) );
  NAND U33975 ( .A(n25326), .B(n25327), .Z(n25322) );
  AND U33976 ( .A(n25328), .B(n25329), .Z(n25251) );
  NAND U33977 ( .A(n25330), .B(n25331), .Z(n25329) );
  NAND U33978 ( .A(n25332), .B(n25333), .Z(n25328) );
  NANDN U33979 ( .A(n25334), .B(n25335), .Z(n25254) );
  ANDN U33980 ( .B(n25336), .A(n25337), .Z(n25248) );
  XNOR U33981 ( .A(n25239), .B(n25338), .Z(n25244) );
  XNOR U33982 ( .A(n25237), .B(n25241), .Z(n25338) );
  AND U33983 ( .A(n25339), .B(n25340), .Z(n25241) );
  NAND U33984 ( .A(n25341), .B(n25342), .Z(n25340) );
  NAND U33985 ( .A(n25343), .B(n25344), .Z(n25339) );
  AND U33986 ( .A(n25345), .B(n25346), .Z(n25237) );
  NAND U33987 ( .A(n25347), .B(n25348), .Z(n25346) );
  NAND U33988 ( .A(n25349), .B(n25350), .Z(n25345) );
  AND U33989 ( .A(n25351), .B(n25352), .Z(n25239) );
  XOR U33990 ( .A(n25319), .B(n25318), .Z(N63140) );
  XNOR U33991 ( .A(n25336), .B(n25337), .Z(n25318) );
  XNOR U33992 ( .A(n25351), .B(n25352), .Z(n25337) );
  XOR U33993 ( .A(n25348), .B(n25347), .Z(n25352) );
  XOR U33994 ( .A(y[4716]), .B(x[4716]), .Z(n25347) );
  XOR U33995 ( .A(n25350), .B(n25349), .Z(n25348) );
  XOR U33996 ( .A(y[4718]), .B(x[4718]), .Z(n25349) );
  XOR U33997 ( .A(y[4717]), .B(x[4717]), .Z(n25350) );
  XOR U33998 ( .A(n25342), .B(n25341), .Z(n25351) );
  XOR U33999 ( .A(n25344), .B(n25343), .Z(n25341) );
  XOR U34000 ( .A(y[4715]), .B(x[4715]), .Z(n25343) );
  XOR U34001 ( .A(y[4714]), .B(x[4714]), .Z(n25344) );
  XOR U34002 ( .A(y[4713]), .B(x[4713]), .Z(n25342) );
  XNOR U34003 ( .A(n25335), .B(n25334), .Z(n25336) );
  XNOR U34004 ( .A(n25331), .B(n25330), .Z(n25334) );
  XOR U34005 ( .A(n25333), .B(n25332), .Z(n25330) );
  XOR U34006 ( .A(y[4712]), .B(x[4712]), .Z(n25332) );
  XOR U34007 ( .A(y[4711]), .B(x[4711]), .Z(n25333) );
  XOR U34008 ( .A(y[4710]), .B(x[4710]), .Z(n25331) );
  XOR U34009 ( .A(n25325), .B(n25324), .Z(n25335) );
  XOR U34010 ( .A(n25327), .B(n25326), .Z(n25324) );
  XOR U34011 ( .A(y[4709]), .B(x[4709]), .Z(n25326) );
  XOR U34012 ( .A(y[4708]), .B(x[4708]), .Z(n25327) );
  XOR U34013 ( .A(y[4707]), .B(x[4707]), .Z(n25325) );
  XNOR U34014 ( .A(n25301), .B(n25302), .Z(n25319) );
  XNOR U34015 ( .A(n25316), .B(n25317), .Z(n25302) );
  XOR U34016 ( .A(n25313), .B(n25312), .Z(n25317) );
  XOR U34017 ( .A(y[4704]), .B(x[4704]), .Z(n25312) );
  XOR U34018 ( .A(n25315), .B(n25314), .Z(n25313) );
  XOR U34019 ( .A(y[4706]), .B(x[4706]), .Z(n25314) );
  XOR U34020 ( .A(y[4705]), .B(x[4705]), .Z(n25315) );
  XOR U34021 ( .A(n25307), .B(n25306), .Z(n25316) );
  XOR U34022 ( .A(n25309), .B(n25308), .Z(n25306) );
  XOR U34023 ( .A(y[4703]), .B(x[4703]), .Z(n25308) );
  XOR U34024 ( .A(y[4702]), .B(x[4702]), .Z(n25309) );
  XOR U34025 ( .A(y[4701]), .B(x[4701]), .Z(n25307) );
  XNOR U34026 ( .A(n25300), .B(n25299), .Z(n25301) );
  XNOR U34027 ( .A(n25296), .B(n25295), .Z(n25299) );
  XOR U34028 ( .A(n25298), .B(n25297), .Z(n25295) );
  XOR U34029 ( .A(y[4700]), .B(x[4700]), .Z(n25297) );
  XOR U34030 ( .A(y[4699]), .B(x[4699]), .Z(n25298) );
  XOR U34031 ( .A(y[4698]), .B(x[4698]), .Z(n25296) );
  XOR U34032 ( .A(n25290), .B(n25289), .Z(n25300) );
  XOR U34033 ( .A(n25292), .B(n25291), .Z(n25289) );
  XOR U34034 ( .A(y[4697]), .B(x[4697]), .Z(n25291) );
  XOR U34035 ( .A(y[4696]), .B(x[4696]), .Z(n25292) );
  XOR U34036 ( .A(y[4695]), .B(x[4695]), .Z(n25290) );
  NAND U34037 ( .A(n25353), .B(n25354), .Z(N63131) );
  NAND U34038 ( .A(n25355), .B(n25356), .Z(n25354) );
  NANDN U34039 ( .A(n25357), .B(n25358), .Z(n25356) );
  NANDN U34040 ( .A(n25358), .B(n25357), .Z(n25353) );
  XOR U34041 ( .A(n25357), .B(n25359), .Z(N63130) );
  XNOR U34042 ( .A(n25355), .B(n25358), .Z(n25359) );
  NAND U34043 ( .A(n25360), .B(n25361), .Z(n25358) );
  NAND U34044 ( .A(n25362), .B(n25363), .Z(n25361) );
  NANDN U34045 ( .A(n25364), .B(n25365), .Z(n25363) );
  NANDN U34046 ( .A(n25365), .B(n25364), .Z(n25360) );
  AND U34047 ( .A(n25366), .B(n25367), .Z(n25355) );
  NAND U34048 ( .A(n25368), .B(n25369), .Z(n25367) );
  NANDN U34049 ( .A(n25370), .B(n25371), .Z(n25369) );
  NANDN U34050 ( .A(n25371), .B(n25370), .Z(n25366) );
  IV U34051 ( .A(n25372), .Z(n25371) );
  AND U34052 ( .A(n25373), .B(n25374), .Z(n25357) );
  NAND U34053 ( .A(n25375), .B(n25376), .Z(n25374) );
  NANDN U34054 ( .A(n25377), .B(n25378), .Z(n25376) );
  NANDN U34055 ( .A(n25378), .B(n25377), .Z(n25373) );
  XOR U34056 ( .A(n25370), .B(n25379), .Z(N63129) );
  XNOR U34057 ( .A(n25368), .B(n25372), .Z(n25379) );
  XOR U34058 ( .A(n25365), .B(n25380), .Z(n25372) );
  XNOR U34059 ( .A(n25362), .B(n25364), .Z(n25380) );
  AND U34060 ( .A(n25381), .B(n25382), .Z(n25364) );
  NANDN U34061 ( .A(n25383), .B(n25384), .Z(n25382) );
  OR U34062 ( .A(n25385), .B(n25386), .Z(n25384) );
  IV U34063 ( .A(n25387), .Z(n25386) );
  NANDN U34064 ( .A(n25387), .B(n25385), .Z(n25381) );
  AND U34065 ( .A(n25388), .B(n25389), .Z(n25362) );
  NAND U34066 ( .A(n25390), .B(n25391), .Z(n25389) );
  NANDN U34067 ( .A(n25392), .B(n25393), .Z(n25391) );
  NANDN U34068 ( .A(n25393), .B(n25392), .Z(n25388) );
  IV U34069 ( .A(n25394), .Z(n25393) );
  NAND U34070 ( .A(n25395), .B(n25396), .Z(n25365) );
  NANDN U34071 ( .A(n25397), .B(n25398), .Z(n25396) );
  NANDN U34072 ( .A(n25399), .B(n25400), .Z(n25398) );
  NANDN U34073 ( .A(n25400), .B(n25399), .Z(n25395) );
  IV U34074 ( .A(n25401), .Z(n25399) );
  AND U34075 ( .A(n25402), .B(n25403), .Z(n25368) );
  NAND U34076 ( .A(n25404), .B(n25405), .Z(n25403) );
  NANDN U34077 ( .A(n25406), .B(n25407), .Z(n25405) );
  NANDN U34078 ( .A(n25407), .B(n25406), .Z(n25402) );
  XOR U34079 ( .A(n25378), .B(n25408), .Z(n25370) );
  XNOR U34080 ( .A(n25375), .B(n25377), .Z(n25408) );
  AND U34081 ( .A(n25409), .B(n25410), .Z(n25377) );
  NANDN U34082 ( .A(n25411), .B(n25412), .Z(n25410) );
  OR U34083 ( .A(n25413), .B(n25414), .Z(n25412) );
  IV U34084 ( .A(n25415), .Z(n25414) );
  NANDN U34085 ( .A(n25415), .B(n25413), .Z(n25409) );
  AND U34086 ( .A(n25416), .B(n25417), .Z(n25375) );
  NAND U34087 ( .A(n25418), .B(n25419), .Z(n25417) );
  NANDN U34088 ( .A(n25420), .B(n25421), .Z(n25419) );
  NANDN U34089 ( .A(n25421), .B(n25420), .Z(n25416) );
  IV U34090 ( .A(n25422), .Z(n25421) );
  NAND U34091 ( .A(n25423), .B(n25424), .Z(n25378) );
  NANDN U34092 ( .A(n25425), .B(n25426), .Z(n25424) );
  NANDN U34093 ( .A(n25427), .B(n25428), .Z(n25426) );
  NANDN U34094 ( .A(n25428), .B(n25427), .Z(n25423) );
  IV U34095 ( .A(n25429), .Z(n25427) );
  XOR U34096 ( .A(n25404), .B(n25430), .Z(N63128) );
  XNOR U34097 ( .A(n25407), .B(n25406), .Z(n25430) );
  XNOR U34098 ( .A(n25418), .B(n25431), .Z(n25406) );
  XNOR U34099 ( .A(n25422), .B(n25420), .Z(n25431) );
  XOR U34100 ( .A(n25428), .B(n25432), .Z(n25420) );
  XNOR U34101 ( .A(n25425), .B(n25429), .Z(n25432) );
  AND U34102 ( .A(n25433), .B(n25434), .Z(n25429) );
  NAND U34103 ( .A(n25435), .B(n25436), .Z(n25434) );
  NAND U34104 ( .A(n25437), .B(n25438), .Z(n25433) );
  AND U34105 ( .A(n25439), .B(n25440), .Z(n25425) );
  NAND U34106 ( .A(n25441), .B(n25442), .Z(n25440) );
  NAND U34107 ( .A(n25443), .B(n25444), .Z(n25439) );
  NANDN U34108 ( .A(n25445), .B(n25446), .Z(n25428) );
  ANDN U34109 ( .B(n25447), .A(n25448), .Z(n25422) );
  XNOR U34110 ( .A(n25413), .B(n25449), .Z(n25418) );
  XNOR U34111 ( .A(n25411), .B(n25415), .Z(n25449) );
  AND U34112 ( .A(n25450), .B(n25451), .Z(n25415) );
  NAND U34113 ( .A(n25452), .B(n25453), .Z(n25451) );
  NAND U34114 ( .A(n25454), .B(n25455), .Z(n25450) );
  AND U34115 ( .A(n25456), .B(n25457), .Z(n25411) );
  NAND U34116 ( .A(n25458), .B(n25459), .Z(n25457) );
  NAND U34117 ( .A(n25460), .B(n25461), .Z(n25456) );
  AND U34118 ( .A(n25462), .B(n25463), .Z(n25413) );
  NAND U34119 ( .A(n25464), .B(n25465), .Z(n25407) );
  XNOR U34120 ( .A(n25390), .B(n25466), .Z(n25404) );
  XNOR U34121 ( .A(n25394), .B(n25392), .Z(n25466) );
  XOR U34122 ( .A(n25400), .B(n25467), .Z(n25392) );
  XNOR U34123 ( .A(n25397), .B(n25401), .Z(n25467) );
  AND U34124 ( .A(n25468), .B(n25469), .Z(n25401) );
  NAND U34125 ( .A(n25470), .B(n25471), .Z(n25469) );
  NAND U34126 ( .A(n25472), .B(n25473), .Z(n25468) );
  AND U34127 ( .A(n25474), .B(n25475), .Z(n25397) );
  NAND U34128 ( .A(n25476), .B(n25477), .Z(n25475) );
  NAND U34129 ( .A(n25478), .B(n25479), .Z(n25474) );
  NANDN U34130 ( .A(n25480), .B(n25481), .Z(n25400) );
  ANDN U34131 ( .B(n25482), .A(n25483), .Z(n25394) );
  XNOR U34132 ( .A(n25385), .B(n25484), .Z(n25390) );
  XNOR U34133 ( .A(n25383), .B(n25387), .Z(n25484) );
  AND U34134 ( .A(n25485), .B(n25486), .Z(n25387) );
  NAND U34135 ( .A(n25487), .B(n25488), .Z(n25486) );
  NAND U34136 ( .A(n25489), .B(n25490), .Z(n25485) );
  AND U34137 ( .A(n25491), .B(n25492), .Z(n25383) );
  NAND U34138 ( .A(n25493), .B(n25494), .Z(n25492) );
  NAND U34139 ( .A(n25495), .B(n25496), .Z(n25491) );
  AND U34140 ( .A(n25497), .B(n25498), .Z(n25385) );
  XOR U34141 ( .A(n25465), .B(n25464), .Z(N63127) );
  XNOR U34142 ( .A(n25482), .B(n25483), .Z(n25464) );
  XNOR U34143 ( .A(n25497), .B(n25498), .Z(n25483) );
  XOR U34144 ( .A(n25494), .B(n25493), .Z(n25498) );
  XOR U34145 ( .A(y[4692]), .B(x[4692]), .Z(n25493) );
  XOR U34146 ( .A(n25496), .B(n25495), .Z(n25494) );
  XOR U34147 ( .A(y[4694]), .B(x[4694]), .Z(n25495) );
  XOR U34148 ( .A(y[4693]), .B(x[4693]), .Z(n25496) );
  XOR U34149 ( .A(n25488), .B(n25487), .Z(n25497) );
  XOR U34150 ( .A(n25490), .B(n25489), .Z(n25487) );
  XOR U34151 ( .A(y[4691]), .B(x[4691]), .Z(n25489) );
  XOR U34152 ( .A(y[4690]), .B(x[4690]), .Z(n25490) );
  XOR U34153 ( .A(y[4689]), .B(x[4689]), .Z(n25488) );
  XNOR U34154 ( .A(n25481), .B(n25480), .Z(n25482) );
  XNOR U34155 ( .A(n25477), .B(n25476), .Z(n25480) );
  XOR U34156 ( .A(n25479), .B(n25478), .Z(n25476) );
  XOR U34157 ( .A(y[4688]), .B(x[4688]), .Z(n25478) );
  XOR U34158 ( .A(y[4687]), .B(x[4687]), .Z(n25479) );
  XOR U34159 ( .A(y[4686]), .B(x[4686]), .Z(n25477) );
  XOR U34160 ( .A(n25471), .B(n25470), .Z(n25481) );
  XOR U34161 ( .A(n25473), .B(n25472), .Z(n25470) );
  XOR U34162 ( .A(y[4685]), .B(x[4685]), .Z(n25472) );
  XOR U34163 ( .A(y[4684]), .B(x[4684]), .Z(n25473) );
  XOR U34164 ( .A(y[4683]), .B(x[4683]), .Z(n25471) );
  XNOR U34165 ( .A(n25447), .B(n25448), .Z(n25465) );
  XNOR U34166 ( .A(n25462), .B(n25463), .Z(n25448) );
  XOR U34167 ( .A(n25459), .B(n25458), .Z(n25463) );
  XOR U34168 ( .A(y[4680]), .B(x[4680]), .Z(n25458) );
  XOR U34169 ( .A(n25461), .B(n25460), .Z(n25459) );
  XOR U34170 ( .A(y[4682]), .B(x[4682]), .Z(n25460) );
  XOR U34171 ( .A(y[4681]), .B(x[4681]), .Z(n25461) );
  XOR U34172 ( .A(n25453), .B(n25452), .Z(n25462) );
  XOR U34173 ( .A(n25455), .B(n25454), .Z(n25452) );
  XOR U34174 ( .A(y[4679]), .B(x[4679]), .Z(n25454) );
  XOR U34175 ( .A(y[4678]), .B(x[4678]), .Z(n25455) );
  XOR U34176 ( .A(y[4677]), .B(x[4677]), .Z(n25453) );
  XNOR U34177 ( .A(n25446), .B(n25445), .Z(n25447) );
  XNOR U34178 ( .A(n25442), .B(n25441), .Z(n25445) );
  XOR U34179 ( .A(n25444), .B(n25443), .Z(n25441) );
  XOR U34180 ( .A(y[4676]), .B(x[4676]), .Z(n25443) );
  XOR U34181 ( .A(y[4675]), .B(x[4675]), .Z(n25444) );
  XOR U34182 ( .A(y[4674]), .B(x[4674]), .Z(n25442) );
  XOR U34183 ( .A(n25436), .B(n25435), .Z(n25446) );
  XOR U34184 ( .A(n25438), .B(n25437), .Z(n25435) );
  XOR U34185 ( .A(y[4673]), .B(x[4673]), .Z(n25437) );
  XOR U34186 ( .A(y[4672]), .B(x[4672]), .Z(n25438) );
  XOR U34187 ( .A(y[4671]), .B(x[4671]), .Z(n25436) );
  NAND U34188 ( .A(n25499), .B(n25500), .Z(N63118) );
  NAND U34189 ( .A(n25501), .B(n25502), .Z(n25500) );
  NANDN U34190 ( .A(n25503), .B(n25504), .Z(n25502) );
  NANDN U34191 ( .A(n25504), .B(n25503), .Z(n25499) );
  XOR U34192 ( .A(n25503), .B(n25505), .Z(N63117) );
  XNOR U34193 ( .A(n25501), .B(n25504), .Z(n25505) );
  NAND U34194 ( .A(n25506), .B(n25507), .Z(n25504) );
  NAND U34195 ( .A(n25508), .B(n25509), .Z(n25507) );
  NANDN U34196 ( .A(n25510), .B(n25511), .Z(n25509) );
  NANDN U34197 ( .A(n25511), .B(n25510), .Z(n25506) );
  AND U34198 ( .A(n25512), .B(n25513), .Z(n25501) );
  NAND U34199 ( .A(n25514), .B(n25515), .Z(n25513) );
  NANDN U34200 ( .A(n25516), .B(n25517), .Z(n25515) );
  NANDN U34201 ( .A(n25517), .B(n25516), .Z(n25512) );
  IV U34202 ( .A(n25518), .Z(n25517) );
  AND U34203 ( .A(n25519), .B(n25520), .Z(n25503) );
  NAND U34204 ( .A(n25521), .B(n25522), .Z(n25520) );
  NANDN U34205 ( .A(n25523), .B(n25524), .Z(n25522) );
  NANDN U34206 ( .A(n25524), .B(n25523), .Z(n25519) );
  XOR U34207 ( .A(n25516), .B(n25525), .Z(N63116) );
  XNOR U34208 ( .A(n25514), .B(n25518), .Z(n25525) );
  XOR U34209 ( .A(n25511), .B(n25526), .Z(n25518) );
  XNOR U34210 ( .A(n25508), .B(n25510), .Z(n25526) );
  AND U34211 ( .A(n25527), .B(n25528), .Z(n25510) );
  NANDN U34212 ( .A(n25529), .B(n25530), .Z(n25528) );
  OR U34213 ( .A(n25531), .B(n25532), .Z(n25530) );
  IV U34214 ( .A(n25533), .Z(n25532) );
  NANDN U34215 ( .A(n25533), .B(n25531), .Z(n25527) );
  AND U34216 ( .A(n25534), .B(n25535), .Z(n25508) );
  NAND U34217 ( .A(n25536), .B(n25537), .Z(n25535) );
  NANDN U34218 ( .A(n25538), .B(n25539), .Z(n25537) );
  NANDN U34219 ( .A(n25539), .B(n25538), .Z(n25534) );
  IV U34220 ( .A(n25540), .Z(n25539) );
  NAND U34221 ( .A(n25541), .B(n25542), .Z(n25511) );
  NANDN U34222 ( .A(n25543), .B(n25544), .Z(n25542) );
  NANDN U34223 ( .A(n25545), .B(n25546), .Z(n25544) );
  NANDN U34224 ( .A(n25546), .B(n25545), .Z(n25541) );
  IV U34225 ( .A(n25547), .Z(n25545) );
  AND U34226 ( .A(n25548), .B(n25549), .Z(n25514) );
  NAND U34227 ( .A(n25550), .B(n25551), .Z(n25549) );
  NANDN U34228 ( .A(n25552), .B(n25553), .Z(n25551) );
  NANDN U34229 ( .A(n25553), .B(n25552), .Z(n25548) );
  XOR U34230 ( .A(n25524), .B(n25554), .Z(n25516) );
  XNOR U34231 ( .A(n25521), .B(n25523), .Z(n25554) );
  AND U34232 ( .A(n25555), .B(n25556), .Z(n25523) );
  NANDN U34233 ( .A(n25557), .B(n25558), .Z(n25556) );
  OR U34234 ( .A(n25559), .B(n25560), .Z(n25558) );
  IV U34235 ( .A(n25561), .Z(n25560) );
  NANDN U34236 ( .A(n25561), .B(n25559), .Z(n25555) );
  AND U34237 ( .A(n25562), .B(n25563), .Z(n25521) );
  NAND U34238 ( .A(n25564), .B(n25565), .Z(n25563) );
  NANDN U34239 ( .A(n25566), .B(n25567), .Z(n25565) );
  NANDN U34240 ( .A(n25567), .B(n25566), .Z(n25562) );
  IV U34241 ( .A(n25568), .Z(n25567) );
  NAND U34242 ( .A(n25569), .B(n25570), .Z(n25524) );
  NANDN U34243 ( .A(n25571), .B(n25572), .Z(n25570) );
  NANDN U34244 ( .A(n25573), .B(n25574), .Z(n25572) );
  NANDN U34245 ( .A(n25574), .B(n25573), .Z(n25569) );
  IV U34246 ( .A(n25575), .Z(n25573) );
  XOR U34247 ( .A(n25550), .B(n25576), .Z(N63115) );
  XNOR U34248 ( .A(n25553), .B(n25552), .Z(n25576) );
  XNOR U34249 ( .A(n25564), .B(n25577), .Z(n25552) );
  XNOR U34250 ( .A(n25568), .B(n25566), .Z(n25577) );
  XOR U34251 ( .A(n25574), .B(n25578), .Z(n25566) );
  XNOR U34252 ( .A(n25571), .B(n25575), .Z(n25578) );
  AND U34253 ( .A(n25579), .B(n25580), .Z(n25575) );
  NAND U34254 ( .A(n25581), .B(n25582), .Z(n25580) );
  NAND U34255 ( .A(n25583), .B(n25584), .Z(n25579) );
  AND U34256 ( .A(n25585), .B(n25586), .Z(n25571) );
  NAND U34257 ( .A(n25587), .B(n25588), .Z(n25586) );
  NAND U34258 ( .A(n25589), .B(n25590), .Z(n25585) );
  NANDN U34259 ( .A(n25591), .B(n25592), .Z(n25574) );
  ANDN U34260 ( .B(n25593), .A(n25594), .Z(n25568) );
  XNOR U34261 ( .A(n25559), .B(n25595), .Z(n25564) );
  XNOR U34262 ( .A(n25557), .B(n25561), .Z(n25595) );
  AND U34263 ( .A(n25596), .B(n25597), .Z(n25561) );
  NAND U34264 ( .A(n25598), .B(n25599), .Z(n25597) );
  NAND U34265 ( .A(n25600), .B(n25601), .Z(n25596) );
  AND U34266 ( .A(n25602), .B(n25603), .Z(n25557) );
  NAND U34267 ( .A(n25604), .B(n25605), .Z(n25603) );
  NAND U34268 ( .A(n25606), .B(n25607), .Z(n25602) );
  AND U34269 ( .A(n25608), .B(n25609), .Z(n25559) );
  NAND U34270 ( .A(n25610), .B(n25611), .Z(n25553) );
  XNOR U34271 ( .A(n25536), .B(n25612), .Z(n25550) );
  XNOR U34272 ( .A(n25540), .B(n25538), .Z(n25612) );
  XOR U34273 ( .A(n25546), .B(n25613), .Z(n25538) );
  XNOR U34274 ( .A(n25543), .B(n25547), .Z(n25613) );
  AND U34275 ( .A(n25614), .B(n25615), .Z(n25547) );
  NAND U34276 ( .A(n25616), .B(n25617), .Z(n25615) );
  NAND U34277 ( .A(n25618), .B(n25619), .Z(n25614) );
  AND U34278 ( .A(n25620), .B(n25621), .Z(n25543) );
  NAND U34279 ( .A(n25622), .B(n25623), .Z(n25621) );
  NAND U34280 ( .A(n25624), .B(n25625), .Z(n25620) );
  NANDN U34281 ( .A(n25626), .B(n25627), .Z(n25546) );
  ANDN U34282 ( .B(n25628), .A(n25629), .Z(n25540) );
  XNOR U34283 ( .A(n25531), .B(n25630), .Z(n25536) );
  XNOR U34284 ( .A(n25529), .B(n25533), .Z(n25630) );
  AND U34285 ( .A(n25631), .B(n25632), .Z(n25533) );
  NAND U34286 ( .A(n25633), .B(n25634), .Z(n25632) );
  NAND U34287 ( .A(n25635), .B(n25636), .Z(n25631) );
  AND U34288 ( .A(n25637), .B(n25638), .Z(n25529) );
  NAND U34289 ( .A(n25639), .B(n25640), .Z(n25638) );
  NAND U34290 ( .A(n25641), .B(n25642), .Z(n25637) );
  AND U34291 ( .A(n25643), .B(n25644), .Z(n25531) );
  XOR U34292 ( .A(n25611), .B(n25610), .Z(N63114) );
  XNOR U34293 ( .A(n25628), .B(n25629), .Z(n25610) );
  XNOR U34294 ( .A(n25643), .B(n25644), .Z(n25629) );
  XOR U34295 ( .A(n25640), .B(n25639), .Z(n25644) );
  XOR U34296 ( .A(y[4668]), .B(x[4668]), .Z(n25639) );
  XOR U34297 ( .A(n25642), .B(n25641), .Z(n25640) );
  XOR U34298 ( .A(y[4670]), .B(x[4670]), .Z(n25641) );
  XOR U34299 ( .A(y[4669]), .B(x[4669]), .Z(n25642) );
  XOR U34300 ( .A(n25634), .B(n25633), .Z(n25643) );
  XOR U34301 ( .A(n25636), .B(n25635), .Z(n25633) );
  XOR U34302 ( .A(y[4667]), .B(x[4667]), .Z(n25635) );
  XOR U34303 ( .A(y[4666]), .B(x[4666]), .Z(n25636) );
  XOR U34304 ( .A(y[4665]), .B(x[4665]), .Z(n25634) );
  XNOR U34305 ( .A(n25627), .B(n25626), .Z(n25628) );
  XNOR U34306 ( .A(n25623), .B(n25622), .Z(n25626) );
  XOR U34307 ( .A(n25625), .B(n25624), .Z(n25622) );
  XOR U34308 ( .A(y[4664]), .B(x[4664]), .Z(n25624) );
  XOR U34309 ( .A(y[4663]), .B(x[4663]), .Z(n25625) );
  XOR U34310 ( .A(y[4662]), .B(x[4662]), .Z(n25623) );
  XOR U34311 ( .A(n25617), .B(n25616), .Z(n25627) );
  XOR U34312 ( .A(n25619), .B(n25618), .Z(n25616) );
  XOR U34313 ( .A(y[4661]), .B(x[4661]), .Z(n25618) );
  XOR U34314 ( .A(y[4660]), .B(x[4660]), .Z(n25619) );
  XOR U34315 ( .A(y[4659]), .B(x[4659]), .Z(n25617) );
  XNOR U34316 ( .A(n25593), .B(n25594), .Z(n25611) );
  XNOR U34317 ( .A(n25608), .B(n25609), .Z(n25594) );
  XOR U34318 ( .A(n25605), .B(n25604), .Z(n25609) );
  XOR U34319 ( .A(y[4656]), .B(x[4656]), .Z(n25604) );
  XOR U34320 ( .A(n25607), .B(n25606), .Z(n25605) );
  XOR U34321 ( .A(y[4658]), .B(x[4658]), .Z(n25606) );
  XOR U34322 ( .A(y[4657]), .B(x[4657]), .Z(n25607) );
  XOR U34323 ( .A(n25599), .B(n25598), .Z(n25608) );
  XOR U34324 ( .A(n25601), .B(n25600), .Z(n25598) );
  XOR U34325 ( .A(y[4655]), .B(x[4655]), .Z(n25600) );
  XOR U34326 ( .A(y[4654]), .B(x[4654]), .Z(n25601) );
  XOR U34327 ( .A(y[4653]), .B(x[4653]), .Z(n25599) );
  XNOR U34328 ( .A(n25592), .B(n25591), .Z(n25593) );
  XNOR U34329 ( .A(n25588), .B(n25587), .Z(n25591) );
  XOR U34330 ( .A(n25590), .B(n25589), .Z(n25587) );
  XOR U34331 ( .A(y[4652]), .B(x[4652]), .Z(n25589) );
  XOR U34332 ( .A(y[4651]), .B(x[4651]), .Z(n25590) );
  XOR U34333 ( .A(y[4650]), .B(x[4650]), .Z(n25588) );
  XOR U34334 ( .A(n25582), .B(n25581), .Z(n25592) );
  XOR U34335 ( .A(n25584), .B(n25583), .Z(n25581) );
  XOR U34336 ( .A(y[4649]), .B(x[4649]), .Z(n25583) );
  XOR U34337 ( .A(y[4648]), .B(x[4648]), .Z(n25584) );
  XOR U34338 ( .A(y[4647]), .B(x[4647]), .Z(n25582) );
  NAND U34339 ( .A(n25645), .B(n25646), .Z(N63105) );
  NAND U34340 ( .A(n25647), .B(n25648), .Z(n25646) );
  NANDN U34341 ( .A(n25649), .B(n25650), .Z(n25648) );
  NANDN U34342 ( .A(n25650), .B(n25649), .Z(n25645) );
  XOR U34343 ( .A(n25649), .B(n25651), .Z(N63104) );
  XNOR U34344 ( .A(n25647), .B(n25650), .Z(n25651) );
  NAND U34345 ( .A(n25652), .B(n25653), .Z(n25650) );
  NAND U34346 ( .A(n25654), .B(n25655), .Z(n25653) );
  NANDN U34347 ( .A(n25656), .B(n25657), .Z(n25655) );
  NANDN U34348 ( .A(n25657), .B(n25656), .Z(n25652) );
  AND U34349 ( .A(n25658), .B(n25659), .Z(n25647) );
  NAND U34350 ( .A(n25660), .B(n25661), .Z(n25659) );
  NANDN U34351 ( .A(n25662), .B(n25663), .Z(n25661) );
  NANDN U34352 ( .A(n25663), .B(n25662), .Z(n25658) );
  IV U34353 ( .A(n25664), .Z(n25663) );
  AND U34354 ( .A(n25665), .B(n25666), .Z(n25649) );
  NAND U34355 ( .A(n25667), .B(n25668), .Z(n25666) );
  NANDN U34356 ( .A(n25669), .B(n25670), .Z(n25668) );
  NANDN U34357 ( .A(n25670), .B(n25669), .Z(n25665) );
  XOR U34358 ( .A(n25662), .B(n25671), .Z(N63103) );
  XNOR U34359 ( .A(n25660), .B(n25664), .Z(n25671) );
  XOR U34360 ( .A(n25657), .B(n25672), .Z(n25664) );
  XNOR U34361 ( .A(n25654), .B(n25656), .Z(n25672) );
  AND U34362 ( .A(n25673), .B(n25674), .Z(n25656) );
  NANDN U34363 ( .A(n25675), .B(n25676), .Z(n25674) );
  OR U34364 ( .A(n25677), .B(n25678), .Z(n25676) );
  IV U34365 ( .A(n25679), .Z(n25678) );
  NANDN U34366 ( .A(n25679), .B(n25677), .Z(n25673) );
  AND U34367 ( .A(n25680), .B(n25681), .Z(n25654) );
  NAND U34368 ( .A(n25682), .B(n25683), .Z(n25681) );
  NANDN U34369 ( .A(n25684), .B(n25685), .Z(n25683) );
  NANDN U34370 ( .A(n25685), .B(n25684), .Z(n25680) );
  IV U34371 ( .A(n25686), .Z(n25685) );
  NAND U34372 ( .A(n25687), .B(n25688), .Z(n25657) );
  NANDN U34373 ( .A(n25689), .B(n25690), .Z(n25688) );
  NANDN U34374 ( .A(n25691), .B(n25692), .Z(n25690) );
  NANDN U34375 ( .A(n25692), .B(n25691), .Z(n25687) );
  IV U34376 ( .A(n25693), .Z(n25691) );
  AND U34377 ( .A(n25694), .B(n25695), .Z(n25660) );
  NAND U34378 ( .A(n25696), .B(n25697), .Z(n25695) );
  NANDN U34379 ( .A(n25698), .B(n25699), .Z(n25697) );
  NANDN U34380 ( .A(n25699), .B(n25698), .Z(n25694) );
  XOR U34381 ( .A(n25670), .B(n25700), .Z(n25662) );
  XNOR U34382 ( .A(n25667), .B(n25669), .Z(n25700) );
  AND U34383 ( .A(n25701), .B(n25702), .Z(n25669) );
  NANDN U34384 ( .A(n25703), .B(n25704), .Z(n25702) );
  OR U34385 ( .A(n25705), .B(n25706), .Z(n25704) );
  IV U34386 ( .A(n25707), .Z(n25706) );
  NANDN U34387 ( .A(n25707), .B(n25705), .Z(n25701) );
  AND U34388 ( .A(n25708), .B(n25709), .Z(n25667) );
  NAND U34389 ( .A(n25710), .B(n25711), .Z(n25709) );
  NANDN U34390 ( .A(n25712), .B(n25713), .Z(n25711) );
  NANDN U34391 ( .A(n25713), .B(n25712), .Z(n25708) );
  IV U34392 ( .A(n25714), .Z(n25713) );
  NAND U34393 ( .A(n25715), .B(n25716), .Z(n25670) );
  NANDN U34394 ( .A(n25717), .B(n25718), .Z(n25716) );
  NANDN U34395 ( .A(n25719), .B(n25720), .Z(n25718) );
  NANDN U34396 ( .A(n25720), .B(n25719), .Z(n25715) );
  IV U34397 ( .A(n25721), .Z(n25719) );
  XOR U34398 ( .A(n25696), .B(n25722), .Z(N63102) );
  XNOR U34399 ( .A(n25699), .B(n25698), .Z(n25722) );
  XNOR U34400 ( .A(n25710), .B(n25723), .Z(n25698) );
  XNOR U34401 ( .A(n25714), .B(n25712), .Z(n25723) );
  XOR U34402 ( .A(n25720), .B(n25724), .Z(n25712) );
  XNOR U34403 ( .A(n25717), .B(n25721), .Z(n25724) );
  AND U34404 ( .A(n25725), .B(n25726), .Z(n25721) );
  NAND U34405 ( .A(n25727), .B(n25728), .Z(n25726) );
  NAND U34406 ( .A(n25729), .B(n25730), .Z(n25725) );
  AND U34407 ( .A(n25731), .B(n25732), .Z(n25717) );
  NAND U34408 ( .A(n25733), .B(n25734), .Z(n25732) );
  NAND U34409 ( .A(n25735), .B(n25736), .Z(n25731) );
  NANDN U34410 ( .A(n25737), .B(n25738), .Z(n25720) );
  ANDN U34411 ( .B(n25739), .A(n25740), .Z(n25714) );
  XNOR U34412 ( .A(n25705), .B(n25741), .Z(n25710) );
  XNOR U34413 ( .A(n25703), .B(n25707), .Z(n25741) );
  AND U34414 ( .A(n25742), .B(n25743), .Z(n25707) );
  NAND U34415 ( .A(n25744), .B(n25745), .Z(n25743) );
  NAND U34416 ( .A(n25746), .B(n25747), .Z(n25742) );
  AND U34417 ( .A(n25748), .B(n25749), .Z(n25703) );
  NAND U34418 ( .A(n25750), .B(n25751), .Z(n25749) );
  NAND U34419 ( .A(n25752), .B(n25753), .Z(n25748) );
  AND U34420 ( .A(n25754), .B(n25755), .Z(n25705) );
  NAND U34421 ( .A(n25756), .B(n25757), .Z(n25699) );
  XNOR U34422 ( .A(n25682), .B(n25758), .Z(n25696) );
  XNOR U34423 ( .A(n25686), .B(n25684), .Z(n25758) );
  XOR U34424 ( .A(n25692), .B(n25759), .Z(n25684) );
  XNOR U34425 ( .A(n25689), .B(n25693), .Z(n25759) );
  AND U34426 ( .A(n25760), .B(n25761), .Z(n25693) );
  NAND U34427 ( .A(n25762), .B(n25763), .Z(n25761) );
  NAND U34428 ( .A(n25764), .B(n25765), .Z(n25760) );
  AND U34429 ( .A(n25766), .B(n25767), .Z(n25689) );
  NAND U34430 ( .A(n25768), .B(n25769), .Z(n25767) );
  NAND U34431 ( .A(n25770), .B(n25771), .Z(n25766) );
  NANDN U34432 ( .A(n25772), .B(n25773), .Z(n25692) );
  ANDN U34433 ( .B(n25774), .A(n25775), .Z(n25686) );
  XNOR U34434 ( .A(n25677), .B(n25776), .Z(n25682) );
  XNOR U34435 ( .A(n25675), .B(n25679), .Z(n25776) );
  AND U34436 ( .A(n25777), .B(n25778), .Z(n25679) );
  NAND U34437 ( .A(n25779), .B(n25780), .Z(n25778) );
  NAND U34438 ( .A(n25781), .B(n25782), .Z(n25777) );
  AND U34439 ( .A(n25783), .B(n25784), .Z(n25675) );
  NAND U34440 ( .A(n25785), .B(n25786), .Z(n25784) );
  NAND U34441 ( .A(n25787), .B(n25788), .Z(n25783) );
  AND U34442 ( .A(n25789), .B(n25790), .Z(n25677) );
  XOR U34443 ( .A(n25757), .B(n25756), .Z(N63101) );
  XNOR U34444 ( .A(n25774), .B(n25775), .Z(n25756) );
  XNOR U34445 ( .A(n25789), .B(n25790), .Z(n25775) );
  XOR U34446 ( .A(n25786), .B(n25785), .Z(n25790) );
  XOR U34447 ( .A(y[4644]), .B(x[4644]), .Z(n25785) );
  XOR U34448 ( .A(n25788), .B(n25787), .Z(n25786) );
  XOR U34449 ( .A(y[4646]), .B(x[4646]), .Z(n25787) );
  XOR U34450 ( .A(y[4645]), .B(x[4645]), .Z(n25788) );
  XOR U34451 ( .A(n25780), .B(n25779), .Z(n25789) );
  XOR U34452 ( .A(n25782), .B(n25781), .Z(n25779) );
  XOR U34453 ( .A(y[4643]), .B(x[4643]), .Z(n25781) );
  XOR U34454 ( .A(y[4642]), .B(x[4642]), .Z(n25782) );
  XOR U34455 ( .A(y[4641]), .B(x[4641]), .Z(n25780) );
  XNOR U34456 ( .A(n25773), .B(n25772), .Z(n25774) );
  XNOR U34457 ( .A(n25769), .B(n25768), .Z(n25772) );
  XOR U34458 ( .A(n25771), .B(n25770), .Z(n25768) );
  XOR U34459 ( .A(y[4640]), .B(x[4640]), .Z(n25770) );
  XOR U34460 ( .A(y[4639]), .B(x[4639]), .Z(n25771) );
  XOR U34461 ( .A(y[4638]), .B(x[4638]), .Z(n25769) );
  XOR U34462 ( .A(n25763), .B(n25762), .Z(n25773) );
  XOR U34463 ( .A(n25765), .B(n25764), .Z(n25762) );
  XOR U34464 ( .A(y[4637]), .B(x[4637]), .Z(n25764) );
  XOR U34465 ( .A(y[4636]), .B(x[4636]), .Z(n25765) );
  XOR U34466 ( .A(y[4635]), .B(x[4635]), .Z(n25763) );
  XNOR U34467 ( .A(n25739), .B(n25740), .Z(n25757) );
  XNOR U34468 ( .A(n25754), .B(n25755), .Z(n25740) );
  XOR U34469 ( .A(n25751), .B(n25750), .Z(n25755) );
  XOR U34470 ( .A(y[4632]), .B(x[4632]), .Z(n25750) );
  XOR U34471 ( .A(n25753), .B(n25752), .Z(n25751) );
  XOR U34472 ( .A(y[4634]), .B(x[4634]), .Z(n25752) );
  XOR U34473 ( .A(y[4633]), .B(x[4633]), .Z(n25753) );
  XOR U34474 ( .A(n25745), .B(n25744), .Z(n25754) );
  XOR U34475 ( .A(n25747), .B(n25746), .Z(n25744) );
  XOR U34476 ( .A(y[4631]), .B(x[4631]), .Z(n25746) );
  XOR U34477 ( .A(y[4630]), .B(x[4630]), .Z(n25747) );
  XOR U34478 ( .A(y[4629]), .B(x[4629]), .Z(n25745) );
  XNOR U34479 ( .A(n25738), .B(n25737), .Z(n25739) );
  XNOR U34480 ( .A(n25734), .B(n25733), .Z(n25737) );
  XOR U34481 ( .A(n25736), .B(n25735), .Z(n25733) );
  XOR U34482 ( .A(y[4628]), .B(x[4628]), .Z(n25735) );
  XOR U34483 ( .A(y[4627]), .B(x[4627]), .Z(n25736) );
  XOR U34484 ( .A(y[4626]), .B(x[4626]), .Z(n25734) );
  XOR U34485 ( .A(n25728), .B(n25727), .Z(n25738) );
  XOR U34486 ( .A(n25730), .B(n25729), .Z(n25727) );
  XOR U34487 ( .A(y[4625]), .B(x[4625]), .Z(n25729) );
  XOR U34488 ( .A(y[4624]), .B(x[4624]), .Z(n25730) );
  XOR U34489 ( .A(y[4623]), .B(x[4623]), .Z(n25728) );
  NAND U34490 ( .A(n25791), .B(n25792), .Z(N63092) );
  NAND U34491 ( .A(n25793), .B(n25794), .Z(n25792) );
  NANDN U34492 ( .A(n25795), .B(n25796), .Z(n25794) );
  NANDN U34493 ( .A(n25796), .B(n25795), .Z(n25791) );
  XOR U34494 ( .A(n25795), .B(n25797), .Z(N63091) );
  XNOR U34495 ( .A(n25793), .B(n25796), .Z(n25797) );
  NAND U34496 ( .A(n25798), .B(n25799), .Z(n25796) );
  NAND U34497 ( .A(n25800), .B(n25801), .Z(n25799) );
  NANDN U34498 ( .A(n25802), .B(n25803), .Z(n25801) );
  NANDN U34499 ( .A(n25803), .B(n25802), .Z(n25798) );
  AND U34500 ( .A(n25804), .B(n25805), .Z(n25793) );
  NAND U34501 ( .A(n25806), .B(n25807), .Z(n25805) );
  NANDN U34502 ( .A(n25808), .B(n25809), .Z(n25807) );
  NANDN U34503 ( .A(n25809), .B(n25808), .Z(n25804) );
  IV U34504 ( .A(n25810), .Z(n25809) );
  AND U34505 ( .A(n25811), .B(n25812), .Z(n25795) );
  NAND U34506 ( .A(n25813), .B(n25814), .Z(n25812) );
  NANDN U34507 ( .A(n25815), .B(n25816), .Z(n25814) );
  NANDN U34508 ( .A(n25816), .B(n25815), .Z(n25811) );
  XOR U34509 ( .A(n25808), .B(n25817), .Z(N63090) );
  XNOR U34510 ( .A(n25806), .B(n25810), .Z(n25817) );
  XOR U34511 ( .A(n25803), .B(n25818), .Z(n25810) );
  XNOR U34512 ( .A(n25800), .B(n25802), .Z(n25818) );
  AND U34513 ( .A(n25819), .B(n25820), .Z(n25802) );
  NANDN U34514 ( .A(n25821), .B(n25822), .Z(n25820) );
  OR U34515 ( .A(n25823), .B(n25824), .Z(n25822) );
  IV U34516 ( .A(n25825), .Z(n25824) );
  NANDN U34517 ( .A(n25825), .B(n25823), .Z(n25819) );
  AND U34518 ( .A(n25826), .B(n25827), .Z(n25800) );
  NAND U34519 ( .A(n25828), .B(n25829), .Z(n25827) );
  NANDN U34520 ( .A(n25830), .B(n25831), .Z(n25829) );
  NANDN U34521 ( .A(n25831), .B(n25830), .Z(n25826) );
  IV U34522 ( .A(n25832), .Z(n25831) );
  NAND U34523 ( .A(n25833), .B(n25834), .Z(n25803) );
  NANDN U34524 ( .A(n25835), .B(n25836), .Z(n25834) );
  NANDN U34525 ( .A(n25837), .B(n25838), .Z(n25836) );
  NANDN U34526 ( .A(n25838), .B(n25837), .Z(n25833) );
  IV U34527 ( .A(n25839), .Z(n25837) );
  AND U34528 ( .A(n25840), .B(n25841), .Z(n25806) );
  NAND U34529 ( .A(n25842), .B(n25843), .Z(n25841) );
  NANDN U34530 ( .A(n25844), .B(n25845), .Z(n25843) );
  NANDN U34531 ( .A(n25845), .B(n25844), .Z(n25840) );
  XOR U34532 ( .A(n25816), .B(n25846), .Z(n25808) );
  XNOR U34533 ( .A(n25813), .B(n25815), .Z(n25846) );
  AND U34534 ( .A(n25847), .B(n25848), .Z(n25815) );
  NANDN U34535 ( .A(n25849), .B(n25850), .Z(n25848) );
  OR U34536 ( .A(n25851), .B(n25852), .Z(n25850) );
  IV U34537 ( .A(n25853), .Z(n25852) );
  NANDN U34538 ( .A(n25853), .B(n25851), .Z(n25847) );
  AND U34539 ( .A(n25854), .B(n25855), .Z(n25813) );
  NAND U34540 ( .A(n25856), .B(n25857), .Z(n25855) );
  NANDN U34541 ( .A(n25858), .B(n25859), .Z(n25857) );
  NANDN U34542 ( .A(n25859), .B(n25858), .Z(n25854) );
  IV U34543 ( .A(n25860), .Z(n25859) );
  NAND U34544 ( .A(n25861), .B(n25862), .Z(n25816) );
  NANDN U34545 ( .A(n25863), .B(n25864), .Z(n25862) );
  NANDN U34546 ( .A(n25865), .B(n25866), .Z(n25864) );
  NANDN U34547 ( .A(n25866), .B(n25865), .Z(n25861) );
  IV U34548 ( .A(n25867), .Z(n25865) );
  XOR U34549 ( .A(n25842), .B(n25868), .Z(N63089) );
  XNOR U34550 ( .A(n25845), .B(n25844), .Z(n25868) );
  XNOR U34551 ( .A(n25856), .B(n25869), .Z(n25844) );
  XNOR U34552 ( .A(n25860), .B(n25858), .Z(n25869) );
  XOR U34553 ( .A(n25866), .B(n25870), .Z(n25858) );
  XNOR U34554 ( .A(n25863), .B(n25867), .Z(n25870) );
  AND U34555 ( .A(n25871), .B(n25872), .Z(n25867) );
  NAND U34556 ( .A(n25873), .B(n25874), .Z(n25872) );
  NAND U34557 ( .A(n25875), .B(n25876), .Z(n25871) );
  AND U34558 ( .A(n25877), .B(n25878), .Z(n25863) );
  NAND U34559 ( .A(n25879), .B(n25880), .Z(n25878) );
  NAND U34560 ( .A(n25881), .B(n25882), .Z(n25877) );
  NANDN U34561 ( .A(n25883), .B(n25884), .Z(n25866) );
  ANDN U34562 ( .B(n25885), .A(n25886), .Z(n25860) );
  XNOR U34563 ( .A(n25851), .B(n25887), .Z(n25856) );
  XNOR U34564 ( .A(n25849), .B(n25853), .Z(n25887) );
  AND U34565 ( .A(n25888), .B(n25889), .Z(n25853) );
  NAND U34566 ( .A(n25890), .B(n25891), .Z(n25889) );
  NAND U34567 ( .A(n25892), .B(n25893), .Z(n25888) );
  AND U34568 ( .A(n25894), .B(n25895), .Z(n25849) );
  NAND U34569 ( .A(n25896), .B(n25897), .Z(n25895) );
  NAND U34570 ( .A(n25898), .B(n25899), .Z(n25894) );
  AND U34571 ( .A(n25900), .B(n25901), .Z(n25851) );
  NAND U34572 ( .A(n25902), .B(n25903), .Z(n25845) );
  XNOR U34573 ( .A(n25828), .B(n25904), .Z(n25842) );
  XNOR U34574 ( .A(n25832), .B(n25830), .Z(n25904) );
  XOR U34575 ( .A(n25838), .B(n25905), .Z(n25830) );
  XNOR U34576 ( .A(n25835), .B(n25839), .Z(n25905) );
  AND U34577 ( .A(n25906), .B(n25907), .Z(n25839) );
  NAND U34578 ( .A(n25908), .B(n25909), .Z(n25907) );
  NAND U34579 ( .A(n25910), .B(n25911), .Z(n25906) );
  AND U34580 ( .A(n25912), .B(n25913), .Z(n25835) );
  NAND U34581 ( .A(n25914), .B(n25915), .Z(n25913) );
  NAND U34582 ( .A(n25916), .B(n25917), .Z(n25912) );
  NANDN U34583 ( .A(n25918), .B(n25919), .Z(n25838) );
  ANDN U34584 ( .B(n25920), .A(n25921), .Z(n25832) );
  XNOR U34585 ( .A(n25823), .B(n25922), .Z(n25828) );
  XNOR U34586 ( .A(n25821), .B(n25825), .Z(n25922) );
  AND U34587 ( .A(n25923), .B(n25924), .Z(n25825) );
  NAND U34588 ( .A(n25925), .B(n25926), .Z(n25924) );
  NAND U34589 ( .A(n25927), .B(n25928), .Z(n25923) );
  AND U34590 ( .A(n25929), .B(n25930), .Z(n25821) );
  NAND U34591 ( .A(n25931), .B(n25932), .Z(n25930) );
  NAND U34592 ( .A(n25933), .B(n25934), .Z(n25929) );
  AND U34593 ( .A(n25935), .B(n25936), .Z(n25823) );
  XOR U34594 ( .A(n25903), .B(n25902), .Z(N63088) );
  XNOR U34595 ( .A(n25920), .B(n25921), .Z(n25902) );
  XNOR U34596 ( .A(n25935), .B(n25936), .Z(n25921) );
  XOR U34597 ( .A(n25932), .B(n25931), .Z(n25936) );
  XOR U34598 ( .A(y[4620]), .B(x[4620]), .Z(n25931) );
  XOR U34599 ( .A(n25934), .B(n25933), .Z(n25932) );
  XOR U34600 ( .A(y[4622]), .B(x[4622]), .Z(n25933) );
  XOR U34601 ( .A(y[4621]), .B(x[4621]), .Z(n25934) );
  XOR U34602 ( .A(n25926), .B(n25925), .Z(n25935) );
  XOR U34603 ( .A(n25928), .B(n25927), .Z(n25925) );
  XOR U34604 ( .A(y[4619]), .B(x[4619]), .Z(n25927) );
  XOR U34605 ( .A(y[4618]), .B(x[4618]), .Z(n25928) );
  XOR U34606 ( .A(y[4617]), .B(x[4617]), .Z(n25926) );
  XNOR U34607 ( .A(n25919), .B(n25918), .Z(n25920) );
  XNOR U34608 ( .A(n25915), .B(n25914), .Z(n25918) );
  XOR U34609 ( .A(n25917), .B(n25916), .Z(n25914) );
  XOR U34610 ( .A(y[4616]), .B(x[4616]), .Z(n25916) );
  XOR U34611 ( .A(y[4615]), .B(x[4615]), .Z(n25917) );
  XOR U34612 ( .A(y[4614]), .B(x[4614]), .Z(n25915) );
  XOR U34613 ( .A(n25909), .B(n25908), .Z(n25919) );
  XOR U34614 ( .A(n25911), .B(n25910), .Z(n25908) );
  XOR U34615 ( .A(y[4613]), .B(x[4613]), .Z(n25910) );
  XOR U34616 ( .A(y[4612]), .B(x[4612]), .Z(n25911) );
  XOR U34617 ( .A(y[4611]), .B(x[4611]), .Z(n25909) );
  XNOR U34618 ( .A(n25885), .B(n25886), .Z(n25903) );
  XNOR U34619 ( .A(n25900), .B(n25901), .Z(n25886) );
  XOR U34620 ( .A(n25897), .B(n25896), .Z(n25901) );
  XOR U34621 ( .A(y[4608]), .B(x[4608]), .Z(n25896) );
  XOR U34622 ( .A(n25899), .B(n25898), .Z(n25897) );
  XOR U34623 ( .A(y[4610]), .B(x[4610]), .Z(n25898) );
  XOR U34624 ( .A(y[4609]), .B(x[4609]), .Z(n25899) );
  XOR U34625 ( .A(n25891), .B(n25890), .Z(n25900) );
  XOR U34626 ( .A(n25893), .B(n25892), .Z(n25890) );
  XOR U34627 ( .A(y[4607]), .B(x[4607]), .Z(n25892) );
  XOR U34628 ( .A(y[4606]), .B(x[4606]), .Z(n25893) );
  XOR U34629 ( .A(y[4605]), .B(x[4605]), .Z(n25891) );
  XNOR U34630 ( .A(n25884), .B(n25883), .Z(n25885) );
  XNOR U34631 ( .A(n25880), .B(n25879), .Z(n25883) );
  XOR U34632 ( .A(n25882), .B(n25881), .Z(n25879) );
  XOR U34633 ( .A(y[4604]), .B(x[4604]), .Z(n25881) );
  XOR U34634 ( .A(y[4603]), .B(x[4603]), .Z(n25882) );
  XOR U34635 ( .A(y[4602]), .B(x[4602]), .Z(n25880) );
  XOR U34636 ( .A(n25874), .B(n25873), .Z(n25884) );
  XOR U34637 ( .A(n25876), .B(n25875), .Z(n25873) );
  XOR U34638 ( .A(y[4601]), .B(x[4601]), .Z(n25875) );
  XOR U34639 ( .A(y[4600]), .B(x[4600]), .Z(n25876) );
  XOR U34640 ( .A(y[4599]), .B(x[4599]), .Z(n25874) );
  NAND U34641 ( .A(n25937), .B(n25938), .Z(N63079) );
  NAND U34642 ( .A(n25939), .B(n25940), .Z(n25938) );
  NANDN U34643 ( .A(n25941), .B(n25942), .Z(n25940) );
  NANDN U34644 ( .A(n25942), .B(n25941), .Z(n25937) );
  XOR U34645 ( .A(n25941), .B(n25943), .Z(N63078) );
  XNOR U34646 ( .A(n25939), .B(n25942), .Z(n25943) );
  NAND U34647 ( .A(n25944), .B(n25945), .Z(n25942) );
  NAND U34648 ( .A(n25946), .B(n25947), .Z(n25945) );
  NANDN U34649 ( .A(n25948), .B(n25949), .Z(n25947) );
  NANDN U34650 ( .A(n25949), .B(n25948), .Z(n25944) );
  AND U34651 ( .A(n25950), .B(n25951), .Z(n25939) );
  NAND U34652 ( .A(n25952), .B(n25953), .Z(n25951) );
  NANDN U34653 ( .A(n25954), .B(n25955), .Z(n25953) );
  NANDN U34654 ( .A(n25955), .B(n25954), .Z(n25950) );
  IV U34655 ( .A(n25956), .Z(n25955) );
  AND U34656 ( .A(n25957), .B(n25958), .Z(n25941) );
  NAND U34657 ( .A(n25959), .B(n25960), .Z(n25958) );
  NANDN U34658 ( .A(n25961), .B(n25962), .Z(n25960) );
  NANDN U34659 ( .A(n25962), .B(n25961), .Z(n25957) );
  XOR U34660 ( .A(n25954), .B(n25963), .Z(N63077) );
  XNOR U34661 ( .A(n25952), .B(n25956), .Z(n25963) );
  XOR U34662 ( .A(n25949), .B(n25964), .Z(n25956) );
  XNOR U34663 ( .A(n25946), .B(n25948), .Z(n25964) );
  AND U34664 ( .A(n25965), .B(n25966), .Z(n25948) );
  NANDN U34665 ( .A(n25967), .B(n25968), .Z(n25966) );
  OR U34666 ( .A(n25969), .B(n25970), .Z(n25968) );
  IV U34667 ( .A(n25971), .Z(n25970) );
  NANDN U34668 ( .A(n25971), .B(n25969), .Z(n25965) );
  AND U34669 ( .A(n25972), .B(n25973), .Z(n25946) );
  NAND U34670 ( .A(n25974), .B(n25975), .Z(n25973) );
  NANDN U34671 ( .A(n25976), .B(n25977), .Z(n25975) );
  NANDN U34672 ( .A(n25977), .B(n25976), .Z(n25972) );
  IV U34673 ( .A(n25978), .Z(n25977) );
  NAND U34674 ( .A(n25979), .B(n25980), .Z(n25949) );
  NANDN U34675 ( .A(n25981), .B(n25982), .Z(n25980) );
  NANDN U34676 ( .A(n25983), .B(n25984), .Z(n25982) );
  NANDN U34677 ( .A(n25984), .B(n25983), .Z(n25979) );
  IV U34678 ( .A(n25985), .Z(n25983) );
  AND U34679 ( .A(n25986), .B(n25987), .Z(n25952) );
  NAND U34680 ( .A(n25988), .B(n25989), .Z(n25987) );
  NANDN U34681 ( .A(n25990), .B(n25991), .Z(n25989) );
  NANDN U34682 ( .A(n25991), .B(n25990), .Z(n25986) );
  XOR U34683 ( .A(n25962), .B(n25992), .Z(n25954) );
  XNOR U34684 ( .A(n25959), .B(n25961), .Z(n25992) );
  AND U34685 ( .A(n25993), .B(n25994), .Z(n25961) );
  NANDN U34686 ( .A(n25995), .B(n25996), .Z(n25994) );
  OR U34687 ( .A(n25997), .B(n25998), .Z(n25996) );
  IV U34688 ( .A(n25999), .Z(n25998) );
  NANDN U34689 ( .A(n25999), .B(n25997), .Z(n25993) );
  AND U34690 ( .A(n26000), .B(n26001), .Z(n25959) );
  NAND U34691 ( .A(n26002), .B(n26003), .Z(n26001) );
  NANDN U34692 ( .A(n26004), .B(n26005), .Z(n26003) );
  NANDN U34693 ( .A(n26005), .B(n26004), .Z(n26000) );
  IV U34694 ( .A(n26006), .Z(n26005) );
  NAND U34695 ( .A(n26007), .B(n26008), .Z(n25962) );
  NANDN U34696 ( .A(n26009), .B(n26010), .Z(n26008) );
  NANDN U34697 ( .A(n26011), .B(n26012), .Z(n26010) );
  NANDN U34698 ( .A(n26012), .B(n26011), .Z(n26007) );
  IV U34699 ( .A(n26013), .Z(n26011) );
  XOR U34700 ( .A(n25988), .B(n26014), .Z(N63076) );
  XNOR U34701 ( .A(n25991), .B(n25990), .Z(n26014) );
  XNOR U34702 ( .A(n26002), .B(n26015), .Z(n25990) );
  XNOR U34703 ( .A(n26006), .B(n26004), .Z(n26015) );
  XOR U34704 ( .A(n26012), .B(n26016), .Z(n26004) );
  XNOR U34705 ( .A(n26009), .B(n26013), .Z(n26016) );
  AND U34706 ( .A(n26017), .B(n26018), .Z(n26013) );
  NAND U34707 ( .A(n26019), .B(n26020), .Z(n26018) );
  NAND U34708 ( .A(n26021), .B(n26022), .Z(n26017) );
  AND U34709 ( .A(n26023), .B(n26024), .Z(n26009) );
  NAND U34710 ( .A(n26025), .B(n26026), .Z(n26024) );
  NAND U34711 ( .A(n26027), .B(n26028), .Z(n26023) );
  NANDN U34712 ( .A(n26029), .B(n26030), .Z(n26012) );
  ANDN U34713 ( .B(n26031), .A(n26032), .Z(n26006) );
  XNOR U34714 ( .A(n25997), .B(n26033), .Z(n26002) );
  XNOR U34715 ( .A(n25995), .B(n25999), .Z(n26033) );
  AND U34716 ( .A(n26034), .B(n26035), .Z(n25999) );
  NAND U34717 ( .A(n26036), .B(n26037), .Z(n26035) );
  NAND U34718 ( .A(n26038), .B(n26039), .Z(n26034) );
  AND U34719 ( .A(n26040), .B(n26041), .Z(n25995) );
  NAND U34720 ( .A(n26042), .B(n26043), .Z(n26041) );
  NAND U34721 ( .A(n26044), .B(n26045), .Z(n26040) );
  AND U34722 ( .A(n26046), .B(n26047), .Z(n25997) );
  NAND U34723 ( .A(n26048), .B(n26049), .Z(n25991) );
  XNOR U34724 ( .A(n25974), .B(n26050), .Z(n25988) );
  XNOR U34725 ( .A(n25978), .B(n25976), .Z(n26050) );
  XOR U34726 ( .A(n25984), .B(n26051), .Z(n25976) );
  XNOR U34727 ( .A(n25981), .B(n25985), .Z(n26051) );
  AND U34728 ( .A(n26052), .B(n26053), .Z(n25985) );
  NAND U34729 ( .A(n26054), .B(n26055), .Z(n26053) );
  NAND U34730 ( .A(n26056), .B(n26057), .Z(n26052) );
  AND U34731 ( .A(n26058), .B(n26059), .Z(n25981) );
  NAND U34732 ( .A(n26060), .B(n26061), .Z(n26059) );
  NAND U34733 ( .A(n26062), .B(n26063), .Z(n26058) );
  NANDN U34734 ( .A(n26064), .B(n26065), .Z(n25984) );
  ANDN U34735 ( .B(n26066), .A(n26067), .Z(n25978) );
  XNOR U34736 ( .A(n25969), .B(n26068), .Z(n25974) );
  XNOR U34737 ( .A(n25967), .B(n25971), .Z(n26068) );
  AND U34738 ( .A(n26069), .B(n26070), .Z(n25971) );
  NAND U34739 ( .A(n26071), .B(n26072), .Z(n26070) );
  NAND U34740 ( .A(n26073), .B(n26074), .Z(n26069) );
  AND U34741 ( .A(n26075), .B(n26076), .Z(n25967) );
  NAND U34742 ( .A(n26077), .B(n26078), .Z(n26076) );
  NAND U34743 ( .A(n26079), .B(n26080), .Z(n26075) );
  AND U34744 ( .A(n26081), .B(n26082), .Z(n25969) );
  XOR U34745 ( .A(n26049), .B(n26048), .Z(N63075) );
  XNOR U34746 ( .A(n26066), .B(n26067), .Z(n26048) );
  XNOR U34747 ( .A(n26081), .B(n26082), .Z(n26067) );
  XOR U34748 ( .A(n26078), .B(n26077), .Z(n26082) );
  XOR U34749 ( .A(y[4596]), .B(x[4596]), .Z(n26077) );
  XOR U34750 ( .A(n26080), .B(n26079), .Z(n26078) );
  XOR U34751 ( .A(y[4598]), .B(x[4598]), .Z(n26079) );
  XOR U34752 ( .A(y[4597]), .B(x[4597]), .Z(n26080) );
  XOR U34753 ( .A(n26072), .B(n26071), .Z(n26081) );
  XOR U34754 ( .A(n26074), .B(n26073), .Z(n26071) );
  XOR U34755 ( .A(y[4595]), .B(x[4595]), .Z(n26073) );
  XOR U34756 ( .A(y[4594]), .B(x[4594]), .Z(n26074) );
  XOR U34757 ( .A(y[4593]), .B(x[4593]), .Z(n26072) );
  XNOR U34758 ( .A(n26065), .B(n26064), .Z(n26066) );
  XNOR U34759 ( .A(n26061), .B(n26060), .Z(n26064) );
  XOR U34760 ( .A(n26063), .B(n26062), .Z(n26060) );
  XOR U34761 ( .A(y[4592]), .B(x[4592]), .Z(n26062) );
  XOR U34762 ( .A(y[4591]), .B(x[4591]), .Z(n26063) );
  XOR U34763 ( .A(y[4590]), .B(x[4590]), .Z(n26061) );
  XOR U34764 ( .A(n26055), .B(n26054), .Z(n26065) );
  XOR U34765 ( .A(n26057), .B(n26056), .Z(n26054) );
  XOR U34766 ( .A(y[4589]), .B(x[4589]), .Z(n26056) );
  XOR U34767 ( .A(y[4588]), .B(x[4588]), .Z(n26057) );
  XOR U34768 ( .A(y[4587]), .B(x[4587]), .Z(n26055) );
  XNOR U34769 ( .A(n26031), .B(n26032), .Z(n26049) );
  XNOR U34770 ( .A(n26046), .B(n26047), .Z(n26032) );
  XOR U34771 ( .A(n26043), .B(n26042), .Z(n26047) );
  XOR U34772 ( .A(y[4584]), .B(x[4584]), .Z(n26042) );
  XOR U34773 ( .A(n26045), .B(n26044), .Z(n26043) );
  XOR U34774 ( .A(y[4586]), .B(x[4586]), .Z(n26044) );
  XOR U34775 ( .A(y[4585]), .B(x[4585]), .Z(n26045) );
  XOR U34776 ( .A(n26037), .B(n26036), .Z(n26046) );
  XOR U34777 ( .A(n26039), .B(n26038), .Z(n26036) );
  XOR U34778 ( .A(y[4583]), .B(x[4583]), .Z(n26038) );
  XOR U34779 ( .A(y[4582]), .B(x[4582]), .Z(n26039) );
  XOR U34780 ( .A(y[4581]), .B(x[4581]), .Z(n26037) );
  XNOR U34781 ( .A(n26030), .B(n26029), .Z(n26031) );
  XNOR U34782 ( .A(n26026), .B(n26025), .Z(n26029) );
  XOR U34783 ( .A(n26028), .B(n26027), .Z(n26025) );
  XOR U34784 ( .A(y[4580]), .B(x[4580]), .Z(n26027) );
  XOR U34785 ( .A(y[4579]), .B(x[4579]), .Z(n26028) );
  XOR U34786 ( .A(y[4578]), .B(x[4578]), .Z(n26026) );
  XOR U34787 ( .A(n26020), .B(n26019), .Z(n26030) );
  XOR U34788 ( .A(n26022), .B(n26021), .Z(n26019) );
  XOR U34789 ( .A(y[4577]), .B(x[4577]), .Z(n26021) );
  XOR U34790 ( .A(y[4576]), .B(x[4576]), .Z(n26022) );
  XOR U34791 ( .A(y[4575]), .B(x[4575]), .Z(n26020) );
  NAND U34792 ( .A(n26083), .B(n26084), .Z(N63066) );
  NAND U34793 ( .A(n26085), .B(n26086), .Z(n26084) );
  NANDN U34794 ( .A(n26087), .B(n26088), .Z(n26086) );
  NANDN U34795 ( .A(n26088), .B(n26087), .Z(n26083) );
  XOR U34796 ( .A(n26087), .B(n26089), .Z(N63065) );
  XNOR U34797 ( .A(n26085), .B(n26088), .Z(n26089) );
  NAND U34798 ( .A(n26090), .B(n26091), .Z(n26088) );
  NAND U34799 ( .A(n26092), .B(n26093), .Z(n26091) );
  NANDN U34800 ( .A(n26094), .B(n26095), .Z(n26093) );
  NANDN U34801 ( .A(n26095), .B(n26094), .Z(n26090) );
  AND U34802 ( .A(n26096), .B(n26097), .Z(n26085) );
  NAND U34803 ( .A(n26098), .B(n26099), .Z(n26097) );
  NANDN U34804 ( .A(n26100), .B(n26101), .Z(n26099) );
  NANDN U34805 ( .A(n26101), .B(n26100), .Z(n26096) );
  IV U34806 ( .A(n26102), .Z(n26101) );
  AND U34807 ( .A(n26103), .B(n26104), .Z(n26087) );
  NAND U34808 ( .A(n26105), .B(n26106), .Z(n26104) );
  NANDN U34809 ( .A(n26107), .B(n26108), .Z(n26106) );
  NANDN U34810 ( .A(n26108), .B(n26107), .Z(n26103) );
  XOR U34811 ( .A(n26100), .B(n26109), .Z(N63064) );
  XNOR U34812 ( .A(n26098), .B(n26102), .Z(n26109) );
  XOR U34813 ( .A(n26095), .B(n26110), .Z(n26102) );
  XNOR U34814 ( .A(n26092), .B(n26094), .Z(n26110) );
  AND U34815 ( .A(n26111), .B(n26112), .Z(n26094) );
  NANDN U34816 ( .A(n26113), .B(n26114), .Z(n26112) );
  OR U34817 ( .A(n26115), .B(n26116), .Z(n26114) );
  IV U34818 ( .A(n26117), .Z(n26116) );
  NANDN U34819 ( .A(n26117), .B(n26115), .Z(n26111) );
  AND U34820 ( .A(n26118), .B(n26119), .Z(n26092) );
  NAND U34821 ( .A(n26120), .B(n26121), .Z(n26119) );
  NANDN U34822 ( .A(n26122), .B(n26123), .Z(n26121) );
  NANDN U34823 ( .A(n26123), .B(n26122), .Z(n26118) );
  IV U34824 ( .A(n26124), .Z(n26123) );
  NAND U34825 ( .A(n26125), .B(n26126), .Z(n26095) );
  NANDN U34826 ( .A(n26127), .B(n26128), .Z(n26126) );
  NANDN U34827 ( .A(n26129), .B(n26130), .Z(n26128) );
  NANDN U34828 ( .A(n26130), .B(n26129), .Z(n26125) );
  IV U34829 ( .A(n26131), .Z(n26129) );
  AND U34830 ( .A(n26132), .B(n26133), .Z(n26098) );
  NAND U34831 ( .A(n26134), .B(n26135), .Z(n26133) );
  NANDN U34832 ( .A(n26136), .B(n26137), .Z(n26135) );
  NANDN U34833 ( .A(n26137), .B(n26136), .Z(n26132) );
  XOR U34834 ( .A(n26108), .B(n26138), .Z(n26100) );
  XNOR U34835 ( .A(n26105), .B(n26107), .Z(n26138) );
  AND U34836 ( .A(n26139), .B(n26140), .Z(n26107) );
  NANDN U34837 ( .A(n26141), .B(n26142), .Z(n26140) );
  OR U34838 ( .A(n26143), .B(n26144), .Z(n26142) );
  IV U34839 ( .A(n26145), .Z(n26144) );
  NANDN U34840 ( .A(n26145), .B(n26143), .Z(n26139) );
  AND U34841 ( .A(n26146), .B(n26147), .Z(n26105) );
  NAND U34842 ( .A(n26148), .B(n26149), .Z(n26147) );
  NANDN U34843 ( .A(n26150), .B(n26151), .Z(n26149) );
  NANDN U34844 ( .A(n26151), .B(n26150), .Z(n26146) );
  IV U34845 ( .A(n26152), .Z(n26151) );
  NAND U34846 ( .A(n26153), .B(n26154), .Z(n26108) );
  NANDN U34847 ( .A(n26155), .B(n26156), .Z(n26154) );
  NANDN U34848 ( .A(n26157), .B(n26158), .Z(n26156) );
  NANDN U34849 ( .A(n26158), .B(n26157), .Z(n26153) );
  IV U34850 ( .A(n26159), .Z(n26157) );
  XOR U34851 ( .A(n26134), .B(n26160), .Z(N63063) );
  XNOR U34852 ( .A(n26137), .B(n26136), .Z(n26160) );
  XNOR U34853 ( .A(n26148), .B(n26161), .Z(n26136) );
  XNOR U34854 ( .A(n26152), .B(n26150), .Z(n26161) );
  XOR U34855 ( .A(n26158), .B(n26162), .Z(n26150) );
  XNOR U34856 ( .A(n26155), .B(n26159), .Z(n26162) );
  AND U34857 ( .A(n26163), .B(n26164), .Z(n26159) );
  NAND U34858 ( .A(n26165), .B(n26166), .Z(n26164) );
  NAND U34859 ( .A(n26167), .B(n26168), .Z(n26163) );
  AND U34860 ( .A(n26169), .B(n26170), .Z(n26155) );
  NAND U34861 ( .A(n26171), .B(n26172), .Z(n26170) );
  NAND U34862 ( .A(n26173), .B(n26174), .Z(n26169) );
  NANDN U34863 ( .A(n26175), .B(n26176), .Z(n26158) );
  ANDN U34864 ( .B(n26177), .A(n26178), .Z(n26152) );
  XNOR U34865 ( .A(n26143), .B(n26179), .Z(n26148) );
  XNOR U34866 ( .A(n26141), .B(n26145), .Z(n26179) );
  AND U34867 ( .A(n26180), .B(n26181), .Z(n26145) );
  NAND U34868 ( .A(n26182), .B(n26183), .Z(n26181) );
  NAND U34869 ( .A(n26184), .B(n26185), .Z(n26180) );
  AND U34870 ( .A(n26186), .B(n26187), .Z(n26141) );
  NAND U34871 ( .A(n26188), .B(n26189), .Z(n26187) );
  NAND U34872 ( .A(n26190), .B(n26191), .Z(n26186) );
  AND U34873 ( .A(n26192), .B(n26193), .Z(n26143) );
  NAND U34874 ( .A(n26194), .B(n26195), .Z(n26137) );
  XNOR U34875 ( .A(n26120), .B(n26196), .Z(n26134) );
  XNOR U34876 ( .A(n26124), .B(n26122), .Z(n26196) );
  XOR U34877 ( .A(n26130), .B(n26197), .Z(n26122) );
  XNOR U34878 ( .A(n26127), .B(n26131), .Z(n26197) );
  AND U34879 ( .A(n26198), .B(n26199), .Z(n26131) );
  NAND U34880 ( .A(n26200), .B(n26201), .Z(n26199) );
  NAND U34881 ( .A(n26202), .B(n26203), .Z(n26198) );
  AND U34882 ( .A(n26204), .B(n26205), .Z(n26127) );
  NAND U34883 ( .A(n26206), .B(n26207), .Z(n26205) );
  NAND U34884 ( .A(n26208), .B(n26209), .Z(n26204) );
  NANDN U34885 ( .A(n26210), .B(n26211), .Z(n26130) );
  ANDN U34886 ( .B(n26212), .A(n26213), .Z(n26124) );
  XNOR U34887 ( .A(n26115), .B(n26214), .Z(n26120) );
  XNOR U34888 ( .A(n26113), .B(n26117), .Z(n26214) );
  AND U34889 ( .A(n26215), .B(n26216), .Z(n26117) );
  NAND U34890 ( .A(n26217), .B(n26218), .Z(n26216) );
  NAND U34891 ( .A(n26219), .B(n26220), .Z(n26215) );
  AND U34892 ( .A(n26221), .B(n26222), .Z(n26113) );
  NAND U34893 ( .A(n26223), .B(n26224), .Z(n26222) );
  NAND U34894 ( .A(n26225), .B(n26226), .Z(n26221) );
  AND U34895 ( .A(n26227), .B(n26228), .Z(n26115) );
  XOR U34896 ( .A(n26195), .B(n26194), .Z(N63062) );
  XNOR U34897 ( .A(n26212), .B(n26213), .Z(n26194) );
  XNOR U34898 ( .A(n26227), .B(n26228), .Z(n26213) );
  XOR U34899 ( .A(n26224), .B(n26223), .Z(n26228) );
  XOR U34900 ( .A(y[4572]), .B(x[4572]), .Z(n26223) );
  XOR U34901 ( .A(n26226), .B(n26225), .Z(n26224) );
  XOR U34902 ( .A(y[4574]), .B(x[4574]), .Z(n26225) );
  XOR U34903 ( .A(y[4573]), .B(x[4573]), .Z(n26226) );
  XOR U34904 ( .A(n26218), .B(n26217), .Z(n26227) );
  XOR U34905 ( .A(n26220), .B(n26219), .Z(n26217) );
  XOR U34906 ( .A(y[4571]), .B(x[4571]), .Z(n26219) );
  XOR U34907 ( .A(y[4570]), .B(x[4570]), .Z(n26220) );
  XOR U34908 ( .A(y[4569]), .B(x[4569]), .Z(n26218) );
  XNOR U34909 ( .A(n26211), .B(n26210), .Z(n26212) );
  XNOR U34910 ( .A(n26207), .B(n26206), .Z(n26210) );
  XOR U34911 ( .A(n26209), .B(n26208), .Z(n26206) );
  XOR U34912 ( .A(y[4568]), .B(x[4568]), .Z(n26208) );
  XOR U34913 ( .A(y[4567]), .B(x[4567]), .Z(n26209) );
  XOR U34914 ( .A(y[4566]), .B(x[4566]), .Z(n26207) );
  XOR U34915 ( .A(n26201), .B(n26200), .Z(n26211) );
  XOR U34916 ( .A(n26203), .B(n26202), .Z(n26200) );
  XOR U34917 ( .A(y[4565]), .B(x[4565]), .Z(n26202) );
  XOR U34918 ( .A(y[4564]), .B(x[4564]), .Z(n26203) );
  XOR U34919 ( .A(y[4563]), .B(x[4563]), .Z(n26201) );
  XNOR U34920 ( .A(n26177), .B(n26178), .Z(n26195) );
  XNOR U34921 ( .A(n26192), .B(n26193), .Z(n26178) );
  XOR U34922 ( .A(n26189), .B(n26188), .Z(n26193) );
  XOR U34923 ( .A(y[4560]), .B(x[4560]), .Z(n26188) );
  XOR U34924 ( .A(n26191), .B(n26190), .Z(n26189) );
  XOR U34925 ( .A(y[4562]), .B(x[4562]), .Z(n26190) );
  XOR U34926 ( .A(y[4561]), .B(x[4561]), .Z(n26191) );
  XOR U34927 ( .A(n26183), .B(n26182), .Z(n26192) );
  XOR U34928 ( .A(n26185), .B(n26184), .Z(n26182) );
  XOR U34929 ( .A(y[4559]), .B(x[4559]), .Z(n26184) );
  XOR U34930 ( .A(y[4558]), .B(x[4558]), .Z(n26185) );
  XOR U34931 ( .A(y[4557]), .B(x[4557]), .Z(n26183) );
  XNOR U34932 ( .A(n26176), .B(n26175), .Z(n26177) );
  XNOR U34933 ( .A(n26172), .B(n26171), .Z(n26175) );
  XOR U34934 ( .A(n26174), .B(n26173), .Z(n26171) );
  XOR U34935 ( .A(y[4556]), .B(x[4556]), .Z(n26173) );
  XOR U34936 ( .A(y[4555]), .B(x[4555]), .Z(n26174) );
  XOR U34937 ( .A(y[4554]), .B(x[4554]), .Z(n26172) );
  XOR U34938 ( .A(n26166), .B(n26165), .Z(n26176) );
  XOR U34939 ( .A(n26168), .B(n26167), .Z(n26165) );
  XOR U34940 ( .A(y[4553]), .B(x[4553]), .Z(n26167) );
  XOR U34941 ( .A(y[4552]), .B(x[4552]), .Z(n26168) );
  XOR U34942 ( .A(y[4551]), .B(x[4551]), .Z(n26166) );
  NAND U34943 ( .A(n26229), .B(n26230), .Z(N63053) );
  NAND U34944 ( .A(n26231), .B(n26232), .Z(n26230) );
  NANDN U34945 ( .A(n26233), .B(n26234), .Z(n26232) );
  NANDN U34946 ( .A(n26234), .B(n26233), .Z(n26229) );
  XOR U34947 ( .A(n26233), .B(n26235), .Z(N63052) );
  XNOR U34948 ( .A(n26231), .B(n26234), .Z(n26235) );
  NAND U34949 ( .A(n26236), .B(n26237), .Z(n26234) );
  NAND U34950 ( .A(n26238), .B(n26239), .Z(n26237) );
  NANDN U34951 ( .A(n26240), .B(n26241), .Z(n26239) );
  NANDN U34952 ( .A(n26241), .B(n26240), .Z(n26236) );
  AND U34953 ( .A(n26242), .B(n26243), .Z(n26231) );
  NAND U34954 ( .A(n26244), .B(n26245), .Z(n26243) );
  NANDN U34955 ( .A(n26246), .B(n26247), .Z(n26245) );
  NANDN U34956 ( .A(n26247), .B(n26246), .Z(n26242) );
  IV U34957 ( .A(n26248), .Z(n26247) );
  AND U34958 ( .A(n26249), .B(n26250), .Z(n26233) );
  NAND U34959 ( .A(n26251), .B(n26252), .Z(n26250) );
  NANDN U34960 ( .A(n26253), .B(n26254), .Z(n26252) );
  NANDN U34961 ( .A(n26254), .B(n26253), .Z(n26249) );
  XOR U34962 ( .A(n26246), .B(n26255), .Z(N63051) );
  XNOR U34963 ( .A(n26244), .B(n26248), .Z(n26255) );
  XOR U34964 ( .A(n26241), .B(n26256), .Z(n26248) );
  XNOR U34965 ( .A(n26238), .B(n26240), .Z(n26256) );
  AND U34966 ( .A(n26257), .B(n26258), .Z(n26240) );
  NANDN U34967 ( .A(n26259), .B(n26260), .Z(n26258) );
  OR U34968 ( .A(n26261), .B(n26262), .Z(n26260) );
  IV U34969 ( .A(n26263), .Z(n26262) );
  NANDN U34970 ( .A(n26263), .B(n26261), .Z(n26257) );
  AND U34971 ( .A(n26264), .B(n26265), .Z(n26238) );
  NAND U34972 ( .A(n26266), .B(n26267), .Z(n26265) );
  NANDN U34973 ( .A(n26268), .B(n26269), .Z(n26267) );
  NANDN U34974 ( .A(n26269), .B(n26268), .Z(n26264) );
  IV U34975 ( .A(n26270), .Z(n26269) );
  NAND U34976 ( .A(n26271), .B(n26272), .Z(n26241) );
  NANDN U34977 ( .A(n26273), .B(n26274), .Z(n26272) );
  NANDN U34978 ( .A(n26275), .B(n26276), .Z(n26274) );
  NANDN U34979 ( .A(n26276), .B(n26275), .Z(n26271) );
  IV U34980 ( .A(n26277), .Z(n26275) );
  AND U34981 ( .A(n26278), .B(n26279), .Z(n26244) );
  NAND U34982 ( .A(n26280), .B(n26281), .Z(n26279) );
  NANDN U34983 ( .A(n26282), .B(n26283), .Z(n26281) );
  NANDN U34984 ( .A(n26283), .B(n26282), .Z(n26278) );
  XOR U34985 ( .A(n26254), .B(n26284), .Z(n26246) );
  XNOR U34986 ( .A(n26251), .B(n26253), .Z(n26284) );
  AND U34987 ( .A(n26285), .B(n26286), .Z(n26253) );
  NANDN U34988 ( .A(n26287), .B(n26288), .Z(n26286) );
  OR U34989 ( .A(n26289), .B(n26290), .Z(n26288) );
  IV U34990 ( .A(n26291), .Z(n26290) );
  NANDN U34991 ( .A(n26291), .B(n26289), .Z(n26285) );
  AND U34992 ( .A(n26292), .B(n26293), .Z(n26251) );
  NAND U34993 ( .A(n26294), .B(n26295), .Z(n26293) );
  NANDN U34994 ( .A(n26296), .B(n26297), .Z(n26295) );
  NANDN U34995 ( .A(n26297), .B(n26296), .Z(n26292) );
  IV U34996 ( .A(n26298), .Z(n26297) );
  NAND U34997 ( .A(n26299), .B(n26300), .Z(n26254) );
  NANDN U34998 ( .A(n26301), .B(n26302), .Z(n26300) );
  NANDN U34999 ( .A(n26303), .B(n26304), .Z(n26302) );
  NANDN U35000 ( .A(n26304), .B(n26303), .Z(n26299) );
  IV U35001 ( .A(n26305), .Z(n26303) );
  XOR U35002 ( .A(n26280), .B(n26306), .Z(N63050) );
  XNOR U35003 ( .A(n26283), .B(n26282), .Z(n26306) );
  XNOR U35004 ( .A(n26294), .B(n26307), .Z(n26282) );
  XNOR U35005 ( .A(n26298), .B(n26296), .Z(n26307) );
  XOR U35006 ( .A(n26304), .B(n26308), .Z(n26296) );
  XNOR U35007 ( .A(n26301), .B(n26305), .Z(n26308) );
  AND U35008 ( .A(n26309), .B(n26310), .Z(n26305) );
  NAND U35009 ( .A(n26311), .B(n26312), .Z(n26310) );
  NAND U35010 ( .A(n26313), .B(n26314), .Z(n26309) );
  AND U35011 ( .A(n26315), .B(n26316), .Z(n26301) );
  NAND U35012 ( .A(n26317), .B(n26318), .Z(n26316) );
  NAND U35013 ( .A(n26319), .B(n26320), .Z(n26315) );
  NANDN U35014 ( .A(n26321), .B(n26322), .Z(n26304) );
  ANDN U35015 ( .B(n26323), .A(n26324), .Z(n26298) );
  XNOR U35016 ( .A(n26289), .B(n26325), .Z(n26294) );
  XNOR U35017 ( .A(n26287), .B(n26291), .Z(n26325) );
  AND U35018 ( .A(n26326), .B(n26327), .Z(n26291) );
  NAND U35019 ( .A(n26328), .B(n26329), .Z(n26327) );
  NAND U35020 ( .A(n26330), .B(n26331), .Z(n26326) );
  AND U35021 ( .A(n26332), .B(n26333), .Z(n26287) );
  NAND U35022 ( .A(n26334), .B(n26335), .Z(n26333) );
  NAND U35023 ( .A(n26336), .B(n26337), .Z(n26332) );
  AND U35024 ( .A(n26338), .B(n26339), .Z(n26289) );
  NAND U35025 ( .A(n26340), .B(n26341), .Z(n26283) );
  XNOR U35026 ( .A(n26266), .B(n26342), .Z(n26280) );
  XNOR U35027 ( .A(n26270), .B(n26268), .Z(n26342) );
  XOR U35028 ( .A(n26276), .B(n26343), .Z(n26268) );
  XNOR U35029 ( .A(n26273), .B(n26277), .Z(n26343) );
  AND U35030 ( .A(n26344), .B(n26345), .Z(n26277) );
  NAND U35031 ( .A(n26346), .B(n26347), .Z(n26345) );
  NAND U35032 ( .A(n26348), .B(n26349), .Z(n26344) );
  AND U35033 ( .A(n26350), .B(n26351), .Z(n26273) );
  NAND U35034 ( .A(n26352), .B(n26353), .Z(n26351) );
  NAND U35035 ( .A(n26354), .B(n26355), .Z(n26350) );
  NANDN U35036 ( .A(n26356), .B(n26357), .Z(n26276) );
  ANDN U35037 ( .B(n26358), .A(n26359), .Z(n26270) );
  XNOR U35038 ( .A(n26261), .B(n26360), .Z(n26266) );
  XNOR U35039 ( .A(n26259), .B(n26263), .Z(n26360) );
  AND U35040 ( .A(n26361), .B(n26362), .Z(n26263) );
  NAND U35041 ( .A(n26363), .B(n26364), .Z(n26362) );
  NAND U35042 ( .A(n26365), .B(n26366), .Z(n26361) );
  AND U35043 ( .A(n26367), .B(n26368), .Z(n26259) );
  NAND U35044 ( .A(n26369), .B(n26370), .Z(n26368) );
  NAND U35045 ( .A(n26371), .B(n26372), .Z(n26367) );
  AND U35046 ( .A(n26373), .B(n26374), .Z(n26261) );
  XOR U35047 ( .A(n26341), .B(n26340), .Z(N63049) );
  XNOR U35048 ( .A(n26358), .B(n26359), .Z(n26340) );
  XNOR U35049 ( .A(n26373), .B(n26374), .Z(n26359) );
  XOR U35050 ( .A(n26370), .B(n26369), .Z(n26374) );
  XOR U35051 ( .A(y[4548]), .B(x[4548]), .Z(n26369) );
  XOR U35052 ( .A(n26372), .B(n26371), .Z(n26370) );
  XOR U35053 ( .A(y[4550]), .B(x[4550]), .Z(n26371) );
  XOR U35054 ( .A(y[4549]), .B(x[4549]), .Z(n26372) );
  XOR U35055 ( .A(n26364), .B(n26363), .Z(n26373) );
  XOR U35056 ( .A(n26366), .B(n26365), .Z(n26363) );
  XOR U35057 ( .A(y[4547]), .B(x[4547]), .Z(n26365) );
  XOR U35058 ( .A(y[4546]), .B(x[4546]), .Z(n26366) );
  XOR U35059 ( .A(y[4545]), .B(x[4545]), .Z(n26364) );
  XNOR U35060 ( .A(n26357), .B(n26356), .Z(n26358) );
  XNOR U35061 ( .A(n26353), .B(n26352), .Z(n26356) );
  XOR U35062 ( .A(n26355), .B(n26354), .Z(n26352) );
  XOR U35063 ( .A(y[4544]), .B(x[4544]), .Z(n26354) );
  XOR U35064 ( .A(y[4543]), .B(x[4543]), .Z(n26355) );
  XOR U35065 ( .A(y[4542]), .B(x[4542]), .Z(n26353) );
  XOR U35066 ( .A(n26347), .B(n26346), .Z(n26357) );
  XOR U35067 ( .A(n26349), .B(n26348), .Z(n26346) );
  XOR U35068 ( .A(y[4541]), .B(x[4541]), .Z(n26348) );
  XOR U35069 ( .A(y[4540]), .B(x[4540]), .Z(n26349) );
  XOR U35070 ( .A(y[4539]), .B(x[4539]), .Z(n26347) );
  XNOR U35071 ( .A(n26323), .B(n26324), .Z(n26341) );
  XNOR U35072 ( .A(n26338), .B(n26339), .Z(n26324) );
  XOR U35073 ( .A(n26335), .B(n26334), .Z(n26339) );
  XOR U35074 ( .A(y[4536]), .B(x[4536]), .Z(n26334) );
  XOR U35075 ( .A(n26337), .B(n26336), .Z(n26335) );
  XOR U35076 ( .A(y[4538]), .B(x[4538]), .Z(n26336) );
  XOR U35077 ( .A(y[4537]), .B(x[4537]), .Z(n26337) );
  XOR U35078 ( .A(n26329), .B(n26328), .Z(n26338) );
  XOR U35079 ( .A(n26331), .B(n26330), .Z(n26328) );
  XOR U35080 ( .A(y[4535]), .B(x[4535]), .Z(n26330) );
  XOR U35081 ( .A(y[4534]), .B(x[4534]), .Z(n26331) );
  XOR U35082 ( .A(y[4533]), .B(x[4533]), .Z(n26329) );
  XNOR U35083 ( .A(n26322), .B(n26321), .Z(n26323) );
  XNOR U35084 ( .A(n26318), .B(n26317), .Z(n26321) );
  XOR U35085 ( .A(n26320), .B(n26319), .Z(n26317) );
  XOR U35086 ( .A(y[4532]), .B(x[4532]), .Z(n26319) );
  XOR U35087 ( .A(y[4531]), .B(x[4531]), .Z(n26320) );
  XOR U35088 ( .A(y[4530]), .B(x[4530]), .Z(n26318) );
  XOR U35089 ( .A(n26312), .B(n26311), .Z(n26322) );
  XOR U35090 ( .A(n26314), .B(n26313), .Z(n26311) );
  XOR U35091 ( .A(y[4529]), .B(x[4529]), .Z(n26313) );
  XOR U35092 ( .A(y[4528]), .B(x[4528]), .Z(n26314) );
  XOR U35093 ( .A(y[4527]), .B(x[4527]), .Z(n26312) );
  NAND U35094 ( .A(n26375), .B(n26376), .Z(N63040) );
  NAND U35095 ( .A(n26377), .B(n26378), .Z(n26376) );
  NANDN U35096 ( .A(n26379), .B(n26380), .Z(n26378) );
  NANDN U35097 ( .A(n26380), .B(n26379), .Z(n26375) );
  XOR U35098 ( .A(n26379), .B(n26381), .Z(N63039) );
  XNOR U35099 ( .A(n26377), .B(n26380), .Z(n26381) );
  NAND U35100 ( .A(n26382), .B(n26383), .Z(n26380) );
  NAND U35101 ( .A(n26384), .B(n26385), .Z(n26383) );
  NANDN U35102 ( .A(n26386), .B(n26387), .Z(n26385) );
  NANDN U35103 ( .A(n26387), .B(n26386), .Z(n26382) );
  AND U35104 ( .A(n26388), .B(n26389), .Z(n26377) );
  NAND U35105 ( .A(n26390), .B(n26391), .Z(n26389) );
  NANDN U35106 ( .A(n26392), .B(n26393), .Z(n26391) );
  NANDN U35107 ( .A(n26393), .B(n26392), .Z(n26388) );
  IV U35108 ( .A(n26394), .Z(n26393) );
  AND U35109 ( .A(n26395), .B(n26396), .Z(n26379) );
  NAND U35110 ( .A(n26397), .B(n26398), .Z(n26396) );
  NANDN U35111 ( .A(n26399), .B(n26400), .Z(n26398) );
  NANDN U35112 ( .A(n26400), .B(n26399), .Z(n26395) );
  XOR U35113 ( .A(n26392), .B(n26401), .Z(N63038) );
  XNOR U35114 ( .A(n26390), .B(n26394), .Z(n26401) );
  XOR U35115 ( .A(n26387), .B(n26402), .Z(n26394) );
  XNOR U35116 ( .A(n26384), .B(n26386), .Z(n26402) );
  AND U35117 ( .A(n26403), .B(n26404), .Z(n26386) );
  NANDN U35118 ( .A(n26405), .B(n26406), .Z(n26404) );
  OR U35119 ( .A(n26407), .B(n26408), .Z(n26406) );
  IV U35120 ( .A(n26409), .Z(n26408) );
  NANDN U35121 ( .A(n26409), .B(n26407), .Z(n26403) );
  AND U35122 ( .A(n26410), .B(n26411), .Z(n26384) );
  NAND U35123 ( .A(n26412), .B(n26413), .Z(n26411) );
  NANDN U35124 ( .A(n26414), .B(n26415), .Z(n26413) );
  NANDN U35125 ( .A(n26415), .B(n26414), .Z(n26410) );
  IV U35126 ( .A(n26416), .Z(n26415) );
  NAND U35127 ( .A(n26417), .B(n26418), .Z(n26387) );
  NANDN U35128 ( .A(n26419), .B(n26420), .Z(n26418) );
  NANDN U35129 ( .A(n26421), .B(n26422), .Z(n26420) );
  NANDN U35130 ( .A(n26422), .B(n26421), .Z(n26417) );
  IV U35131 ( .A(n26423), .Z(n26421) );
  AND U35132 ( .A(n26424), .B(n26425), .Z(n26390) );
  NAND U35133 ( .A(n26426), .B(n26427), .Z(n26425) );
  NANDN U35134 ( .A(n26428), .B(n26429), .Z(n26427) );
  NANDN U35135 ( .A(n26429), .B(n26428), .Z(n26424) );
  XOR U35136 ( .A(n26400), .B(n26430), .Z(n26392) );
  XNOR U35137 ( .A(n26397), .B(n26399), .Z(n26430) );
  AND U35138 ( .A(n26431), .B(n26432), .Z(n26399) );
  NANDN U35139 ( .A(n26433), .B(n26434), .Z(n26432) );
  OR U35140 ( .A(n26435), .B(n26436), .Z(n26434) );
  IV U35141 ( .A(n26437), .Z(n26436) );
  NANDN U35142 ( .A(n26437), .B(n26435), .Z(n26431) );
  AND U35143 ( .A(n26438), .B(n26439), .Z(n26397) );
  NAND U35144 ( .A(n26440), .B(n26441), .Z(n26439) );
  NANDN U35145 ( .A(n26442), .B(n26443), .Z(n26441) );
  NANDN U35146 ( .A(n26443), .B(n26442), .Z(n26438) );
  IV U35147 ( .A(n26444), .Z(n26443) );
  NAND U35148 ( .A(n26445), .B(n26446), .Z(n26400) );
  NANDN U35149 ( .A(n26447), .B(n26448), .Z(n26446) );
  NANDN U35150 ( .A(n26449), .B(n26450), .Z(n26448) );
  NANDN U35151 ( .A(n26450), .B(n26449), .Z(n26445) );
  IV U35152 ( .A(n26451), .Z(n26449) );
  XOR U35153 ( .A(n26426), .B(n26452), .Z(N63037) );
  XNOR U35154 ( .A(n26429), .B(n26428), .Z(n26452) );
  XNOR U35155 ( .A(n26440), .B(n26453), .Z(n26428) );
  XNOR U35156 ( .A(n26444), .B(n26442), .Z(n26453) );
  XOR U35157 ( .A(n26450), .B(n26454), .Z(n26442) );
  XNOR U35158 ( .A(n26447), .B(n26451), .Z(n26454) );
  AND U35159 ( .A(n26455), .B(n26456), .Z(n26451) );
  NAND U35160 ( .A(n26457), .B(n26458), .Z(n26456) );
  NAND U35161 ( .A(n26459), .B(n26460), .Z(n26455) );
  AND U35162 ( .A(n26461), .B(n26462), .Z(n26447) );
  NAND U35163 ( .A(n26463), .B(n26464), .Z(n26462) );
  NAND U35164 ( .A(n26465), .B(n26466), .Z(n26461) );
  NANDN U35165 ( .A(n26467), .B(n26468), .Z(n26450) );
  ANDN U35166 ( .B(n26469), .A(n26470), .Z(n26444) );
  XNOR U35167 ( .A(n26435), .B(n26471), .Z(n26440) );
  XNOR U35168 ( .A(n26433), .B(n26437), .Z(n26471) );
  AND U35169 ( .A(n26472), .B(n26473), .Z(n26437) );
  NAND U35170 ( .A(n26474), .B(n26475), .Z(n26473) );
  NAND U35171 ( .A(n26476), .B(n26477), .Z(n26472) );
  AND U35172 ( .A(n26478), .B(n26479), .Z(n26433) );
  NAND U35173 ( .A(n26480), .B(n26481), .Z(n26479) );
  NAND U35174 ( .A(n26482), .B(n26483), .Z(n26478) );
  AND U35175 ( .A(n26484), .B(n26485), .Z(n26435) );
  NAND U35176 ( .A(n26486), .B(n26487), .Z(n26429) );
  XNOR U35177 ( .A(n26412), .B(n26488), .Z(n26426) );
  XNOR U35178 ( .A(n26416), .B(n26414), .Z(n26488) );
  XOR U35179 ( .A(n26422), .B(n26489), .Z(n26414) );
  XNOR U35180 ( .A(n26419), .B(n26423), .Z(n26489) );
  AND U35181 ( .A(n26490), .B(n26491), .Z(n26423) );
  NAND U35182 ( .A(n26492), .B(n26493), .Z(n26491) );
  NAND U35183 ( .A(n26494), .B(n26495), .Z(n26490) );
  AND U35184 ( .A(n26496), .B(n26497), .Z(n26419) );
  NAND U35185 ( .A(n26498), .B(n26499), .Z(n26497) );
  NAND U35186 ( .A(n26500), .B(n26501), .Z(n26496) );
  NANDN U35187 ( .A(n26502), .B(n26503), .Z(n26422) );
  ANDN U35188 ( .B(n26504), .A(n26505), .Z(n26416) );
  XNOR U35189 ( .A(n26407), .B(n26506), .Z(n26412) );
  XNOR U35190 ( .A(n26405), .B(n26409), .Z(n26506) );
  AND U35191 ( .A(n26507), .B(n26508), .Z(n26409) );
  NAND U35192 ( .A(n26509), .B(n26510), .Z(n26508) );
  NAND U35193 ( .A(n26511), .B(n26512), .Z(n26507) );
  AND U35194 ( .A(n26513), .B(n26514), .Z(n26405) );
  NAND U35195 ( .A(n26515), .B(n26516), .Z(n26514) );
  NAND U35196 ( .A(n26517), .B(n26518), .Z(n26513) );
  AND U35197 ( .A(n26519), .B(n26520), .Z(n26407) );
  XOR U35198 ( .A(n26487), .B(n26486), .Z(N63036) );
  XNOR U35199 ( .A(n26504), .B(n26505), .Z(n26486) );
  XNOR U35200 ( .A(n26519), .B(n26520), .Z(n26505) );
  XOR U35201 ( .A(n26516), .B(n26515), .Z(n26520) );
  XOR U35202 ( .A(y[4524]), .B(x[4524]), .Z(n26515) );
  XOR U35203 ( .A(n26518), .B(n26517), .Z(n26516) );
  XOR U35204 ( .A(y[4526]), .B(x[4526]), .Z(n26517) );
  XOR U35205 ( .A(y[4525]), .B(x[4525]), .Z(n26518) );
  XOR U35206 ( .A(n26510), .B(n26509), .Z(n26519) );
  XOR U35207 ( .A(n26512), .B(n26511), .Z(n26509) );
  XOR U35208 ( .A(y[4523]), .B(x[4523]), .Z(n26511) );
  XOR U35209 ( .A(y[4522]), .B(x[4522]), .Z(n26512) );
  XOR U35210 ( .A(y[4521]), .B(x[4521]), .Z(n26510) );
  XNOR U35211 ( .A(n26503), .B(n26502), .Z(n26504) );
  XNOR U35212 ( .A(n26499), .B(n26498), .Z(n26502) );
  XOR U35213 ( .A(n26501), .B(n26500), .Z(n26498) );
  XOR U35214 ( .A(y[4520]), .B(x[4520]), .Z(n26500) );
  XOR U35215 ( .A(y[4519]), .B(x[4519]), .Z(n26501) );
  XOR U35216 ( .A(y[4518]), .B(x[4518]), .Z(n26499) );
  XOR U35217 ( .A(n26493), .B(n26492), .Z(n26503) );
  XOR U35218 ( .A(n26495), .B(n26494), .Z(n26492) );
  XOR U35219 ( .A(y[4517]), .B(x[4517]), .Z(n26494) );
  XOR U35220 ( .A(y[4516]), .B(x[4516]), .Z(n26495) );
  XOR U35221 ( .A(y[4515]), .B(x[4515]), .Z(n26493) );
  XNOR U35222 ( .A(n26469), .B(n26470), .Z(n26487) );
  XNOR U35223 ( .A(n26484), .B(n26485), .Z(n26470) );
  XOR U35224 ( .A(n26481), .B(n26480), .Z(n26485) );
  XOR U35225 ( .A(y[4512]), .B(x[4512]), .Z(n26480) );
  XOR U35226 ( .A(n26483), .B(n26482), .Z(n26481) );
  XOR U35227 ( .A(y[4514]), .B(x[4514]), .Z(n26482) );
  XOR U35228 ( .A(y[4513]), .B(x[4513]), .Z(n26483) );
  XOR U35229 ( .A(n26475), .B(n26474), .Z(n26484) );
  XOR U35230 ( .A(n26477), .B(n26476), .Z(n26474) );
  XOR U35231 ( .A(y[4511]), .B(x[4511]), .Z(n26476) );
  XOR U35232 ( .A(y[4510]), .B(x[4510]), .Z(n26477) );
  XOR U35233 ( .A(y[4509]), .B(x[4509]), .Z(n26475) );
  XNOR U35234 ( .A(n26468), .B(n26467), .Z(n26469) );
  XNOR U35235 ( .A(n26464), .B(n26463), .Z(n26467) );
  XOR U35236 ( .A(n26466), .B(n26465), .Z(n26463) );
  XOR U35237 ( .A(y[4508]), .B(x[4508]), .Z(n26465) );
  XOR U35238 ( .A(y[4507]), .B(x[4507]), .Z(n26466) );
  XOR U35239 ( .A(y[4506]), .B(x[4506]), .Z(n26464) );
  XOR U35240 ( .A(n26458), .B(n26457), .Z(n26468) );
  XOR U35241 ( .A(n26460), .B(n26459), .Z(n26457) );
  XOR U35242 ( .A(y[4505]), .B(x[4505]), .Z(n26459) );
  XOR U35243 ( .A(y[4504]), .B(x[4504]), .Z(n26460) );
  XOR U35244 ( .A(y[4503]), .B(x[4503]), .Z(n26458) );
  NAND U35245 ( .A(n26521), .B(n26522), .Z(N63027) );
  NAND U35246 ( .A(n26523), .B(n26524), .Z(n26522) );
  NANDN U35247 ( .A(n26525), .B(n26526), .Z(n26524) );
  NANDN U35248 ( .A(n26526), .B(n26525), .Z(n26521) );
  XOR U35249 ( .A(n26525), .B(n26527), .Z(N63026) );
  XNOR U35250 ( .A(n26523), .B(n26526), .Z(n26527) );
  NAND U35251 ( .A(n26528), .B(n26529), .Z(n26526) );
  NAND U35252 ( .A(n26530), .B(n26531), .Z(n26529) );
  NANDN U35253 ( .A(n26532), .B(n26533), .Z(n26531) );
  NANDN U35254 ( .A(n26533), .B(n26532), .Z(n26528) );
  AND U35255 ( .A(n26534), .B(n26535), .Z(n26523) );
  NAND U35256 ( .A(n26536), .B(n26537), .Z(n26535) );
  NANDN U35257 ( .A(n26538), .B(n26539), .Z(n26537) );
  NANDN U35258 ( .A(n26539), .B(n26538), .Z(n26534) );
  IV U35259 ( .A(n26540), .Z(n26539) );
  AND U35260 ( .A(n26541), .B(n26542), .Z(n26525) );
  NAND U35261 ( .A(n26543), .B(n26544), .Z(n26542) );
  NANDN U35262 ( .A(n26545), .B(n26546), .Z(n26544) );
  NANDN U35263 ( .A(n26546), .B(n26545), .Z(n26541) );
  XOR U35264 ( .A(n26538), .B(n26547), .Z(N63025) );
  XNOR U35265 ( .A(n26536), .B(n26540), .Z(n26547) );
  XOR U35266 ( .A(n26533), .B(n26548), .Z(n26540) );
  XNOR U35267 ( .A(n26530), .B(n26532), .Z(n26548) );
  AND U35268 ( .A(n26549), .B(n26550), .Z(n26532) );
  NANDN U35269 ( .A(n26551), .B(n26552), .Z(n26550) );
  OR U35270 ( .A(n26553), .B(n26554), .Z(n26552) );
  IV U35271 ( .A(n26555), .Z(n26554) );
  NANDN U35272 ( .A(n26555), .B(n26553), .Z(n26549) );
  AND U35273 ( .A(n26556), .B(n26557), .Z(n26530) );
  NAND U35274 ( .A(n26558), .B(n26559), .Z(n26557) );
  NANDN U35275 ( .A(n26560), .B(n26561), .Z(n26559) );
  NANDN U35276 ( .A(n26561), .B(n26560), .Z(n26556) );
  IV U35277 ( .A(n26562), .Z(n26561) );
  NAND U35278 ( .A(n26563), .B(n26564), .Z(n26533) );
  NANDN U35279 ( .A(n26565), .B(n26566), .Z(n26564) );
  NANDN U35280 ( .A(n26567), .B(n26568), .Z(n26566) );
  NANDN U35281 ( .A(n26568), .B(n26567), .Z(n26563) );
  IV U35282 ( .A(n26569), .Z(n26567) );
  AND U35283 ( .A(n26570), .B(n26571), .Z(n26536) );
  NAND U35284 ( .A(n26572), .B(n26573), .Z(n26571) );
  NANDN U35285 ( .A(n26574), .B(n26575), .Z(n26573) );
  NANDN U35286 ( .A(n26575), .B(n26574), .Z(n26570) );
  XOR U35287 ( .A(n26546), .B(n26576), .Z(n26538) );
  XNOR U35288 ( .A(n26543), .B(n26545), .Z(n26576) );
  AND U35289 ( .A(n26577), .B(n26578), .Z(n26545) );
  NANDN U35290 ( .A(n26579), .B(n26580), .Z(n26578) );
  OR U35291 ( .A(n26581), .B(n26582), .Z(n26580) );
  IV U35292 ( .A(n26583), .Z(n26582) );
  NANDN U35293 ( .A(n26583), .B(n26581), .Z(n26577) );
  AND U35294 ( .A(n26584), .B(n26585), .Z(n26543) );
  NAND U35295 ( .A(n26586), .B(n26587), .Z(n26585) );
  NANDN U35296 ( .A(n26588), .B(n26589), .Z(n26587) );
  NANDN U35297 ( .A(n26589), .B(n26588), .Z(n26584) );
  IV U35298 ( .A(n26590), .Z(n26589) );
  NAND U35299 ( .A(n26591), .B(n26592), .Z(n26546) );
  NANDN U35300 ( .A(n26593), .B(n26594), .Z(n26592) );
  NANDN U35301 ( .A(n26595), .B(n26596), .Z(n26594) );
  NANDN U35302 ( .A(n26596), .B(n26595), .Z(n26591) );
  IV U35303 ( .A(n26597), .Z(n26595) );
  XOR U35304 ( .A(n26572), .B(n26598), .Z(N63024) );
  XNOR U35305 ( .A(n26575), .B(n26574), .Z(n26598) );
  XNOR U35306 ( .A(n26586), .B(n26599), .Z(n26574) );
  XNOR U35307 ( .A(n26590), .B(n26588), .Z(n26599) );
  XOR U35308 ( .A(n26596), .B(n26600), .Z(n26588) );
  XNOR U35309 ( .A(n26593), .B(n26597), .Z(n26600) );
  AND U35310 ( .A(n26601), .B(n26602), .Z(n26597) );
  NAND U35311 ( .A(n26603), .B(n26604), .Z(n26602) );
  NAND U35312 ( .A(n26605), .B(n26606), .Z(n26601) );
  AND U35313 ( .A(n26607), .B(n26608), .Z(n26593) );
  NAND U35314 ( .A(n26609), .B(n26610), .Z(n26608) );
  NAND U35315 ( .A(n26611), .B(n26612), .Z(n26607) );
  NANDN U35316 ( .A(n26613), .B(n26614), .Z(n26596) );
  ANDN U35317 ( .B(n26615), .A(n26616), .Z(n26590) );
  XNOR U35318 ( .A(n26581), .B(n26617), .Z(n26586) );
  XNOR U35319 ( .A(n26579), .B(n26583), .Z(n26617) );
  AND U35320 ( .A(n26618), .B(n26619), .Z(n26583) );
  NAND U35321 ( .A(n26620), .B(n26621), .Z(n26619) );
  NAND U35322 ( .A(n26622), .B(n26623), .Z(n26618) );
  AND U35323 ( .A(n26624), .B(n26625), .Z(n26579) );
  NAND U35324 ( .A(n26626), .B(n26627), .Z(n26625) );
  NAND U35325 ( .A(n26628), .B(n26629), .Z(n26624) );
  AND U35326 ( .A(n26630), .B(n26631), .Z(n26581) );
  NAND U35327 ( .A(n26632), .B(n26633), .Z(n26575) );
  XNOR U35328 ( .A(n26558), .B(n26634), .Z(n26572) );
  XNOR U35329 ( .A(n26562), .B(n26560), .Z(n26634) );
  XOR U35330 ( .A(n26568), .B(n26635), .Z(n26560) );
  XNOR U35331 ( .A(n26565), .B(n26569), .Z(n26635) );
  AND U35332 ( .A(n26636), .B(n26637), .Z(n26569) );
  NAND U35333 ( .A(n26638), .B(n26639), .Z(n26637) );
  NAND U35334 ( .A(n26640), .B(n26641), .Z(n26636) );
  AND U35335 ( .A(n26642), .B(n26643), .Z(n26565) );
  NAND U35336 ( .A(n26644), .B(n26645), .Z(n26643) );
  NAND U35337 ( .A(n26646), .B(n26647), .Z(n26642) );
  NANDN U35338 ( .A(n26648), .B(n26649), .Z(n26568) );
  ANDN U35339 ( .B(n26650), .A(n26651), .Z(n26562) );
  XNOR U35340 ( .A(n26553), .B(n26652), .Z(n26558) );
  XNOR U35341 ( .A(n26551), .B(n26555), .Z(n26652) );
  AND U35342 ( .A(n26653), .B(n26654), .Z(n26555) );
  NAND U35343 ( .A(n26655), .B(n26656), .Z(n26654) );
  NAND U35344 ( .A(n26657), .B(n26658), .Z(n26653) );
  AND U35345 ( .A(n26659), .B(n26660), .Z(n26551) );
  NAND U35346 ( .A(n26661), .B(n26662), .Z(n26660) );
  NAND U35347 ( .A(n26663), .B(n26664), .Z(n26659) );
  AND U35348 ( .A(n26665), .B(n26666), .Z(n26553) );
  XOR U35349 ( .A(n26633), .B(n26632), .Z(N63023) );
  XNOR U35350 ( .A(n26650), .B(n26651), .Z(n26632) );
  XNOR U35351 ( .A(n26665), .B(n26666), .Z(n26651) );
  XOR U35352 ( .A(n26662), .B(n26661), .Z(n26666) );
  XOR U35353 ( .A(y[4500]), .B(x[4500]), .Z(n26661) );
  XOR U35354 ( .A(n26664), .B(n26663), .Z(n26662) );
  XOR U35355 ( .A(y[4502]), .B(x[4502]), .Z(n26663) );
  XOR U35356 ( .A(y[4501]), .B(x[4501]), .Z(n26664) );
  XOR U35357 ( .A(n26656), .B(n26655), .Z(n26665) );
  XOR U35358 ( .A(n26658), .B(n26657), .Z(n26655) );
  XOR U35359 ( .A(y[4499]), .B(x[4499]), .Z(n26657) );
  XOR U35360 ( .A(y[4498]), .B(x[4498]), .Z(n26658) );
  XOR U35361 ( .A(y[4497]), .B(x[4497]), .Z(n26656) );
  XNOR U35362 ( .A(n26649), .B(n26648), .Z(n26650) );
  XNOR U35363 ( .A(n26645), .B(n26644), .Z(n26648) );
  XOR U35364 ( .A(n26647), .B(n26646), .Z(n26644) );
  XOR U35365 ( .A(y[4496]), .B(x[4496]), .Z(n26646) );
  XOR U35366 ( .A(y[4495]), .B(x[4495]), .Z(n26647) );
  XOR U35367 ( .A(y[4494]), .B(x[4494]), .Z(n26645) );
  XOR U35368 ( .A(n26639), .B(n26638), .Z(n26649) );
  XOR U35369 ( .A(n26641), .B(n26640), .Z(n26638) );
  XOR U35370 ( .A(y[4493]), .B(x[4493]), .Z(n26640) );
  XOR U35371 ( .A(y[4492]), .B(x[4492]), .Z(n26641) );
  XOR U35372 ( .A(y[4491]), .B(x[4491]), .Z(n26639) );
  XNOR U35373 ( .A(n26615), .B(n26616), .Z(n26633) );
  XNOR U35374 ( .A(n26630), .B(n26631), .Z(n26616) );
  XOR U35375 ( .A(n26627), .B(n26626), .Z(n26631) );
  XOR U35376 ( .A(y[4488]), .B(x[4488]), .Z(n26626) );
  XOR U35377 ( .A(n26629), .B(n26628), .Z(n26627) );
  XOR U35378 ( .A(y[4490]), .B(x[4490]), .Z(n26628) );
  XOR U35379 ( .A(y[4489]), .B(x[4489]), .Z(n26629) );
  XOR U35380 ( .A(n26621), .B(n26620), .Z(n26630) );
  XOR U35381 ( .A(n26623), .B(n26622), .Z(n26620) );
  XOR U35382 ( .A(y[4487]), .B(x[4487]), .Z(n26622) );
  XOR U35383 ( .A(y[4486]), .B(x[4486]), .Z(n26623) );
  XOR U35384 ( .A(y[4485]), .B(x[4485]), .Z(n26621) );
  XNOR U35385 ( .A(n26614), .B(n26613), .Z(n26615) );
  XNOR U35386 ( .A(n26610), .B(n26609), .Z(n26613) );
  XOR U35387 ( .A(n26612), .B(n26611), .Z(n26609) );
  XOR U35388 ( .A(y[4484]), .B(x[4484]), .Z(n26611) );
  XOR U35389 ( .A(y[4483]), .B(x[4483]), .Z(n26612) );
  XOR U35390 ( .A(y[4482]), .B(x[4482]), .Z(n26610) );
  XOR U35391 ( .A(n26604), .B(n26603), .Z(n26614) );
  XOR U35392 ( .A(n26606), .B(n26605), .Z(n26603) );
  XOR U35393 ( .A(y[4481]), .B(x[4481]), .Z(n26605) );
  XOR U35394 ( .A(y[4480]), .B(x[4480]), .Z(n26606) );
  XOR U35395 ( .A(y[4479]), .B(x[4479]), .Z(n26604) );
  NAND U35396 ( .A(n26667), .B(n26668), .Z(N63014) );
  NAND U35397 ( .A(n26669), .B(n26670), .Z(n26668) );
  NANDN U35398 ( .A(n26671), .B(n26672), .Z(n26670) );
  NANDN U35399 ( .A(n26672), .B(n26671), .Z(n26667) );
  XOR U35400 ( .A(n26671), .B(n26673), .Z(N63013) );
  XNOR U35401 ( .A(n26669), .B(n26672), .Z(n26673) );
  NAND U35402 ( .A(n26674), .B(n26675), .Z(n26672) );
  NAND U35403 ( .A(n26676), .B(n26677), .Z(n26675) );
  NANDN U35404 ( .A(n26678), .B(n26679), .Z(n26677) );
  NANDN U35405 ( .A(n26679), .B(n26678), .Z(n26674) );
  AND U35406 ( .A(n26680), .B(n26681), .Z(n26669) );
  NAND U35407 ( .A(n26682), .B(n26683), .Z(n26681) );
  NANDN U35408 ( .A(n26684), .B(n26685), .Z(n26683) );
  NANDN U35409 ( .A(n26685), .B(n26684), .Z(n26680) );
  IV U35410 ( .A(n26686), .Z(n26685) );
  AND U35411 ( .A(n26687), .B(n26688), .Z(n26671) );
  NAND U35412 ( .A(n26689), .B(n26690), .Z(n26688) );
  NANDN U35413 ( .A(n26691), .B(n26692), .Z(n26690) );
  NANDN U35414 ( .A(n26692), .B(n26691), .Z(n26687) );
  XOR U35415 ( .A(n26684), .B(n26693), .Z(N63012) );
  XNOR U35416 ( .A(n26682), .B(n26686), .Z(n26693) );
  XOR U35417 ( .A(n26679), .B(n26694), .Z(n26686) );
  XNOR U35418 ( .A(n26676), .B(n26678), .Z(n26694) );
  AND U35419 ( .A(n26695), .B(n26696), .Z(n26678) );
  NANDN U35420 ( .A(n26697), .B(n26698), .Z(n26696) );
  OR U35421 ( .A(n26699), .B(n26700), .Z(n26698) );
  IV U35422 ( .A(n26701), .Z(n26700) );
  NANDN U35423 ( .A(n26701), .B(n26699), .Z(n26695) );
  AND U35424 ( .A(n26702), .B(n26703), .Z(n26676) );
  NAND U35425 ( .A(n26704), .B(n26705), .Z(n26703) );
  NANDN U35426 ( .A(n26706), .B(n26707), .Z(n26705) );
  NANDN U35427 ( .A(n26707), .B(n26706), .Z(n26702) );
  IV U35428 ( .A(n26708), .Z(n26707) );
  NAND U35429 ( .A(n26709), .B(n26710), .Z(n26679) );
  NANDN U35430 ( .A(n26711), .B(n26712), .Z(n26710) );
  NANDN U35431 ( .A(n26713), .B(n26714), .Z(n26712) );
  NANDN U35432 ( .A(n26714), .B(n26713), .Z(n26709) );
  IV U35433 ( .A(n26715), .Z(n26713) );
  AND U35434 ( .A(n26716), .B(n26717), .Z(n26682) );
  NAND U35435 ( .A(n26718), .B(n26719), .Z(n26717) );
  NANDN U35436 ( .A(n26720), .B(n26721), .Z(n26719) );
  NANDN U35437 ( .A(n26721), .B(n26720), .Z(n26716) );
  XOR U35438 ( .A(n26692), .B(n26722), .Z(n26684) );
  XNOR U35439 ( .A(n26689), .B(n26691), .Z(n26722) );
  AND U35440 ( .A(n26723), .B(n26724), .Z(n26691) );
  NANDN U35441 ( .A(n26725), .B(n26726), .Z(n26724) );
  OR U35442 ( .A(n26727), .B(n26728), .Z(n26726) );
  IV U35443 ( .A(n26729), .Z(n26728) );
  NANDN U35444 ( .A(n26729), .B(n26727), .Z(n26723) );
  AND U35445 ( .A(n26730), .B(n26731), .Z(n26689) );
  NAND U35446 ( .A(n26732), .B(n26733), .Z(n26731) );
  NANDN U35447 ( .A(n26734), .B(n26735), .Z(n26733) );
  NANDN U35448 ( .A(n26735), .B(n26734), .Z(n26730) );
  IV U35449 ( .A(n26736), .Z(n26735) );
  NAND U35450 ( .A(n26737), .B(n26738), .Z(n26692) );
  NANDN U35451 ( .A(n26739), .B(n26740), .Z(n26738) );
  NANDN U35452 ( .A(n26741), .B(n26742), .Z(n26740) );
  NANDN U35453 ( .A(n26742), .B(n26741), .Z(n26737) );
  IV U35454 ( .A(n26743), .Z(n26741) );
  XOR U35455 ( .A(n26718), .B(n26744), .Z(N63011) );
  XNOR U35456 ( .A(n26721), .B(n26720), .Z(n26744) );
  XNOR U35457 ( .A(n26732), .B(n26745), .Z(n26720) );
  XNOR U35458 ( .A(n26736), .B(n26734), .Z(n26745) );
  XOR U35459 ( .A(n26742), .B(n26746), .Z(n26734) );
  XNOR U35460 ( .A(n26739), .B(n26743), .Z(n26746) );
  AND U35461 ( .A(n26747), .B(n26748), .Z(n26743) );
  NAND U35462 ( .A(n26749), .B(n26750), .Z(n26748) );
  NAND U35463 ( .A(n26751), .B(n26752), .Z(n26747) );
  AND U35464 ( .A(n26753), .B(n26754), .Z(n26739) );
  NAND U35465 ( .A(n26755), .B(n26756), .Z(n26754) );
  NAND U35466 ( .A(n26757), .B(n26758), .Z(n26753) );
  NANDN U35467 ( .A(n26759), .B(n26760), .Z(n26742) );
  ANDN U35468 ( .B(n26761), .A(n26762), .Z(n26736) );
  XNOR U35469 ( .A(n26727), .B(n26763), .Z(n26732) );
  XNOR U35470 ( .A(n26725), .B(n26729), .Z(n26763) );
  AND U35471 ( .A(n26764), .B(n26765), .Z(n26729) );
  NAND U35472 ( .A(n26766), .B(n26767), .Z(n26765) );
  NAND U35473 ( .A(n26768), .B(n26769), .Z(n26764) );
  AND U35474 ( .A(n26770), .B(n26771), .Z(n26725) );
  NAND U35475 ( .A(n26772), .B(n26773), .Z(n26771) );
  NAND U35476 ( .A(n26774), .B(n26775), .Z(n26770) );
  AND U35477 ( .A(n26776), .B(n26777), .Z(n26727) );
  NAND U35478 ( .A(n26778), .B(n26779), .Z(n26721) );
  XNOR U35479 ( .A(n26704), .B(n26780), .Z(n26718) );
  XNOR U35480 ( .A(n26708), .B(n26706), .Z(n26780) );
  XOR U35481 ( .A(n26714), .B(n26781), .Z(n26706) );
  XNOR U35482 ( .A(n26711), .B(n26715), .Z(n26781) );
  AND U35483 ( .A(n26782), .B(n26783), .Z(n26715) );
  NAND U35484 ( .A(n26784), .B(n26785), .Z(n26783) );
  NAND U35485 ( .A(n26786), .B(n26787), .Z(n26782) );
  AND U35486 ( .A(n26788), .B(n26789), .Z(n26711) );
  NAND U35487 ( .A(n26790), .B(n26791), .Z(n26789) );
  NAND U35488 ( .A(n26792), .B(n26793), .Z(n26788) );
  NANDN U35489 ( .A(n26794), .B(n26795), .Z(n26714) );
  ANDN U35490 ( .B(n26796), .A(n26797), .Z(n26708) );
  XNOR U35491 ( .A(n26699), .B(n26798), .Z(n26704) );
  XNOR U35492 ( .A(n26697), .B(n26701), .Z(n26798) );
  AND U35493 ( .A(n26799), .B(n26800), .Z(n26701) );
  NAND U35494 ( .A(n26801), .B(n26802), .Z(n26800) );
  NAND U35495 ( .A(n26803), .B(n26804), .Z(n26799) );
  AND U35496 ( .A(n26805), .B(n26806), .Z(n26697) );
  NAND U35497 ( .A(n26807), .B(n26808), .Z(n26806) );
  NAND U35498 ( .A(n26809), .B(n26810), .Z(n26805) );
  AND U35499 ( .A(n26811), .B(n26812), .Z(n26699) );
  XOR U35500 ( .A(n26779), .B(n26778), .Z(N63010) );
  XNOR U35501 ( .A(n26796), .B(n26797), .Z(n26778) );
  XNOR U35502 ( .A(n26811), .B(n26812), .Z(n26797) );
  XOR U35503 ( .A(n26808), .B(n26807), .Z(n26812) );
  XOR U35504 ( .A(y[4476]), .B(x[4476]), .Z(n26807) );
  XOR U35505 ( .A(n26810), .B(n26809), .Z(n26808) );
  XOR U35506 ( .A(y[4478]), .B(x[4478]), .Z(n26809) );
  XOR U35507 ( .A(y[4477]), .B(x[4477]), .Z(n26810) );
  XOR U35508 ( .A(n26802), .B(n26801), .Z(n26811) );
  XOR U35509 ( .A(n26804), .B(n26803), .Z(n26801) );
  XOR U35510 ( .A(y[4475]), .B(x[4475]), .Z(n26803) );
  XOR U35511 ( .A(y[4474]), .B(x[4474]), .Z(n26804) );
  XOR U35512 ( .A(y[4473]), .B(x[4473]), .Z(n26802) );
  XNOR U35513 ( .A(n26795), .B(n26794), .Z(n26796) );
  XNOR U35514 ( .A(n26791), .B(n26790), .Z(n26794) );
  XOR U35515 ( .A(n26793), .B(n26792), .Z(n26790) );
  XOR U35516 ( .A(y[4472]), .B(x[4472]), .Z(n26792) );
  XOR U35517 ( .A(y[4471]), .B(x[4471]), .Z(n26793) );
  XOR U35518 ( .A(y[4470]), .B(x[4470]), .Z(n26791) );
  XOR U35519 ( .A(n26785), .B(n26784), .Z(n26795) );
  XOR U35520 ( .A(n26787), .B(n26786), .Z(n26784) );
  XOR U35521 ( .A(y[4469]), .B(x[4469]), .Z(n26786) );
  XOR U35522 ( .A(y[4468]), .B(x[4468]), .Z(n26787) );
  XOR U35523 ( .A(y[4467]), .B(x[4467]), .Z(n26785) );
  XNOR U35524 ( .A(n26761), .B(n26762), .Z(n26779) );
  XNOR U35525 ( .A(n26776), .B(n26777), .Z(n26762) );
  XOR U35526 ( .A(n26773), .B(n26772), .Z(n26777) );
  XOR U35527 ( .A(y[4464]), .B(x[4464]), .Z(n26772) );
  XOR U35528 ( .A(n26775), .B(n26774), .Z(n26773) );
  XOR U35529 ( .A(y[4466]), .B(x[4466]), .Z(n26774) );
  XOR U35530 ( .A(y[4465]), .B(x[4465]), .Z(n26775) );
  XOR U35531 ( .A(n26767), .B(n26766), .Z(n26776) );
  XOR U35532 ( .A(n26769), .B(n26768), .Z(n26766) );
  XOR U35533 ( .A(y[4463]), .B(x[4463]), .Z(n26768) );
  XOR U35534 ( .A(y[4462]), .B(x[4462]), .Z(n26769) );
  XOR U35535 ( .A(y[4461]), .B(x[4461]), .Z(n26767) );
  XNOR U35536 ( .A(n26760), .B(n26759), .Z(n26761) );
  XNOR U35537 ( .A(n26756), .B(n26755), .Z(n26759) );
  XOR U35538 ( .A(n26758), .B(n26757), .Z(n26755) );
  XOR U35539 ( .A(y[4460]), .B(x[4460]), .Z(n26757) );
  XOR U35540 ( .A(y[4459]), .B(x[4459]), .Z(n26758) );
  XOR U35541 ( .A(y[4458]), .B(x[4458]), .Z(n26756) );
  XOR U35542 ( .A(n26750), .B(n26749), .Z(n26760) );
  XOR U35543 ( .A(n26752), .B(n26751), .Z(n26749) );
  XOR U35544 ( .A(y[4457]), .B(x[4457]), .Z(n26751) );
  XOR U35545 ( .A(y[4456]), .B(x[4456]), .Z(n26752) );
  XOR U35546 ( .A(y[4455]), .B(x[4455]), .Z(n26750) );
  NAND U35547 ( .A(n26813), .B(n26814), .Z(N63001) );
  NAND U35548 ( .A(n26815), .B(n26816), .Z(n26814) );
  NANDN U35549 ( .A(n26817), .B(n26818), .Z(n26816) );
  NANDN U35550 ( .A(n26818), .B(n26817), .Z(n26813) );
  XOR U35551 ( .A(n26817), .B(n26819), .Z(N63000) );
  XNOR U35552 ( .A(n26815), .B(n26818), .Z(n26819) );
  NAND U35553 ( .A(n26820), .B(n26821), .Z(n26818) );
  NAND U35554 ( .A(n26822), .B(n26823), .Z(n26821) );
  NANDN U35555 ( .A(n26824), .B(n26825), .Z(n26823) );
  NANDN U35556 ( .A(n26825), .B(n26824), .Z(n26820) );
  AND U35557 ( .A(n26826), .B(n26827), .Z(n26815) );
  NAND U35558 ( .A(n26828), .B(n26829), .Z(n26827) );
  NANDN U35559 ( .A(n26830), .B(n26831), .Z(n26829) );
  NANDN U35560 ( .A(n26831), .B(n26830), .Z(n26826) );
  IV U35561 ( .A(n26832), .Z(n26831) );
  AND U35562 ( .A(n26833), .B(n26834), .Z(n26817) );
  NAND U35563 ( .A(n26835), .B(n26836), .Z(n26834) );
  NANDN U35564 ( .A(n26837), .B(n26838), .Z(n26836) );
  NANDN U35565 ( .A(n26838), .B(n26837), .Z(n26833) );
  XOR U35566 ( .A(n26830), .B(n26839), .Z(N62999) );
  XNOR U35567 ( .A(n26828), .B(n26832), .Z(n26839) );
  XOR U35568 ( .A(n26825), .B(n26840), .Z(n26832) );
  XNOR U35569 ( .A(n26822), .B(n26824), .Z(n26840) );
  AND U35570 ( .A(n26841), .B(n26842), .Z(n26824) );
  NANDN U35571 ( .A(n26843), .B(n26844), .Z(n26842) );
  OR U35572 ( .A(n26845), .B(n26846), .Z(n26844) );
  IV U35573 ( .A(n26847), .Z(n26846) );
  NANDN U35574 ( .A(n26847), .B(n26845), .Z(n26841) );
  AND U35575 ( .A(n26848), .B(n26849), .Z(n26822) );
  NAND U35576 ( .A(n26850), .B(n26851), .Z(n26849) );
  NANDN U35577 ( .A(n26852), .B(n26853), .Z(n26851) );
  NANDN U35578 ( .A(n26853), .B(n26852), .Z(n26848) );
  IV U35579 ( .A(n26854), .Z(n26853) );
  NAND U35580 ( .A(n26855), .B(n26856), .Z(n26825) );
  NANDN U35581 ( .A(n26857), .B(n26858), .Z(n26856) );
  NANDN U35582 ( .A(n26859), .B(n26860), .Z(n26858) );
  NANDN U35583 ( .A(n26860), .B(n26859), .Z(n26855) );
  IV U35584 ( .A(n26861), .Z(n26859) );
  AND U35585 ( .A(n26862), .B(n26863), .Z(n26828) );
  NAND U35586 ( .A(n26864), .B(n26865), .Z(n26863) );
  NANDN U35587 ( .A(n26866), .B(n26867), .Z(n26865) );
  NANDN U35588 ( .A(n26867), .B(n26866), .Z(n26862) );
  XOR U35589 ( .A(n26838), .B(n26868), .Z(n26830) );
  XNOR U35590 ( .A(n26835), .B(n26837), .Z(n26868) );
  AND U35591 ( .A(n26869), .B(n26870), .Z(n26837) );
  NANDN U35592 ( .A(n26871), .B(n26872), .Z(n26870) );
  OR U35593 ( .A(n26873), .B(n26874), .Z(n26872) );
  IV U35594 ( .A(n26875), .Z(n26874) );
  NANDN U35595 ( .A(n26875), .B(n26873), .Z(n26869) );
  AND U35596 ( .A(n26876), .B(n26877), .Z(n26835) );
  NAND U35597 ( .A(n26878), .B(n26879), .Z(n26877) );
  NANDN U35598 ( .A(n26880), .B(n26881), .Z(n26879) );
  NANDN U35599 ( .A(n26881), .B(n26880), .Z(n26876) );
  IV U35600 ( .A(n26882), .Z(n26881) );
  NAND U35601 ( .A(n26883), .B(n26884), .Z(n26838) );
  NANDN U35602 ( .A(n26885), .B(n26886), .Z(n26884) );
  NANDN U35603 ( .A(n26887), .B(n26888), .Z(n26886) );
  NANDN U35604 ( .A(n26888), .B(n26887), .Z(n26883) );
  IV U35605 ( .A(n26889), .Z(n26887) );
  XOR U35606 ( .A(n26864), .B(n26890), .Z(N62998) );
  XNOR U35607 ( .A(n26867), .B(n26866), .Z(n26890) );
  XNOR U35608 ( .A(n26878), .B(n26891), .Z(n26866) );
  XNOR U35609 ( .A(n26882), .B(n26880), .Z(n26891) );
  XOR U35610 ( .A(n26888), .B(n26892), .Z(n26880) );
  XNOR U35611 ( .A(n26885), .B(n26889), .Z(n26892) );
  AND U35612 ( .A(n26893), .B(n26894), .Z(n26889) );
  NAND U35613 ( .A(n26895), .B(n26896), .Z(n26894) );
  NAND U35614 ( .A(n26897), .B(n26898), .Z(n26893) );
  AND U35615 ( .A(n26899), .B(n26900), .Z(n26885) );
  NAND U35616 ( .A(n26901), .B(n26902), .Z(n26900) );
  NAND U35617 ( .A(n26903), .B(n26904), .Z(n26899) );
  NANDN U35618 ( .A(n26905), .B(n26906), .Z(n26888) );
  ANDN U35619 ( .B(n26907), .A(n26908), .Z(n26882) );
  XNOR U35620 ( .A(n26873), .B(n26909), .Z(n26878) );
  XNOR U35621 ( .A(n26871), .B(n26875), .Z(n26909) );
  AND U35622 ( .A(n26910), .B(n26911), .Z(n26875) );
  NAND U35623 ( .A(n26912), .B(n26913), .Z(n26911) );
  NAND U35624 ( .A(n26914), .B(n26915), .Z(n26910) );
  AND U35625 ( .A(n26916), .B(n26917), .Z(n26871) );
  NAND U35626 ( .A(n26918), .B(n26919), .Z(n26917) );
  NAND U35627 ( .A(n26920), .B(n26921), .Z(n26916) );
  AND U35628 ( .A(n26922), .B(n26923), .Z(n26873) );
  NAND U35629 ( .A(n26924), .B(n26925), .Z(n26867) );
  XNOR U35630 ( .A(n26850), .B(n26926), .Z(n26864) );
  XNOR U35631 ( .A(n26854), .B(n26852), .Z(n26926) );
  XOR U35632 ( .A(n26860), .B(n26927), .Z(n26852) );
  XNOR U35633 ( .A(n26857), .B(n26861), .Z(n26927) );
  AND U35634 ( .A(n26928), .B(n26929), .Z(n26861) );
  NAND U35635 ( .A(n26930), .B(n26931), .Z(n26929) );
  NAND U35636 ( .A(n26932), .B(n26933), .Z(n26928) );
  AND U35637 ( .A(n26934), .B(n26935), .Z(n26857) );
  NAND U35638 ( .A(n26936), .B(n26937), .Z(n26935) );
  NAND U35639 ( .A(n26938), .B(n26939), .Z(n26934) );
  NANDN U35640 ( .A(n26940), .B(n26941), .Z(n26860) );
  ANDN U35641 ( .B(n26942), .A(n26943), .Z(n26854) );
  XNOR U35642 ( .A(n26845), .B(n26944), .Z(n26850) );
  XNOR U35643 ( .A(n26843), .B(n26847), .Z(n26944) );
  AND U35644 ( .A(n26945), .B(n26946), .Z(n26847) );
  NAND U35645 ( .A(n26947), .B(n26948), .Z(n26946) );
  NAND U35646 ( .A(n26949), .B(n26950), .Z(n26945) );
  AND U35647 ( .A(n26951), .B(n26952), .Z(n26843) );
  NAND U35648 ( .A(n26953), .B(n26954), .Z(n26952) );
  NAND U35649 ( .A(n26955), .B(n26956), .Z(n26951) );
  AND U35650 ( .A(n26957), .B(n26958), .Z(n26845) );
  XOR U35651 ( .A(n26925), .B(n26924), .Z(N62997) );
  XNOR U35652 ( .A(n26942), .B(n26943), .Z(n26924) );
  XNOR U35653 ( .A(n26957), .B(n26958), .Z(n26943) );
  XOR U35654 ( .A(n26954), .B(n26953), .Z(n26958) );
  XOR U35655 ( .A(y[4452]), .B(x[4452]), .Z(n26953) );
  XOR U35656 ( .A(n26956), .B(n26955), .Z(n26954) );
  XOR U35657 ( .A(y[4454]), .B(x[4454]), .Z(n26955) );
  XOR U35658 ( .A(y[4453]), .B(x[4453]), .Z(n26956) );
  XOR U35659 ( .A(n26948), .B(n26947), .Z(n26957) );
  XOR U35660 ( .A(n26950), .B(n26949), .Z(n26947) );
  XOR U35661 ( .A(y[4451]), .B(x[4451]), .Z(n26949) );
  XOR U35662 ( .A(y[4450]), .B(x[4450]), .Z(n26950) );
  XOR U35663 ( .A(y[4449]), .B(x[4449]), .Z(n26948) );
  XNOR U35664 ( .A(n26941), .B(n26940), .Z(n26942) );
  XNOR U35665 ( .A(n26937), .B(n26936), .Z(n26940) );
  XOR U35666 ( .A(n26939), .B(n26938), .Z(n26936) );
  XOR U35667 ( .A(y[4448]), .B(x[4448]), .Z(n26938) );
  XOR U35668 ( .A(y[4447]), .B(x[4447]), .Z(n26939) );
  XOR U35669 ( .A(y[4446]), .B(x[4446]), .Z(n26937) );
  XOR U35670 ( .A(n26931), .B(n26930), .Z(n26941) );
  XOR U35671 ( .A(n26933), .B(n26932), .Z(n26930) );
  XOR U35672 ( .A(y[4445]), .B(x[4445]), .Z(n26932) );
  XOR U35673 ( .A(y[4444]), .B(x[4444]), .Z(n26933) );
  XOR U35674 ( .A(y[4443]), .B(x[4443]), .Z(n26931) );
  XNOR U35675 ( .A(n26907), .B(n26908), .Z(n26925) );
  XNOR U35676 ( .A(n26922), .B(n26923), .Z(n26908) );
  XOR U35677 ( .A(n26919), .B(n26918), .Z(n26923) );
  XOR U35678 ( .A(y[4440]), .B(x[4440]), .Z(n26918) );
  XOR U35679 ( .A(n26921), .B(n26920), .Z(n26919) );
  XOR U35680 ( .A(y[4442]), .B(x[4442]), .Z(n26920) );
  XOR U35681 ( .A(y[4441]), .B(x[4441]), .Z(n26921) );
  XOR U35682 ( .A(n26913), .B(n26912), .Z(n26922) );
  XOR U35683 ( .A(n26915), .B(n26914), .Z(n26912) );
  XOR U35684 ( .A(y[4439]), .B(x[4439]), .Z(n26914) );
  XOR U35685 ( .A(y[4438]), .B(x[4438]), .Z(n26915) );
  XOR U35686 ( .A(y[4437]), .B(x[4437]), .Z(n26913) );
  XNOR U35687 ( .A(n26906), .B(n26905), .Z(n26907) );
  XNOR U35688 ( .A(n26902), .B(n26901), .Z(n26905) );
  XOR U35689 ( .A(n26904), .B(n26903), .Z(n26901) );
  XOR U35690 ( .A(y[4436]), .B(x[4436]), .Z(n26903) );
  XOR U35691 ( .A(y[4435]), .B(x[4435]), .Z(n26904) );
  XOR U35692 ( .A(y[4434]), .B(x[4434]), .Z(n26902) );
  XOR U35693 ( .A(n26896), .B(n26895), .Z(n26906) );
  XOR U35694 ( .A(n26898), .B(n26897), .Z(n26895) );
  XOR U35695 ( .A(y[4433]), .B(x[4433]), .Z(n26897) );
  XOR U35696 ( .A(y[4432]), .B(x[4432]), .Z(n26898) );
  XOR U35697 ( .A(y[4431]), .B(x[4431]), .Z(n26896) );
  NAND U35698 ( .A(n26959), .B(n26960), .Z(N62988) );
  NAND U35699 ( .A(n26961), .B(n26962), .Z(n26960) );
  NANDN U35700 ( .A(n26963), .B(n26964), .Z(n26962) );
  NANDN U35701 ( .A(n26964), .B(n26963), .Z(n26959) );
  XOR U35702 ( .A(n26963), .B(n26965), .Z(N62987) );
  XNOR U35703 ( .A(n26961), .B(n26964), .Z(n26965) );
  NAND U35704 ( .A(n26966), .B(n26967), .Z(n26964) );
  NAND U35705 ( .A(n26968), .B(n26969), .Z(n26967) );
  NANDN U35706 ( .A(n26970), .B(n26971), .Z(n26969) );
  NANDN U35707 ( .A(n26971), .B(n26970), .Z(n26966) );
  AND U35708 ( .A(n26972), .B(n26973), .Z(n26961) );
  NAND U35709 ( .A(n26974), .B(n26975), .Z(n26973) );
  NANDN U35710 ( .A(n26976), .B(n26977), .Z(n26975) );
  NANDN U35711 ( .A(n26977), .B(n26976), .Z(n26972) );
  IV U35712 ( .A(n26978), .Z(n26977) );
  AND U35713 ( .A(n26979), .B(n26980), .Z(n26963) );
  NAND U35714 ( .A(n26981), .B(n26982), .Z(n26980) );
  NANDN U35715 ( .A(n26983), .B(n26984), .Z(n26982) );
  NANDN U35716 ( .A(n26984), .B(n26983), .Z(n26979) );
  XOR U35717 ( .A(n26976), .B(n26985), .Z(N62986) );
  XNOR U35718 ( .A(n26974), .B(n26978), .Z(n26985) );
  XOR U35719 ( .A(n26971), .B(n26986), .Z(n26978) );
  XNOR U35720 ( .A(n26968), .B(n26970), .Z(n26986) );
  AND U35721 ( .A(n26987), .B(n26988), .Z(n26970) );
  NANDN U35722 ( .A(n26989), .B(n26990), .Z(n26988) );
  OR U35723 ( .A(n26991), .B(n26992), .Z(n26990) );
  IV U35724 ( .A(n26993), .Z(n26992) );
  NANDN U35725 ( .A(n26993), .B(n26991), .Z(n26987) );
  AND U35726 ( .A(n26994), .B(n26995), .Z(n26968) );
  NAND U35727 ( .A(n26996), .B(n26997), .Z(n26995) );
  NANDN U35728 ( .A(n26998), .B(n26999), .Z(n26997) );
  NANDN U35729 ( .A(n26999), .B(n26998), .Z(n26994) );
  IV U35730 ( .A(n27000), .Z(n26999) );
  NAND U35731 ( .A(n27001), .B(n27002), .Z(n26971) );
  NANDN U35732 ( .A(n27003), .B(n27004), .Z(n27002) );
  NANDN U35733 ( .A(n27005), .B(n27006), .Z(n27004) );
  NANDN U35734 ( .A(n27006), .B(n27005), .Z(n27001) );
  IV U35735 ( .A(n27007), .Z(n27005) );
  AND U35736 ( .A(n27008), .B(n27009), .Z(n26974) );
  NAND U35737 ( .A(n27010), .B(n27011), .Z(n27009) );
  NANDN U35738 ( .A(n27012), .B(n27013), .Z(n27011) );
  NANDN U35739 ( .A(n27013), .B(n27012), .Z(n27008) );
  XOR U35740 ( .A(n26984), .B(n27014), .Z(n26976) );
  XNOR U35741 ( .A(n26981), .B(n26983), .Z(n27014) );
  AND U35742 ( .A(n27015), .B(n27016), .Z(n26983) );
  NANDN U35743 ( .A(n27017), .B(n27018), .Z(n27016) );
  OR U35744 ( .A(n27019), .B(n27020), .Z(n27018) );
  IV U35745 ( .A(n27021), .Z(n27020) );
  NANDN U35746 ( .A(n27021), .B(n27019), .Z(n27015) );
  AND U35747 ( .A(n27022), .B(n27023), .Z(n26981) );
  NAND U35748 ( .A(n27024), .B(n27025), .Z(n27023) );
  NANDN U35749 ( .A(n27026), .B(n27027), .Z(n27025) );
  NANDN U35750 ( .A(n27027), .B(n27026), .Z(n27022) );
  IV U35751 ( .A(n27028), .Z(n27027) );
  NAND U35752 ( .A(n27029), .B(n27030), .Z(n26984) );
  NANDN U35753 ( .A(n27031), .B(n27032), .Z(n27030) );
  NANDN U35754 ( .A(n27033), .B(n27034), .Z(n27032) );
  NANDN U35755 ( .A(n27034), .B(n27033), .Z(n27029) );
  IV U35756 ( .A(n27035), .Z(n27033) );
  XOR U35757 ( .A(n27010), .B(n27036), .Z(N62985) );
  XNOR U35758 ( .A(n27013), .B(n27012), .Z(n27036) );
  XNOR U35759 ( .A(n27024), .B(n27037), .Z(n27012) );
  XNOR U35760 ( .A(n27028), .B(n27026), .Z(n27037) );
  XOR U35761 ( .A(n27034), .B(n27038), .Z(n27026) );
  XNOR U35762 ( .A(n27031), .B(n27035), .Z(n27038) );
  AND U35763 ( .A(n27039), .B(n27040), .Z(n27035) );
  NAND U35764 ( .A(n27041), .B(n27042), .Z(n27040) );
  NAND U35765 ( .A(n27043), .B(n27044), .Z(n27039) );
  AND U35766 ( .A(n27045), .B(n27046), .Z(n27031) );
  NAND U35767 ( .A(n27047), .B(n27048), .Z(n27046) );
  NAND U35768 ( .A(n27049), .B(n27050), .Z(n27045) );
  NANDN U35769 ( .A(n27051), .B(n27052), .Z(n27034) );
  ANDN U35770 ( .B(n27053), .A(n27054), .Z(n27028) );
  XNOR U35771 ( .A(n27019), .B(n27055), .Z(n27024) );
  XNOR U35772 ( .A(n27017), .B(n27021), .Z(n27055) );
  AND U35773 ( .A(n27056), .B(n27057), .Z(n27021) );
  NAND U35774 ( .A(n27058), .B(n27059), .Z(n27057) );
  NAND U35775 ( .A(n27060), .B(n27061), .Z(n27056) );
  AND U35776 ( .A(n27062), .B(n27063), .Z(n27017) );
  NAND U35777 ( .A(n27064), .B(n27065), .Z(n27063) );
  NAND U35778 ( .A(n27066), .B(n27067), .Z(n27062) );
  AND U35779 ( .A(n27068), .B(n27069), .Z(n27019) );
  NAND U35780 ( .A(n27070), .B(n27071), .Z(n27013) );
  XNOR U35781 ( .A(n26996), .B(n27072), .Z(n27010) );
  XNOR U35782 ( .A(n27000), .B(n26998), .Z(n27072) );
  XOR U35783 ( .A(n27006), .B(n27073), .Z(n26998) );
  XNOR U35784 ( .A(n27003), .B(n27007), .Z(n27073) );
  AND U35785 ( .A(n27074), .B(n27075), .Z(n27007) );
  NAND U35786 ( .A(n27076), .B(n27077), .Z(n27075) );
  NAND U35787 ( .A(n27078), .B(n27079), .Z(n27074) );
  AND U35788 ( .A(n27080), .B(n27081), .Z(n27003) );
  NAND U35789 ( .A(n27082), .B(n27083), .Z(n27081) );
  NAND U35790 ( .A(n27084), .B(n27085), .Z(n27080) );
  NANDN U35791 ( .A(n27086), .B(n27087), .Z(n27006) );
  ANDN U35792 ( .B(n27088), .A(n27089), .Z(n27000) );
  XNOR U35793 ( .A(n26991), .B(n27090), .Z(n26996) );
  XNOR U35794 ( .A(n26989), .B(n26993), .Z(n27090) );
  AND U35795 ( .A(n27091), .B(n27092), .Z(n26993) );
  NAND U35796 ( .A(n27093), .B(n27094), .Z(n27092) );
  NAND U35797 ( .A(n27095), .B(n27096), .Z(n27091) );
  AND U35798 ( .A(n27097), .B(n27098), .Z(n26989) );
  NAND U35799 ( .A(n27099), .B(n27100), .Z(n27098) );
  NAND U35800 ( .A(n27101), .B(n27102), .Z(n27097) );
  AND U35801 ( .A(n27103), .B(n27104), .Z(n26991) );
  XOR U35802 ( .A(n27071), .B(n27070), .Z(N62984) );
  XNOR U35803 ( .A(n27088), .B(n27089), .Z(n27070) );
  XNOR U35804 ( .A(n27103), .B(n27104), .Z(n27089) );
  XOR U35805 ( .A(n27100), .B(n27099), .Z(n27104) );
  XOR U35806 ( .A(y[4428]), .B(x[4428]), .Z(n27099) );
  XOR U35807 ( .A(n27102), .B(n27101), .Z(n27100) );
  XOR U35808 ( .A(y[4430]), .B(x[4430]), .Z(n27101) );
  XOR U35809 ( .A(y[4429]), .B(x[4429]), .Z(n27102) );
  XOR U35810 ( .A(n27094), .B(n27093), .Z(n27103) );
  XOR U35811 ( .A(n27096), .B(n27095), .Z(n27093) );
  XOR U35812 ( .A(y[4427]), .B(x[4427]), .Z(n27095) );
  XOR U35813 ( .A(y[4426]), .B(x[4426]), .Z(n27096) );
  XOR U35814 ( .A(y[4425]), .B(x[4425]), .Z(n27094) );
  XNOR U35815 ( .A(n27087), .B(n27086), .Z(n27088) );
  XNOR U35816 ( .A(n27083), .B(n27082), .Z(n27086) );
  XOR U35817 ( .A(n27085), .B(n27084), .Z(n27082) );
  XOR U35818 ( .A(y[4424]), .B(x[4424]), .Z(n27084) );
  XOR U35819 ( .A(y[4423]), .B(x[4423]), .Z(n27085) );
  XOR U35820 ( .A(y[4422]), .B(x[4422]), .Z(n27083) );
  XOR U35821 ( .A(n27077), .B(n27076), .Z(n27087) );
  XOR U35822 ( .A(n27079), .B(n27078), .Z(n27076) );
  XOR U35823 ( .A(y[4421]), .B(x[4421]), .Z(n27078) );
  XOR U35824 ( .A(y[4420]), .B(x[4420]), .Z(n27079) );
  XOR U35825 ( .A(y[4419]), .B(x[4419]), .Z(n27077) );
  XNOR U35826 ( .A(n27053), .B(n27054), .Z(n27071) );
  XNOR U35827 ( .A(n27068), .B(n27069), .Z(n27054) );
  XOR U35828 ( .A(n27065), .B(n27064), .Z(n27069) );
  XOR U35829 ( .A(y[4416]), .B(x[4416]), .Z(n27064) );
  XOR U35830 ( .A(n27067), .B(n27066), .Z(n27065) );
  XOR U35831 ( .A(y[4418]), .B(x[4418]), .Z(n27066) );
  XOR U35832 ( .A(y[4417]), .B(x[4417]), .Z(n27067) );
  XOR U35833 ( .A(n27059), .B(n27058), .Z(n27068) );
  XOR U35834 ( .A(n27061), .B(n27060), .Z(n27058) );
  XOR U35835 ( .A(y[4415]), .B(x[4415]), .Z(n27060) );
  XOR U35836 ( .A(y[4414]), .B(x[4414]), .Z(n27061) );
  XOR U35837 ( .A(y[4413]), .B(x[4413]), .Z(n27059) );
  XNOR U35838 ( .A(n27052), .B(n27051), .Z(n27053) );
  XNOR U35839 ( .A(n27048), .B(n27047), .Z(n27051) );
  XOR U35840 ( .A(n27050), .B(n27049), .Z(n27047) );
  XOR U35841 ( .A(y[4412]), .B(x[4412]), .Z(n27049) );
  XOR U35842 ( .A(y[4411]), .B(x[4411]), .Z(n27050) );
  XOR U35843 ( .A(y[4410]), .B(x[4410]), .Z(n27048) );
  XOR U35844 ( .A(n27042), .B(n27041), .Z(n27052) );
  XOR U35845 ( .A(n27044), .B(n27043), .Z(n27041) );
  XOR U35846 ( .A(y[4409]), .B(x[4409]), .Z(n27043) );
  XOR U35847 ( .A(y[4408]), .B(x[4408]), .Z(n27044) );
  XOR U35848 ( .A(y[4407]), .B(x[4407]), .Z(n27042) );
  NAND U35849 ( .A(n27105), .B(n27106), .Z(N62975) );
  NAND U35850 ( .A(n27107), .B(n27108), .Z(n27106) );
  NANDN U35851 ( .A(n27109), .B(n27110), .Z(n27108) );
  NANDN U35852 ( .A(n27110), .B(n27109), .Z(n27105) );
  XOR U35853 ( .A(n27109), .B(n27111), .Z(N62974) );
  XNOR U35854 ( .A(n27107), .B(n27110), .Z(n27111) );
  NAND U35855 ( .A(n27112), .B(n27113), .Z(n27110) );
  NAND U35856 ( .A(n27114), .B(n27115), .Z(n27113) );
  NANDN U35857 ( .A(n27116), .B(n27117), .Z(n27115) );
  NANDN U35858 ( .A(n27117), .B(n27116), .Z(n27112) );
  AND U35859 ( .A(n27118), .B(n27119), .Z(n27107) );
  NAND U35860 ( .A(n27120), .B(n27121), .Z(n27119) );
  NANDN U35861 ( .A(n27122), .B(n27123), .Z(n27121) );
  NANDN U35862 ( .A(n27123), .B(n27122), .Z(n27118) );
  IV U35863 ( .A(n27124), .Z(n27123) );
  AND U35864 ( .A(n27125), .B(n27126), .Z(n27109) );
  NAND U35865 ( .A(n27127), .B(n27128), .Z(n27126) );
  NANDN U35866 ( .A(n27129), .B(n27130), .Z(n27128) );
  NANDN U35867 ( .A(n27130), .B(n27129), .Z(n27125) );
  XOR U35868 ( .A(n27122), .B(n27131), .Z(N62973) );
  XNOR U35869 ( .A(n27120), .B(n27124), .Z(n27131) );
  XOR U35870 ( .A(n27117), .B(n27132), .Z(n27124) );
  XNOR U35871 ( .A(n27114), .B(n27116), .Z(n27132) );
  AND U35872 ( .A(n27133), .B(n27134), .Z(n27116) );
  NANDN U35873 ( .A(n27135), .B(n27136), .Z(n27134) );
  OR U35874 ( .A(n27137), .B(n27138), .Z(n27136) );
  IV U35875 ( .A(n27139), .Z(n27138) );
  NANDN U35876 ( .A(n27139), .B(n27137), .Z(n27133) );
  AND U35877 ( .A(n27140), .B(n27141), .Z(n27114) );
  NAND U35878 ( .A(n27142), .B(n27143), .Z(n27141) );
  NANDN U35879 ( .A(n27144), .B(n27145), .Z(n27143) );
  NANDN U35880 ( .A(n27145), .B(n27144), .Z(n27140) );
  IV U35881 ( .A(n27146), .Z(n27145) );
  NAND U35882 ( .A(n27147), .B(n27148), .Z(n27117) );
  NANDN U35883 ( .A(n27149), .B(n27150), .Z(n27148) );
  NANDN U35884 ( .A(n27151), .B(n27152), .Z(n27150) );
  NANDN U35885 ( .A(n27152), .B(n27151), .Z(n27147) );
  IV U35886 ( .A(n27153), .Z(n27151) );
  AND U35887 ( .A(n27154), .B(n27155), .Z(n27120) );
  NAND U35888 ( .A(n27156), .B(n27157), .Z(n27155) );
  NANDN U35889 ( .A(n27158), .B(n27159), .Z(n27157) );
  NANDN U35890 ( .A(n27159), .B(n27158), .Z(n27154) );
  XOR U35891 ( .A(n27130), .B(n27160), .Z(n27122) );
  XNOR U35892 ( .A(n27127), .B(n27129), .Z(n27160) );
  AND U35893 ( .A(n27161), .B(n27162), .Z(n27129) );
  NANDN U35894 ( .A(n27163), .B(n27164), .Z(n27162) );
  OR U35895 ( .A(n27165), .B(n27166), .Z(n27164) );
  IV U35896 ( .A(n27167), .Z(n27166) );
  NANDN U35897 ( .A(n27167), .B(n27165), .Z(n27161) );
  AND U35898 ( .A(n27168), .B(n27169), .Z(n27127) );
  NAND U35899 ( .A(n27170), .B(n27171), .Z(n27169) );
  NANDN U35900 ( .A(n27172), .B(n27173), .Z(n27171) );
  NANDN U35901 ( .A(n27173), .B(n27172), .Z(n27168) );
  IV U35902 ( .A(n27174), .Z(n27173) );
  NAND U35903 ( .A(n27175), .B(n27176), .Z(n27130) );
  NANDN U35904 ( .A(n27177), .B(n27178), .Z(n27176) );
  NANDN U35905 ( .A(n27179), .B(n27180), .Z(n27178) );
  NANDN U35906 ( .A(n27180), .B(n27179), .Z(n27175) );
  IV U35907 ( .A(n27181), .Z(n27179) );
  XOR U35908 ( .A(n27156), .B(n27182), .Z(N62972) );
  XNOR U35909 ( .A(n27159), .B(n27158), .Z(n27182) );
  XNOR U35910 ( .A(n27170), .B(n27183), .Z(n27158) );
  XNOR U35911 ( .A(n27174), .B(n27172), .Z(n27183) );
  XOR U35912 ( .A(n27180), .B(n27184), .Z(n27172) );
  XNOR U35913 ( .A(n27177), .B(n27181), .Z(n27184) );
  AND U35914 ( .A(n27185), .B(n27186), .Z(n27181) );
  NAND U35915 ( .A(n27187), .B(n27188), .Z(n27186) );
  NAND U35916 ( .A(n27189), .B(n27190), .Z(n27185) );
  AND U35917 ( .A(n27191), .B(n27192), .Z(n27177) );
  NAND U35918 ( .A(n27193), .B(n27194), .Z(n27192) );
  NAND U35919 ( .A(n27195), .B(n27196), .Z(n27191) );
  NANDN U35920 ( .A(n27197), .B(n27198), .Z(n27180) );
  ANDN U35921 ( .B(n27199), .A(n27200), .Z(n27174) );
  XNOR U35922 ( .A(n27165), .B(n27201), .Z(n27170) );
  XNOR U35923 ( .A(n27163), .B(n27167), .Z(n27201) );
  AND U35924 ( .A(n27202), .B(n27203), .Z(n27167) );
  NAND U35925 ( .A(n27204), .B(n27205), .Z(n27203) );
  NAND U35926 ( .A(n27206), .B(n27207), .Z(n27202) );
  AND U35927 ( .A(n27208), .B(n27209), .Z(n27163) );
  NAND U35928 ( .A(n27210), .B(n27211), .Z(n27209) );
  NAND U35929 ( .A(n27212), .B(n27213), .Z(n27208) );
  AND U35930 ( .A(n27214), .B(n27215), .Z(n27165) );
  NAND U35931 ( .A(n27216), .B(n27217), .Z(n27159) );
  XNOR U35932 ( .A(n27142), .B(n27218), .Z(n27156) );
  XNOR U35933 ( .A(n27146), .B(n27144), .Z(n27218) );
  XOR U35934 ( .A(n27152), .B(n27219), .Z(n27144) );
  XNOR U35935 ( .A(n27149), .B(n27153), .Z(n27219) );
  AND U35936 ( .A(n27220), .B(n27221), .Z(n27153) );
  NAND U35937 ( .A(n27222), .B(n27223), .Z(n27221) );
  NAND U35938 ( .A(n27224), .B(n27225), .Z(n27220) );
  AND U35939 ( .A(n27226), .B(n27227), .Z(n27149) );
  NAND U35940 ( .A(n27228), .B(n27229), .Z(n27227) );
  NAND U35941 ( .A(n27230), .B(n27231), .Z(n27226) );
  NANDN U35942 ( .A(n27232), .B(n27233), .Z(n27152) );
  ANDN U35943 ( .B(n27234), .A(n27235), .Z(n27146) );
  XNOR U35944 ( .A(n27137), .B(n27236), .Z(n27142) );
  XNOR U35945 ( .A(n27135), .B(n27139), .Z(n27236) );
  AND U35946 ( .A(n27237), .B(n27238), .Z(n27139) );
  NAND U35947 ( .A(n27239), .B(n27240), .Z(n27238) );
  NAND U35948 ( .A(n27241), .B(n27242), .Z(n27237) );
  AND U35949 ( .A(n27243), .B(n27244), .Z(n27135) );
  NAND U35950 ( .A(n27245), .B(n27246), .Z(n27244) );
  NAND U35951 ( .A(n27247), .B(n27248), .Z(n27243) );
  AND U35952 ( .A(n27249), .B(n27250), .Z(n27137) );
  XOR U35953 ( .A(n27217), .B(n27216), .Z(N62971) );
  XNOR U35954 ( .A(n27234), .B(n27235), .Z(n27216) );
  XNOR U35955 ( .A(n27249), .B(n27250), .Z(n27235) );
  XOR U35956 ( .A(n27246), .B(n27245), .Z(n27250) );
  XOR U35957 ( .A(y[4404]), .B(x[4404]), .Z(n27245) );
  XOR U35958 ( .A(n27248), .B(n27247), .Z(n27246) );
  XOR U35959 ( .A(y[4406]), .B(x[4406]), .Z(n27247) );
  XOR U35960 ( .A(y[4405]), .B(x[4405]), .Z(n27248) );
  XOR U35961 ( .A(n27240), .B(n27239), .Z(n27249) );
  XOR U35962 ( .A(n27242), .B(n27241), .Z(n27239) );
  XOR U35963 ( .A(y[4403]), .B(x[4403]), .Z(n27241) );
  XOR U35964 ( .A(y[4402]), .B(x[4402]), .Z(n27242) );
  XOR U35965 ( .A(y[4401]), .B(x[4401]), .Z(n27240) );
  XNOR U35966 ( .A(n27233), .B(n27232), .Z(n27234) );
  XNOR U35967 ( .A(n27229), .B(n27228), .Z(n27232) );
  XOR U35968 ( .A(n27231), .B(n27230), .Z(n27228) );
  XOR U35969 ( .A(y[4400]), .B(x[4400]), .Z(n27230) );
  XOR U35970 ( .A(y[4399]), .B(x[4399]), .Z(n27231) );
  XOR U35971 ( .A(y[4398]), .B(x[4398]), .Z(n27229) );
  XOR U35972 ( .A(n27223), .B(n27222), .Z(n27233) );
  XOR U35973 ( .A(n27225), .B(n27224), .Z(n27222) );
  XOR U35974 ( .A(y[4397]), .B(x[4397]), .Z(n27224) );
  XOR U35975 ( .A(y[4396]), .B(x[4396]), .Z(n27225) );
  XOR U35976 ( .A(y[4395]), .B(x[4395]), .Z(n27223) );
  XNOR U35977 ( .A(n27199), .B(n27200), .Z(n27217) );
  XNOR U35978 ( .A(n27214), .B(n27215), .Z(n27200) );
  XOR U35979 ( .A(n27211), .B(n27210), .Z(n27215) );
  XOR U35980 ( .A(y[4392]), .B(x[4392]), .Z(n27210) );
  XOR U35981 ( .A(n27213), .B(n27212), .Z(n27211) );
  XOR U35982 ( .A(y[4394]), .B(x[4394]), .Z(n27212) );
  XOR U35983 ( .A(y[4393]), .B(x[4393]), .Z(n27213) );
  XOR U35984 ( .A(n27205), .B(n27204), .Z(n27214) );
  XOR U35985 ( .A(n27207), .B(n27206), .Z(n27204) );
  XOR U35986 ( .A(y[4391]), .B(x[4391]), .Z(n27206) );
  XOR U35987 ( .A(y[4390]), .B(x[4390]), .Z(n27207) );
  XOR U35988 ( .A(y[4389]), .B(x[4389]), .Z(n27205) );
  XNOR U35989 ( .A(n27198), .B(n27197), .Z(n27199) );
  XNOR U35990 ( .A(n27194), .B(n27193), .Z(n27197) );
  XOR U35991 ( .A(n27196), .B(n27195), .Z(n27193) );
  XOR U35992 ( .A(y[4388]), .B(x[4388]), .Z(n27195) );
  XOR U35993 ( .A(y[4387]), .B(x[4387]), .Z(n27196) );
  XOR U35994 ( .A(y[4386]), .B(x[4386]), .Z(n27194) );
  XOR U35995 ( .A(n27188), .B(n27187), .Z(n27198) );
  XOR U35996 ( .A(n27190), .B(n27189), .Z(n27187) );
  XOR U35997 ( .A(y[4385]), .B(x[4385]), .Z(n27189) );
  XOR U35998 ( .A(y[4384]), .B(x[4384]), .Z(n27190) );
  XOR U35999 ( .A(y[4383]), .B(x[4383]), .Z(n27188) );
  NAND U36000 ( .A(n27251), .B(n27252), .Z(N62962) );
  NAND U36001 ( .A(n27253), .B(n27254), .Z(n27252) );
  NANDN U36002 ( .A(n27255), .B(n27256), .Z(n27254) );
  NANDN U36003 ( .A(n27256), .B(n27255), .Z(n27251) );
  XOR U36004 ( .A(n27255), .B(n27257), .Z(N62961) );
  XNOR U36005 ( .A(n27253), .B(n27256), .Z(n27257) );
  NAND U36006 ( .A(n27258), .B(n27259), .Z(n27256) );
  NAND U36007 ( .A(n27260), .B(n27261), .Z(n27259) );
  NANDN U36008 ( .A(n27262), .B(n27263), .Z(n27261) );
  NANDN U36009 ( .A(n27263), .B(n27262), .Z(n27258) );
  AND U36010 ( .A(n27264), .B(n27265), .Z(n27253) );
  NAND U36011 ( .A(n27266), .B(n27267), .Z(n27265) );
  NANDN U36012 ( .A(n27268), .B(n27269), .Z(n27267) );
  NANDN U36013 ( .A(n27269), .B(n27268), .Z(n27264) );
  IV U36014 ( .A(n27270), .Z(n27269) );
  AND U36015 ( .A(n27271), .B(n27272), .Z(n27255) );
  NAND U36016 ( .A(n27273), .B(n27274), .Z(n27272) );
  NANDN U36017 ( .A(n27275), .B(n27276), .Z(n27274) );
  NANDN U36018 ( .A(n27276), .B(n27275), .Z(n27271) );
  XOR U36019 ( .A(n27268), .B(n27277), .Z(N62960) );
  XNOR U36020 ( .A(n27266), .B(n27270), .Z(n27277) );
  XOR U36021 ( .A(n27263), .B(n27278), .Z(n27270) );
  XNOR U36022 ( .A(n27260), .B(n27262), .Z(n27278) );
  AND U36023 ( .A(n27279), .B(n27280), .Z(n27262) );
  NANDN U36024 ( .A(n27281), .B(n27282), .Z(n27280) );
  OR U36025 ( .A(n27283), .B(n27284), .Z(n27282) );
  IV U36026 ( .A(n27285), .Z(n27284) );
  NANDN U36027 ( .A(n27285), .B(n27283), .Z(n27279) );
  AND U36028 ( .A(n27286), .B(n27287), .Z(n27260) );
  NAND U36029 ( .A(n27288), .B(n27289), .Z(n27287) );
  NANDN U36030 ( .A(n27290), .B(n27291), .Z(n27289) );
  NANDN U36031 ( .A(n27291), .B(n27290), .Z(n27286) );
  IV U36032 ( .A(n27292), .Z(n27291) );
  NAND U36033 ( .A(n27293), .B(n27294), .Z(n27263) );
  NANDN U36034 ( .A(n27295), .B(n27296), .Z(n27294) );
  NANDN U36035 ( .A(n27297), .B(n27298), .Z(n27296) );
  NANDN U36036 ( .A(n27298), .B(n27297), .Z(n27293) );
  IV U36037 ( .A(n27299), .Z(n27297) );
  AND U36038 ( .A(n27300), .B(n27301), .Z(n27266) );
  NAND U36039 ( .A(n27302), .B(n27303), .Z(n27301) );
  NANDN U36040 ( .A(n27304), .B(n27305), .Z(n27303) );
  NANDN U36041 ( .A(n27305), .B(n27304), .Z(n27300) );
  XOR U36042 ( .A(n27276), .B(n27306), .Z(n27268) );
  XNOR U36043 ( .A(n27273), .B(n27275), .Z(n27306) );
  AND U36044 ( .A(n27307), .B(n27308), .Z(n27275) );
  NANDN U36045 ( .A(n27309), .B(n27310), .Z(n27308) );
  OR U36046 ( .A(n27311), .B(n27312), .Z(n27310) );
  IV U36047 ( .A(n27313), .Z(n27312) );
  NANDN U36048 ( .A(n27313), .B(n27311), .Z(n27307) );
  AND U36049 ( .A(n27314), .B(n27315), .Z(n27273) );
  NAND U36050 ( .A(n27316), .B(n27317), .Z(n27315) );
  NANDN U36051 ( .A(n27318), .B(n27319), .Z(n27317) );
  NANDN U36052 ( .A(n27319), .B(n27318), .Z(n27314) );
  IV U36053 ( .A(n27320), .Z(n27319) );
  NAND U36054 ( .A(n27321), .B(n27322), .Z(n27276) );
  NANDN U36055 ( .A(n27323), .B(n27324), .Z(n27322) );
  NANDN U36056 ( .A(n27325), .B(n27326), .Z(n27324) );
  NANDN U36057 ( .A(n27326), .B(n27325), .Z(n27321) );
  IV U36058 ( .A(n27327), .Z(n27325) );
  XOR U36059 ( .A(n27302), .B(n27328), .Z(N62959) );
  XNOR U36060 ( .A(n27305), .B(n27304), .Z(n27328) );
  XNOR U36061 ( .A(n27316), .B(n27329), .Z(n27304) );
  XNOR U36062 ( .A(n27320), .B(n27318), .Z(n27329) );
  XOR U36063 ( .A(n27326), .B(n27330), .Z(n27318) );
  XNOR U36064 ( .A(n27323), .B(n27327), .Z(n27330) );
  AND U36065 ( .A(n27331), .B(n27332), .Z(n27327) );
  NAND U36066 ( .A(n27333), .B(n27334), .Z(n27332) );
  NAND U36067 ( .A(n27335), .B(n27336), .Z(n27331) );
  AND U36068 ( .A(n27337), .B(n27338), .Z(n27323) );
  NAND U36069 ( .A(n27339), .B(n27340), .Z(n27338) );
  NAND U36070 ( .A(n27341), .B(n27342), .Z(n27337) );
  NANDN U36071 ( .A(n27343), .B(n27344), .Z(n27326) );
  ANDN U36072 ( .B(n27345), .A(n27346), .Z(n27320) );
  XNOR U36073 ( .A(n27311), .B(n27347), .Z(n27316) );
  XNOR U36074 ( .A(n27309), .B(n27313), .Z(n27347) );
  AND U36075 ( .A(n27348), .B(n27349), .Z(n27313) );
  NAND U36076 ( .A(n27350), .B(n27351), .Z(n27349) );
  NAND U36077 ( .A(n27352), .B(n27353), .Z(n27348) );
  AND U36078 ( .A(n27354), .B(n27355), .Z(n27309) );
  NAND U36079 ( .A(n27356), .B(n27357), .Z(n27355) );
  NAND U36080 ( .A(n27358), .B(n27359), .Z(n27354) );
  AND U36081 ( .A(n27360), .B(n27361), .Z(n27311) );
  NAND U36082 ( .A(n27362), .B(n27363), .Z(n27305) );
  XNOR U36083 ( .A(n27288), .B(n27364), .Z(n27302) );
  XNOR U36084 ( .A(n27292), .B(n27290), .Z(n27364) );
  XOR U36085 ( .A(n27298), .B(n27365), .Z(n27290) );
  XNOR U36086 ( .A(n27295), .B(n27299), .Z(n27365) );
  AND U36087 ( .A(n27366), .B(n27367), .Z(n27299) );
  NAND U36088 ( .A(n27368), .B(n27369), .Z(n27367) );
  NAND U36089 ( .A(n27370), .B(n27371), .Z(n27366) );
  AND U36090 ( .A(n27372), .B(n27373), .Z(n27295) );
  NAND U36091 ( .A(n27374), .B(n27375), .Z(n27373) );
  NAND U36092 ( .A(n27376), .B(n27377), .Z(n27372) );
  NANDN U36093 ( .A(n27378), .B(n27379), .Z(n27298) );
  ANDN U36094 ( .B(n27380), .A(n27381), .Z(n27292) );
  XNOR U36095 ( .A(n27283), .B(n27382), .Z(n27288) );
  XNOR U36096 ( .A(n27281), .B(n27285), .Z(n27382) );
  AND U36097 ( .A(n27383), .B(n27384), .Z(n27285) );
  NAND U36098 ( .A(n27385), .B(n27386), .Z(n27384) );
  NAND U36099 ( .A(n27387), .B(n27388), .Z(n27383) );
  AND U36100 ( .A(n27389), .B(n27390), .Z(n27281) );
  NAND U36101 ( .A(n27391), .B(n27392), .Z(n27390) );
  NAND U36102 ( .A(n27393), .B(n27394), .Z(n27389) );
  AND U36103 ( .A(n27395), .B(n27396), .Z(n27283) );
  XOR U36104 ( .A(n27363), .B(n27362), .Z(N62958) );
  XNOR U36105 ( .A(n27380), .B(n27381), .Z(n27362) );
  XNOR U36106 ( .A(n27395), .B(n27396), .Z(n27381) );
  XOR U36107 ( .A(n27392), .B(n27391), .Z(n27396) );
  XOR U36108 ( .A(y[4380]), .B(x[4380]), .Z(n27391) );
  XOR U36109 ( .A(n27394), .B(n27393), .Z(n27392) );
  XOR U36110 ( .A(y[4382]), .B(x[4382]), .Z(n27393) );
  XOR U36111 ( .A(y[4381]), .B(x[4381]), .Z(n27394) );
  XOR U36112 ( .A(n27386), .B(n27385), .Z(n27395) );
  XOR U36113 ( .A(n27388), .B(n27387), .Z(n27385) );
  XOR U36114 ( .A(y[4379]), .B(x[4379]), .Z(n27387) );
  XOR U36115 ( .A(y[4378]), .B(x[4378]), .Z(n27388) );
  XOR U36116 ( .A(y[4377]), .B(x[4377]), .Z(n27386) );
  XNOR U36117 ( .A(n27379), .B(n27378), .Z(n27380) );
  XNOR U36118 ( .A(n27375), .B(n27374), .Z(n27378) );
  XOR U36119 ( .A(n27377), .B(n27376), .Z(n27374) );
  XOR U36120 ( .A(y[4376]), .B(x[4376]), .Z(n27376) );
  XOR U36121 ( .A(y[4375]), .B(x[4375]), .Z(n27377) );
  XOR U36122 ( .A(y[4374]), .B(x[4374]), .Z(n27375) );
  XOR U36123 ( .A(n27369), .B(n27368), .Z(n27379) );
  XOR U36124 ( .A(n27371), .B(n27370), .Z(n27368) );
  XOR U36125 ( .A(y[4373]), .B(x[4373]), .Z(n27370) );
  XOR U36126 ( .A(y[4372]), .B(x[4372]), .Z(n27371) );
  XOR U36127 ( .A(y[4371]), .B(x[4371]), .Z(n27369) );
  XNOR U36128 ( .A(n27345), .B(n27346), .Z(n27363) );
  XNOR U36129 ( .A(n27360), .B(n27361), .Z(n27346) );
  XOR U36130 ( .A(n27357), .B(n27356), .Z(n27361) );
  XOR U36131 ( .A(y[4368]), .B(x[4368]), .Z(n27356) );
  XOR U36132 ( .A(n27359), .B(n27358), .Z(n27357) );
  XOR U36133 ( .A(y[4370]), .B(x[4370]), .Z(n27358) );
  XOR U36134 ( .A(y[4369]), .B(x[4369]), .Z(n27359) );
  XOR U36135 ( .A(n27351), .B(n27350), .Z(n27360) );
  XOR U36136 ( .A(n27353), .B(n27352), .Z(n27350) );
  XOR U36137 ( .A(y[4367]), .B(x[4367]), .Z(n27352) );
  XOR U36138 ( .A(y[4366]), .B(x[4366]), .Z(n27353) );
  XOR U36139 ( .A(y[4365]), .B(x[4365]), .Z(n27351) );
  XNOR U36140 ( .A(n27344), .B(n27343), .Z(n27345) );
  XNOR U36141 ( .A(n27340), .B(n27339), .Z(n27343) );
  XOR U36142 ( .A(n27342), .B(n27341), .Z(n27339) );
  XOR U36143 ( .A(y[4364]), .B(x[4364]), .Z(n27341) );
  XOR U36144 ( .A(y[4363]), .B(x[4363]), .Z(n27342) );
  XOR U36145 ( .A(y[4362]), .B(x[4362]), .Z(n27340) );
  XOR U36146 ( .A(n27334), .B(n27333), .Z(n27344) );
  XOR U36147 ( .A(n27336), .B(n27335), .Z(n27333) );
  XOR U36148 ( .A(y[4361]), .B(x[4361]), .Z(n27335) );
  XOR U36149 ( .A(y[4360]), .B(x[4360]), .Z(n27336) );
  XOR U36150 ( .A(y[4359]), .B(x[4359]), .Z(n27334) );
  NAND U36151 ( .A(n27397), .B(n27398), .Z(N62949) );
  NAND U36152 ( .A(n27399), .B(n27400), .Z(n27398) );
  NANDN U36153 ( .A(n27401), .B(n27402), .Z(n27400) );
  NANDN U36154 ( .A(n27402), .B(n27401), .Z(n27397) );
  XOR U36155 ( .A(n27401), .B(n27403), .Z(N62948) );
  XNOR U36156 ( .A(n27399), .B(n27402), .Z(n27403) );
  NAND U36157 ( .A(n27404), .B(n27405), .Z(n27402) );
  NAND U36158 ( .A(n27406), .B(n27407), .Z(n27405) );
  NANDN U36159 ( .A(n27408), .B(n27409), .Z(n27407) );
  NANDN U36160 ( .A(n27409), .B(n27408), .Z(n27404) );
  AND U36161 ( .A(n27410), .B(n27411), .Z(n27399) );
  NAND U36162 ( .A(n27412), .B(n27413), .Z(n27411) );
  NANDN U36163 ( .A(n27414), .B(n27415), .Z(n27413) );
  NANDN U36164 ( .A(n27415), .B(n27414), .Z(n27410) );
  IV U36165 ( .A(n27416), .Z(n27415) );
  AND U36166 ( .A(n27417), .B(n27418), .Z(n27401) );
  NAND U36167 ( .A(n27419), .B(n27420), .Z(n27418) );
  NANDN U36168 ( .A(n27421), .B(n27422), .Z(n27420) );
  NANDN U36169 ( .A(n27422), .B(n27421), .Z(n27417) );
  XOR U36170 ( .A(n27414), .B(n27423), .Z(N62947) );
  XNOR U36171 ( .A(n27412), .B(n27416), .Z(n27423) );
  XOR U36172 ( .A(n27409), .B(n27424), .Z(n27416) );
  XNOR U36173 ( .A(n27406), .B(n27408), .Z(n27424) );
  AND U36174 ( .A(n27425), .B(n27426), .Z(n27408) );
  NANDN U36175 ( .A(n27427), .B(n27428), .Z(n27426) );
  OR U36176 ( .A(n27429), .B(n27430), .Z(n27428) );
  IV U36177 ( .A(n27431), .Z(n27430) );
  NANDN U36178 ( .A(n27431), .B(n27429), .Z(n27425) );
  AND U36179 ( .A(n27432), .B(n27433), .Z(n27406) );
  NAND U36180 ( .A(n27434), .B(n27435), .Z(n27433) );
  NANDN U36181 ( .A(n27436), .B(n27437), .Z(n27435) );
  NANDN U36182 ( .A(n27437), .B(n27436), .Z(n27432) );
  IV U36183 ( .A(n27438), .Z(n27437) );
  NAND U36184 ( .A(n27439), .B(n27440), .Z(n27409) );
  NANDN U36185 ( .A(n27441), .B(n27442), .Z(n27440) );
  NANDN U36186 ( .A(n27443), .B(n27444), .Z(n27442) );
  NANDN U36187 ( .A(n27444), .B(n27443), .Z(n27439) );
  IV U36188 ( .A(n27445), .Z(n27443) );
  AND U36189 ( .A(n27446), .B(n27447), .Z(n27412) );
  NAND U36190 ( .A(n27448), .B(n27449), .Z(n27447) );
  NANDN U36191 ( .A(n27450), .B(n27451), .Z(n27449) );
  NANDN U36192 ( .A(n27451), .B(n27450), .Z(n27446) );
  XOR U36193 ( .A(n27422), .B(n27452), .Z(n27414) );
  XNOR U36194 ( .A(n27419), .B(n27421), .Z(n27452) );
  AND U36195 ( .A(n27453), .B(n27454), .Z(n27421) );
  NANDN U36196 ( .A(n27455), .B(n27456), .Z(n27454) );
  OR U36197 ( .A(n27457), .B(n27458), .Z(n27456) );
  IV U36198 ( .A(n27459), .Z(n27458) );
  NANDN U36199 ( .A(n27459), .B(n27457), .Z(n27453) );
  AND U36200 ( .A(n27460), .B(n27461), .Z(n27419) );
  NAND U36201 ( .A(n27462), .B(n27463), .Z(n27461) );
  NANDN U36202 ( .A(n27464), .B(n27465), .Z(n27463) );
  NANDN U36203 ( .A(n27465), .B(n27464), .Z(n27460) );
  IV U36204 ( .A(n27466), .Z(n27465) );
  NAND U36205 ( .A(n27467), .B(n27468), .Z(n27422) );
  NANDN U36206 ( .A(n27469), .B(n27470), .Z(n27468) );
  NANDN U36207 ( .A(n27471), .B(n27472), .Z(n27470) );
  NANDN U36208 ( .A(n27472), .B(n27471), .Z(n27467) );
  IV U36209 ( .A(n27473), .Z(n27471) );
  XOR U36210 ( .A(n27448), .B(n27474), .Z(N62946) );
  XNOR U36211 ( .A(n27451), .B(n27450), .Z(n27474) );
  XNOR U36212 ( .A(n27462), .B(n27475), .Z(n27450) );
  XNOR U36213 ( .A(n27466), .B(n27464), .Z(n27475) );
  XOR U36214 ( .A(n27472), .B(n27476), .Z(n27464) );
  XNOR U36215 ( .A(n27469), .B(n27473), .Z(n27476) );
  AND U36216 ( .A(n27477), .B(n27478), .Z(n27473) );
  NAND U36217 ( .A(n27479), .B(n27480), .Z(n27478) );
  NAND U36218 ( .A(n27481), .B(n27482), .Z(n27477) );
  AND U36219 ( .A(n27483), .B(n27484), .Z(n27469) );
  NAND U36220 ( .A(n27485), .B(n27486), .Z(n27484) );
  NAND U36221 ( .A(n27487), .B(n27488), .Z(n27483) );
  NANDN U36222 ( .A(n27489), .B(n27490), .Z(n27472) );
  ANDN U36223 ( .B(n27491), .A(n27492), .Z(n27466) );
  XNOR U36224 ( .A(n27457), .B(n27493), .Z(n27462) );
  XNOR U36225 ( .A(n27455), .B(n27459), .Z(n27493) );
  AND U36226 ( .A(n27494), .B(n27495), .Z(n27459) );
  NAND U36227 ( .A(n27496), .B(n27497), .Z(n27495) );
  NAND U36228 ( .A(n27498), .B(n27499), .Z(n27494) );
  AND U36229 ( .A(n27500), .B(n27501), .Z(n27455) );
  NAND U36230 ( .A(n27502), .B(n27503), .Z(n27501) );
  NAND U36231 ( .A(n27504), .B(n27505), .Z(n27500) );
  AND U36232 ( .A(n27506), .B(n27507), .Z(n27457) );
  NAND U36233 ( .A(n27508), .B(n27509), .Z(n27451) );
  XNOR U36234 ( .A(n27434), .B(n27510), .Z(n27448) );
  XNOR U36235 ( .A(n27438), .B(n27436), .Z(n27510) );
  XOR U36236 ( .A(n27444), .B(n27511), .Z(n27436) );
  XNOR U36237 ( .A(n27441), .B(n27445), .Z(n27511) );
  AND U36238 ( .A(n27512), .B(n27513), .Z(n27445) );
  NAND U36239 ( .A(n27514), .B(n27515), .Z(n27513) );
  NAND U36240 ( .A(n27516), .B(n27517), .Z(n27512) );
  AND U36241 ( .A(n27518), .B(n27519), .Z(n27441) );
  NAND U36242 ( .A(n27520), .B(n27521), .Z(n27519) );
  NAND U36243 ( .A(n27522), .B(n27523), .Z(n27518) );
  NANDN U36244 ( .A(n27524), .B(n27525), .Z(n27444) );
  ANDN U36245 ( .B(n27526), .A(n27527), .Z(n27438) );
  XNOR U36246 ( .A(n27429), .B(n27528), .Z(n27434) );
  XNOR U36247 ( .A(n27427), .B(n27431), .Z(n27528) );
  AND U36248 ( .A(n27529), .B(n27530), .Z(n27431) );
  NAND U36249 ( .A(n27531), .B(n27532), .Z(n27530) );
  NAND U36250 ( .A(n27533), .B(n27534), .Z(n27529) );
  AND U36251 ( .A(n27535), .B(n27536), .Z(n27427) );
  NAND U36252 ( .A(n27537), .B(n27538), .Z(n27536) );
  NAND U36253 ( .A(n27539), .B(n27540), .Z(n27535) );
  AND U36254 ( .A(n27541), .B(n27542), .Z(n27429) );
  XOR U36255 ( .A(n27509), .B(n27508), .Z(N62945) );
  XNOR U36256 ( .A(n27526), .B(n27527), .Z(n27508) );
  XNOR U36257 ( .A(n27541), .B(n27542), .Z(n27527) );
  XOR U36258 ( .A(n27538), .B(n27537), .Z(n27542) );
  XOR U36259 ( .A(y[4356]), .B(x[4356]), .Z(n27537) );
  XOR U36260 ( .A(n27540), .B(n27539), .Z(n27538) );
  XOR U36261 ( .A(y[4358]), .B(x[4358]), .Z(n27539) );
  XOR U36262 ( .A(y[4357]), .B(x[4357]), .Z(n27540) );
  XOR U36263 ( .A(n27532), .B(n27531), .Z(n27541) );
  XOR U36264 ( .A(n27534), .B(n27533), .Z(n27531) );
  XOR U36265 ( .A(y[4355]), .B(x[4355]), .Z(n27533) );
  XOR U36266 ( .A(y[4354]), .B(x[4354]), .Z(n27534) );
  XOR U36267 ( .A(y[4353]), .B(x[4353]), .Z(n27532) );
  XNOR U36268 ( .A(n27525), .B(n27524), .Z(n27526) );
  XNOR U36269 ( .A(n27521), .B(n27520), .Z(n27524) );
  XOR U36270 ( .A(n27523), .B(n27522), .Z(n27520) );
  XOR U36271 ( .A(y[4352]), .B(x[4352]), .Z(n27522) );
  XOR U36272 ( .A(y[4351]), .B(x[4351]), .Z(n27523) );
  XOR U36273 ( .A(y[4350]), .B(x[4350]), .Z(n27521) );
  XOR U36274 ( .A(n27515), .B(n27514), .Z(n27525) );
  XOR U36275 ( .A(n27517), .B(n27516), .Z(n27514) );
  XOR U36276 ( .A(y[4349]), .B(x[4349]), .Z(n27516) );
  XOR U36277 ( .A(y[4348]), .B(x[4348]), .Z(n27517) );
  XOR U36278 ( .A(y[4347]), .B(x[4347]), .Z(n27515) );
  XNOR U36279 ( .A(n27491), .B(n27492), .Z(n27509) );
  XNOR U36280 ( .A(n27506), .B(n27507), .Z(n27492) );
  XOR U36281 ( .A(n27503), .B(n27502), .Z(n27507) );
  XOR U36282 ( .A(y[4344]), .B(x[4344]), .Z(n27502) );
  XOR U36283 ( .A(n27505), .B(n27504), .Z(n27503) );
  XOR U36284 ( .A(y[4346]), .B(x[4346]), .Z(n27504) );
  XOR U36285 ( .A(y[4345]), .B(x[4345]), .Z(n27505) );
  XOR U36286 ( .A(n27497), .B(n27496), .Z(n27506) );
  XOR U36287 ( .A(n27499), .B(n27498), .Z(n27496) );
  XOR U36288 ( .A(y[4343]), .B(x[4343]), .Z(n27498) );
  XOR U36289 ( .A(y[4342]), .B(x[4342]), .Z(n27499) );
  XOR U36290 ( .A(y[4341]), .B(x[4341]), .Z(n27497) );
  XNOR U36291 ( .A(n27490), .B(n27489), .Z(n27491) );
  XNOR U36292 ( .A(n27486), .B(n27485), .Z(n27489) );
  XOR U36293 ( .A(n27488), .B(n27487), .Z(n27485) );
  XOR U36294 ( .A(y[4340]), .B(x[4340]), .Z(n27487) );
  XOR U36295 ( .A(y[4339]), .B(x[4339]), .Z(n27488) );
  XOR U36296 ( .A(y[4338]), .B(x[4338]), .Z(n27486) );
  XOR U36297 ( .A(n27480), .B(n27479), .Z(n27490) );
  XOR U36298 ( .A(n27482), .B(n27481), .Z(n27479) );
  XOR U36299 ( .A(y[4337]), .B(x[4337]), .Z(n27481) );
  XOR U36300 ( .A(y[4336]), .B(x[4336]), .Z(n27482) );
  XOR U36301 ( .A(y[4335]), .B(x[4335]), .Z(n27480) );
  NAND U36302 ( .A(n27543), .B(n27544), .Z(N62936) );
  NAND U36303 ( .A(n27545), .B(n27546), .Z(n27544) );
  NANDN U36304 ( .A(n27547), .B(n27548), .Z(n27546) );
  NANDN U36305 ( .A(n27548), .B(n27547), .Z(n27543) );
  XOR U36306 ( .A(n27547), .B(n27549), .Z(N62935) );
  XNOR U36307 ( .A(n27545), .B(n27548), .Z(n27549) );
  NAND U36308 ( .A(n27550), .B(n27551), .Z(n27548) );
  NAND U36309 ( .A(n27552), .B(n27553), .Z(n27551) );
  NANDN U36310 ( .A(n27554), .B(n27555), .Z(n27553) );
  NANDN U36311 ( .A(n27555), .B(n27554), .Z(n27550) );
  AND U36312 ( .A(n27556), .B(n27557), .Z(n27545) );
  NAND U36313 ( .A(n27558), .B(n27559), .Z(n27557) );
  NANDN U36314 ( .A(n27560), .B(n27561), .Z(n27559) );
  NANDN U36315 ( .A(n27561), .B(n27560), .Z(n27556) );
  IV U36316 ( .A(n27562), .Z(n27561) );
  AND U36317 ( .A(n27563), .B(n27564), .Z(n27547) );
  NAND U36318 ( .A(n27565), .B(n27566), .Z(n27564) );
  NANDN U36319 ( .A(n27567), .B(n27568), .Z(n27566) );
  NANDN U36320 ( .A(n27568), .B(n27567), .Z(n27563) );
  XOR U36321 ( .A(n27560), .B(n27569), .Z(N62934) );
  XNOR U36322 ( .A(n27558), .B(n27562), .Z(n27569) );
  XOR U36323 ( .A(n27555), .B(n27570), .Z(n27562) );
  XNOR U36324 ( .A(n27552), .B(n27554), .Z(n27570) );
  AND U36325 ( .A(n27571), .B(n27572), .Z(n27554) );
  NANDN U36326 ( .A(n27573), .B(n27574), .Z(n27572) );
  OR U36327 ( .A(n27575), .B(n27576), .Z(n27574) );
  IV U36328 ( .A(n27577), .Z(n27576) );
  NANDN U36329 ( .A(n27577), .B(n27575), .Z(n27571) );
  AND U36330 ( .A(n27578), .B(n27579), .Z(n27552) );
  NAND U36331 ( .A(n27580), .B(n27581), .Z(n27579) );
  NANDN U36332 ( .A(n27582), .B(n27583), .Z(n27581) );
  NANDN U36333 ( .A(n27583), .B(n27582), .Z(n27578) );
  IV U36334 ( .A(n27584), .Z(n27583) );
  NAND U36335 ( .A(n27585), .B(n27586), .Z(n27555) );
  NANDN U36336 ( .A(n27587), .B(n27588), .Z(n27586) );
  NANDN U36337 ( .A(n27589), .B(n27590), .Z(n27588) );
  NANDN U36338 ( .A(n27590), .B(n27589), .Z(n27585) );
  IV U36339 ( .A(n27591), .Z(n27589) );
  AND U36340 ( .A(n27592), .B(n27593), .Z(n27558) );
  NAND U36341 ( .A(n27594), .B(n27595), .Z(n27593) );
  NANDN U36342 ( .A(n27596), .B(n27597), .Z(n27595) );
  NANDN U36343 ( .A(n27597), .B(n27596), .Z(n27592) );
  XOR U36344 ( .A(n27568), .B(n27598), .Z(n27560) );
  XNOR U36345 ( .A(n27565), .B(n27567), .Z(n27598) );
  AND U36346 ( .A(n27599), .B(n27600), .Z(n27567) );
  NANDN U36347 ( .A(n27601), .B(n27602), .Z(n27600) );
  OR U36348 ( .A(n27603), .B(n27604), .Z(n27602) );
  IV U36349 ( .A(n27605), .Z(n27604) );
  NANDN U36350 ( .A(n27605), .B(n27603), .Z(n27599) );
  AND U36351 ( .A(n27606), .B(n27607), .Z(n27565) );
  NAND U36352 ( .A(n27608), .B(n27609), .Z(n27607) );
  NANDN U36353 ( .A(n27610), .B(n27611), .Z(n27609) );
  NANDN U36354 ( .A(n27611), .B(n27610), .Z(n27606) );
  IV U36355 ( .A(n27612), .Z(n27611) );
  NAND U36356 ( .A(n27613), .B(n27614), .Z(n27568) );
  NANDN U36357 ( .A(n27615), .B(n27616), .Z(n27614) );
  NANDN U36358 ( .A(n27617), .B(n27618), .Z(n27616) );
  NANDN U36359 ( .A(n27618), .B(n27617), .Z(n27613) );
  IV U36360 ( .A(n27619), .Z(n27617) );
  XOR U36361 ( .A(n27594), .B(n27620), .Z(N62933) );
  XNOR U36362 ( .A(n27597), .B(n27596), .Z(n27620) );
  XNOR U36363 ( .A(n27608), .B(n27621), .Z(n27596) );
  XNOR U36364 ( .A(n27612), .B(n27610), .Z(n27621) );
  XOR U36365 ( .A(n27618), .B(n27622), .Z(n27610) );
  XNOR U36366 ( .A(n27615), .B(n27619), .Z(n27622) );
  AND U36367 ( .A(n27623), .B(n27624), .Z(n27619) );
  NAND U36368 ( .A(n27625), .B(n27626), .Z(n27624) );
  NAND U36369 ( .A(n27627), .B(n27628), .Z(n27623) );
  AND U36370 ( .A(n27629), .B(n27630), .Z(n27615) );
  NAND U36371 ( .A(n27631), .B(n27632), .Z(n27630) );
  NAND U36372 ( .A(n27633), .B(n27634), .Z(n27629) );
  NANDN U36373 ( .A(n27635), .B(n27636), .Z(n27618) );
  ANDN U36374 ( .B(n27637), .A(n27638), .Z(n27612) );
  XNOR U36375 ( .A(n27603), .B(n27639), .Z(n27608) );
  XNOR U36376 ( .A(n27601), .B(n27605), .Z(n27639) );
  AND U36377 ( .A(n27640), .B(n27641), .Z(n27605) );
  NAND U36378 ( .A(n27642), .B(n27643), .Z(n27641) );
  NAND U36379 ( .A(n27644), .B(n27645), .Z(n27640) );
  AND U36380 ( .A(n27646), .B(n27647), .Z(n27601) );
  NAND U36381 ( .A(n27648), .B(n27649), .Z(n27647) );
  NAND U36382 ( .A(n27650), .B(n27651), .Z(n27646) );
  AND U36383 ( .A(n27652), .B(n27653), .Z(n27603) );
  NAND U36384 ( .A(n27654), .B(n27655), .Z(n27597) );
  XNOR U36385 ( .A(n27580), .B(n27656), .Z(n27594) );
  XNOR U36386 ( .A(n27584), .B(n27582), .Z(n27656) );
  XOR U36387 ( .A(n27590), .B(n27657), .Z(n27582) );
  XNOR U36388 ( .A(n27587), .B(n27591), .Z(n27657) );
  AND U36389 ( .A(n27658), .B(n27659), .Z(n27591) );
  NAND U36390 ( .A(n27660), .B(n27661), .Z(n27659) );
  NAND U36391 ( .A(n27662), .B(n27663), .Z(n27658) );
  AND U36392 ( .A(n27664), .B(n27665), .Z(n27587) );
  NAND U36393 ( .A(n27666), .B(n27667), .Z(n27665) );
  NAND U36394 ( .A(n27668), .B(n27669), .Z(n27664) );
  NANDN U36395 ( .A(n27670), .B(n27671), .Z(n27590) );
  ANDN U36396 ( .B(n27672), .A(n27673), .Z(n27584) );
  XNOR U36397 ( .A(n27575), .B(n27674), .Z(n27580) );
  XNOR U36398 ( .A(n27573), .B(n27577), .Z(n27674) );
  AND U36399 ( .A(n27675), .B(n27676), .Z(n27577) );
  NAND U36400 ( .A(n27677), .B(n27678), .Z(n27676) );
  NAND U36401 ( .A(n27679), .B(n27680), .Z(n27675) );
  AND U36402 ( .A(n27681), .B(n27682), .Z(n27573) );
  NAND U36403 ( .A(n27683), .B(n27684), .Z(n27682) );
  NAND U36404 ( .A(n27685), .B(n27686), .Z(n27681) );
  AND U36405 ( .A(n27687), .B(n27688), .Z(n27575) );
  XOR U36406 ( .A(n27655), .B(n27654), .Z(N62932) );
  XNOR U36407 ( .A(n27672), .B(n27673), .Z(n27654) );
  XNOR U36408 ( .A(n27687), .B(n27688), .Z(n27673) );
  XOR U36409 ( .A(n27684), .B(n27683), .Z(n27688) );
  XOR U36410 ( .A(y[4332]), .B(x[4332]), .Z(n27683) );
  XOR U36411 ( .A(n27686), .B(n27685), .Z(n27684) );
  XOR U36412 ( .A(y[4334]), .B(x[4334]), .Z(n27685) );
  XOR U36413 ( .A(y[4333]), .B(x[4333]), .Z(n27686) );
  XOR U36414 ( .A(n27678), .B(n27677), .Z(n27687) );
  XOR U36415 ( .A(n27680), .B(n27679), .Z(n27677) );
  XOR U36416 ( .A(y[4331]), .B(x[4331]), .Z(n27679) );
  XOR U36417 ( .A(y[4330]), .B(x[4330]), .Z(n27680) );
  XOR U36418 ( .A(y[4329]), .B(x[4329]), .Z(n27678) );
  XNOR U36419 ( .A(n27671), .B(n27670), .Z(n27672) );
  XNOR U36420 ( .A(n27667), .B(n27666), .Z(n27670) );
  XOR U36421 ( .A(n27669), .B(n27668), .Z(n27666) );
  XOR U36422 ( .A(y[4328]), .B(x[4328]), .Z(n27668) );
  XOR U36423 ( .A(y[4327]), .B(x[4327]), .Z(n27669) );
  XOR U36424 ( .A(y[4326]), .B(x[4326]), .Z(n27667) );
  XOR U36425 ( .A(n27661), .B(n27660), .Z(n27671) );
  XOR U36426 ( .A(n27663), .B(n27662), .Z(n27660) );
  XOR U36427 ( .A(y[4325]), .B(x[4325]), .Z(n27662) );
  XOR U36428 ( .A(y[4324]), .B(x[4324]), .Z(n27663) );
  XOR U36429 ( .A(y[4323]), .B(x[4323]), .Z(n27661) );
  XNOR U36430 ( .A(n27637), .B(n27638), .Z(n27655) );
  XNOR U36431 ( .A(n27652), .B(n27653), .Z(n27638) );
  XOR U36432 ( .A(n27649), .B(n27648), .Z(n27653) );
  XOR U36433 ( .A(y[4320]), .B(x[4320]), .Z(n27648) );
  XOR U36434 ( .A(n27651), .B(n27650), .Z(n27649) );
  XOR U36435 ( .A(y[4322]), .B(x[4322]), .Z(n27650) );
  XOR U36436 ( .A(y[4321]), .B(x[4321]), .Z(n27651) );
  XOR U36437 ( .A(n27643), .B(n27642), .Z(n27652) );
  XOR U36438 ( .A(n27645), .B(n27644), .Z(n27642) );
  XOR U36439 ( .A(y[4319]), .B(x[4319]), .Z(n27644) );
  XOR U36440 ( .A(y[4318]), .B(x[4318]), .Z(n27645) );
  XOR U36441 ( .A(y[4317]), .B(x[4317]), .Z(n27643) );
  XNOR U36442 ( .A(n27636), .B(n27635), .Z(n27637) );
  XNOR U36443 ( .A(n27632), .B(n27631), .Z(n27635) );
  XOR U36444 ( .A(n27634), .B(n27633), .Z(n27631) );
  XOR U36445 ( .A(y[4316]), .B(x[4316]), .Z(n27633) );
  XOR U36446 ( .A(y[4315]), .B(x[4315]), .Z(n27634) );
  XOR U36447 ( .A(y[4314]), .B(x[4314]), .Z(n27632) );
  XOR U36448 ( .A(n27626), .B(n27625), .Z(n27636) );
  XOR U36449 ( .A(n27628), .B(n27627), .Z(n27625) );
  XOR U36450 ( .A(y[4313]), .B(x[4313]), .Z(n27627) );
  XOR U36451 ( .A(y[4312]), .B(x[4312]), .Z(n27628) );
  XOR U36452 ( .A(y[4311]), .B(x[4311]), .Z(n27626) );
  NAND U36453 ( .A(n27689), .B(n27690), .Z(N62923) );
  NAND U36454 ( .A(n27691), .B(n27692), .Z(n27690) );
  NANDN U36455 ( .A(n27693), .B(n27694), .Z(n27692) );
  NANDN U36456 ( .A(n27694), .B(n27693), .Z(n27689) );
  XOR U36457 ( .A(n27693), .B(n27695), .Z(N62922) );
  XNOR U36458 ( .A(n27691), .B(n27694), .Z(n27695) );
  NAND U36459 ( .A(n27696), .B(n27697), .Z(n27694) );
  NAND U36460 ( .A(n27698), .B(n27699), .Z(n27697) );
  NANDN U36461 ( .A(n27700), .B(n27701), .Z(n27699) );
  NANDN U36462 ( .A(n27701), .B(n27700), .Z(n27696) );
  AND U36463 ( .A(n27702), .B(n27703), .Z(n27691) );
  NAND U36464 ( .A(n27704), .B(n27705), .Z(n27703) );
  NANDN U36465 ( .A(n27706), .B(n27707), .Z(n27705) );
  NANDN U36466 ( .A(n27707), .B(n27706), .Z(n27702) );
  IV U36467 ( .A(n27708), .Z(n27707) );
  AND U36468 ( .A(n27709), .B(n27710), .Z(n27693) );
  NAND U36469 ( .A(n27711), .B(n27712), .Z(n27710) );
  NANDN U36470 ( .A(n27713), .B(n27714), .Z(n27712) );
  NANDN U36471 ( .A(n27714), .B(n27713), .Z(n27709) );
  XOR U36472 ( .A(n27706), .B(n27715), .Z(N62921) );
  XNOR U36473 ( .A(n27704), .B(n27708), .Z(n27715) );
  XOR U36474 ( .A(n27701), .B(n27716), .Z(n27708) );
  XNOR U36475 ( .A(n27698), .B(n27700), .Z(n27716) );
  AND U36476 ( .A(n27717), .B(n27718), .Z(n27700) );
  NANDN U36477 ( .A(n27719), .B(n27720), .Z(n27718) );
  OR U36478 ( .A(n27721), .B(n27722), .Z(n27720) );
  IV U36479 ( .A(n27723), .Z(n27722) );
  NANDN U36480 ( .A(n27723), .B(n27721), .Z(n27717) );
  AND U36481 ( .A(n27724), .B(n27725), .Z(n27698) );
  NAND U36482 ( .A(n27726), .B(n27727), .Z(n27725) );
  NANDN U36483 ( .A(n27728), .B(n27729), .Z(n27727) );
  NANDN U36484 ( .A(n27729), .B(n27728), .Z(n27724) );
  IV U36485 ( .A(n27730), .Z(n27729) );
  NAND U36486 ( .A(n27731), .B(n27732), .Z(n27701) );
  NANDN U36487 ( .A(n27733), .B(n27734), .Z(n27732) );
  NANDN U36488 ( .A(n27735), .B(n27736), .Z(n27734) );
  NANDN U36489 ( .A(n27736), .B(n27735), .Z(n27731) );
  IV U36490 ( .A(n27737), .Z(n27735) );
  AND U36491 ( .A(n27738), .B(n27739), .Z(n27704) );
  NAND U36492 ( .A(n27740), .B(n27741), .Z(n27739) );
  NANDN U36493 ( .A(n27742), .B(n27743), .Z(n27741) );
  NANDN U36494 ( .A(n27743), .B(n27742), .Z(n27738) );
  XOR U36495 ( .A(n27714), .B(n27744), .Z(n27706) );
  XNOR U36496 ( .A(n27711), .B(n27713), .Z(n27744) );
  AND U36497 ( .A(n27745), .B(n27746), .Z(n27713) );
  NANDN U36498 ( .A(n27747), .B(n27748), .Z(n27746) );
  OR U36499 ( .A(n27749), .B(n27750), .Z(n27748) );
  IV U36500 ( .A(n27751), .Z(n27750) );
  NANDN U36501 ( .A(n27751), .B(n27749), .Z(n27745) );
  AND U36502 ( .A(n27752), .B(n27753), .Z(n27711) );
  NAND U36503 ( .A(n27754), .B(n27755), .Z(n27753) );
  NANDN U36504 ( .A(n27756), .B(n27757), .Z(n27755) );
  NANDN U36505 ( .A(n27757), .B(n27756), .Z(n27752) );
  IV U36506 ( .A(n27758), .Z(n27757) );
  NAND U36507 ( .A(n27759), .B(n27760), .Z(n27714) );
  NANDN U36508 ( .A(n27761), .B(n27762), .Z(n27760) );
  NANDN U36509 ( .A(n27763), .B(n27764), .Z(n27762) );
  NANDN U36510 ( .A(n27764), .B(n27763), .Z(n27759) );
  IV U36511 ( .A(n27765), .Z(n27763) );
  XOR U36512 ( .A(n27740), .B(n27766), .Z(N62920) );
  XNOR U36513 ( .A(n27743), .B(n27742), .Z(n27766) );
  XNOR U36514 ( .A(n27754), .B(n27767), .Z(n27742) );
  XNOR U36515 ( .A(n27758), .B(n27756), .Z(n27767) );
  XOR U36516 ( .A(n27764), .B(n27768), .Z(n27756) );
  XNOR U36517 ( .A(n27761), .B(n27765), .Z(n27768) );
  AND U36518 ( .A(n27769), .B(n27770), .Z(n27765) );
  NAND U36519 ( .A(n27771), .B(n27772), .Z(n27770) );
  NAND U36520 ( .A(n27773), .B(n27774), .Z(n27769) );
  AND U36521 ( .A(n27775), .B(n27776), .Z(n27761) );
  NAND U36522 ( .A(n27777), .B(n27778), .Z(n27776) );
  NAND U36523 ( .A(n27779), .B(n27780), .Z(n27775) );
  NANDN U36524 ( .A(n27781), .B(n27782), .Z(n27764) );
  ANDN U36525 ( .B(n27783), .A(n27784), .Z(n27758) );
  XNOR U36526 ( .A(n27749), .B(n27785), .Z(n27754) );
  XNOR U36527 ( .A(n27747), .B(n27751), .Z(n27785) );
  AND U36528 ( .A(n27786), .B(n27787), .Z(n27751) );
  NAND U36529 ( .A(n27788), .B(n27789), .Z(n27787) );
  NAND U36530 ( .A(n27790), .B(n27791), .Z(n27786) );
  AND U36531 ( .A(n27792), .B(n27793), .Z(n27747) );
  NAND U36532 ( .A(n27794), .B(n27795), .Z(n27793) );
  NAND U36533 ( .A(n27796), .B(n27797), .Z(n27792) );
  AND U36534 ( .A(n27798), .B(n27799), .Z(n27749) );
  NAND U36535 ( .A(n27800), .B(n27801), .Z(n27743) );
  XNOR U36536 ( .A(n27726), .B(n27802), .Z(n27740) );
  XNOR U36537 ( .A(n27730), .B(n27728), .Z(n27802) );
  XOR U36538 ( .A(n27736), .B(n27803), .Z(n27728) );
  XNOR U36539 ( .A(n27733), .B(n27737), .Z(n27803) );
  AND U36540 ( .A(n27804), .B(n27805), .Z(n27737) );
  NAND U36541 ( .A(n27806), .B(n27807), .Z(n27805) );
  NAND U36542 ( .A(n27808), .B(n27809), .Z(n27804) );
  AND U36543 ( .A(n27810), .B(n27811), .Z(n27733) );
  NAND U36544 ( .A(n27812), .B(n27813), .Z(n27811) );
  NAND U36545 ( .A(n27814), .B(n27815), .Z(n27810) );
  NANDN U36546 ( .A(n27816), .B(n27817), .Z(n27736) );
  ANDN U36547 ( .B(n27818), .A(n27819), .Z(n27730) );
  XNOR U36548 ( .A(n27721), .B(n27820), .Z(n27726) );
  XNOR U36549 ( .A(n27719), .B(n27723), .Z(n27820) );
  AND U36550 ( .A(n27821), .B(n27822), .Z(n27723) );
  NAND U36551 ( .A(n27823), .B(n27824), .Z(n27822) );
  NAND U36552 ( .A(n27825), .B(n27826), .Z(n27821) );
  AND U36553 ( .A(n27827), .B(n27828), .Z(n27719) );
  NAND U36554 ( .A(n27829), .B(n27830), .Z(n27828) );
  NAND U36555 ( .A(n27831), .B(n27832), .Z(n27827) );
  AND U36556 ( .A(n27833), .B(n27834), .Z(n27721) );
  XOR U36557 ( .A(n27801), .B(n27800), .Z(N62919) );
  XNOR U36558 ( .A(n27818), .B(n27819), .Z(n27800) );
  XNOR U36559 ( .A(n27833), .B(n27834), .Z(n27819) );
  XOR U36560 ( .A(n27830), .B(n27829), .Z(n27834) );
  XOR U36561 ( .A(y[4308]), .B(x[4308]), .Z(n27829) );
  XOR U36562 ( .A(n27832), .B(n27831), .Z(n27830) );
  XOR U36563 ( .A(y[4310]), .B(x[4310]), .Z(n27831) );
  XOR U36564 ( .A(y[4309]), .B(x[4309]), .Z(n27832) );
  XOR U36565 ( .A(n27824), .B(n27823), .Z(n27833) );
  XOR U36566 ( .A(n27826), .B(n27825), .Z(n27823) );
  XOR U36567 ( .A(y[4307]), .B(x[4307]), .Z(n27825) );
  XOR U36568 ( .A(y[4306]), .B(x[4306]), .Z(n27826) );
  XOR U36569 ( .A(y[4305]), .B(x[4305]), .Z(n27824) );
  XNOR U36570 ( .A(n27817), .B(n27816), .Z(n27818) );
  XNOR U36571 ( .A(n27813), .B(n27812), .Z(n27816) );
  XOR U36572 ( .A(n27815), .B(n27814), .Z(n27812) );
  XOR U36573 ( .A(y[4304]), .B(x[4304]), .Z(n27814) );
  XOR U36574 ( .A(y[4303]), .B(x[4303]), .Z(n27815) );
  XOR U36575 ( .A(y[4302]), .B(x[4302]), .Z(n27813) );
  XOR U36576 ( .A(n27807), .B(n27806), .Z(n27817) );
  XOR U36577 ( .A(n27809), .B(n27808), .Z(n27806) );
  XOR U36578 ( .A(y[4301]), .B(x[4301]), .Z(n27808) );
  XOR U36579 ( .A(y[4300]), .B(x[4300]), .Z(n27809) );
  XOR U36580 ( .A(y[4299]), .B(x[4299]), .Z(n27807) );
  XNOR U36581 ( .A(n27783), .B(n27784), .Z(n27801) );
  XNOR U36582 ( .A(n27798), .B(n27799), .Z(n27784) );
  XOR U36583 ( .A(n27795), .B(n27794), .Z(n27799) );
  XOR U36584 ( .A(y[4296]), .B(x[4296]), .Z(n27794) );
  XOR U36585 ( .A(n27797), .B(n27796), .Z(n27795) );
  XOR U36586 ( .A(y[4298]), .B(x[4298]), .Z(n27796) );
  XOR U36587 ( .A(y[4297]), .B(x[4297]), .Z(n27797) );
  XOR U36588 ( .A(n27789), .B(n27788), .Z(n27798) );
  XOR U36589 ( .A(n27791), .B(n27790), .Z(n27788) );
  XOR U36590 ( .A(y[4295]), .B(x[4295]), .Z(n27790) );
  XOR U36591 ( .A(y[4294]), .B(x[4294]), .Z(n27791) );
  XOR U36592 ( .A(y[4293]), .B(x[4293]), .Z(n27789) );
  XNOR U36593 ( .A(n27782), .B(n27781), .Z(n27783) );
  XNOR U36594 ( .A(n27778), .B(n27777), .Z(n27781) );
  XOR U36595 ( .A(n27780), .B(n27779), .Z(n27777) );
  XOR U36596 ( .A(y[4292]), .B(x[4292]), .Z(n27779) );
  XOR U36597 ( .A(y[4291]), .B(x[4291]), .Z(n27780) );
  XOR U36598 ( .A(y[4290]), .B(x[4290]), .Z(n27778) );
  XOR U36599 ( .A(n27772), .B(n27771), .Z(n27782) );
  XOR U36600 ( .A(n27774), .B(n27773), .Z(n27771) );
  XOR U36601 ( .A(y[4289]), .B(x[4289]), .Z(n27773) );
  XOR U36602 ( .A(y[4288]), .B(x[4288]), .Z(n27774) );
  XOR U36603 ( .A(y[4287]), .B(x[4287]), .Z(n27772) );
  NAND U36604 ( .A(n27835), .B(n27836), .Z(N62910) );
  NAND U36605 ( .A(n27837), .B(n27838), .Z(n27836) );
  NANDN U36606 ( .A(n27839), .B(n27840), .Z(n27838) );
  NANDN U36607 ( .A(n27840), .B(n27839), .Z(n27835) );
  XOR U36608 ( .A(n27839), .B(n27841), .Z(N62909) );
  XNOR U36609 ( .A(n27837), .B(n27840), .Z(n27841) );
  NAND U36610 ( .A(n27842), .B(n27843), .Z(n27840) );
  NAND U36611 ( .A(n27844), .B(n27845), .Z(n27843) );
  NANDN U36612 ( .A(n27846), .B(n27847), .Z(n27845) );
  NANDN U36613 ( .A(n27847), .B(n27846), .Z(n27842) );
  AND U36614 ( .A(n27848), .B(n27849), .Z(n27837) );
  NAND U36615 ( .A(n27850), .B(n27851), .Z(n27849) );
  NANDN U36616 ( .A(n27852), .B(n27853), .Z(n27851) );
  NANDN U36617 ( .A(n27853), .B(n27852), .Z(n27848) );
  IV U36618 ( .A(n27854), .Z(n27853) );
  AND U36619 ( .A(n27855), .B(n27856), .Z(n27839) );
  NAND U36620 ( .A(n27857), .B(n27858), .Z(n27856) );
  NANDN U36621 ( .A(n27859), .B(n27860), .Z(n27858) );
  NANDN U36622 ( .A(n27860), .B(n27859), .Z(n27855) );
  XOR U36623 ( .A(n27852), .B(n27861), .Z(N62908) );
  XNOR U36624 ( .A(n27850), .B(n27854), .Z(n27861) );
  XOR U36625 ( .A(n27847), .B(n27862), .Z(n27854) );
  XNOR U36626 ( .A(n27844), .B(n27846), .Z(n27862) );
  AND U36627 ( .A(n27863), .B(n27864), .Z(n27846) );
  NANDN U36628 ( .A(n27865), .B(n27866), .Z(n27864) );
  OR U36629 ( .A(n27867), .B(n27868), .Z(n27866) );
  IV U36630 ( .A(n27869), .Z(n27868) );
  NANDN U36631 ( .A(n27869), .B(n27867), .Z(n27863) );
  AND U36632 ( .A(n27870), .B(n27871), .Z(n27844) );
  NAND U36633 ( .A(n27872), .B(n27873), .Z(n27871) );
  NANDN U36634 ( .A(n27874), .B(n27875), .Z(n27873) );
  NANDN U36635 ( .A(n27875), .B(n27874), .Z(n27870) );
  IV U36636 ( .A(n27876), .Z(n27875) );
  NAND U36637 ( .A(n27877), .B(n27878), .Z(n27847) );
  NANDN U36638 ( .A(n27879), .B(n27880), .Z(n27878) );
  NANDN U36639 ( .A(n27881), .B(n27882), .Z(n27880) );
  NANDN U36640 ( .A(n27882), .B(n27881), .Z(n27877) );
  IV U36641 ( .A(n27883), .Z(n27881) );
  AND U36642 ( .A(n27884), .B(n27885), .Z(n27850) );
  NAND U36643 ( .A(n27886), .B(n27887), .Z(n27885) );
  NANDN U36644 ( .A(n27888), .B(n27889), .Z(n27887) );
  NANDN U36645 ( .A(n27889), .B(n27888), .Z(n27884) );
  XOR U36646 ( .A(n27860), .B(n27890), .Z(n27852) );
  XNOR U36647 ( .A(n27857), .B(n27859), .Z(n27890) );
  AND U36648 ( .A(n27891), .B(n27892), .Z(n27859) );
  NANDN U36649 ( .A(n27893), .B(n27894), .Z(n27892) );
  OR U36650 ( .A(n27895), .B(n27896), .Z(n27894) );
  IV U36651 ( .A(n27897), .Z(n27896) );
  NANDN U36652 ( .A(n27897), .B(n27895), .Z(n27891) );
  AND U36653 ( .A(n27898), .B(n27899), .Z(n27857) );
  NAND U36654 ( .A(n27900), .B(n27901), .Z(n27899) );
  NANDN U36655 ( .A(n27902), .B(n27903), .Z(n27901) );
  NANDN U36656 ( .A(n27903), .B(n27902), .Z(n27898) );
  IV U36657 ( .A(n27904), .Z(n27903) );
  NAND U36658 ( .A(n27905), .B(n27906), .Z(n27860) );
  NANDN U36659 ( .A(n27907), .B(n27908), .Z(n27906) );
  NANDN U36660 ( .A(n27909), .B(n27910), .Z(n27908) );
  NANDN U36661 ( .A(n27910), .B(n27909), .Z(n27905) );
  IV U36662 ( .A(n27911), .Z(n27909) );
  XOR U36663 ( .A(n27886), .B(n27912), .Z(N62907) );
  XNOR U36664 ( .A(n27889), .B(n27888), .Z(n27912) );
  XNOR U36665 ( .A(n27900), .B(n27913), .Z(n27888) );
  XNOR U36666 ( .A(n27904), .B(n27902), .Z(n27913) );
  XOR U36667 ( .A(n27910), .B(n27914), .Z(n27902) );
  XNOR U36668 ( .A(n27907), .B(n27911), .Z(n27914) );
  AND U36669 ( .A(n27915), .B(n27916), .Z(n27911) );
  NAND U36670 ( .A(n27917), .B(n27918), .Z(n27916) );
  NAND U36671 ( .A(n27919), .B(n27920), .Z(n27915) );
  AND U36672 ( .A(n27921), .B(n27922), .Z(n27907) );
  NAND U36673 ( .A(n27923), .B(n27924), .Z(n27922) );
  NAND U36674 ( .A(n27925), .B(n27926), .Z(n27921) );
  NANDN U36675 ( .A(n27927), .B(n27928), .Z(n27910) );
  ANDN U36676 ( .B(n27929), .A(n27930), .Z(n27904) );
  XNOR U36677 ( .A(n27895), .B(n27931), .Z(n27900) );
  XNOR U36678 ( .A(n27893), .B(n27897), .Z(n27931) );
  AND U36679 ( .A(n27932), .B(n27933), .Z(n27897) );
  NAND U36680 ( .A(n27934), .B(n27935), .Z(n27933) );
  NAND U36681 ( .A(n27936), .B(n27937), .Z(n27932) );
  AND U36682 ( .A(n27938), .B(n27939), .Z(n27893) );
  NAND U36683 ( .A(n27940), .B(n27941), .Z(n27939) );
  NAND U36684 ( .A(n27942), .B(n27943), .Z(n27938) );
  AND U36685 ( .A(n27944), .B(n27945), .Z(n27895) );
  NAND U36686 ( .A(n27946), .B(n27947), .Z(n27889) );
  XNOR U36687 ( .A(n27872), .B(n27948), .Z(n27886) );
  XNOR U36688 ( .A(n27876), .B(n27874), .Z(n27948) );
  XOR U36689 ( .A(n27882), .B(n27949), .Z(n27874) );
  XNOR U36690 ( .A(n27879), .B(n27883), .Z(n27949) );
  AND U36691 ( .A(n27950), .B(n27951), .Z(n27883) );
  NAND U36692 ( .A(n27952), .B(n27953), .Z(n27951) );
  NAND U36693 ( .A(n27954), .B(n27955), .Z(n27950) );
  AND U36694 ( .A(n27956), .B(n27957), .Z(n27879) );
  NAND U36695 ( .A(n27958), .B(n27959), .Z(n27957) );
  NAND U36696 ( .A(n27960), .B(n27961), .Z(n27956) );
  NANDN U36697 ( .A(n27962), .B(n27963), .Z(n27882) );
  ANDN U36698 ( .B(n27964), .A(n27965), .Z(n27876) );
  XNOR U36699 ( .A(n27867), .B(n27966), .Z(n27872) );
  XNOR U36700 ( .A(n27865), .B(n27869), .Z(n27966) );
  AND U36701 ( .A(n27967), .B(n27968), .Z(n27869) );
  NAND U36702 ( .A(n27969), .B(n27970), .Z(n27968) );
  NAND U36703 ( .A(n27971), .B(n27972), .Z(n27967) );
  AND U36704 ( .A(n27973), .B(n27974), .Z(n27865) );
  NAND U36705 ( .A(n27975), .B(n27976), .Z(n27974) );
  NAND U36706 ( .A(n27977), .B(n27978), .Z(n27973) );
  AND U36707 ( .A(n27979), .B(n27980), .Z(n27867) );
  XOR U36708 ( .A(n27947), .B(n27946), .Z(N62906) );
  XNOR U36709 ( .A(n27964), .B(n27965), .Z(n27946) );
  XNOR U36710 ( .A(n27979), .B(n27980), .Z(n27965) );
  XOR U36711 ( .A(n27976), .B(n27975), .Z(n27980) );
  XOR U36712 ( .A(y[4284]), .B(x[4284]), .Z(n27975) );
  XOR U36713 ( .A(n27978), .B(n27977), .Z(n27976) );
  XOR U36714 ( .A(y[4286]), .B(x[4286]), .Z(n27977) );
  XOR U36715 ( .A(y[4285]), .B(x[4285]), .Z(n27978) );
  XOR U36716 ( .A(n27970), .B(n27969), .Z(n27979) );
  XOR U36717 ( .A(n27972), .B(n27971), .Z(n27969) );
  XOR U36718 ( .A(y[4283]), .B(x[4283]), .Z(n27971) );
  XOR U36719 ( .A(y[4282]), .B(x[4282]), .Z(n27972) );
  XOR U36720 ( .A(y[4281]), .B(x[4281]), .Z(n27970) );
  XNOR U36721 ( .A(n27963), .B(n27962), .Z(n27964) );
  XNOR U36722 ( .A(n27959), .B(n27958), .Z(n27962) );
  XOR U36723 ( .A(n27961), .B(n27960), .Z(n27958) );
  XOR U36724 ( .A(y[4280]), .B(x[4280]), .Z(n27960) );
  XOR U36725 ( .A(y[4279]), .B(x[4279]), .Z(n27961) );
  XOR U36726 ( .A(y[4278]), .B(x[4278]), .Z(n27959) );
  XOR U36727 ( .A(n27953), .B(n27952), .Z(n27963) );
  XOR U36728 ( .A(n27955), .B(n27954), .Z(n27952) );
  XOR U36729 ( .A(y[4277]), .B(x[4277]), .Z(n27954) );
  XOR U36730 ( .A(y[4276]), .B(x[4276]), .Z(n27955) );
  XOR U36731 ( .A(y[4275]), .B(x[4275]), .Z(n27953) );
  XNOR U36732 ( .A(n27929), .B(n27930), .Z(n27947) );
  XNOR U36733 ( .A(n27944), .B(n27945), .Z(n27930) );
  XOR U36734 ( .A(n27941), .B(n27940), .Z(n27945) );
  XOR U36735 ( .A(y[4272]), .B(x[4272]), .Z(n27940) );
  XOR U36736 ( .A(n27943), .B(n27942), .Z(n27941) );
  XOR U36737 ( .A(y[4274]), .B(x[4274]), .Z(n27942) );
  XOR U36738 ( .A(y[4273]), .B(x[4273]), .Z(n27943) );
  XOR U36739 ( .A(n27935), .B(n27934), .Z(n27944) );
  XOR U36740 ( .A(n27937), .B(n27936), .Z(n27934) );
  XOR U36741 ( .A(y[4271]), .B(x[4271]), .Z(n27936) );
  XOR U36742 ( .A(y[4270]), .B(x[4270]), .Z(n27937) );
  XOR U36743 ( .A(y[4269]), .B(x[4269]), .Z(n27935) );
  XNOR U36744 ( .A(n27928), .B(n27927), .Z(n27929) );
  XNOR U36745 ( .A(n27924), .B(n27923), .Z(n27927) );
  XOR U36746 ( .A(n27926), .B(n27925), .Z(n27923) );
  XOR U36747 ( .A(y[4268]), .B(x[4268]), .Z(n27925) );
  XOR U36748 ( .A(y[4267]), .B(x[4267]), .Z(n27926) );
  XOR U36749 ( .A(y[4266]), .B(x[4266]), .Z(n27924) );
  XOR U36750 ( .A(n27918), .B(n27917), .Z(n27928) );
  XOR U36751 ( .A(n27920), .B(n27919), .Z(n27917) );
  XOR U36752 ( .A(y[4265]), .B(x[4265]), .Z(n27919) );
  XOR U36753 ( .A(y[4264]), .B(x[4264]), .Z(n27920) );
  XOR U36754 ( .A(y[4263]), .B(x[4263]), .Z(n27918) );
  NAND U36755 ( .A(n27981), .B(n27982), .Z(N62897) );
  NAND U36756 ( .A(n27983), .B(n27984), .Z(n27982) );
  NANDN U36757 ( .A(n27985), .B(n27986), .Z(n27984) );
  NANDN U36758 ( .A(n27986), .B(n27985), .Z(n27981) );
  XOR U36759 ( .A(n27985), .B(n27987), .Z(N62896) );
  XNOR U36760 ( .A(n27983), .B(n27986), .Z(n27987) );
  NAND U36761 ( .A(n27988), .B(n27989), .Z(n27986) );
  NAND U36762 ( .A(n27990), .B(n27991), .Z(n27989) );
  NANDN U36763 ( .A(n27992), .B(n27993), .Z(n27991) );
  NANDN U36764 ( .A(n27993), .B(n27992), .Z(n27988) );
  AND U36765 ( .A(n27994), .B(n27995), .Z(n27983) );
  NAND U36766 ( .A(n27996), .B(n27997), .Z(n27995) );
  NANDN U36767 ( .A(n27998), .B(n27999), .Z(n27997) );
  NANDN U36768 ( .A(n27999), .B(n27998), .Z(n27994) );
  IV U36769 ( .A(n28000), .Z(n27999) );
  AND U36770 ( .A(n28001), .B(n28002), .Z(n27985) );
  NAND U36771 ( .A(n28003), .B(n28004), .Z(n28002) );
  NANDN U36772 ( .A(n28005), .B(n28006), .Z(n28004) );
  NANDN U36773 ( .A(n28006), .B(n28005), .Z(n28001) );
  XOR U36774 ( .A(n27998), .B(n28007), .Z(N62895) );
  XNOR U36775 ( .A(n27996), .B(n28000), .Z(n28007) );
  XOR U36776 ( .A(n27993), .B(n28008), .Z(n28000) );
  XNOR U36777 ( .A(n27990), .B(n27992), .Z(n28008) );
  AND U36778 ( .A(n28009), .B(n28010), .Z(n27992) );
  NANDN U36779 ( .A(n28011), .B(n28012), .Z(n28010) );
  OR U36780 ( .A(n28013), .B(n28014), .Z(n28012) );
  IV U36781 ( .A(n28015), .Z(n28014) );
  NANDN U36782 ( .A(n28015), .B(n28013), .Z(n28009) );
  AND U36783 ( .A(n28016), .B(n28017), .Z(n27990) );
  NAND U36784 ( .A(n28018), .B(n28019), .Z(n28017) );
  NANDN U36785 ( .A(n28020), .B(n28021), .Z(n28019) );
  NANDN U36786 ( .A(n28021), .B(n28020), .Z(n28016) );
  IV U36787 ( .A(n28022), .Z(n28021) );
  NAND U36788 ( .A(n28023), .B(n28024), .Z(n27993) );
  NANDN U36789 ( .A(n28025), .B(n28026), .Z(n28024) );
  NANDN U36790 ( .A(n28027), .B(n28028), .Z(n28026) );
  NANDN U36791 ( .A(n28028), .B(n28027), .Z(n28023) );
  IV U36792 ( .A(n28029), .Z(n28027) );
  AND U36793 ( .A(n28030), .B(n28031), .Z(n27996) );
  NAND U36794 ( .A(n28032), .B(n28033), .Z(n28031) );
  NANDN U36795 ( .A(n28034), .B(n28035), .Z(n28033) );
  NANDN U36796 ( .A(n28035), .B(n28034), .Z(n28030) );
  XOR U36797 ( .A(n28006), .B(n28036), .Z(n27998) );
  XNOR U36798 ( .A(n28003), .B(n28005), .Z(n28036) );
  AND U36799 ( .A(n28037), .B(n28038), .Z(n28005) );
  NANDN U36800 ( .A(n28039), .B(n28040), .Z(n28038) );
  OR U36801 ( .A(n28041), .B(n28042), .Z(n28040) );
  IV U36802 ( .A(n28043), .Z(n28042) );
  NANDN U36803 ( .A(n28043), .B(n28041), .Z(n28037) );
  AND U36804 ( .A(n28044), .B(n28045), .Z(n28003) );
  NAND U36805 ( .A(n28046), .B(n28047), .Z(n28045) );
  NANDN U36806 ( .A(n28048), .B(n28049), .Z(n28047) );
  NANDN U36807 ( .A(n28049), .B(n28048), .Z(n28044) );
  IV U36808 ( .A(n28050), .Z(n28049) );
  NAND U36809 ( .A(n28051), .B(n28052), .Z(n28006) );
  NANDN U36810 ( .A(n28053), .B(n28054), .Z(n28052) );
  NANDN U36811 ( .A(n28055), .B(n28056), .Z(n28054) );
  NANDN U36812 ( .A(n28056), .B(n28055), .Z(n28051) );
  IV U36813 ( .A(n28057), .Z(n28055) );
  XOR U36814 ( .A(n28032), .B(n28058), .Z(N62894) );
  XNOR U36815 ( .A(n28035), .B(n28034), .Z(n28058) );
  XNOR U36816 ( .A(n28046), .B(n28059), .Z(n28034) );
  XNOR U36817 ( .A(n28050), .B(n28048), .Z(n28059) );
  XOR U36818 ( .A(n28056), .B(n28060), .Z(n28048) );
  XNOR U36819 ( .A(n28053), .B(n28057), .Z(n28060) );
  AND U36820 ( .A(n28061), .B(n28062), .Z(n28057) );
  NAND U36821 ( .A(n28063), .B(n28064), .Z(n28062) );
  NAND U36822 ( .A(n28065), .B(n28066), .Z(n28061) );
  AND U36823 ( .A(n28067), .B(n28068), .Z(n28053) );
  NAND U36824 ( .A(n28069), .B(n28070), .Z(n28068) );
  NAND U36825 ( .A(n28071), .B(n28072), .Z(n28067) );
  NANDN U36826 ( .A(n28073), .B(n28074), .Z(n28056) );
  ANDN U36827 ( .B(n28075), .A(n28076), .Z(n28050) );
  XNOR U36828 ( .A(n28041), .B(n28077), .Z(n28046) );
  XNOR U36829 ( .A(n28039), .B(n28043), .Z(n28077) );
  AND U36830 ( .A(n28078), .B(n28079), .Z(n28043) );
  NAND U36831 ( .A(n28080), .B(n28081), .Z(n28079) );
  NAND U36832 ( .A(n28082), .B(n28083), .Z(n28078) );
  AND U36833 ( .A(n28084), .B(n28085), .Z(n28039) );
  NAND U36834 ( .A(n28086), .B(n28087), .Z(n28085) );
  NAND U36835 ( .A(n28088), .B(n28089), .Z(n28084) );
  AND U36836 ( .A(n28090), .B(n28091), .Z(n28041) );
  NAND U36837 ( .A(n28092), .B(n28093), .Z(n28035) );
  XNOR U36838 ( .A(n28018), .B(n28094), .Z(n28032) );
  XNOR U36839 ( .A(n28022), .B(n28020), .Z(n28094) );
  XOR U36840 ( .A(n28028), .B(n28095), .Z(n28020) );
  XNOR U36841 ( .A(n28025), .B(n28029), .Z(n28095) );
  AND U36842 ( .A(n28096), .B(n28097), .Z(n28029) );
  NAND U36843 ( .A(n28098), .B(n28099), .Z(n28097) );
  NAND U36844 ( .A(n28100), .B(n28101), .Z(n28096) );
  AND U36845 ( .A(n28102), .B(n28103), .Z(n28025) );
  NAND U36846 ( .A(n28104), .B(n28105), .Z(n28103) );
  NAND U36847 ( .A(n28106), .B(n28107), .Z(n28102) );
  NANDN U36848 ( .A(n28108), .B(n28109), .Z(n28028) );
  ANDN U36849 ( .B(n28110), .A(n28111), .Z(n28022) );
  XNOR U36850 ( .A(n28013), .B(n28112), .Z(n28018) );
  XNOR U36851 ( .A(n28011), .B(n28015), .Z(n28112) );
  AND U36852 ( .A(n28113), .B(n28114), .Z(n28015) );
  NAND U36853 ( .A(n28115), .B(n28116), .Z(n28114) );
  NAND U36854 ( .A(n28117), .B(n28118), .Z(n28113) );
  AND U36855 ( .A(n28119), .B(n28120), .Z(n28011) );
  NAND U36856 ( .A(n28121), .B(n28122), .Z(n28120) );
  NAND U36857 ( .A(n28123), .B(n28124), .Z(n28119) );
  AND U36858 ( .A(n28125), .B(n28126), .Z(n28013) );
  XOR U36859 ( .A(n28093), .B(n28092), .Z(N62893) );
  XNOR U36860 ( .A(n28110), .B(n28111), .Z(n28092) );
  XNOR U36861 ( .A(n28125), .B(n28126), .Z(n28111) );
  XOR U36862 ( .A(n28122), .B(n28121), .Z(n28126) );
  XOR U36863 ( .A(y[4260]), .B(x[4260]), .Z(n28121) );
  XOR U36864 ( .A(n28124), .B(n28123), .Z(n28122) );
  XOR U36865 ( .A(y[4262]), .B(x[4262]), .Z(n28123) );
  XOR U36866 ( .A(y[4261]), .B(x[4261]), .Z(n28124) );
  XOR U36867 ( .A(n28116), .B(n28115), .Z(n28125) );
  XOR U36868 ( .A(n28118), .B(n28117), .Z(n28115) );
  XOR U36869 ( .A(y[4259]), .B(x[4259]), .Z(n28117) );
  XOR U36870 ( .A(y[4258]), .B(x[4258]), .Z(n28118) );
  XOR U36871 ( .A(y[4257]), .B(x[4257]), .Z(n28116) );
  XNOR U36872 ( .A(n28109), .B(n28108), .Z(n28110) );
  XNOR U36873 ( .A(n28105), .B(n28104), .Z(n28108) );
  XOR U36874 ( .A(n28107), .B(n28106), .Z(n28104) );
  XOR U36875 ( .A(y[4256]), .B(x[4256]), .Z(n28106) );
  XOR U36876 ( .A(y[4255]), .B(x[4255]), .Z(n28107) );
  XOR U36877 ( .A(y[4254]), .B(x[4254]), .Z(n28105) );
  XOR U36878 ( .A(n28099), .B(n28098), .Z(n28109) );
  XOR U36879 ( .A(n28101), .B(n28100), .Z(n28098) );
  XOR U36880 ( .A(y[4253]), .B(x[4253]), .Z(n28100) );
  XOR U36881 ( .A(y[4252]), .B(x[4252]), .Z(n28101) );
  XOR U36882 ( .A(y[4251]), .B(x[4251]), .Z(n28099) );
  XNOR U36883 ( .A(n28075), .B(n28076), .Z(n28093) );
  XNOR U36884 ( .A(n28090), .B(n28091), .Z(n28076) );
  XOR U36885 ( .A(n28087), .B(n28086), .Z(n28091) );
  XOR U36886 ( .A(y[4248]), .B(x[4248]), .Z(n28086) );
  XOR U36887 ( .A(n28089), .B(n28088), .Z(n28087) );
  XOR U36888 ( .A(y[4250]), .B(x[4250]), .Z(n28088) );
  XOR U36889 ( .A(y[4249]), .B(x[4249]), .Z(n28089) );
  XOR U36890 ( .A(n28081), .B(n28080), .Z(n28090) );
  XOR U36891 ( .A(n28083), .B(n28082), .Z(n28080) );
  XOR U36892 ( .A(y[4247]), .B(x[4247]), .Z(n28082) );
  XOR U36893 ( .A(y[4246]), .B(x[4246]), .Z(n28083) );
  XOR U36894 ( .A(y[4245]), .B(x[4245]), .Z(n28081) );
  XNOR U36895 ( .A(n28074), .B(n28073), .Z(n28075) );
  XNOR U36896 ( .A(n28070), .B(n28069), .Z(n28073) );
  XOR U36897 ( .A(n28072), .B(n28071), .Z(n28069) );
  XOR U36898 ( .A(y[4244]), .B(x[4244]), .Z(n28071) );
  XOR U36899 ( .A(y[4243]), .B(x[4243]), .Z(n28072) );
  XOR U36900 ( .A(y[4242]), .B(x[4242]), .Z(n28070) );
  XOR U36901 ( .A(n28064), .B(n28063), .Z(n28074) );
  XOR U36902 ( .A(n28066), .B(n28065), .Z(n28063) );
  XOR U36903 ( .A(y[4241]), .B(x[4241]), .Z(n28065) );
  XOR U36904 ( .A(y[4240]), .B(x[4240]), .Z(n28066) );
  XOR U36905 ( .A(y[4239]), .B(x[4239]), .Z(n28064) );
  NAND U36906 ( .A(n28127), .B(n28128), .Z(N62884) );
  NAND U36907 ( .A(n28129), .B(n28130), .Z(n28128) );
  NANDN U36908 ( .A(n28131), .B(n28132), .Z(n28130) );
  NANDN U36909 ( .A(n28132), .B(n28131), .Z(n28127) );
  XOR U36910 ( .A(n28131), .B(n28133), .Z(N62883) );
  XNOR U36911 ( .A(n28129), .B(n28132), .Z(n28133) );
  NAND U36912 ( .A(n28134), .B(n28135), .Z(n28132) );
  NAND U36913 ( .A(n28136), .B(n28137), .Z(n28135) );
  NANDN U36914 ( .A(n28138), .B(n28139), .Z(n28137) );
  NANDN U36915 ( .A(n28139), .B(n28138), .Z(n28134) );
  AND U36916 ( .A(n28140), .B(n28141), .Z(n28129) );
  NAND U36917 ( .A(n28142), .B(n28143), .Z(n28141) );
  NANDN U36918 ( .A(n28144), .B(n28145), .Z(n28143) );
  NANDN U36919 ( .A(n28145), .B(n28144), .Z(n28140) );
  IV U36920 ( .A(n28146), .Z(n28145) );
  AND U36921 ( .A(n28147), .B(n28148), .Z(n28131) );
  NAND U36922 ( .A(n28149), .B(n28150), .Z(n28148) );
  NANDN U36923 ( .A(n28151), .B(n28152), .Z(n28150) );
  NANDN U36924 ( .A(n28152), .B(n28151), .Z(n28147) );
  XOR U36925 ( .A(n28144), .B(n28153), .Z(N62882) );
  XNOR U36926 ( .A(n28142), .B(n28146), .Z(n28153) );
  XOR U36927 ( .A(n28139), .B(n28154), .Z(n28146) );
  XNOR U36928 ( .A(n28136), .B(n28138), .Z(n28154) );
  AND U36929 ( .A(n28155), .B(n28156), .Z(n28138) );
  NANDN U36930 ( .A(n28157), .B(n28158), .Z(n28156) );
  OR U36931 ( .A(n28159), .B(n28160), .Z(n28158) );
  IV U36932 ( .A(n28161), .Z(n28160) );
  NANDN U36933 ( .A(n28161), .B(n28159), .Z(n28155) );
  AND U36934 ( .A(n28162), .B(n28163), .Z(n28136) );
  NAND U36935 ( .A(n28164), .B(n28165), .Z(n28163) );
  NANDN U36936 ( .A(n28166), .B(n28167), .Z(n28165) );
  NANDN U36937 ( .A(n28167), .B(n28166), .Z(n28162) );
  IV U36938 ( .A(n28168), .Z(n28167) );
  NAND U36939 ( .A(n28169), .B(n28170), .Z(n28139) );
  NANDN U36940 ( .A(n28171), .B(n28172), .Z(n28170) );
  NANDN U36941 ( .A(n28173), .B(n28174), .Z(n28172) );
  NANDN U36942 ( .A(n28174), .B(n28173), .Z(n28169) );
  IV U36943 ( .A(n28175), .Z(n28173) );
  AND U36944 ( .A(n28176), .B(n28177), .Z(n28142) );
  NAND U36945 ( .A(n28178), .B(n28179), .Z(n28177) );
  NANDN U36946 ( .A(n28180), .B(n28181), .Z(n28179) );
  NANDN U36947 ( .A(n28181), .B(n28180), .Z(n28176) );
  XOR U36948 ( .A(n28152), .B(n28182), .Z(n28144) );
  XNOR U36949 ( .A(n28149), .B(n28151), .Z(n28182) );
  AND U36950 ( .A(n28183), .B(n28184), .Z(n28151) );
  NANDN U36951 ( .A(n28185), .B(n28186), .Z(n28184) );
  OR U36952 ( .A(n28187), .B(n28188), .Z(n28186) );
  IV U36953 ( .A(n28189), .Z(n28188) );
  NANDN U36954 ( .A(n28189), .B(n28187), .Z(n28183) );
  AND U36955 ( .A(n28190), .B(n28191), .Z(n28149) );
  NAND U36956 ( .A(n28192), .B(n28193), .Z(n28191) );
  NANDN U36957 ( .A(n28194), .B(n28195), .Z(n28193) );
  NANDN U36958 ( .A(n28195), .B(n28194), .Z(n28190) );
  IV U36959 ( .A(n28196), .Z(n28195) );
  NAND U36960 ( .A(n28197), .B(n28198), .Z(n28152) );
  NANDN U36961 ( .A(n28199), .B(n28200), .Z(n28198) );
  NANDN U36962 ( .A(n28201), .B(n28202), .Z(n28200) );
  NANDN U36963 ( .A(n28202), .B(n28201), .Z(n28197) );
  IV U36964 ( .A(n28203), .Z(n28201) );
  XOR U36965 ( .A(n28178), .B(n28204), .Z(N62881) );
  XNOR U36966 ( .A(n28181), .B(n28180), .Z(n28204) );
  XNOR U36967 ( .A(n28192), .B(n28205), .Z(n28180) );
  XNOR U36968 ( .A(n28196), .B(n28194), .Z(n28205) );
  XOR U36969 ( .A(n28202), .B(n28206), .Z(n28194) );
  XNOR U36970 ( .A(n28199), .B(n28203), .Z(n28206) );
  AND U36971 ( .A(n28207), .B(n28208), .Z(n28203) );
  NAND U36972 ( .A(n28209), .B(n28210), .Z(n28208) );
  NAND U36973 ( .A(n28211), .B(n28212), .Z(n28207) );
  AND U36974 ( .A(n28213), .B(n28214), .Z(n28199) );
  NAND U36975 ( .A(n28215), .B(n28216), .Z(n28214) );
  NAND U36976 ( .A(n28217), .B(n28218), .Z(n28213) );
  NANDN U36977 ( .A(n28219), .B(n28220), .Z(n28202) );
  ANDN U36978 ( .B(n28221), .A(n28222), .Z(n28196) );
  XNOR U36979 ( .A(n28187), .B(n28223), .Z(n28192) );
  XNOR U36980 ( .A(n28185), .B(n28189), .Z(n28223) );
  AND U36981 ( .A(n28224), .B(n28225), .Z(n28189) );
  NAND U36982 ( .A(n28226), .B(n28227), .Z(n28225) );
  NAND U36983 ( .A(n28228), .B(n28229), .Z(n28224) );
  AND U36984 ( .A(n28230), .B(n28231), .Z(n28185) );
  NAND U36985 ( .A(n28232), .B(n28233), .Z(n28231) );
  NAND U36986 ( .A(n28234), .B(n28235), .Z(n28230) );
  AND U36987 ( .A(n28236), .B(n28237), .Z(n28187) );
  NAND U36988 ( .A(n28238), .B(n28239), .Z(n28181) );
  XNOR U36989 ( .A(n28164), .B(n28240), .Z(n28178) );
  XNOR U36990 ( .A(n28168), .B(n28166), .Z(n28240) );
  XOR U36991 ( .A(n28174), .B(n28241), .Z(n28166) );
  XNOR U36992 ( .A(n28171), .B(n28175), .Z(n28241) );
  AND U36993 ( .A(n28242), .B(n28243), .Z(n28175) );
  NAND U36994 ( .A(n28244), .B(n28245), .Z(n28243) );
  NAND U36995 ( .A(n28246), .B(n28247), .Z(n28242) );
  AND U36996 ( .A(n28248), .B(n28249), .Z(n28171) );
  NAND U36997 ( .A(n28250), .B(n28251), .Z(n28249) );
  NAND U36998 ( .A(n28252), .B(n28253), .Z(n28248) );
  NANDN U36999 ( .A(n28254), .B(n28255), .Z(n28174) );
  ANDN U37000 ( .B(n28256), .A(n28257), .Z(n28168) );
  XNOR U37001 ( .A(n28159), .B(n28258), .Z(n28164) );
  XNOR U37002 ( .A(n28157), .B(n28161), .Z(n28258) );
  AND U37003 ( .A(n28259), .B(n28260), .Z(n28161) );
  NAND U37004 ( .A(n28261), .B(n28262), .Z(n28260) );
  NAND U37005 ( .A(n28263), .B(n28264), .Z(n28259) );
  AND U37006 ( .A(n28265), .B(n28266), .Z(n28157) );
  NAND U37007 ( .A(n28267), .B(n28268), .Z(n28266) );
  NAND U37008 ( .A(n28269), .B(n28270), .Z(n28265) );
  AND U37009 ( .A(n28271), .B(n28272), .Z(n28159) );
  XOR U37010 ( .A(n28239), .B(n28238), .Z(N62880) );
  XNOR U37011 ( .A(n28256), .B(n28257), .Z(n28238) );
  XNOR U37012 ( .A(n28271), .B(n28272), .Z(n28257) );
  XOR U37013 ( .A(n28268), .B(n28267), .Z(n28272) );
  XOR U37014 ( .A(y[4236]), .B(x[4236]), .Z(n28267) );
  XOR U37015 ( .A(n28270), .B(n28269), .Z(n28268) );
  XOR U37016 ( .A(y[4238]), .B(x[4238]), .Z(n28269) );
  XOR U37017 ( .A(y[4237]), .B(x[4237]), .Z(n28270) );
  XOR U37018 ( .A(n28262), .B(n28261), .Z(n28271) );
  XOR U37019 ( .A(n28264), .B(n28263), .Z(n28261) );
  XOR U37020 ( .A(y[4235]), .B(x[4235]), .Z(n28263) );
  XOR U37021 ( .A(y[4234]), .B(x[4234]), .Z(n28264) );
  XOR U37022 ( .A(y[4233]), .B(x[4233]), .Z(n28262) );
  XNOR U37023 ( .A(n28255), .B(n28254), .Z(n28256) );
  XNOR U37024 ( .A(n28251), .B(n28250), .Z(n28254) );
  XOR U37025 ( .A(n28253), .B(n28252), .Z(n28250) );
  XOR U37026 ( .A(y[4232]), .B(x[4232]), .Z(n28252) );
  XOR U37027 ( .A(y[4231]), .B(x[4231]), .Z(n28253) );
  XOR U37028 ( .A(y[4230]), .B(x[4230]), .Z(n28251) );
  XOR U37029 ( .A(n28245), .B(n28244), .Z(n28255) );
  XOR U37030 ( .A(n28247), .B(n28246), .Z(n28244) );
  XOR U37031 ( .A(y[4229]), .B(x[4229]), .Z(n28246) );
  XOR U37032 ( .A(y[4228]), .B(x[4228]), .Z(n28247) );
  XOR U37033 ( .A(y[4227]), .B(x[4227]), .Z(n28245) );
  XNOR U37034 ( .A(n28221), .B(n28222), .Z(n28239) );
  XNOR U37035 ( .A(n28236), .B(n28237), .Z(n28222) );
  XOR U37036 ( .A(n28233), .B(n28232), .Z(n28237) );
  XOR U37037 ( .A(y[4224]), .B(x[4224]), .Z(n28232) );
  XOR U37038 ( .A(n28235), .B(n28234), .Z(n28233) );
  XOR U37039 ( .A(y[4226]), .B(x[4226]), .Z(n28234) );
  XOR U37040 ( .A(y[4225]), .B(x[4225]), .Z(n28235) );
  XOR U37041 ( .A(n28227), .B(n28226), .Z(n28236) );
  XOR U37042 ( .A(n28229), .B(n28228), .Z(n28226) );
  XOR U37043 ( .A(y[4223]), .B(x[4223]), .Z(n28228) );
  XOR U37044 ( .A(y[4222]), .B(x[4222]), .Z(n28229) );
  XOR U37045 ( .A(y[4221]), .B(x[4221]), .Z(n28227) );
  XNOR U37046 ( .A(n28220), .B(n28219), .Z(n28221) );
  XNOR U37047 ( .A(n28216), .B(n28215), .Z(n28219) );
  XOR U37048 ( .A(n28218), .B(n28217), .Z(n28215) );
  XOR U37049 ( .A(y[4220]), .B(x[4220]), .Z(n28217) );
  XOR U37050 ( .A(y[4219]), .B(x[4219]), .Z(n28218) );
  XOR U37051 ( .A(y[4218]), .B(x[4218]), .Z(n28216) );
  XOR U37052 ( .A(n28210), .B(n28209), .Z(n28220) );
  XOR U37053 ( .A(n28212), .B(n28211), .Z(n28209) );
  XOR U37054 ( .A(y[4217]), .B(x[4217]), .Z(n28211) );
  XOR U37055 ( .A(y[4216]), .B(x[4216]), .Z(n28212) );
  XOR U37056 ( .A(y[4215]), .B(x[4215]), .Z(n28210) );
  NAND U37057 ( .A(n28273), .B(n28274), .Z(N62871) );
  NAND U37058 ( .A(n28275), .B(n28276), .Z(n28274) );
  NANDN U37059 ( .A(n28277), .B(n28278), .Z(n28276) );
  NANDN U37060 ( .A(n28278), .B(n28277), .Z(n28273) );
  XOR U37061 ( .A(n28277), .B(n28279), .Z(N62870) );
  XNOR U37062 ( .A(n28275), .B(n28278), .Z(n28279) );
  NAND U37063 ( .A(n28280), .B(n28281), .Z(n28278) );
  NAND U37064 ( .A(n28282), .B(n28283), .Z(n28281) );
  NANDN U37065 ( .A(n28284), .B(n28285), .Z(n28283) );
  NANDN U37066 ( .A(n28285), .B(n28284), .Z(n28280) );
  AND U37067 ( .A(n28286), .B(n28287), .Z(n28275) );
  NAND U37068 ( .A(n28288), .B(n28289), .Z(n28287) );
  NANDN U37069 ( .A(n28290), .B(n28291), .Z(n28289) );
  NANDN U37070 ( .A(n28291), .B(n28290), .Z(n28286) );
  IV U37071 ( .A(n28292), .Z(n28291) );
  AND U37072 ( .A(n28293), .B(n28294), .Z(n28277) );
  NAND U37073 ( .A(n28295), .B(n28296), .Z(n28294) );
  NANDN U37074 ( .A(n28297), .B(n28298), .Z(n28296) );
  NANDN U37075 ( .A(n28298), .B(n28297), .Z(n28293) );
  XOR U37076 ( .A(n28290), .B(n28299), .Z(N62869) );
  XNOR U37077 ( .A(n28288), .B(n28292), .Z(n28299) );
  XOR U37078 ( .A(n28285), .B(n28300), .Z(n28292) );
  XNOR U37079 ( .A(n28282), .B(n28284), .Z(n28300) );
  AND U37080 ( .A(n28301), .B(n28302), .Z(n28284) );
  NANDN U37081 ( .A(n28303), .B(n28304), .Z(n28302) );
  OR U37082 ( .A(n28305), .B(n28306), .Z(n28304) );
  IV U37083 ( .A(n28307), .Z(n28306) );
  NANDN U37084 ( .A(n28307), .B(n28305), .Z(n28301) );
  AND U37085 ( .A(n28308), .B(n28309), .Z(n28282) );
  NAND U37086 ( .A(n28310), .B(n28311), .Z(n28309) );
  NANDN U37087 ( .A(n28312), .B(n28313), .Z(n28311) );
  NANDN U37088 ( .A(n28313), .B(n28312), .Z(n28308) );
  IV U37089 ( .A(n28314), .Z(n28313) );
  NAND U37090 ( .A(n28315), .B(n28316), .Z(n28285) );
  NANDN U37091 ( .A(n28317), .B(n28318), .Z(n28316) );
  NANDN U37092 ( .A(n28319), .B(n28320), .Z(n28318) );
  NANDN U37093 ( .A(n28320), .B(n28319), .Z(n28315) );
  IV U37094 ( .A(n28321), .Z(n28319) );
  AND U37095 ( .A(n28322), .B(n28323), .Z(n28288) );
  NAND U37096 ( .A(n28324), .B(n28325), .Z(n28323) );
  NANDN U37097 ( .A(n28326), .B(n28327), .Z(n28325) );
  NANDN U37098 ( .A(n28327), .B(n28326), .Z(n28322) );
  XOR U37099 ( .A(n28298), .B(n28328), .Z(n28290) );
  XNOR U37100 ( .A(n28295), .B(n28297), .Z(n28328) );
  AND U37101 ( .A(n28329), .B(n28330), .Z(n28297) );
  NANDN U37102 ( .A(n28331), .B(n28332), .Z(n28330) );
  OR U37103 ( .A(n28333), .B(n28334), .Z(n28332) );
  IV U37104 ( .A(n28335), .Z(n28334) );
  NANDN U37105 ( .A(n28335), .B(n28333), .Z(n28329) );
  AND U37106 ( .A(n28336), .B(n28337), .Z(n28295) );
  NAND U37107 ( .A(n28338), .B(n28339), .Z(n28337) );
  NANDN U37108 ( .A(n28340), .B(n28341), .Z(n28339) );
  NANDN U37109 ( .A(n28341), .B(n28340), .Z(n28336) );
  IV U37110 ( .A(n28342), .Z(n28341) );
  NAND U37111 ( .A(n28343), .B(n28344), .Z(n28298) );
  NANDN U37112 ( .A(n28345), .B(n28346), .Z(n28344) );
  NANDN U37113 ( .A(n28347), .B(n28348), .Z(n28346) );
  NANDN U37114 ( .A(n28348), .B(n28347), .Z(n28343) );
  IV U37115 ( .A(n28349), .Z(n28347) );
  XOR U37116 ( .A(n28324), .B(n28350), .Z(N62868) );
  XNOR U37117 ( .A(n28327), .B(n28326), .Z(n28350) );
  XNOR U37118 ( .A(n28338), .B(n28351), .Z(n28326) );
  XNOR U37119 ( .A(n28342), .B(n28340), .Z(n28351) );
  XOR U37120 ( .A(n28348), .B(n28352), .Z(n28340) );
  XNOR U37121 ( .A(n28345), .B(n28349), .Z(n28352) );
  AND U37122 ( .A(n28353), .B(n28354), .Z(n28349) );
  NAND U37123 ( .A(n28355), .B(n28356), .Z(n28354) );
  NAND U37124 ( .A(n28357), .B(n28358), .Z(n28353) );
  AND U37125 ( .A(n28359), .B(n28360), .Z(n28345) );
  NAND U37126 ( .A(n28361), .B(n28362), .Z(n28360) );
  NAND U37127 ( .A(n28363), .B(n28364), .Z(n28359) );
  NANDN U37128 ( .A(n28365), .B(n28366), .Z(n28348) );
  ANDN U37129 ( .B(n28367), .A(n28368), .Z(n28342) );
  XNOR U37130 ( .A(n28333), .B(n28369), .Z(n28338) );
  XNOR U37131 ( .A(n28331), .B(n28335), .Z(n28369) );
  AND U37132 ( .A(n28370), .B(n28371), .Z(n28335) );
  NAND U37133 ( .A(n28372), .B(n28373), .Z(n28371) );
  NAND U37134 ( .A(n28374), .B(n28375), .Z(n28370) );
  AND U37135 ( .A(n28376), .B(n28377), .Z(n28331) );
  NAND U37136 ( .A(n28378), .B(n28379), .Z(n28377) );
  NAND U37137 ( .A(n28380), .B(n28381), .Z(n28376) );
  AND U37138 ( .A(n28382), .B(n28383), .Z(n28333) );
  NAND U37139 ( .A(n28384), .B(n28385), .Z(n28327) );
  XNOR U37140 ( .A(n28310), .B(n28386), .Z(n28324) );
  XNOR U37141 ( .A(n28314), .B(n28312), .Z(n28386) );
  XOR U37142 ( .A(n28320), .B(n28387), .Z(n28312) );
  XNOR U37143 ( .A(n28317), .B(n28321), .Z(n28387) );
  AND U37144 ( .A(n28388), .B(n28389), .Z(n28321) );
  NAND U37145 ( .A(n28390), .B(n28391), .Z(n28389) );
  NAND U37146 ( .A(n28392), .B(n28393), .Z(n28388) );
  AND U37147 ( .A(n28394), .B(n28395), .Z(n28317) );
  NAND U37148 ( .A(n28396), .B(n28397), .Z(n28395) );
  NAND U37149 ( .A(n28398), .B(n28399), .Z(n28394) );
  NANDN U37150 ( .A(n28400), .B(n28401), .Z(n28320) );
  ANDN U37151 ( .B(n28402), .A(n28403), .Z(n28314) );
  XNOR U37152 ( .A(n28305), .B(n28404), .Z(n28310) );
  XNOR U37153 ( .A(n28303), .B(n28307), .Z(n28404) );
  AND U37154 ( .A(n28405), .B(n28406), .Z(n28307) );
  NAND U37155 ( .A(n28407), .B(n28408), .Z(n28406) );
  NAND U37156 ( .A(n28409), .B(n28410), .Z(n28405) );
  AND U37157 ( .A(n28411), .B(n28412), .Z(n28303) );
  NAND U37158 ( .A(n28413), .B(n28414), .Z(n28412) );
  NAND U37159 ( .A(n28415), .B(n28416), .Z(n28411) );
  AND U37160 ( .A(n28417), .B(n28418), .Z(n28305) );
  XOR U37161 ( .A(n28385), .B(n28384), .Z(N62867) );
  XNOR U37162 ( .A(n28402), .B(n28403), .Z(n28384) );
  XNOR U37163 ( .A(n28417), .B(n28418), .Z(n28403) );
  XOR U37164 ( .A(n28414), .B(n28413), .Z(n28418) );
  XOR U37165 ( .A(y[4212]), .B(x[4212]), .Z(n28413) );
  XOR U37166 ( .A(n28416), .B(n28415), .Z(n28414) );
  XOR U37167 ( .A(y[4214]), .B(x[4214]), .Z(n28415) );
  XOR U37168 ( .A(y[4213]), .B(x[4213]), .Z(n28416) );
  XOR U37169 ( .A(n28408), .B(n28407), .Z(n28417) );
  XOR U37170 ( .A(n28410), .B(n28409), .Z(n28407) );
  XOR U37171 ( .A(y[4211]), .B(x[4211]), .Z(n28409) );
  XOR U37172 ( .A(y[4210]), .B(x[4210]), .Z(n28410) );
  XOR U37173 ( .A(y[4209]), .B(x[4209]), .Z(n28408) );
  XNOR U37174 ( .A(n28401), .B(n28400), .Z(n28402) );
  XNOR U37175 ( .A(n28397), .B(n28396), .Z(n28400) );
  XOR U37176 ( .A(n28399), .B(n28398), .Z(n28396) );
  XOR U37177 ( .A(y[4208]), .B(x[4208]), .Z(n28398) );
  XOR U37178 ( .A(y[4207]), .B(x[4207]), .Z(n28399) );
  XOR U37179 ( .A(y[4206]), .B(x[4206]), .Z(n28397) );
  XOR U37180 ( .A(n28391), .B(n28390), .Z(n28401) );
  XOR U37181 ( .A(n28393), .B(n28392), .Z(n28390) );
  XOR U37182 ( .A(y[4205]), .B(x[4205]), .Z(n28392) );
  XOR U37183 ( .A(y[4204]), .B(x[4204]), .Z(n28393) );
  XOR U37184 ( .A(y[4203]), .B(x[4203]), .Z(n28391) );
  XNOR U37185 ( .A(n28367), .B(n28368), .Z(n28385) );
  XNOR U37186 ( .A(n28382), .B(n28383), .Z(n28368) );
  XOR U37187 ( .A(n28379), .B(n28378), .Z(n28383) );
  XOR U37188 ( .A(y[4200]), .B(x[4200]), .Z(n28378) );
  XOR U37189 ( .A(n28381), .B(n28380), .Z(n28379) );
  XOR U37190 ( .A(y[4202]), .B(x[4202]), .Z(n28380) );
  XOR U37191 ( .A(y[4201]), .B(x[4201]), .Z(n28381) );
  XOR U37192 ( .A(n28373), .B(n28372), .Z(n28382) );
  XOR U37193 ( .A(n28375), .B(n28374), .Z(n28372) );
  XOR U37194 ( .A(y[4199]), .B(x[4199]), .Z(n28374) );
  XOR U37195 ( .A(y[4198]), .B(x[4198]), .Z(n28375) );
  XOR U37196 ( .A(y[4197]), .B(x[4197]), .Z(n28373) );
  XNOR U37197 ( .A(n28366), .B(n28365), .Z(n28367) );
  XNOR U37198 ( .A(n28362), .B(n28361), .Z(n28365) );
  XOR U37199 ( .A(n28364), .B(n28363), .Z(n28361) );
  XOR U37200 ( .A(y[4196]), .B(x[4196]), .Z(n28363) );
  XOR U37201 ( .A(y[4195]), .B(x[4195]), .Z(n28364) );
  XOR U37202 ( .A(y[4194]), .B(x[4194]), .Z(n28362) );
  XOR U37203 ( .A(n28356), .B(n28355), .Z(n28366) );
  XOR U37204 ( .A(n28358), .B(n28357), .Z(n28355) );
  XOR U37205 ( .A(y[4193]), .B(x[4193]), .Z(n28357) );
  XOR U37206 ( .A(y[4192]), .B(x[4192]), .Z(n28358) );
  XOR U37207 ( .A(y[4191]), .B(x[4191]), .Z(n28356) );
  NAND U37208 ( .A(n28419), .B(n28420), .Z(N62858) );
  NAND U37209 ( .A(n28421), .B(n28422), .Z(n28420) );
  NANDN U37210 ( .A(n28423), .B(n28424), .Z(n28422) );
  NANDN U37211 ( .A(n28424), .B(n28423), .Z(n28419) );
  XOR U37212 ( .A(n28423), .B(n28425), .Z(N62857) );
  XNOR U37213 ( .A(n28421), .B(n28424), .Z(n28425) );
  NAND U37214 ( .A(n28426), .B(n28427), .Z(n28424) );
  NAND U37215 ( .A(n28428), .B(n28429), .Z(n28427) );
  NANDN U37216 ( .A(n28430), .B(n28431), .Z(n28429) );
  NANDN U37217 ( .A(n28431), .B(n28430), .Z(n28426) );
  AND U37218 ( .A(n28432), .B(n28433), .Z(n28421) );
  NAND U37219 ( .A(n28434), .B(n28435), .Z(n28433) );
  NANDN U37220 ( .A(n28436), .B(n28437), .Z(n28435) );
  NANDN U37221 ( .A(n28437), .B(n28436), .Z(n28432) );
  IV U37222 ( .A(n28438), .Z(n28437) );
  AND U37223 ( .A(n28439), .B(n28440), .Z(n28423) );
  NAND U37224 ( .A(n28441), .B(n28442), .Z(n28440) );
  NANDN U37225 ( .A(n28443), .B(n28444), .Z(n28442) );
  NANDN U37226 ( .A(n28444), .B(n28443), .Z(n28439) );
  XOR U37227 ( .A(n28436), .B(n28445), .Z(N62856) );
  XNOR U37228 ( .A(n28434), .B(n28438), .Z(n28445) );
  XOR U37229 ( .A(n28431), .B(n28446), .Z(n28438) );
  XNOR U37230 ( .A(n28428), .B(n28430), .Z(n28446) );
  AND U37231 ( .A(n28447), .B(n28448), .Z(n28430) );
  NANDN U37232 ( .A(n28449), .B(n28450), .Z(n28448) );
  OR U37233 ( .A(n28451), .B(n28452), .Z(n28450) );
  IV U37234 ( .A(n28453), .Z(n28452) );
  NANDN U37235 ( .A(n28453), .B(n28451), .Z(n28447) );
  AND U37236 ( .A(n28454), .B(n28455), .Z(n28428) );
  NAND U37237 ( .A(n28456), .B(n28457), .Z(n28455) );
  NANDN U37238 ( .A(n28458), .B(n28459), .Z(n28457) );
  NANDN U37239 ( .A(n28459), .B(n28458), .Z(n28454) );
  IV U37240 ( .A(n28460), .Z(n28459) );
  NAND U37241 ( .A(n28461), .B(n28462), .Z(n28431) );
  NANDN U37242 ( .A(n28463), .B(n28464), .Z(n28462) );
  NANDN U37243 ( .A(n28465), .B(n28466), .Z(n28464) );
  NANDN U37244 ( .A(n28466), .B(n28465), .Z(n28461) );
  IV U37245 ( .A(n28467), .Z(n28465) );
  AND U37246 ( .A(n28468), .B(n28469), .Z(n28434) );
  NAND U37247 ( .A(n28470), .B(n28471), .Z(n28469) );
  NANDN U37248 ( .A(n28472), .B(n28473), .Z(n28471) );
  NANDN U37249 ( .A(n28473), .B(n28472), .Z(n28468) );
  XOR U37250 ( .A(n28444), .B(n28474), .Z(n28436) );
  XNOR U37251 ( .A(n28441), .B(n28443), .Z(n28474) );
  AND U37252 ( .A(n28475), .B(n28476), .Z(n28443) );
  NANDN U37253 ( .A(n28477), .B(n28478), .Z(n28476) );
  OR U37254 ( .A(n28479), .B(n28480), .Z(n28478) );
  IV U37255 ( .A(n28481), .Z(n28480) );
  NANDN U37256 ( .A(n28481), .B(n28479), .Z(n28475) );
  AND U37257 ( .A(n28482), .B(n28483), .Z(n28441) );
  NAND U37258 ( .A(n28484), .B(n28485), .Z(n28483) );
  NANDN U37259 ( .A(n28486), .B(n28487), .Z(n28485) );
  NANDN U37260 ( .A(n28487), .B(n28486), .Z(n28482) );
  IV U37261 ( .A(n28488), .Z(n28487) );
  NAND U37262 ( .A(n28489), .B(n28490), .Z(n28444) );
  NANDN U37263 ( .A(n28491), .B(n28492), .Z(n28490) );
  NANDN U37264 ( .A(n28493), .B(n28494), .Z(n28492) );
  NANDN U37265 ( .A(n28494), .B(n28493), .Z(n28489) );
  IV U37266 ( .A(n28495), .Z(n28493) );
  XOR U37267 ( .A(n28470), .B(n28496), .Z(N62855) );
  XNOR U37268 ( .A(n28473), .B(n28472), .Z(n28496) );
  XNOR U37269 ( .A(n28484), .B(n28497), .Z(n28472) );
  XNOR U37270 ( .A(n28488), .B(n28486), .Z(n28497) );
  XOR U37271 ( .A(n28494), .B(n28498), .Z(n28486) );
  XNOR U37272 ( .A(n28491), .B(n28495), .Z(n28498) );
  AND U37273 ( .A(n28499), .B(n28500), .Z(n28495) );
  NAND U37274 ( .A(n28501), .B(n28502), .Z(n28500) );
  NAND U37275 ( .A(n28503), .B(n28504), .Z(n28499) );
  AND U37276 ( .A(n28505), .B(n28506), .Z(n28491) );
  NAND U37277 ( .A(n28507), .B(n28508), .Z(n28506) );
  NAND U37278 ( .A(n28509), .B(n28510), .Z(n28505) );
  NANDN U37279 ( .A(n28511), .B(n28512), .Z(n28494) );
  ANDN U37280 ( .B(n28513), .A(n28514), .Z(n28488) );
  XNOR U37281 ( .A(n28479), .B(n28515), .Z(n28484) );
  XNOR U37282 ( .A(n28477), .B(n28481), .Z(n28515) );
  AND U37283 ( .A(n28516), .B(n28517), .Z(n28481) );
  NAND U37284 ( .A(n28518), .B(n28519), .Z(n28517) );
  NAND U37285 ( .A(n28520), .B(n28521), .Z(n28516) );
  AND U37286 ( .A(n28522), .B(n28523), .Z(n28477) );
  NAND U37287 ( .A(n28524), .B(n28525), .Z(n28523) );
  NAND U37288 ( .A(n28526), .B(n28527), .Z(n28522) );
  AND U37289 ( .A(n28528), .B(n28529), .Z(n28479) );
  NAND U37290 ( .A(n28530), .B(n28531), .Z(n28473) );
  XNOR U37291 ( .A(n28456), .B(n28532), .Z(n28470) );
  XNOR U37292 ( .A(n28460), .B(n28458), .Z(n28532) );
  XOR U37293 ( .A(n28466), .B(n28533), .Z(n28458) );
  XNOR U37294 ( .A(n28463), .B(n28467), .Z(n28533) );
  AND U37295 ( .A(n28534), .B(n28535), .Z(n28467) );
  NAND U37296 ( .A(n28536), .B(n28537), .Z(n28535) );
  NAND U37297 ( .A(n28538), .B(n28539), .Z(n28534) );
  AND U37298 ( .A(n28540), .B(n28541), .Z(n28463) );
  NAND U37299 ( .A(n28542), .B(n28543), .Z(n28541) );
  NAND U37300 ( .A(n28544), .B(n28545), .Z(n28540) );
  NANDN U37301 ( .A(n28546), .B(n28547), .Z(n28466) );
  ANDN U37302 ( .B(n28548), .A(n28549), .Z(n28460) );
  XNOR U37303 ( .A(n28451), .B(n28550), .Z(n28456) );
  XNOR U37304 ( .A(n28449), .B(n28453), .Z(n28550) );
  AND U37305 ( .A(n28551), .B(n28552), .Z(n28453) );
  NAND U37306 ( .A(n28553), .B(n28554), .Z(n28552) );
  NAND U37307 ( .A(n28555), .B(n28556), .Z(n28551) );
  AND U37308 ( .A(n28557), .B(n28558), .Z(n28449) );
  NAND U37309 ( .A(n28559), .B(n28560), .Z(n28558) );
  NAND U37310 ( .A(n28561), .B(n28562), .Z(n28557) );
  AND U37311 ( .A(n28563), .B(n28564), .Z(n28451) );
  XOR U37312 ( .A(n28531), .B(n28530), .Z(N62854) );
  XNOR U37313 ( .A(n28548), .B(n28549), .Z(n28530) );
  XNOR U37314 ( .A(n28563), .B(n28564), .Z(n28549) );
  XOR U37315 ( .A(n28560), .B(n28559), .Z(n28564) );
  XOR U37316 ( .A(y[4188]), .B(x[4188]), .Z(n28559) );
  XOR U37317 ( .A(n28562), .B(n28561), .Z(n28560) );
  XOR U37318 ( .A(y[4190]), .B(x[4190]), .Z(n28561) );
  XOR U37319 ( .A(y[4189]), .B(x[4189]), .Z(n28562) );
  XOR U37320 ( .A(n28554), .B(n28553), .Z(n28563) );
  XOR U37321 ( .A(n28556), .B(n28555), .Z(n28553) );
  XOR U37322 ( .A(y[4187]), .B(x[4187]), .Z(n28555) );
  XOR U37323 ( .A(y[4186]), .B(x[4186]), .Z(n28556) );
  XOR U37324 ( .A(y[4185]), .B(x[4185]), .Z(n28554) );
  XNOR U37325 ( .A(n28547), .B(n28546), .Z(n28548) );
  XNOR U37326 ( .A(n28543), .B(n28542), .Z(n28546) );
  XOR U37327 ( .A(n28545), .B(n28544), .Z(n28542) );
  XOR U37328 ( .A(y[4184]), .B(x[4184]), .Z(n28544) );
  XOR U37329 ( .A(y[4183]), .B(x[4183]), .Z(n28545) );
  XOR U37330 ( .A(y[4182]), .B(x[4182]), .Z(n28543) );
  XOR U37331 ( .A(n28537), .B(n28536), .Z(n28547) );
  XOR U37332 ( .A(n28539), .B(n28538), .Z(n28536) );
  XOR U37333 ( .A(y[4181]), .B(x[4181]), .Z(n28538) );
  XOR U37334 ( .A(y[4180]), .B(x[4180]), .Z(n28539) );
  XOR U37335 ( .A(y[4179]), .B(x[4179]), .Z(n28537) );
  XNOR U37336 ( .A(n28513), .B(n28514), .Z(n28531) );
  XNOR U37337 ( .A(n28528), .B(n28529), .Z(n28514) );
  XOR U37338 ( .A(n28525), .B(n28524), .Z(n28529) );
  XOR U37339 ( .A(y[4176]), .B(x[4176]), .Z(n28524) );
  XOR U37340 ( .A(n28527), .B(n28526), .Z(n28525) );
  XOR U37341 ( .A(y[4178]), .B(x[4178]), .Z(n28526) );
  XOR U37342 ( .A(y[4177]), .B(x[4177]), .Z(n28527) );
  XOR U37343 ( .A(n28519), .B(n28518), .Z(n28528) );
  XOR U37344 ( .A(n28521), .B(n28520), .Z(n28518) );
  XOR U37345 ( .A(y[4175]), .B(x[4175]), .Z(n28520) );
  XOR U37346 ( .A(y[4174]), .B(x[4174]), .Z(n28521) );
  XOR U37347 ( .A(y[4173]), .B(x[4173]), .Z(n28519) );
  XNOR U37348 ( .A(n28512), .B(n28511), .Z(n28513) );
  XNOR U37349 ( .A(n28508), .B(n28507), .Z(n28511) );
  XOR U37350 ( .A(n28510), .B(n28509), .Z(n28507) );
  XOR U37351 ( .A(y[4172]), .B(x[4172]), .Z(n28509) );
  XOR U37352 ( .A(y[4171]), .B(x[4171]), .Z(n28510) );
  XOR U37353 ( .A(y[4170]), .B(x[4170]), .Z(n28508) );
  XOR U37354 ( .A(n28502), .B(n28501), .Z(n28512) );
  XOR U37355 ( .A(n28504), .B(n28503), .Z(n28501) );
  XOR U37356 ( .A(y[4169]), .B(x[4169]), .Z(n28503) );
  XOR U37357 ( .A(y[4168]), .B(x[4168]), .Z(n28504) );
  XOR U37358 ( .A(y[4167]), .B(x[4167]), .Z(n28502) );
  NAND U37359 ( .A(n28565), .B(n28566), .Z(N62845) );
  NAND U37360 ( .A(n28567), .B(n28568), .Z(n28566) );
  NANDN U37361 ( .A(n28569), .B(n28570), .Z(n28568) );
  NANDN U37362 ( .A(n28570), .B(n28569), .Z(n28565) );
  XOR U37363 ( .A(n28569), .B(n28571), .Z(N62844) );
  XNOR U37364 ( .A(n28567), .B(n28570), .Z(n28571) );
  NAND U37365 ( .A(n28572), .B(n28573), .Z(n28570) );
  NAND U37366 ( .A(n28574), .B(n28575), .Z(n28573) );
  NANDN U37367 ( .A(n28576), .B(n28577), .Z(n28575) );
  NANDN U37368 ( .A(n28577), .B(n28576), .Z(n28572) );
  AND U37369 ( .A(n28578), .B(n28579), .Z(n28567) );
  NAND U37370 ( .A(n28580), .B(n28581), .Z(n28579) );
  NANDN U37371 ( .A(n28582), .B(n28583), .Z(n28581) );
  NANDN U37372 ( .A(n28583), .B(n28582), .Z(n28578) );
  IV U37373 ( .A(n28584), .Z(n28583) );
  AND U37374 ( .A(n28585), .B(n28586), .Z(n28569) );
  NAND U37375 ( .A(n28587), .B(n28588), .Z(n28586) );
  NANDN U37376 ( .A(n28589), .B(n28590), .Z(n28588) );
  NANDN U37377 ( .A(n28590), .B(n28589), .Z(n28585) );
  XOR U37378 ( .A(n28582), .B(n28591), .Z(N62843) );
  XNOR U37379 ( .A(n28580), .B(n28584), .Z(n28591) );
  XOR U37380 ( .A(n28577), .B(n28592), .Z(n28584) );
  XNOR U37381 ( .A(n28574), .B(n28576), .Z(n28592) );
  AND U37382 ( .A(n28593), .B(n28594), .Z(n28576) );
  NANDN U37383 ( .A(n28595), .B(n28596), .Z(n28594) );
  OR U37384 ( .A(n28597), .B(n28598), .Z(n28596) );
  IV U37385 ( .A(n28599), .Z(n28598) );
  NANDN U37386 ( .A(n28599), .B(n28597), .Z(n28593) );
  AND U37387 ( .A(n28600), .B(n28601), .Z(n28574) );
  NAND U37388 ( .A(n28602), .B(n28603), .Z(n28601) );
  NANDN U37389 ( .A(n28604), .B(n28605), .Z(n28603) );
  NANDN U37390 ( .A(n28605), .B(n28604), .Z(n28600) );
  IV U37391 ( .A(n28606), .Z(n28605) );
  NAND U37392 ( .A(n28607), .B(n28608), .Z(n28577) );
  NANDN U37393 ( .A(n28609), .B(n28610), .Z(n28608) );
  NANDN U37394 ( .A(n28611), .B(n28612), .Z(n28610) );
  NANDN U37395 ( .A(n28612), .B(n28611), .Z(n28607) );
  IV U37396 ( .A(n28613), .Z(n28611) );
  AND U37397 ( .A(n28614), .B(n28615), .Z(n28580) );
  NAND U37398 ( .A(n28616), .B(n28617), .Z(n28615) );
  NANDN U37399 ( .A(n28618), .B(n28619), .Z(n28617) );
  NANDN U37400 ( .A(n28619), .B(n28618), .Z(n28614) );
  XOR U37401 ( .A(n28590), .B(n28620), .Z(n28582) );
  XNOR U37402 ( .A(n28587), .B(n28589), .Z(n28620) );
  AND U37403 ( .A(n28621), .B(n28622), .Z(n28589) );
  NANDN U37404 ( .A(n28623), .B(n28624), .Z(n28622) );
  OR U37405 ( .A(n28625), .B(n28626), .Z(n28624) );
  IV U37406 ( .A(n28627), .Z(n28626) );
  NANDN U37407 ( .A(n28627), .B(n28625), .Z(n28621) );
  AND U37408 ( .A(n28628), .B(n28629), .Z(n28587) );
  NAND U37409 ( .A(n28630), .B(n28631), .Z(n28629) );
  NANDN U37410 ( .A(n28632), .B(n28633), .Z(n28631) );
  NANDN U37411 ( .A(n28633), .B(n28632), .Z(n28628) );
  IV U37412 ( .A(n28634), .Z(n28633) );
  NAND U37413 ( .A(n28635), .B(n28636), .Z(n28590) );
  NANDN U37414 ( .A(n28637), .B(n28638), .Z(n28636) );
  NANDN U37415 ( .A(n28639), .B(n28640), .Z(n28638) );
  NANDN U37416 ( .A(n28640), .B(n28639), .Z(n28635) );
  IV U37417 ( .A(n28641), .Z(n28639) );
  XOR U37418 ( .A(n28616), .B(n28642), .Z(N62842) );
  XNOR U37419 ( .A(n28619), .B(n28618), .Z(n28642) );
  XNOR U37420 ( .A(n28630), .B(n28643), .Z(n28618) );
  XNOR U37421 ( .A(n28634), .B(n28632), .Z(n28643) );
  XOR U37422 ( .A(n28640), .B(n28644), .Z(n28632) );
  XNOR U37423 ( .A(n28637), .B(n28641), .Z(n28644) );
  AND U37424 ( .A(n28645), .B(n28646), .Z(n28641) );
  NAND U37425 ( .A(n28647), .B(n28648), .Z(n28646) );
  NAND U37426 ( .A(n28649), .B(n28650), .Z(n28645) );
  AND U37427 ( .A(n28651), .B(n28652), .Z(n28637) );
  NAND U37428 ( .A(n28653), .B(n28654), .Z(n28652) );
  NAND U37429 ( .A(n28655), .B(n28656), .Z(n28651) );
  NANDN U37430 ( .A(n28657), .B(n28658), .Z(n28640) );
  ANDN U37431 ( .B(n28659), .A(n28660), .Z(n28634) );
  XNOR U37432 ( .A(n28625), .B(n28661), .Z(n28630) );
  XNOR U37433 ( .A(n28623), .B(n28627), .Z(n28661) );
  AND U37434 ( .A(n28662), .B(n28663), .Z(n28627) );
  NAND U37435 ( .A(n28664), .B(n28665), .Z(n28663) );
  NAND U37436 ( .A(n28666), .B(n28667), .Z(n28662) );
  AND U37437 ( .A(n28668), .B(n28669), .Z(n28623) );
  NAND U37438 ( .A(n28670), .B(n28671), .Z(n28669) );
  NAND U37439 ( .A(n28672), .B(n28673), .Z(n28668) );
  AND U37440 ( .A(n28674), .B(n28675), .Z(n28625) );
  NAND U37441 ( .A(n28676), .B(n28677), .Z(n28619) );
  XNOR U37442 ( .A(n28602), .B(n28678), .Z(n28616) );
  XNOR U37443 ( .A(n28606), .B(n28604), .Z(n28678) );
  XOR U37444 ( .A(n28612), .B(n28679), .Z(n28604) );
  XNOR U37445 ( .A(n28609), .B(n28613), .Z(n28679) );
  AND U37446 ( .A(n28680), .B(n28681), .Z(n28613) );
  NAND U37447 ( .A(n28682), .B(n28683), .Z(n28681) );
  NAND U37448 ( .A(n28684), .B(n28685), .Z(n28680) );
  AND U37449 ( .A(n28686), .B(n28687), .Z(n28609) );
  NAND U37450 ( .A(n28688), .B(n28689), .Z(n28687) );
  NAND U37451 ( .A(n28690), .B(n28691), .Z(n28686) );
  NANDN U37452 ( .A(n28692), .B(n28693), .Z(n28612) );
  ANDN U37453 ( .B(n28694), .A(n28695), .Z(n28606) );
  XNOR U37454 ( .A(n28597), .B(n28696), .Z(n28602) );
  XNOR U37455 ( .A(n28595), .B(n28599), .Z(n28696) );
  AND U37456 ( .A(n28697), .B(n28698), .Z(n28599) );
  NAND U37457 ( .A(n28699), .B(n28700), .Z(n28698) );
  NAND U37458 ( .A(n28701), .B(n28702), .Z(n28697) );
  AND U37459 ( .A(n28703), .B(n28704), .Z(n28595) );
  NAND U37460 ( .A(n28705), .B(n28706), .Z(n28704) );
  NAND U37461 ( .A(n28707), .B(n28708), .Z(n28703) );
  AND U37462 ( .A(n28709), .B(n28710), .Z(n28597) );
  XOR U37463 ( .A(n28677), .B(n28676), .Z(N62841) );
  XNOR U37464 ( .A(n28694), .B(n28695), .Z(n28676) );
  XNOR U37465 ( .A(n28709), .B(n28710), .Z(n28695) );
  XOR U37466 ( .A(n28706), .B(n28705), .Z(n28710) );
  XOR U37467 ( .A(y[4164]), .B(x[4164]), .Z(n28705) );
  XOR U37468 ( .A(n28708), .B(n28707), .Z(n28706) );
  XOR U37469 ( .A(y[4166]), .B(x[4166]), .Z(n28707) );
  XOR U37470 ( .A(y[4165]), .B(x[4165]), .Z(n28708) );
  XOR U37471 ( .A(n28700), .B(n28699), .Z(n28709) );
  XOR U37472 ( .A(n28702), .B(n28701), .Z(n28699) );
  XOR U37473 ( .A(y[4163]), .B(x[4163]), .Z(n28701) );
  XOR U37474 ( .A(y[4162]), .B(x[4162]), .Z(n28702) );
  XOR U37475 ( .A(y[4161]), .B(x[4161]), .Z(n28700) );
  XNOR U37476 ( .A(n28693), .B(n28692), .Z(n28694) );
  XNOR U37477 ( .A(n28689), .B(n28688), .Z(n28692) );
  XOR U37478 ( .A(n28691), .B(n28690), .Z(n28688) );
  XOR U37479 ( .A(y[4160]), .B(x[4160]), .Z(n28690) );
  XOR U37480 ( .A(y[4159]), .B(x[4159]), .Z(n28691) );
  XOR U37481 ( .A(y[4158]), .B(x[4158]), .Z(n28689) );
  XOR U37482 ( .A(n28683), .B(n28682), .Z(n28693) );
  XOR U37483 ( .A(n28685), .B(n28684), .Z(n28682) );
  XOR U37484 ( .A(y[4157]), .B(x[4157]), .Z(n28684) );
  XOR U37485 ( .A(y[4156]), .B(x[4156]), .Z(n28685) );
  XOR U37486 ( .A(y[4155]), .B(x[4155]), .Z(n28683) );
  XNOR U37487 ( .A(n28659), .B(n28660), .Z(n28677) );
  XNOR U37488 ( .A(n28674), .B(n28675), .Z(n28660) );
  XOR U37489 ( .A(n28671), .B(n28670), .Z(n28675) );
  XOR U37490 ( .A(y[4152]), .B(x[4152]), .Z(n28670) );
  XOR U37491 ( .A(n28673), .B(n28672), .Z(n28671) );
  XOR U37492 ( .A(y[4154]), .B(x[4154]), .Z(n28672) );
  XOR U37493 ( .A(y[4153]), .B(x[4153]), .Z(n28673) );
  XOR U37494 ( .A(n28665), .B(n28664), .Z(n28674) );
  XOR U37495 ( .A(n28667), .B(n28666), .Z(n28664) );
  XOR U37496 ( .A(y[4151]), .B(x[4151]), .Z(n28666) );
  XOR U37497 ( .A(y[4150]), .B(x[4150]), .Z(n28667) );
  XOR U37498 ( .A(y[4149]), .B(x[4149]), .Z(n28665) );
  XNOR U37499 ( .A(n28658), .B(n28657), .Z(n28659) );
  XNOR U37500 ( .A(n28654), .B(n28653), .Z(n28657) );
  XOR U37501 ( .A(n28656), .B(n28655), .Z(n28653) );
  XOR U37502 ( .A(y[4148]), .B(x[4148]), .Z(n28655) );
  XOR U37503 ( .A(y[4147]), .B(x[4147]), .Z(n28656) );
  XOR U37504 ( .A(y[4146]), .B(x[4146]), .Z(n28654) );
  XOR U37505 ( .A(n28648), .B(n28647), .Z(n28658) );
  XOR U37506 ( .A(n28650), .B(n28649), .Z(n28647) );
  XOR U37507 ( .A(y[4145]), .B(x[4145]), .Z(n28649) );
  XOR U37508 ( .A(y[4144]), .B(x[4144]), .Z(n28650) );
  XOR U37509 ( .A(y[4143]), .B(x[4143]), .Z(n28648) );
  NAND U37510 ( .A(n28711), .B(n28712), .Z(N62832) );
  NAND U37511 ( .A(n28713), .B(n28714), .Z(n28712) );
  NANDN U37512 ( .A(n28715), .B(n28716), .Z(n28714) );
  NANDN U37513 ( .A(n28716), .B(n28715), .Z(n28711) );
  XOR U37514 ( .A(n28715), .B(n28717), .Z(N62831) );
  XNOR U37515 ( .A(n28713), .B(n28716), .Z(n28717) );
  NAND U37516 ( .A(n28718), .B(n28719), .Z(n28716) );
  NAND U37517 ( .A(n28720), .B(n28721), .Z(n28719) );
  NANDN U37518 ( .A(n28722), .B(n28723), .Z(n28721) );
  NANDN U37519 ( .A(n28723), .B(n28722), .Z(n28718) );
  AND U37520 ( .A(n28724), .B(n28725), .Z(n28713) );
  NAND U37521 ( .A(n28726), .B(n28727), .Z(n28725) );
  NANDN U37522 ( .A(n28728), .B(n28729), .Z(n28727) );
  NANDN U37523 ( .A(n28729), .B(n28728), .Z(n28724) );
  IV U37524 ( .A(n28730), .Z(n28729) );
  AND U37525 ( .A(n28731), .B(n28732), .Z(n28715) );
  NAND U37526 ( .A(n28733), .B(n28734), .Z(n28732) );
  NANDN U37527 ( .A(n28735), .B(n28736), .Z(n28734) );
  NANDN U37528 ( .A(n28736), .B(n28735), .Z(n28731) );
  XOR U37529 ( .A(n28728), .B(n28737), .Z(N62830) );
  XNOR U37530 ( .A(n28726), .B(n28730), .Z(n28737) );
  XOR U37531 ( .A(n28723), .B(n28738), .Z(n28730) );
  XNOR U37532 ( .A(n28720), .B(n28722), .Z(n28738) );
  AND U37533 ( .A(n28739), .B(n28740), .Z(n28722) );
  NANDN U37534 ( .A(n28741), .B(n28742), .Z(n28740) );
  OR U37535 ( .A(n28743), .B(n28744), .Z(n28742) );
  IV U37536 ( .A(n28745), .Z(n28744) );
  NANDN U37537 ( .A(n28745), .B(n28743), .Z(n28739) );
  AND U37538 ( .A(n28746), .B(n28747), .Z(n28720) );
  NAND U37539 ( .A(n28748), .B(n28749), .Z(n28747) );
  NANDN U37540 ( .A(n28750), .B(n28751), .Z(n28749) );
  NANDN U37541 ( .A(n28751), .B(n28750), .Z(n28746) );
  IV U37542 ( .A(n28752), .Z(n28751) );
  NAND U37543 ( .A(n28753), .B(n28754), .Z(n28723) );
  NANDN U37544 ( .A(n28755), .B(n28756), .Z(n28754) );
  NANDN U37545 ( .A(n28757), .B(n28758), .Z(n28756) );
  NANDN U37546 ( .A(n28758), .B(n28757), .Z(n28753) );
  IV U37547 ( .A(n28759), .Z(n28757) );
  AND U37548 ( .A(n28760), .B(n28761), .Z(n28726) );
  NAND U37549 ( .A(n28762), .B(n28763), .Z(n28761) );
  NANDN U37550 ( .A(n28764), .B(n28765), .Z(n28763) );
  NANDN U37551 ( .A(n28765), .B(n28764), .Z(n28760) );
  XOR U37552 ( .A(n28736), .B(n28766), .Z(n28728) );
  XNOR U37553 ( .A(n28733), .B(n28735), .Z(n28766) );
  AND U37554 ( .A(n28767), .B(n28768), .Z(n28735) );
  NANDN U37555 ( .A(n28769), .B(n28770), .Z(n28768) );
  OR U37556 ( .A(n28771), .B(n28772), .Z(n28770) );
  IV U37557 ( .A(n28773), .Z(n28772) );
  NANDN U37558 ( .A(n28773), .B(n28771), .Z(n28767) );
  AND U37559 ( .A(n28774), .B(n28775), .Z(n28733) );
  NAND U37560 ( .A(n28776), .B(n28777), .Z(n28775) );
  NANDN U37561 ( .A(n28778), .B(n28779), .Z(n28777) );
  NANDN U37562 ( .A(n28779), .B(n28778), .Z(n28774) );
  IV U37563 ( .A(n28780), .Z(n28779) );
  NAND U37564 ( .A(n28781), .B(n28782), .Z(n28736) );
  NANDN U37565 ( .A(n28783), .B(n28784), .Z(n28782) );
  NANDN U37566 ( .A(n28785), .B(n28786), .Z(n28784) );
  NANDN U37567 ( .A(n28786), .B(n28785), .Z(n28781) );
  IV U37568 ( .A(n28787), .Z(n28785) );
  XOR U37569 ( .A(n28762), .B(n28788), .Z(N62829) );
  XNOR U37570 ( .A(n28765), .B(n28764), .Z(n28788) );
  XNOR U37571 ( .A(n28776), .B(n28789), .Z(n28764) );
  XNOR U37572 ( .A(n28780), .B(n28778), .Z(n28789) );
  XOR U37573 ( .A(n28786), .B(n28790), .Z(n28778) );
  XNOR U37574 ( .A(n28783), .B(n28787), .Z(n28790) );
  AND U37575 ( .A(n28791), .B(n28792), .Z(n28787) );
  NAND U37576 ( .A(n28793), .B(n28794), .Z(n28792) );
  NAND U37577 ( .A(n28795), .B(n28796), .Z(n28791) );
  AND U37578 ( .A(n28797), .B(n28798), .Z(n28783) );
  NAND U37579 ( .A(n28799), .B(n28800), .Z(n28798) );
  NAND U37580 ( .A(n28801), .B(n28802), .Z(n28797) );
  NANDN U37581 ( .A(n28803), .B(n28804), .Z(n28786) );
  ANDN U37582 ( .B(n28805), .A(n28806), .Z(n28780) );
  XNOR U37583 ( .A(n28771), .B(n28807), .Z(n28776) );
  XNOR U37584 ( .A(n28769), .B(n28773), .Z(n28807) );
  AND U37585 ( .A(n28808), .B(n28809), .Z(n28773) );
  NAND U37586 ( .A(n28810), .B(n28811), .Z(n28809) );
  NAND U37587 ( .A(n28812), .B(n28813), .Z(n28808) );
  AND U37588 ( .A(n28814), .B(n28815), .Z(n28769) );
  NAND U37589 ( .A(n28816), .B(n28817), .Z(n28815) );
  NAND U37590 ( .A(n28818), .B(n28819), .Z(n28814) );
  AND U37591 ( .A(n28820), .B(n28821), .Z(n28771) );
  NAND U37592 ( .A(n28822), .B(n28823), .Z(n28765) );
  XNOR U37593 ( .A(n28748), .B(n28824), .Z(n28762) );
  XNOR U37594 ( .A(n28752), .B(n28750), .Z(n28824) );
  XOR U37595 ( .A(n28758), .B(n28825), .Z(n28750) );
  XNOR U37596 ( .A(n28755), .B(n28759), .Z(n28825) );
  AND U37597 ( .A(n28826), .B(n28827), .Z(n28759) );
  NAND U37598 ( .A(n28828), .B(n28829), .Z(n28827) );
  NAND U37599 ( .A(n28830), .B(n28831), .Z(n28826) );
  AND U37600 ( .A(n28832), .B(n28833), .Z(n28755) );
  NAND U37601 ( .A(n28834), .B(n28835), .Z(n28833) );
  NAND U37602 ( .A(n28836), .B(n28837), .Z(n28832) );
  NANDN U37603 ( .A(n28838), .B(n28839), .Z(n28758) );
  ANDN U37604 ( .B(n28840), .A(n28841), .Z(n28752) );
  XNOR U37605 ( .A(n28743), .B(n28842), .Z(n28748) );
  XNOR U37606 ( .A(n28741), .B(n28745), .Z(n28842) );
  AND U37607 ( .A(n28843), .B(n28844), .Z(n28745) );
  NAND U37608 ( .A(n28845), .B(n28846), .Z(n28844) );
  NAND U37609 ( .A(n28847), .B(n28848), .Z(n28843) );
  AND U37610 ( .A(n28849), .B(n28850), .Z(n28741) );
  NAND U37611 ( .A(n28851), .B(n28852), .Z(n28850) );
  NAND U37612 ( .A(n28853), .B(n28854), .Z(n28849) );
  AND U37613 ( .A(n28855), .B(n28856), .Z(n28743) );
  XOR U37614 ( .A(n28823), .B(n28822), .Z(N62828) );
  XNOR U37615 ( .A(n28840), .B(n28841), .Z(n28822) );
  XNOR U37616 ( .A(n28855), .B(n28856), .Z(n28841) );
  XOR U37617 ( .A(n28852), .B(n28851), .Z(n28856) );
  XOR U37618 ( .A(y[4140]), .B(x[4140]), .Z(n28851) );
  XOR U37619 ( .A(n28854), .B(n28853), .Z(n28852) );
  XOR U37620 ( .A(y[4142]), .B(x[4142]), .Z(n28853) );
  XOR U37621 ( .A(y[4141]), .B(x[4141]), .Z(n28854) );
  XOR U37622 ( .A(n28846), .B(n28845), .Z(n28855) );
  XOR U37623 ( .A(n28848), .B(n28847), .Z(n28845) );
  XOR U37624 ( .A(y[4139]), .B(x[4139]), .Z(n28847) );
  XOR U37625 ( .A(y[4138]), .B(x[4138]), .Z(n28848) );
  XOR U37626 ( .A(y[4137]), .B(x[4137]), .Z(n28846) );
  XNOR U37627 ( .A(n28839), .B(n28838), .Z(n28840) );
  XNOR U37628 ( .A(n28835), .B(n28834), .Z(n28838) );
  XOR U37629 ( .A(n28837), .B(n28836), .Z(n28834) );
  XOR U37630 ( .A(y[4136]), .B(x[4136]), .Z(n28836) );
  XOR U37631 ( .A(y[4135]), .B(x[4135]), .Z(n28837) );
  XOR U37632 ( .A(y[4134]), .B(x[4134]), .Z(n28835) );
  XOR U37633 ( .A(n28829), .B(n28828), .Z(n28839) );
  XOR U37634 ( .A(n28831), .B(n28830), .Z(n28828) );
  XOR U37635 ( .A(y[4133]), .B(x[4133]), .Z(n28830) );
  XOR U37636 ( .A(y[4132]), .B(x[4132]), .Z(n28831) );
  XOR U37637 ( .A(y[4131]), .B(x[4131]), .Z(n28829) );
  XNOR U37638 ( .A(n28805), .B(n28806), .Z(n28823) );
  XNOR U37639 ( .A(n28820), .B(n28821), .Z(n28806) );
  XOR U37640 ( .A(n28817), .B(n28816), .Z(n28821) );
  XOR U37641 ( .A(y[4128]), .B(x[4128]), .Z(n28816) );
  XOR U37642 ( .A(n28819), .B(n28818), .Z(n28817) );
  XOR U37643 ( .A(y[4130]), .B(x[4130]), .Z(n28818) );
  XOR U37644 ( .A(y[4129]), .B(x[4129]), .Z(n28819) );
  XOR U37645 ( .A(n28811), .B(n28810), .Z(n28820) );
  XOR U37646 ( .A(n28813), .B(n28812), .Z(n28810) );
  XOR U37647 ( .A(y[4127]), .B(x[4127]), .Z(n28812) );
  XOR U37648 ( .A(y[4126]), .B(x[4126]), .Z(n28813) );
  XOR U37649 ( .A(y[4125]), .B(x[4125]), .Z(n28811) );
  XNOR U37650 ( .A(n28804), .B(n28803), .Z(n28805) );
  XNOR U37651 ( .A(n28800), .B(n28799), .Z(n28803) );
  XOR U37652 ( .A(n28802), .B(n28801), .Z(n28799) );
  XOR U37653 ( .A(y[4124]), .B(x[4124]), .Z(n28801) );
  XOR U37654 ( .A(y[4123]), .B(x[4123]), .Z(n28802) );
  XOR U37655 ( .A(y[4122]), .B(x[4122]), .Z(n28800) );
  XOR U37656 ( .A(n28794), .B(n28793), .Z(n28804) );
  XOR U37657 ( .A(n28796), .B(n28795), .Z(n28793) );
  XOR U37658 ( .A(y[4121]), .B(x[4121]), .Z(n28795) );
  XOR U37659 ( .A(y[4120]), .B(x[4120]), .Z(n28796) );
  XOR U37660 ( .A(y[4119]), .B(x[4119]), .Z(n28794) );
  NAND U37661 ( .A(n28857), .B(n28858), .Z(N62819) );
  NAND U37662 ( .A(n28859), .B(n28860), .Z(n28858) );
  NANDN U37663 ( .A(n28861), .B(n28862), .Z(n28860) );
  NANDN U37664 ( .A(n28862), .B(n28861), .Z(n28857) );
  XOR U37665 ( .A(n28861), .B(n28863), .Z(N62818) );
  XNOR U37666 ( .A(n28859), .B(n28862), .Z(n28863) );
  NAND U37667 ( .A(n28864), .B(n28865), .Z(n28862) );
  NAND U37668 ( .A(n28866), .B(n28867), .Z(n28865) );
  NANDN U37669 ( .A(n28868), .B(n28869), .Z(n28867) );
  NANDN U37670 ( .A(n28869), .B(n28868), .Z(n28864) );
  AND U37671 ( .A(n28870), .B(n28871), .Z(n28859) );
  NAND U37672 ( .A(n28872), .B(n28873), .Z(n28871) );
  NANDN U37673 ( .A(n28874), .B(n28875), .Z(n28873) );
  NANDN U37674 ( .A(n28875), .B(n28874), .Z(n28870) );
  IV U37675 ( .A(n28876), .Z(n28875) );
  AND U37676 ( .A(n28877), .B(n28878), .Z(n28861) );
  NAND U37677 ( .A(n28879), .B(n28880), .Z(n28878) );
  NANDN U37678 ( .A(n28881), .B(n28882), .Z(n28880) );
  NANDN U37679 ( .A(n28882), .B(n28881), .Z(n28877) );
  XOR U37680 ( .A(n28874), .B(n28883), .Z(N62817) );
  XNOR U37681 ( .A(n28872), .B(n28876), .Z(n28883) );
  XOR U37682 ( .A(n28869), .B(n28884), .Z(n28876) );
  XNOR U37683 ( .A(n28866), .B(n28868), .Z(n28884) );
  AND U37684 ( .A(n28885), .B(n28886), .Z(n28868) );
  NANDN U37685 ( .A(n28887), .B(n28888), .Z(n28886) );
  OR U37686 ( .A(n28889), .B(n28890), .Z(n28888) );
  IV U37687 ( .A(n28891), .Z(n28890) );
  NANDN U37688 ( .A(n28891), .B(n28889), .Z(n28885) );
  AND U37689 ( .A(n28892), .B(n28893), .Z(n28866) );
  NAND U37690 ( .A(n28894), .B(n28895), .Z(n28893) );
  NANDN U37691 ( .A(n28896), .B(n28897), .Z(n28895) );
  NANDN U37692 ( .A(n28897), .B(n28896), .Z(n28892) );
  IV U37693 ( .A(n28898), .Z(n28897) );
  NAND U37694 ( .A(n28899), .B(n28900), .Z(n28869) );
  NANDN U37695 ( .A(n28901), .B(n28902), .Z(n28900) );
  NANDN U37696 ( .A(n28903), .B(n28904), .Z(n28902) );
  NANDN U37697 ( .A(n28904), .B(n28903), .Z(n28899) );
  IV U37698 ( .A(n28905), .Z(n28903) );
  AND U37699 ( .A(n28906), .B(n28907), .Z(n28872) );
  NAND U37700 ( .A(n28908), .B(n28909), .Z(n28907) );
  NANDN U37701 ( .A(n28910), .B(n28911), .Z(n28909) );
  NANDN U37702 ( .A(n28911), .B(n28910), .Z(n28906) );
  XOR U37703 ( .A(n28882), .B(n28912), .Z(n28874) );
  XNOR U37704 ( .A(n28879), .B(n28881), .Z(n28912) );
  AND U37705 ( .A(n28913), .B(n28914), .Z(n28881) );
  NANDN U37706 ( .A(n28915), .B(n28916), .Z(n28914) );
  OR U37707 ( .A(n28917), .B(n28918), .Z(n28916) );
  IV U37708 ( .A(n28919), .Z(n28918) );
  NANDN U37709 ( .A(n28919), .B(n28917), .Z(n28913) );
  AND U37710 ( .A(n28920), .B(n28921), .Z(n28879) );
  NAND U37711 ( .A(n28922), .B(n28923), .Z(n28921) );
  NANDN U37712 ( .A(n28924), .B(n28925), .Z(n28923) );
  NANDN U37713 ( .A(n28925), .B(n28924), .Z(n28920) );
  IV U37714 ( .A(n28926), .Z(n28925) );
  NAND U37715 ( .A(n28927), .B(n28928), .Z(n28882) );
  NANDN U37716 ( .A(n28929), .B(n28930), .Z(n28928) );
  NANDN U37717 ( .A(n28931), .B(n28932), .Z(n28930) );
  NANDN U37718 ( .A(n28932), .B(n28931), .Z(n28927) );
  IV U37719 ( .A(n28933), .Z(n28931) );
  XOR U37720 ( .A(n28908), .B(n28934), .Z(N62816) );
  XNOR U37721 ( .A(n28911), .B(n28910), .Z(n28934) );
  XNOR U37722 ( .A(n28922), .B(n28935), .Z(n28910) );
  XNOR U37723 ( .A(n28926), .B(n28924), .Z(n28935) );
  XOR U37724 ( .A(n28932), .B(n28936), .Z(n28924) );
  XNOR U37725 ( .A(n28929), .B(n28933), .Z(n28936) );
  AND U37726 ( .A(n28937), .B(n28938), .Z(n28933) );
  NAND U37727 ( .A(n28939), .B(n28940), .Z(n28938) );
  NAND U37728 ( .A(n28941), .B(n28942), .Z(n28937) );
  AND U37729 ( .A(n28943), .B(n28944), .Z(n28929) );
  NAND U37730 ( .A(n28945), .B(n28946), .Z(n28944) );
  NAND U37731 ( .A(n28947), .B(n28948), .Z(n28943) );
  NANDN U37732 ( .A(n28949), .B(n28950), .Z(n28932) );
  ANDN U37733 ( .B(n28951), .A(n28952), .Z(n28926) );
  XNOR U37734 ( .A(n28917), .B(n28953), .Z(n28922) );
  XNOR U37735 ( .A(n28915), .B(n28919), .Z(n28953) );
  AND U37736 ( .A(n28954), .B(n28955), .Z(n28919) );
  NAND U37737 ( .A(n28956), .B(n28957), .Z(n28955) );
  NAND U37738 ( .A(n28958), .B(n28959), .Z(n28954) );
  AND U37739 ( .A(n28960), .B(n28961), .Z(n28915) );
  NAND U37740 ( .A(n28962), .B(n28963), .Z(n28961) );
  NAND U37741 ( .A(n28964), .B(n28965), .Z(n28960) );
  AND U37742 ( .A(n28966), .B(n28967), .Z(n28917) );
  NAND U37743 ( .A(n28968), .B(n28969), .Z(n28911) );
  XNOR U37744 ( .A(n28894), .B(n28970), .Z(n28908) );
  XNOR U37745 ( .A(n28898), .B(n28896), .Z(n28970) );
  XOR U37746 ( .A(n28904), .B(n28971), .Z(n28896) );
  XNOR U37747 ( .A(n28901), .B(n28905), .Z(n28971) );
  AND U37748 ( .A(n28972), .B(n28973), .Z(n28905) );
  NAND U37749 ( .A(n28974), .B(n28975), .Z(n28973) );
  NAND U37750 ( .A(n28976), .B(n28977), .Z(n28972) );
  AND U37751 ( .A(n28978), .B(n28979), .Z(n28901) );
  NAND U37752 ( .A(n28980), .B(n28981), .Z(n28979) );
  NAND U37753 ( .A(n28982), .B(n28983), .Z(n28978) );
  NANDN U37754 ( .A(n28984), .B(n28985), .Z(n28904) );
  ANDN U37755 ( .B(n28986), .A(n28987), .Z(n28898) );
  XNOR U37756 ( .A(n28889), .B(n28988), .Z(n28894) );
  XNOR U37757 ( .A(n28887), .B(n28891), .Z(n28988) );
  AND U37758 ( .A(n28989), .B(n28990), .Z(n28891) );
  NAND U37759 ( .A(n28991), .B(n28992), .Z(n28990) );
  NAND U37760 ( .A(n28993), .B(n28994), .Z(n28989) );
  AND U37761 ( .A(n28995), .B(n28996), .Z(n28887) );
  NAND U37762 ( .A(n28997), .B(n28998), .Z(n28996) );
  NAND U37763 ( .A(n28999), .B(n29000), .Z(n28995) );
  AND U37764 ( .A(n29001), .B(n29002), .Z(n28889) );
  XOR U37765 ( .A(n28969), .B(n28968), .Z(N62815) );
  XNOR U37766 ( .A(n28986), .B(n28987), .Z(n28968) );
  XNOR U37767 ( .A(n29001), .B(n29002), .Z(n28987) );
  XOR U37768 ( .A(n28998), .B(n28997), .Z(n29002) );
  XOR U37769 ( .A(y[4116]), .B(x[4116]), .Z(n28997) );
  XOR U37770 ( .A(n29000), .B(n28999), .Z(n28998) );
  XOR U37771 ( .A(y[4118]), .B(x[4118]), .Z(n28999) );
  XOR U37772 ( .A(y[4117]), .B(x[4117]), .Z(n29000) );
  XOR U37773 ( .A(n28992), .B(n28991), .Z(n29001) );
  XOR U37774 ( .A(n28994), .B(n28993), .Z(n28991) );
  XOR U37775 ( .A(y[4115]), .B(x[4115]), .Z(n28993) );
  XOR U37776 ( .A(y[4114]), .B(x[4114]), .Z(n28994) );
  XOR U37777 ( .A(y[4113]), .B(x[4113]), .Z(n28992) );
  XNOR U37778 ( .A(n28985), .B(n28984), .Z(n28986) );
  XNOR U37779 ( .A(n28981), .B(n28980), .Z(n28984) );
  XOR U37780 ( .A(n28983), .B(n28982), .Z(n28980) );
  XOR U37781 ( .A(y[4112]), .B(x[4112]), .Z(n28982) );
  XOR U37782 ( .A(y[4111]), .B(x[4111]), .Z(n28983) );
  XOR U37783 ( .A(y[4110]), .B(x[4110]), .Z(n28981) );
  XOR U37784 ( .A(n28975), .B(n28974), .Z(n28985) );
  XOR U37785 ( .A(n28977), .B(n28976), .Z(n28974) );
  XOR U37786 ( .A(y[4109]), .B(x[4109]), .Z(n28976) );
  XOR U37787 ( .A(y[4108]), .B(x[4108]), .Z(n28977) );
  XOR U37788 ( .A(y[4107]), .B(x[4107]), .Z(n28975) );
  XNOR U37789 ( .A(n28951), .B(n28952), .Z(n28969) );
  XNOR U37790 ( .A(n28966), .B(n28967), .Z(n28952) );
  XOR U37791 ( .A(n28963), .B(n28962), .Z(n28967) );
  XOR U37792 ( .A(y[4104]), .B(x[4104]), .Z(n28962) );
  XOR U37793 ( .A(n28965), .B(n28964), .Z(n28963) );
  XOR U37794 ( .A(y[4106]), .B(x[4106]), .Z(n28964) );
  XOR U37795 ( .A(y[4105]), .B(x[4105]), .Z(n28965) );
  XOR U37796 ( .A(n28957), .B(n28956), .Z(n28966) );
  XOR U37797 ( .A(n28959), .B(n28958), .Z(n28956) );
  XOR U37798 ( .A(y[4103]), .B(x[4103]), .Z(n28958) );
  XOR U37799 ( .A(y[4102]), .B(x[4102]), .Z(n28959) );
  XOR U37800 ( .A(y[4101]), .B(x[4101]), .Z(n28957) );
  XNOR U37801 ( .A(n28950), .B(n28949), .Z(n28951) );
  XNOR U37802 ( .A(n28946), .B(n28945), .Z(n28949) );
  XOR U37803 ( .A(n28948), .B(n28947), .Z(n28945) );
  XOR U37804 ( .A(y[4100]), .B(x[4100]), .Z(n28947) );
  XOR U37805 ( .A(y[4099]), .B(x[4099]), .Z(n28948) );
  XOR U37806 ( .A(y[4098]), .B(x[4098]), .Z(n28946) );
  XOR U37807 ( .A(n28940), .B(n28939), .Z(n28950) );
  XOR U37808 ( .A(n28942), .B(n28941), .Z(n28939) );
  XOR U37809 ( .A(y[4097]), .B(x[4097]), .Z(n28941) );
  XOR U37810 ( .A(y[4096]), .B(x[4096]), .Z(n28942) );
  XOR U37811 ( .A(y[4095]), .B(x[4095]), .Z(n28940) );
  NAND U37812 ( .A(n29003), .B(n29004), .Z(N62806) );
  NAND U37813 ( .A(n29005), .B(n29006), .Z(n29004) );
  NANDN U37814 ( .A(n29007), .B(n29008), .Z(n29006) );
  NANDN U37815 ( .A(n29008), .B(n29007), .Z(n29003) );
  XOR U37816 ( .A(n29007), .B(n29009), .Z(N62805) );
  XNOR U37817 ( .A(n29005), .B(n29008), .Z(n29009) );
  NAND U37818 ( .A(n29010), .B(n29011), .Z(n29008) );
  NAND U37819 ( .A(n29012), .B(n29013), .Z(n29011) );
  NANDN U37820 ( .A(n29014), .B(n29015), .Z(n29013) );
  NANDN U37821 ( .A(n29015), .B(n29014), .Z(n29010) );
  AND U37822 ( .A(n29016), .B(n29017), .Z(n29005) );
  NAND U37823 ( .A(n29018), .B(n29019), .Z(n29017) );
  NANDN U37824 ( .A(n29020), .B(n29021), .Z(n29019) );
  NANDN U37825 ( .A(n29021), .B(n29020), .Z(n29016) );
  IV U37826 ( .A(n29022), .Z(n29021) );
  AND U37827 ( .A(n29023), .B(n29024), .Z(n29007) );
  NAND U37828 ( .A(n29025), .B(n29026), .Z(n29024) );
  NANDN U37829 ( .A(n29027), .B(n29028), .Z(n29026) );
  NANDN U37830 ( .A(n29028), .B(n29027), .Z(n29023) );
  XOR U37831 ( .A(n29020), .B(n29029), .Z(N62804) );
  XNOR U37832 ( .A(n29018), .B(n29022), .Z(n29029) );
  XOR U37833 ( .A(n29015), .B(n29030), .Z(n29022) );
  XNOR U37834 ( .A(n29012), .B(n29014), .Z(n29030) );
  AND U37835 ( .A(n29031), .B(n29032), .Z(n29014) );
  NANDN U37836 ( .A(n29033), .B(n29034), .Z(n29032) );
  OR U37837 ( .A(n29035), .B(n29036), .Z(n29034) );
  IV U37838 ( .A(n29037), .Z(n29036) );
  NANDN U37839 ( .A(n29037), .B(n29035), .Z(n29031) );
  AND U37840 ( .A(n29038), .B(n29039), .Z(n29012) );
  NAND U37841 ( .A(n29040), .B(n29041), .Z(n29039) );
  NANDN U37842 ( .A(n29042), .B(n29043), .Z(n29041) );
  NANDN U37843 ( .A(n29043), .B(n29042), .Z(n29038) );
  IV U37844 ( .A(n29044), .Z(n29043) );
  NAND U37845 ( .A(n29045), .B(n29046), .Z(n29015) );
  NANDN U37846 ( .A(n29047), .B(n29048), .Z(n29046) );
  NANDN U37847 ( .A(n29049), .B(n29050), .Z(n29048) );
  NANDN U37848 ( .A(n29050), .B(n29049), .Z(n29045) );
  IV U37849 ( .A(n29051), .Z(n29049) );
  AND U37850 ( .A(n29052), .B(n29053), .Z(n29018) );
  NAND U37851 ( .A(n29054), .B(n29055), .Z(n29053) );
  NANDN U37852 ( .A(n29056), .B(n29057), .Z(n29055) );
  NANDN U37853 ( .A(n29057), .B(n29056), .Z(n29052) );
  XOR U37854 ( .A(n29028), .B(n29058), .Z(n29020) );
  XNOR U37855 ( .A(n29025), .B(n29027), .Z(n29058) );
  AND U37856 ( .A(n29059), .B(n29060), .Z(n29027) );
  NANDN U37857 ( .A(n29061), .B(n29062), .Z(n29060) );
  OR U37858 ( .A(n29063), .B(n29064), .Z(n29062) );
  IV U37859 ( .A(n29065), .Z(n29064) );
  NANDN U37860 ( .A(n29065), .B(n29063), .Z(n29059) );
  AND U37861 ( .A(n29066), .B(n29067), .Z(n29025) );
  NAND U37862 ( .A(n29068), .B(n29069), .Z(n29067) );
  NANDN U37863 ( .A(n29070), .B(n29071), .Z(n29069) );
  NANDN U37864 ( .A(n29071), .B(n29070), .Z(n29066) );
  IV U37865 ( .A(n29072), .Z(n29071) );
  NAND U37866 ( .A(n29073), .B(n29074), .Z(n29028) );
  NANDN U37867 ( .A(n29075), .B(n29076), .Z(n29074) );
  NANDN U37868 ( .A(n29077), .B(n29078), .Z(n29076) );
  NANDN U37869 ( .A(n29078), .B(n29077), .Z(n29073) );
  IV U37870 ( .A(n29079), .Z(n29077) );
  XOR U37871 ( .A(n29054), .B(n29080), .Z(N62803) );
  XNOR U37872 ( .A(n29057), .B(n29056), .Z(n29080) );
  XNOR U37873 ( .A(n29068), .B(n29081), .Z(n29056) );
  XNOR U37874 ( .A(n29072), .B(n29070), .Z(n29081) );
  XOR U37875 ( .A(n29078), .B(n29082), .Z(n29070) );
  XNOR U37876 ( .A(n29075), .B(n29079), .Z(n29082) );
  AND U37877 ( .A(n29083), .B(n29084), .Z(n29079) );
  NAND U37878 ( .A(n29085), .B(n29086), .Z(n29084) );
  NAND U37879 ( .A(n29087), .B(n29088), .Z(n29083) );
  AND U37880 ( .A(n29089), .B(n29090), .Z(n29075) );
  NAND U37881 ( .A(n29091), .B(n29092), .Z(n29090) );
  NAND U37882 ( .A(n29093), .B(n29094), .Z(n29089) );
  NANDN U37883 ( .A(n29095), .B(n29096), .Z(n29078) );
  ANDN U37884 ( .B(n29097), .A(n29098), .Z(n29072) );
  XNOR U37885 ( .A(n29063), .B(n29099), .Z(n29068) );
  XNOR U37886 ( .A(n29061), .B(n29065), .Z(n29099) );
  AND U37887 ( .A(n29100), .B(n29101), .Z(n29065) );
  NAND U37888 ( .A(n29102), .B(n29103), .Z(n29101) );
  NAND U37889 ( .A(n29104), .B(n29105), .Z(n29100) );
  AND U37890 ( .A(n29106), .B(n29107), .Z(n29061) );
  NAND U37891 ( .A(n29108), .B(n29109), .Z(n29107) );
  NAND U37892 ( .A(n29110), .B(n29111), .Z(n29106) );
  AND U37893 ( .A(n29112), .B(n29113), .Z(n29063) );
  NAND U37894 ( .A(n29114), .B(n29115), .Z(n29057) );
  XNOR U37895 ( .A(n29040), .B(n29116), .Z(n29054) );
  XNOR U37896 ( .A(n29044), .B(n29042), .Z(n29116) );
  XOR U37897 ( .A(n29050), .B(n29117), .Z(n29042) );
  XNOR U37898 ( .A(n29047), .B(n29051), .Z(n29117) );
  AND U37899 ( .A(n29118), .B(n29119), .Z(n29051) );
  NAND U37900 ( .A(n29120), .B(n29121), .Z(n29119) );
  NAND U37901 ( .A(n29122), .B(n29123), .Z(n29118) );
  AND U37902 ( .A(n29124), .B(n29125), .Z(n29047) );
  NAND U37903 ( .A(n29126), .B(n29127), .Z(n29125) );
  NAND U37904 ( .A(n29128), .B(n29129), .Z(n29124) );
  NANDN U37905 ( .A(n29130), .B(n29131), .Z(n29050) );
  ANDN U37906 ( .B(n29132), .A(n29133), .Z(n29044) );
  XNOR U37907 ( .A(n29035), .B(n29134), .Z(n29040) );
  XNOR U37908 ( .A(n29033), .B(n29037), .Z(n29134) );
  AND U37909 ( .A(n29135), .B(n29136), .Z(n29037) );
  NAND U37910 ( .A(n29137), .B(n29138), .Z(n29136) );
  NAND U37911 ( .A(n29139), .B(n29140), .Z(n29135) );
  AND U37912 ( .A(n29141), .B(n29142), .Z(n29033) );
  NAND U37913 ( .A(n29143), .B(n29144), .Z(n29142) );
  NAND U37914 ( .A(n29145), .B(n29146), .Z(n29141) );
  AND U37915 ( .A(n29147), .B(n29148), .Z(n29035) );
  XOR U37916 ( .A(n29115), .B(n29114), .Z(N62802) );
  XNOR U37917 ( .A(n29132), .B(n29133), .Z(n29114) );
  XNOR U37918 ( .A(n29147), .B(n29148), .Z(n29133) );
  XOR U37919 ( .A(n29144), .B(n29143), .Z(n29148) );
  XOR U37920 ( .A(y[4092]), .B(x[4092]), .Z(n29143) );
  XOR U37921 ( .A(n29146), .B(n29145), .Z(n29144) );
  XOR U37922 ( .A(y[4094]), .B(x[4094]), .Z(n29145) );
  XOR U37923 ( .A(y[4093]), .B(x[4093]), .Z(n29146) );
  XOR U37924 ( .A(n29138), .B(n29137), .Z(n29147) );
  XOR U37925 ( .A(n29140), .B(n29139), .Z(n29137) );
  XOR U37926 ( .A(y[4091]), .B(x[4091]), .Z(n29139) );
  XOR U37927 ( .A(y[4090]), .B(x[4090]), .Z(n29140) );
  XOR U37928 ( .A(y[4089]), .B(x[4089]), .Z(n29138) );
  XNOR U37929 ( .A(n29131), .B(n29130), .Z(n29132) );
  XNOR U37930 ( .A(n29127), .B(n29126), .Z(n29130) );
  XOR U37931 ( .A(n29129), .B(n29128), .Z(n29126) );
  XOR U37932 ( .A(y[4088]), .B(x[4088]), .Z(n29128) );
  XOR U37933 ( .A(y[4087]), .B(x[4087]), .Z(n29129) );
  XOR U37934 ( .A(y[4086]), .B(x[4086]), .Z(n29127) );
  XOR U37935 ( .A(n29121), .B(n29120), .Z(n29131) );
  XOR U37936 ( .A(n29123), .B(n29122), .Z(n29120) );
  XOR U37937 ( .A(y[4085]), .B(x[4085]), .Z(n29122) );
  XOR U37938 ( .A(y[4084]), .B(x[4084]), .Z(n29123) );
  XOR U37939 ( .A(y[4083]), .B(x[4083]), .Z(n29121) );
  XNOR U37940 ( .A(n29097), .B(n29098), .Z(n29115) );
  XNOR U37941 ( .A(n29112), .B(n29113), .Z(n29098) );
  XOR U37942 ( .A(n29109), .B(n29108), .Z(n29113) );
  XOR U37943 ( .A(y[4080]), .B(x[4080]), .Z(n29108) );
  XOR U37944 ( .A(n29111), .B(n29110), .Z(n29109) );
  XOR U37945 ( .A(y[4082]), .B(x[4082]), .Z(n29110) );
  XOR U37946 ( .A(y[4081]), .B(x[4081]), .Z(n29111) );
  XOR U37947 ( .A(n29103), .B(n29102), .Z(n29112) );
  XOR U37948 ( .A(n29105), .B(n29104), .Z(n29102) );
  XOR U37949 ( .A(y[4079]), .B(x[4079]), .Z(n29104) );
  XOR U37950 ( .A(y[4078]), .B(x[4078]), .Z(n29105) );
  XOR U37951 ( .A(y[4077]), .B(x[4077]), .Z(n29103) );
  XNOR U37952 ( .A(n29096), .B(n29095), .Z(n29097) );
  XNOR U37953 ( .A(n29092), .B(n29091), .Z(n29095) );
  XOR U37954 ( .A(n29094), .B(n29093), .Z(n29091) );
  XOR U37955 ( .A(y[4076]), .B(x[4076]), .Z(n29093) );
  XOR U37956 ( .A(y[4075]), .B(x[4075]), .Z(n29094) );
  XOR U37957 ( .A(y[4074]), .B(x[4074]), .Z(n29092) );
  XOR U37958 ( .A(n29086), .B(n29085), .Z(n29096) );
  XOR U37959 ( .A(n29088), .B(n29087), .Z(n29085) );
  XOR U37960 ( .A(y[4073]), .B(x[4073]), .Z(n29087) );
  XOR U37961 ( .A(y[4072]), .B(x[4072]), .Z(n29088) );
  XOR U37962 ( .A(y[4071]), .B(x[4071]), .Z(n29086) );
  NAND U37963 ( .A(n29149), .B(n29150), .Z(N62793) );
  NAND U37964 ( .A(n29151), .B(n29152), .Z(n29150) );
  NANDN U37965 ( .A(n29153), .B(n29154), .Z(n29152) );
  NANDN U37966 ( .A(n29154), .B(n29153), .Z(n29149) );
  XOR U37967 ( .A(n29153), .B(n29155), .Z(N62792) );
  XNOR U37968 ( .A(n29151), .B(n29154), .Z(n29155) );
  NAND U37969 ( .A(n29156), .B(n29157), .Z(n29154) );
  NAND U37970 ( .A(n29158), .B(n29159), .Z(n29157) );
  NANDN U37971 ( .A(n29160), .B(n29161), .Z(n29159) );
  NANDN U37972 ( .A(n29161), .B(n29160), .Z(n29156) );
  AND U37973 ( .A(n29162), .B(n29163), .Z(n29151) );
  NAND U37974 ( .A(n29164), .B(n29165), .Z(n29163) );
  NANDN U37975 ( .A(n29166), .B(n29167), .Z(n29165) );
  NANDN U37976 ( .A(n29167), .B(n29166), .Z(n29162) );
  IV U37977 ( .A(n29168), .Z(n29167) );
  AND U37978 ( .A(n29169), .B(n29170), .Z(n29153) );
  NAND U37979 ( .A(n29171), .B(n29172), .Z(n29170) );
  NANDN U37980 ( .A(n29173), .B(n29174), .Z(n29172) );
  NANDN U37981 ( .A(n29174), .B(n29173), .Z(n29169) );
  XOR U37982 ( .A(n29166), .B(n29175), .Z(N62791) );
  XNOR U37983 ( .A(n29164), .B(n29168), .Z(n29175) );
  XOR U37984 ( .A(n29161), .B(n29176), .Z(n29168) );
  XNOR U37985 ( .A(n29158), .B(n29160), .Z(n29176) );
  AND U37986 ( .A(n29177), .B(n29178), .Z(n29160) );
  NANDN U37987 ( .A(n29179), .B(n29180), .Z(n29178) );
  OR U37988 ( .A(n29181), .B(n29182), .Z(n29180) );
  IV U37989 ( .A(n29183), .Z(n29182) );
  NANDN U37990 ( .A(n29183), .B(n29181), .Z(n29177) );
  AND U37991 ( .A(n29184), .B(n29185), .Z(n29158) );
  NAND U37992 ( .A(n29186), .B(n29187), .Z(n29185) );
  NANDN U37993 ( .A(n29188), .B(n29189), .Z(n29187) );
  NANDN U37994 ( .A(n29189), .B(n29188), .Z(n29184) );
  IV U37995 ( .A(n29190), .Z(n29189) );
  NAND U37996 ( .A(n29191), .B(n29192), .Z(n29161) );
  NANDN U37997 ( .A(n29193), .B(n29194), .Z(n29192) );
  NANDN U37998 ( .A(n29195), .B(n29196), .Z(n29194) );
  NANDN U37999 ( .A(n29196), .B(n29195), .Z(n29191) );
  IV U38000 ( .A(n29197), .Z(n29195) );
  AND U38001 ( .A(n29198), .B(n29199), .Z(n29164) );
  NAND U38002 ( .A(n29200), .B(n29201), .Z(n29199) );
  NANDN U38003 ( .A(n29202), .B(n29203), .Z(n29201) );
  NANDN U38004 ( .A(n29203), .B(n29202), .Z(n29198) );
  XOR U38005 ( .A(n29174), .B(n29204), .Z(n29166) );
  XNOR U38006 ( .A(n29171), .B(n29173), .Z(n29204) );
  AND U38007 ( .A(n29205), .B(n29206), .Z(n29173) );
  NANDN U38008 ( .A(n29207), .B(n29208), .Z(n29206) );
  OR U38009 ( .A(n29209), .B(n29210), .Z(n29208) );
  IV U38010 ( .A(n29211), .Z(n29210) );
  NANDN U38011 ( .A(n29211), .B(n29209), .Z(n29205) );
  AND U38012 ( .A(n29212), .B(n29213), .Z(n29171) );
  NAND U38013 ( .A(n29214), .B(n29215), .Z(n29213) );
  NANDN U38014 ( .A(n29216), .B(n29217), .Z(n29215) );
  NANDN U38015 ( .A(n29217), .B(n29216), .Z(n29212) );
  IV U38016 ( .A(n29218), .Z(n29217) );
  NAND U38017 ( .A(n29219), .B(n29220), .Z(n29174) );
  NANDN U38018 ( .A(n29221), .B(n29222), .Z(n29220) );
  NANDN U38019 ( .A(n29223), .B(n29224), .Z(n29222) );
  NANDN U38020 ( .A(n29224), .B(n29223), .Z(n29219) );
  IV U38021 ( .A(n29225), .Z(n29223) );
  XOR U38022 ( .A(n29200), .B(n29226), .Z(N62790) );
  XNOR U38023 ( .A(n29203), .B(n29202), .Z(n29226) );
  XNOR U38024 ( .A(n29214), .B(n29227), .Z(n29202) );
  XNOR U38025 ( .A(n29218), .B(n29216), .Z(n29227) );
  XOR U38026 ( .A(n29224), .B(n29228), .Z(n29216) );
  XNOR U38027 ( .A(n29221), .B(n29225), .Z(n29228) );
  AND U38028 ( .A(n29229), .B(n29230), .Z(n29225) );
  NAND U38029 ( .A(n29231), .B(n29232), .Z(n29230) );
  NAND U38030 ( .A(n29233), .B(n29234), .Z(n29229) );
  AND U38031 ( .A(n29235), .B(n29236), .Z(n29221) );
  NAND U38032 ( .A(n29237), .B(n29238), .Z(n29236) );
  NAND U38033 ( .A(n29239), .B(n29240), .Z(n29235) );
  NANDN U38034 ( .A(n29241), .B(n29242), .Z(n29224) );
  ANDN U38035 ( .B(n29243), .A(n29244), .Z(n29218) );
  XNOR U38036 ( .A(n29209), .B(n29245), .Z(n29214) );
  XNOR U38037 ( .A(n29207), .B(n29211), .Z(n29245) );
  AND U38038 ( .A(n29246), .B(n29247), .Z(n29211) );
  NAND U38039 ( .A(n29248), .B(n29249), .Z(n29247) );
  NAND U38040 ( .A(n29250), .B(n29251), .Z(n29246) );
  AND U38041 ( .A(n29252), .B(n29253), .Z(n29207) );
  NAND U38042 ( .A(n29254), .B(n29255), .Z(n29253) );
  NAND U38043 ( .A(n29256), .B(n29257), .Z(n29252) );
  AND U38044 ( .A(n29258), .B(n29259), .Z(n29209) );
  NAND U38045 ( .A(n29260), .B(n29261), .Z(n29203) );
  XNOR U38046 ( .A(n29186), .B(n29262), .Z(n29200) );
  XNOR U38047 ( .A(n29190), .B(n29188), .Z(n29262) );
  XOR U38048 ( .A(n29196), .B(n29263), .Z(n29188) );
  XNOR U38049 ( .A(n29193), .B(n29197), .Z(n29263) );
  AND U38050 ( .A(n29264), .B(n29265), .Z(n29197) );
  NAND U38051 ( .A(n29266), .B(n29267), .Z(n29265) );
  NAND U38052 ( .A(n29268), .B(n29269), .Z(n29264) );
  AND U38053 ( .A(n29270), .B(n29271), .Z(n29193) );
  NAND U38054 ( .A(n29272), .B(n29273), .Z(n29271) );
  NAND U38055 ( .A(n29274), .B(n29275), .Z(n29270) );
  NANDN U38056 ( .A(n29276), .B(n29277), .Z(n29196) );
  ANDN U38057 ( .B(n29278), .A(n29279), .Z(n29190) );
  XNOR U38058 ( .A(n29181), .B(n29280), .Z(n29186) );
  XNOR U38059 ( .A(n29179), .B(n29183), .Z(n29280) );
  AND U38060 ( .A(n29281), .B(n29282), .Z(n29183) );
  NAND U38061 ( .A(n29283), .B(n29284), .Z(n29282) );
  NAND U38062 ( .A(n29285), .B(n29286), .Z(n29281) );
  AND U38063 ( .A(n29287), .B(n29288), .Z(n29179) );
  NAND U38064 ( .A(n29289), .B(n29290), .Z(n29288) );
  NAND U38065 ( .A(n29291), .B(n29292), .Z(n29287) );
  AND U38066 ( .A(n29293), .B(n29294), .Z(n29181) );
  XOR U38067 ( .A(n29261), .B(n29260), .Z(N62789) );
  XNOR U38068 ( .A(n29278), .B(n29279), .Z(n29260) );
  XNOR U38069 ( .A(n29293), .B(n29294), .Z(n29279) );
  XOR U38070 ( .A(n29290), .B(n29289), .Z(n29294) );
  XOR U38071 ( .A(y[4068]), .B(x[4068]), .Z(n29289) );
  XOR U38072 ( .A(n29292), .B(n29291), .Z(n29290) );
  XOR U38073 ( .A(y[4070]), .B(x[4070]), .Z(n29291) );
  XOR U38074 ( .A(y[4069]), .B(x[4069]), .Z(n29292) );
  XOR U38075 ( .A(n29284), .B(n29283), .Z(n29293) );
  XOR U38076 ( .A(n29286), .B(n29285), .Z(n29283) );
  XOR U38077 ( .A(y[4067]), .B(x[4067]), .Z(n29285) );
  XOR U38078 ( .A(y[4066]), .B(x[4066]), .Z(n29286) );
  XOR U38079 ( .A(y[4065]), .B(x[4065]), .Z(n29284) );
  XNOR U38080 ( .A(n29277), .B(n29276), .Z(n29278) );
  XNOR U38081 ( .A(n29273), .B(n29272), .Z(n29276) );
  XOR U38082 ( .A(n29275), .B(n29274), .Z(n29272) );
  XOR U38083 ( .A(y[4064]), .B(x[4064]), .Z(n29274) );
  XOR U38084 ( .A(y[4063]), .B(x[4063]), .Z(n29275) );
  XOR U38085 ( .A(y[4062]), .B(x[4062]), .Z(n29273) );
  XOR U38086 ( .A(n29267), .B(n29266), .Z(n29277) );
  XOR U38087 ( .A(n29269), .B(n29268), .Z(n29266) );
  XOR U38088 ( .A(y[4061]), .B(x[4061]), .Z(n29268) );
  XOR U38089 ( .A(y[4060]), .B(x[4060]), .Z(n29269) );
  XOR U38090 ( .A(y[4059]), .B(x[4059]), .Z(n29267) );
  XNOR U38091 ( .A(n29243), .B(n29244), .Z(n29261) );
  XNOR U38092 ( .A(n29258), .B(n29259), .Z(n29244) );
  XOR U38093 ( .A(n29255), .B(n29254), .Z(n29259) );
  XOR U38094 ( .A(y[4056]), .B(x[4056]), .Z(n29254) );
  XOR U38095 ( .A(n29257), .B(n29256), .Z(n29255) );
  XOR U38096 ( .A(y[4058]), .B(x[4058]), .Z(n29256) );
  XOR U38097 ( .A(y[4057]), .B(x[4057]), .Z(n29257) );
  XOR U38098 ( .A(n29249), .B(n29248), .Z(n29258) );
  XOR U38099 ( .A(n29251), .B(n29250), .Z(n29248) );
  XOR U38100 ( .A(y[4055]), .B(x[4055]), .Z(n29250) );
  XOR U38101 ( .A(y[4054]), .B(x[4054]), .Z(n29251) );
  XOR U38102 ( .A(y[4053]), .B(x[4053]), .Z(n29249) );
  XNOR U38103 ( .A(n29242), .B(n29241), .Z(n29243) );
  XNOR U38104 ( .A(n29238), .B(n29237), .Z(n29241) );
  XOR U38105 ( .A(n29240), .B(n29239), .Z(n29237) );
  XOR U38106 ( .A(y[4052]), .B(x[4052]), .Z(n29239) );
  XOR U38107 ( .A(y[4051]), .B(x[4051]), .Z(n29240) );
  XOR U38108 ( .A(y[4050]), .B(x[4050]), .Z(n29238) );
  XOR U38109 ( .A(n29232), .B(n29231), .Z(n29242) );
  XOR U38110 ( .A(n29234), .B(n29233), .Z(n29231) );
  XOR U38111 ( .A(y[4049]), .B(x[4049]), .Z(n29233) );
  XOR U38112 ( .A(y[4048]), .B(x[4048]), .Z(n29234) );
  XOR U38113 ( .A(y[4047]), .B(x[4047]), .Z(n29232) );
  NAND U38114 ( .A(n29295), .B(n29296), .Z(N62780) );
  NAND U38115 ( .A(n29297), .B(n29298), .Z(n29296) );
  NANDN U38116 ( .A(n29299), .B(n29300), .Z(n29298) );
  NANDN U38117 ( .A(n29300), .B(n29299), .Z(n29295) );
  XOR U38118 ( .A(n29299), .B(n29301), .Z(N62779) );
  XNOR U38119 ( .A(n29297), .B(n29300), .Z(n29301) );
  NAND U38120 ( .A(n29302), .B(n29303), .Z(n29300) );
  NAND U38121 ( .A(n29304), .B(n29305), .Z(n29303) );
  NANDN U38122 ( .A(n29306), .B(n29307), .Z(n29305) );
  NANDN U38123 ( .A(n29307), .B(n29306), .Z(n29302) );
  AND U38124 ( .A(n29308), .B(n29309), .Z(n29297) );
  NAND U38125 ( .A(n29310), .B(n29311), .Z(n29309) );
  NANDN U38126 ( .A(n29312), .B(n29313), .Z(n29311) );
  NANDN U38127 ( .A(n29313), .B(n29312), .Z(n29308) );
  IV U38128 ( .A(n29314), .Z(n29313) );
  AND U38129 ( .A(n29315), .B(n29316), .Z(n29299) );
  NAND U38130 ( .A(n29317), .B(n29318), .Z(n29316) );
  NANDN U38131 ( .A(n29319), .B(n29320), .Z(n29318) );
  NANDN U38132 ( .A(n29320), .B(n29319), .Z(n29315) );
  XOR U38133 ( .A(n29312), .B(n29321), .Z(N62778) );
  XNOR U38134 ( .A(n29310), .B(n29314), .Z(n29321) );
  XOR U38135 ( .A(n29307), .B(n29322), .Z(n29314) );
  XNOR U38136 ( .A(n29304), .B(n29306), .Z(n29322) );
  AND U38137 ( .A(n29323), .B(n29324), .Z(n29306) );
  NANDN U38138 ( .A(n29325), .B(n29326), .Z(n29324) );
  OR U38139 ( .A(n29327), .B(n29328), .Z(n29326) );
  IV U38140 ( .A(n29329), .Z(n29328) );
  NANDN U38141 ( .A(n29329), .B(n29327), .Z(n29323) );
  AND U38142 ( .A(n29330), .B(n29331), .Z(n29304) );
  NAND U38143 ( .A(n29332), .B(n29333), .Z(n29331) );
  NANDN U38144 ( .A(n29334), .B(n29335), .Z(n29333) );
  NANDN U38145 ( .A(n29335), .B(n29334), .Z(n29330) );
  IV U38146 ( .A(n29336), .Z(n29335) );
  NAND U38147 ( .A(n29337), .B(n29338), .Z(n29307) );
  NANDN U38148 ( .A(n29339), .B(n29340), .Z(n29338) );
  NANDN U38149 ( .A(n29341), .B(n29342), .Z(n29340) );
  NANDN U38150 ( .A(n29342), .B(n29341), .Z(n29337) );
  IV U38151 ( .A(n29343), .Z(n29341) );
  AND U38152 ( .A(n29344), .B(n29345), .Z(n29310) );
  NAND U38153 ( .A(n29346), .B(n29347), .Z(n29345) );
  NANDN U38154 ( .A(n29348), .B(n29349), .Z(n29347) );
  NANDN U38155 ( .A(n29349), .B(n29348), .Z(n29344) );
  XOR U38156 ( .A(n29320), .B(n29350), .Z(n29312) );
  XNOR U38157 ( .A(n29317), .B(n29319), .Z(n29350) );
  AND U38158 ( .A(n29351), .B(n29352), .Z(n29319) );
  NANDN U38159 ( .A(n29353), .B(n29354), .Z(n29352) );
  OR U38160 ( .A(n29355), .B(n29356), .Z(n29354) );
  IV U38161 ( .A(n29357), .Z(n29356) );
  NANDN U38162 ( .A(n29357), .B(n29355), .Z(n29351) );
  AND U38163 ( .A(n29358), .B(n29359), .Z(n29317) );
  NAND U38164 ( .A(n29360), .B(n29361), .Z(n29359) );
  NANDN U38165 ( .A(n29362), .B(n29363), .Z(n29361) );
  NANDN U38166 ( .A(n29363), .B(n29362), .Z(n29358) );
  IV U38167 ( .A(n29364), .Z(n29363) );
  NAND U38168 ( .A(n29365), .B(n29366), .Z(n29320) );
  NANDN U38169 ( .A(n29367), .B(n29368), .Z(n29366) );
  NANDN U38170 ( .A(n29369), .B(n29370), .Z(n29368) );
  NANDN U38171 ( .A(n29370), .B(n29369), .Z(n29365) );
  IV U38172 ( .A(n29371), .Z(n29369) );
  XOR U38173 ( .A(n29346), .B(n29372), .Z(N62777) );
  XNOR U38174 ( .A(n29349), .B(n29348), .Z(n29372) );
  XNOR U38175 ( .A(n29360), .B(n29373), .Z(n29348) );
  XNOR U38176 ( .A(n29364), .B(n29362), .Z(n29373) );
  XOR U38177 ( .A(n29370), .B(n29374), .Z(n29362) );
  XNOR U38178 ( .A(n29367), .B(n29371), .Z(n29374) );
  AND U38179 ( .A(n29375), .B(n29376), .Z(n29371) );
  NAND U38180 ( .A(n29377), .B(n29378), .Z(n29376) );
  NAND U38181 ( .A(n29379), .B(n29380), .Z(n29375) );
  AND U38182 ( .A(n29381), .B(n29382), .Z(n29367) );
  NAND U38183 ( .A(n29383), .B(n29384), .Z(n29382) );
  NAND U38184 ( .A(n29385), .B(n29386), .Z(n29381) );
  NANDN U38185 ( .A(n29387), .B(n29388), .Z(n29370) );
  ANDN U38186 ( .B(n29389), .A(n29390), .Z(n29364) );
  XNOR U38187 ( .A(n29355), .B(n29391), .Z(n29360) );
  XNOR U38188 ( .A(n29353), .B(n29357), .Z(n29391) );
  AND U38189 ( .A(n29392), .B(n29393), .Z(n29357) );
  NAND U38190 ( .A(n29394), .B(n29395), .Z(n29393) );
  NAND U38191 ( .A(n29396), .B(n29397), .Z(n29392) );
  AND U38192 ( .A(n29398), .B(n29399), .Z(n29353) );
  NAND U38193 ( .A(n29400), .B(n29401), .Z(n29399) );
  NAND U38194 ( .A(n29402), .B(n29403), .Z(n29398) );
  AND U38195 ( .A(n29404), .B(n29405), .Z(n29355) );
  NAND U38196 ( .A(n29406), .B(n29407), .Z(n29349) );
  XNOR U38197 ( .A(n29332), .B(n29408), .Z(n29346) );
  XNOR U38198 ( .A(n29336), .B(n29334), .Z(n29408) );
  XOR U38199 ( .A(n29342), .B(n29409), .Z(n29334) );
  XNOR U38200 ( .A(n29339), .B(n29343), .Z(n29409) );
  AND U38201 ( .A(n29410), .B(n29411), .Z(n29343) );
  NAND U38202 ( .A(n29412), .B(n29413), .Z(n29411) );
  NAND U38203 ( .A(n29414), .B(n29415), .Z(n29410) );
  AND U38204 ( .A(n29416), .B(n29417), .Z(n29339) );
  NAND U38205 ( .A(n29418), .B(n29419), .Z(n29417) );
  NAND U38206 ( .A(n29420), .B(n29421), .Z(n29416) );
  NANDN U38207 ( .A(n29422), .B(n29423), .Z(n29342) );
  ANDN U38208 ( .B(n29424), .A(n29425), .Z(n29336) );
  XNOR U38209 ( .A(n29327), .B(n29426), .Z(n29332) );
  XNOR U38210 ( .A(n29325), .B(n29329), .Z(n29426) );
  AND U38211 ( .A(n29427), .B(n29428), .Z(n29329) );
  NAND U38212 ( .A(n29429), .B(n29430), .Z(n29428) );
  NAND U38213 ( .A(n29431), .B(n29432), .Z(n29427) );
  AND U38214 ( .A(n29433), .B(n29434), .Z(n29325) );
  NAND U38215 ( .A(n29435), .B(n29436), .Z(n29434) );
  NAND U38216 ( .A(n29437), .B(n29438), .Z(n29433) );
  AND U38217 ( .A(n29439), .B(n29440), .Z(n29327) );
  XOR U38218 ( .A(n29407), .B(n29406), .Z(N62776) );
  XNOR U38219 ( .A(n29424), .B(n29425), .Z(n29406) );
  XNOR U38220 ( .A(n29439), .B(n29440), .Z(n29425) );
  XOR U38221 ( .A(n29436), .B(n29435), .Z(n29440) );
  XOR U38222 ( .A(y[4044]), .B(x[4044]), .Z(n29435) );
  XOR U38223 ( .A(n29438), .B(n29437), .Z(n29436) );
  XOR U38224 ( .A(y[4046]), .B(x[4046]), .Z(n29437) );
  XOR U38225 ( .A(y[4045]), .B(x[4045]), .Z(n29438) );
  XOR U38226 ( .A(n29430), .B(n29429), .Z(n29439) );
  XOR U38227 ( .A(n29432), .B(n29431), .Z(n29429) );
  XOR U38228 ( .A(y[4043]), .B(x[4043]), .Z(n29431) );
  XOR U38229 ( .A(y[4042]), .B(x[4042]), .Z(n29432) );
  XOR U38230 ( .A(y[4041]), .B(x[4041]), .Z(n29430) );
  XNOR U38231 ( .A(n29423), .B(n29422), .Z(n29424) );
  XNOR U38232 ( .A(n29419), .B(n29418), .Z(n29422) );
  XOR U38233 ( .A(n29421), .B(n29420), .Z(n29418) );
  XOR U38234 ( .A(y[4040]), .B(x[4040]), .Z(n29420) );
  XOR U38235 ( .A(y[4039]), .B(x[4039]), .Z(n29421) );
  XOR U38236 ( .A(y[4038]), .B(x[4038]), .Z(n29419) );
  XOR U38237 ( .A(n29413), .B(n29412), .Z(n29423) );
  XOR U38238 ( .A(n29415), .B(n29414), .Z(n29412) );
  XOR U38239 ( .A(y[4037]), .B(x[4037]), .Z(n29414) );
  XOR U38240 ( .A(y[4036]), .B(x[4036]), .Z(n29415) );
  XOR U38241 ( .A(y[4035]), .B(x[4035]), .Z(n29413) );
  XNOR U38242 ( .A(n29389), .B(n29390), .Z(n29407) );
  XNOR U38243 ( .A(n29404), .B(n29405), .Z(n29390) );
  XOR U38244 ( .A(n29401), .B(n29400), .Z(n29405) );
  XOR U38245 ( .A(y[4032]), .B(x[4032]), .Z(n29400) );
  XOR U38246 ( .A(n29403), .B(n29402), .Z(n29401) );
  XOR U38247 ( .A(y[4034]), .B(x[4034]), .Z(n29402) );
  XOR U38248 ( .A(y[4033]), .B(x[4033]), .Z(n29403) );
  XOR U38249 ( .A(n29395), .B(n29394), .Z(n29404) );
  XOR U38250 ( .A(n29397), .B(n29396), .Z(n29394) );
  XOR U38251 ( .A(y[4031]), .B(x[4031]), .Z(n29396) );
  XOR U38252 ( .A(y[4030]), .B(x[4030]), .Z(n29397) );
  XOR U38253 ( .A(y[4029]), .B(x[4029]), .Z(n29395) );
  XNOR U38254 ( .A(n29388), .B(n29387), .Z(n29389) );
  XNOR U38255 ( .A(n29384), .B(n29383), .Z(n29387) );
  XOR U38256 ( .A(n29386), .B(n29385), .Z(n29383) );
  XOR U38257 ( .A(y[4028]), .B(x[4028]), .Z(n29385) );
  XOR U38258 ( .A(y[4027]), .B(x[4027]), .Z(n29386) );
  XOR U38259 ( .A(y[4026]), .B(x[4026]), .Z(n29384) );
  XOR U38260 ( .A(n29378), .B(n29377), .Z(n29388) );
  XOR U38261 ( .A(n29380), .B(n29379), .Z(n29377) );
  XOR U38262 ( .A(y[4025]), .B(x[4025]), .Z(n29379) );
  XOR U38263 ( .A(y[4024]), .B(x[4024]), .Z(n29380) );
  XOR U38264 ( .A(y[4023]), .B(x[4023]), .Z(n29378) );
  NAND U38265 ( .A(n29441), .B(n29442), .Z(N62767) );
  NAND U38266 ( .A(n29443), .B(n29444), .Z(n29442) );
  NANDN U38267 ( .A(n29445), .B(n29446), .Z(n29444) );
  NANDN U38268 ( .A(n29446), .B(n29445), .Z(n29441) );
  XOR U38269 ( .A(n29445), .B(n29447), .Z(N62766) );
  XNOR U38270 ( .A(n29443), .B(n29446), .Z(n29447) );
  NAND U38271 ( .A(n29448), .B(n29449), .Z(n29446) );
  NAND U38272 ( .A(n29450), .B(n29451), .Z(n29449) );
  NANDN U38273 ( .A(n29452), .B(n29453), .Z(n29451) );
  NANDN U38274 ( .A(n29453), .B(n29452), .Z(n29448) );
  AND U38275 ( .A(n29454), .B(n29455), .Z(n29443) );
  NAND U38276 ( .A(n29456), .B(n29457), .Z(n29455) );
  NANDN U38277 ( .A(n29458), .B(n29459), .Z(n29457) );
  NANDN U38278 ( .A(n29459), .B(n29458), .Z(n29454) );
  IV U38279 ( .A(n29460), .Z(n29459) );
  AND U38280 ( .A(n29461), .B(n29462), .Z(n29445) );
  NAND U38281 ( .A(n29463), .B(n29464), .Z(n29462) );
  NANDN U38282 ( .A(n29465), .B(n29466), .Z(n29464) );
  NANDN U38283 ( .A(n29466), .B(n29465), .Z(n29461) );
  XOR U38284 ( .A(n29458), .B(n29467), .Z(N62765) );
  XNOR U38285 ( .A(n29456), .B(n29460), .Z(n29467) );
  XOR U38286 ( .A(n29453), .B(n29468), .Z(n29460) );
  XNOR U38287 ( .A(n29450), .B(n29452), .Z(n29468) );
  AND U38288 ( .A(n29469), .B(n29470), .Z(n29452) );
  NANDN U38289 ( .A(n29471), .B(n29472), .Z(n29470) );
  OR U38290 ( .A(n29473), .B(n29474), .Z(n29472) );
  IV U38291 ( .A(n29475), .Z(n29474) );
  NANDN U38292 ( .A(n29475), .B(n29473), .Z(n29469) );
  AND U38293 ( .A(n29476), .B(n29477), .Z(n29450) );
  NAND U38294 ( .A(n29478), .B(n29479), .Z(n29477) );
  NANDN U38295 ( .A(n29480), .B(n29481), .Z(n29479) );
  NANDN U38296 ( .A(n29481), .B(n29480), .Z(n29476) );
  IV U38297 ( .A(n29482), .Z(n29481) );
  NAND U38298 ( .A(n29483), .B(n29484), .Z(n29453) );
  NANDN U38299 ( .A(n29485), .B(n29486), .Z(n29484) );
  NANDN U38300 ( .A(n29487), .B(n29488), .Z(n29486) );
  NANDN U38301 ( .A(n29488), .B(n29487), .Z(n29483) );
  IV U38302 ( .A(n29489), .Z(n29487) );
  AND U38303 ( .A(n29490), .B(n29491), .Z(n29456) );
  NAND U38304 ( .A(n29492), .B(n29493), .Z(n29491) );
  NANDN U38305 ( .A(n29494), .B(n29495), .Z(n29493) );
  NANDN U38306 ( .A(n29495), .B(n29494), .Z(n29490) );
  XOR U38307 ( .A(n29466), .B(n29496), .Z(n29458) );
  XNOR U38308 ( .A(n29463), .B(n29465), .Z(n29496) );
  AND U38309 ( .A(n29497), .B(n29498), .Z(n29465) );
  NANDN U38310 ( .A(n29499), .B(n29500), .Z(n29498) );
  OR U38311 ( .A(n29501), .B(n29502), .Z(n29500) );
  IV U38312 ( .A(n29503), .Z(n29502) );
  NANDN U38313 ( .A(n29503), .B(n29501), .Z(n29497) );
  AND U38314 ( .A(n29504), .B(n29505), .Z(n29463) );
  NAND U38315 ( .A(n29506), .B(n29507), .Z(n29505) );
  NANDN U38316 ( .A(n29508), .B(n29509), .Z(n29507) );
  NANDN U38317 ( .A(n29509), .B(n29508), .Z(n29504) );
  IV U38318 ( .A(n29510), .Z(n29509) );
  NAND U38319 ( .A(n29511), .B(n29512), .Z(n29466) );
  NANDN U38320 ( .A(n29513), .B(n29514), .Z(n29512) );
  NANDN U38321 ( .A(n29515), .B(n29516), .Z(n29514) );
  NANDN U38322 ( .A(n29516), .B(n29515), .Z(n29511) );
  IV U38323 ( .A(n29517), .Z(n29515) );
  XOR U38324 ( .A(n29492), .B(n29518), .Z(N62764) );
  XNOR U38325 ( .A(n29495), .B(n29494), .Z(n29518) );
  XNOR U38326 ( .A(n29506), .B(n29519), .Z(n29494) );
  XNOR U38327 ( .A(n29510), .B(n29508), .Z(n29519) );
  XOR U38328 ( .A(n29516), .B(n29520), .Z(n29508) );
  XNOR U38329 ( .A(n29513), .B(n29517), .Z(n29520) );
  AND U38330 ( .A(n29521), .B(n29522), .Z(n29517) );
  NAND U38331 ( .A(n29523), .B(n29524), .Z(n29522) );
  NAND U38332 ( .A(n29525), .B(n29526), .Z(n29521) );
  AND U38333 ( .A(n29527), .B(n29528), .Z(n29513) );
  NAND U38334 ( .A(n29529), .B(n29530), .Z(n29528) );
  NAND U38335 ( .A(n29531), .B(n29532), .Z(n29527) );
  NANDN U38336 ( .A(n29533), .B(n29534), .Z(n29516) );
  ANDN U38337 ( .B(n29535), .A(n29536), .Z(n29510) );
  XNOR U38338 ( .A(n29501), .B(n29537), .Z(n29506) );
  XNOR U38339 ( .A(n29499), .B(n29503), .Z(n29537) );
  AND U38340 ( .A(n29538), .B(n29539), .Z(n29503) );
  NAND U38341 ( .A(n29540), .B(n29541), .Z(n29539) );
  NAND U38342 ( .A(n29542), .B(n29543), .Z(n29538) );
  AND U38343 ( .A(n29544), .B(n29545), .Z(n29499) );
  NAND U38344 ( .A(n29546), .B(n29547), .Z(n29545) );
  NAND U38345 ( .A(n29548), .B(n29549), .Z(n29544) );
  AND U38346 ( .A(n29550), .B(n29551), .Z(n29501) );
  NAND U38347 ( .A(n29552), .B(n29553), .Z(n29495) );
  XNOR U38348 ( .A(n29478), .B(n29554), .Z(n29492) );
  XNOR U38349 ( .A(n29482), .B(n29480), .Z(n29554) );
  XOR U38350 ( .A(n29488), .B(n29555), .Z(n29480) );
  XNOR U38351 ( .A(n29485), .B(n29489), .Z(n29555) );
  AND U38352 ( .A(n29556), .B(n29557), .Z(n29489) );
  NAND U38353 ( .A(n29558), .B(n29559), .Z(n29557) );
  NAND U38354 ( .A(n29560), .B(n29561), .Z(n29556) );
  AND U38355 ( .A(n29562), .B(n29563), .Z(n29485) );
  NAND U38356 ( .A(n29564), .B(n29565), .Z(n29563) );
  NAND U38357 ( .A(n29566), .B(n29567), .Z(n29562) );
  NANDN U38358 ( .A(n29568), .B(n29569), .Z(n29488) );
  ANDN U38359 ( .B(n29570), .A(n29571), .Z(n29482) );
  XNOR U38360 ( .A(n29473), .B(n29572), .Z(n29478) );
  XNOR U38361 ( .A(n29471), .B(n29475), .Z(n29572) );
  AND U38362 ( .A(n29573), .B(n29574), .Z(n29475) );
  NAND U38363 ( .A(n29575), .B(n29576), .Z(n29574) );
  NAND U38364 ( .A(n29577), .B(n29578), .Z(n29573) );
  AND U38365 ( .A(n29579), .B(n29580), .Z(n29471) );
  NAND U38366 ( .A(n29581), .B(n29582), .Z(n29580) );
  NAND U38367 ( .A(n29583), .B(n29584), .Z(n29579) );
  AND U38368 ( .A(n29585), .B(n29586), .Z(n29473) );
  XOR U38369 ( .A(n29553), .B(n29552), .Z(N62763) );
  XNOR U38370 ( .A(n29570), .B(n29571), .Z(n29552) );
  XNOR U38371 ( .A(n29585), .B(n29586), .Z(n29571) );
  XOR U38372 ( .A(n29582), .B(n29581), .Z(n29586) );
  XOR U38373 ( .A(y[4020]), .B(x[4020]), .Z(n29581) );
  XOR U38374 ( .A(n29584), .B(n29583), .Z(n29582) );
  XOR U38375 ( .A(y[4022]), .B(x[4022]), .Z(n29583) );
  XOR U38376 ( .A(y[4021]), .B(x[4021]), .Z(n29584) );
  XOR U38377 ( .A(n29576), .B(n29575), .Z(n29585) );
  XOR U38378 ( .A(n29578), .B(n29577), .Z(n29575) );
  XOR U38379 ( .A(y[4019]), .B(x[4019]), .Z(n29577) );
  XOR U38380 ( .A(y[4018]), .B(x[4018]), .Z(n29578) );
  XOR U38381 ( .A(y[4017]), .B(x[4017]), .Z(n29576) );
  XNOR U38382 ( .A(n29569), .B(n29568), .Z(n29570) );
  XNOR U38383 ( .A(n29565), .B(n29564), .Z(n29568) );
  XOR U38384 ( .A(n29567), .B(n29566), .Z(n29564) );
  XOR U38385 ( .A(y[4016]), .B(x[4016]), .Z(n29566) );
  XOR U38386 ( .A(y[4015]), .B(x[4015]), .Z(n29567) );
  XOR U38387 ( .A(y[4014]), .B(x[4014]), .Z(n29565) );
  XOR U38388 ( .A(n29559), .B(n29558), .Z(n29569) );
  XOR U38389 ( .A(n29561), .B(n29560), .Z(n29558) );
  XOR U38390 ( .A(y[4013]), .B(x[4013]), .Z(n29560) );
  XOR U38391 ( .A(y[4012]), .B(x[4012]), .Z(n29561) );
  XOR U38392 ( .A(y[4011]), .B(x[4011]), .Z(n29559) );
  XNOR U38393 ( .A(n29535), .B(n29536), .Z(n29553) );
  XNOR U38394 ( .A(n29550), .B(n29551), .Z(n29536) );
  XOR U38395 ( .A(n29547), .B(n29546), .Z(n29551) );
  XOR U38396 ( .A(y[4008]), .B(x[4008]), .Z(n29546) );
  XOR U38397 ( .A(n29549), .B(n29548), .Z(n29547) );
  XOR U38398 ( .A(y[4010]), .B(x[4010]), .Z(n29548) );
  XOR U38399 ( .A(y[4009]), .B(x[4009]), .Z(n29549) );
  XOR U38400 ( .A(n29541), .B(n29540), .Z(n29550) );
  XOR U38401 ( .A(n29543), .B(n29542), .Z(n29540) );
  XOR U38402 ( .A(y[4007]), .B(x[4007]), .Z(n29542) );
  XOR U38403 ( .A(y[4006]), .B(x[4006]), .Z(n29543) );
  XOR U38404 ( .A(y[4005]), .B(x[4005]), .Z(n29541) );
  XNOR U38405 ( .A(n29534), .B(n29533), .Z(n29535) );
  XNOR U38406 ( .A(n29530), .B(n29529), .Z(n29533) );
  XOR U38407 ( .A(n29532), .B(n29531), .Z(n29529) );
  XOR U38408 ( .A(y[4004]), .B(x[4004]), .Z(n29531) );
  XOR U38409 ( .A(y[4003]), .B(x[4003]), .Z(n29532) );
  XOR U38410 ( .A(y[4002]), .B(x[4002]), .Z(n29530) );
  XOR U38411 ( .A(n29524), .B(n29523), .Z(n29534) );
  XOR U38412 ( .A(n29526), .B(n29525), .Z(n29523) );
  XOR U38413 ( .A(y[4001]), .B(x[4001]), .Z(n29525) );
  XOR U38414 ( .A(y[4000]), .B(x[4000]), .Z(n29526) );
  XOR U38415 ( .A(y[3999]), .B(x[3999]), .Z(n29524) );
  NAND U38416 ( .A(n29587), .B(n29588), .Z(N62754) );
  NAND U38417 ( .A(n29589), .B(n29590), .Z(n29588) );
  NANDN U38418 ( .A(n29591), .B(n29592), .Z(n29590) );
  NANDN U38419 ( .A(n29592), .B(n29591), .Z(n29587) );
  XOR U38420 ( .A(n29591), .B(n29593), .Z(N62753) );
  XNOR U38421 ( .A(n29589), .B(n29592), .Z(n29593) );
  NAND U38422 ( .A(n29594), .B(n29595), .Z(n29592) );
  NAND U38423 ( .A(n29596), .B(n29597), .Z(n29595) );
  NANDN U38424 ( .A(n29598), .B(n29599), .Z(n29597) );
  NANDN U38425 ( .A(n29599), .B(n29598), .Z(n29594) );
  AND U38426 ( .A(n29600), .B(n29601), .Z(n29589) );
  NAND U38427 ( .A(n29602), .B(n29603), .Z(n29601) );
  NANDN U38428 ( .A(n29604), .B(n29605), .Z(n29603) );
  NANDN U38429 ( .A(n29605), .B(n29604), .Z(n29600) );
  IV U38430 ( .A(n29606), .Z(n29605) );
  AND U38431 ( .A(n29607), .B(n29608), .Z(n29591) );
  NAND U38432 ( .A(n29609), .B(n29610), .Z(n29608) );
  NANDN U38433 ( .A(n29611), .B(n29612), .Z(n29610) );
  NANDN U38434 ( .A(n29612), .B(n29611), .Z(n29607) );
  XOR U38435 ( .A(n29604), .B(n29613), .Z(N62752) );
  XNOR U38436 ( .A(n29602), .B(n29606), .Z(n29613) );
  XOR U38437 ( .A(n29599), .B(n29614), .Z(n29606) );
  XNOR U38438 ( .A(n29596), .B(n29598), .Z(n29614) );
  AND U38439 ( .A(n29615), .B(n29616), .Z(n29598) );
  NANDN U38440 ( .A(n29617), .B(n29618), .Z(n29616) );
  OR U38441 ( .A(n29619), .B(n29620), .Z(n29618) );
  IV U38442 ( .A(n29621), .Z(n29620) );
  NANDN U38443 ( .A(n29621), .B(n29619), .Z(n29615) );
  AND U38444 ( .A(n29622), .B(n29623), .Z(n29596) );
  NAND U38445 ( .A(n29624), .B(n29625), .Z(n29623) );
  NANDN U38446 ( .A(n29626), .B(n29627), .Z(n29625) );
  NANDN U38447 ( .A(n29627), .B(n29626), .Z(n29622) );
  IV U38448 ( .A(n29628), .Z(n29627) );
  NAND U38449 ( .A(n29629), .B(n29630), .Z(n29599) );
  NANDN U38450 ( .A(n29631), .B(n29632), .Z(n29630) );
  NANDN U38451 ( .A(n29633), .B(n29634), .Z(n29632) );
  NANDN U38452 ( .A(n29634), .B(n29633), .Z(n29629) );
  IV U38453 ( .A(n29635), .Z(n29633) );
  AND U38454 ( .A(n29636), .B(n29637), .Z(n29602) );
  NAND U38455 ( .A(n29638), .B(n29639), .Z(n29637) );
  NANDN U38456 ( .A(n29640), .B(n29641), .Z(n29639) );
  NANDN U38457 ( .A(n29641), .B(n29640), .Z(n29636) );
  XOR U38458 ( .A(n29612), .B(n29642), .Z(n29604) );
  XNOR U38459 ( .A(n29609), .B(n29611), .Z(n29642) );
  AND U38460 ( .A(n29643), .B(n29644), .Z(n29611) );
  NANDN U38461 ( .A(n29645), .B(n29646), .Z(n29644) );
  OR U38462 ( .A(n29647), .B(n29648), .Z(n29646) );
  IV U38463 ( .A(n29649), .Z(n29648) );
  NANDN U38464 ( .A(n29649), .B(n29647), .Z(n29643) );
  AND U38465 ( .A(n29650), .B(n29651), .Z(n29609) );
  NAND U38466 ( .A(n29652), .B(n29653), .Z(n29651) );
  NANDN U38467 ( .A(n29654), .B(n29655), .Z(n29653) );
  NANDN U38468 ( .A(n29655), .B(n29654), .Z(n29650) );
  IV U38469 ( .A(n29656), .Z(n29655) );
  NAND U38470 ( .A(n29657), .B(n29658), .Z(n29612) );
  NANDN U38471 ( .A(n29659), .B(n29660), .Z(n29658) );
  NANDN U38472 ( .A(n29661), .B(n29662), .Z(n29660) );
  NANDN U38473 ( .A(n29662), .B(n29661), .Z(n29657) );
  IV U38474 ( .A(n29663), .Z(n29661) );
  XOR U38475 ( .A(n29638), .B(n29664), .Z(N62751) );
  XNOR U38476 ( .A(n29641), .B(n29640), .Z(n29664) );
  XNOR U38477 ( .A(n29652), .B(n29665), .Z(n29640) );
  XNOR U38478 ( .A(n29656), .B(n29654), .Z(n29665) );
  XOR U38479 ( .A(n29662), .B(n29666), .Z(n29654) );
  XNOR U38480 ( .A(n29659), .B(n29663), .Z(n29666) );
  AND U38481 ( .A(n29667), .B(n29668), .Z(n29663) );
  NAND U38482 ( .A(n29669), .B(n29670), .Z(n29668) );
  NAND U38483 ( .A(n29671), .B(n29672), .Z(n29667) );
  AND U38484 ( .A(n29673), .B(n29674), .Z(n29659) );
  NAND U38485 ( .A(n29675), .B(n29676), .Z(n29674) );
  NAND U38486 ( .A(n29677), .B(n29678), .Z(n29673) );
  NANDN U38487 ( .A(n29679), .B(n29680), .Z(n29662) );
  ANDN U38488 ( .B(n29681), .A(n29682), .Z(n29656) );
  XNOR U38489 ( .A(n29647), .B(n29683), .Z(n29652) );
  XNOR U38490 ( .A(n29645), .B(n29649), .Z(n29683) );
  AND U38491 ( .A(n29684), .B(n29685), .Z(n29649) );
  NAND U38492 ( .A(n29686), .B(n29687), .Z(n29685) );
  NAND U38493 ( .A(n29688), .B(n29689), .Z(n29684) );
  AND U38494 ( .A(n29690), .B(n29691), .Z(n29645) );
  NAND U38495 ( .A(n29692), .B(n29693), .Z(n29691) );
  NAND U38496 ( .A(n29694), .B(n29695), .Z(n29690) );
  AND U38497 ( .A(n29696), .B(n29697), .Z(n29647) );
  NAND U38498 ( .A(n29698), .B(n29699), .Z(n29641) );
  XNOR U38499 ( .A(n29624), .B(n29700), .Z(n29638) );
  XNOR U38500 ( .A(n29628), .B(n29626), .Z(n29700) );
  XOR U38501 ( .A(n29634), .B(n29701), .Z(n29626) );
  XNOR U38502 ( .A(n29631), .B(n29635), .Z(n29701) );
  AND U38503 ( .A(n29702), .B(n29703), .Z(n29635) );
  NAND U38504 ( .A(n29704), .B(n29705), .Z(n29703) );
  NAND U38505 ( .A(n29706), .B(n29707), .Z(n29702) );
  AND U38506 ( .A(n29708), .B(n29709), .Z(n29631) );
  NAND U38507 ( .A(n29710), .B(n29711), .Z(n29709) );
  NAND U38508 ( .A(n29712), .B(n29713), .Z(n29708) );
  NANDN U38509 ( .A(n29714), .B(n29715), .Z(n29634) );
  ANDN U38510 ( .B(n29716), .A(n29717), .Z(n29628) );
  XNOR U38511 ( .A(n29619), .B(n29718), .Z(n29624) );
  XNOR U38512 ( .A(n29617), .B(n29621), .Z(n29718) );
  AND U38513 ( .A(n29719), .B(n29720), .Z(n29621) );
  NAND U38514 ( .A(n29721), .B(n29722), .Z(n29720) );
  NAND U38515 ( .A(n29723), .B(n29724), .Z(n29719) );
  AND U38516 ( .A(n29725), .B(n29726), .Z(n29617) );
  NAND U38517 ( .A(n29727), .B(n29728), .Z(n29726) );
  NAND U38518 ( .A(n29729), .B(n29730), .Z(n29725) );
  AND U38519 ( .A(n29731), .B(n29732), .Z(n29619) );
  XOR U38520 ( .A(n29699), .B(n29698), .Z(N62750) );
  XNOR U38521 ( .A(n29716), .B(n29717), .Z(n29698) );
  XNOR U38522 ( .A(n29731), .B(n29732), .Z(n29717) );
  XOR U38523 ( .A(n29728), .B(n29727), .Z(n29732) );
  XOR U38524 ( .A(y[3996]), .B(x[3996]), .Z(n29727) );
  XOR U38525 ( .A(n29730), .B(n29729), .Z(n29728) );
  XOR U38526 ( .A(y[3998]), .B(x[3998]), .Z(n29729) );
  XOR U38527 ( .A(y[3997]), .B(x[3997]), .Z(n29730) );
  XOR U38528 ( .A(n29722), .B(n29721), .Z(n29731) );
  XOR U38529 ( .A(n29724), .B(n29723), .Z(n29721) );
  XOR U38530 ( .A(y[3995]), .B(x[3995]), .Z(n29723) );
  XOR U38531 ( .A(y[3994]), .B(x[3994]), .Z(n29724) );
  XOR U38532 ( .A(y[3993]), .B(x[3993]), .Z(n29722) );
  XNOR U38533 ( .A(n29715), .B(n29714), .Z(n29716) );
  XNOR U38534 ( .A(n29711), .B(n29710), .Z(n29714) );
  XOR U38535 ( .A(n29713), .B(n29712), .Z(n29710) );
  XOR U38536 ( .A(y[3992]), .B(x[3992]), .Z(n29712) );
  XOR U38537 ( .A(y[3991]), .B(x[3991]), .Z(n29713) );
  XOR U38538 ( .A(y[3990]), .B(x[3990]), .Z(n29711) );
  XOR U38539 ( .A(n29705), .B(n29704), .Z(n29715) );
  XOR U38540 ( .A(n29707), .B(n29706), .Z(n29704) );
  XOR U38541 ( .A(y[3989]), .B(x[3989]), .Z(n29706) );
  XOR U38542 ( .A(y[3988]), .B(x[3988]), .Z(n29707) );
  XOR U38543 ( .A(y[3987]), .B(x[3987]), .Z(n29705) );
  XNOR U38544 ( .A(n29681), .B(n29682), .Z(n29699) );
  XNOR U38545 ( .A(n29696), .B(n29697), .Z(n29682) );
  XOR U38546 ( .A(n29693), .B(n29692), .Z(n29697) );
  XOR U38547 ( .A(y[3984]), .B(x[3984]), .Z(n29692) );
  XOR U38548 ( .A(n29695), .B(n29694), .Z(n29693) );
  XOR U38549 ( .A(y[3986]), .B(x[3986]), .Z(n29694) );
  XOR U38550 ( .A(y[3985]), .B(x[3985]), .Z(n29695) );
  XOR U38551 ( .A(n29687), .B(n29686), .Z(n29696) );
  XOR U38552 ( .A(n29689), .B(n29688), .Z(n29686) );
  XOR U38553 ( .A(y[3983]), .B(x[3983]), .Z(n29688) );
  XOR U38554 ( .A(y[3982]), .B(x[3982]), .Z(n29689) );
  XOR U38555 ( .A(y[3981]), .B(x[3981]), .Z(n29687) );
  XNOR U38556 ( .A(n29680), .B(n29679), .Z(n29681) );
  XNOR U38557 ( .A(n29676), .B(n29675), .Z(n29679) );
  XOR U38558 ( .A(n29678), .B(n29677), .Z(n29675) );
  XOR U38559 ( .A(y[3980]), .B(x[3980]), .Z(n29677) );
  XOR U38560 ( .A(y[3979]), .B(x[3979]), .Z(n29678) );
  XOR U38561 ( .A(y[3978]), .B(x[3978]), .Z(n29676) );
  XOR U38562 ( .A(n29670), .B(n29669), .Z(n29680) );
  XOR U38563 ( .A(n29672), .B(n29671), .Z(n29669) );
  XOR U38564 ( .A(y[3977]), .B(x[3977]), .Z(n29671) );
  XOR U38565 ( .A(y[3976]), .B(x[3976]), .Z(n29672) );
  XOR U38566 ( .A(y[3975]), .B(x[3975]), .Z(n29670) );
  NAND U38567 ( .A(n29733), .B(n29734), .Z(N62741) );
  NAND U38568 ( .A(n29735), .B(n29736), .Z(n29734) );
  NANDN U38569 ( .A(n29737), .B(n29738), .Z(n29736) );
  NANDN U38570 ( .A(n29738), .B(n29737), .Z(n29733) );
  XOR U38571 ( .A(n29737), .B(n29739), .Z(N62740) );
  XNOR U38572 ( .A(n29735), .B(n29738), .Z(n29739) );
  NAND U38573 ( .A(n29740), .B(n29741), .Z(n29738) );
  NAND U38574 ( .A(n29742), .B(n29743), .Z(n29741) );
  NANDN U38575 ( .A(n29744), .B(n29745), .Z(n29743) );
  NANDN U38576 ( .A(n29745), .B(n29744), .Z(n29740) );
  AND U38577 ( .A(n29746), .B(n29747), .Z(n29735) );
  NAND U38578 ( .A(n29748), .B(n29749), .Z(n29747) );
  NANDN U38579 ( .A(n29750), .B(n29751), .Z(n29749) );
  NANDN U38580 ( .A(n29751), .B(n29750), .Z(n29746) );
  IV U38581 ( .A(n29752), .Z(n29751) );
  AND U38582 ( .A(n29753), .B(n29754), .Z(n29737) );
  NAND U38583 ( .A(n29755), .B(n29756), .Z(n29754) );
  NANDN U38584 ( .A(n29757), .B(n29758), .Z(n29756) );
  NANDN U38585 ( .A(n29758), .B(n29757), .Z(n29753) );
  XOR U38586 ( .A(n29750), .B(n29759), .Z(N62739) );
  XNOR U38587 ( .A(n29748), .B(n29752), .Z(n29759) );
  XOR U38588 ( .A(n29745), .B(n29760), .Z(n29752) );
  XNOR U38589 ( .A(n29742), .B(n29744), .Z(n29760) );
  AND U38590 ( .A(n29761), .B(n29762), .Z(n29744) );
  NANDN U38591 ( .A(n29763), .B(n29764), .Z(n29762) );
  OR U38592 ( .A(n29765), .B(n29766), .Z(n29764) );
  IV U38593 ( .A(n29767), .Z(n29766) );
  NANDN U38594 ( .A(n29767), .B(n29765), .Z(n29761) );
  AND U38595 ( .A(n29768), .B(n29769), .Z(n29742) );
  NAND U38596 ( .A(n29770), .B(n29771), .Z(n29769) );
  NANDN U38597 ( .A(n29772), .B(n29773), .Z(n29771) );
  NANDN U38598 ( .A(n29773), .B(n29772), .Z(n29768) );
  IV U38599 ( .A(n29774), .Z(n29773) );
  NAND U38600 ( .A(n29775), .B(n29776), .Z(n29745) );
  NANDN U38601 ( .A(n29777), .B(n29778), .Z(n29776) );
  NANDN U38602 ( .A(n29779), .B(n29780), .Z(n29778) );
  NANDN U38603 ( .A(n29780), .B(n29779), .Z(n29775) );
  IV U38604 ( .A(n29781), .Z(n29779) );
  AND U38605 ( .A(n29782), .B(n29783), .Z(n29748) );
  NAND U38606 ( .A(n29784), .B(n29785), .Z(n29783) );
  NANDN U38607 ( .A(n29786), .B(n29787), .Z(n29785) );
  NANDN U38608 ( .A(n29787), .B(n29786), .Z(n29782) );
  XOR U38609 ( .A(n29758), .B(n29788), .Z(n29750) );
  XNOR U38610 ( .A(n29755), .B(n29757), .Z(n29788) );
  AND U38611 ( .A(n29789), .B(n29790), .Z(n29757) );
  NANDN U38612 ( .A(n29791), .B(n29792), .Z(n29790) );
  OR U38613 ( .A(n29793), .B(n29794), .Z(n29792) );
  IV U38614 ( .A(n29795), .Z(n29794) );
  NANDN U38615 ( .A(n29795), .B(n29793), .Z(n29789) );
  AND U38616 ( .A(n29796), .B(n29797), .Z(n29755) );
  NAND U38617 ( .A(n29798), .B(n29799), .Z(n29797) );
  NANDN U38618 ( .A(n29800), .B(n29801), .Z(n29799) );
  NANDN U38619 ( .A(n29801), .B(n29800), .Z(n29796) );
  IV U38620 ( .A(n29802), .Z(n29801) );
  NAND U38621 ( .A(n29803), .B(n29804), .Z(n29758) );
  NANDN U38622 ( .A(n29805), .B(n29806), .Z(n29804) );
  NANDN U38623 ( .A(n29807), .B(n29808), .Z(n29806) );
  NANDN U38624 ( .A(n29808), .B(n29807), .Z(n29803) );
  IV U38625 ( .A(n29809), .Z(n29807) );
  XOR U38626 ( .A(n29784), .B(n29810), .Z(N62738) );
  XNOR U38627 ( .A(n29787), .B(n29786), .Z(n29810) );
  XNOR U38628 ( .A(n29798), .B(n29811), .Z(n29786) );
  XNOR U38629 ( .A(n29802), .B(n29800), .Z(n29811) );
  XOR U38630 ( .A(n29808), .B(n29812), .Z(n29800) );
  XNOR U38631 ( .A(n29805), .B(n29809), .Z(n29812) );
  AND U38632 ( .A(n29813), .B(n29814), .Z(n29809) );
  NAND U38633 ( .A(n29815), .B(n29816), .Z(n29814) );
  NAND U38634 ( .A(n29817), .B(n29818), .Z(n29813) );
  AND U38635 ( .A(n29819), .B(n29820), .Z(n29805) );
  NAND U38636 ( .A(n29821), .B(n29822), .Z(n29820) );
  NAND U38637 ( .A(n29823), .B(n29824), .Z(n29819) );
  NANDN U38638 ( .A(n29825), .B(n29826), .Z(n29808) );
  ANDN U38639 ( .B(n29827), .A(n29828), .Z(n29802) );
  XNOR U38640 ( .A(n29793), .B(n29829), .Z(n29798) );
  XNOR U38641 ( .A(n29791), .B(n29795), .Z(n29829) );
  AND U38642 ( .A(n29830), .B(n29831), .Z(n29795) );
  NAND U38643 ( .A(n29832), .B(n29833), .Z(n29831) );
  NAND U38644 ( .A(n29834), .B(n29835), .Z(n29830) );
  AND U38645 ( .A(n29836), .B(n29837), .Z(n29791) );
  NAND U38646 ( .A(n29838), .B(n29839), .Z(n29837) );
  NAND U38647 ( .A(n29840), .B(n29841), .Z(n29836) );
  AND U38648 ( .A(n29842), .B(n29843), .Z(n29793) );
  NAND U38649 ( .A(n29844), .B(n29845), .Z(n29787) );
  XNOR U38650 ( .A(n29770), .B(n29846), .Z(n29784) );
  XNOR U38651 ( .A(n29774), .B(n29772), .Z(n29846) );
  XOR U38652 ( .A(n29780), .B(n29847), .Z(n29772) );
  XNOR U38653 ( .A(n29777), .B(n29781), .Z(n29847) );
  AND U38654 ( .A(n29848), .B(n29849), .Z(n29781) );
  NAND U38655 ( .A(n29850), .B(n29851), .Z(n29849) );
  NAND U38656 ( .A(n29852), .B(n29853), .Z(n29848) );
  AND U38657 ( .A(n29854), .B(n29855), .Z(n29777) );
  NAND U38658 ( .A(n29856), .B(n29857), .Z(n29855) );
  NAND U38659 ( .A(n29858), .B(n29859), .Z(n29854) );
  NANDN U38660 ( .A(n29860), .B(n29861), .Z(n29780) );
  ANDN U38661 ( .B(n29862), .A(n29863), .Z(n29774) );
  XNOR U38662 ( .A(n29765), .B(n29864), .Z(n29770) );
  XNOR U38663 ( .A(n29763), .B(n29767), .Z(n29864) );
  AND U38664 ( .A(n29865), .B(n29866), .Z(n29767) );
  NAND U38665 ( .A(n29867), .B(n29868), .Z(n29866) );
  NAND U38666 ( .A(n29869), .B(n29870), .Z(n29865) );
  AND U38667 ( .A(n29871), .B(n29872), .Z(n29763) );
  NAND U38668 ( .A(n29873), .B(n29874), .Z(n29872) );
  NAND U38669 ( .A(n29875), .B(n29876), .Z(n29871) );
  AND U38670 ( .A(n29877), .B(n29878), .Z(n29765) );
  XOR U38671 ( .A(n29845), .B(n29844), .Z(N62737) );
  XNOR U38672 ( .A(n29862), .B(n29863), .Z(n29844) );
  XNOR U38673 ( .A(n29877), .B(n29878), .Z(n29863) );
  XOR U38674 ( .A(n29874), .B(n29873), .Z(n29878) );
  XOR U38675 ( .A(y[3972]), .B(x[3972]), .Z(n29873) );
  XOR U38676 ( .A(n29876), .B(n29875), .Z(n29874) );
  XOR U38677 ( .A(y[3974]), .B(x[3974]), .Z(n29875) );
  XOR U38678 ( .A(y[3973]), .B(x[3973]), .Z(n29876) );
  XOR U38679 ( .A(n29868), .B(n29867), .Z(n29877) );
  XOR U38680 ( .A(n29870), .B(n29869), .Z(n29867) );
  XOR U38681 ( .A(y[3971]), .B(x[3971]), .Z(n29869) );
  XOR U38682 ( .A(y[3970]), .B(x[3970]), .Z(n29870) );
  XOR U38683 ( .A(y[3969]), .B(x[3969]), .Z(n29868) );
  XNOR U38684 ( .A(n29861), .B(n29860), .Z(n29862) );
  XNOR U38685 ( .A(n29857), .B(n29856), .Z(n29860) );
  XOR U38686 ( .A(n29859), .B(n29858), .Z(n29856) );
  XOR U38687 ( .A(y[3968]), .B(x[3968]), .Z(n29858) );
  XOR U38688 ( .A(y[3967]), .B(x[3967]), .Z(n29859) );
  XOR U38689 ( .A(y[3966]), .B(x[3966]), .Z(n29857) );
  XOR U38690 ( .A(n29851), .B(n29850), .Z(n29861) );
  XOR U38691 ( .A(n29853), .B(n29852), .Z(n29850) );
  XOR U38692 ( .A(y[3965]), .B(x[3965]), .Z(n29852) );
  XOR U38693 ( .A(y[3964]), .B(x[3964]), .Z(n29853) );
  XOR U38694 ( .A(y[3963]), .B(x[3963]), .Z(n29851) );
  XNOR U38695 ( .A(n29827), .B(n29828), .Z(n29845) );
  XNOR U38696 ( .A(n29842), .B(n29843), .Z(n29828) );
  XOR U38697 ( .A(n29839), .B(n29838), .Z(n29843) );
  XOR U38698 ( .A(y[3960]), .B(x[3960]), .Z(n29838) );
  XOR U38699 ( .A(n29841), .B(n29840), .Z(n29839) );
  XOR U38700 ( .A(y[3962]), .B(x[3962]), .Z(n29840) );
  XOR U38701 ( .A(y[3961]), .B(x[3961]), .Z(n29841) );
  XOR U38702 ( .A(n29833), .B(n29832), .Z(n29842) );
  XOR U38703 ( .A(n29835), .B(n29834), .Z(n29832) );
  XOR U38704 ( .A(y[3959]), .B(x[3959]), .Z(n29834) );
  XOR U38705 ( .A(y[3958]), .B(x[3958]), .Z(n29835) );
  XOR U38706 ( .A(y[3957]), .B(x[3957]), .Z(n29833) );
  XNOR U38707 ( .A(n29826), .B(n29825), .Z(n29827) );
  XNOR U38708 ( .A(n29822), .B(n29821), .Z(n29825) );
  XOR U38709 ( .A(n29824), .B(n29823), .Z(n29821) );
  XOR U38710 ( .A(y[3956]), .B(x[3956]), .Z(n29823) );
  XOR U38711 ( .A(y[3955]), .B(x[3955]), .Z(n29824) );
  XOR U38712 ( .A(y[3954]), .B(x[3954]), .Z(n29822) );
  XOR U38713 ( .A(n29816), .B(n29815), .Z(n29826) );
  XOR U38714 ( .A(n29818), .B(n29817), .Z(n29815) );
  XOR U38715 ( .A(y[3953]), .B(x[3953]), .Z(n29817) );
  XOR U38716 ( .A(y[3952]), .B(x[3952]), .Z(n29818) );
  XOR U38717 ( .A(y[3951]), .B(x[3951]), .Z(n29816) );
  NAND U38718 ( .A(n29879), .B(n29880), .Z(N62728) );
  NAND U38719 ( .A(n29881), .B(n29882), .Z(n29880) );
  NANDN U38720 ( .A(n29883), .B(n29884), .Z(n29882) );
  NANDN U38721 ( .A(n29884), .B(n29883), .Z(n29879) );
  XOR U38722 ( .A(n29883), .B(n29885), .Z(N62727) );
  XNOR U38723 ( .A(n29881), .B(n29884), .Z(n29885) );
  NAND U38724 ( .A(n29886), .B(n29887), .Z(n29884) );
  NAND U38725 ( .A(n29888), .B(n29889), .Z(n29887) );
  NANDN U38726 ( .A(n29890), .B(n29891), .Z(n29889) );
  NANDN U38727 ( .A(n29891), .B(n29890), .Z(n29886) );
  AND U38728 ( .A(n29892), .B(n29893), .Z(n29881) );
  NAND U38729 ( .A(n29894), .B(n29895), .Z(n29893) );
  NANDN U38730 ( .A(n29896), .B(n29897), .Z(n29895) );
  NANDN U38731 ( .A(n29897), .B(n29896), .Z(n29892) );
  IV U38732 ( .A(n29898), .Z(n29897) );
  AND U38733 ( .A(n29899), .B(n29900), .Z(n29883) );
  NAND U38734 ( .A(n29901), .B(n29902), .Z(n29900) );
  NANDN U38735 ( .A(n29903), .B(n29904), .Z(n29902) );
  NANDN U38736 ( .A(n29904), .B(n29903), .Z(n29899) );
  XOR U38737 ( .A(n29896), .B(n29905), .Z(N62726) );
  XNOR U38738 ( .A(n29894), .B(n29898), .Z(n29905) );
  XOR U38739 ( .A(n29891), .B(n29906), .Z(n29898) );
  XNOR U38740 ( .A(n29888), .B(n29890), .Z(n29906) );
  AND U38741 ( .A(n29907), .B(n29908), .Z(n29890) );
  NANDN U38742 ( .A(n29909), .B(n29910), .Z(n29908) );
  OR U38743 ( .A(n29911), .B(n29912), .Z(n29910) );
  IV U38744 ( .A(n29913), .Z(n29912) );
  NANDN U38745 ( .A(n29913), .B(n29911), .Z(n29907) );
  AND U38746 ( .A(n29914), .B(n29915), .Z(n29888) );
  NAND U38747 ( .A(n29916), .B(n29917), .Z(n29915) );
  NANDN U38748 ( .A(n29918), .B(n29919), .Z(n29917) );
  NANDN U38749 ( .A(n29919), .B(n29918), .Z(n29914) );
  IV U38750 ( .A(n29920), .Z(n29919) );
  NAND U38751 ( .A(n29921), .B(n29922), .Z(n29891) );
  NANDN U38752 ( .A(n29923), .B(n29924), .Z(n29922) );
  NANDN U38753 ( .A(n29925), .B(n29926), .Z(n29924) );
  NANDN U38754 ( .A(n29926), .B(n29925), .Z(n29921) );
  IV U38755 ( .A(n29927), .Z(n29925) );
  AND U38756 ( .A(n29928), .B(n29929), .Z(n29894) );
  NAND U38757 ( .A(n29930), .B(n29931), .Z(n29929) );
  NANDN U38758 ( .A(n29932), .B(n29933), .Z(n29931) );
  NANDN U38759 ( .A(n29933), .B(n29932), .Z(n29928) );
  XOR U38760 ( .A(n29904), .B(n29934), .Z(n29896) );
  XNOR U38761 ( .A(n29901), .B(n29903), .Z(n29934) );
  AND U38762 ( .A(n29935), .B(n29936), .Z(n29903) );
  NANDN U38763 ( .A(n29937), .B(n29938), .Z(n29936) );
  OR U38764 ( .A(n29939), .B(n29940), .Z(n29938) );
  IV U38765 ( .A(n29941), .Z(n29940) );
  NANDN U38766 ( .A(n29941), .B(n29939), .Z(n29935) );
  AND U38767 ( .A(n29942), .B(n29943), .Z(n29901) );
  NAND U38768 ( .A(n29944), .B(n29945), .Z(n29943) );
  NANDN U38769 ( .A(n29946), .B(n29947), .Z(n29945) );
  NANDN U38770 ( .A(n29947), .B(n29946), .Z(n29942) );
  IV U38771 ( .A(n29948), .Z(n29947) );
  NAND U38772 ( .A(n29949), .B(n29950), .Z(n29904) );
  NANDN U38773 ( .A(n29951), .B(n29952), .Z(n29950) );
  NANDN U38774 ( .A(n29953), .B(n29954), .Z(n29952) );
  NANDN U38775 ( .A(n29954), .B(n29953), .Z(n29949) );
  IV U38776 ( .A(n29955), .Z(n29953) );
  XOR U38777 ( .A(n29930), .B(n29956), .Z(N62725) );
  XNOR U38778 ( .A(n29933), .B(n29932), .Z(n29956) );
  XNOR U38779 ( .A(n29944), .B(n29957), .Z(n29932) );
  XNOR U38780 ( .A(n29948), .B(n29946), .Z(n29957) );
  XOR U38781 ( .A(n29954), .B(n29958), .Z(n29946) );
  XNOR U38782 ( .A(n29951), .B(n29955), .Z(n29958) );
  AND U38783 ( .A(n29959), .B(n29960), .Z(n29955) );
  NAND U38784 ( .A(n29961), .B(n29962), .Z(n29960) );
  NAND U38785 ( .A(n29963), .B(n29964), .Z(n29959) );
  AND U38786 ( .A(n29965), .B(n29966), .Z(n29951) );
  NAND U38787 ( .A(n29967), .B(n29968), .Z(n29966) );
  NAND U38788 ( .A(n29969), .B(n29970), .Z(n29965) );
  NANDN U38789 ( .A(n29971), .B(n29972), .Z(n29954) );
  ANDN U38790 ( .B(n29973), .A(n29974), .Z(n29948) );
  XNOR U38791 ( .A(n29939), .B(n29975), .Z(n29944) );
  XNOR U38792 ( .A(n29937), .B(n29941), .Z(n29975) );
  AND U38793 ( .A(n29976), .B(n29977), .Z(n29941) );
  NAND U38794 ( .A(n29978), .B(n29979), .Z(n29977) );
  NAND U38795 ( .A(n29980), .B(n29981), .Z(n29976) );
  AND U38796 ( .A(n29982), .B(n29983), .Z(n29937) );
  NAND U38797 ( .A(n29984), .B(n29985), .Z(n29983) );
  NAND U38798 ( .A(n29986), .B(n29987), .Z(n29982) );
  AND U38799 ( .A(n29988), .B(n29989), .Z(n29939) );
  NAND U38800 ( .A(n29990), .B(n29991), .Z(n29933) );
  XNOR U38801 ( .A(n29916), .B(n29992), .Z(n29930) );
  XNOR U38802 ( .A(n29920), .B(n29918), .Z(n29992) );
  XOR U38803 ( .A(n29926), .B(n29993), .Z(n29918) );
  XNOR U38804 ( .A(n29923), .B(n29927), .Z(n29993) );
  AND U38805 ( .A(n29994), .B(n29995), .Z(n29927) );
  NAND U38806 ( .A(n29996), .B(n29997), .Z(n29995) );
  NAND U38807 ( .A(n29998), .B(n29999), .Z(n29994) );
  AND U38808 ( .A(n30000), .B(n30001), .Z(n29923) );
  NAND U38809 ( .A(n30002), .B(n30003), .Z(n30001) );
  NAND U38810 ( .A(n30004), .B(n30005), .Z(n30000) );
  NANDN U38811 ( .A(n30006), .B(n30007), .Z(n29926) );
  ANDN U38812 ( .B(n30008), .A(n30009), .Z(n29920) );
  XNOR U38813 ( .A(n29911), .B(n30010), .Z(n29916) );
  XNOR U38814 ( .A(n29909), .B(n29913), .Z(n30010) );
  AND U38815 ( .A(n30011), .B(n30012), .Z(n29913) );
  NAND U38816 ( .A(n30013), .B(n30014), .Z(n30012) );
  NAND U38817 ( .A(n30015), .B(n30016), .Z(n30011) );
  AND U38818 ( .A(n30017), .B(n30018), .Z(n29909) );
  NAND U38819 ( .A(n30019), .B(n30020), .Z(n30018) );
  NAND U38820 ( .A(n30021), .B(n30022), .Z(n30017) );
  AND U38821 ( .A(n30023), .B(n30024), .Z(n29911) );
  XOR U38822 ( .A(n29991), .B(n29990), .Z(N62724) );
  XNOR U38823 ( .A(n30008), .B(n30009), .Z(n29990) );
  XNOR U38824 ( .A(n30023), .B(n30024), .Z(n30009) );
  XOR U38825 ( .A(n30020), .B(n30019), .Z(n30024) );
  XOR U38826 ( .A(y[3948]), .B(x[3948]), .Z(n30019) );
  XOR U38827 ( .A(n30022), .B(n30021), .Z(n30020) );
  XOR U38828 ( .A(y[3950]), .B(x[3950]), .Z(n30021) );
  XOR U38829 ( .A(y[3949]), .B(x[3949]), .Z(n30022) );
  XOR U38830 ( .A(n30014), .B(n30013), .Z(n30023) );
  XOR U38831 ( .A(n30016), .B(n30015), .Z(n30013) );
  XOR U38832 ( .A(y[3947]), .B(x[3947]), .Z(n30015) );
  XOR U38833 ( .A(y[3946]), .B(x[3946]), .Z(n30016) );
  XOR U38834 ( .A(y[3945]), .B(x[3945]), .Z(n30014) );
  XNOR U38835 ( .A(n30007), .B(n30006), .Z(n30008) );
  XNOR U38836 ( .A(n30003), .B(n30002), .Z(n30006) );
  XOR U38837 ( .A(n30005), .B(n30004), .Z(n30002) );
  XOR U38838 ( .A(y[3944]), .B(x[3944]), .Z(n30004) );
  XOR U38839 ( .A(y[3943]), .B(x[3943]), .Z(n30005) );
  XOR U38840 ( .A(y[3942]), .B(x[3942]), .Z(n30003) );
  XOR U38841 ( .A(n29997), .B(n29996), .Z(n30007) );
  XOR U38842 ( .A(n29999), .B(n29998), .Z(n29996) );
  XOR U38843 ( .A(y[3941]), .B(x[3941]), .Z(n29998) );
  XOR U38844 ( .A(y[3940]), .B(x[3940]), .Z(n29999) );
  XOR U38845 ( .A(y[3939]), .B(x[3939]), .Z(n29997) );
  XNOR U38846 ( .A(n29973), .B(n29974), .Z(n29991) );
  XNOR U38847 ( .A(n29988), .B(n29989), .Z(n29974) );
  XOR U38848 ( .A(n29985), .B(n29984), .Z(n29989) );
  XOR U38849 ( .A(y[3936]), .B(x[3936]), .Z(n29984) );
  XOR U38850 ( .A(n29987), .B(n29986), .Z(n29985) );
  XOR U38851 ( .A(y[3938]), .B(x[3938]), .Z(n29986) );
  XOR U38852 ( .A(y[3937]), .B(x[3937]), .Z(n29987) );
  XOR U38853 ( .A(n29979), .B(n29978), .Z(n29988) );
  XOR U38854 ( .A(n29981), .B(n29980), .Z(n29978) );
  XOR U38855 ( .A(y[3935]), .B(x[3935]), .Z(n29980) );
  XOR U38856 ( .A(y[3934]), .B(x[3934]), .Z(n29981) );
  XOR U38857 ( .A(y[3933]), .B(x[3933]), .Z(n29979) );
  XNOR U38858 ( .A(n29972), .B(n29971), .Z(n29973) );
  XNOR U38859 ( .A(n29968), .B(n29967), .Z(n29971) );
  XOR U38860 ( .A(n29970), .B(n29969), .Z(n29967) );
  XOR U38861 ( .A(y[3932]), .B(x[3932]), .Z(n29969) );
  XOR U38862 ( .A(y[3931]), .B(x[3931]), .Z(n29970) );
  XOR U38863 ( .A(y[3930]), .B(x[3930]), .Z(n29968) );
  XOR U38864 ( .A(n29962), .B(n29961), .Z(n29972) );
  XOR U38865 ( .A(n29964), .B(n29963), .Z(n29961) );
  XOR U38866 ( .A(y[3929]), .B(x[3929]), .Z(n29963) );
  XOR U38867 ( .A(y[3928]), .B(x[3928]), .Z(n29964) );
  XOR U38868 ( .A(y[3927]), .B(x[3927]), .Z(n29962) );
  NAND U38869 ( .A(n30025), .B(n30026), .Z(N62715) );
  NAND U38870 ( .A(n30027), .B(n30028), .Z(n30026) );
  NANDN U38871 ( .A(n30029), .B(n30030), .Z(n30028) );
  NANDN U38872 ( .A(n30030), .B(n30029), .Z(n30025) );
  XOR U38873 ( .A(n30029), .B(n30031), .Z(N62714) );
  XNOR U38874 ( .A(n30027), .B(n30030), .Z(n30031) );
  NAND U38875 ( .A(n30032), .B(n30033), .Z(n30030) );
  NAND U38876 ( .A(n30034), .B(n30035), .Z(n30033) );
  NANDN U38877 ( .A(n30036), .B(n30037), .Z(n30035) );
  NANDN U38878 ( .A(n30037), .B(n30036), .Z(n30032) );
  AND U38879 ( .A(n30038), .B(n30039), .Z(n30027) );
  NAND U38880 ( .A(n30040), .B(n30041), .Z(n30039) );
  NANDN U38881 ( .A(n30042), .B(n30043), .Z(n30041) );
  NANDN U38882 ( .A(n30043), .B(n30042), .Z(n30038) );
  IV U38883 ( .A(n30044), .Z(n30043) );
  AND U38884 ( .A(n30045), .B(n30046), .Z(n30029) );
  NAND U38885 ( .A(n30047), .B(n30048), .Z(n30046) );
  NANDN U38886 ( .A(n30049), .B(n30050), .Z(n30048) );
  NANDN U38887 ( .A(n30050), .B(n30049), .Z(n30045) );
  XOR U38888 ( .A(n30042), .B(n30051), .Z(N62713) );
  XNOR U38889 ( .A(n30040), .B(n30044), .Z(n30051) );
  XOR U38890 ( .A(n30037), .B(n30052), .Z(n30044) );
  XNOR U38891 ( .A(n30034), .B(n30036), .Z(n30052) );
  AND U38892 ( .A(n30053), .B(n30054), .Z(n30036) );
  NANDN U38893 ( .A(n30055), .B(n30056), .Z(n30054) );
  OR U38894 ( .A(n30057), .B(n30058), .Z(n30056) );
  IV U38895 ( .A(n30059), .Z(n30058) );
  NANDN U38896 ( .A(n30059), .B(n30057), .Z(n30053) );
  AND U38897 ( .A(n30060), .B(n30061), .Z(n30034) );
  NAND U38898 ( .A(n30062), .B(n30063), .Z(n30061) );
  NANDN U38899 ( .A(n30064), .B(n30065), .Z(n30063) );
  NANDN U38900 ( .A(n30065), .B(n30064), .Z(n30060) );
  IV U38901 ( .A(n30066), .Z(n30065) );
  NAND U38902 ( .A(n30067), .B(n30068), .Z(n30037) );
  NANDN U38903 ( .A(n30069), .B(n30070), .Z(n30068) );
  NANDN U38904 ( .A(n30071), .B(n30072), .Z(n30070) );
  NANDN U38905 ( .A(n30072), .B(n30071), .Z(n30067) );
  IV U38906 ( .A(n30073), .Z(n30071) );
  AND U38907 ( .A(n30074), .B(n30075), .Z(n30040) );
  NAND U38908 ( .A(n30076), .B(n30077), .Z(n30075) );
  NANDN U38909 ( .A(n30078), .B(n30079), .Z(n30077) );
  NANDN U38910 ( .A(n30079), .B(n30078), .Z(n30074) );
  XOR U38911 ( .A(n30050), .B(n30080), .Z(n30042) );
  XNOR U38912 ( .A(n30047), .B(n30049), .Z(n30080) );
  AND U38913 ( .A(n30081), .B(n30082), .Z(n30049) );
  NANDN U38914 ( .A(n30083), .B(n30084), .Z(n30082) );
  OR U38915 ( .A(n30085), .B(n30086), .Z(n30084) );
  IV U38916 ( .A(n30087), .Z(n30086) );
  NANDN U38917 ( .A(n30087), .B(n30085), .Z(n30081) );
  AND U38918 ( .A(n30088), .B(n30089), .Z(n30047) );
  NAND U38919 ( .A(n30090), .B(n30091), .Z(n30089) );
  NANDN U38920 ( .A(n30092), .B(n30093), .Z(n30091) );
  NANDN U38921 ( .A(n30093), .B(n30092), .Z(n30088) );
  IV U38922 ( .A(n30094), .Z(n30093) );
  NAND U38923 ( .A(n30095), .B(n30096), .Z(n30050) );
  NANDN U38924 ( .A(n30097), .B(n30098), .Z(n30096) );
  NANDN U38925 ( .A(n30099), .B(n30100), .Z(n30098) );
  NANDN U38926 ( .A(n30100), .B(n30099), .Z(n30095) );
  IV U38927 ( .A(n30101), .Z(n30099) );
  XOR U38928 ( .A(n30076), .B(n30102), .Z(N62712) );
  XNOR U38929 ( .A(n30079), .B(n30078), .Z(n30102) );
  XNOR U38930 ( .A(n30090), .B(n30103), .Z(n30078) );
  XNOR U38931 ( .A(n30094), .B(n30092), .Z(n30103) );
  XOR U38932 ( .A(n30100), .B(n30104), .Z(n30092) );
  XNOR U38933 ( .A(n30097), .B(n30101), .Z(n30104) );
  AND U38934 ( .A(n30105), .B(n30106), .Z(n30101) );
  NAND U38935 ( .A(n30107), .B(n30108), .Z(n30106) );
  NAND U38936 ( .A(n30109), .B(n30110), .Z(n30105) );
  AND U38937 ( .A(n30111), .B(n30112), .Z(n30097) );
  NAND U38938 ( .A(n30113), .B(n30114), .Z(n30112) );
  NAND U38939 ( .A(n30115), .B(n30116), .Z(n30111) );
  NANDN U38940 ( .A(n30117), .B(n30118), .Z(n30100) );
  ANDN U38941 ( .B(n30119), .A(n30120), .Z(n30094) );
  XNOR U38942 ( .A(n30085), .B(n30121), .Z(n30090) );
  XNOR U38943 ( .A(n30083), .B(n30087), .Z(n30121) );
  AND U38944 ( .A(n30122), .B(n30123), .Z(n30087) );
  NAND U38945 ( .A(n30124), .B(n30125), .Z(n30123) );
  NAND U38946 ( .A(n30126), .B(n30127), .Z(n30122) );
  AND U38947 ( .A(n30128), .B(n30129), .Z(n30083) );
  NAND U38948 ( .A(n30130), .B(n30131), .Z(n30129) );
  NAND U38949 ( .A(n30132), .B(n30133), .Z(n30128) );
  AND U38950 ( .A(n30134), .B(n30135), .Z(n30085) );
  NAND U38951 ( .A(n30136), .B(n30137), .Z(n30079) );
  XNOR U38952 ( .A(n30062), .B(n30138), .Z(n30076) );
  XNOR U38953 ( .A(n30066), .B(n30064), .Z(n30138) );
  XOR U38954 ( .A(n30072), .B(n30139), .Z(n30064) );
  XNOR U38955 ( .A(n30069), .B(n30073), .Z(n30139) );
  AND U38956 ( .A(n30140), .B(n30141), .Z(n30073) );
  NAND U38957 ( .A(n30142), .B(n30143), .Z(n30141) );
  NAND U38958 ( .A(n30144), .B(n30145), .Z(n30140) );
  AND U38959 ( .A(n30146), .B(n30147), .Z(n30069) );
  NAND U38960 ( .A(n30148), .B(n30149), .Z(n30147) );
  NAND U38961 ( .A(n30150), .B(n30151), .Z(n30146) );
  NANDN U38962 ( .A(n30152), .B(n30153), .Z(n30072) );
  ANDN U38963 ( .B(n30154), .A(n30155), .Z(n30066) );
  XNOR U38964 ( .A(n30057), .B(n30156), .Z(n30062) );
  XNOR U38965 ( .A(n30055), .B(n30059), .Z(n30156) );
  AND U38966 ( .A(n30157), .B(n30158), .Z(n30059) );
  NAND U38967 ( .A(n30159), .B(n30160), .Z(n30158) );
  NAND U38968 ( .A(n30161), .B(n30162), .Z(n30157) );
  AND U38969 ( .A(n30163), .B(n30164), .Z(n30055) );
  NAND U38970 ( .A(n30165), .B(n30166), .Z(n30164) );
  NAND U38971 ( .A(n30167), .B(n30168), .Z(n30163) );
  AND U38972 ( .A(n30169), .B(n30170), .Z(n30057) );
  XOR U38973 ( .A(n30137), .B(n30136), .Z(N62711) );
  XNOR U38974 ( .A(n30154), .B(n30155), .Z(n30136) );
  XNOR U38975 ( .A(n30169), .B(n30170), .Z(n30155) );
  XOR U38976 ( .A(n30166), .B(n30165), .Z(n30170) );
  XOR U38977 ( .A(y[3924]), .B(x[3924]), .Z(n30165) );
  XOR U38978 ( .A(n30168), .B(n30167), .Z(n30166) );
  XOR U38979 ( .A(y[3926]), .B(x[3926]), .Z(n30167) );
  XOR U38980 ( .A(y[3925]), .B(x[3925]), .Z(n30168) );
  XOR U38981 ( .A(n30160), .B(n30159), .Z(n30169) );
  XOR U38982 ( .A(n30162), .B(n30161), .Z(n30159) );
  XOR U38983 ( .A(y[3923]), .B(x[3923]), .Z(n30161) );
  XOR U38984 ( .A(y[3922]), .B(x[3922]), .Z(n30162) );
  XOR U38985 ( .A(y[3921]), .B(x[3921]), .Z(n30160) );
  XNOR U38986 ( .A(n30153), .B(n30152), .Z(n30154) );
  XNOR U38987 ( .A(n30149), .B(n30148), .Z(n30152) );
  XOR U38988 ( .A(n30151), .B(n30150), .Z(n30148) );
  XOR U38989 ( .A(y[3920]), .B(x[3920]), .Z(n30150) );
  XOR U38990 ( .A(y[3919]), .B(x[3919]), .Z(n30151) );
  XOR U38991 ( .A(y[3918]), .B(x[3918]), .Z(n30149) );
  XOR U38992 ( .A(n30143), .B(n30142), .Z(n30153) );
  XOR U38993 ( .A(n30145), .B(n30144), .Z(n30142) );
  XOR U38994 ( .A(y[3917]), .B(x[3917]), .Z(n30144) );
  XOR U38995 ( .A(y[3916]), .B(x[3916]), .Z(n30145) );
  XOR U38996 ( .A(y[3915]), .B(x[3915]), .Z(n30143) );
  XNOR U38997 ( .A(n30119), .B(n30120), .Z(n30137) );
  XNOR U38998 ( .A(n30134), .B(n30135), .Z(n30120) );
  XOR U38999 ( .A(n30131), .B(n30130), .Z(n30135) );
  XOR U39000 ( .A(y[3912]), .B(x[3912]), .Z(n30130) );
  XOR U39001 ( .A(n30133), .B(n30132), .Z(n30131) );
  XOR U39002 ( .A(y[3914]), .B(x[3914]), .Z(n30132) );
  XOR U39003 ( .A(y[3913]), .B(x[3913]), .Z(n30133) );
  XOR U39004 ( .A(n30125), .B(n30124), .Z(n30134) );
  XOR U39005 ( .A(n30127), .B(n30126), .Z(n30124) );
  XOR U39006 ( .A(y[3911]), .B(x[3911]), .Z(n30126) );
  XOR U39007 ( .A(y[3910]), .B(x[3910]), .Z(n30127) );
  XOR U39008 ( .A(y[3909]), .B(x[3909]), .Z(n30125) );
  XNOR U39009 ( .A(n30118), .B(n30117), .Z(n30119) );
  XNOR U39010 ( .A(n30114), .B(n30113), .Z(n30117) );
  XOR U39011 ( .A(n30116), .B(n30115), .Z(n30113) );
  XOR U39012 ( .A(y[3908]), .B(x[3908]), .Z(n30115) );
  XOR U39013 ( .A(y[3907]), .B(x[3907]), .Z(n30116) );
  XOR U39014 ( .A(y[3906]), .B(x[3906]), .Z(n30114) );
  XOR U39015 ( .A(n30108), .B(n30107), .Z(n30118) );
  XOR U39016 ( .A(n30110), .B(n30109), .Z(n30107) );
  XOR U39017 ( .A(y[3905]), .B(x[3905]), .Z(n30109) );
  XOR U39018 ( .A(y[3904]), .B(x[3904]), .Z(n30110) );
  XOR U39019 ( .A(y[3903]), .B(x[3903]), .Z(n30108) );
  NAND U39020 ( .A(n30171), .B(n30172), .Z(N62702) );
  NAND U39021 ( .A(n30173), .B(n30174), .Z(n30172) );
  NANDN U39022 ( .A(n30175), .B(n30176), .Z(n30174) );
  NANDN U39023 ( .A(n30176), .B(n30175), .Z(n30171) );
  XOR U39024 ( .A(n30175), .B(n30177), .Z(N62701) );
  XNOR U39025 ( .A(n30173), .B(n30176), .Z(n30177) );
  NAND U39026 ( .A(n30178), .B(n30179), .Z(n30176) );
  NAND U39027 ( .A(n30180), .B(n30181), .Z(n30179) );
  NANDN U39028 ( .A(n30182), .B(n30183), .Z(n30181) );
  NANDN U39029 ( .A(n30183), .B(n30182), .Z(n30178) );
  AND U39030 ( .A(n30184), .B(n30185), .Z(n30173) );
  NAND U39031 ( .A(n30186), .B(n30187), .Z(n30185) );
  NANDN U39032 ( .A(n30188), .B(n30189), .Z(n30187) );
  NANDN U39033 ( .A(n30189), .B(n30188), .Z(n30184) );
  IV U39034 ( .A(n30190), .Z(n30189) );
  AND U39035 ( .A(n30191), .B(n30192), .Z(n30175) );
  NAND U39036 ( .A(n30193), .B(n30194), .Z(n30192) );
  NANDN U39037 ( .A(n30195), .B(n30196), .Z(n30194) );
  NANDN U39038 ( .A(n30196), .B(n30195), .Z(n30191) );
  XOR U39039 ( .A(n30188), .B(n30197), .Z(N62700) );
  XNOR U39040 ( .A(n30186), .B(n30190), .Z(n30197) );
  XOR U39041 ( .A(n30183), .B(n30198), .Z(n30190) );
  XNOR U39042 ( .A(n30180), .B(n30182), .Z(n30198) );
  AND U39043 ( .A(n30199), .B(n30200), .Z(n30182) );
  NANDN U39044 ( .A(n30201), .B(n30202), .Z(n30200) );
  OR U39045 ( .A(n30203), .B(n30204), .Z(n30202) );
  IV U39046 ( .A(n30205), .Z(n30204) );
  NANDN U39047 ( .A(n30205), .B(n30203), .Z(n30199) );
  AND U39048 ( .A(n30206), .B(n30207), .Z(n30180) );
  NAND U39049 ( .A(n30208), .B(n30209), .Z(n30207) );
  NANDN U39050 ( .A(n30210), .B(n30211), .Z(n30209) );
  NANDN U39051 ( .A(n30211), .B(n30210), .Z(n30206) );
  IV U39052 ( .A(n30212), .Z(n30211) );
  NAND U39053 ( .A(n30213), .B(n30214), .Z(n30183) );
  NANDN U39054 ( .A(n30215), .B(n30216), .Z(n30214) );
  NANDN U39055 ( .A(n30217), .B(n30218), .Z(n30216) );
  NANDN U39056 ( .A(n30218), .B(n30217), .Z(n30213) );
  IV U39057 ( .A(n30219), .Z(n30217) );
  AND U39058 ( .A(n30220), .B(n30221), .Z(n30186) );
  NAND U39059 ( .A(n30222), .B(n30223), .Z(n30221) );
  NANDN U39060 ( .A(n30224), .B(n30225), .Z(n30223) );
  NANDN U39061 ( .A(n30225), .B(n30224), .Z(n30220) );
  XOR U39062 ( .A(n30196), .B(n30226), .Z(n30188) );
  XNOR U39063 ( .A(n30193), .B(n30195), .Z(n30226) );
  AND U39064 ( .A(n30227), .B(n30228), .Z(n30195) );
  NANDN U39065 ( .A(n30229), .B(n30230), .Z(n30228) );
  OR U39066 ( .A(n30231), .B(n30232), .Z(n30230) );
  IV U39067 ( .A(n30233), .Z(n30232) );
  NANDN U39068 ( .A(n30233), .B(n30231), .Z(n30227) );
  AND U39069 ( .A(n30234), .B(n30235), .Z(n30193) );
  NAND U39070 ( .A(n30236), .B(n30237), .Z(n30235) );
  NANDN U39071 ( .A(n30238), .B(n30239), .Z(n30237) );
  NANDN U39072 ( .A(n30239), .B(n30238), .Z(n30234) );
  IV U39073 ( .A(n30240), .Z(n30239) );
  NAND U39074 ( .A(n30241), .B(n30242), .Z(n30196) );
  NANDN U39075 ( .A(n30243), .B(n30244), .Z(n30242) );
  NANDN U39076 ( .A(n30245), .B(n30246), .Z(n30244) );
  NANDN U39077 ( .A(n30246), .B(n30245), .Z(n30241) );
  IV U39078 ( .A(n30247), .Z(n30245) );
  XOR U39079 ( .A(n30222), .B(n30248), .Z(N62699) );
  XNOR U39080 ( .A(n30225), .B(n30224), .Z(n30248) );
  XNOR U39081 ( .A(n30236), .B(n30249), .Z(n30224) );
  XNOR U39082 ( .A(n30240), .B(n30238), .Z(n30249) );
  XOR U39083 ( .A(n30246), .B(n30250), .Z(n30238) );
  XNOR U39084 ( .A(n30243), .B(n30247), .Z(n30250) );
  AND U39085 ( .A(n30251), .B(n30252), .Z(n30247) );
  NAND U39086 ( .A(n30253), .B(n30254), .Z(n30252) );
  NAND U39087 ( .A(n30255), .B(n30256), .Z(n30251) );
  AND U39088 ( .A(n30257), .B(n30258), .Z(n30243) );
  NAND U39089 ( .A(n30259), .B(n30260), .Z(n30258) );
  NAND U39090 ( .A(n30261), .B(n30262), .Z(n30257) );
  NANDN U39091 ( .A(n30263), .B(n30264), .Z(n30246) );
  ANDN U39092 ( .B(n30265), .A(n30266), .Z(n30240) );
  XNOR U39093 ( .A(n30231), .B(n30267), .Z(n30236) );
  XNOR U39094 ( .A(n30229), .B(n30233), .Z(n30267) );
  AND U39095 ( .A(n30268), .B(n30269), .Z(n30233) );
  NAND U39096 ( .A(n30270), .B(n30271), .Z(n30269) );
  NAND U39097 ( .A(n30272), .B(n30273), .Z(n30268) );
  AND U39098 ( .A(n30274), .B(n30275), .Z(n30229) );
  NAND U39099 ( .A(n30276), .B(n30277), .Z(n30275) );
  NAND U39100 ( .A(n30278), .B(n30279), .Z(n30274) );
  AND U39101 ( .A(n30280), .B(n30281), .Z(n30231) );
  NAND U39102 ( .A(n30282), .B(n30283), .Z(n30225) );
  XNOR U39103 ( .A(n30208), .B(n30284), .Z(n30222) );
  XNOR U39104 ( .A(n30212), .B(n30210), .Z(n30284) );
  XOR U39105 ( .A(n30218), .B(n30285), .Z(n30210) );
  XNOR U39106 ( .A(n30215), .B(n30219), .Z(n30285) );
  AND U39107 ( .A(n30286), .B(n30287), .Z(n30219) );
  NAND U39108 ( .A(n30288), .B(n30289), .Z(n30287) );
  NAND U39109 ( .A(n30290), .B(n30291), .Z(n30286) );
  AND U39110 ( .A(n30292), .B(n30293), .Z(n30215) );
  NAND U39111 ( .A(n30294), .B(n30295), .Z(n30293) );
  NAND U39112 ( .A(n30296), .B(n30297), .Z(n30292) );
  NANDN U39113 ( .A(n30298), .B(n30299), .Z(n30218) );
  ANDN U39114 ( .B(n30300), .A(n30301), .Z(n30212) );
  XNOR U39115 ( .A(n30203), .B(n30302), .Z(n30208) );
  XNOR U39116 ( .A(n30201), .B(n30205), .Z(n30302) );
  AND U39117 ( .A(n30303), .B(n30304), .Z(n30205) );
  NAND U39118 ( .A(n30305), .B(n30306), .Z(n30304) );
  NAND U39119 ( .A(n30307), .B(n30308), .Z(n30303) );
  AND U39120 ( .A(n30309), .B(n30310), .Z(n30201) );
  NAND U39121 ( .A(n30311), .B(n30312), .Z(n30310) );
  NAND U39122 ( .A(n30313), .B(n30314), .Z(n30309) );
  AND U39123 ( .A(n30315), .B(n30316), .Z(n30203) );
  XOR U39124 ( .A(n30283), .B(n30282), .Z(N62698) );
  XNOR U39125 ( .A(n30300), .B(n30301), .Z(n30282) );
  XNOR U39126 ( .A(n30315), .B(n30316), .Z(n30301) );
  XOR U39127 ( .A(n30312), .B(n30311), .Z(n30316) );
  XOR U39128 ( .A(y[3900]), .B(x[3900]), .Z(n30311) );
  XOR U39129 ( .A(n30314), .B(n30313), .Z(n30312) );
  XOR U39130 ( .A(y[3902]), .B(x[3902]), .Z(n30313) );
  XOR U39131 ( .A(y[3901]), .B(x[3901]), .Z(n30314) );
  XOR U39132 ( .A(n30306), .B(n30305), .Z(n30315) );
  XOR U39133 ( .A(n30308), .B(n30307), .Z(n30305) );
  XOR U39134 ( .A(y[3899]), .B(x[3899]), .Z(n30307) );
  XOR U39135 ( .A(y[3898]), .B(x[3898]), .Z(n30308) );
  XOR U39136 ( .A(y[3897]), .B(x[3897]), .Z(n30306) );
  XNOR U39137 ( .A(n30299), .B(n30298), .Z(n30300) );
  XNOR U39138 ( .A(n30295), .B(n30294), .Z(n30298) );
  XOR U39139 ( .A(n30297), .B(n30296), .Z(n30294) );
  XOR U39140 ( .A(y[3896]), .B(x[3896]), .Z(n30296) );
  XOR U39141 ( .A(y[3895]), .B(x[3895]), .Z(n30297) );
  XOR U39142 ( .A(y[3894]), .B(x[3894]), .Z(n30295) );
  XOR U39143 ( .A(n30289), .B(n30288), .Z(n30299) );
  XOR U39144 ( .A(n30291), .B(n30290), .Z(n30288) );
  XOR U39145 ( .A(y[3893]), .B(x[3893]), .Z(n30290) );
  XOR U39146 ( .A(y[3892]), .B(x[3892]), .Z(n30291) );
  XOR U39147 ( .A(y[3891]), .B(x[3891]), .Z(n30289) );
  XNOR U39148 ( .A(n30265), .B(n30266), .Z(n30283) );
  XNOR U39149 ( .A(n30280), .B(n30281), .Z(n30266) );
  XOR U39150 ( .A(n30277), .B(n30276), .Z(n30281) );
  XOR U39151 ( .A(y[3888]), .B(x[3888]), .Z(n30276) );
  XOR U39152 ( .A(n30279), .B(n30278), .Z(n30277) );
  XOR U39153 ( .A(y[3890]), .B(x[3890]), .Z(n30278) );
  XOR U39154 ( .A(y[3889]), .B(x[3889]), .Z(n30279) );
  XOR U39155 ( .A(n30271), .B(n30270), .Z(n30280) );
  XOR U39156 ( .A(n30273), .B(n30272), .Z(n30270) );
  XOR U39157 ( .A(y[3887]), .B(x[3887]), .Z(n30272) );
  XOR U39158 ( .A(y[3886]), .B(x[3886]), .Z(n30273) );
  XOR U39159 ( .A(y[3885]), .B(x[3885]), .Z(n30271) );
  XNOR U39160 ( .A(n30264), .B(n30263), .Z(n30265) );
  XNOR U39161 ( .A(n30260), .B(n30259), .Z(n30263) );
  XOR U39162 ( .A(n30262), .B(n30261), .Z(n30259) );
  XOR U39163 ( .A(y[3884]), .B(x[3884]), .Z(n30261) );
  XOR U39164 ( .A(y[3883]), .B(x[3883]), .Z(n30262) );
  XOR U39165 ( .A(y[3882]), .B(x[3882]), .Z(n30260) );
  XOR U39166 ( .A(n30254), .B(n30253), .Z(n30264) );
  XOR U39167 ( .A(n30256), .B(n30255), .Z(n30253) );
  XOR U39168 ( .A(y[3881]), .B(x[3881]), .Z(n30255) );
  XOR U39169 ( .A(y[3880]), .B(x[3880]), .Z(n30256) );
  XOR U39170 ( .A(y[3879]), .B(x[3879]), .Z(n30254) );
  NAND U39171 ( .A(n30317), .B(n30318), .Z(N62689) );
  NAND U39172 ( .A(n30319), .B(n30320), .Z(n30318) );
  NANDN U39173 ( .A(n30321), .B(n30322), .Z(n30320) );
  NANDN U39174 ( .A(n30322), .B(n30321), .Z(n30317) );
  XOR U39175 ( .A(n30321), .B(n30323), .Z(N62688) );
  XNOR U39176 ( .A(n30319), .B(n30322), .Z(n30323) );
  NAND U39177 ( .A(n30324), .B(n30325), .Z(n30322) );
  NAND U39178 ( .A(n30326), .B(n30327), .Z(n30325) );
  NANDN U39179 ( .A(n30328), .B(n30329), .Z(n30327) );
  NANDN U39180 ( .A(n30329), .B(n30328), .Z(n30324) );
  AND U39181 ( .A(n30330), .B(n30331), .Z(n30319) );
  NAND U39182 ( .A(n30332), .B(n30333), .Z(n30331) );
  NANDN U39183 ( .A(n30334), .B(n30335), .Z(n30333) );
  NANDN U39184 ( .A(n30335), .B(n30334), .Z(n30330) );
  IV U39185 ( .A(n30336), .Z(n30335) );
  AND U39186 ( .A(n30337), .B(n30338), .Z(n30321) );
  NAND U39187 ( .A(n30339), .B(n30340), .Z(n30338) );
  NANDN U39188 ( .A(n30341), .B(n30342), .Z(n30340) );
  NANDN U39189 ( .A(n30342), .B(n30341), .Z(n30337) );
  XOR U39190 ( .A(n30334), .B(n30343), .Z(N62687) );
  XNOR U39191 ( .A(n30332), .B(n30336), .Z(n30343) );
  XOR U39192 ( .A(n30329), .B(n30344), .Z(n30336) );
  XNOR U39193 ( .A(n30326), .B(n30328), .Z(n30344) );
  AND U39194 ( .A(n30345), .B(n30346), .Z(n30328) );
  NANDN U39195 ( .A(n30347), .B(n30348), .Z(n30346) );
  OR U39196 ( .A(n30349), .B(n30350), .Z(n30348) );
  IV U39197 ( .A(n30351), .Z(n30350) );
  NANDN U39198 ( .A(n30351), .B(n30349), .Z(n30345) );
  AND U39199 ( .A(n30352), .B(n30353), .Z(n30326) );
  NAND U39200 ( .A(n30354), .B(n30355), .Z(n30353) );
  NANDN U39201 ( .A(n30356), .B(n30357), .Z(n30355) );
  NANDN U39202 ( .A(n30357), .B(n30356), .Z(n30352) );
  IV U39203 ( .A(n30358), .Z(n30357) );
  NAND U39204 ( .A(n30359), .B(n30360), .Z(n30329) );
  NANDN U39205 ( .A(n30361), .B(n30362), .Z(n30360) );
  NANDN U39206 ( .A(n30363), .B(n30364), .Z(n30362) );
  NANDN U39207 ( .A(n30364), .B(n30363), .Z(n30359) );
  IV U39208 ( .A(n30365), .Z(n30363) );
  AND U39209 ( .A(n30366), .B(n30367), .Z(n30332) );
  NAND U39210 ( .A(n30368), .B(n30369), .Z(n30367) );
  NANDN U39211 ( .A(n30370), .B(n30371), .Z(n30369) );
  NANDN U39212 ( .A(n30371), .B(n30370), .Z(n30366) );
  XOR U39213 ( .A(n30342), .B(n30372), .Z(n30334) );
  XNOR U39214 ( .A(n30339), .B(n30341), .Z(n30372) );
  AND U39215 ( .A(n30373), .B(n30374), .Z(n30341) );
  NANDN U39216 ( .A(n30375), .B(n30376), .Z(n30374) );
  OR U39217 ( .A(n30377), .B(n30378), .Z(n30376) );
  IV U39218 ( .A(n30379), .Z(n30378) );
  NANDN U39219 ( .A(n30379), .B(n30377), .Z(n30373) );
  AND U39220 ( .A(n30380), .B(n30381), .Z(n30339) );
  NAND U39221 ( .A(n30382), .B(n30383), .Z(n30381) );
  NANDN U39222 ( .A(n30384), .B(n30385), .Z(n30383) );
  NANDN U39223 ( .A(n30385), .B(n30384), .Z(n30380) );
  IV U39224 ( .A(n30386), .Z(n30385) );
  NAND U39225 ( .A(n30387), .B(n30388), .Z(n30342) );
  NANDN U39226 ( .A(n30389), .B(n30390), .Z(n30388) );
  NANDN U39227 ( .A(n30391), .B(n30392), .Z(n30390) );
  NANDN U39228 ( .A(n30392), .B(n30391), .Z(n30387) );
  IV U39229 ( .A(n30393), .Z(n30391) );
  XOR U39230 ( .A(n30368), .B(n30394), .Z(N62686) );
  XNOR U39231 ( .A(n30371), .B(n30370), .Z(n30394) );
  XNOR U39232 ( .A(n30382), .B(n30395), .Z(n30370) );
  XNOR U39233 ( .A(n30386), .B(n30384), .Z(n30395) );
  XOR U39234 ( .A(n30392), .B(n30396), .Z(n30384) );
  XNOR U39235 ( .A(n30389), .B(n30393), .Z(n30396) );
  AND U39236 ( .A(n30397), .B(n30398), .Z(n30393) );
  NAND U39237 ( .A(n30399), .B(n30400), .Z(n30398) );
  NAND U39238 ( .A(n30401), .B(n30402), .Z(n30397) );
  AND U39239 ( .A(n30403), .B(n30404), .Z(n30389) );
  NAND U39240 ( .A(n30405), .B(n30406), .Z(n30404) );
  NAND U39241 ( .A(n30407), .B(n30408), .Z(n30403) );
  NANDN U39242 ( .A(n30409), .B(n30410), .Z(n30392) );
  ANDN U39243 ( .B(n30411), .A(n30412), .Z(n30386) );
  XNOR U39244 ( .A(n30377), .B(n30413), .Z(n30382) );
  XNOR U39245 ( .A(n30375), .B(n30379), .Z(n30413) );
  AND U39246 ( .A(n30414), .B(n30415), .Z(n30379) );
  NAND U39247 ( .A(n30416), .B(n30417), .Z(n30415) );
  NAND U39248 ( .A(n30418), .B(n30419), .Z(n30414) );
  AND U39249 ( .A(n30420), .B(n30421), .Z(n30375) );
  NAND U39250 ( .A(n30422), .B(n30423), .Z(n30421) );
  NAND U39251 ( .A(n30424), .B(n30425), .Z(n30420) );
  AND U39252 ( .A(n30426), .B(n30427), .Z(n30377) );
  NAND U39253 ( .A(n30428), .B(n30429), .Z(n30371) );
  XNOR U39254 ( .A(n30354), .B(n30430), .Z(n30368) );
  XNOR U39255 ( .A(n30358), .B(n30356), .Z(n30430) );
  XOR U39256 ( .A(n30364), .B(n30431), .Z(n30356) );
  XNOR U39257 ( .A(n30361), .B(n30365), .Z(n30431) );
  AND U39258 ( .A(n30432), .B(n30433), .Z(n30365) );
  NAND U39259 ( .A(n30434), .B(n30435), .Z(n30433) );
  NAND U39260 ( .A(n30436), .B(n30437), .Z(n30432) );
  AND U39261 ( .A(n30438), .B(n30439), .Z(n30361) );
  NAND U39262 ( .A(n30440), .B(n30441), .Z(n30439) );
  NAND U39263 ( .A(n30442), .B(n30443), .Z(n30438) );
  NANDN U39264 ( .A(n30444), .B(n30445), .Z(n30364) );
  ANDN U39265 ( .B(n30446), .A(n30447), .Z(n30358) );
  XNOR U39266 ( .A(n30349), .B(n30448), .Z(n30354) );
  XNOR U39267 ( .A(n30347), .B(n30351), .Z(n30448) );
  AND U39268 ( .A(n30449), .B(n30450), .Z(n30351) );
  NAND U39269 ( .A(n30451), .B(n30452), .Z(n30450) );
  NAND U39270 ( .A(n30453), .B(n30454), .Z(n30449) );
  AND U39271 ( .A(n30455), .B(n30456), .Z(n30347) );
  NAND U39272 ( .A(n30457), .B(n30458), .Z(n30456) );
  NAND U39273 ( .A(n30459), .B(n30460), .Z(n30455) );
  AND U39274 ( .A(n30461), .B(n30462), .Z(n30349) );
  XOR U39275 ( .A(n30429), .B(n30428), .Z(N62685) );
  XNOR U39276 ( .A(n30446), .B(n30447), .Z(n30428) );
  XNOR U39277 ( .A(n30461), .B(n30462), .Z(n30447) );
  XOR U39278 ( .A(n30458), .B(n30457), .Z(n30462) );
  XOR U39279 ( .A(y[3876]), .B(x[3876]), .Z(n30457) );
  XOR U39280 ( .A(n30460), .B(n30459), .Z(n30458) );
  XOR U39281 ( .A(y[3878]), .B(x[3878]), .Z(n30459) );
  XOR U39282 ( .A(y[3877]), .B(x[3877]), .Z(n30460) );
  XOR U39283 ( .A(n30452), .B(n30451), .Z(n30461) );
  XOR U39284 ( .A(n30454), .B(n30453), .Z(n30451) );
  XOR U39285 ( .A(y[3875]), .B(x[3875]), .Z(n30453) );
  XOR U39286 ( .A(y[3874]), .B(x[3874]), .Z(n30454) );
  XOR U39287 ( .A(y[3873]), .B(x[3873]), .Z(n30452) );
  XNOR U39288 ( .A(n30445), .B(n30444), .Z(n30446) );
  XNOR U39289 ( .A(n30441), .B(n30440), .Z(n30444) );
  XOR U39290 ( .A(n30443), .B(n30442), .Z(n30440) );
  XOR U39291 ( .A(y[3872]), .B(x[3872]), .Z(n30442) );
  XOR U39292 ( .A(y[3871]), .B(x[3871]), .Z(n30443) );
  XOR U39293 ( .A(y[3870]), .B(x[3870]), .Z(n30441) );
  XOR U39294 ( .A(n30435), .B(n30434), .Z(n30445) );
  XOR U39295 ( .A(n30437), .B(n30436), .Z(n30434) );
  XOR U39296 ( .A(y[3869]), .B(x[3869]), .Z(n30436) );
  XOR U39297 ( .A(y[3868]), .B(x[3868]), .Z(n30437) );
  XOR U39298 ( .A(y[3867]), .B(x[3867]), .Z(n30435) );
  XNOR U39299 ( .A(n30411), .B(n30412), .Z(n30429) );
  XNOR U39300 ( .A(n30426), .B(n30427), .Z(n30412) );
  XOR U39301 ( .A(n30423), .B(n30422), .Z(n30427) );
  XOR U39302 ( .A(y[3864]), .B(x[3864]), .Z(n30422) );
  XOR U39303 ( .A(n30425), .B(n30424), .Z(n30423) );
  XOR U39304 ( .A(y[3866]), .B(x[3866]), .Z(n30424) );
  XOR U39305 ( .A(y[3865]), .B(x[3865]), .Z(n30425) );
  XOR U39306 ( .A(n30417), .B(n30416), .Z(n30426) );
  XOR U39307 ( .A(n30419), .B(n30418), .Z(n30416) );
  XOR U39308 ( .A(y[3863]), .B(x[3863]), .Z(n30418) );
  XOR U39309 ( .A(y[3862]), .B(x[3862]), .Z(n30419) );
  XOR U39310 ( .A(y[3861]), .B(x[3861]), .Z(n30417) );
  XNOR U39311 ( .A(n30410), .B(n30409), .Z(n30411) );
  XNOR U39312 ( .A(n30406), .B(n30405), .Z(n30409) );
  XOR U39313 ( .A(n30408), .B(n30407), .Z(n30405) );
  XOR U39314 ( .A(y[3860]), .B(x[3860]), .Z(n30407) );
  XOR U39315 ( .A(y[3859]), .B(x[3859]), .Z(n30408) );
  XOR U39316 ( .A(y[3858]), .B(x[3858]), .Z(n30406) );
  XOR U39317 ( .A(n30400), .B(n30399), .Z(n30410) );
  XOR U39318 ( .A(n30402), .B(n30401), .Z(n30399) );
  XOR U39319 ( .A(y[3857]), .B(x[3857]), .Z(n30401) );
  XOR U39320 ( .A(y[3856]), .B(x[3856]), .Z(n30402) );
  XOR U39321 ( .A(y[3855]), .B(x[3855]), .Z(n30400) );
  NAND U39322 ( .A(n30463), .B(n30464), .Z(N62676) );
  NAND U39323 ( .A(n30465), .B(n30466), .Z(n30464) );
  NANDN U39324 ( .A(n30467), .B(n30468), .Z(n30466) );
  NANDN U39325 ( .A(n30468), .B(n30467), .Z(n30463) );
  XOR U39326 ( .A(n30467), .B(n30469), .Z(N62675) );
  XNOR U39327 ( .A(n30465), .B(n30468), .Z(n30469) );
  NAND U39328 ( .A(n30470), .B(n30471), .Z(n30468) );
  NAND U39329 ( .A(n30472), .B(n30473), .Z(n30471) );
  NANDN U39330 ( .A(n30474), .B(n30475), .Z(n30473) );
  NANDN U39331 ( .A(n30475), .B(n30474), .Z(n30470) );
  AND U39332 ( .A(n30476), .B(n30477), .Z(n30465) );
  NAND U39333 ( .A(n30478), .B(n30479), .Z(n30477) );
  NANDN U39334 ( .A(n30480), .B(n30481), .Z(n30479) );
  NANDN U39335 ( .A(n30481), .B(n30480), .Z(n30476) );
  IV U39336 ( .A(n30482), .Z(n30481) );
  AND U39337 ( .A(n30483), .B(n30484), .Z(n30467) );
  NAND U39338 ( .A(n30485), .B(n30486), .Z(n30484) );
  NANDN U39339 ( .A(n30487), .B(n30488), .Z(n30486) );
  NANDN U39340 ( .A(n30488), .B(n30487), .Z(n30483) );
  XOR U39341 ( .A(n30480), .B(n30489), .Z(N62674) );
  XNOR U39342 ( .A(n30478), .B(n30482), .Z(n30489) );
  XOR U39343 ( .A(n30475), .B(n30490), .Z(n30482) );
  XNOR U39344 ( .A(n30472), .B(n30474), .Z(n30490) );
  AND U39345 ( .A(n30491), .B(n30492), .Z(n30474) );
  NANDN U39346 ( .A(n30493), .B(n30494), .Z(n30492) );
  OR U39347 ( .A(n30495), .B(n30496), .Z(n30494) );
  IV U39348 ( .A(n30497), .Z(n30496) );
  NANDN U39349 ( .A(n30497), .B(n30495), .Z(n30491) );
  AND U39350 ( .A(n30498), .B(n30499), .Z(n30472) );
  NAND U39351 ( .A(n30500), .B(n30501), .Z(n30499) );
  NANDN U39352 ( .A(n30502), .B(n30503), .Z(n30501) );
  NANDN U39353 ( .A(n30503), .B(n30502), .Z(n30498) );
  IV U39354 ( .A(n30504), .Z(n30503) );
  NAND U39355 ( .A(n30505), .B(n30506), .Z(n30475) );
  NANDN U39356 ( .A(n30507), .B(n30508), .Z(n30506) );
  NANDN U39357 ( .A(n30509), .B(n30510), .Z(n30508) );
  NANDN U39358 ( .A(n30510), .B(n30509), .Z(n30505) );
  IV U39359 ( .A(n30511), .Z(n30509) );
  AND U39360 ( .A(n30512), .B(n30513), .Z(n30478) );
  NAND U39361 ( .A(n30514), .B(n30515), .Z(n30513) );
  NANDN U39362 ( .A(n30516), .B(n30517), .Z(n30515) );
  NANDN U39363 ( .A(n30517), .B(n30516), .Z(n30512) );
  XOR U39364 ( .A(n30488), .B(n30518), .Z(n30480) );
  XNOR U39365 ( .A(n30485), .B(n30487), .Z(n30518) );
  AND U39366 ( .A(n30519), .B(n30520), .Z(n30487) );
  NANDN U39367 ( .A(n30521), .B(n30522), .Z(n30520) );
  OR U39368 ( .A(n30523), .B(n30524), .Z(n30522) );
  IV U39369 ( .A(n30525), .Z(n30524) );
  NANDN U39370 ( .A(n30525), .B(n30523), .Z(n30519) );
  AND U39371 ( .A(n30526), .B(n30527), .Z(n30485) );
  NAND U39372 ( .A(n30528), .B(n30529), .Z(n30527) );
  NANDN U39373 ( .A(n30530), .B(n30531), .Z(n30529) );
  NANDN U39374 ( .A(n30531), .B(n30530), .Z(n30526) );
  IV U39375 ( .A(n30532), .Z(n30531) );
  NAND U39376 ( .A(n30533), .B(n30534), .Z(n30488) );
  NANDN U39377 ( .A(n30535), .B(n30536), .Z(n30534) );
  NANDN U39378 ( .A(n30537), .B(n30538), .Z(n30536) );
  NANDN U39379 ( .A(n30538), .B(n30537), .Z(n30533) );
  IV U39380 ( .A(n30539), .Z(n30537) );
  XOR U39381 ( .A(n30514), .B(n30540), .Z(N62673) );
  XNOR U39382 ( .A(n30517), .B(n30516), .Z(n30540) );
  XNOR U39383 ( .A(n30528), .B(n30541), .Z(n30516) );
  XNOR U39384 ( .A(n30532), .B(n30530), .Z(n30541) );
  XOR U39385 ( .A(n30538), .B(n30542), .Z(n30530) );
  XNOR U39386 ( .A(n30535), .B(n30539), .Z(n30542) );
  AND U39387 ( .A(n30543), .B(n30544), .Z(n30539) );
  NAND U39388 ( .A(n30545), .B(n30546), .Z(n30544) );
  NAND U39389 ( .A(n30547), .B(n30548), .Z(n30543) );
  AND U39390 ( .A(n30549), .B(n30550), .Z(n30535) );
  NAND U39391 ( .A(n30551), .B(n30552), .Z(n30550) );
  NAND U39392 ( .A(n30553), .B(n30554), .Z(n30549) );
  NANDN U39393 ( .A(n30555), .B(n30556), .Z(n30538) );
  ANDN U39394 ( .B(n30557), .A(n30558), .Z(n30532) );
  XNOR U39395 ( .A(n30523), .B(n30559), .Z(n30528) );
  XNOR U39396 ( .A(n30521), .B(n30525), .Z(n30559) );
  AND U39397 ( .A(n30560), .B(n30561), .Z(n30525) );
  NAND U39398 ( .A(n30562), .B(n30563), .Z(n30561) );
  NAND U39399 ( .A(n30564), .B(n30565), .Z(n30560) );
  AND U39400 ( .A(n30566), .B(n30567), .Z(n30521) );
  NAND U39401 ( .A(n30568), .B(n30569), .Z(n30567) );
  NAND U39402 ( .A(n30570), .B(n30571), .Z(n30566) );
  AND U39403 ( .A(n30572), .B(n30573), .Z(n30523) );
  NAND U39404 ( .A(n30574), .B(n30575), .Z(n30517) );
  XNOR U39405 ( .A(n30500), .B(n30576), .Z(n30514) );
  XNOR U39406 ( .A(n30504), .B(n30502), .Z(n30576) );
  XOR U39407 ( .A(n30510), .B(n30577), .Z(n30502) );
  XNOR U39408 ( .A(n30507), .B(n30511), .Z(n30577) );
  AND U39409 ( .A(n30578), .B(n30579), .Z(n30511) );
  NAND U39410 ( .A(n30580), .B(n30581), .Z(n30579) );
  NAND U39411 ( .A(n30582), .B(n30583), .Z(n30578) );
  AND U39412 ( .A(n30584), .B(n30585), .Z(n30507) );
  NAND U39413 ( .A(n30586), .B(n30587), .Z(n30585) );
  NAND U39414 ( .A(n30588), .B(n30589), .Z(n30584) );
  NANDN U39415 ( .A(n30590), .B(n30591), .Z(n30510) );
  ANDN U39416 ( .B(n30592), .A(n30593), .Z(n30504) );
  XNOR U39417 ( .A(n30495), .B(n30594), .Z(n30500) );
  XNOR U39418 ( .A(n30493), .B(n30497), .Z(n30594) );
  AND U39419 ( .A(n30595), .B(n30596), .Z(n30497) );
  NAND U39420 ( .A(n30597), .B(n30598), .Z(n30596) );
  NAND U39421 ( .A(n30599), .B(n30600), .Z(n30595) );
  AND U39422 ( .A(n30601), .B(n30602), .Z(n30493) );
  NAND U39423 ( .A(n30603), .B(n30604), .Z(n30602) );
  NAND U39424 ( .A(n30605), .B(n30606), .Z(n30601) );
  AND U39425 ( .A(n30607), .B(n30608), .Z(n30495) );
  XOR U39426 ( .A(n30575), .B(n30574), .Z(N62672) );
  XNOR U39427 ( .A(n30592), .B(n30593), .Z(n30574) );
  XNOR U39428 ( .A(n30607), .B(n30608), .Z(n30593) );
  XOR U39429 ( .A(n30604), .B(n30603), .Z(n30608) );
  XOR U39430 ( .A(y[3852]), .B(x[3852]), .Z(n30603) );
  XOR U39431 ( .A(n30606), .B(n30605), .Z(n30604) );
  XOR U39432 ( .A(y[3854]), .B(x[3854]), .Z(n30605) );
  XOR U39433 ( .A(y[3853]), .B(x[3853]), .Z(n30606) );
  XOR U39434 ( .A(n30598), .B(n30597), .Z(n30607) );
  XOR U39435 ( .A(n30600), .B(n30599), .Z(n30597) );
  XOR U39436 ( .A(y[3851]), .B(x[3851]), .Z(n30599) );
  XOR U39437 ( .A(y[3850]), .B(x[3850]), .Z(n30600) );
  XOR U39438 ( .A(y[3849]), .B(x[3849]), .Z(n30598) );
  XNOR U39439 ( .A(n30591), .B(n30590), .Z(n30592) );
  XNOR U39440 ( .A(n30587), .B(n30586), .Z(n30590) );
  XOR U39441 ( .A(n30589), .B(n30588), .Z(n30586) );
  XOR U39442 ( .A(y[3848]), .B(x[3848]), .Z(n30588) );
  XOR U39443 ( .A(y[3847]), .B(x[3847]), .Z(n30589) );
  XOR U39444 ( .A(y[3846]), .B(x[3846]), .Z(n30587) );
  XOR U39445 ( .A(n30581), .B(n30580), .Z(n30591) );
  XOR U39446 ( .A(n30583), .B(n30582), .Z(n30580) );
  XOR U39447 ( .A(y[3845]), .B(x[3845]), .Z(n30582) );
  XOR U39448 ( .A(y[3844]), .B(x[3844]), .Z(n30583) );
  XOR U39449 ( .A(y[3843]), .B(x[3843]), .Z(n30581) );
  XNOR U39450 ( .A(n30557), .B(n30558), .Z(n30575) );
  XNOR U39451 ( .A(n30572), .B(n30573), .Z(n30558) );
  XOR U39452 ( .A(n30569), .B(n30568), .Z(n30573) );
  XOR U39453 ( .A(y[3840]), .B(x[3840]), .Z(n30568) );
  XOR U39454 ( .A(n30571), .B(n30570), .Z(n30569) );
  XOR U39455 ( .A(y[3842]), .B(x[3842]), .Z(n30570) );
  XOR U39456 ( .A(y[3841]), .B(x[3841]), .Z(n30571) );
  XOR U39457 ( .A(n30563), .B(n30562), .Z(n30572) );
  XOR U39458 ( .A(n30565), .B(n30564), .Z(n30562) );
  XOR U39459 ( .A(y[3839]), .B(x[3839]), .Z(n30564) );
  XOR U39460 ( .A(y[3838]), .B(x[3838]), .Z(n30565) );
  XOR U39461 ( .A(y[3837]), .B(x[3837]), .Z(n30563) );
  XNOR U39462 ( .A(n30556), .B(n30555), .Z(n30557) );
  XNOR U39463 ( .A(n30552), .B(n30551), .Z(n30555) );
  XOR U39464 ( .A(n30554), .B(n30553), .Z(n30551) );
  XOR U39465 ( .A(y[3836]), .B(x[3836]), .Z(n30553) );
  XOR U39466 ( .A(y[3835]), .B(x[3835]), .Z(n30554) );
  XOR U39467 ( .A(y[3834]), .B(x[3834]), .Z(n30552) );
  XOR U39468 ( .A(n30546), .B(n30545), .Z(n30556) );
  XOR U39469 ( .A(n30548), .B(n30547), .Z(n30545) );
  XOR U39470 ( .A(y[3833]), .B(x[3833]), .Z(n30547) );
  XOR U39471 ( .A(y[3832]), .B(x[3832]), .Z(n30548) );
  XOR U39472 ( .A(y[3831]), .B(x[3831]), .Z(n30546) );
  NAND U39473 ( .A(n30609), .B(n30610), .Z(N62663) );
  NAND U39474 ( .A(n30611), .B(n30612), .Z(n30610) );
  NANDN U39475 ( .A(n30613), .B(n30614), .Z(n30612) );
  NANDN U39476 ( .A(n30614), .B(n30613), .Z(n30609) );
  XOR U39477 ( .A(n30613), .B(n30615), .Z(N62662) );
  XNOR U39478 ( .A(n30611), .B(n30614), .Z(n30615) );
  NAND U39479 ( .A(n30616), .B(n30617), .Z(n30614) );
  NAND U39480 ( .A(n30618), .B(n30619), .Z(n30617) );
  NANDN U39481 ( .A(n30620), .B(n30621), .Z(n30619) );
  NANDN U39482 ( .A(n30621), .B(n30620), .Z(n30616) );
  AND U39483 ( .A(n30622), .B(n30623), .Z(n30611) );
  NAND U39484 ( .A(n30624), .B(n30625), .Z(n30623) );
  NANDN U39485 ( .A(n30626), .B(n30627), .Z(n30625) );
  NANDN U39486 ( .A(n30627), .B(n30626), .Z(n30622) );
  IV U39487 ( .A(n30628), .Z(n30627) );
  AND U39488 ( .A(n30629), .B(n30630), .Z(n30613) );
  NAND U39489 ( .A(n30631), .B(n30632), .Z(n30630) );
  NANDN U39490 ( .A(n30633), .B(n30634), .Z(n30632) );
  NANDN U39491 ( .A(n30634), .B(n30633), .Z(n30629) );
  XOR U39492 ( .A(n30626), .B(n30635), .Z(N62661) );
  XNOR U39493 ( .A(n30624), .B(n30628), .Z(n30635) );
  XOR U39494 ( .A(n30621), .B(n30636), .Z(n30628) );
  XNOR U39495 ( .A(n30618), .B(n30620), .Z(n30636) );
  AND U39496 ( .A(n30637), .B(n30638), .Z(n30620) );
  NANDN U39497 ( .A(n30639), .B(n30640), .Z(n30638) );
  OR U39498 ( .A(n30641), .B(n30642), .Z(n30640) );
  IV U39499 ( .A(n30643), .Z(n30642) );
  NANDN U39500 ( .A(n30643), .B(n30641), .Z(n30637) );
  AND U39501 ( .A(n30644), .B(n30645), .Z(n30618) );
  NAND U39502 ( .A(n30646), .B(n30647), .Z(n30645) );
  NANDN U39503 ( .A(n30648), .B(n30649), .Z(n30647) );
  NANDN U39504 ( .A(n30649), .B(n30648), .Z(n30644) );
  IV U39505 ( .A(n30650), .Z(n30649) );
  NAND U39506 ( .A(n30651), .B(n30652), .Z(n30621) );
  NANDN U39507 ( .A(n30653), .B(n30654), .Z(n30652) );
  NANDN U39508 ( .A(n30655), .B(n30656), .Z(n30654) );
  NANDN U39509 ( .A(n30656), .B(n30655), .Z(n30651) );
  IV U39510 ( .A(n30657), .Z(n30655) );
  AND U39511 ( .A(n30658), .B(n30659), .Z(n30624) );
  NAND U39512 ( .A(n30660), .B(n30661), .Z(n30659) );
  NANDN U39513 ( .A(n30662), .B(n30663), .Z(n30661) );
  NANDN U39514 ( .A(n30663), .B(n30662), .Z(n30658) );
  XOR U39515 ( .A(n30634), .B(n30664), .Z(n30626) );
  XNOR U39516 ( .A(n30631), .B(n30633), .Z(n30664) );
  AND U39517 ( .A(n30665), .B(n30666), .Z(n30633) );
  NANDN U39518 ( .A(n30667), .B(n30668), .Z(n30666) );
  OR U39519 ( .A(n30669), .B(n30670), .Z(n30668) );
  IV U39520 ( .A(n30671), .Z(n30670) );
  NANDN U39521 ( .A(n30671), .B(n30669), .Z(n30665) );
  AND U39522 ( .A(n30672), .B(n30673), .Z(n30631) );
  NAND U39523 ( .A(n30674), .B(n30675), .Z(n30673) );
  NANDN U39524 ( .A(n30676), .B(n30677), .Z(n30675) );
  NANDN U39525 ( .A(n30677), .B(n30676), .Z(n30672) );
  IV U39526 ( .A(n30678), .Z(n30677) );
  NAND U39527 ( .A(n30679), .B(n30680), .Z(n30634) );
  NANDN U39528 ( .A(n30681), .B(n30682), .Z(n30680) );
  NANDN U39529 ( .A(n30683), .B(n30684), .Z(n30682) );
  NANDN U39530 ( .A(n30684), .B(n30683), .Z(n30679) );
  IV U39531 ( .A(n30685), .Z(n30683) );
  XOR U39532 ( .A(n30660), .B(n30686), .Z(N62660) );
  XNOR U39533 ( .A(n30663), .B(n30662), .Z(n30686) );
  XNOR U39534 ( .A(n30674), .B(n30687), .Z(n30662) );
  XNOR U39535 ( .A(n30678), .B(n30676), .Z(n30687) );
  XOR U39536 ( .A(n30684), .B(n30688), .Z(n30676) );
  XNOR U39537 ( .A(n30681), .B(n30685), .Z(n30688) );
  AND U39538 ( .A(n30689), .B(n30690), .Z(n30685) );
  NAND U39539 ( .A(n30691), .B(n30692), .Z(n30690) );
  NAND U39540 ( .A(n30693), .B(n30694), .Z(n30689) );
  AND U39541 ( .A(n30695), .B(n30696), .Z(n30681) );
  NAND U39542 ( .A(n30697), .B(n30698), .Z(n30696) );
  NAND U39543 ( .A(n30699), .B(n30700), .Z(n30695) );
  NANDN U39544 ( .A(n30701), .B(n30702), .Z(n30684) );
  ANDN U39545 ( .B(n30703), .A(n30704), .Z(n30678) );
  XNOR U39546 ( .A(n30669), .B(n30705), .Z(n30674) );
  XNOR U39547 ( .A(n30667), .B(n30671), .Z(n30705) );
  AND U39548 ( .A(n30706), .B(n30707), .Z(n30671) );
  NAND U39549 ( .A(n30708), .B(n30709), .Z(n30707) );
  NAND U39550 ( .A(n30710), .B(n30711), .Z(n30706) );
  AND U39551 ( .A(n30712), .B(n30713), .Z(n30667) );
  NAND U39552 ( .A(n30714), .B(n30715), .Z(n30713) );
  NAND U39553 ( .A(n30716), .B(n30717), .Z(n30712) );
  AND U39554 ( .A(n30718), .B(n30719), .Z(n30669) );
  NAND U39555 ( .A(n30720), .B(n30721), .Z(n30663) );
  XNOR U39556 ( .A(n30646), .B(n30722), .Z(n30660) );
  XNOR U39557 ( .A(n30650), .B(n30648), .Z(n30722) );
  XOR U39558 ( .A(n30656), .B(n30723), .Z(n30648) );
  XNOR U39559 ( .A(n30653), .B(n30657), .Z(n30723) );
  AND U39560 ( .A(n30724), .B(n30725), .Z(n30657) );
  NAND U39561 ( .A(n30726), .B(n30727), .Z(n30725) );
  NAND U39562 ( .A(n30728), .B(n30729), .Z(n30724) );
  AND U39563 ( .A(n30730), .B(n30731), .Z(n30653) );
  NAND U39564 ( .A(n30732), .B(n30733), .Z(n30731) );
  NAND U39565 ( .A(n30734), .B(n30735), .Z(n30730) );
  NANDN U39566 ( .A(n30736), .B(n30737), .Z(n30656) );
  ANDN U39567 ( .B(n30738), .A(n30739), .Z(n30650) );
  XNOR U39568 ( .A(n30641), .B(n30740), .Z(n30646) );
  XNOR U39569 ( .A(n30639), .B(n30643), .Z(n30740) );
  AND U39570 ( .A(n30741), .B(n30742), .Z(n30643) );
  NAND U39571 ( .A(n30743), .B(n30744), .Z(n30742) );
  NAND U39572 ( .A(n30745), .B(n30746), .Z(n30741) );
  AND U39573 ( .A(n30747), .B(n30748), .Z(n30639) );
  NAND U39574 ( .A(n30749), .B(n30750), .Z(n30748) );
  NAND U39575 ( .A(n30751), .B(n30752), .Z(n30747) );
  AND U39576 ( .A(n30753), .B(n30754), .Z(n30641) );
  XOR U39577 ( .A(n30721), .B(n30720), .Z(N62659) );
  XNOR U39578 ( .A(n30738), .B(n30739), .Z(n30720) );
  XNOR U39579 ( .A(n30753), .B(n30754), .Z(n30739) );
  XOR U39580 ( .A(n30750), .B(n30749), .Z(n30754) );
  XOR U39581 ( .A(y[3828]), .B(x[3828]), .Z(n30749) );
  XOR U39582 ( .A(n30752), .B(n30751), .Z(n30750) );
  XOR U39583 ( .A(y[3830]), .B(x[3830]), .Z(n30751) );
  XOR U39584 ( .A(y[3829]), .B(x[3829]), .Z(n30752) );
  XOR U39585 ( .A(n30744), .B(n30743), .Z(n30753) );
  XOR U39586 ( .A(n30746), .B(n30745), .Z(n30743) );
  XOR U39587 ( .A(y[3827]), .B(x[3827]), .Z(n30745) );
  XOR U39588 ( .A(y[3826]), .B(x[3826]), .Z(n30746) );
  XOR U39589 ( .A(y[3825]), .B(x[3825]), .Z(n30744) );
  XNOR U39590 ( .A(n30737), .B(n30736), .Z(n30738) );
  XNOR U39591 ( .A(n30733), .B(n30732), .Z(n30736) );
  XOR U39592 ( .A(n30735), .B(n30734), .Z(n30732) );
  XOR U39593 ( .A(y[3824]), .B(x[3824]), .Z(n30734) );
  XOR U39594 ( .A(y[3823]), .B(x[3823]), .Z(n30735) );
  XOR U39595 ( .A(y[3822]), .B(x[3822]), .Z(n30733) );
  XOR U39596 ( .A(n30727), .B(n30726), .Z(n30737) );
  XOR U39597 ( .A(n30729), .B(n30728), .Z(n30726) );
  XOR U39598 ( .A(y[3821]), .B(x[3821]), .Z(n30728) );
  XOR U39599 ( .A(y[3820]), .B(x[3820]), .Z(n30729) );
  XOR U39600 ( .A(y[3819]), .B(x[3819]), .Z(n30727) );
  XNOR U39601 ( .A(n30703), .B(n30704), .Z(n30721) );
  XNOR U39602 ( .A(n30718), .B(n30719), .Z(n30704) );
  XOR U39603 ( .A(n30715), .B(n30714), .Z(n30719) );
  XOR U39604 ( .A(y[3816]), .B(x[3816]), .Z(n30714) );
  XOR U39605 ( .A(n30717), .B(n30716), .Z(n30715) );
  XOR U39606 ( .A(y[3818]), .B(x[3818]), .Z(n30716) );
  XOR U39607 ( .A(y[3817]), .B(x[3817]), .Z(n30717) );
  XOR U39608 ( .A(n30709), .B(n30708), .Z(n30718) );
  XOR U39609 ( .A(n30711), .B(n30710), .Z(n30708) );
  XOR U39610 ( .A(y[3815]), .B(x[3815]), .Z(n30710) );
  XOR U39611 ( .A(y[3814]), .B(x[3814]), .Z(n30711) );
  XOR U39612 ( .A(y[3813]), .B(x[3813]), .Z(n30709) );
  XNOR U39613 ( .A(n30702), .B(n30701), .Z(n30703) );
  XNOR U39614 ( .A(n30698), .B(n30697), .Z(n30701) );
  XOR U39615 ( .A(n30700), .B(n30699), .Z(n30697) );
  XOR U39616 ( .A(y[3812]), .B(x[3812]), .Z(n30699) );
  XOR U39617 ( .A(y[3811]), .B(x[3811]), .Z(n30700) );
  XOR U39618 ( .A(y[3810]), .B(x[3810]), .Z(n30698) );
  XOR U39619 ( .A(n30692), .B(n30691), .Z(n30702) );
  XOR U39620 ( .A(n30694), .B(n30693), .Z(n30691) );
  XOR U39621 ( .A(y[3809]), .B(x[3809]), .Z(n30693) );
  XOR U39622 ( .A(y[3808]), .B(x[3808]), .Z(n30694) );
  XOR U39623 ( .A(y[3807]), .B(x[3807]), .Z(n30692) );
  NAND U39624 ( .A(n30755), .B(n30756), .Z(N62650) );
  NAND U39625 ( .A(n30757), .B(n30758), .Z(n30756) );
  NANDN U39626 ( .A(n30759), .B(n30760), .Z(n30758) );
  NANDN U39627 ( .A(n30760), .B(n30759), .Z(n30755) );
  XOR U39628 ( .A(n30759), .B(n30761), .Z(N62649) );
  XNOR U39629 ( .A(n30757), .B(n30760), .Z(n30761) );
  NAND U39630 ( .A(n30762), .B(n30763), .Z(n30760) );
  NAND U39631 ( .A(n30764), .B(n30765), .Z(n30763) );
  NANDN U39632 ( .A(n30766), .B(n30767), .Z(n30765) );
  NANDN U39633 ( .A(n30767), .B(n30766), .Z(n30762) );
  AND U39634 ( .A(n30768), .B(n30769), .Z(n30757) );
  NAND U39635 ( .A(n30770), .B(n30771), .Z(n30769) );
  NANDN U39636 ( .A(n30772), .B(n30773), .Z(n30771) );
  NANDN U39637 ( .A(n30773), .B(n30772), .Z(n30768) );
  IV U39638 ( .A(n30774), .Z(n30773) );
  AND U39639 ( .A(n30775), .B(n30776), .Z(n30759) );
  NAND U39640 ( .A(n30777), .B(n30778), .Z(n30776) );
  NANDN U39641 ( .A(n30779), .B(n30780), .Z(n30778) );
  NANDN U39642 ( .A(n30780), .B(n30779), .Z(n30775) );
  XOR U39643 ( .A(n30772), .B(n30781), .Z(N62648) );
  XNOR U39644 ( .A(n30770), .B(n30774), .Z(n30781) );
  XOR U39645 ( .A(n30767), .B(n30782), .Z(n30774) );
  XNOR U39646 ( .A(n30764), .B(n30766), .Z(n30782) );
  AND U39647 ( .A(n30783), .B(n30784), .Z(n30766) );
  NANDN U39648 ( .A(n30785), .B(n30786), .Z(n30784) );
  OR U39649 ( .A(n30787), .B(n30788), .Z(n30786) );
  IV U39650 ( .A(n30789), .Z(n30788) );
  NANDN U39651 ( .A(n30789), .B(n30787), .Z(n30783) );
  AND U39652 ( .A(n30790), .B(n30791), .Z(n30764) );
  NAND U39653 ( .A(n30792), .B(n30793), .Z(n30791) );
  NANDN U39654 ( .A(n30794), .B(n30795), .Z(n30793) );
  NANDN U39655 ( .A(n30795), .B(n30794), .Z(n30790) );
  IV U39656 ( .A(n30796), .Z(n30795) );
  NAND U39657 ( .A(n30797), .B(n30798), .Z(n30767) );
  NANDN U39658 ( .A(n30799), .B(n30800), .Z(n30798) );
  NANDN U39659 ( .A(n30801), .B(n30802), .Z(n30800) );
  NANDN U39660 ( .A(n30802), .B(n30801), .Z(n30797) );
  IV U39661 ( .A(n30803), .Z(n30801) );
  AND U39662 ( .A(n30804), .B(n30805), .Z(n30770) );
  NAND U39663 ( .A(n30806), .B(n30807), .Z(n30805) );
  NANDN U39664 ( .A(n30808), .B(n30809), .Z(n30807) );
  NANDN U39665 ( .A(n30809), .B(n30808), .Z(n30804) );
  XOR U39666 ( .A(n30780), .B(n30810), .Z(n30772) );
  XNOR U39667 ( .A(n30777), .B(n30779), .Z(n30810) );
  AND U39668 ( .A(n30811), .B(n30812), .Z(n30779) );
  NANDN U39669 ( .A(n30813), .B(n30814), .Z(n30812) );
  OR U39670 ( .A(n30815), .B(n30816), .Z(n30814) );
  IV U39671 ( .A(n30817), .Z(n30816) );
  NANDN U39672 ( .A(n30817), .B(n30815), .Z(n30811) );
  AND U39673 ( .A(n30818), .B(n30819), .Z(n30777) );
  NAND U39674 ( .A(n30820), .B(n30821), .Z(n30819) );
  NANDN U39675 ( .A(n30822), .B(n30823), .Z(n30821) );
  NANDN U39676 ( .A(n30823), .B(n30822), .Z(n30818) );
  IV U39677 ( .A(n30824), .Z(n30823) );
  NAND U39678 ( .A(n30825), .B(n30826), .Z(n30780) );
  NANDN U39679 ( .A(n30827), .B(n30828), .Z(n30826) );
  NANDN U39680 ( .A(n30829), .B(n30830), .Z(n30828) );
  NANDN U39681 ( .A(n30830), .B(n30829), .Z(n30825) );
  IV U39682 ( .A(n30831), .Z(n30829) );
  XOR U39683 ( .A(n30806), .B(n30832), .Z(N62647) );
  XNOR U39684 ( .A(n30809), .B(n30808), .Z(n30832) );
  XNOR U39685 ( .A(n30820), .B(n30833), .Z(n30808) );
  XNOR U39686 ( .A(n30824), .B(n30822), .Z(n30833) );
  XOR U39687 ( .A(n30830), .B(n30834), .Z(n30822) );
  XNOR U39688 ( .A(n30827), .B(n30831), .Z(n30834) );
  AND U39689 ( .A(n30835), .B(n30836), .Z(n30831) );
  NAND U39690 ( .A(n30837), .B(n30838), .Z(n30836) );
  NAND U39691 ( .A(n30839), .B(n30840), .Z(n30835) );
  AND U39692 ( .A(n30841), .B(n30842), .Z(n30827) );
  NAND U39693 ( .A(n30843), .B(n30844), .Z(n30842) );
  NAND U39694 ( .A(n30845), .B(n30846), .Z(n30841) );
  NANDN U39695 ( .A(n30847), .B(n30848), .Z(n30830) );
  ANDN U39696 ( .B(n30849), .A(n30850), .Z(n30824) );
  XNOR U39697 ( .A(n30815), .B(n30851), .Z(n30820) );
  XNOR U39698 ( .A(n30813), .B(n30817), .Z(n30851) );
  AND U39699 ( .A(n30852), .B(n30853), .Z(n30817) );
  NAND U39700 ( .A(n30854), .B(n30855), .Z(n30853) );
  NAND U39701 ( .A(n30856), .B(n30857), .Z(n30852) );
  AND U39702 ( .A(n30858), .B(n30859), .Z(n30813) );
  NAND U39703 ( .A(n30860), .B(n30861), .Z(n30859) );
  NAND U39704 ( .A(n30862), .B(n30863), .Z(n30858) );
  AND U39705 ( .A(n30864), .B(n30865), .Z(n30815) );
  NAND U39706 ( .A(n30866), .B(n30867), .Z(n30809) );
  XNOR U39707 ( .A(n30792), .B(n30868), .Z(n30806) );
  XNOR U39708 ( .A(n30796), .B(n30794), .Z(n30868) );
  XOR U39709 ( .A(n30802), .B(n30869), .Z(n30794) );
  XNOR U39710 ( .A(n30799), .B(n30803), .Z(n30869) );
  AND U39711 ( .A(n30870), .B(n30871), .Z(n30803) );
  NAND U39712 ( .A(n30872), .B(n30873), .Z(n30871) );
  NAND U39713 ( .A(n30874), .B(n30875), .Z(n30870) );
  AND U39714 ( .A(n30876), .B(n30877), .Z(n30799) );
  NAND U39715 ( .A(n30878), .B(n30879), .Z(n30877) );
  NAND U39716 ( .A(n30880), .B(n30881), .Z(n30876) );
  NANDN U39717 ( .A(n30882), .B(n30883), .Z(n30802) );
  ANDN U39718 ( .B(n30884), .A(n30885), .Z(n30796) );
  XNOR U39719 ( .A(n30787), .B(n30886), .Z(n30792) );
  XNOR U39720 ( .A(n30785), .B(n30789), .Z(n30886) );
  AND U39721 ( .A(n30887), .B(n30888), .Z(n30789) );
  NAND U39722 ( .A(n30889), .B(n30890), .Z(n30888) );
  NAND U39723 ( .A(n30891), .B(n30892), .Z(n30887) );
  AND U39724 ( .A(n30893), .B(n30894), .Z(n30785) );
  NAND U39725 ( .A(n30895), .B(n30896), .Z(n30894) );
  NAND U39726 ( .A(n30897), .B(n30898), .Z(n30893) );
  AND U39727 ( .A(n30899), .B(n30900), .Z(n30787) );
  XOR U39728 ( .A(n30867), .B(n30866), .Z(N62646) );
  XNOR U39729 ( .A(n30884), .B(n30885), .Z(n30866) );
  XNOR U39730 ( .A(n30899), .B(n30900), .Z(n30885) );
  XOR U39731 ( .A(n30896), .B(n30895), .Z(n30900) );
  XOR U39732 ( .A(y[3804]), .B(x[3804]), .Z(n30895) );
  XOR U39733 ( .A(n30898), .B(n30897), .Z(n30896) );
  XOR U39734 ( .A(y[3806]), .B(x[3806]), .Z(n30897) );
  XOR U39735 ( .A(y[3805]), .B(x[3805]), .Z(n30898) );
  XOR U39736 ( .A(n30890), .B(n30889), .Z(n30899) );
  XOR U39737 ( .A(n30892), .B(n30891), .Z(n30889) );
  XOR U39738 ( .A(y[3803]), .B(x[3803]), .Z(n30891) );
  XOR U39739 ( .A(y[3802]), .B(x[3802]), .Z(n30892) );
  XOR U39740 ( .A(y[3801]), .B(x[3801]), .Z(n30890) );
  XNOR U39741 ( .A(n30883), .B(n30882), .Z(n30884) );
  XNOR U39742 ( .A(n30879), .B(n30878), .Z(n30882) );
  XOR U39743 ( .A(n30881), .B(n30880), .Z(n30878) );
  XOR U39744 ( .A(y[3800]), .B(x[3800]), .Z(n30880) );
  XOR U39745 ( .A(y[3799]), .B(x[3799]), .Z(n30881) );
  XOR U39746 ( .A(y[3798]), .B(x[3798]), .Z(n30879) );
  XOR U39747 ( .A(n30873), .B(n30872), .Z(n30883) );
  XOR U39748 ( .A(n30875), .B(n30874), .Z(n30872) );
  XOR U39749 ( .A(y[3797]), .B(x[3797]), .Z(n30874) );
  XOR U39750 ( .A(y[3796]), .B(x[3796]), .Z(n30875) );
  XOR U39751 ( .A(y[3795]), .B(x[3795]), .Z(n30873) );
  XNOR U39752 ( .A(n30849), .B(n30850), .Z(n30867) );
  XNOR U39753 ( .A(n30864), .B(n30865), .Z(n30850) );
  XOR U39754 ( .A(n30861), .B(n30860), .Z(n30865) );
  XOR U39755 ( .A(y[3792]), .B(x[3792]), .Z(n30860) );
  XOR U39756 ( .A(n30863), .B(n30862), .Z(n30861) );
  XOR U39757 ( .A(y[3794]), .B(x[3794]), .Z(n30862) );
  XOR U39758 ( .A(y[3793]), .B(x[3793]), .Z(n30863) );
  XOR U39759 ( .A(n30855), .B(n30854), .Z(n30864) );
  XOR U39760 ( .A(n30857), .B(n30856), .Z(n30854) );
  XOR U39761 ( .A(y[3791]), .B(x[3791]), .Z(n30856) );
  XOR U39762 ( .A(y[3790]), .B(x[3790]), .Z(n30857) );
  XOR U39763 ( .A(y[3789]), .B(x[3789]), .Z(n30855) );
  XNOR U39764 ( .A(n30848), .B(n30847), .Z(n30849) );
  XNOR U39765 ( .A(n30844), .B(n30843), .Z(n30847) );
  XOR U39766 ( .A(n30846), .B(n30845), .Z(n30843) );
  XOR U39767 ( .A(y[3788]), .B(x[3788]), .Z(n30845) );
  XOR U39768 ( .A(y[3787]), .B(x[3787]), .Z(n30846) );
  XOR U39769 ( .A(y[3786]), .B(x[3786]), .Z(n30844) );
  XOR U39770 ( .A(n30838), .B(n30837), .Z(n30848) );
  XOR U39771 ( .A(n30840), .B(n30839), .Z(n30837) );
  XOR U39772 ( .A(y[3785]), .B(x[3785]), .Z(n30839) );
  XOR U39773 ( .A(y[3784]), .B(x[3784]), .Z(n30840) );
  XOR U39774 ( .A(y[3783]), .B(x[3783]), .Z(n30838) );
  NAND U39775 ( .A(n30901), .B(n30902), .Z(N62637) );
  NAND U39776 ( .A(n30903), .B(n30904), .Z(n30902) );
  NANDN U39777 ( .A(n30905), .B(n30906), .Z(n30904) );
  NANDN U39778 ( .A(n30906), .B(n30905), .Z(n30901) );
  XOR U39779 ( .A(n30905), .B(n30907), .Z(N62636) );
  XNOR U39780 ( .A(n30903), .B(n30906), .Z(n30907) );
  NAND U39781 ( .A(n30908), .B(n30909), .Z(n30906) );
  NAND U39782 ( .A(n30910), .B(n30911), .Z(n30909) );
  NANDN U39783 ( .A(n30912), .B(n30913), .Z(n30911) );
  NANDN U39784 ( .A(n30913), .B(n30912), .Z(n30908) );
  AND U39785 ( .A(n30914), .B(n30915), .Z(n30903) );
  NAND U39786 ( .A(n30916), .B(n30917), .Z(n30915) );
  NANDN U39787 ( .A(n30918), .B(n30919), .Z(n30917) );
  NANDN U39788 ( .A(n30919), .B(n30918), .Z(n30914) );
  IV U39789 ( .A(n30920), .Z(n30919) );
  AND U39790 ( .A(n30921), .B(n30922), .Z(n30905) );
  NAND U39791 ( .A(n30923), .B(n30924), .Z(n30922) );
  NANDN U39792 ( .A(n30925), .B(n30926), .Z(n30924) );
  NANDN U39793 ( .A(n30926), .B(n30925), .Z(n30921) );
  XOR U39794 ( .A(n30918), .B(n30927), .Z(N62635) );
  XNOR U39795 ( .A(n30916), .B(n30920), .Z(n30927) );
  XOR U39796 ( .A(n30913), .B(n30928), .Z(n30920) );
  XNOR U39797 ( .A(n30910), .B(n30912), .Z(n30928) );
  AND U39798 ( .A(n30929), .B(n30930), .Z(n30912) );
  NANDN U39799 ( .A(n30931), .B(n30932), .Z(n30930) );
  OR U39800 ( .A(n30933), .B(n30934), .Z(n30932) );
  IV U39801 ( .A(n30935), .Z(n30934) );
  NANDN U39802 ( .A(n30935), .B(n30933), .Z(n30929) );
  AND U39803 ( .A(n30936), .B(n30937), .Z(n30910) );
  NAND U39804 ( .A(n30938), .B(n30939), .Z(n30937) );
  NANDN U39805 ( .A(n30940), .B(n30941), .Z(n30939) );
  NANDN U39806 ( .A(n30941), .B(n30940), .Z(n30936) );
  IV U39807 ( .A(n30942), .Z(n30941) );
  NAND U39808 ( .A(n30943), .B(n30944), .Z(n30913) );
  NANDN U39809 ( .A(n30945), .B(n30946), .Z(n30944) );
  NANDN U39810 ( .A(n30947), .B(n30948), .Z(n30946) );
  NANDN U39811 ( .A(n30948), .B(n30947), .Z(n30943) );
  IV U39812 ( .A(n30949), .Z(n30947) );
  AND U39813 ( .A(n30950), .B(n30951), .Z(n30916) );
  NAND U39814 ( .A(n30952), .B(n30953), .Z(n30951) );
  NANDN U39815 ( .A(n30954), .B(n30955), .Z(n30953) );
  NANDN U39816 ( .A(n30955), .B(n30954), .Z(n30950) );
  XOR U39817 ( .A(n30926), .B(n30956), .Z(n30918) );
  XNOR U39818 ( .A(n30923), .B(n30925), .Z(n30956) );
  AND U39819 ( .A(n30957), .B(n30958), .Z(n30925) );
  NANDN U39820 ( .A(n30959), .B(n30960), .Z(n30958) );
  OR U39821 ( .A(n30961), .B(n30962), .Z(n30960) );
  IV U39822 ( .A(n30963), .Z(n30962) );
  NANDN U39823 ( .A(n30963), .B(n30961), .Z(n30957) );
  AND U39824 ( .A(n30964), .B(n30965), .Z(n30923) );
  NAND U39825 ( .A(n30966), .B(n30967), .Z(n30965) );
  NANDN U39826 ( .A(n30968), .B(n30969), .Z(n30967) );
  NANDN U39827 ( .A(n30969), .B(n30968), .Z(n30964) );
  IV U39828 ( .A(n30970), .Z(n30969) );
  NAND U39829 ( .A(n30971), .B(n30972), .Z(n30926) );
  NANDN U39830 ( .A(n30973), .B(n30974), .Z(n30972) );
  NANDN U39831 ( .A(n30975), .B(n30976), .Z(n30974) );
  NANDN U39832 ( .A(n30976), .B(n30975), .Z(n30971) );
  IV U39833 ( .A(n30977), .Z(n30975) );
  XOR U39834 ( .A(n30952), .B(n30978), .Z(N62634) );
  XNOR U39835 ( .A(n30955), .B(n30954), .Z(n30978) );
  XNOR U39836 ( .A(n30966), .B(n30979), .Z(n30954) );
  XNOR U39837 ( .A(n30970), .B(n30968), .Z(n30979) );
  XOR U39838 ( .A(n30976), .B(n30980), .Z(n30968) );
  XNOR U39839 ( .A(n30973), .B(n30977), .Z(n30980) );
  AND U39840 ( .A(n30981), .B(n30982), .Z(n30977) );
  NAND U39841 ( .A(n30983), .B(n30984), .Z(n30982) );
  NAND U39842 ( .A(n30985), .B(n30986), .Z(n30981) );
  AND U39843 ( .A(n30987), .B(n30988), .Z(n30973) );
  NAND U39844 ( .A(n30989), .B(n30990), .Z(n30988) );
  NAND U39845 ( .A(n30991), .B(n30992), .Z(n30987) );
  NANDN U39846 ( .A(n30993), .B(n30994), .Z(n30976) );
  ANDN U39847 ( .B(n30995), .A(n30996), .Z(n30970) );
  XNOR U39848 ( .A(n30961), .B(n30997), .Z(n30966) );
  XNOR U39849 ( .A(n30959), .B(n30963), .Z(n30997) );
  AND U39850 ( .A(n30998), .B(n30999), .Z(n30963) );
  NAND U39851 ( .A(n31000), .B(n31001), .Z(n30999) );
  NAND U39852 ( .A(n31002), .B(n31003), .Z(n30998) );
  AND U39853 ( .A(n31004), .B(n31005), .Z(n30959) );
  NAND U39854 ( .A(n31006), .B(n31007), .Z(n31005) );
  NAND U39855 ( .A(n31008), .B(n31009), .Z(n31004) );
  AND U39856 ( .A(n31010), .B(n31011), .Z(n30961) );
  NAND U39857 ( .A(n31012), .B(n31013), .Z(n30955) );
  XNOR U39858 ( .A(n30938), .B(n31014), .Z(n30952) );
  XNOR U39859 ( .A(n30942), .B(n30940), .Z(n31014) );
  XOR U39860 ( .A(n30948), .B(n31015), .Z(n30940) );
  XNOR U39861 ( .A(n30945), .B(n30949), .Z(n31015) );
  AND U39862 ( .A(n31016), .B(n31017), .Z(n30949) );
  NAND U39863 ( .A(n31018), .B(n31019), .Z(n31017) );
  NAND U39864 ( .A(n31020), .B(n31021), .Z(n31016) );
  AND U39865 ( .A(n31022), .B(n31023), .Z(n30945) );
  NAND U39866 ( .A(n31024), .B(n31025), .Z(n31023) );
  NAND U39867 ( .A(n31026), .B(n31027), .Z(n31022) );
  NANDN U39868 ( .A(n31028), .B(n31029), .Z(n30948) );
  ANDN U39869 ( .B(n31030), .A(n31031), .Z(n30942) );
  XNOR U39870 ( .A(n30933), .B(n31032), .Z(n30938) );
  XNOR U39871 ( .A(n30931), .B(n30935), .Z(n31032) );
  AND U39872 ( .A(n31033), .B(n31034), .Z(n30935) );
  NAND U39873 ( .A(n31035), .B(n31036), .Z(n31034) );
  NAND U39874 ( .A(n31037), .B(n31038), .Z(n31033) );
  AND U39875 ( .A(n31039), .B(n31040), .Z(n30931) );
  NAND U39876 ( .A(n31041), .B(n31042), .Z(n31040) );
  NAND U39877 ( .A(n31043), .B(n31044), .Z(n31039) );
  AND U39878 ( .A(n31045), .B(n31046), .Z(n30933) );
  XOR U39879 ( .A(n31013), .B(n31012), .Z(N62633) );
  XNOR U39880 ( .A(n31030), .B(n31031), .Z(n31012) );
  XNOR U39881 ( .A(n31045), .B(n31046), .Z(n31031) );
  XOR U39882 ( .A(n31042), .B(n31041), .Z(n31046) );
  XOR U39883 ( .A(y[3780]), .B(x[3780]), .Z(n31041) );
  XOR U39884 ( .A(n31044), .B(n31043), .Z(n31042) );
  XOR U39885 ( .A(y[3782]), .B(x[3782]), .Z(n31043) );
  XOR U39886 ( .A(y[3781]), .B(x[3781]), .Z(n31044) );
  XOR U39887 ( .A(n31036), .B(n31035), .Z(n31045) );
  XOR U39888 ( .A(n31038), .B(n31037), .Z(n31035) );
  XOR U39889 ( .A(y[3779]), .B(x[3779]), .Z(n31037) );
  XOR U39890 ( .A(y[3778]), .B(x[3778]), .Z(n31038) );
  XOR U39891 ( .A(y[3777]), .B(x[3777]), .Z(n31036) );
  XNOR U39892 ( .A(n31029), .B(n31028), .Z(n31030) );
  XNOR U39893 ( .A(n31025), .B(n31024), .Z(n31028) );
  XOR U39894 ( .A(n31027), .B(n31026), .Z(n31024) );
  XOR U39895 ( .A(y[3776]), .B(x[3776]), .Z(n31026) );
  XOR U39896 ( .A(y[3775]), .B(x[3775]), .Z(n31027) );
  XOR U39897 ( .A(y[3774]), .B(x[3774]), .Z(n31025) );
  XOR U39898 ( .A(n31019), .B(n31018), .Z(n31029) );
  XOR U39899 ( .A(n31021), .B(n31020), .Z(n31018) );
  XOR U39900 ( .A(y[3773]), .B(x[3773]), .Z(n31020) );
  XOR U39901 ( .A(y[3772]), .B(x[3772]), .Z(n31021) );
  XOR U39902 ( .A(y[3771]), .B(x[3771]), .Z(n31019) );
  XNOR U39903 ( .A(n30995), .B(n30996), .Z(n31013) );
  XNOR U39904 ( .A(n31010), .B(n31011), .Z(n30996) );
  XOR U39905 ( .A(n31007), .B(n31006), .Z(n31011) );
  XOR U39906 ( .A(y[3768]), .B(x[3768]), .Z(n31006) );
  XOR U39907 ( .A(n31009), .B(n31008), .Z(n31007) );
  XOR U39908 ( .A(y[3770]), .B(x[3770]), .Z(n31008) );
  XOR U39909 ( .A(y[3769]), .B(x[3769]), .Z(n31009) );
  XOR U39910 ( .A(n31001), .B(n31000), .Z(n31010) );
  XOR U39911 ( .A(n31003), .B(n31002), .Z(n31000) );
  XOR U39912 ( .A(y[3767]), .B(x[3767]), .Z(n31002) );
  XOR U39913 ( .A(y[3766]), .B(x[3766]), .Z(n31003) );
  XOR U39914 ( .A(y[3765]), .B(x[3765]), .Z(n31001) );
  XNOR U39915 ( .A(n30994), .B(n30993), .Z(n30995) );
  XNOR U39916 ( .A(n30990), .B(n30989), .Z(n30993) );
  XOR U39917 ( .A(n30992), .B(n30991), .Z(n30989) );
  XOR U39918 ( .A(y[3764]), .B(x[3764]), .Z(n30991) );
  XOR U39919 ( .A(y[3763]), .B(x[3763]), .Z(n30992) );
  XOR U39920 ( .A(y[3762]), .B(x[3762]), .Z(n30990) );
  XOR U39921 ( .A(n30984), .B(n30983), .Z(n30994) );
  XOR U39922 ( .A(n30986), .B(n30985), .Z(n30983) );
  XOR U39923 ( .A(y[3761]), .B(x[3761]), .Z(n30985) );
  XOR U39924 ( .A(y[3760]), .B(x[3760]), .Z(n30986) );
  XOR U39925 ( .A(y[3759]), .B(x[3759]), .Z(n30984) );
  NAND U39926 ( .A(n31047), .B(n31048), .Z(N62624) );
  NAND U39927 ( .A(n31049), .B(n31050), .Z(n31048) );
  NANDN U39928 ( .A(n31051), .B(n31052), .Z(n31050) );
  NANDN U39929 ( .A(n31052), .B(n31051), .Z(n31047) );
  XOR U39930 ( .A(n31051), .B(n31053), .Z(N62623) );
  XNOR U39931 ( .A(n31049), .B(n31052), .Z(n31053) );
  NAND U39932 ( .A(n31054), .B(n31055), .Z(n31052) );
  NAND U39933 ( .A(n31056), .B(n31057), .Z(n31055) );
  NANDN U39934 ( .A(n31058), .B(n31059), .Z(n31057) );
  NANDN U39935 ( .A(n31059), .B(n31058), .Z(n31054) );
  AND U39936 ( .A(n31060), .B(n31061), .Z(n31049) );
  NAND U39937 ( .A(n31062), .B(n31063), .Z(n31061) );
  NANDN U39938 ( .A(n31064), .B(n31065), .Z(n31063) );
  NANDN U39939 ( .A(n31065), .B(n31064), .Z(n31060) );
  IV U39940 ( .A(n31066), .Z(n31065) );
  AND U39941 ( .A(n31067), .B(n31068), .Z(n31051) );
  NAND U39942 ( .A(n31069), .B(n31070), .Z(n31068) );
  NANDN U39943 ( .A(n31071), .B(n31072), .Z(n31070) );
  NANDN U39944 ( .A(n31072), .B(n31071), .Z(n31067) );
  XOR U39945 ( .A(n31064), .B(n31073), .Z(N62622) );
  XNOR U39946 ( .A(n31062), .B(n31066), .Z(n31073) );
  XOR U39947 ( .A(n31059), .B(n31074), .Z(n31066) );
  XNOR U39948 ( .A(n31056), .B(n31058), .Z(n31074) );
  AND U39949 ( .A(n31075), .B(n31076), .Z(n31058) );
  NANDN U39950 ( .A(n31077), .B(n31078), .Z(n31076) );
  OR U39951 ( .A(n31079), .B(n31080), .Z(n31078) );
  IV U39952 ( .A(n31081), .Z(n31080) );
  NANDN U39953 ( .A(n31081), .B(n31079), .Z(n31075) );
  AND U39954 ( .A(n31082), .B(n31083), .Z(n31056) );
  NAND U39955 ( .A(n31084), .B(n31085), .Z(n31083) );
  NANDN U39956 ( .A(n31086), .B(n31087), .Z(n31085) );
  NANDN U39957 ( .A(n31087), .B(n31086), .Z(n31082) );
  IV U39958 ( .A(n31088), .Z(n31087) );
  NAND U39959 ( .A(n31089), .B(n31090), .Z(n31059) );
  NANDN U39960 ( .A(n31091), .B(n31092), .Z(n31090) );
  NANDN U39961 ( .A(n31093), .B(n31094), .Z(n31092) );
  NANDN U39962 ( .A(n31094), .B(n31093), .Z(n31089) );
  IV U39963 ( .A(n31095), .Z(n31093) );
  AND U39964 ( .A(n31096), .B(n31097), .Z(n31062) );
  NAND U39965 ( .A(n31098), .B(n31099), .Z(n31097) );
  NANDN U39966 ( .A(n31100), .B(n31101), .Z(n31099) );
  NANDN U39967 ( .A(n31101), .B(n31100), .Z(n31096) );
  XOR U39968 ( .A(n31072), .B(n31102), .Z(n31064) );
  XNOR U39969 ( .A(n31069), .B(n31071), .Z(n31102) );
  AND U39970 ( .A(n31103), .B(n31104), .Z(n31071) );
  NANDN U39971 ( .A(n31105), .B(n31106), .Z(n31104) );
  OR U39972 ( .A(n31107), .B(n31108), .Z(n31106) );
  IV U39973 ( .A(n31109), .Z(n31108) );
  NANDN U39974 ( .A(n31109), .B(n31107), .Z(n31103) );
  AND U39975 ( .A(n31110), .B(n31111), .Z(n31069) );
  NAND U39976 ( .A(n31112), .B(n31113), .Z(n31111) );
  NANDN U39977 ( .A(n31114), .B(n31115), .Z(n31113) );
  NANDN U39978 ( .A(n31115), .B(n31114), .Z(n31110) );
  IV U39979 ( .A(n31116), .Z(n31115) );
  NAND U39980 ( .A(n31117), .B(n31118), .Z(n31072) );
  NANDN U39981 ( .A(n31119), .B(n31120), .Z(n31118) );
  NANDN U39982 ( .A(n31121), .B(n31122), .Z(n31120) );
  NANDN U39983 ( .A(n31122), .B(n31121), .Z(n31117) );
  IV U39984 ( .A(n31123), .Z(n31121) );
  XOR U39985 ( .A(n31098), .B(n31124), .Z(N62621) );
  XNOR U39986 ( .A(n31101), .B(n31100), .Z(n31124) );
  XNOR U39987 ( .A(n31112), .B(n31125), .Z(n31100) );
  XNOR U39988 ( .A(n31116), .B(n31114), .Z(n31125) );
  XOR U39989 ( .A(n31122), .B(n31126), .Z(n31114) );
  XNOR U39990 ( .A(n31119), .B(n31123), .Z(n31126) );
  AND U39991 ( .A(n31127), .B(n31128), .Z(n31123) );
  NAND U39992 ( .A(n31129), .B(n31130), .Z(n31128) );
  NAND U39993 ( .A(n31131), .B(n31132), .Z(n31127) );
  AND U39994 ( .A(n31133), .B(n31134), .Z(n31119) );
  NAND U39995 ( .A(n31135), .B(n31136), .Z(n31134) );
  NAND U39996 ( .A(n31137), .B(n31138), .Z(n31133) );
  NANDN U39997 ( .A(n31139), .B(n31140), .Z(n31122) );
  ANDN U39998 ( .B(n31141), .A(n31142), .Z(n31116) );
  XNOR U39999 ( .A(n31107), .B(n31143), .Z(n31112) );
  XNOR U40000 ( .A(n31105), .B(n31109), .Z(n31143) );
  AND U40001 ( .A(n31144), .B(n31145), .Z(n31109) );
  NAND U40002 ( .A(n31146), .B(n31147), .Z(n31145) );
  NAND U40003 ( .A(n31148), .B(n31149), .Z(n31144) );
  AND U40004 ( .A(n31150), .B(n31151), .Z(n31105) );
  NAND U40005 ( .A(n31152), .B(n31153), .Z(n31151) );
  NAND U40006 ( .A(n31154), .B(n31155), .Z(n31150) );
  AND U40007 ( .A(n31156), .B(n31157), .Z(n31107) );
  NAND U40008 ( .A(n31158), .B(n31159), .Z(n31101) );
  XNOR U40009 ( .A(n31084), .B(n31160), .Z(n31098) );
  XNOR U40010 ( .A(n31088), .B(n31086), .Z(n31160) );
  XOR U40011 ( .A(n31094), .B(n31161), .Z(n31086) );
  XNOR U40012 ( .A(n31091), .B(n31095), .Z(n31161) );
  AND U40013 ( .A(n31162), .B(n31163), .Z(n31095) );
  NAND U40014 ( .A(n31164), .B(n31165), .Z(n31163) );
  NAND U40015 ( .A(n31166), .B(n31167), .Z(n31162) );
  AND U40016 ( .A(n31168), .B(n31169), .Z(n31091) );
  NAND U40017 ( .A(n31170), .B(n31171), .Z(n31169) );
  NAND U40018 ( .A(n31172), .B(n31173), .Z(n31168) );
  NANDN U40019 ( .A(n31174), .B(n31175), .Z(n31094) );
  ANDN U40020 ( .B(n31176), .A(n31177), .Z(n31088) );
  XNOR U40021 ( .A(n31079), .B(n31178), .Z(n31084) );
  XNOR U40022 ( .A(n31077), .B(n31081), .Z(n31178) );
  AND U40023 ( .A(n31179), .B(n31180), .Z(n31081) );
  NAND U40024 ( .A(n31181), .B(n31182), .Z(n31180) );
  NAND U40025 ( .A(n31183), .B(n31184), .Z(n31179) );
  AND U40026 ( .A(n31185), .B(n31186), .Z(n31077) );
  NAND U40027 ( .A(n31187), .B(n31188), .Z(n31186) );
  NAND U40028 ( .A(n31189), .B(n31190), .Z(n31185) );
  AND U40029 ( .A(n31191), .B(n31192), .Z(n31079) );
  XOR U40030 ( .A(n31159), .B(n31158), .Z(N62620) );
  XNOR U40031 ( .A(n31176), .B(n31177), .Z(n31158) );
  XNOR U40032 ( .A(n31191), .B(n31192), .Z(n31177) );
  XOR U40033 ( .A(n31188), .B(n31187), .Z(n31192) );
  XOR U40034 ( .A(y[3756]), .B(x[3756]), .Z(n31187) );
  XOR U40035 ( .A(n31190), .B(n31189), .Z(n31188) );
  XOR U40036 ( .A(y[3758]), .B(x[3758]), .Z(n31189) );
  XOR U40037 ( .A(y[3757]), .B(x[3757]), .Z(n31190) );
  XOR U40038 ( .A(n31182), .B(n31181), .Z(n31191) );
  XOR U40039 ( .A(n31184), .B(n31183), .Z(n31181) );
  XOR U40040 ( .A(y[3755]), .B(x[3755]), .Z(n31183) );
  XOR U40041 ( .A(y[3754]), .B(x[3754]), .Z(n31184) );
  XOR U40042 ( .A(y[3753]), .B(x[3753]), .Z(n31182) );
  XNOR U40043 ( .A(n31175), .B(n31174), .Z(n31176) );
  XNOR U40044 ( .A(n31171), .B(n31170), .Z(n31174) );
  XOR U40045 ( .A(n31173), .B(n31172), .Z(n31170) );
  XOR U40046 ( .A(y[3752]), .B(x[3752]), .Z(n31172) );
  XOR U40047 ( .A(y[3751]), .B(x[3751]), .Z(n31173) );
  XOR U40048 ( .A(y[3750]), .B(x[3750]), .Z(n31171) );
  XOR U40049 ( .A(n31165), .B(n31164), .Z(n31175) );
  XOR U40050 ( .A(n31167), .B(n31166), .Z(n31164) );
  XOR U40051 ( .A(y[3749]), .B(x[3749]), .Z(n31166) );
  XOR U40052 ( .A(y[3748]), .B(x[3748]), .Z(n31167) );
  XOR U40053 ( .A(y[3747]), .B(x[3747]), .Z(n31165) );
  XNOR U40054 ( .A(n31141), .B(n31142), .Z(n31159) );
  XNOR U40055 ( .A(n31156), .B(n31157), .Z(n31142) );
  XOR U40056 ( .A(n31153), .B(n31152), .Z(n31157) );
  XOR U40057 ( .A(y[3744]), .B(x[3744]), .Z(n31152) );
  XOR U40058 ( .A(n31155), .B(n31154), .Z(n31153) );
  XOR U40059 ( .A(y[3746]), .B(x[3746]), .Z(n31154) );
  XOR U40060 ( .A(y[3745]), .B(x[3745]), .Z(n31155) );
  XOR U40061 ( .A(n31147), .B(n31146), .Z(n31156) );
  XOR U40062 ( .A(n31149), .B(n31148), .Z(n31146) );
  XOR U40063 ( .A(y[3743]), .B(x[3743]), .Z(n31148) );
  XOR U40064 ( .A(y[3742]), .B(x[3742]), .Z(n31149) );
  XOR U40065 ( .A(y[3741]), .B(x[3741]), .Z(n31147) );
  XNOR U40066 ( .A(n31140), .B(n31139), .Z(n31141) );
  XNOR U40067 ( .A(n31136), .B(n31135), .Z(n31139) );
  XOR U40068 ( .A(n31138), .B(n31137), .Z(n31135) );
  XOR U40069 ( .A(y[3740]), .B(x[3740]), .Z(n31137) );
  XOR U40070 ( .A(y[3739]), .B(x[3739]), .Z(n31138) );
  XOR U40071 ( .A(y[3738]), .B(x[3738]), .Z(n31136) );
  XOR U40072 ( .A(n31130), .B(n31129), .Z(n31140) );
  XOR U40073 ( .A(n31132), .B(n31131), .Z(n31129) );
  XOR U40074 ( .A(y[3737]), .B(x[3737]), .Z(n31131) );
  XOR U40075 ( .A(y[3736]), .B(x[3736]), .Z(n31132) );
  XOR U40076 ( .A(y[3735]), .B(x[3735]), .Z(n31130) );
  NAND U40077 ( .A(n31193), .B(n31194), .Z(N62611) );
  NAND U40078 ( .A(n31195), .B(n31196), .Z(n31194) );
  NANDN U40079 ( .A(n31197), .B(n31198), .Z(n31196) );
  NANDN U40080 ( .A(n31198), .B(n31197), .Z(n31193) );
  XOR U40081 ( .A(n31197), .B(n31199), .Z(N62610) );
  XNOR U40082 ( .A(n31195), .B(n31198), .Z(n31199) );
  NAND U40083 ( .A(n31200), .B(n31201), .Z(n31198) );
  NAND U40084 ( .A(n31202), .B(n31203), .Z(n31201) );
  NANDN U40085 ( .A(n31204), .B(n31205), .Z(n31203) );
  NANDN U40086 ( .A(n31205), .B(n31204), .Z(n31200) );
  AND U40087 ( .A(n31206), .B(n31207), .Z(n31195) );
  NAND U40088 ( .A(n31208), .B(n31209), .Z(n31207) );
  NANDN U40089 ( .A(n31210), .B(n31211), .Z(n31209) );
  NANDN U40090 ( .A(n31211), .B(n31210), .Z(n31206) );
  IV U40091 ( .A(n31212), .Z(n31211) );
  AND U40092 ( .A(n31213), .B(n31214), .Z(n31197) );
  NAND U40093 ( .A(n31215), .B(n31216), .Z(n31214) );
  NANDN U40094 ( .A(n31217), .B(n31218), .Z(n31216) );
  NANDN U40095 ( .A(n31218), .B(n31217), .Z(n31213) );
  XOR U40096 ( .A(n31210), .B(n31219), .Z(N62609) );
  XNOR U40097 ( .A(n31208), .B(n31212), .Z(n31219) );
  XOR U40098 ( .A(n31205), .B(n31220), .Z(n31212) );
  XNOR U40099 ( .A(n31202), .B(n31204), .Z(n31220) );
  AND U40100 ( .A(n31221), .B(n31222), .Z(n31204) );
  NANDN U40101 ( .A(n31223), .B(n31224), .Z(n31222) );
  OR U40102 ( .A(n31225), .B(n31226), .Z(n31224) );
  IV U40103 ( .A(n31227), .Z(n31226) );
  NANDN U40104 ( .A(n31227), .B(n31225), .Z(n31221) );
  AND U40105 ( .A(n31228), .B(n31229), .Z(n31202) );
  NAND U40106 ( .A(n31230), .B(n31231), .Z(n31229) );
  NANDN U40107 ( .A(n31232), .B(n31233), .Z(n31231) );
  NANDN U40108 ( .A(n31233), .B(n31232), .Z(n31228) );
  IV U40109 ( .A(n31234), .Z(n31233) );
  NAND U40110 ( .A(n31235), .B(n31236), .Z(n31205) );
  NANDN U40111 ( .A(n31237), .B(n31238), .Z(n31236) );
  NANDN U40112 ( .A(n31239), .B(n31240), .Z(n31238) );
  NANDN U40113 ( .A(n31240), .B(n31239), .Z(n31235) );
  IV U40114 ( .A(n31241), .Z(n31239) );
  AND U40115 ( .A(n31242), .B(n31243), .Z(n31208) );
  NAND U40116 ( .A(n31244), .B(n31245), .Z(n31243) );
  NANDN U40117 ( .A(n31246), .B(n31247), .Z(n31245) );
  NANDN U40118 ( .A(n31247), .B(n31246), .Z(n31242) );
  XOR U40119 ( .A(n31218), .B(n31248), .Z(n31210) );
  XNOR U40120 ( .A(n31215), .B(n31217), .Z(n31248) );
  AND U40121 ( .A(n31249), .B(n31250), .Z(n31217) );
  NANDN U40122 ( .A(n31251), .B(n31252), .Z(n31250) );
  OR U40123 ( .A(n31253), .B(n31254), .Z(n31252) );
  IV U40124 ( .A(n31255), .Z(n31254) );
  NANDN U40125 ( .A(n31255), .B(n31253), .Z(n31249) );
  AND U40126 ( .A(n31256), .B(n31257), .Z(n31215) );
  NAND U40127 ( .A(n31258), .B(n31259), .Z(n31257) );
  NANDN U40128 ( .A(n31260), .B(n31261), .Z(n31259) );
  NANDN U40129 ( .A(n31261), .B(n31260), .Z(n31256) );
  IV U40130 ( .A(n31262), .Z(n31261) );
  NAND U40131 ( .A(n31263), .B(n31264), .Z(n31218) );
  NANDN U40132 ( .A(n31265), .B(n31266), .Z(n31264) );
  NANDN U40133 ( .A(n31267), .B(n31268), .Z(n31266) );
  NANDN U40134 ( .A(n31268), .B(n31267), .Z(n31263) );
  IV U40135 ( .A(n31269), .Z(n31267) );
  XOR U40136 ( .A(n31244), .B(n31270), .Z(N62608) );
  XNOR U40137 ( .A(n31247), .B(n31246), .Z(n31270) );
  XNOR U40138 ( .A(n31258), .B(n31271), .Z(n31246) );
  XNOR U40139 ( .A(n31262), .B(n31260), .Z(n31271) );
  XOR U40140 ( .A(n31268), .B(n31272), .Z(n31260) );
  XNOR U40141 ( .A(n31265), .B(n31269), .Z(n31272) );
  AND U40142 ( .A(n31273), .B(n31274), .Z(n31269) );
  NAND U40143 ( .A(n31275), .B(n31276), .Z(n31274) );
  NAND U40144 ( .A(n31277), .B(n31278), .Z(n31273) );
  AND U40145 ( .A(n31279), .B(n31280), .Z(n31265) );
  NAND U40146 ( .A(n31281), .B(n31282), .Z(n31280) );
  NAND U40147 ( .A(n31283), .B(n31284), .Z(n31279) );
  NANDN U40148 ( .A(n31285), .B(n31286), .Z(n31268) );
  ANDN U40149 ( .B(n31287), .A(n31288), .Z(n31262) );
  XNOR U40150 ( .A(n31253), .B(n31289), .Z(n31258) );
  XNOR U40151 ( .A(n31251), .B(n31255), .Z(n31289) );
  AND U40152 ( .A(n31290), .B(n31291), .Z(n31255) );
  NAND U40153 ( .A(n31292), .B(n31293), .Z(n31291) );
  NAND U40154 ( .A(n31294), .B(n31295), .Z(n31290) );
  AND U40155 ( .A(n31296), .B(n31297), .Z(n31251) );
  NAND U40156 ( .A(n31298), .B(n31299), .Z(n31297) );
  NAND U40157 ( .A(n31300), .B(n31301), .Z(n31296) );
  AND U40158 ( .A(n31302), .B(n31303), .Z(n31253) );
  NAND U40159 ( .A(n31304), .B(n31305), .Z(n31247) );
  XNOR U40160 ( .A(n31230), .B(n31306), .Z(n31244) );
  XNOR U40161 ( .A(n31234), .B(n31232), .Z(n31306) );
  XOR U40162 ( .A(n31240), .B(n31307), .Z(n31232) );
  XNOR U40163 ( .A(n31237), .B(n31241), .Z(n31307) );
  AND U40164 ( .A(n31308), .B(n31309), .Z(n31241) );
  NAND U40165 ( .A(n31310), .B(n31311), .Z(n31309) );
  NAND U40166 ( .A(n31312), .B(n31313), .Z(n31308) );
  AND U40167 ( .A(n31314), .B(n31315), .Z(n31237) );
  NAND U40168 ( .A(n31316), .B(n31317), .Z(n31315) );
  NAND U40169 ( .A(n31318), .B(n31319), .Z(n31314) );
  NANDN U40170 ( .A(n31320), .B(n31321), .Z(n31240) );
  ANDN U40171 ( .B(n31322), .A(n31323), .Z(n31234) );
  XNOR U40172 ( .A(n31225), .B(n31324), .Z(n31230) );
  XNOR U40173 ( .A(n31223), .B(n31227), .Z(n31324) );
  AND U40174 ( .A(n31325), .B(n31326), .Z(n31227) );
  NAND U40175 ( .A(n31327), .B(n31328), .Z(n31326) );
  NAND U40176 ( .A(n31329), .B(n31330), .Z(n31325) );
  AND U40177 ( .A(n31331), .B(n31332), .Z(n31223) );
  NAND U40178 ( .A(n31333), .B(n31334), .Z(n31332) );
  NAND U40179 ( .A(n31335), .B(n31336), .Z(n31331) );
  AND U40180 ( .A(n31337), .B(n31338), .Z(n31225) );
  XOR U40181 ( .A(n31305), .B(n31304), .Z(N62607) );
  XNOR U40182 ( .A(n31322), .B(n31323), .Z(n31304) );
  XNOR U40183 ( .A(n31337), .B(n31338), .Z(n31323) );
  XOR U40184 ( .A(n31334), .B(n31333), .Z(n31338) );
  XOR U40185 ( .A(y[3732]), .B(x[3732]), .Z(n31333) );
  XOR U40186 ( .A(n31336), .B(n31335), .Z(n31334) );
  XOR U40187 ( .A(y[3734]), .B(x[3734]), .Z(n31335) );
  XOR U40188 ( .A(y[3733]), .B(x[3733]), .Z(n31336) );
  XOR U40189 ( .A(n31328), .B(n31327), .Z(n31337) );
  XOR U40190 ( .A(n31330), .B(n31329), .Z(n31327) );
  XOR U40191 ( .A(y[3731]), .B(x[3731]), .Z(n31329) );
  XOR U40192 ( .A(y[3730]), .B(x[3730]), .Z(n31330) );
  XOR U40193 ( .A(y[3729]), .B(x[3729]), .Z(n31328) );
  XNOR U40194 ( .A(n31321), .B(n31320), .Z(n31322) );
  XNOR U40195 ( .A(n31317), .B(n31316), .Z(n31320) );
  XOR U40196 ( .A(n31319), .B(n31318), .Z(n31316) );
  XOR U40197 ( .A(y[3728]), .B(x[3728]), .Z(n31318) );
  XOR U40198 ( .A(y[3727]), .B(x[3727]), .Z(n31319) );
  XOR U40199 ( .A(y[3726]), .B(x[3726]), .Z(n31317) );
  XOR U40200 ( .A(n31311), .B(n31310), .Z(n31321) );
  XOR U40201 ( .A(n31313), .B(n31312), .Z(n31310) );
  XOR U40202 ( .A(y[3725]), .B(x[3725]), .Z(n31312) );
  XOR U40203 ( .A(y[3724]), .B(x[3724]), .Z(n31313) );
  XOR U40204 ( .A(y[3723]), .B(x[3723]), .Z(n31311) );
  XNOR U40205 ( .A(n31287), .B(n31288), .Z(n31305) );
  XNOR U40206 ( .A(n31302), .B(n31303), .Z(n31288) );
  XOR U40207 ( .A(n31299), .B(n31298), .Z(n31303) );
  XOR U40208 ( .A(y[3720]), .B(x[3720]), .Z(n31298) );
  XOR U40209 ( .A(n31301), .B(n31300), .Z(n31299) );
  XOR U40210 ( .A(y[3722]), .B(x[3722]), .Z(n31300) );
  XOR U40211 ( .A(y[3721]), .B(x[3721]), .Z(n31301) );
  XOR U40212 ( .A(n31293), .B(n31292), .Z(n31302) );
  XOR U40213 ( .A(n31295), .B(n31294), .Z(n31292) );
  XOR U40214 ( .A(y[3719]), .B(x[3719]), .Z(n31294) );
  XOR U40215 ( .A(y[3718]), .B(x[3718]), .Z(n31295) );
  XOR U40216 ( .A(y[3717]), .B(x[3717]), .Z(n31293) );
  XNOR U40217 ( .A(n31286), .B(n31285), .Z(n31287) );
  XNOR U40218 ( .A(n31282), .B(n31281), .Z(n31285) );
  XOR U40219 ( .A(n31284), .B(n31283), .Z(n31281) );
  XOR U40220 ( .A(y[3716]), .B(x[3716]), .Z(n31283) );
  XOR U40221 ( .A(y[3715]), .B(x[3715]), .Z(n31284) );
  XOR U40222 ( .A(y[3714]), .B(x[3714]), .Z(n31282) );
  XOR U40223 ( .A(n31276), .B(n31275), .Z(n31286) );
  XOR U40224 ( .A(n31278), .B(n31277), .Z(n31275) );
  XOR U40225 ( .A(y[3713]), .B(x[3713]), .Z(n31277) );
  XOR U40226 ( .A(y[3712]), .B(x[3712]), .Z(n31278) );
  XOR U40227 ( .A(y[3711]), .B(x[3711]), .Z(n31276) );
  NAND U40228 ( .A(n31339), .B(n31340), .Z(N62598) );
  NAND U40229 ( .A(n31341), .B(n31342), .Z(n31340) );
  NANDN U40230 ( .A(n31343), .B(n31344), .Z(n31342) );
  NANDN U40231 ( .A(n31344), .B(n31343), .Z(n31339) );
  XOR U40232 ( .A(n31343), .B(n31345), .Z(N62597) );
  XNOR U40233 ( .A(n31341), .B(n31344), .Z(n31345) );
  NAND U40234 ( .A(n31346), .B(n31347), .Z(n31344) );
  NAND U40235 ( .A(n31348), .B(n31349), .Z(n31347) );
  NANDN U40236 ( .A(n31350), .B(n31351), .Z(n31349) );
  NANDN U40237 ( .A(n31351), .B(n31350), .Z(n31346) );
  AND U40238 ( .A(n31352), .B(n31353), .Z(n31341) );
  NAND U40239 ( .A(n31354), .B(n31355), .Z(n31353) );
  NANDN U40240 ( .A(n31356), .B(n31357), .Z(n31355) );
  NANDN U40241 ( .A(n31357), .B(n31356), .Z(n31352) );
  IV U40242 ( .A(n31358), .Z(n31357) );
  AND U40243 ( .A(n31359), .B(n31360), .Z(n31343) );
  NAND U40244 ( .A(n31361), .B(n31362), .Z(n31360) );
  NANDN U40245 ( .A(n31363), .B(n31364), .Z(n31362) );
  NANDN U40246 ( .A(n31364), .B(n31363), .Z(n31359) );
  XOR U40247 ( .A(n31356), .B(n31365), .Z(N62596) );
  XNOR U40248 ( .A(n31354), .B(n31358), .Z(n31365) );
  XOR U40249 ( .A(n31351), .B(n31366), .Z(n31358) );
  XNOR U40250 ( .A(n31348), .B(n31350), .Z(n31366) );
  AND U40251 ( .A(n31367), .B(n31368), .Z(n31350) );
  NANDN U40252 ( .A(n31369), .B(n31370), .Z(n31368) );
  OR U40253 ( .A(n31371), .B(n31372), .Z(n31370) );
  IV U40254 ( .A(n31373), .Z(n31372) );
  NANDN U40255 ( .A(n31373), .B(n31371), .Z(n31367) );
  AND U40256 ( .A(n31374), .B(n31375), .Z(n31348) );
  NAND U40257 ( .A(n31376), .B(n31377), .Z(n31375) );
  NANDN U40258 ( .A(n31378), .B(n31379), .Z(n31377) );
  NANDN U40259 ( .A(n31379), .B(n31378), .Z(n31374) );
  IV U40260 ( .A(n31380), .Z(n31379) );
  NAND U40261 ( .A(n31381), .B(n31382), .Z(n31351) );
  NANDN U40262 ( .A(n31383), .B(n31384), .Z(n31382) );
  NANDN U40263 ( .A(n31385), .B(n31386), .Z(n31384) );
  NANDN U40264 ( .A(n31386), .B(n31385), .Z(n31381) );
  IV U40265 ( .A(n31387), .Z(n31385) );
  AND U40266 ( .A(n31388), .B(n31389), .Z(n31354) );
  NAND U40267 ( .A(n31390), .B(n31391), .Z(n31389) );
  NANDN U40268 ( .A(n31392), .B(n31393), .Z(n31391) );
  NANDN U40269 ( .A(n31393), .B(n31392), .Z(n31388) );
  XOR U40270 ( .A(n31364), .B(n31394), .Z(n31356) );
  XNOR U40271 ( .A(n31361), .B(n31363), .Z(n31394) );
  AND U40272 ( .A(n31395), .B(n31396), .Z(n31363) );
  NANDN U40273 ( .A(n31397), .B(n31398), .Z(n31396) );
  OR U40274 ( .A(n31399), .B(n31400), .Z(n31398) );
  IV U40275 ( .A(n31401), .Z(n31400) );
  NANDN U40276 ( .A(n31401), .B(n31399), .Z(n31395) );
  AND U40277 ( .A(n31402), .B(n31403), .Z(n31361) );
  NAND U40278 ( .A(n31404), .B(n31405), .Z(n31403) );
  NANDN U40279 ( .A(n31406), .B(n31407), .Z(n31405) );
  NANDN U40280 ( .A(n31407), .B(n31406), .Z(n31402) );
  IV U40281 ( .A(n31408), .Z(n31407) );
  NAND U40282 ( .A(n31409), .B(n31410), .Z(n31364) );
  NANDN U40283 ( .A(n31411), .B(n31412), .Z(n31410) );
  NANDN U40284 ( .A(n31413), .B(n31414), .Z(n31412) );
  NANDN U40285 ( .A(n31414), .B(n31413), .Z(n31409) );
  IV U40286 ( .A(n31415), .Z(n31413) );
  XOR U40287 ( .A(n31390), .B(n31416), .Z(N62595) );
  XNOR U40288 ( .A(n31393), .B(n31392), .Z(n31416) );
  XNOR U40289 ( .A(n31404), .B(n31417), .Z(n31392) );
  XNOR U40290 ( .A(n31408), .B(n31406), .Z(n31417) );
  XOR U40291 ( .A(n31414), .B(n31418), .Z(n31406) );
  XNOR U40292 ( .A(n31411), .B(n31415), .Z(n31418) );
  AND U40293 ( .A(n31419), .B(n31420), .Z(n31415) );
  NAND U40294 ( .A(n31421), .B(n31422), .Z(n31420) );
  NAND U40295 ( .A(n31423), .B(n31424), .Z(n31419) );
  AND U40296 ( .A(n31425), .B(n31426), .Z(n31411) );
  NAND U40297 ( .A(n31427), .B(n31428), .Z(n31426) );
  NAND U40298 ( .A(n31429), .B(n31430), .Z(n31425) );
  NANDN U40299 ( .A(n31431), .B(n31432), .Z(n31414) );
  ANDN U40300 ( .B(n31433), .A(n31434), .Z(n31408) );
  XNOR U40301 ( .A(n31399), .B(n31435), .Z(n31404) );
  XNOR U40302 ( .A(n31397), .B(n31401), .Z(n31435) );
  AND U40303 ( .A(n31436), .B(n31437), .Z(n31401) );
  NAND U40304 ( .A(n31438), .B(n31439), .Z(n31437) );
  NAND U40305 ( .A(n31440), .B(n31441), .Z(n31436) );
  AND U40306 ( .A(n31442), .B(n31443), .Z(n31397) );
  NAND U40307 ( .A(n31444), .B(n31445), .Z(n31443) );
  NAND U40308 ( .A(n31446), .B(n31447), .Z(n31442) );
  AND U40309 ( .A(n31448), .B(n31449), .Z(n31399) );
  NAND U40310 ( .A(n31450), .B(n31451), .Z(n31393) );
  XNOR U40311 ( .A(n31376), .B(n31452), .Z(n31390) );
  XNOR U40312 ( .A(n31380), .B(n31378), .Z(n31452) );
  XOR U40313 ( .A(n31386), .B(n31453), .Z(n31378) );
  XNOR U40314 ( .A(n31383), .B(n31387), .Z(n31453) );
  AND U40315 ( .A(n31454), .B(n31455), .Z(n31387) );
  NAND U40316 ( .A(n31456), .B(n31457), .Z(n31455) );
  NAND U40317 ( .A(n31458), .B(n31459), .Z(n31454) );
  AND U40318 ( .A(n31460), .B(n31461), .Z(n31383) );
  NAND U40319 ( .A(n31462), .B(n31463), .Z(n31461) );
  NAND U40320 ( .A(n31464), .B(n31465), .Z(n31460) );
  NANDN U40321 ( .A(n31466), .B(n31467), .Z(n31386) );
  ANDN U40322 ( .B(n31468), .A(n31469), .Z(n31380) );
  XNOR U40323 ( .A(n31371), .B(n31470), .Z(n31376) );
  XNOR U40324 ( .A(n31369), .B(n31373), .Z(n31470) );
  AND U40325 ( .A(n31471), .B(n31472), .Z(n31373) );
  NAND U40326 ( .A(n31473), .B(n31474), .Z(n31472) );
  NAND U40327 ( .A(n31475), .B(n31476), .Z(n31471) );
  AND U40328 ( .A(n31477), .B(n31478), .Z(n31369) );
  NAND U40329 ( .A(n31479), .B(n31480), .Z(n31478) );
  NAND U40330 ( .A(n31481), .B(n31482), .Z(n31477) );
  AND U40331 ( .A(n31483), .B(n31484), .Z(n31371) );
  XOR U40332 ( .A(n31451), .B(n31450), .Z(N62594) );
  XNOR U40333 ( .A(n31468), .B(n31469), .Z(n31450) );
  XNOR U40334 ( .A(n31483), .B(n31484), .Z(n31469) );
  XOR U40335 ( .A(n31480), .B(n31479), .Z(n31484) );
  XOR U40336 ( .A(y[3708]), .B(x[3708]), .Z(n31479) );
  XOR U40337 ( .A(n31482), .B(n31481), .Z(n31480) );
  XOR U40338 ( .A(y[3710]), .B(x[3710]), .Z(n31481) );
  XOR U40339 ( .A(y[3709]), .B(x[3709]), .Z(n31482) );
  XOR U40340 ( .A(n31474), .B(n31473), .Z(n31483) );
  XOR U40341 ( .A(n31476), .B(n31475), .Z(n31473) );
  XOR U40342 ( .A(y[3707]), .B(x[3707]), .Z(n31475) );
  XOR U40343 ( .A(y[3706]), .B(x[3706]), .Z(n31476) );
  XOR U40344 ( .A(y[3705]), .B(x[3705]), .Z(n31474) );
  XNOR U40345 ( .A(n31467), .B(n31466), .Z(n31468) );
  XNOR U40346 ( .A(n31463), .B(n31462), .Z(n31466) );
  XOR U40347 ( .A(n31465), .B(n31464), .Z(n31462) );
  XOR U40348 ( .A(y[3704]), .B(x[3704]), .Z(n31464) );
  XOR U40349 ( .A(y[3703]), .B(x[3703]), .Z(n31465) );
  XOR U40350 ( .A(y[3702]), .B(x[3702]), .Z(n31463) );
  XOR U40351 ( .A(n31457), .B(n31456), .Z(n31467) );
  XOR U40352 ( .A(n31459), .B(n31458), .Z(n31456) );
  XOR U40353 ( .A(y[3701]), .B(x[3701]), .Z(n31458) );
  XOR U40354 ( .A(y[3700]), .B(x[3700]), .Z(n31459) );
  XOR U40355 ( .A(y[3699]), .B(x[3699]), .Z(n31457) );
  XNOR U40356 ( .A(n31433), .B(n31434), .Z(n31451) );
  XNOR U40357 ( .A(n31448), .B(n31449), .Z(n31434) );
  XOR U40358 ( .A(n31445), .B(n31444), .Z(n31449) );
  XOR U40359 ( .A(y[3696]), .B(x[3696]), .Z(n31444) );
  XOR U40360 ( .A(n31447), .B(n31446), .Z(n31445) );
  XOR U40361 ( .A(y[3698]), .B(x[3698]), .Z(n31446) );
  XOR U40362 ( .A(y[3697]), .B(x[3697]), .Z(n31447) );
  XOR U40363 ( .A(n31439), .B(n31438), .Z(n31448) );
  XOR U40364 ( .A(n31441), .B(n31440), .Z(n31438) );
  XOR U40365 ( .A(y[3695]), .B(x[3695]), .Z(n31440) );
  XOR U40366 ( .A(y[3694]), .B(x[3694]), .Z(n31441) );
  XOR U40367 ( .A(y[3693]), .B(x[3693]), .Z(n31439) );
  XNOR U40368 ( .A(n31432), .B(n31431), .Z(n31433) );
  XNOR U40369 ( .A(n31428), .B(n31427), .Z(n31431) );
  XOR U40370 ( .A(n31430), .B(n31429), .Z(n31427) );
  XOR U40371 ( .A(y[3692]), .B(x[3692]), .Z(n31429) );
  XOR U40372 ( .A(y[3691]), .B(x[3691]), .Z(n31430) );
  XOR U40373 ( .A(y[3690]), .B(x[3690]), .Z(n31428) );
  XOR U40374 ( .A(n31422), .B(n31421), .Z(n31432) );
  XOR U40375 ( .A(n31424), .B(n31423), .Z(n31421) );
  XOR U40376 ( .A(y[3689]), .B(x[3689]), .Z(n31423) );
  XOR U40377 ( .A(y[3688]), .B(x[3688]), .Z(n31424) );
  XOR U40378 ( .A(y[3687]), .B(x[3687]), .Z(n31422) );
  NAND U40379 ( .A(n31485), .B(n31486), .Z(N62585) );
  NAND U40380 ( .A(n31487), .B(n31488), .Z(n31486) );
  NANDN U40381 ( .A(n31489), .B(n31490), .Z(n31488) );
  NANDN U40382 ( .A(n31490), .B(n31489), .Z(n31485) );
  XOR U40383 ( .A(n31489), .B(n31491), .Z(N62584) );
  XNOR U40384 ( .A(n31487), .B(n31490), .Z(n31491) );
  NAND U40385 ( .A(n31492), .B(n31493), .Z(n31490) );
  NAND U40386 ( .A(n31494), .B(n31495), .Z(n31493) );
  NANDN U40387 ( .A(n31496), .B(n31497), .Z(n31495) );
  NANDN U40388 ( .A(n31497), .B(n31496), .Z(n31492) );
  AND U40389 ( .A(n31498), .B(n31499), .Z(n31487) );
  NAND U40390 ( .A(n31500), .B(n31501), .Z(n31499) );
  NANDN U40391 ( .A(n31502), .B(n31503), .Z(n31501) );
  NANDN U40392 ( .A(n31503), .B(n31502), .Z(n31498) );
  IV U40393 ( .A(n31504), .Z(n31503) );
  AND U40394 ( .A(n31505), .B(n31506), .Z(n31489) );
  NAND U40395 ( .A(n31507), .B(n31508), .Z(n31506) );
  NANDN U40396 ( .A(n31509), .B(n31510), .Z(n31508) );
  NANDN U40397 ( .A(n31510), .B(n31509), .Z(n31505) );
  XOR U40398 ( .A(n31502), .B(n31511), .Z(N62583) );
  XNOR U40399 ( .A(n31500), .B(n31504), .Z(n31511) );
  XOR U40400 ( .A(n31497), .B(n31512), .Z(n31504) );
  XNOR U40401 ( .A(n31494), .B(n31496), .Z(n31512) );
  AND U40402 ( .A(n31513), .B(n31514), .Z(n31496) );
  NANDN U40403 ( .A(n31515), .B(n31516), .Z(n31514) );
  OR U40404 ( .A(n31517), .B(n31518), .Z(n31516) );
  IV U40405 ( .A(n31519), .Z(n31518) );
  NANDN U40406 ( .A(n31519), .B(n31517), .Z(n31513) );
  AND U40407 ( .A(n31520), .B(n31521), .Z(n31494) );
  NAND U40408 ( .A(n31522), .B(n31523), .Z(n31521) );
  NANDN U40409 ( .A(n31524), .B(n31525), .Z(n31523) );
  NANDN U40410 ( .A(n31525), .B(n31524), .Z(n31520) );
  IV U40411 ( .A(n31526), .Z(n31525) );
  NAND U40412 ( .A(n31527), .B(n31528), .Z(n31497) );
  NANDN U40413 ( .A(n31529), .B(n31530), .Z(n31528) );
  NANDN U40414 ( .A(n31531), .B(n31532), .Z(n31530) );
  NANDN U40415 ( .A(n31532), .B(n31531), .Z(n31527) );
  IV U40416 ( .A(n31533), .Z(n31531) );
  AND U40417 ( .A(n31534), .B(n31535), .Z(n31500) );
  NAND U40418 ( .A(n31536), .B(n31537), .Z(n31535) );
  NANDN U40419 ( .A(n31538), .B(n31539), .Z(n31537) );
  NANDN U40420 ( .A(n31539), .B(n31538), .Z(n31534) );
  XOR U40421 ( .A(n31510), .B(n31540), .Z(n31502) );
  XNOR U40422 ( .A(n31507), .B(n31509), .Z(n31540) );
  AND U40423 ( .A(n31541), .B(n31542), .Z(n31509) );
  NANDN U40424 ( .A(n31543), .B(n31544), .Z(n31542) );
  OR U40425 ( .A(n31545), .B(n31546), .Z(n31544) );
  IV U40426 ( .A(n31547), .Z(n31546) );
  NANDN U40427 ( .A(n31547), .B(n31545), .Z(n31541) );
  AND U40428 ( .A(n31548), .B(n31549), .Z(n31507) );
  NAND U40429 ( .A(n31550), .B(n31551), .Z(n31549) );
  NANDN U40430 ( .A(n31552), .B(n31553), .Z(n31551) );
  NANDN U40431 ( .A(n31553), .B(n31552), .Z(n31548) );
  IV U40432 ( .A(n31554), .Z(n31553) );
  NAND U40433 ( .A(n31555), .B(n31556), .Z(n31510) );
  NANDN U40434 ( .A(n31557), .B(n31558), .Z(n31556) );
  NANDN U40435 ( .A(n31559), .B(n31560), .Z(n31558) );
  NANDN U40436 ( .A(n31560), .B(n31559), .Z(n31555) );
  IV U40437 ( .A(n31561), .Z(n31559) );
  XOR U40438 ( .A(n31536), .B(n31562), .Z(N62582) );
  XNOR U40439 ( .A(n31539), .B(n31538), .Z(n31562) );
  XNOR U40440 ( .A(n31550), .B(n31563), .Z(n31538) );
  XNOR U40441 ( .A(n31554), .B(n31552), .Z(n31563) );
  XOR U40442 ( .A(n31560), .B(n31564), .Z(n31552) );
  XNOR U40443 ( .A(n31557), .B(n31561), .Z(n31564) );
  AND U40444 ( .A(n31565), .B(n31566), .Z(n31561) );
  NAND U40445 ( .A(n31567), .B(n31568), .Z(n31566) );
  NAND U40446 ( .A(n31569), .B(n31570), .Z(n31565) );
  AND U40447 ( .A(n31571), .B(n31572), .Z(n31557) );
  NAND U40448 ( .A(n31573), .B(n31574), .Z(n31572) );
  NAND U40449 ( .A(n31575), .B(n31576), .Z(n31571) );
  NANDN U40450 ( .A(n31577), .B(n31578), .Z(n31560) );
  ANDN U40451 ( .B(n31579), .A(n31580), .Z(n31554) );
  XNOR U40452 ( .A(n31545), .B(n31581), .Z(n31550) );
  XNOR U40453 ( .A(n31543), .B(n31547), .Z(n31581) );
  AND U40454 ( .A(n31582), .B(n31583), .Z(n31547) );
  NAND U40455 ( .A(n31584), .B(n31585), .Z(n31583) );
  NAND U40456 ( .A(n31586), .B(n31587), .Z(n31582) );
  AND U40457 ( .A(n31588), .B(n31589), .Z(n31543) );
  NAND U40458 ( .A(n31590), .B(n31591), .Z(n31589) );
  NAND U40459 ( .A(n31592), .B(n31593), .Z(n31588) );
  AND U40460 ( .A(n31594), .B(n31595), .Z(n31545) );
  NAND U40461 ( .A(n31596), .B(n31597), .Z(n31539) );
  XNOR U40462 ( .A(n31522), .B(n31598), .Z(n31536) );
  XNOR U40463 ( .A(n31526), .B(n31524), .Z(n31598) );
  XOR U40464 ( .A(n31532), .B(n31599), .Z(n31524) );
  XNOR U40465 ( .A(n31529), .B(n31533), .Z(n31599) );
  AND U40466 ( .A(n31600), .B(n31601), .Z(n31533) );
  NAND U40467 ( .A(n31602), .B(n31603), .Z(n31601) );
  NAND U40468 ( .A(n31604), .B(n31605), .Z(n31600) );
  AND U40469 ( .A(n31606), .B(n31607), .Z(n31529) );
  NAND U40470 ( .A(n31608), .B(n31609), .Z(n31607) );
  NAND U40471 ( .A(n31610), .B(n31611), .Z(n31606) );
  NANDN U40472 ( .A(n31612), .B(n31613), .Z(n31532) );
  ANDN U40473 ( .B(n31614), .A(n31615), .Z(n31526) );
  XNOR U40474 ( .A(n31517), .B(n31616), .Z(n31522) );
  XNOR U40475 ( .A(n31515), .B(n31519), .Z(n31616) );
  AND U40476 ( .A(n31617), .B(n31618), .Z(n31519) );
  NAND U40477 ( .A(n31619), .B(n31620), .Z(n31618) );
  NAND U40478 ( .A(n31621), .B(n31622), .Z(n31617) );
  AND U40479 ( .A(n31623), .B(n31624), .Z(n31515) );
  NAND U40480 ( .A(n31625), .B(n31626), .Z(n31624) );
  NAND U40481 ( .A(n31627), .B(n31628), .Z(n31623) );
  AND U40482 ( .A(n31629), .B(n31630), .Z(n31517) );
  XOR U40483 ( .A(n31597), .B(n31596), .Z(N62581) );
  XNOR U40484 ( .A(n31614), .B(n31615), .Z(n31596) );
  XNOR U40485 ( .A(n31629), .B(n31630), .Z(n31615) );
  XOR U40486 ( .A(n31626), .B(n31625), .Z(n31630) );
  XOR U40487 ( .A(y[3684]), .B(x[3684]), .Z(n31625) );
  XOR U40488 ( .A(n31628), .B(n31627), .Z(n31626) );
  XOR U40489 ( .A(y[3686]), .B(x[3686]), .Z(n31627) );
  XOR U40490 ( .A(y[3685]), .B(x[3685]), .Z(n31628) );
  XOR U40491 ( .A(n31620), .B(n31619), .Z(n31629) );
  XOR U40492 ( .A(n31622), .B(n31621), .Z(n31619) );
  XOR U40493 ( .A(y[3683]), .B(x[3683]), .Z(n31621) );
  XOR U40494 ( .A(y[3682]), .B(x[3682]), .Z(n31622) );
  XOR U40495 ( .A(y[3681]), .B(x[3681]), .Z(n31620) );
  XNOR U40496 ( .A(n31613), .B(n31612), .Z(n31614) );
  XNOR U40497 ( .A(n31609), .B(n31608), .Z(n31612) );
  XOR U40498 ( .A(n31611), .B(n31610), .Z(n31608) );
  XOR U40499 ( .A(y[3680]), .B(x[3680]), .Z(n31610) );
  XOR U40500 ( .A(y[3679]), .B(x[3679]), .Z(n31611) );
  XOR U40501 ( .A(y[3678]), .B(x[3678]), .Z(n31609) );
  XOR U40502 ( .A(n31603), .B(n31602), .Z(n31613) );
  XOR U40503 ( .A(n31605), .B(n31604), .Z(n31602) );
  XOR U40504 ( .A(y[3677]), .B(x[3677]), .Z(n31604) );
  XOR U40505 ( .A(y[3676]), .B(x[3676]), .Z(n31605) );
  XOR U40506 ( .A(y[3675]), .B(x[3675]), .Z(n31603) );
  XNOR U40507 ( .A(n31579), .B(n31580), .Z(n31597) );
  XNOR U40508 ( .A(n31594), .B(n31595), .Z(n31580) );
  XOR U40509 ( .A(n31591), .B(n31590), .Z(n31595) );
  XOR U40510 ( .A(y[3672]), .B(x[3672]), .Z(n31590) );
  XOR U40511 ( .A(n31593), .B(n31592), .Z(n31591) );
  XOR U40512 ( .A(y[3674]), .B(x[3674]), .Z(n31592) );
  XOR U40513 ( .A(y[3673]), .B(x[3673]), .Z(n31593) );
  XOR U40514 ( .A(n31585), .B(n31584), .Z(n31594) );
  XOR U40515 ( .A(n31587), .B(n31586), .Z(n31584) );
  XOR U40516 ( .A(y[3671]), .B(x[3671]), .Z(n31586) );
  XOR U40517 ( .A(y[3670]), .B(x[3670]), .Z(n31587) );
  XOR U40518 ( .A(y[3669]), .B(x[3669]), .Z(n31585) );
  XNOR U40519 ( .A(n31578), .B(n31577), .Z(n31579) );
  XNOR U40520 ( .A(n31574), .B(n31573), .Z(n31577) );
  XOR U40521 ( .A(n31576), .B(n31575), .Z(n31573) );
  XOR U40522 ( .A(y[3668]), .B(x[3668]), .Z(n31575) );
  XOR U40523 ( .A(y[3667]), .B(x[3667]), .Z(n31576) );
  XOR U40524 ( .A(y[3666]), .B(x[3666]), .Z(n31574) );
  XOR U40525 ( .A(n31568), .B(n31567), .Z(n31578) );
  XOR U40526 ( .A(n31570), .B(n31569), .Z(n31567) );
  XOR U40527 ( .A(y[3665]), .B(x[3665]), .Z(n31569) );
  XOR U40528 ( .A(y[3664]), .B(x[3664]), .Z(n31570) );
  XOR U40529 ( .A(y[3663]), .B(x[3663]), .Z(n31568) );
  NAND U40530 ( .A(n31631), .B(n31632), .Z(N62572) );
  NAND U40531 ( .A(n31633), .B(n31634), .Z(n31632) );
  NANDN U40532 ( .A(n31635), .B(n31636), .Z(n31634) );
  NANDN U40533 ( .A(n31636), .B(n31635), .Z(n31631) );
  XOR U40534 ( .A(n31635), .B(n31637), .Z(N62571) );
  XNOR U40535 ( .A(n31633), .B(n31636), .Z(n31637) );
  NAND U40536 ( .A(n31638), .B(n31639), .Z(n31636) );
  NAND U40537 ( .A(n31640), .B(n31641), .Z(n31639) );
  NANDN U40538 ( .A(n31642), .B(n31643), .Z(n31641) );
  NANDN U40539 ( .A(n31643), .B(n31642), .Z(n31638) );
  AND U40540 ( .A(n31644), .B(n31645), .Z(n31633) );
  NAND U40541 ( .A(n31646), .B(n31647), .Z(n31645) );
  NANDN U40542 ( .A(n31648), .B(n31649), .Z(n31647) );
  NANDN U40543 ( .A(n31649), .B(n31648), .Z(n31644) );
  IV U40544 ( .A(n31650), .Z(n31649) );
  AND U40545 ( .A(n31651), .B(n31652), .Z(n31635) );
  NAND U40546 ( .A(n31653), .B(n31654), .Z(n31652) );
  NANDN U40547 ( .A(n31655), .B(n31656), .Z(n31654) );
  NANDN U40548 ( .A(n31656), .B(n31655), .Z(n31651) );
  XOR U40549 ( .A(n31648), .B(n31657), .Z(N62570) );
  XNOR U40550 ( .A(n31646), .B(n31650), .Z(n31657) );
  XOR U40551 ( .A(n31643), .B(n31658), .Z(n31650) );
  XNOR U40552 ( .A(n31640), .B(n31642), .Z(n31658) );
  AND U40553 ( .A(n31659), .B(n31660), .Z(n31642) );
  NANDN U40554 ( .A(n31661), .B(n31662), .Z(n31660) );
  OR U40555 ( .A(n31663), .B(n31664), .Z(n31662) );
  IV U40556 ( .A(n31665), .Z(n31664) );
  NANDN U40557 ( .A(n31665), .B(n31663), .Z(n31659) );
  AND U40558 ( .A(n31666), .B(n31667), .Z(n31640) );
  NAND U40559 ( .A(n31668), .B(n31669), .Z(n31667) );
  NANDN U40560 ( .A(n31670), .B(n31671), .Z(n31669) );
  NANDN U40561 ( .A(n31671), .B(n31670), .Z(n31666) );
  IV U40562 ( .A(n31672), .Z(n31671) );
  NAND U40563 ( .A(n31673), .B(n31674), .Z(n31643) );
  NANDN U40564 ( .A(n31675), .B(n31676), .Z(n31674) );
  NANDN U40565 ( .A(n31677), .B(n31678), .Z(n31676) );
  NANDN U40566 ( .A(n31678), .B(n31677), .Z(n31673) );
  IV U40567 ( .A(n31679), .Z(n31677) );
  AND U40568 ( .A(n31680), .B(n31681), .Z(n31646) );
  NAND U40569 ( .A(n31682), .B(n31683), .Z(n31681) );
  NANDN U40570 ( .A(n31684), .B(n31685), .Z(n31683) );
  NANDN U40571 ( .A(n31685), .B(n31684), .Z(n31680) );
  XOR U40572 ( .A(n31656), .B(n31686), .Z(n31648) );
  XNOR U40573 ( .A(n31653), .B(n31655), .Z(n31686) );
  AND U40574 ( .A(n31687), .B(n31688), .Z(n31655) );
  NANDN U40575 ( .A(n31689), .B(n31690), .Z(n31688) );
  OR U40576 ( .A(n31691), .B(n31692), .Z(n31690) );
  IV U40577 ( .A(n31693), .Z(n31692) );
  NANDN U40578 ( .A(n31693), .B(n31691), .Z(n31687) );
  AND U40579 ( .A(n31694), .B(n31695), .Z(n31653) );
  NAND U40580 ( .A(n31696), .B(n31697), .Z(n31695) );
  NANDN U40581 ( .A(n31698), .B(n31699), .Z(n31697) );
  NANDN U40582 ( .A(n31699), .B(n31698), .Z(n31694) );
  IV U40583 ( .A(n31700), .Z(n31699) );
  NAND U40584 ( .A(n31701), .B(n31702), .Z(n31656) );
  NANDN U40585 ( .A(n31703), .B(n31704), .Z(n31702) );
  NANDN U40586 ( .A(n31705), .B(n31706), .Z(n31704) );
  NANDN U40587 ( .A(n31706), .B(n31705), .Z(n31701) );
  IV U40588 ( .A(n31707), .Z(n31705) );
  XOR U40589 ( .A(n31682), .B(n31708), .Z(N62569) );
  XNOR U40590 ( .A(n31685), .B(n31684), .Z(n31708) );
  XNOR U40591 ( .A(n31696), .B(n31709), .Z(n31684) );
  XNOR U40592 ( .A(n31700), .B(n31698), .Z(n31709) );
  XOR U40593 ( .A(n31706), .B(n31710), .Z(n31698) );
  XNOR U40594 ( .A(n31703), .B(n31707), .Z(n31710) );
  AND U40595 ( .A(n31711), .B(n31712), .Z(n31707) );
  NAND U40596 ( .A(n31713), .B(n31714), .Z(n31712) );
  NAND U40597 ( .A(n31715), .B(n31716), .Z(n31711) );
  AND U40598 ( .A(n31717), .B(n31718), .Z(n31703) );
  NAND U40599 ( .A(n31719), .B(n31720), .Z(n31718) );
  NAND U40600 ( .A(n31721), .B(n31722), .Z(n31717) );
  NANDN U40601 ( .A(n31723), .B(n31724), .Z(n31706) );
  ANDN U40602 ( .B(n31725), .A(n31726), .Z(n31700) );
  XNOR U40603 ( .A(n31691), .B(n31727), .Z(n31696) );
  XNOR U40604 ( .A(n31689), .B(n31693), .Z(n31727) );
  AND U40605 ( .A(n31728), .B(n31729), .Z(n31693) );
  NAND U40606 ( .A(n31730), .B(n31731), .Z(n31729) );
  NAND U40607 ( .A(n31732), .B(n31733), .Z(n31728) );
  AND U40608 ( .A(n31734), .B(n31735), .Z(n31689) );
  NAND U40609 ( .A(n31736), .B(n31737), .Z(n31735) );
  NAND U40610 ( .A(n31738), .B(n31739), .Z(n31734) );
  AND U40611 ( .A(n31740), .B(n31741), .Z(n31691) );
  NAND U40612 ( .A(n31742), .B(n31743), .Z(n31685) );
  XNOR U40613 ( .A(n31668), .B(n31744), .Z(n31682) );
  XNOR U40614 ( .A(n31672), .B(n31670), .Z(n31744) );
  XOR U40615 ( .A(n31678), .B(n31745), .Z(n31670) );
  XNOR U40616 ( .A(n31675), .B(n31679), .Z(n31745) );
  AND U40617 ( .A(n31746), .B(n31747), .Z(n31679) );
  NAND U40618 ( .A(n31748), .B(n31749), .Z(n31747) );
  NAND U40619 ( .A(n31750), .B(n31751), .Z(n31746) );
  AND U40620 ( .A(n31752), .B(n31753), .Z(n31675) );
  NAND U40621 ( .A(n31754), .B(n31755), .Z(n31753) );
  NAND U40622 ( .A(n31756), .B(n31757), .Z(n31752) );
  NANDN U40623 ( .A(n31758), .B(n31759), .Z(n31678) );
  ANDN U40624 ( .B(n31760), .A(n31761), .Z(n31672) );
  XNOR U40625 ( .A(n31663), .B(n31762), .Z(n31668) );
  XNOR U40626 ( .A(n31661), .B(n31665), .Z(n31762) );
  AND U40627 ( .A(n31763), .B(n31764), .Z(n31665) );
  NAND U40628 ( .A(n31765), .B(n31766), .Z(n31764) );
  NAND U40629 ( .A(n31767), .B(n31768), .Z(n31763) );
  AND U40630 ( .A(n31769), .B(n31770), .Z(n31661) );
  NAND U40631 ( .A(n31771), .B(n31772), .Z(n31770) );
  NAND U40632 ( .A(n31773), .B(n31774), .Z(n31769) );
  AND U40633 ( .A(n31775), .B(n31776), .Z(n31663) );
  XOR U40634 ( .A(n31743), .B(n31742), .Z(N62568) );
  XNOR U40635 ( .A(n31760), .B(n31761), .Z(n31742) );
  XNOR U40636 ( .A(n31775), .B(n31776), .Z(n31761) );
  XOR U40637 ( .A(n31772), .B(n31771), .Z(n31776) );
  XOR U40638 ( .A(y[3660]), .B(x[3660]), .Z(n31771) );
  XOR U40639 ( .A(n31774), .B(n31773), .Z(n31772) );
  XOR U40640 ( .A(y[3662]), .B(x[3662]), .Z(n31773) );
  XOR U40641 ( .A(y[3661]), .B(x[3661]), .Z(n31774) );
  XOR U40642 ( .A(n31766), .B(n31765), .Z(n31775) );
  XOR U40643 ( .A(n31768), .B(n31767), .Z(n31765) );
  XOR U40644 ( .A(y[3659]), .B(x[3659]), .Z(n31767) );
  XOR U40645 ( .A(y[3658]), .B(x[3658]), .Z(n31768) );
  XOR U40646 ( .A(y[3657]), .B(x[3657]), .Z(n31766) );
  XNOR U40647 ( .A(n31759), .B(n31758), .Z(n31760) );
  XNOR U40648 ( .A(n31755), .B(n31754), .Z(n31758) );
  XOR U40649 ( .A(n31757), .B(n31756), .Z(n31754) );
  XOR U40650 ( .A(y[3656]), .B(x[3656]), .Z(n31756) );
  XOR U40651 ( .A(y[3655]), .B(x[3655]), .Z(n31757) );
  XOR U40652 ( .A(y[3654]), .B(x[3654]), .Z(n31755) );
  XOR U40653 ( .A(n31749), .B(n31748), .Z(n31759) );
  XOR U40654 ( .A(n31751), .B(n31750), .Z(n31748) );
  XOR U40655 ( .A(y[3653]), .B(x[3653]), .Z(n31750) );
  XOR U40656 ( .A(y[3652]), .B(x[3652]), .Z(n31751) );
  XOR U40657 ( .A(y[3651]), .B(x[3651]), .Z(n31749) );
  XNOR U40658 ( .A(n31725), .B(n31726), .Z(n31743) );
  XNOR U40659 ( .A(n31740), .B(n31741), .Z(n31726) );
  XOR U40660 ( .A(n31737), .B(n31736), .Z(n31741) );
  XOR U40661 ( .A(y[3648]), .B(x[3648]), .Z(n31736) );
  XOR U40662 ( .A(n31739), .B(n31738), .Z(n31737) );
  XOR U40663 ( .A(y[3650]), .B(x[3650]), .Z(n31738) );
  XOR U40664 ( .A(y[3649]), .B(x[3649]), .Z(n31739) );
  XOR U40665 ( .A(n31731), .B(n31730), .Z(n31740) );
  XOR U40666 ( .A(n31733), .B(n31732), .Z(n31730) );
  XOR U40667 ( .A(y[3647]), .B(x[3647]), .Z(n31732) );
  XOR U40668 ( .A(y[3646]), .B(x[3646]), .Z(n31733) );
  XOR U40669 ( .A(y[3645]), .B(x[3645]), .Z(n31731) );
  XNOR U40670 ( .A(n31724), .B(n31723), .Z(n31725) );
  XNOR U40671 ( .A(n31720), .B(n31719), .Z(n31723) );
  XOR U40672 ( .A(n31722), .B(n31721), .Z(n31719) );
  XOR U40673 ( .A(y[3644]), .B(x[3644]), .Z(n31721) );
  XOR U40674 ( .A(y[3643]), .B(x[3643]), .Z(n31722) );
  XOR U40675 ( .A(y[3642]), .B(x[3642]), .Z(n31720) );
  XOR U40676 ( .A(n31714), .B(n31713), .Z(n31724) );
  XOR U40677 ( .A(n31716), .B(n31715), .Z(n31713) );
  XOR U40678 ( .A(y[3641]), .B(x[3641]), .Z(n31715) );
  XOR U40679 ( .A(y[3640]), .B(x[3640]), .Z(n31716) );
  XOR U40680 ( .A(y[3639]), .B(x[3639]), .Z(n31714) );
  NAND U40681 ( .A(n31777), .B(n31778), .Z(N62559) );
  NAND U40682 ( .A(n31779), .B(n31780), .Z(n31778) );
  NANDN U40683 ( .A(n31781), .B(n31782), .Z(n31780) );
  NANDN U40684 ( .A(n31782), .B(n31781), .Z(n31777) );
  XOR U40685 ( .A(n31781), .B(n31783), .Z(N62558) );
  XNOR U40686 ( .A(n31779), .B(n31782), .Z(n31783) );
  NAND U40687 ( .A(n31784), .B(n31785), .Z(n31782) );
  NAND U40688 ( .A(n31786), .B(n31787), .Z(n31785) );
  NANDN U40689 ( .A(n31788), .B(n31789), .Z(n31787) );
  NANDN U40690 ( .A(n31789), .B(n31788), .Z(n31784) );
  AND U40691 ( .A(n31790), .B(n31791), .Z(n31779) );
  NAND U40692 ( .A(n31792), .B(n31793), .Z(n31791) );
  NANDN U40693 ( .A(n31794), .B(n31795), .Z(n31793) );
  NANDN U40694 ( .A(n31795), .B(n31794), .Z(n31790) );
  IV U40695 ( .A(n31796), .Z(n31795) );
  AND U40696 ( .A(n31797), .B(n31798), .Z(n31781) );
  NAND U40697 ( .A(n31799), .B(n31800), .Z(n31798) );
  NANDN U40698 ( .A(n31801), .B(n31802), .Z(n31800) );
  NANDN U40699 ( .A(n31802), .B(n31801), .Z(n31797) );
  XOR U40700 ( .A(n31794), .B(n31803), .Z(N62557) );
  XNOR U40701 ( .A(n31792), .B(n31796), .Z(n31803) );
  XOR U40702 ( .A(n31789), .B(n31804), .Z(n31796) );
  XNOR U40703 ( .A(n31786), .B(n31788), .Z(n31804) );
  AND U40704 ( .A(n31805), .B(n31806), .Z(n31788) );
  NANDN U40705 ( .A(n31807), .B(n31808), .Z(n31806) );
  OR U40706 ( .A(n31809), .B(n31810), .Z(n31808) );
  IV U40707 ( .A(n31811), .Z(n31810) );
  NANDN U40708 ( .A(n31811), .B(n31809), .Z(n31805) );
  AND U40709 ( .A(n31812), .B(n31813), .Z(n31786) );
  NAND U40710 ( .A(n31814), .B(n31815), .Z(n31813) );
  NANDN U40711 ( .A(n31816), .B(n31817), .Z(n31815) );
  NANDN U40712 ( .A(n31817), .B(n31816), .Z(n31812) );
  IV U40713 ( .A(n31818), .Z(n31817) );
  NAND U40714 ( .A(n31819), .B(n31820), .Z(n31789) );
  NANDN U40715 ( .A(n31821), .B(n31822), .Z(n31820) );
  NANDN U40716 ( .A(n31823), .B(n31824), .Z(n31822) );
  NANDN U40717 ( .A(n31824), .B(n31823), .Z(n31819) );
  IV U40718 ( .A(n31825), .Z(n31823) );
  AND U40719 ( .A(n31826), .B(n31827), .Z(n31792) );
  NAND U40720 ( .A(n31828), .B(n31829), .Z(n31827) );
  NANDN U40721 ( .A(n31830), .B(n31831), .Z(n31829) );
  NANDN U40722 ( .A(n31831), .B(n31830), .Z(n31826) );
  XOR U40723 ( .A(n31802), .B(n31832), .Z(n31794) );
  XNOR U40724 ( .A(n31799), .B(n31801), .Z(n31832) );
  AND U40725 ( .A(n31833), .B(n31834), .Z(n31801) );
  NANDN U40726 ( .A(n31835), .B(n31836), .Z(n31834) );
  OR U40727 ( .A(n31837), .B(n31838), .Z(n31836) );
  IV U40728 ( .A(n31839), .Z(n31838) );
  NANDN U40729 ( .A(n31839), .B(n31837), .Z(n31833) );
  AND U40730 ( .A(n31840), .B(n31841), .Z(n31799) );
  NAND U40731 ( .A(n31842), .B(n31843), .Z(n31841) );
  NANDN U40732 ( .A(n31844), .B(n31845), .Z(n31843) );
  NANDN U40733 ( .A(n31845), .B(n31844), .Z(n31840) );
  IV U40734 ( .A(n31846), .Z(n31845) );
  NAND U40735 ( .A(n31847), .B(n31848), .Z(n31802) );
  NANDN U40736 ( .A(n31849), .B(n31850), .Z(n31848) );
  NANDN U40737 ( .A(n31851), .B(n31852), .Z(n31850) );
  NANDN U40738 ( .A(n31852), .B(n31851), .Z(n31847) );
  IV U40739 ( .A(n31853), .Z(n31851) );
  XOR U40740 ( .A(n31828), .B(n31854), .Z(N62556) );
  XNOR U40741 ( .A(n31831), .B(n31830), .Z(n31854) );
  XNOR U40742 ( .A(n31842), .B(n31855), .Z(n31830) );
  XNOR U40743 ( .A(n31846), .B(n31844), .Z(n31855) );
  XOR U40744 ( .A(n31852), .B(n31856), .Z(n31844) );
  XNOR U40745 ( .A(n31849), .B(n31853), .Z(n31856) );
  AND U40746 ( .A(n31857), .B(n31858), .Z(n31853) );
  NAND U40747 ( .A(n31859), .B(n31860), .Z(n31858) );
  NAND U40748 ( .A(n31861), .B(n31862), .Z(n31857) );
  AND U40749 ( .A(n31863), .B(n31864), .Z(n31849) );
  NAND U40750 ( .A(n31865), .B(n31866), .Z(n31864) );
  NAND U40751 ( .A(n31867), .B(n31868), .Z(n31863) );
  NANDN U40752 ( .A(n31869), .B(n31870), .Z(n31852) );
  ANDN U40753 ( .B(n31871), .A(n31872), .Z(n31846) );
  XNOR U40754 ( .A(n31837), .B(n31873), .Z(n31842) );
  XNOR U40755 ( .A(n31835), .B(n31839), .Z(n31873) );
  AND U40756 ( .A(n31874), .B(n31875), .Z(n31839) );
  NAND U40757 ( .A(n31876), .B(n31877), .Z(n31875) );
  NAND U40758 ( .A(n31878), .B(n31879), .Z(n31874) );
  AND U40759 ( .A(n31880), .B(n31881), .Z(n31835) );
  NAND U40760 ( .A(n31882), .B(n31883), .Z(n31881) );
  NAND U40761 ( .A(n31884), .B(n31885), .Z(n31880) );
  AND U40762 ( .A(n31886), .B(n31887), .Z(n31837) );
  NAND U40763 ( .A(n31888), .B(n31889), .Z(n31831) );
  XNOR U40764 ( .A(n31814), .B(n31890), .Z(n31828) );
  XNOR U40765 ( .A(n31818), .B(n31816), .Z(n31890) );
  XOR U40766 ( .A(n31824), .B(n31891), .Z(n31816) );
  XNOR U40767 ( .A(n31821), .B(n31825), .Z(n31891) );
  AND U40768 ( .A(n31892), .B(n31893), .Z(n31825) );
  NAND U40769 ( .A(n31894), .B(n31895), .Z(n31893) );
  NAND U40770 ( .A(n31896), .B(n31897), .Z(n31892) );
  AND U40771 ( .A(n31898), .B(n31899), .Z(n31821) );
  NAND U40772 ( .A(n31900), .B(n31901), .Z(n31899) );
  NAND U40773 ( .A(n31902), .B(n31903), .Z(n31898) );
  NANDN U40774 ( .A(n31904), .B(n31905), .Z(n31824) );
  ANDN U40775 ( .B(n31906), .A(n31907), .Z(n31818) );
  XNOR U40776 ( .A(n31809), .B(n31908), .Z(n31814) );
  XNOR U40777 ( .A(n31807), .B(n31811), .Z(n31908) );
  AND U40778 ( .A(n31909), .B(n31910), .Z(n31811) );
  NAND U40779 ( .A(n31911), .B(n31912), .Z(n31910) );
  NAND U40780 ( .A(n31913), .B(n31914), .Z(n31909) );
  AND U40781 ( .A(n31915), .B(n31916), .Z(n31807) );
  NAND U40782 ( .A(n31917), .B(n31918), .Z(n31916) );
  NAND U40783 ( .A(n31919), .B(n31920), .Z(n31915) );
  AND U40784 ( .A(n31921), .B(n31922), .Z(n31809) );
  XOR U40785 ( .A(n31889), .B(n31888), .Z(N62555) );
  XNOR U40786 ( .A(n31906), .B(n31907), .Z(n31888) );
  XNOR U40787 ( .A(n31921), .B(n31922), .Z(n31907) );
  XOR U40788 ( .A(n31918), .B(n31917), .Z(n31922) );
  XOR U40789 ( .A(y[3636]), .B(x[3636]), .Z(n31917) );
  XOR U40790 ( .A(n31920), .B(n31919), .Z(n31918) );
  XOR U40791 ( .A(y[3638]), .B(x[3638]), .Z(n31919) );
  XOR U40792 ( .A(y[3637]), .B(x[3637]), .Z(n31920) );
  XOR U40793 ( .A(n31912), .B(n31911), .Z(n31921) );
  XOR U40794 ( .A(n31914), .B(n31913), .Z(n31911) );
  XOR U40795 ( .A(y[3635]), .B(x[3635]), .Z(n31913) );
  XOR U40796 ( .A(y[3634]), .B(x[3634]), .Z(n31914) );
  XOR U40797 ( .A(y[3633]), .B(x[3633]), .Z(n31912) );
  XNOR U40798 ( .A(n31905), .B(n31904), .Z(n31906) );
  XNOR U40799 ( .A(n31901), .B(n31900), .Z(n31904) );
  XOR U40800 ( .A(n31903), .B(n31902), .Z(n31900) );
  XOR U40801 ( .A(y[3632]), .B(x[3632]), .Z(n31902) );
  XOR U40802 ( .A(y[3631]), .B(x[3631]), .Z(n31903) );
  XOR U40803 ( .A(y[3630]), .B(x[3630]), .Z(n31901) );
  XOR U40804 ( .A(n31895), .B(n31894), .Z(n31905) );
  XOR U40805 ( .A(n31897), .B(n31896), .Z(n31894) );
  XOR U40806 ( .A(y[3629]), .B(x[3629]), .Z(n31896) );
  XOR U40807 ( .A(y[3628]), .B(x[3628]), .Z(n31897) );
  XOR U40808 ( .A(y[3627]), .B(x[3627]), .Z(n31895) );
  XNOR U40809 ( .A(n31871), .B(n31872), .Z(n31889) );
  XNOR U40810 ( .A(n31886), .B(n31887), .Z(n31872) );
  XOR U40811 ( .A(n31883), .B(n31882), .Z(n31887) );
  XOR U40812 ( .A(y[3624]), .B(x[3624]), .Z(n31882) );
  XOR U40813 ( .A(n31885), .B(n31884), .Z(n31883) );
  XOR U40814 ( .A(y[3626]), .B(x[3626]), .Z(n31884) );
  XOR U40815 ( .A(y[3625]), .B(x[3625]), .Z(n31885) );
  XOR U40816 ( .A(n31877), .B(n31876), .Z(n31886) );
  XOR U40817 ( .A(n31879), .B(n31878), .Z(n31876) );
  XOR U40818 ( .A(y[3623]), .B(x[3623]), .Z(n31878) );
  XOR U40819 ( .A(y[3622]), .B(x[3622]), .Z(n31879) );
  XOR U40820 ( .A(y[3621]), .B(x[3621]), .Z(n31877) );
  XNOR U40821 ( .A(n31870), .B(n31869), .Z(n31871) );
  XNOR U40822 ( .A(n31866), .B(n31865), .Z(n31869) );
  XOR U40823 ( .A(n31868), .B(n31867), .Z(n31865) );
  XOR U40824 ( .A(y[3620]), .B(x[3620]), .Z(n31867) );
  XOR U40825 ( .A(y[3619]), .B(x[3619]), .Z(n31868) );
  XOR U40826 ( .A(y[3618]), .B(x[3618]), .Z(n31866) );
  XOR U40827 ( .A(n31860), .B(n31859), .Z(n31870) );
  XOR U40828 ( .A(n31862), .B(n31861), .Z(n31859) );
  XOR U40829 ( .A(y[3617]), .B(x[3617]), .Z(n31861) );
  XOR U40830 ( .A(y[3616]), .B(x[3616]), .Z(n31862) );
  XOR U40831 ( .A(y[3615]), .B(x[3615]), .Z(n31860) );
  NAND U40832 ( .A(n31923), .B(n31924), .Z(N62546) );
  NAND U40833 ( .A(n31925), .B(n31926), .Z(n31924) );
  NANDN U40834 ( .A(n31927), .B(n31928), .Z(n31926) );
  NANDN U40835 ( .A(n31928), .B(n31927), .Z(n31923) );
  XOR U40836 ( .A(n31927), .B(n31929), .Z(N62545) );
  XNOR U40837 ( .A(n31925), .B(n31928), .Z(n31929) );
  NAND U40838 ( .A(n31930), .B(n31931), .Z(n31928) );
  NAND U40839 ( .A(n31932), .B(n31933), .Z(n31931) );
  NANDN U40840 ( .A(n31934), .B(n31935), .Z(n31933) );
  NANDN U40841 ( .A(n31935), .B(n31934), .Z(n31930) );
  AND U40842 ( .A(n31936), .B(n31937), .Z(n31925) );
  NAND U40843 ( .A(n31938), .B(n31939), .Z(n31937) );
  NANDN U40844 ( .A(n31940), .B(n31941), .Z(n31939) );
  NANDN U40845 ( .A(n31941), .B(n31940), .Z(n31936) );
  IV U40846 ( .A(n31942), .Z(n31941) );
  AND U40847 ( .A(n31943), .B(n31944), .Z(n31927) );
  NAND U40848 ( .A(n31945), .B(n31946), .Z(n31944) );
  NANDN U40849 ( .A(n31947), .B(n31948), .Z(n31946) );
  NANDN U40850 ( .A(n31948), .B(n31947), .Z(n31943) );
  XOR U40851 ( .A(n31940), .B(n31949), .Z(N62544) );
  XNOR U40852 ( .A(n31938), .B(n31942), .Z(n31949) );
  XOR U40853 ( .A(n31935), .B(n31950), .Z(n31942) );
  XNOR U40854 ( .A(n31932), .B(n31934), .Z(n31950) );
  AND U40855 ( .A(n31951), .B(n31952), .Z(n31934) );
  NANDN U40856 ( .A(n31953), .B(n31954), .Z(n31952) );
  OR U40857 ( .A(n31955), .B(n31956), .Z(n31954) );
  IV U40858 ( .A(n31957), .Z(n31956) );
  NANDN U40859 ( .A(n31957), .B(n31955), .Z(n31951) );
  AND U40860 ( .A(n31958), .B(n31959), .Z(n31932) );
  NAND U40861 ( .A(n31960), .B(n31961), .Z(n31959) );
  NANDN U40862 ( .A(n31962), .B(n31963), .Z(n31961) );
  NANDN U40863 ( .A(n31963), .B(n31962), .Z(n31958) );
  IV U40864 ( .A(n31964), .Z(n31963) );
  NAND U40865 ( .A(n31965), .B(n31966), .Z(n31935) );
  NANDN U40866 ( .A(n31967), .B(n31968), .Z(n31966) );
  NANDN U40867 ( .A(n31969), .B(n31970), .Z(n31968) );
  NANDN U40868 ( .A(n31970), .B(n31969), .Z(n31965) );
  IV U40869 ( .A(n31971), .Z(n31969) );
  AND U40870 ( .A(n31972), .B(n31973), .Z(n31938) );
  NAND U40871 ( .A(n31974), .B(n31975), .Z(n31973) );
  NANDN U40872 ( .A(n31976), .B(n31977), .Z(n31975) );
  NANDN U40873 ( .A(n31977), .B(n31976), .Z(n31972) );
  XOR U40874 ( .A(n31948), .B(n31978), .Z(n31940) );
  XNOR U40875 ( .A(n31945), .B(n31947), .Z(n31978) );
  AND U40876 ( .A(n31979), .B(n31980), .Z(n31947) );
  NANDN U40877 ( .A(n31981), .B(n31982), .Z(n31980) );
  OR U40878 ( .A(n31983), .B(n31984), .Z(n31982) );
  IV U40879 ( .A(n31985), .Z(n31984) );
  NANDN U40880 ( .A(n31985), .B(n31983), .Z(n31979) );
  AND U40881 ( .A(n31986), .B(n31987), .Z(n31945) );
  NAND U40882 ( .A(n31988), .B(n31989), .Z(n31987) );
  NANDN U40883 ( .A(n31990), .B(n31991), .Z(n31989) );
  NANDN U40884 ( .A(n31991), .B(n31990), .Z(n31986) );
  IV U40885 ( .A(n31992), .Z(n31991) );
  NAND U40886 ( .A(n31993), .B(n31994), .Z(n31948) );
  NANDN U40887 ( .A(n31995), .B(n31996), .Z(n31994) );
  NANDN U40888 ( .A(n31997), .B(n31998), .Z(n31996) );
  NANDN U40889 ( .A(n31998), .B(n31997), .Z(n31993) );
  IV U40890 ( .A(n31999), .Z(n31997) );
  XOR U40891 ( .A(n31974), .B(n32000), .Z(N62543) );
  XNOR U40892 ( .A(n31977), .B(n31976), .Z(n32000) );
  XNOR U40893 ( .A(n31988), .B(n32001), .Z(n31976) );
  XNOR U40894 ( .A(n31992), .B(n31990), .Z(n32001) );
  XOR U40895 ( .A(n31998), .B(n32002), .Z(n31990) );
  XNOR U40896 ( .A(n31995), .B(n31999), .Z(n32002) );
  AND U40897 ( .A(n32003), .B(n32004), .Z(n31999) );
  NAND U40898 ( .A(n32005), .B(n32006), .Z(n32004) );
  NAND U40899 ( .A(n32007), .B(n32008), .Z(n32003) );
  AND U40900 ( .A(n32009), .B(n32010), .Z(n31995) );
  NAND U40901 ( .A(n32011), .B(n32012), .Z(n32010) );
  NAND U40902 ( .A(n32013), .B(n32014), .Z(n32009) );
  NANDN U40903 ( .A(n32015), .B(n32016), .Z(n31998) );
  ANDN U40904 ( .B(n32017), .A(n32018), .Z(n31992) );
  XNOR U40905 ( .A(n31983), .B(n32019), .Z(n31988) );
  XNOR U40906 ( .A(n31981), .B(n31985), .Z(n32019) );
  AND U40907 ( .A(n32020), .B(n32021), .Z(n31985) );
  NAND U40908 ( .A(n32022), .B(n32023), .Z(n32021) );
  NAND U40909 ( .A(n32024), .B(n32025), .Z(n32020) );
  AND U40910 ( .A(n32026), .B(n32027), .Z(n31981) );
  NAND U40911 ( .A(n32028), .B(n32029), .Z(n32027) );
  NAND U40912 ( .A(n32030), .B(n32031), .Z(n32026) );
  AND U40913 ( .A(n32032), .B(n32033), .Z(n31983) );
  NAND U40914 ( .A(n32034), .B(n32035), .Z(n31977) );
  XNOR U40915 ( .A(n31960), .B(n32036), .Z(n31974) );
  XNOR U40916 ( .A(n31964), .B(n31962), .Z(n32036) );
  XOR U40917 ( .A(n31970), .B(n32037), .Z(n31962) );
  XNOR U40918 ( .A(n31967), .B(n31971), .Z(n32037) );
  AND U40919 ( .A(n32038), .B(n32039), .Z(n31971) );
  NAND U40920 ( .A(n32040), .B(n32041), .Z(n32039) );
  NAND U40921 ( .A(n32042), .B(n32043), .Z(n32038) );
  AND U40922 ( .A(n32044), .B(n32045), .Z(n31967) );
  NAND U40923 ( .A(n32046), .B(n32047), .Z(n32045) );
  NAND U40924 ( .A(n32048), .B(n32049), .Z(n32044) );
  NANDN U40925 ( .A(n32050), .B(n32051), .Z(n31970) );
  ANDN U40926 ( .B(n32052), .A(n32053), .Z(n31964) );
  XNOR U40927 ( .A(n31955), .B(n32054), .Z(n31960) );
  XNOR U40928 ( .A(n31953), .B(n31957), .Z(n32054) );
  AND U40929 ( .A(n32055), .B(n32056), .Z(n31957) );
  NAND U40930 ( .A(n32057), .B(n32058), .Z(n32056) );
  NAND U40931 ( .A(n32059), .B(n32060), .Z(n32055) );
  AND U40932 ( .A(n32061), .B(n32062), .Z(n31953) );
  NAND U40933 ( .A(n32063), .B(n32064), .Z(n32062) );
  NAND U40934 ( .A(n32065), .B(n32066), .Z(n32061) );
  AND U40935 ( .A(n32067), .B(n32068), .Z(n31955) );
  XOR U40936 ( .A(n32035), .B(n32034), .Z(N62542) );
  XNOR U40937 ( .A(n32052), .B(n32053), .Z(n32034) );
  XNOR U40938 ( .A(n32067), .B(n32068), .Z(n32053) );
  XOR U40939 ( .A(n32064), .B(n32063), .Z(n32068) );
  XOR U40940 ( .A(y[3612]), .B(x[3612]), .Z(n32063) );
  XOR U40941 ( .A(n32066), .B(n32065), .Z(n32064) );
  XOR U40942 ( .A(y[3614]), .B(x[3614]), .Z(n32065) );
  XOR U40943 ( .A(y[3613]), .B(x[3613]), .Z(n32066) );
  XOR U40944 ( .A(n32058), .B(n32057), .Z(n32067) );
  XOR U40945 ( .A(n32060), .B(n32059), .Z(n32057) );
  XOR U40946 ( .A(y[3611]), .B(x[3611]), .Z(n32059) );
  XOR U40947 ( .A(y[3610]), .B(x[3610]), .Z(n32060) );
  XOR U40948 ( .A(y[3609]), .B(x[3609]), .Z(n32058) );
  XNOR U40949 ( .A(n32051), .B(n32050), .Z(n32052) );
  XNOR U40950 ( .A(n32047), .B(n32046), .Z(n32050) );
  XOR U40951 ( .A(n32049), .B(n32048), .Z(n32046) );
  XOR U40952 ( .A(y[3608]), .B(x[3608]), .Z(n32048) );
  XOR U40953 ( .A(y[3607]), .B(x[3607]), .Z(n32049) );
  XOR U40954 ( .A(y[3606]), .B(x[3606]), .Z(n32047) );
  XOR U40955 ( .A(n32041), .B(n32040), .Z(n32051) );
  XOR U40956 ( .A(n32043), .B(n32042), .Z(n32040) );
  XOR U40957 ( .A(y[3605]), .B(x[3605]), .Z(n32042) );
  XOR U40958 ( .A(y[3604]), .B(x[3604]), .Z(n32043) );
  XOR U40959 ( .A(y[3603]), .B(x[3603]), .Z(n32041) );
  XNOR U40960 ( .A(n32017), .B(n32018), .Z(n32035) );
  XNOR U40961 ( .A(n32032), .B(n32033), .Z(n32018) );
  XOR U40962 ( .A(n32029), .B(n32028), .Z(n32033) );
  XOR U40963 ( .A(y[3600]), .B(x[3600]), .Z(n32028) );
  XOR U40964 ( .A(n32031), .B(n32030), .Z(n32029) );
  XOR U40965 ( .A(y[3602]), .B(x[3602]), .Z(n32030) );
  XOR U40966 ( .A(y[3601]), .B(x[3601]), .Z(n32031) );
  XOR U40967 ( .A(n32023), .B(n32022), .Z(n32032) );
  XOR U40968 ( .A(n32025), .B(n32024), .Z(n32022) );
  XOR U40969 ( .A(y[3599]), .B(x[3599]), .Z(n32024) );
  XOR U40970 ( .A(y[3598]), .B(x[3598]), .Z(n32025) );
  XOR U40971 ( .A(y[3597]), .B(x[3597]), .Z(n32023) );
  XNOR U40972 ( .A(n32016), .B(n32015), .Z(n32017) );
  XNOR U40973 ( .A(n32012), .B(n32011), .Z(n32015) );
  XOR U40974 ( .A(n32014), .B(n32013), .Z(n32011) );
  XOR U40975 ( .A(y[3596]), .B(x[3596]), .Z(n32013) );
  XOR U40976 ( .A(y[3595]), .B(x[3595]), .Z(n32014) );
  XOR U40977 ( .A(y[3594]), .B(x[3594]), .Z(n32012) );
  XOR U40978 ( .A(n32006), .B(n32005), .Z(n32016) );
  XOR U40979 ( .A(n32008), .B(n32007), .Z(n32005) );
  XOR U40980 ( .A(y[3593]), .B(x[3593]), .Z(n32007) );
  XOR U40981 ( .A(y[3592]), .B(x[3592]), .Z(n32008) );
  XOR U40982 ( .A(y[3591]), .B(x[3591]), .Z(n32006) );
  NAND U40983 ( .A(n32069), .B(n32070), .Z(N62533) );
  NAND U40984 ( .A(n32071), .B(n32072), .Z(n32070) );
  NANDN U40985 ( .A(n32073), .B(n32074), .Z(n32072) );
  NANDN U40986 ( .A(n32074), .B(n32073), .Z(n32069) );
  XOR U40987 ( .A(n32073), .B(n32075), .Z(N62532) );
  XNOR U40988 ( .A(n32071), .B(n32074), .Z(n32075) );
  NAND U40989 ( .A(n32076), .B(n32077), .Z(n32074) );
  NAND U40990 ( .A(n32078), .B(n32079), .Z(n32077) );
  NANDN U40991 ( .A(n32080), .B(n32081), .Z(n32079) );
  NANDN U40992 ( .A(n32081), .B(n32080), .Z(n32076) );
  AND U40993 ( .A(n32082), .B(n32083), .Z(n32071) );
  NAND U40994 ( .A(n32084), .B(n32085), .Z(n32083) );
  NANDN U40995 ( .A(n32086), .B(n32087), .Z(n32085) );
  NANDN U40996 ( .A(n32087), .B(n32086), .Z(n32082) );
  IV U40997 ( .A(n32088), .Z(n32087) );
  AND U40998 ( .A(n32089), .B(n32090), .Z(n32073) );
  NAND U40999 ( .A(n32091), .B(n32092), .Z(n32090) );
  NANDN U41000 ( .A(n32093), .B(n32094), .Z(n32092) );
  NANDN U41001 ( .A(n32094), .B(n32093), .Z(n32089) );
  XOR U41002 ( .A(n32086), .B(n32095), .Z(N62531) );
  XNOR U41003 ( .A(n32084), .B(n32088), .Z(n32095) );
  XOR U41004 ( .A(n32081), .B(n32096), .Z(n32088) );
  XNOR U41005 ( .A(n32078), .B(n32080), .Z(n32096) );
  AND U41006 ( .A(n32097), .B(n32098), .Z(n32080) );
  NANDN U41007 ( .A(n32099), .B(n32100), .Z(n32098) );
  OR U41008 ( .A(n32101), .B(n32102), .Z(n32100) );
  IV U41009 ( .A(n32103), .Z(n32102) );
  NANDN U41010 ( .A(n32103), .B(n32101), .Z(n32097) );
  AND U41011 ( .A(n32104), .B(n32105), .Z(n32078) );
  NAND U41012 ( .A(n32106), .B(n32107), .Z(n32105) );
  NANDN U41013 ( .A(n32108), .B(n32109), .Z(n32107) );
  NANDN U41014 ( .A(n32109), .B(n32108), .Z(n32104) );
  IV U41015 ( .A(n32110), .Z(n32109) );
  NAND U41016 ( .A(n32111), .B(n32112), .Z(n32081) );
  NANDN U41017 ( .A(n32113), .B(n32114), .Z(n32112) );
  NANDN U41018 ( .A(n32115), .B(n32116), .Z(n32114) );
  NANDN U41019 ( .A(n32116), .B(n32115), .Z(n32111) );
  IV U41020 ( .A(n32117), .Z(n32115) );
  AND U41021 ( .A(n32118), .B(n32119), .Z(n32084) );
  NAND U41022 ( .A(n32120), .B(n32121), .Z(n32119) );
  NANDN U41023 ( .A(n32122), .B(n32123), .Z(n32121) );
  NANDN U41024 ( .A(n32123), .B(n32122), .Z(n32118) );
  XOR U41025 ( .A(n32094), .B(n32124), .Z(n32086) );
  XNOR U41026 ( .A(n32091), .B(n32093), .Z(n32124) );
  AND U41027 ( .A(n32125), .B(n32126), .Z(n32093) );
  NANDN U41028 ( .A(n32127), .B(n32128), .Z(n32126) );
  OR U41029 ( .A(n32129), .B(n32130), .Z(n32128) );
  IV U41030 ( .A(n32131), .Z(n32130) );
  NANDN U41031 ( .A(n32131), .B(n32129), .Z(n32125) );
  AND U41032 ( .A(n32132), .B(n32133), .Z(n32091) );
  NAND U41033 ( .A(n32134), .B(n32135), .Z(n32133) );
  NANDN U41034 ( .A(n32136), .B(n32137), .Z(n32135) );
  NANDN U41035 ( .A(n32137), .B(n32136), .Z(n32132) );
  IV U41036 ( .A(n32138), .Z(n32137) );
  NAND U41037 ( .A(n32139), .B(n32140), .Z(n32094) );
  NANDN U41038 ( .A(n32141), .B(n32142), .Z(n32140) );
  NANDN U41039 ( .A(n32143), .B(n32144), .Z(n32142) );
  NANDN U41040 ( .A(n32144), .B(n32143), .Z(n32139) );
  IV U41041 ( .A(n32145), .Z(n32143) );
  XOR U41042 ( .A(n32120), .B(n32146), .Z(N62530) );
  XNOR U41043 ( .A(n32123), .B(n32122), .Z(n32146) );
  XNOR U41044 ( .A(n32134), .B(n32147), .Z(n32122) );
  XNOR U41045 ( .A(n32138), .B(n32136), .Z(n32147) );
  XOR U41046 ( .A(n32144), .B(n32148), .Z(n32136) );
  XNOR U41047 ( .A(n32141), .B(n32145), .Z(n32148) );
  AND U41048 ( .A(n32149), .B(n32150), .Z(n32145) );
  NAND U41049 ( .A(n32151), .B(n32152), .Z(n32150) );
  NAND U41050 ( .A(n32153), .B(n32154), .Z(n32149) );
  AND U41051 ( .A(n32155), .B(n32156), .Z(n32141) );
  NAND U41052 ( .A(n32157), .B(n32158), .Z(n32156) );
  NAND U41053 ( .A(n32159), .B(n32160), .Z(n32155) );
  NANDN U41054 ( .A(n32161), .B(n32162), .Z(n32144) );
  ANDN U41055 ( .B(n32163), .A(n32164), .Z(n32138) );
  XNOR U41056 ( .A(n32129), .B(n32165), .Z(n32134) );
  XNOR U41057 ( .A(n32127), .B(n32131), .Z(n32165) );
  AND U41058 ( .A(n32166), .B(n32167), .Z(n32131) );
  NAND U41059 ( .A(n32168), .B(n32169), .Z(n32167) );
  NAND U41060 ( .A(n32170), .B(n32171), .Z(n32166) );
  AND U41061 ( .A(n32172), .B(n32173), .Z(n32127) );
  NAND U41062 ( .A(n32174), .B(n32175), .Z(n32173) );
  NAND U41063 ( .A(n32176), .B(n32177), .Z(n32172) );
  AND U41064 ( .A(n32178), .B(n32179), .Z(n32129) );
  NAND U41065 ( .A(n32180), .B(n32181), .Z(n32123) );
  XNOR U41066 ( .A(n32106), .B(n32182), .Z(n32120) );
  XNOR U41067 ( .A(n32110), .B(n32108), .Z(n32182) );
  XOR U41068 ( .A(n32116), .B(n32183), .Z(n32108) );
  XNOR U41069 ( .A(n32113), .B(n32117), .Z(n32183) );
  AND U41070 ( .A(n32184), .B(n32185), .Z(n32117) );
  NAND U41071 ( .A(n32186), .B(n32187), .Z(n32185) );
  NAND U41072 ( .A(n32188), .B(n32189), .Z(n32184) );
  AND U41073 ( .A(n32190), .B(n32191), .Z(n32113) );
  NAND U41074 ( .A(n32192), .B(n32193), .Z(n32191) );
  NAND U41075 ( .A(n32194), .B(n32195), .Z(n32190) );
  NANDN U41076 ( .A(n32196), .B(n32197), .Z(n32116) );
  ANDN U41077 ( .B(n32198), .A(n32199), .Z(n32110) );
  XNOR U41078 ( .A(n32101), .B(n32200), .Z(n32106) );
  XNOR U41079 ( .A(n32099), .B(n32103), .Z(n32200) );
  AND U41080 ( .A(n32201), .B(n32202), .Z(n32103) );
  NAND U41081 ( .A(n32203), .B(n32204), .Z(n32202) );
  NAND U41082 ( .A(n32205), .B(n32206), .Z(n32201) );
  AND U41083 ( .A(n32207), .B(n32208), .Z(n32099) );
  NAND U41084 ( .A(n32209), .B(n32210), .Z(n32208) );
  NAND U41085 ( .A(n32211), .B(n32212), .Z(n32207) );
  AND U41086 ( .A(n32213), .B(n32214), .Z(n32101) );
  XOR U41087 ( .A(n32181), .B(n32180), .Z(N62529) );
  XNOR U41088 ( .A(n32198), .B(n32199), .Z(n32180) );
  XNOR U41089 ( .A(n32213), .B(n32214), .Z(n32199) );
  XOR U41090 ( .A(n32210), .B(n32209), .Z(n32214) );
  XOR U41091 ( .A(y[3588]), .B(x[3588]), .Z(n32209) );
  XOR U41092 ( .A(n32212), .B(n32211), .Z(n32210) );
  XOR U41093 ( .A(y[3590]), .B(x[3590]), .Z(n32211) );
  XOR U41094 ( .A(y[3589]), .B(x[3589]), .Z(n32212) );
  XOR U41095 ( .A(n32204), .B(n32203), .Z(n32213) );
  XOR U41096 ( .A(n32206), .B(n32205), .Z(n32203) );
  XOR U41097 ( .A(y[3587]), .B(x[3587]), .Z(n32205) );
  XOR U41098 ( .A(y[3586]), .B(x[3586]), .Z(n32206) );
  XOR U41099 ( .A(y[3585]), .B(x[3585]), .Z(n32204) );
  XNOR U41100 ( .A(n32197), .B(n32196), .Z(n32198) );
  XNOR U41101 ( .A(n32193), .B(n32192), .Z(n32196) );
  XOR U41102 ( .A(n32195), .B(n32194), .Z(n32192) );
  XOR U41103 ( .A(y[3584]), .B(x[3584]), .Z(n32194) );
  XOR U41104 ( .A(y[3583]), .B(x[3583]), .Z(n32195) );
  XOR U41105 ( .A(y[3582]), .B(x[3582]), .Z(n32193) );
  XOR U41106 ( .A(n32187), .B(n32186), .Z(n32197) );
  XOR U41107 ( .A(n32189), .B(n32188), .Z(n32186) );
  XOR U41108 ( .A(y[3581]), .B(x[3581]), .Z(n32188) );
  XOR U41109 ( .A(y[3580]), .B(x[3580]), .Z(n32189) );
  XOR U41110 ( .A(y[3579]), .B(x[3579]), .Z(n32187) );
  XNOR U41111 ( .A(n32163), .B(n32164), .Z(n32181) );
  XNOR U41112 ( .A(n32178), .B(n32179), .Z(n32164) );
  XOR U41113 ( .A(n32175), .B(n32174), .Z(n32179) );
  XOR U41114 ( .A(y[3576]), .B(x[3576]), .Z(n32174) );
  XOR U41115 ( .A(n32177), .B(n32176), .Z(n32175) );
  XOR U41116 ( .A(y[3578]), .B(x[3578]), .Z(n32176) );
  XOR U41117 ( .A(y[3577]), .B(x[3577]), .Z(n32177) );
  XOR U41118 ( .A(n32169), .B(n32168), .Z(n32178) );
  XOR U41119 ( .A(n32171), .B(n32170), .Z(n32168) );
  XOR U41120 ( .A(y[3575]), .B(x[3575]), .Z(n32170) );
  XOR U41121 ( .A(y[3574]), .B(x[3574]), .Z(n32171) );
  XOR U41122 ( .A(y[3573]), .B(x[3573]), .Z(n32169) );
  XNOR U41123 ( .A(n32162), .B(n32161), .Z(n32163) );
  XNOR U41124 ( .A(n32158), .B(n32157), .Z(n32161) );
  XOR U41125 ( .A(n32160), .B(n32159), .Z(n32157) );
  XOR U41126 ( .A(y[3572]), .B(x[3572]), .Z(n32159) );
  XOR U41127 ( .A(y[3571]), .B(x[3571]), .Z(n32160) );
  XOR U41128 ( .A(y[3570]), .B(x[3570]), .Z(n32158) );
  XOR U41129 ( .A(n32152), .B(n32151), .Z(n32162) );
  XOR U41130 ( .A(n32154), .B(n32153), .Z(n32151) );
  XOR U41131 ( .A(y[3569]), .B(x[3569]), .Z(n32153) );
  XOR U41132 ( .A(y[3568]), .B(x[3568]), .Z(n32154) );
  XOR U41133 ( .A(y[3567]), .B(x[3567]), .Z(n32152) );
  NAND U41134 ( .A(n32215), .B(n32216), .Z(N62520) );
  NAND U41135 ( .A(n32217), .B(n32218), .Z(n32216) );
  NANDN U41136 ( .A(n32219), .B(n32220), .Z(n32218) );
  NANDN U41137 ( .A(n32220), .B(n32219), .Z(n32215) );
  XOR U41138 ( .A(n32219), .B(n32221), .Z(N62519) );
  XNOR U41139 ( .A(n32217), .B(n32220), .Z(n32221) );
  NAND U41140 ( .A(n32222), .B(n32223), .Z(n32220) );
  NAND U41141 ( .A(n32224), .B(n32225), .Z(n32223) );
  NANDN U41142 ( .A(n32226), .B(n32227), .Z(n32225) );
  NANDN U41143 ( .A(n32227), .B(n32226), .Z(n32222) );
  AND U41144 ( .A(n32228), .B(n32229), .Z(n32217) );
  NAND U41145 ( .A(n32230), .B(n32231), .Z(n32229) );
  NANDN U41146 ( .A(n32232), .B(n32233), .Z(n32231) );
  NANDN U41147 ( .A(n32233), .B(n32232), .Z(n32228) );
  IV U41148 ( .A(n32234), .Z(n32233) );
  AND U41149 ( .A(n32235), .B(n32236), .Z(n32219) );
  NAND U41150 ( .A(n32237), .B(n32238), .Z(n32236) );
  NANDN U41151 ( .A(n32239), .B(n32240), .Z(n32238) );
  NANDN U41152 ( .A(n32240), .B(n32239), .Z(n32235) );
  XOR U41153 ( .A(n32232), .B(n32241), .Z(N62518) );
  XNOR U41154 ( .A(n32230), .B(n32234), .Z(n32241) );
  XOR U41155 ( .A(n32227), .B(n32242), .Z(n32234) );
  XNOR U41156 ( .A(n32224), .B(n32226), .Z(n32242) );
  AND U41157 ( .A(n32243), .B(n32244), .Z(n32226) );
  NANDN U41158 ( .A(n32245), .B(n32246), .Z(n32244) );
  OR U41159 ( .A(n32247), .B(n32248), .Z(n32246) );
  IV U41160 ( .A(n32249), .Z(n32248) );
  NANDN U41161 ( .A(n32249), .B(n32247), .Z(n32243) );
  AND U41162 ( .A(n32250), .B(n32251), .Z(n32224) );
  NAND U41163 ( .A(n32252), .B(n32253), .Z(n32251) );
  NANDN U41164 ( .A(n32254), .B(n32255), .Z(n32253) );
  NANDN U41165 ( .A(n32255), .B(n32254), .Z(n32250) );
  IV U41166 ( .A(n32256), .Z(n32255) );
  NAND U41167 ( .A(n32257), .B(n32258), .Z(n32227) );
  NANDN U41168 ( .A(n32259), .B(n32260), .Z(n32258) );
  NANDN U41169 ( .A(n32261), .B(n32262), .Z(n32260) );
  NANDN U41170 ( .A(n32262), .B(n32261), .Z(n32257) );
  IV U41171 ( .A(n32263), .Z(n32261) );
  AND U41172 ( .A(n32264), .B(n32265), .Z(n32230) );
  NAND U41173 ( .A(n32266), .B(n32267), .Z(n32265) );
  NANDN U41174 ( .A(n32268), .B(n32269), .Z(n32267) );
  NANDN U41175 ( .A(n32269), .B(n32268), .Z(n32264) );
  XOR U41176 ( .A(n32240), .B(n32270), .Z(n32232) );
  XNOR U41177 ( .A(n32237), .B(n32239), .Z(n32270) );
  AND U41178 ( .A(n32271), .B(n32272), .Z(n32239) );
  NANDN U41179 ( .A(n32273), .B(n32274), .Z(n32272) );
  OR U41180 ( .A(n32275), .B(n32276), .Z(n32274) );
  IV U41181 ( .A(n32277), .Z(n32276) );
  NANDN U41182 ( .A(n32277), .B(n32275), .Z(n32271) );
  AND U41183 ( .A(n32278), .B(n32279), .Z(n32237) );
  NAND U41184 ( .A(n32280), .B(n32281), .Z(n32279) );
  NANDN U41185 ( .A(n32282), .B(n32283), .Z(n32281) );
  NANDN U41186 ( .A(n32283), .B(n32282), .Z(n32278) );
  IV U41187 ( .A(n32284), .Z(n32283) );
  NAND U41188 ( .A(n32285), .B(n32286), .Z(n32240) );
  NANDN U41189 ( .A(n32287), .B(n32288), .Z(n32286) );
  NANDN U41190 ( .A(n32289), .B(n32290), .Z(n32288) );
  NANDN U41191 ( .A(n32290), .B(n32289), .Z(n32285) );
  IV U41192 ( .A(n32291), .Z(n32289) );
  XOR U41193 ( .A(n32266), .B(n32292), .Z(N62517) );
  XNOR U41194 ( .A(n32269), .B(n32268), .Z(n32292) );
  XNOR U41195 ( .A(n32280), .B(n32293), .Z(n32268) );
  XNOR U41196 ( .A(n32284), .B(n32282), .Z(n32293) );
  XOR U41197 ( .A(n32290), .B(n32294), .Z(n32282) );
  XNOR U41198 ( .A(n32287), .B(n32291), .Z(n32294) );
  AND U41199 ( .A(n32295), .B(n32296), .Z(n32291) );
  NAND U41200 ( .A(n32297), .B(n32298), .Z(n32296) );
  NAND U41201 ( .A(n32299), .B(n32300), .Z(n32295) );
  AND U41202 ( .A(n32301), .B(n32302), .Z(n32287) );
  NAND U41203 ( .A(n32303), .B(n32304), .Z(n32302) );
  NAND U41204 ( .A(n32305), .B(n32306), .Z(n32301) );
  NANDN U41205 ( .A(n32307), .B(n32308), .Z(n32290) );
  ANDN U41206 ( .B(n32309), .A(n32310), .Z(n32284) );
  XNOR U41207 ( .A(n32275), .B(n32311), .Z(n32280) );
  XNOR U41208 ( .A(n32273), .B(n32277), .Z(n32311) );
  AND U41209 ( .A(n32312), .B(n32313), .Z(n32277) );
  NAND U41210 ( .A(n32314), .B(n32315), .Z(n32313) );
  NAND U41211 ( .A(n32316), .B(n32317), .Z(n32312) );
  AND U41212 ( .A(n32318), .B(n32319), .Z(n32273) );
  NAND U41213 ( .A(n32320), .B(n32321), .Z(n32319) );
  NAND U41214 ( .A(n32322), .B(n32323), .Z(n32318) );
  AND U41215 ( .A(n32324), .B(n32325), .Z(n32275) );
  NAND U41216 ( .A(n32326), .B(n32327), .Z(n32269) );
  XNOR U41217 ( .A(n32252), .B(n32328), .Z(n32266) );
  XNOR U41218 ( .A(n32256), .B(n32254), .Z(n32328) );
  XOR U41219 ( .A(n32262), .B(n32329), .Z(n32254) );
  XNOR U41220 ( .A(n32259), .B(n32263), .Z(n32329) );
  AND U41221 ( .A(n32330), .B(n32331), .Z(n32263) );
  NAND U41222 ( .A(n32332), .B(n32333), .Z(n32331) );
  NAND U41223 ( .A(n32334), .B(n32335), .Z(n32330) );
  AND U41224 ( .A(n32336), .B(n32337), .Z(n32259) );
  NAND U41225 ( .A(n32338), .B(n32339), .Z(n32337) );
  NAND U41226 ( .A(n32340), .B(n32341), .Z(n32336) );
  NANDN U41227 ( .A(n32342), .B(n32343), .Z(n32262) );
  ANDN U41228 ( .B(n32344), .A(n32345), .Z(n32256) );
  XNOR U41229 ( .A(n32247), .B(n32346), .Z(n32252) );
  XNOR U41230 ( .A(n32245), .B(n32249), .Z(n32346) );
  AND U41231 ( .A(n32347), .B(n32348), .Z(n32249) );
  NAND U41232 ( .A(n32349), .B(n32350), .Z(n32348) );
  NAND U41233 ( .A(n32351), .B(n32352), .Z(n32347) );
  AND U41234 ( .A(n32353), .B(n32354), .Z(n32245) );
  NAND U41235 ( .A(n32355), .B(n32356), .Z(n32354) );
  NAND U41236 ( .A(n32357), .B(n32358), .Z(n32353) );
  AND U41237 ( .A(n32359), .B(n32360), .Z(n32247) );
  XOR U41238 ( .A(n32327), .B(n32326), .Z(N62516) );
  XNOR U41239 ( .A(n32344), .B(n32345), .Z(n32326) );
  XNOR U41240 ( .A(n32359), .B(n32360), .Z(n32345) );
  XOR U41241 ( .A(n32356), .B(n32355), .Z(n32360) );
  XOR U41242 ( .A(y[3564]), .B(x[3564]), .Z(n32355) );
  XOR U41243 ( .A(n32358), .B(n32357), .Z(n32356) );
  XOR U41244 ( .A(y[3566]), .B(x[3566]), .Z(n32357) );
  XOR U41245 ( .A(y[3565]), .B(x[3565]), .Z(n32358) );
  XOR U41246 ( .A(n32350), .B(n32349), .Z(n32359) );
  XOR U41247 ( .A(n32352), .B(n32351), .Z(n32349) );
  XOR U41248 ( .A(y[3563]), .B(x[3563]), .Z(n32351) );
  XOR U41249 ( .A(y[3562]), .B(x[3562]), .Z(n32352) );
  XOR U41250 ( .A(y[3561]), .B(x[3561]), .Z(n32350) );
  XNOR U41251 ( .A(n32343), .B(n32342), .Z(n32344) );
  XNOR U41252 ( .A(n32339), .B(n32338), .Z(n32342) );
  XOR U41253 ( .A(n32341), .B(n32340), .Z(n32338) );
  XOR U41254 ( .A(y[3560]), .B(x[3560]), .Z(n32340) );
  XOR U41255 ( .A(y[3559]), .B(x[3559]), .Z(n32341) );
  XOR U41256 ( .A(y[3558]), .B(x[3558]), .Z(n32339) );
  XOR U41257 ( .A(n32333), .B(n32332), .Z(n32343) );
  XOR U41258 ( .A(n32335), .B(n32334), .Z(n32332) );
  XOR U41259 ( .A(y[3557]), .B(x[3557]), .Z(n32334) );
  XOR U41260 ( .A(y[3556]), .B(x[3556]), .Z(n32335) );
  XOR U41261 ( .A(y[3555]), .B(x[3555]), .Z(n32333) );
  XNOR U41262 ( .A(n32309), .B(n32310), .Z(n32327) );
  XNOR U41263 ( .A(n32324), .B(n32325), .Z(n32310) );
  XOR U41264 ( .A(n32321), .B(n32320), .Z(n32325) );
  XOR U41265 ( .A(y[3552]), .B(x[3552]), .Z(n32320) );
  XOR U41266 ( .A(n32323), .B(n32322), .Z(n32321) );
  XOR U41267 ( .A(y[3554]), .B(x[3554]), .Z(n32322) );
  XOR U41268 ( .A(y[3553]), .B(x[3553]), .Z(n32323) );
  XOR U41269 ( .A(n32315), .B(n32314), .Z(n32324) );
  XOR U41270 ( .A(n32317), .B(n32316), .Z(n32314) );
  XOR U41271 ( .A(y[3551]), .B(x[3551]), .Z(n32316) );
  XOR U41272 ( .A(y[3550]), .B(x[3550]), .Z(n32317) );
  XOR U41273 ( .A(y[3549]), .B(x[3549]), .Z(n32315) );
  XNOR U41274 ( .A(n32308), .B(n32307), .Z(n32309) );
  XNOR U41275 ( .A(n32304), .B(n32303), .Z(n32307) );
  XOR U41276 ( .A(n32306), .B(n32305), .Z(n32303) );
  XOR U41277 ( .A(y[3548]), .B(x[3548]), .Z(n32305) );
  XOR U41278 ( .A(y[3547]), .B(x[3547]), .Z(n32306) );
  XOR U41279 ( .A(y[3546]), .B(x[3546]), .Z(n32304) );
  XOR U41280 ( .A(n32298), .B(n32297), .Z(n32308) );
  XOR U41281 ( .A(n32300), .B(n32299), .Z(n32297) );
  XOR U41282 ( .A(y[3545]), .B(x[3545]), .Z(n32299) );
  XOR U41283 ( .A(y[3544]), .B(x[3544]), .Z(n32300) );
  XOR U41284 ( .A(y[3543]), .B(x[3543]), .Z(n32298) );
  NAND U41285 ( .A(n32361), .B(n32362), .Z(N62507) );
  NAND U41286 ( .A(n32363), .B(n32364), .Z(n32362) );
  NANDN U41287 ( .A(n32365), .B(n32366), .Z(n32364) );
  NANDN U41288 ( .A(n32366), .B(n32365), .Z(n32361) );
  XOR U41289 ( .A(n32365), .B(n32367), .Z(N62506) );
  XNOR U41290 ( .A(n32363), .B(n32366), .Z(n32367) );
  NAND U41291 ( .A(n32368), .B(n32369), .Z(n32366) );
  NAND U41292 ( .A(n32370), .B(n32371), .Z(n32369) );
  NANDN U41293 ( .A(n32372), .B(n32373), .Z(n32371) );
  NANDN U41294 ( .A(n32373), .B(n32372), .Z(n32368) );
  AND U41295 ( .A(n32374), .B(n32375), .Z(n32363) );
  NAND U41296 ( .A(n32376), .B(n32377), .Z(n32375) );
  NANDN U41297 ( .A(n32378), .B(n32379), .Z(n32377) );
  NANDN U41298 ( .A(n32379), .B(n32378), .Z(n32374) );
  IV U41299 ( .A(n32380), .Z(n32379) );
  AND U41300 ( .A(n32381), .B(n32382), .Z(n32365) );
  NAND U41301 ( .A(n32383), .B(n32384), .Z(n32382) );
  NANDN U41302 ( .A(n32385), .B(n32386), .Z(n32384) );
  NANDN U41303 ( .A(n32386), .B(n32385), .Z(n32381) );
  XOR U41304 ( .A(n32378), .B(n32387), .Z(N62505) );
  XNOR U41305 ( .A(n32376), .B(n32380), .Z(n32387) );
  XOR U41306 ( .A(n32373), .B(n32388), .Z(n32380) );
  XNOR U41307 ( .A(n32370), .B(n32372), .Z(n32388) );
  AND U41308 ( .A(n32389), .B(n32390), .Z(n32372) );
  NANDN U41309 ( .A(n32391), .B(n32392), .Z(n32390) );
  OR U41310 ( .A(n32393), .B(n32394), .Z(n32392) );
  IV U41311 ( .A(n32395), .Z(n32394) );
  NANDN U41312 ( .A(n32395), .B(n32393), .Z(n32389) );
  AND U41313 ( .A(n32396), .B(n32397), .Z(n32370) );
  NAND U41314 ( .A(n32398), .B(n32399), .Z(n32397) );
  NANDN U41315 ( .A(n32400), .B(n32401), .Z(n32399) );
  NANDN U41316 ( .A(n32401), .B(n32400), .Z(n32396) );
  IV U41317 ( .A(n32402), .Z(n32401) );
  NAND U41318 ( .A(n32403), .B(n32404), .Z(n32373) );
  NANDN U41319 ( .A(n32405), .B(n32406), .Z(n32404) );
  NANDN U41320 ( .A(n32407), .B(n32408), .Z(n32406) );
  NANDN U41321 ( .A(n32408), .B(n32407), .Z(n32403) );
  IV U41322 ( .A(n32409), .Z(n32407) );
  AND U41323 ( .A(n32410), .B(n32411), .Z(n32376) );
  NAND U41324 ( .A(n32412), .B(n32413), .Z(n32411) );
  NANDN U41325 ( .A(n32414), .B(n32415), .Z(n32413) );
  NANDN U41326 ( .A(n32415), .B(n32414), .Z(n32410) );
  XOR U41327 ( .A(n32386), .B(n32416), .Z(n32378) );
  XNOR U41328 ( .A(n32383), .B(n32385), .Z(n32416) );
  AND U41329 ( .A(n32417), .B(n32418), .Z(n32385) );
  NANDN U41330 ( .A(n32419), .B(n32420), .Z(n32418) );
  OR U41331 ( .A(n32421), .B(n32422), .Z(n32420) );
  IV U41332 ( .A(n32423), .Z(n32422) );
  NANDN U41333 ( .A(n32423), .B(n32421), .Z(n32417) );
  AND U41334 ( .A(n32424), .B(n32425), .Z(n32383) );
  NAND U41335 ( .A(n32426), .B(n32427), .Z(n32425) );
  NANDN U41336 ( .A(n32428), .B(n32429), .Z(n32427) );
  NANDN U41337 ( .A(n32429), .B(n32428), .Z(n32424) );
  IV U41338 ( .A(n32430), .Z(n32429) );
  NAND U41339 ( .A(n32431), .B(n32432), .Z(n32386) );
  NANDN U41340 ( .A(n32433), .B(n32434), .Z(n32432) );
  NANDN U41341 ( .A(n32435), .B(n32436), .Z(n32434) );
  NANDN U41342 ( .A(n32436), .B(n32435), .Z(n32431) );
  IV U41343 ( .A(n32437), .Z(n32435) );
  XOR U41344 ( .A(n32412), .B(n32438), .Z(N62504) );
  XNOR U41345 ( .A(n32415), .B(n32414), .Z(n32438) );
  XNOR U41346 ( .A(n32426), .B(n32439), .Z(n32414) );
  XNOR U41347 ( .A(n32430), .B(n32428), .Z(n32439) );
  XOR U41348 ( .A(n32436), .B(n32440), .Z(n32428) );
  XNOR U41349 ( .A(n32433), .B(n32437), .Z(n32440) );
  AND U41350 ( .A(n32441), .B(n32442), .Z(n32437) );
  NAND U41351 ( .A(n32443), .B(n32444), .Z(n32442) );
  NAND U41352 ( .A(n32445), .B(n32446), .Z(n32441) );
  AND U41353 ( .A(n32447), .B(n32448), .Z(n32433) );
  NAND U41354 ( .A(n32449), .B(n32450), .Z(n32448) );
  NAND U41355 ( .A(n32451), .B(n32452), .Z(n32447) );
  NANDN U41356 ( .A(n32453), .B(n32454), .Z(n32436) );
  ANDN U41357 ( .B(n32455), .A(n32456), .Z(n32430) );
  XNOR U41358 ( .A(n32421), .B(n32457), .Z(n32426) );
  XNOR U41359 ( .A(n32419), .B(n32423), .Z(n32457) );
  AND U41360 ( .A(n32458), .B(n32459), .Z(n32423) );
  NAND U41361 ( .A(n32460), .B(n32461), .Z(n32459) );
  NAND U41362 ( .A(n32462), .B(n32463), .Z(n32458) );
  AND U41363 ( .A(n32464), .B(n32465), .Z(n32419) );
  NAND U41364 ( .A(n32466), .B(n32467), .Z(n32465) );
  NAND U41365 ( .A(n32468), .B(n32469), .Z(n32464) );
  AND U41366 ( .A(n32470), .B(n32471), .Z(n32421) );
  NAND U41367 ( .A(n32472), .B(n32473), .Z(n32415) );
  XNOR U41368 ( .A(n32398), .B(n32474), .Z(n32412) );
  XNOR U41369 ( .A(n32402), .B(n32400), .Z(n32474) );
  XOR U41370 ( .A(n32408), .B(n32475), .Z(n32400) );
  XNOR U41371 ( .A(n32405), .B(n32409), .Z(n32475) );
  AND U41372 ( .A(n32476), .B(n32477), .Z(n32409) );
  NAND U41373 ( .A(n32478), .B(n32479), .Z(n32477) );
  NAND U41374 ( .A(n32480), .B(n32481), .Z(n32476) );
  AND U41375 ( .A(n32482), .B(n32483), .Z(n32405) );
  NAND U41376 ( .A(n32484), .B(n32485), .Z(n32483) );
  NAND U41377 ( .A(n32486), .B(n32487), .Z(n32482) );
  NANDN U41378 ( .A(n32488), .B(n32489), .Z(n32408) );
  ANDN U41379 ( .B(n32490), .A(n32491), .Z(n32402) );
  XNOR U41380 ( .A(n32393), .B(n32492), .Z(n32398) );
  XNOR U41381 ( .A(n32391), .B(n32395), .Z(n32492) );
  AND U41382 ( .A(n32493), .B(n32494), .Z(n32395) );
  NAND U41383 ( .A(n32495), .B(n32496), .Z(n32494) );
  NAND U41384 ( .A(n32497), .B(n32498), .Z(n32493) );
  AND U41385 ( .A(n32499), .B(n32500), .Z(n32391) );
  NAND U41386 ( .A(n32501), .B(n32502), .Z(n32500) );
  NAND U41387 ( .A(n32503), .B(n32504), .Z(n32499) );
  AND U41388 ( .A(n32505), .B(n32506), .Z(n32393) );
  XOR U41389 ( .A(n32473), .B(n32472), .Z(N62503) );
  XNOR U41390 ( .A(n32490), .B(n32491), .Z(n32472) );
  XNOR U41391 ( .A(n32505), .B(n32506), .Z(n32491) );
  XOR U41392 ( .A(n32502), .B(n32501), .Z(n32506) );
  XOR U41393 ( .A(y[3540]), .B(x[3540]), .Z(n32501) );
  XOR U41394 ( .A(n32504), .B(n32503), .Z(n32502) );
  XOR U41395 ( .A(y[3542]), .B(x[3542]), .Z(n32503) );
  XOR U41396 ( .A(y[3541]), .B(x[3541]), .Z(n32504) );
  XOR U41397 ( .A(n32496), .B(n32495), .Z(n32505) );
  XOR U41398 ( .A(n32498), .B(n32497), .Z(n32495) );
  XOR U41399 ( .A(y[3539]), .B(x[3539]), .Z(n32497) );
  XOR U41400 ( .A(y[3538]), .B(x[3538]), .Z(n32498) );
  XOR U41401 ( .A(y[3537]), .B(x[3537]), .Z(n32496) );
  XNOR U41402 ( .A(n32489), .B(n32488), .Z(n32490) );
  XNOR U41403 ( .A(n32485), .B(n32484), .Z(n32488) );
  XOR U41404 ( .A(n32487), .B(n32486), .Z(n32484) );
  XOR U41405 ( .A(y[3536]), .B(x[3536]), .Z(n32486) );
  XOR U41406 ( .A(y[3535]), .B(x[3535]), .Z(n32487) );
  XOR U41407 ( .A(y[3534]), .B(x[3534]), .Z(n32485) );
  XOR U41408 ( .A(n32479), .B(n32478), .Z(n32489) );
  XOR U41409 ( .A(n32481), .B(n32480), .Z(n32478) );
  XOR U41410 ( .A(y[3533]), .B(x[3533]), .Z(n32480) );
  XOR U41411 ( .A(y[3532]), .B(x[3532]), .Z(n32481) );
  XOR U41412 ( .A(y[3531]), .B(x[3531]), .Z(n32479) );
  XNOR U41413 ( .A(n32455), .B(n32456), .Z(n32473) );
  XNOR U41414 ( .A(n32470), .B(n32471), .Z(n32456) );
  XOR U41415 ( .A(n32467), .B(n32466), .Z(n32471) );
  XOR U41416 ( .A(y[3528]), .B(x[3528]), .Z(n32466) );
  XOR U41417 ( .A(n32469), .B(n32468), .Z(n32467) );
  XOR U41418 ( .A(y[3530]), .B(x[3530]), .Z(n32468) );
  XOR U41419 ( .A(y[3529]), .B(x[3529]), .Z(n32469) );
  XOR U41420 ( .A(n32461), .B(n32460), .Z(n32470) );
  XOR U41421 ( .A(n32463), .B(n32462), .Z(n32460) );
  XOR U41422 ( .A(y[3527]), .B(x[3527]), .Z(n32462) );
  XOR U41423 ( .A(y[3526]), .B(x[3526]), .Z(n32463) );
  XOR U41424 ( .A(y[3525]), .B(x[3525]), .Z(n32461) );
  XNOR U41425 ( .A(n32454), .B(n32453), .Z(n32455) );
  XNOR U41426 ( .A(n32450), .B(n32449), .Z(n32453) );
  XOR U41427 ( .A(n32452), .B(n32451), .Z(n32449) );
  XOR U41428 ( .A(y[3524]), .B(x[3524]), .Z(n32451) );
  XOR U41429 ( .A(y[3523]), .B(x[3523]), .Z(n32452) );
  XOR U41430 ( .A(y[3522]), .B(x[3522]), .Z(n32450) );
  XOR U41431 ( .A(n32444), .B(n32443), .Z(n32454) );
  XOR U41432 ( .A(n32446), .B(n32445), .Z(n32443) );
  XOR U41433 ( .A(y[3521]), .B(x[3521]), .Z(n32445) );
  XOR U41434 ( .A(y[3520]), .B(x[3520]), .Z(n32446) );
  XOR U41435 ( .A(y[3519]), .B(x[3519]), .Z(n32444) );
  NAND U41436 ( .A(n32507), .B(n32508), .Z(N62494) );
  NAND U41437 ( .A(n32509), .B(n32510), .Z(n32508) );
  NANDN U41438 ( .A(n32511), .B(n32512), .Z(n32510) );
  NANDN U41439 ( .A(n32512), .B(n32511), .Z(n32507) );
  XOR U41440 ( .A(n32511), .B(n32513), .Z(N62493) );
  XNOR U41441 ( .A(n32509), .B(n32512), .Z(n32513) );
  NAND U41442 ( .A(n32514), .B(n32515), .Z(n32512) );
  NAND U41443 ( .A(n32516), .B(n32517), .Z(n32515) );
  NANDN U41444 ( .A(n32518), .B(n32519), .Z(n32517) );
  NANDN U41445 ( .A(n32519), .B(n32518), .Z(n32514) );
  AND U41446 ( .A(n32520), .B(n32521), .Z(n32509) );
  NAND U41447 ( .A(n32522), .B(n32523), .Z(n32521) );
  NANDN U41448 ( .A(n32524), .B(n32525), .Z(n32523) );
  NANDN U41449 ( .A(n32525), .B(n32524), .Z(n32520) );
  IV U41450 ( .A(n32526), .Z(n32525) );
  AND U41451 ( .A(n32527), .B(n32528), .Z(n32511) );
  NAND U41452 ( .A(n32529), .B(n32530), .Z(n32528) );
  NANDN U41453 ( .A(n32531), .B(n32532), .Z(n32530) );
  NANDN U41454 ( .A(n32532), .B(n32531), .Z(n32527) );
  XOR U41455 ( .A(n32524), .B(n32533), .Z(N62492) );
  XNOR U41456 ( .A(n32522), .B(n32526), .Z(n32533) );
  XOR U41457 ( .A(n32519), .B(n32534), .Z(n32526) );
  XNOR U41458 ( .A(n32516), .B(n32518), .Z(n32534) );
  AND U41459 ( .A(n32535), .B(n32536), .Z(n32518) );
  NANDN U41460 ( .A(n32537), .B(n32538), .Z(n32536) );
  OR U41461 ( .A(n32539), .B(n32540), .Z(n32538) );
  IV U41462 ( .A(n32541), .Z(n32540) );
  NANDN U41463 ( .A(n32541), .B(n32539), .Z(n32535) );
  AND U41464 ( .A(n32542), .B(n32543), .Z(n32516) );
  NAND U41465 ( .A(n32544), .B(n32545), .Z(n32543) );
  NANDN U41466 ( .A(n32546), .B(n32547), .Z(n32545) );
  NANDN U41467 ( .A(n32547), .B(n32546), .Z(n32542) );
  IV U41468 ( .A(n32548), .Z(n32547) );
  NAND U41469 ( .A(n32549), .B(n32550), .Z(n32519) );
  NANDN U41470 ( .A(n32551), .B(n32552), .Z(n32550) );
  NANDN U41471 ( .A(n32553), .B(n32554), .Z(n32552) );
  NANDN U41472 ( .A(n32554), .B(n32553), .Z(n32549) );
  IV U41473 ( .A(n32555), .Z(n32553) );
  AND U41474 ( .A(n32556), .B(n32557), .Z(n32522) );
  NAND U41475 ( .A(n32558), .B(n32559), .Z(n32557) );
  NANDN U41476 ( .A(n32560), .B(n32561), .Z(n32559) );
  NANDN U41477 ( .A(n32561), .B(n32560), .Z(n32556) );
  XOR U41478 ( .A(n32532), .B(n32562), .Z(n32524) );
  XNOR U41479 ( .A(n32529), .B(n32531), .Z(n32562) );
  AND U41480 ( .A(n32563), .B(n32564), .Z(n32531) );
  NANDN U41481 ( .A(n32565), .B(n32566), .Z(n32564) );
  OR U41482 ( .A(n32567), .B(n32568), .Z(n32566) );
  IV U41483 ( .A(n32569), .Z(n32568) );
  NANDN U41484 ( .A(n32569), .B(n32567), .Z(n32563) );
  AND U41485 ( .A(n32570), .B(n32571), .Z(n32529) );
  NAND U41486 ( .A(n32572), .B(n32573), .Z(n32571) );
  NANDN U41487 ( .A(n32574), .B(n32575), .Z(n32573) );
  NANDN U41488 ( .A(n32575), .B(n32574), .Z(n32570) );
  IV U41489 ( .A(n32576), .Z(n32575) );
  NAND U41490 ( .A(n32577), .B(n32578), .Z(n32532) );
  NANDN U41491 ( .A(n32579), .B(n32580), .Z(n32578) );
  NANDN U41492 ( .A(n32581), .B(n32582), .Z(n32580) );
  NANDN U41493 ( .A(n32582), .B(n32581), .Z(n32577) );
  IV U41494 ( .A(n32583), .Z(n32581) );
  XOR U41495 ( .A(n32558), .B(n32584), .Z(N62491) );
  XNOR U41496 ( .A(n32561), .B(n32560), .Z(n32584) );
  XNOR U41497 ( .A(n32572), .B(n32585), .Z(n32560) );
  XNOR U41498 ( .A(n32576), .B(n32574), .Z(n32585) );
  XOR U41499 ( .A(n32582), .B(n32586), .Z(n32574) );
  XNOR U41500 ( .A(n32579), .B(n32583), .Z(n32586) );
  AND U41501 ( .A(n32587), .B(n32588), .Z(n32583) );
  NAND U41502 ( .A(n32589), .B(n32590), .Z(n32588) );
  NAND U41503 ( .A(n32591), .B(n32592), .Z(n32587) );
  AND U41504 ( .A(n32593), .B(n32594), .Z(n32579) );
  NAND U41505 ( .A(n32595), .B(n32596), .Z(n32594) );
  NAND U41506 ( .A(n32597), .B(n32598), .Z(n32593) );
  NANDN U41507 ( .A(n32599), .B(n32600), .Z(n32582) );
  ANDN U41508 ( .B(n32601), .A(n32602), .Z(n32576) );
  XNOR U41509 ( .A(n32567), .B(n32603), .Z(n32572) );
  XNOR U41510 ( .A(n32565), .B(n32569), .Z(n32603) );
  AND U41511 ( .A(n32604), .B(n32605), .Z(n32569) );
  NAND U41512 ( .A(n32606), .B(n32607), .Z(n32605) );
  NAND U41513 ( .A(n32608), .B(n32609), .Z(n32604) );
  AND U41514 ( .A(n32610), .B(n32611), .Z(n32565) );
  NAND U41515 ( .A(n32612), .B(n32613), .Z(n32611) );
  NAND U41516 ( .A(n32614), .B(n32615), .Z(n32610) );
  AND U41517 ( .A(n32616), .B(n32617), .Z(n32567) );
  NAND U41518 ( .A(n32618), .B(n32619), .Z(n32561) );
  XNOR U41519 ( .A(n32544), .B(n32620), .Z(n32558) );
  XNOR U41520 ( .A(n32548), .B(n32546), .Z(n32620) );
  XOR U41521 ( .A(n32554), .B(n32621), .Z(n32546) );
  XNOR U41522 ( .A(n32551), .B(n32555), .Z(n32621) );
  AND U41523 ( .A(n32622), .B(n32623), .Z(n32555) );
  NAND U41524 ( .A(n32624), .B(n32625), .Z(n32623) );
  NAND U41525 ( .A(n32626), .B(n32627), .Z(n32622) );
  AND U41526 ( .A(n32628), .B(n32629), .Z(n32551) );
  NAND U41527 ( .A(n32630), .B(n32631), .Z(n32629) );
  NAND U41528 ( .A(n32632), .B(n32633), .Z(n32628) );
  NANDN U41529 ( .A(n32634), .B(n32635), .Z(n32554) );
  ANDN U41530 ( .B(n32636), .A(n32637), .Z(n32548) );
  XNOR U41531 ( .A(n32539), .B(n32638), .Z(n32544) );
  XNOR U41532 ( .A(n32537), .B(n32541), .Z(n32638) );
  AND U41533 ( .A(n32639), .B(n32640), .Z(n32541) );
  NAND U41534 ( .A(n32641), .B(n32642), .Z(n32640) );
  NAND U41535 ( .A(n32643), .B(n32644), .Z(n32639) );
  AND U41536 ( .A(n32645), .B(n32646), .Z(n32537) );
  NAND U41537 ( .A(n32647), .B(n32648), .Z(n32646) );
  NAND U41538 ( .A(n32649), .B(n32650), .Z(n32645) );
  AND U41539 ( .A(n32651), .B(n32652), .Z(n32539) );
  XOR U41540 ( .A(n32619), .B(n32618), .Z(N62490) );
  XNOR U41541 ( .A(n32636), .B(n32637), .Z(n32618) );
  XNOR U41542 ( .A(n32651), .B(n32652), .Z(n32637) );
  XOR U41543 ( .A(n32648), .B(n32647), .Z(n32652) );
  XOR U41544 ( .A(y[3516]), .B(x[3516]), .Z(n32647) );
  XOR U41545 ( .A(n32650), .B(n32649), .Z(n32648) );
  XOR U41546 ( .A(y[3518]), .B(x[3518]), .Z(n32649) );
  XOR U41547 ( .A(y[3517]), .B(x[3517]), .Z(n32650) );
  XOR U41548 ( .A(n32642), .B(n32641), .Z(n32651) );
  XOR U41549 ( .A(n32644), .B(n32643), .Z(n32641) );
  XOR U41550 ( .A(y[3515]), .B(x[3515]), .Z(n32643) );
  XOR U41551 ( .A(y[3514]), .B(x[3514]), .Z(n32644) );
  XOR U41552 ( .A(y[3513]), .B(x[3513]), .Z(n32642) );
  XNOR U41553 ( .A(n32635), .B(n32634), .Z(n32636) );
  XNOR U41554 ( .A(n32631), .B(n32630), .Z(n32634) );
  XOR U41555 ( .A(n32633), .B(n32632), .Z(n32630) );
  XOR U41556 ( .A(y[3512]), .B(x[3512]), .Z(n32632) );
  XOR U41557 ( .A(y[3511]), .B(x[3511]), .Z(n32633) );
  XOR U41558 ( .A(y[3510]), .B(x[3510]), .Z(n32631) );
  XOR U41559 ( .A(n32625), .B(n32624), .Z(n32635) );
  XOR U41560 ( .A(n32627), .B(n32626), .Z(n32624) );
  XOR U41561 ( .A(y[3509]), .B(x[3509]), .Z(n32626) );
  XOR U41562 ( .A(y[3508]), .B(x[3508]), .Z(n32627) );
  XOR U41563 ( .A(y[3507]), .B(x[3507]), .Z(n32625) );
  XNOR U41564 ( .A(n32601), .B(n32602), .Z(n32619) );
  XNOR U41565 ( .A(n32616), .B(n32617), .Z(n32602) );
  XOR U41566 ( .A(n32613), .B(n32612), .Z(n32617) );
  XOR U41567 ( .A(y[3504]), .B(x[3504]), .Z(n32612) );
  XOR U41568 ( .A(n32615), .B(n32614), .Z(n32613) );
  XOR U41569 ( .A(y[3506]), .B(x[3506]), .Z(n32614) );
  XOR U41570 ( .A(y[3505]), .B(x[3505]), .Z(n32615) );
  XOR U41571 ( .A(n32607), .B(n32606), .Z(n32616) );
  XOR U41572 ( .A(n32609), .B(n32608), .Z(n32606) );
  XOR U41573 ( .A(y[3503]), .B(x[3503]), .Z(n32608) );
  XOR U41574 ( .A(y[3502]), .B(x[3502]), .Z(n32609) );
  XOR U41575 ( .A(y[3501]), .B(x[3501]), .Z(n32607) );
  XNOR U41576 ( .A(n32600), .B(n32599), .Z(n32601) );
  XNOR U41577 ( .A(n32596), .B(n32595), .Z(n32599) );
  XOR U41578 ( .A(n32598), .B(n32597), .Z(n32595) );
  XOR U41579 ( .A(y[3500]), .B(x[3500]), .Z(n32597) );
  XOR U41580 ( .A(y[3499]), .B(x[3499]), .Z(n32598) );
  XOR U41581 ( .A(y[3498]), .B(x[3498]), .Z(n32596) );
  XOR U41582 ( .A(n32590), .B(n32589), .Z(n32600) );
  XOR U41583 ( .A(n32592), .B(n32591), .Z(n32589) );
  XOR U41584 ( .A(y[3497]), .B(x[3497]), .Z(n32591) );
  XOR U41585 ( .A(y[3496]), .B(x[3496]), .Z(n32592) );
  XOR U41586 ( .A(y[3495]), .B(x[3495]), .Z(n32590) );
  NAND U41587 ( .A(n32653), .B(n32654), .Z(N62481) );
  NAND U41588 ( .A(n32655), .B(n32656), .Z(n32654) );
  NANDN U41589 ( .A(n32657), .B(n32658), .Z(n32656) );
  NANDN U41590 ( .A(n32658), .B(n32657), .Z(n32653) );
  XOR U41591 ( .A(n32657), .B(n32659), .Z(N62480) );
  XNOR U41592 ( .A(n32655), .B(n32658), .Z(n32659) );
  NAND U41593 ( .A(n32660), .B(n32661), .Z(n32658) );
  NAND U41594 ( .A(n32662), .B(n32663), .Z(n32661) );
  NANDN U41595 ( .A(n32664), .B(n32665), .Z(n32663) );
  NANDN U41596 ( .A(n32665), .B(n32664), .Z(n32660) );
  AND U41597 ( .A(n32666), .B(n32667), .Z(n32655) );
  NAND U41598 ( .A(n32668), .B(n32669), .Z(n32667) );
  NANDN U41599 ( .A(n32670), .B(n32671), .Z(n32669) );
  NANDN U41600 ( .A(n32671), .B(n32670), .Z(n32666) );
  IV U41601 ( .A(n32672), .Z(n32671) );
  AND U41602 ( .A(n32673), .B(n32674), .Z(n32657) );
  NAND U41603 ( .A(n32675), .B(n32676), .Z(n32674) );
  NANDN U41604 ( .A(n32677), .B(n32678), .Z(n32676) );
  NANDN U41605 ( .A(n32678), .B(n32677), .Z(n32673) );
  XOR U41606 ( .A(n32670), .B(n32679), .Z(N62479) );
  XNOR U41607 ( .A(n32668), .B(n32672), .Z(n32679) );
  XOR U41608 ( .A(n32665), .B(n32680), .Z(n32672) );
  XNOR U41609 ( .A(n32662), .B(n32664), .Z(n32680) );
  AND U41610 ( .A(n32681), .B(n32682), .Z(n32664) );
  NANDN U41611 ( .A(n32683), .B(n32684), .Z(n32682) );
  OR U41612 ( .A(n32685), .B(n32686), .Z(n32684) );
  IV U41613 ( .A(n32687), .Z(n32686) );
  NANDN U41614 ( .A(n32687), .B(n32685), .Z(n32681) );
  AND U41615 ( .A(n32688), .B(n32689), .Z(n32662) );
  NAND U41616 ( .A(n32690), .B(n32691), .Z(n32689) );
  NANDN U41617 ( .A(n32692), .B(n32693), .Z(n32691) );
  NANDN U41618 ( .A(n32693), .B(n32692), .Z(n32688) );
  IV U41619 ( .A(n32694), .Z(n32693) );
  NAND U41620 ( .A(n32695), .B(n32696), .Z(n32665) );
  NANDN U41621 ( .A(n32697), .B(n32698), .Z(n32696) );
  NANDN U41622 ( .A(n32699), .B(n32700), .Z(n32698) );
  NANDN U41623 ( .A(n32700), .B(n32699), .Z(n32695) );
  IV U41624 ( .A(n32701), .Z(n32699) );
  AND U41625 ( .A(n32702), .B(n32703), .Z(n32668) );
  NAND U41626 ( .A(n32704), .B(n32705), .Z(n32703) );
  NANDN U41627 ( .A(n32706), .B(n32707), .Z(n32705) );
  NANDN U41628 ( .A(n32707), .B(n32706), .Z(n32702) );
  XOR U41629 ( .A(n32678), .B(n32708), .Z(n32670) );
  XNOR U41630 ( .A(n32675), .B(n32677), .Z(n32708) );
  AND U41631 ( .A(n32709), .B(n32710), .Z(n32677) );
  NANDN U41632 ( .A(n32711), .B(n32712), .Z(n32710) );
  OR U41633 ( .A(n32713), .B(n32714), .Z(n32712) );
  IV U41634 ( .A(n32715), .Z(n32714) );
  NANDN U41635 ( .A(n32715), .B(n32713), .Z(n32709) );
  AND U41636 ( .A(n32716), .B(n32717), .Z(n32675) );
  NAND U41637 ( .A(n32718), .B(n32719), .Z(n32717) );
  NANDN U41638 ( .A(n32720), .B(n32721), .Z(n32719) );
  NANDN U41639 ( .A(n32721), .B(n32720), .Z(n32716) );
  IV U41640 ( .A(n32722), .Z(n32721) );
  NAND U41641 ( .A(n32723), .B(n32724), .Z(n32678) );
  NANDN U41642 ( .A(n32725), .B(n32726), .Z(n32724) );
  NANDN U41643 ( .A(n32727), .B(n32728), .Z(n32726) );
  NANDN U41644 ( .A(n32728), .B(n32727), .Z(n32723) );
  IV U41645 ( .A(n32729), .Z(n32727) );
  XOR U41646 ( .A(n32704), .B(n32730), .Z(N62478) );
  XNOR U41647 ( .A(n32707), .B(n32706), .Z(n32730) );
  XNOR U41648 ( .A(n32718), .B(n32731), .Z(n32706) );
  XNOR U41649 ( .A(n32722), .B(n32720), .Z(n32731) );
  XOR U41650 ( .A(n32728), .B(n32732), .Z(n32720) );
  XNOR U41651 ( .A(n32725), .B(n32729), .Z(n32732) );
  AND U41652 ( .A(n32733), .B(n32734), .Z(n32729) );
  NAND U41653 ( .A(n32735), .B(n32736), .Z(n32734) );
  NAND U41654 ( .A(n32737), .B(n32738), .Z(n32733) );
  AND U41655 ( .A(n32739), .B(n32740), .Z(n32725) );
  NAND U41656 ( .A(n32741), .B(n32742), .Z(n32740) );
  NAND U41657 ( .A(n32743), .B(n32744), .Z(n32739) );
  NANDN U41658 ( .A(n32745), .B(n32746), .Z(n32728) );
  ANDN U41659 ( .B(n32747), .A(n32748), .Z(n32722) );
  XNOR U41660 ( .A(n32713), .B(n32749), .Z(n32718) );
  XNOR U41661 ( .A(n32711), .B(n32715), .Z(n32749) );
  AND U41662 ( .A(n32750), .B(n32751), .Z(n32715) );
  NAND U41663 ( .A(n32752), .B(n32753), .Z(n32751) );
  NAND U41664 ( .A(n32754), .B(n32755), .Z(n32750) );
  AND U41665 ( .A(n32756), .B(n32757), .Z(n32711) );
  NAND U41666 ( .A(n32758), .B(n32759), .Z(n32757) );
  NAND U41667 ( .A(n32760), .B(n32761), .Z(n32756) );
  AND U41668 ( .A(n32762), .B(n32763), .Z(n32713) );
  NAND U41669 ( .A(n32764), .B(n32765), .Z(n32707) );
  XNOR U41670 ( .A(n32690), .B(n32766), .Z(n32704) );
  XNOR U41671 ( .A(n32694), .B(n32692), .Z(n32766) );
  XOR U41672 ( .A(n32700), .B(n32767), .Z(n32692) );
  XNOR U41673 ( .A(n32697), .B(n32701), .Z(n32767) );
  AND U41674 ( .A(n32768), .B(n32769), .Z(n32701) );
  NAND U41675 ( .A(n32770), .B(n32771), .Z(n32769) );
  NAND U41676 ( .A(n32772), .B(n32773), .Z(n32768) );
  AND U41677 ( .A(n32774), .B(n32775), .Z(n32697) );
  NAND U41678 ( .A(n32776), .B(n32777), .Z(n32775) );
  NAND U41679 ( .A(n32778), .B(n32779), .Z(n32774) );
  NANDN U41680 ( .A(n32780), .B(n32781), .Z(n32700) );
  ANDN U41681 ( .B(n32782), .A(n32783), .Z(n32694) );
  XNOR U41682 ( .A(n32685), .B(n32784), .Z(n32690) );
  XNOR U41683 ( .A(n32683), .B(n32687), .Z(n32784) );
  AND U41684 ( .A(n32785), .B(n32786), .Z(n32687) );
  NAND U41685 ( .A(n32787), .B(n32788), .Z(n32786) );
  NAND U41686 ( .A(n32789), .B(n32790), .Z(n32785) );
  AND U41687 ( .A(n32791), .B(n32792), .Z(n32683) );
  NAND U41688 ( .A(n32793), .B(n32794), .Z(n32792) );
  NAND U41689 ( .A(n32795), .B(n32796), .Z(n32791) );
  AND U41690 ( .A(n32797), .B(n32798), .Z(n32685) );
  XOR U41691 ( .A(n32765), .B(n32764), .Z(N62477) );
  XNOR U41692 ( .A(n32782), .B(n32783), .Z(n32764) );
  XNOR U41693 ( .A(n32797), .B(n32798), .Z(n32783) );
  XOR U41694 ( .A(n32794), .B(n32793), .Z(n32798) );
  XOR U41695 ( .A(y[3492]), .B(x[3492]), .Z(n32793) );
  XOR U41696 ( .A(n32796), .B(n32795), .Z(n32794) );
  XOR U41697 ( .A(y[3494]), .B(x[3494]), .Z(n32795) );
  XOR U41698 ( .A(y[3493]), .B(x[3493]), .Z(n32796) );
  XOR U41699 ( .A(n32788), .B(n32787), .Z(n32797) );
  XOR U41700 ( .A(n32790), .B(n32789), .Z(n32787) );
  XOR U41701 ( .A(y[3491]), .B(x[3491]), .Z(n32789) );
  XOR U41702 ( .A(y[3490]), .B(x[3490]), .Z(n32790) );
  XOR U41703 ( .A(y[3489]), .B(x[3489]), .Z(n32788) );
  XNOR U41704 ( .A(n32781), .B(n32780), .Z(n32782) );
  XNOR U41705 ( .A(n32777), .B(n32776), .Z(n32780) );
  XOR U41706 ( .A(n32779), .B(n32778), .Z(n32776) );
  XOR U41707 ( .A(y[3488]), .B(x[3488]), .Z(n32778) );
  XOR U41708 ( .A(y[3487]), .B(x[3487]), .Z(n32779) );
  XOR U41709 ( .A(y[3486]), .B(x[3486]), .Z(n32777) );
  XOR U41710 ( .A(n32771), .B(n32770), .Z(n32781) );
  XOR U41711 ( .A(n32773), .B(n32772), .Z(n32770) );
  XOR U41712 ( .A(y[3485]), .B(x[3485]), .Z(n32772) );
  XOR U41713 ( .A(y[3484]), .B(x[3484]), .Z(n32773) );
  XOR U41714 ( .A(y[3483]), .B(x[3483]), .Z(n32771) );
  XNOR U41715 ( .A(n32747), .B(n32748), .Z(n32765) );
  XNOR U41716 ( .A(n32762), .B(n32763), .Z(n32748) );
  XOR U41717 ( .A(n32759), .B(n32758), .Z(n32763) );
  XOR U41718 ( .A(y[3480]), .B(x[3480]), .Z(n32758) );
  XOR U41719 ( .A(n32761), .B(n32760), .Z(n32759) );
  XOR U41720 ( .A(y[3482]), .B(x[3482]), .Z(n32760) );
  XOR U41721 ( .A(y[3481]), .B(x[3481]), .Z(n32761) );
  XOR U41722 ( .A(n32753), .B(n32752), .Z(n32762) );
  XOR U41723 ( .A(n32755), .B(n32754), .Z(n32752) );
  XOR U41724 ( .A(y[3479]), .B(x[3479]), .Z(n32754) );
  XOR U41725 ( .A(y[3478]), .B(x[3478]), .Z(n32755) );
  XOR U41726 ( .A(y[3477]), .B(x[3477]), .Z(n32753) );
  XNOR U41727 ( .A(n32746), .B(n32745), .Z(n32747) );
  XNOR U41728 ( .A(n32742), .B(n32741), .Z(n32745) );
  XOR U41729 ( .A(n32744), .B(n32743), .Z(n32741) );
  XOR U41730 ( .A(y[3476]), .B(x[3476]), .Z(n32743) );
  XOR U41731 ( .A(y[3475]), .B(x[3475]), .Z(n32744) );
  XOR U41732 ( .A(y[3474]), .B(x[3474]), .Z(n32742) );
  XOR U41733 ( .A(n32736), .B(n32735), .Z(n32746) );
  XOR U41734 ( .A(n32738), .B(n32737), .Z(n32735) );
  XOR U41735 ( .A(y[3473]), .B(x[3473]), .Z(n32737) );
  XOR U41736 ( .A(y[3472]), .B(x[3472]), .Z(n32738) );
  XOR U41737 ( .A(y[3471]), .B(x[3471]), .Z(n32736) );
  NAND U41738 ( .A(n32799), .B(n32800), .Z(N62468) );
  NAND U41739 ( .A(n32801), .B(n32802), .Z(n32800) );
  NANDN U41740 ( .A(n32803), .B(n32804), .Z(n32802) );
  NANDN U41741 ( .A(n32804), .B(n32803), .Z(n32799) );
  XOR U41742 ( .A(n32803), .B(n32805), .Z(N62467) );
  XNOR U41743 ( .A(n32801), .B(n32804), .Z(n32805) );
  NAND U41744 ( .A(n32806), .B(n32807), .Z(n32804) );
  NAND U41745 ( .A(n32808), .B(n32809), .Z(n32807) );
  NANDN U41746 ( .A(n32810), .B(n32811), .Z(n32809) );
  NANDN U41747 ( .A(n32811), .B(n32810), .Z(n32806) );
  AND U41748 ( .A(n32812), .B(n32813), .Z(n32801) );
  NAND U41749 ( .A(n32814), .B(n32815), .Z(n32813) );
  NANDN U41750 ( .A(n32816), .B(n32817), .Z(n32815) );
  NANDN U41751 ( .A(n32817), .B(n32816), .Z(n32812) );
  IV U41752 ( .A(n32818), .Z(n32817) );
  AND U41753 ( .A(n32819), .B(n32820), .Z(n32803) );
  NAND U41754 ( .A(n32821), .B(n32822), .Z(n32820) );
  NANDN U41755 ( .A(n32823), .B(n32824), .Z(n32822) );
  NANDN U41756 ( .A(n32824), .B(n32823), .Z(n32819) );
  XOR U41757 ( .A(n32816), .B(n32825), .Z(N62466) );
  XNOR U41758 ( .A(n32814), .B(n32818), .Z(n32825) );
  XOR U41759 ( .A(n32811), .B(n32826), .Z(n32818) );
  XNOR U41760 ( .A(n32808), .B(n32810), .Z(n32826) );
  AND U41761 ( .A(n32827), .B(n32828), .Z(n32810) );
  NANDN U41762 ( .A(n32829), .B(n32830), .Z(n32828) );
  OR U41763 ( .A(n32831), .B(n32832), .Z(n32830) );
  IV U41764 ( .A(n32833), .Z(n32832) );
  NANDN U41765 ( .A(n32833), .B(n32831), .Z(n32827) );
  AND U41766 ( .A(n32834), .B(n32835), .Z(n32808) );
  NAND U41767 ( .A(n32836), .B(n32837), .Z(n32835) );
  NANDN U41768 ( .A(n32838), .B(n32839), .Z(n32837) );
  NANDN U41769 ( .A(n32839), .B(n32838), .Z(n32834) );
  IV U41770 ( .A(n32840), .Z(n32839) );
  NAND U41771 ( .A(n32841), .B(n32842), .Z(n32811) );
  NANDN U41772 ( .A(n32843), .B(n32844), .Z(n32842) );
  NANDN U41773 ( .A(n32845), .B(n32846), .Z(n32844) );
  NANDN U41774 ( .A(n32846), .B(n32845), .Z(n32841) );
  IV U41775 ( .A(n32847), .Z(n32845) );
  AND U41776 ( .A(n32848), .B(n32849), .Z(n32814) );
  NAND U41777 ( .A(n32850), .B(n32851), .Z(n32849) );
  NANDN U41778 ( .A(n32852), .B(n32853), .Z(n32851) );
  NANDN U41779 ( .A(n32853), .B(n32852), .Z(n32848) );
  XOR U41780 ( .A(n32824), .B(n32854), .Z(n32816) );
  XNOR U41781 ( .A(n32821), .B(n32823), .Z(n32854) );
  AND U41782 ( .A(n32855), .B(n32856), .Z(n32823) );
  NANDN U41783 ( .A(n32857), .B(n32858), .Z(n32856) );
  OR U41784 ( .A(n32859), .B(n32860), .Z(n32858) );
  IV U41785 ( .A(n32861), .Z(n32860) );
  NANDN U41786 ( .A(n32861), .B(n32859), .Z(n32855) );
  AND U41787 ( .A(n32862), .B(n32863), .Z(n32821) );
  NAND U41788 ( .A(n32864), .B(n32865), .Z(n32863) );
  NANDN U41789 ( .A(n32866), .B(n32867), .Z(n32865) );
  NANDN U41790 ( .A(n32867), .B(n32866), .Z(n32862) );
  IV U41791 ( .A(n32868), .Z(n32867) );
  NAND U41792 ( .A(n32869), .B(n32870), .Z(n32824) );
  NANDN U41793 ( .A(n32871), .B(n32872), .Z(n32870) );
  NANDN U41794 ( .A(n32873), .B(n32874), .Z(n32872) );
  NANDN U41795 ( .A(n32874), .B(n32873), .Z(n32869) );
  IV U41796 ( .A(n32875), .Z(n32873) );
  XOR U41797 ( .A(n32850), .B(n32876), .Z(N62465) );
  XNOR U41798 ( .A(n32853), .B(n32852), .Z(n32876) );
  XNOR U41799 ( .A(n32864), .B(n32877), .Z(n32852) );
  XNOR U41800 ( .A(n32868), .B(n32866), .Z(n32877) );
  XOR U41801 ( .A(n32874), .B(n32878), .Z(n32866) );
  XNOR U41802 ( .A(n32871), .B(n32875), .Z(n32878) );
  AND U41803 ( .A(n32879), .B(n32880), .Z(n32875) );
  NAND U41804 ( .A(n32881), .B(n32882), .Z(n32880) );
  NAND U41805 ( .A(n32883), .B(n32884), .Z(n32879) );
  AND U41806 ( .A(n32885), .B(n32886), .Z(n32871) );
  NAND U41807 ( .A(n32887), .B(n32888), .Z(n32886) );
  NAND U41808 ( .A(n32889), .B(n32890), .Z(n32885) );
  NANDN U41809 ( .A(n32891), .B(n32892), .Z(n32874) );
  ANDN U41810 ( .B(n32893), .A(n32894), .Z(n32868) );
  XNOR U41811 ( .A(n32859), .B(n32895), .Z(n32864) );
  XNOR U41812 ( .A(n32857), .B(n32861), .Z(n32895) );
  AND U41813 ( .A(n32896), .B(n32897), .Z(n32861) );
  NAND U41814 ( .A(n32898), .B(n32899), .Z(n32897) );
  NAND U41815 ( .A(n32900), .B(n32901), .Z(n32896) );
  AND U41816 ( .A(n32902), .B(n32903), .Z(n32857) );
  NAND U41817 ( .A(n32904), .B(n32905), .Z(n32903) );
  NAND U41818 ( .A(n32906), .B(n32907), .Z(n32902) );
  AND U41819 ( .A(n32908), .B(n32909), .Z(n32859) );
  NAND U41820 ( .A(n32910), .B(n32911), .Z(n32853) );
  XNOR U41821 ( .A(n32836), .B(n32912), .Z(n32850) );
  XNOR U41822 ( .A(n32840), .B(n32838), .Z(n32912) );
  XOR U41823 ( .A(n32846), .B(n32913), .Z(n32838) );
  XNOR U41824 ( .A(n32843), .B(n32847), .Z(n32913) );
  AND U41825 ( .A(n32914), .B(n32915), .Z(n32847) );
  NAND U41826 ( .A(n32916), .B(n32917), .Z(n32915) );
  NAND U41827 ( .A(n32918), .B(n32919), .Z(n32914) );
  AND U41828 ( .A(n32920), .B(n32921), .Z(n32843) );
  NAND U41829 ( .A(n32922), .B(n32923), .Z(n32921) );
  NAND U41830 ( .A(n32924), .B(n32925), .Z(n32920) );
  NANDN U41831 ( .A(n32926), .B(n32927), .Z(n32846) );
  ANDN U41832 ( .B(n32928), .A(n32929), .Z(n32840) );
  XNOR U41833 ( .A(n32831), .B(n32930), .Z(n32836) );
  XNOR U41834 ( .A(n32829), .B(n32833), .Z(n32930) );
  AND U41835 ( .A(n32931), .B(n32932), .Z(n32833) );
  NAND U41836 ( .A(n32933), .B(n32934), .Z(n32932) );
  NAND U41837 ( .A(n32935), .B(n32936), .Z(n32931) );
  AND U41838 ( .A(n32937), .B(n32938), .Z(n32829) );
  NAND U41839 ( .A(n32939), .B(n32940), .Z(n32938) );
  NAND U41840 ( .A(n32941), .B(n32942), .Z(n32937) );
  AND U41841 ( .A(n32943), .B(n32944), .Z(n32831) );
  XOR U41842 ( .A(n32911), .B(n32910), .Z(N62464) );
  XNOR U41843 ( .A(n32928), .B(n32929), .Z(n32910) );
  XNOR U41844 ( .A(n32943), .B(n32944), .Z(n32929) );
  XOR U41845 ( .A(n32940), .B(n32939), .Z(n32944) );
  XOR U41846 ( .A(y[3468]), .B(x[3468]), .Z(n32939) );
  XOR U41847 ( .A(n32942), .B(n32941), .Z(n32940) );
  XOR U41848 ( .A(y[3470]), .B(x[3470]), .Z(n32941) );
  XOR U41849 ( .A(y[3469]), .B(x[3469]), .Z(n32942) );
  XOR U41850 ( .A(n32934), .B(n32933), .Z(n32943) );
  XOR U41851 ( .A(n32936), .B(n32935), .Z(n32933) );
  XOR U41852 ( .A(y[3467]), .B(x[3467]), .Z(n32935) );
  XOR U41853 ( .A(y[3466]), .B(x[3466]), .Z(n32936) );
  XOR U41854 ( .A(y[3465]), .B(x[3465]), .Z(n32934) );
  XNOR U41855 ( .A(n32927), .B(n32926), .Z(n32928) );
  XNOR U41856 ( .A(n32923), .B(n32922), .Z(n32926) );
  XOR U41857 ( .A(n32925), .B(n32924), .Z(n32922) );
  XOR U41858 ( .A(y[3464]), .B(x[3464]), .Z(n32924) );
  XOR U41859 ( .A(y[3463]), .B(x[3463]), .Z(n32925) );
  XOR U41860 ( .A(y[3462]), .B(x[3462]), .Z(n32923) );
  XOR U41861 ( .A(n32917), .B(n32916), .Z(n32927) );
  XOR U41862 ( .A(n32919), .B(n32918), .Z(n32916) );
  XOR U41863 ( .A(y[3461]), .B(x[3461]), .Z(n32918) );
  XOR U41864 ( .A(y[3460]), .B(x[3460]), .Z(n32919) );
  XOR U41865 ( .A(y[3459]), .B(x[3459]), .Z(n32917) );
  XNOR U41866 ( .A(n32893), .B(n32894), .Z(n32911) );
  XNOR U41867 ( .A(n32908), .B(n32909), .Z(n32894) );
  XOR U41868 ( .A(n32905), .B(n32904), .Z(n32909) );
  XOR U41869 ( .A(y[3456]), .B(x[3456]), .Z(n32904) );
  XOR U41870 ( .A(n32907), .B(n32906), .Z(n32905) );
  XOR U41871 ( .A(y[3458]), .B(x[3458]), .Z(n32906) );
  XOR U41872 ( .A(y[3457]), .B(x[3457]), .Z(n32907) );
  XOR U41873 ( .A(n32899), .B(n32898), .Z(n32908) );
  XOR U41874 ( .A(n32901), .B(n32900), .Z(n32898) );
  XOR U41875 ( .A(y[3455]), .B(x[3455]), .Z(n32900) );
  XOR U41876 ( .A(y[3454]), .B(x[3454]), .Z(n32901) );
  XOR U41877 ( .A(y[3453]), .B(x[3453]), .Z(n32899) );
  XNOR U41878 ( .A(n32892), .B(n32891), .Z(n32893) );
  XNOR U41879 ( .A(n32888), .B(n32887), .Z(n32891) );
  XOR U41880 ( .A(n32890), .B(n32889), .Z(n32887) );
  XOR U41881 ( .A(y[3452]), .B(x[3452]), .Z(n32889) );
  XOR U41882 ( .A(y[3451]), .B(x[3451]), .Z(n32890) );
  XOR U41883 ( .A(y[3450]), .B(x[3450]), .Z(n32888) );
  XOR U41884 ( .A(n32882), .B(n32881), .Z(n32892) );
  XOR U41885 ( .A(n32884), .B(n32883), .Z(n32881) );
  XOR U41886 ( .A(y[3449]), .B(x[3449]), .Z(n32883) );
  XOR U41887 ( .A(y[3448]), .B(x[3448]), .Z(n32884) );
  XOR U41888 ( .A(y[3447]), .B(x[3447]), .Z(n32882) );
  NAND U41889 ( .A(n32945), .B(n32946), .Z(N62455) );
  NAND U41890 ( .A(n32947), .B(n32948), .Z(n32946) );
  NANDN U41891 ( .A(n32949), .B(n32950), .Z(n32948) );
  NANDN U41892 ( .A(n32950), .B(n32949), .Z(n32945) );
  XOR U41893 ( .A(n32949), .B(n32951), .Z(N62454) );
  XNOR U41894 ( .A(n32947), .B(n32950), .Z(n32951) );
  NAND U41895 ( .A(n32952), .B(n32953), .Z(n32950) );
  NAND U41896 ( .A(n32954), .B(n32955), .Z(n32953) );
  NANDN U41897 ( .A(n32956), .B(n32957), .Z(n32955) );
  NANDN U41898 ( .A(n32957), .B(n32956), .Z(n32952) );
  AND U41899 ( .A(n32958), .B(n32959), .Z(n32947) );
  NAND U41900 ( .A(n32960), .B(n32961), .Z(n32959) );
  NANDN U41901 ( .A(n32962), .B(n32963), .Z(n32961) );
  NANDN U41902 ( .A(n32963), .B(n32962), .Z(n32958) );
  IV U41903 ( .A(n32964), .Z(n32963) );
  AND U41904 ( .A(n32965), .B(n32966), .Z(n32949) );
  NAND U41905 ( .A(n32967), .B(n32968), .Z(n32966) );
  NANDN U41906 ( .A(n32969), .B(n32970), .Z(n32968) );
  NANDN U41907 ( .A(n32970), .B(n32969), .Z(n32965) );
  XOR U41908 ( .A(n32962), .B(n32971), .Z(N62453) );
  XNOR U41909 ( .A(n32960), .B(n32964), .Z(n32971) );
  XOR U41910 ( .A(n32957), .B(n32972), .Z(n32964) );
  XNOR U41911 ( .A(n32954), .B(n32956), .Z(n32972) );
  AND U41912 ( .A(n32973), .B(n32974), .Z(n32956) );
  NANDN U41913 ( .A(n32975), .B(n32976), .Z(n32974) );
  OR U41914 ( .A(n32977), .B(n32978), .Z(n32976) );
  IV U41915 ( .A(n32979), .Z(n32978) );
  NANDN U41916 ( .A(n32979), .B(n32977), .Z(n32973) );
  AND U41917 ( .A(n32980), .B(n32981), .Z(n32954) );
  NAND U41918 ( .A(n32982), .B(n32983), .Z(n32981) );
  NANDN U41919 ( .A(n32984), .B(n32985), .Z(n32983) );
  NANDN U41920 ( .A(n32985), .B(n32984), .Z(n32980) );
  IV U41921 ( .A(n32986), .Z(n32985) );
  NAND U41922 ( .A(n32987), .B(n32988), .Z(n32957) );
  NANDN U41923 ( .A(n32989), .B(n32990), .Z(n32988) );
  NANDN U41924 ( .A(n32991), .B(n32992), .Z(n32990) );
  NANDN U41925 ( .A(n32992), .B(n32991), .Z(n32987) );
  IV U41926 ( .A(n32993), .Z(n32991) );
  AND U41927 ( .A(n32994), .B(n32995), .Z(n32960) );
  NAND U41928 ( .A(n32996), .B(n32997), .Z(n32995) );
  NANDN U41929 ( .A(n32998), .B(n32999), .Z(n32997) );
  NANDN U41930 ( .A(n32999), .B(n32998), .Z(n32994) );
  XOR U41931 ( .A(n32970), .B(n33000), .Z(n32962) );
  XNOR U41932 ( .A(n32967), .B(n32969), .Z(n33000) );
  AND U41933 ( .A(n33001), .B(n33002), .Z(n32969) );
  NANDN U41934 ( .A(n33003), .B(n33004), .Z(n33002) );
  OR U41935 ( .A(n33005), .B(n33006), .Z(n33004) );
  IV U41936 ( .A(n33007), .Z(n33006) );
  NANDN U41937 ( .A(n33007), .B(n33005), .Z(n33001) );
  AND U41938 ( .A(n33008), .B(n33009), .Z(n32967) );
  NAND U41939 ( .A(n33010), .B(n33011), .Z(n33009) );
  NANDN U41940 ( .A(n33012), .B(n33013), .Z(n33011) );
  NANDN U41941 ( .A(n33013), .B(n33012), .Z(n33008) );
  IV U41942 ( .A(n33014), .Z(n33013) );
  NAND U41943 ( .A(n33015), .B(n33016), .Z(n32970) );
  NANDN U41944 ( .A(n33017), .B(n33018), .Z(n33016) );
  NANDN U41945 ( .A(n33019), .B(n33020), .Z(n33018) );
  NANDN U41946 ( .A(n33020), .B(n33019), .Z(n33015) );
  IV U41947 ( .A(n33021), .Z(n33019) );
  XOR U41948 ( .A(n32996), .B(n33022), .Z(N62452) );
  XNOR U41949 ( .A(n32999), .B(n32998), .Z(n33022) );
  XNOR U41950 ( .A(n33010), .B(n33023), .Z(n32998) );
  XNOR U41951 ( .A(n33014), .B(n33012), .Z(n33023) );
  XOR U41952 ( .A(n33020), .B(n33024), .Z(n33012) );
  XNOR U41953 ( .A(n33017), .B(n33021), .Z(n33024) );
  AND U41954 ( .A(n33025), .B(n33026), .Z(n33021) );
  NAND U41955 ( .A(n33027), .B(n33028), .Z(n33026) );
  NAND U41956 ( .A(n33029), .B(n33030), .Z(n33025) );
  AND U41957 ( .A(n33031), .B(n33032), .Z(n33017) );
  NAND U41958 ( .A(n33033), .B(n33034), .Z(n33032) );
  NAND U41959 ( .A(n33035), .B(n33036), .Z(n33031) );
  NANDN U41960 ( .A(n33037), .B(n33038), .Z(n33020) );
  ANDN U41961 ( .B(n33039), .A(n33040), .Z(n33014) );
  XNOR U41962 ( .A(n33005), .B(n33041), .Z(n33010) );
  XNOR U41963 ( .A(n33003), .B(n33007), .Z(n33041) );
  AND U41964 ( .A(n33042), .B(n33043), .Z(n33007) );
  NAND U41965 ( .A(n33044), .B(n33045), .Z(n33043) );
  NAND U41966 ( .A(n33046), .B(n33047), .Z(n33042) );
  AND U41967 ( .A(n33048), .B(n33049), .Z(n33003) );
  NAND U41968 ( .A(n33050), .B(n33051), .Z(n33049) );
  NAND U41969 ( .A(n33052), .B(n33053), .Z(n33048) );
  AND U41970 ( .A(n33054), .B(n33055), .Z(n33005) );
  NAND U41971 ( .A(n33056), .B(n33057), .Z(n32999) );
  XNOR U41972 ( .A(n32982), .B(n33058), .Z(n32996) );
  XNOR U41973 ( .A(n32986), .B(n32984), .Z(n33058) );
  XOR U41974 ( .A(n32992), .B(n33059), .Z(n32984) );
  XNOR U41975 ( .A(n32989), .B(n32993), .Z(n33059) );
  AND U41976 ( .A(n33060), .B(n33061), .Z(n32993) );
  NAND U41977 ( .A(n33062), .B(n33063), .Z(n33061) );
  NAND U41978 ( .A(n33064), .B(n33065), .Z(n33060) );
  AND U41979 ( .A(n33066), .B(n33067), .Z(n32989) );
  NAND U41980 ( .A(n33068), .B(n33069), .Z(n33067) );
  NAND U41981 ( .A(n33070), .B(n33071), .Z(n33066) );
  NANDN U41982 ( .A(n33072), .B(n33073), .Z(n32992) );
  ANDN U41983 ( .B(n33074), .A(n33075), .Z(n32986) );
  XNOR U41984 ( .A(n32977), .B(n33076), .Z(n32982) );
  XNOR U41985 ( .A(n32975), .B(n32979), .Z(n33076) );
  AND U41986 ( .A(n33077), .B(n33078), .Z(n32979) );
  NAND U41987 ( .A(n33079), .B(n33080), .Z(n33078) );
  NAND U41988 ( .A(n33081), .B(n33082), .Z(n33077) );
  AND U41989 ( .A(n33083), .B(n33084), .Z(n32975) );
  NAND U41990 ( .A(n33085), .B(n33086), .Z(n33084) );
  NAND U41991 ( .A(n33087), .B(n33088), .Z(n33083) );
  AND U41992 ( .A(n33089), .B(n33090), .Z(n32977) );
  XOR U41993 ( .A(n33057), .B(n33056), .Z(N62451) );
  XNOR U41994 ( .A(n33074), .B(n33075), .Z(n33056) );
  XNOR U41995 ( .A(n33089), .B(n33090), .Z(n33075) );
  XOR U41996 ( .A(n33086), .B(n33085), .Z(n33090) );
  XOR U41997 ( .A(y[3444]), .B(x[3444]), .Z(n33085) );
  XOR U41998 ( .A(n33088), .B(n33087), .Z(n33086) );
  XOR U41999 ( .A(y[3446]), .B(x[3446]), .Z(n33087) );
  XOR U42000 ( .A(y[3445]), .B(x[3445]), .Z(n33088) );
  XOR U42001 ( .A(n33080), .B(n33079), .Z(n33089) );
  XOR U42002 ( .A(n33082), .B(n33081), .Z(n33079) );
  XOR U42003 ( .A(y[3443]), .B(x[3443]), .Z(n33081) );
  XOR U42004 ( .A(y[3442]), .B(x[3442]), .Z(n33082) );
  XOR U42005 ( .A(y[3441]), .B(x[3441]), .Z(n33080) );
  XNOR U42006 ( .A(n33073), .B(n33072), .Z(n33074) );
  XNOR U42007 ( .A(n33069), .B(n33068), .Z(n33072) );
  XOR U42008 ( .A(n33071), .B(n33070), .Z(n33068) );
  XOR U42009 ( .A(y[3440]), .B(x[3440]), .Z(n33070) );
  XOR U42010 ( .A(y[3439]), .B(x[3439]), .Z(n33071) );
  XOR U42011 ( .A(y[3438]), .B(x[3438]), .Z(n33069) );
  XOR U42012 ( .A(n33063), .B(n33062), .Z(n33073) );
  XOR U42013 ( .A(n33065), .B(n33064), .Z(n33062) );
  XOR U42014 ( .A(y[3437]), .B(x[3437]), .Z(n33064) );
  XOR U42015 ( .A(y[3436]), .B(x[3436]), .Z(n33065) );
  XOR U42016 ( .A(y[3435]), .B(x[3435]), .Z(n33063) );
  XNOR U42017 ( .A(n33039), .B(n33040), .Z(n33057) );
  XNOR U42018 ( .A(n33054), .B(n33055), .Z(n33040) );
  XOR U42019 ( .A(n33051), .B(n33050), .Z(n33055) );
  XOR U42020 ( .A(y[3432]), .B(x[3432]), .Z(n33050) );
  XOR U42021 ( .A(n33053), .B(n33052), .Z(n33051) );
  XOR U42022 ( .A(y[3434]), .B(x[3434]), .Z(n33052) );
  XOR U42023 ( .A(y[3433]), .B(x[3433]), .Z(n33053) );
  XOR U42024 ( .A(n33045), .B(n33044), .Z(n33054) );
  XOR U42025 ( .A(n33047), .B(n33046), .Z(n33044) );
  XOR U42026 ( .A(y[3431]), .B(x[3431]), .Z(n33046) );
  XOR U42027 ( .A(y[3430]), .B(x[3430]), .Z(n33047) );
  XOR U42028 ( .A(y[3429]), .B(x[3429]), .Z(n33045) );
  XNOR U42029 ( .A(n33038), .B(n33037), .Z(n33039) );
  XNOR U42030 ( .A(n33034), .B(n33033), .Z(n33037) );
  XOR U42031 ( .A(n33036), .B(n33035), .Z(n33033) );
  XOR U42032 ( .A(y[3428]), .B(x[3428]), .Z(n33035) );
  XOR U42033 ( .A(y[3427]), .B(x[3427]), .Z(n33036) );
  XOR U42034 ( .A(y[3426]), .B(x[3426]), .Z(n33034) );
  XOR U42035 ( .A(n33028), .B(n33027), .Z(n33038) );
  XOR U42036 ( .A(n33030), .B(n33029), .Z(n33027) );
  XOR U42037 ( .A(y[3425]), .B(x[3425]), .Z(n33029) );
  XOR U42038 ( .A(y[3424]), .B(x[3424]), .Z(n33030) );
  XOR U42039 ( .A(y[3423]), .B(x[3423]), .Z(n33028) );
  NAND U42040 ( .A(n33091), .B(n33092), .Z(N62442) );
  NAND U42041 ( .A(n33093), .B(n33094), .Z(n33092) );
  NANDN U42042 ( .A(n33095), .B(n33096), .Z(n33094) );
  NANDN U42043 ( .A(n33096), .B(n33095), .Z(n33091) );
  XOR U42044 ( .A(n33095), .B(n33097), .Z(N62441) );
  XNOR U42045 ( .A(n33093), .B(n33096), .Z(n33097) );
  NAND U42046 ( .A(n33098), .B(n33099), .Z(n33096) );
  NAND U42047 ( .A(n33100), .B(n33101), .Z(n33099) );
  NANDN U42048 ( .A(n33102), .B(n33103), .Z(n33101) );
  NANDN U42049 ( .A(n33103), .B(n33102), .Z(n33098) );
  AND U42050 ( .A(n33104), .B(n33105), .Z(n33093) );
  NAND U42051 ( .A(n33106), .B(n33107), .Z(n33105) );
  NANDN U42052 ( .A(n33108), .B(n33109), .Z(n33107) );
  NANDN U42053 ( .A(n33109), .B(n33108), .Z(n33104) );
  IV U42054 ( .A(n33110), .Z(n33109) );
  AND U42055 ( .A(n33111), .B(n33112), .Z(n33095) );
  NAND U42056 ( .A(n33113), .B(n33114), .Z(n33112) );
  NANDN U42057 ( .A(n33115), .B(n33116), .Z(n33114) );
  NANDN U42058 ( .A(n33116), .B(n33115), .Z(n33111) );
  XOR U42059 ( .A(n33108), .B(n33117), .Z(N62440) );
  XNOR U42060 ( .A(n33106), .B(n33110), .Z(n33117) );
  XOR U42061 ( .A(n33103), .B(n33118), .Z(n33110) );
  XNOR U42062 ( .A(n33100), .B(n33102), .Z(n33118) );
  AND U42063 ( .A(n33119), .B(n33120), .Z(n33102) );
  NANDN U42064 ( .A(n33121), .B(n33122), .Z(n33120) );
  OR U42065 ( .A(n33123), .B(n33124), .Z(n33122) );
  IV U42066 ( .A(n33125), .Z(n33124) );
  NANDN U42067 ( .A(n33125), .B(n33123), .Z(n33119) );
  AND U42068 ( .A(n33126), .B(n33127), .Z(n33100) );
  NAND U42069 ( .A(n33128), .B(n33129), .Z(n33127) );
  NANDN U42070 ( .A(n33130), .B(n33131), .Z(n33129) );
  NANDN U42071 ( .A(n33131), .B(n33130), .Z(n33126) );
  IV U42072 ( .A(n33132), .Z(n33131) );
  NAND U42073 ( .A(n33133), .B(n33134), .Z(n33103) );
  NANDN U42074 ( .A(n33135), .B(n33136), .Z(n33134) );
  NANDN U42075 ( .A(n33137), .B(n33138), .Z(n33136) );
  NANDN U42076 ( .A(n33138), .B(n33137), .Z(n33133) );
  IV U42077 ( .A(n33139), .Z(n33137) );
  AND U42078 ( .A(n33140), .B(n33141), .Z(n33106) );
  NAND U42079 ( .A(n33142), .B(n33143), .Z(n33141) );
  NANDN U42080 ( .A(n33144), .B(n33145), .Z(n33143) );
  NANDN U42081 ( .A(n33145), .B(n33144), .Z(n33140) );
  XOR U42082 ( .A(n33116), .B(n33146), .Z(n33108) );
  XNOR U42083 ( .A(n33113), .B(n33115), .Z(n33146) );
  AND U42084 ( .A(n33147), .B(n33148), .Z(n33115) );
  NANDN U42085 ( .A(n33149), .B(n33150), .Z(n33148) );
  OR U42086 ( .A(n33151), .B(n33152), .Z(n33150) );
  IV U42087 ( .A(n33153), .Z(n33152) );
  NANDN U42088 ( .A(n33153), .B(n33151), .Z(n33147) );
  AND U42089 ( .A(n33154), .B(n33155), .Z(n33113) );
  NAND U42090 ( .A(n33156), .B(n33157), .Z(n33155) );
  NANDN U42091 ( .A(n33158), .B(n33159), .Z(n33157) );
  NANDN U42092 ( .A(n33159), .B(n33158), .Z(n33154) );
  IV U42093 ( .A(n33160), .Z(n33159) );
  NAND U42094 ( .A(n33161), .B(n33162), .Z(n33116) );
  NANDN U42095 ( .A(n33163), .B(n33164), .Z(n33162) );
  NANDN U42096 ( .A(n33165), .B(n33166), .Z(n33164) );
  NANDN U42097 ( .A(n33166), .B(n33165), .Z(n33161) );
  IV U42098 ( .A(n33167), .Z(n33165) );
  XOR U42099 ( .A(n33142), .B(n33168), .Z(N62439) );
  XNOR U42100 ( .A(n33145), .B(n33144), .Z(n33168) );
  XNOR U42101 ( .A(n33156), .B(n33169), .Z(n33144) );
  XNOR U42102 ( .A(n33160), .B(n33158), .Z(n33169) );
  XOR U42103 ( .A(n33166), .B(n33170), .Z(n33158) );
  XNOR U42104 ( .A(n33163), .B(n33167), .Z(n33170) );
  AND U42105 ( .A(n33171), .B(n33172), .Z(n33167) );
  NAND U42106 ( .A(n33173), .B(n33174), .Z(n33172) );
  NAND U42107 ( .A(n33175), .B(n33176), .Z(n33171) );
  AND U42108 ( .A(n33177), .B(n33178), .Z(n33163) );
  NAND U42109 ( .A(n33179), .B(n33180), .Z(n33178) );
  NAND U42110 ( .A(n33181), .B(n33182), .Z(n33177) );
  NANDN U42111 ( .A(n33183), .B(n33184), .Z(n33166) );
  ANDN U42112 ( .B(n33185), .A(n33186), .Z(n33160) );
  XNOR U42113 ( .A(n33151), .B(n33187), .Z(n33156) );
  XNOR U42114 ( .A(n33149), .B(n33153), .Z(n33187) );
  AND U42115 ( .A(n33188), .B(n33189), .Z(n33153) );
  NAND U42116 ( .A(n33190), .B(n33191), .Z(n33189) );
  NAND U42117 ( .A(n33192), .B(n33193), .Z(n33188) );
  AND U42118 ( .A(n33194), .B(n33195), .Z(n33149) );
  NAND U42119 ( .A(n33196), .B(n33197), .Z(n33195) );
  NAND U42120 ( .A(n33198), .B(n33199), .Z(n33194) );
  AND U42121 ( .A(n33200), .B(n33201), .Z(n33151) );
  NAND U42122 ( .A(n33202), .B(n33203), .Z(n33145) );
  XNOR U42123 ( .A(n33128), .B(n33204), .Z(n33142) );
  XNOR U42124 ( .A(n33132), .B(n33130), .Z(n33204) );
  XOR U42125 ( .A(n33138), .B(n33205), .Z(n33130) );
  XNOR U42126 ( .A(n33135), .B(n33139), .Z(n33205) );
  AND U42127 ( .A(n33206), .B(n33207), .Z(n33139) );
  NAND U42128 ( .A(n33208), .B(n33209), .Z(n33207) );
  NAND U42129 ( .A(n33210), .B(n33211), .Z(n33206) );
  AND U42130 ( .A(n33212), .B(n33213), .Z(n33135) );
  NAND U42131 ( .A(n33214), .B(n33215), .Z(n33213) );
  NAND U42132 ( .A(n33216), .B(n33217), .Z(n33212) );
  NANDN U42133 ( .A(n33218), .B(n33219), .Z(n33138) );
  ANDN U42134 ( .B(n33220), .A(n33221), .Z(n33132) );
  XNOR U42135 ( .A(n33123), .B(n33222), .Z(n33128) );
  XNOR U42136 ( .A(n33121), .B(n33125), .Z(n33222) );
  AND U42137 ( .A(n33223), .B(n33224), .Z(n33125) );
  NAND U42138 ( .A(n33225), .B(n33226), .Z(n33224) );
  NAND U42139 ( .A(n33227), .B(n33228), .Z(n33223) );
  AND U42140 ( .A(n33229), .B(n33230), .Z(n33121) );
  NAND U42141 ( .A(n33231), .B(n33232), .Z(n33230) );
  NAND U42142 ( .A(n33233), .B(n33234), .Z(n33229) );
  AND U42143 ( .A(n33235), .B(n33236), .Z(n33123) );
  XOR U42144 ( .A(n33203), .B(n33202), .Z(N62438) );
  XNOR U42145 ( .A(n33220), .B(n33221), .Z(n33202) );
  XNOR U42146 ( .A(n33235), .B(n33236), .Z(n33221) );
  XOR U42147 ( .A(n33232), .B(n33231), .Z(n33236) );
  XOR U42148 ( .A(y[3420]), .B(x[3420]), .Z(n33231) );
  XOR U42149 ( .A(n33234), .B(n33233), .Z(n33232) );
  XOR U42150 ( .A(y[3422]), .B(x[3422]), .Z(n33233) );
  XOR U42151 ( .A(y[3421]), .B(x[3421]), .Z(n33234) );
  XOR U42152 ( .A(n33226), .B(n33225), .Z(n33235) );
  XOR U42153 ( .A(n33228), .B(n33227), .Z(n33225) );
  XOR U42154 ( .A(y[3419]), .B(x[3419]), .Z(n33227) );
  XOR U42155 ( .A(y[3418]), .B(x[3418]), .Z(n33228) );
  XOR U42156 ( .A(y[3417]), .B(x[3417]), .Z(n33226) );
  XNOR U42157 ( .A(n33219), .B(n33218), .Z(n33220) );
  XNOR U42158 ( .A(n33215), .B(n33214), .Z(n33218) );
  XOR U42159 ( .A(n33217), .B(n33216), .Z(n33214) );
  XOR U42160 ( .A(y[3416]), .B(x[3416]), .Z(n33216) );
  XOR U42161 ( .A(y[3415]), .B(x[3415]), .Z(n33217) );
  XOR U42162 ( .A(y[3414]), .B(x[3414]), .Z(n33215) );
  XOR U42163 ( .A(n33209), .B(n33208), .Z(n33219) );
  XOR U42164 ( .A(n33211), .B(n33210), .Z(n33208) );
  XOR U42165 ( .A(y[3413]), .B(x[3413]), .Z(n33210) );
  XOR U42166 ( .A(y[3412]), .B(x[3412]), .Z(n33211) );
  XOR U42167 ( .A(y[3411]), .B(x[3411]), .Z(n33209) );
  XNOR U42168 ( .A(n33185), .B(n33186), .Z(n33203) );
  XNOR U42169 ( .A(n33200), .B(n33201), .Z(n33186) );
  XOR U42170 ( .A(n33197), .B(n33196), .Z(n33201) );
  XOR U42171 ( .A(y[3408]), .B(x[3408]), .Z(n33196) );
  XOR U42172 ( .A(n33199), .B(n33198), .Z(n33197) );
  XOR U42173 ( .A(y[3410]), .B(x[3410]), .Z(n33198) );
  XOR U42174 ( .A(y[3409]), .B(x[3409]), .Z(n33199) );
  XOR U42175 ( .A(n33191), .B(n33190), .Z(n33200) );
  XOR U42176 ( .A(n33193), .B(n33192), .Z(n33190) );
  XOR U42177 ( .A(y[3407]), .B(x[3407]), .Z(n33192) );
  XOR U42178 ( .A(y[3406]), .B(x[3406]), .Z(n33193) );
  XOR U42179 ( .A(y[3405]), .B(x[3405]), .Z(n33191) );
  XNOR U42180 ( .A(n33184), .B(n33183), .Z(n33185) );
  XNOR U42181 ( .A(n33180), .B(n33179), .Z(n33183) );
  XOR U42182 ( .A(n33182), .B(n33181), .Z(n33179) );
  XOR U42183 ( .A(y[3404]), .B(x[3404]), .Z(n33181) );
  XOR U42184 ( .A(y[3403]), .B(x[3403]), .Z(n33182) );
  XOR U42185 ( .A(y[3402]), .B(x[3402]), .Z(n33180) );
  XOR U42186 ( .A(n33174), .B(n33173), .Z(n33184) );
  XOR U42187 ( .A(n33176), .B(n33175), .Z(n33173) );
  XOR U42188 ( .A(y[3401]), .B(x[3401]), .Z(n33175) );
  XOR U42189 ( .A(y[3400]), .B(x[3400]), .Z(n33176) );
  XOR U42190 ( .A(y[3399]), .B(x[3399]), .Z(n33174) );
  NAND U42191 ( .A(n33237), .B(n33238), .Z(N62429) );
  NAND U42192 ( .A(n33239), .B(n33240), .Z(n33238) );
  NANDN U42193 ( .A(n33241), .B(n33242), .Z(n33240) );
  NANDN U42194 ( .A(n33242), .B(n33241), .Z(n33237) );
  XOR U42195 ( .A(n33241), .B(n33243), .Z(N62428) );
  XNOR U42196 ( .A(n33239), .B(n33242), .Z(n33243) );
  NAND U42197 ( .A(n33244), .B(n33245), .Z(n33242) );
  NAND U42198 ( .A(n33246), .B(n33247), .Z(n33245) );
  NANDN U42199 ( .A(n33248), .B(n33249), .Z(n33247) );
  NANDN U42200 ( .A(n33249), .B(n33248), .Z(n33244) );
  AND U42201 ( .A(n33250), .B(n33251), .Z(n33239) );
  NAND U42202 ( .A(n33252), .B(n33253), .Z(n33251) );
  NANDN U42203 ( .A(n33254), .B(n33255), .Z(n33253) );
  NANDN U42204 ( .A(n33255), .B(n33254), .Z(n33250) );
  IV U42205 ( .A(n33256), .Z(n33255) );
  AND U42206 ( .A(n33257), .B(n33258), .Z(n33241) );
  NAND U42207 ( .A(n33259), .B(n33260), .Z(n33258) );
  NANDN U42208 ( .A(n33261), .B(n33262), .Z(n33260) );
  NANDN U42209 ( .A(n33262), .B(n33261), .Z(n33257) );
  XOR U42210 ( .A(n33254), .B(n33263), .Z(N62427) );
  XNOR U42211 ( .A(n33252), .B(n33256), .Z(n33263) );
  XOR U42212 ( .A(n33249), .B(n33264), .Z(n33256) );
  XNOR U42213 ( .A(n33246), .B(n33248), .Z(n33264) );
  AND U42214 ( .A(n33265), .B(n33266), .Z(n33248) );
  NANDN U42215 ( .A(n33267), .B(n33268), .Z(n33266) );
  OR U42216 ( .A(n33269), .B(n33270), .Z(n33268) );
  IV U42217 ( .A(n33271), .Z(n33270) );
  NANDN U42218 ( .A(n33271), .B(n33269), .Z(n33265) );
  AND U42219 ( .A(n33272), .B(n33273), .Z(n33246) );
  NAND U42220 ( .A(n33274), .B(n33275), .Z(n33273) );
  NANDN U42221 ( .A(n33276), .B(n33277), .Z(n33275) );
  NANDN U42222 ( .A(n33277), .B(n33276), .Z(n33272) );
  IV U42223 ( .A(n33278), .Z(n33277) );
  NAND U42224 ( .A(n33279), .B(n33280), .Z(n33249) );
  NANDN U42225 ( .A(n33281), .B(n33282), .Z(n33280) );
  NANDN U42226 ( .A(n33283), .B(n33284), .Z(n33282) );
  NANDN U42227 ( .A(n33284), .B(n33283), .Z(n33279) );
  IV U42228 ( .A(n33285), .Z(n33283) );
  AND U42229 ( .A(n33286), .B(n33287), .Z(n33252) );
  NAND U42230 ( .A(n33288), .B(n33289), .Z(n33287) );
  NANDN U42231 ( .A(n33290), .B(n33291), .Z(n33289) );
  NANDN U42232 ( .A(n33291), .B(n33290), .Z(n33286) );
  XOR U42233 ( .A(n33262), .B(n33292), .Z(n33254) );
  XNOR U42234 ( .A(n33259), .B(n33261), .Z(n33292) );
  AND U42235 ( .A(n33293), .B(n33294), .Z(n33261) );
  NANDN U42236 ( .A(n33295), .B(n33296), .Z(n33294) );
  OR U42237 ( .A(n33297), .B(n33298), .Z(n33296) );
  IV U42238 ( .A(n33299), .Z(n33298) );
  NANDN U42239 ( .A(n33299), .B(n33297), .Z(n33293) );
  AND U42240 ( .A(n33300), .B(n33301), .Z(n33259) );
  NAND U42241 ( .A(n33302), .B(n33303), .Z(n33301) );
  NANDN U42242 ( .A(n33304), .B(n33305), .Z(n33303) );
  NANDN U42243 ( .A(n33305), .B(n33304), .Z(n33300) );
  IV U42244 ( .A(n33306), .Z(n33305) );
  NAND U42245 ( .A(n33307), .B(n33308), .Z(n33262) );
  NANDN U42246 ( .A(n33309), .B(n33310), .Z(n33308) );
  NANDN U42247 ( .A(n33311), .B(n33312), .Z(n33310) );
  NANDN U42248 ( .A(n33312), .B(n33311), .Z(n33307) );
  IV U42249 ( .A(n33313), .Z(n33311) );
  XOR U42250 ( .A(n33288), .B(n33314), .Z(N62426) );
  XNOR U42251 ( .A(n33291), .B(n33290), .Z(n33314) );
  XNOR U42252 ( .A(n33302), .B(n33315), .Z(n33290) );
  XNOR U42253 ( .A(n33306), .B(n33304), .Z(n33315) );
  XOR U42254 ( .A(n33312), .B(n33316), .Z(n33304) );
  XNOR U42255 ( .A(n33309), .B(n33313), .Z(n33316) );
  AND U42256 ( .A(n33317), .B(n33318), .Z(n33313) );
  NAND U42257 ( .A(n33319), .B(n33320), .Z(n33318) );
  NAND U42258 ( .A(n33321), .B(n33322), .Z(n33317) );
  AND U42259 ( .A(n33323), .B(n33324), .Z(n33309) );
  NAND U42260 ( .A(n33325), .B(n33326), .Z(n33324) );
  NAND U42261 ( .A(n33327), .B(n33328), .Z(n33323) );
  NANDN U42262 ( .A(n33329), .B(n33330), .Z(n33312) );
  ANDN U42263 ( .B(n33331), .A(n33332), .Z(n33306) );
  XNOR U42264 ( .A(n33297), .B(n33333), .Z(n33302) );
  XNOR U42265 ( .A(n33295), .B(n33299), .Z(n33333) );
  AND U42266 ( .A(n33334), .B(n33335), .Z(n33299) );
  NAND U42267 ( .A(n33336), .B(n33337), .Z(n33335) );
  NAND U42268 ( .A(n33338), .B(n33339), .Z(n33334) );
  AND U42269 ( .A(n33340), .B(n33341), .Z(n33295) );
  NAND U42270 ( .A(n33342), .B(n33343), .Z(n33341) );
  NAND U42271 ( .A(n33344), .B(n33345), .Z(n33340) );
  AND U42272 ( .A(n33346), .B(n33347), .Z(n33297) );
  NAND U42273 ( .A(n33348), .B(n33349), .Z(n33291) );
  XNOR U42274 ( .A(n33274), .B(n33350), .Z(n33288) );
  XNOR U42275 ( .A(n33278), .B(n33276), .Z(n33350) );
  XOR U42276 ( .A(n33284), .B(n33351), .Z(n33276) );
  XNOR U42277 ( .A(n33281), .B(n33285), .Z(n33351) );
  AND U42278 ( .A(n33352), .B(n33353), .Z(n33285) );
  NAND U42279 ( .A(n33354), .B(n33355), .Z(n33353) );
  NAND U42280 ( .A(n33356), .B(n33357), .Z(n33352) );
  AND U42281 ( .A(n33358), .B(n33359), .Z(n33281) );
  NAND U42282 ( .A(n33360), .B(n33361), .Z(n33359) );
  NAND U42283 ( .A(n33362), .B(n33363), .Z(n33358) );
  NANDN U42284 ( .A(n33364), .B(n33365), .Z(n33284) );
  ANDN U42285 ( .B(n33366), .A(n33367), .Z(n33278) );
  XNOR U42286 ( .A(n33269), .B(n33368), .Z(n33274) );
  XNOR U42287 ( .A(n33267), .B(n33271), .Z(n33368) );
  AND U42288 ( .A(n33369), .B(n33370), .Z(n33271) );
  NAND U42289 ( .A(n33371), .B(n33372), .Z(n33370) );
  NAND U42290 ( .A(n33373), .B(n33374), .Z(n33369) );
  AND U42291 ( .A(n33375), .B(n33376), .Z(n33267) );
  NAND U42292 ( .A(n33377), .B(n33378), .Z(n33376) );
  NAND U42293 ( .A(n33379), .B(n33380), .Z(n33375) );
  AND U42294 ( .A(n33381), .B(n33382), .Z(n33269) );
  XOR U42295 ( .A(n33349), .B(n33348), .Z(N62425) );
  XNOR U42296 ( .A(n33366), .B(n33367), .Z(n33348) );
  XNOR U42297 ( .A(n33381), .B(n33382), .Z(n33367) );
  XOR U42298 ( .A(n33378), .B(n33377), .Z(n33382) );
  XOR U42299 ( .A(y[3396]), .B(x[3396]), .Z(n33377) );
  XOR U42300 ( .A(n33380), .B(n33379), .Z(n33378) );
  XOR U42301 ( .A(y[3398]), .B(x[3398]), .Z(n33379) );
  XOR U42302 ( .A(y[3397]), .B(x[3397]), .Z(n33380) );
  XOR U42303 ( .A(n33372), .B(n33371), .Z(n33381) );
  XOR U42304 ( .A(n33374), .B(n33373), .Z(n33371) );
  XOR U42305 ( .A(y[3395]), .B(x[3395]), .Z(n33373) );
  XOR U42306 ( .A(y[3394]), .B(x[3394]), .Z(n33374) );
  XOR U42307 ( .A(y[3393]), .B(x[3393]), .Z(n33372) );
  XNOR U42308 ( .A(n33365), .B(n33364), .Z(n33366) );
  XNOR U42309 ( .A(n33361), .B(n33360), .Z(n33364) );
  XOR U42310 ( .A(n33363), .B(n33362), .Z(n33360) );
  XOR U42311 ( .A(y[3392]), .B(x[3392]), .Z(n33362) );
  XOR U42312 ( .A(y[3391]), .B(x[3391]), .Z(n33363) );
  XOR U42313 ( .A(y[3390]), .B(x[3390]), .Z(n33361) );
  XOR U42314 ( .A(n33355), .B(n33354), .Z(n33365) );
  XOR U42315 ( .A(n33357), .B(n33356), .Z(n33354) );
  XOR U42316 ( .A(y[3389]), .B(x[3389]), .Z(n33356) );
  XOR U42317 ( .A(y[3388]), .B(x[3388]), .Z(n33357) );
  XOR U42318 ( .A(y[3387]), .B(x[3387]), .Z(n33355) );
  XNOR U42319 ( .A(n33331), .B(n33332), .Z(n33349) );
  XNOR U42320 ( .A(n33346), .B(n33347), .Z(n33332) );
  XOR U42321 ( .A(n33343), .B(n33342), .Z(n33347) );
  XOR U42322 ( .A(y[3384]), .B(x[3384]), .Z(n33342) );
  XOR U42323 ( .A(n33345), .B(n33344), .Z(n33343) );
  XOR U42324 ( .A(y[3386]), .B(x[3386]), .Z(n33344) );
  XOR U42325 ( .A(y[3385]), .B(x[3385]), .Z(n33345) );
  XOR U42326 ( .A(n33337), .B(n33336), .Z(n33346) );
  XOR U42327 ( .A(n33339), .B(n33338), .Z(n33336) );
  XOR U42328 ( .A(y[3383]), .B(x[3383]), .Z(n33338) );
  XOR U42329 ( .A(y[3382]), .B(x[3382]), .Z(n33339) );
  XOR U42330 ( .A(y[3381]), .B(x[3381]), .Z(n33337) );
  XNOR U42331 ( .A(n33330), .B(n33329), .Z(n33331) );
  XNOR U42332 ( .A(n33326), .B(n33325), .Z(n33329) );
  XOR U42333 ( .A(n33328), .B(n33327), .Z(n33325) );
  XOR U42334 ( .A(y[3380]), .B(x[3380]), .Z(n33327) );
  XOR U42335 ( .A(y[3379]), .B(x[3379]), .Z(n33328) );
  XOR U42336 ( .A(y[3378]), .B(x[3378]), .Z(n33326) );
  XOR U42337 ( .A(n33320), .B(n33319), .Z(n33330) );
  XOR U42338 ( .A(n33322), .B(n33321), .Z(n33319) );
  XOR U42339 ( .A(y[3377]), .B(x[3377]), .Z(n33321) );
  XOR U42340 ( .A(y[3376]), .B(x[3376]), .Z(n33322) );
  XOR U42341 ( .A(y[3375]), .B(x[3375]), .Z(n33320) );
  NAND U42342 ( .A(n33383), .B(n33384), .Z(N62416) );
  NAND U42343 ( .A(n33385), .B(n33386), .Z(n33384) );
  NANDN U42344 ( .A(n33387), .B(n33388), .Z(n33386) );
  NANDN U42345 ( .A(n33388), .B(n33387), .Z(n33383) );
  XOR U42346 ( .A(n33387), .B(n33389), .Z(N62415) );
  XNOR U42347 ( .A(n33385), .B(n33388), .Z(n33389) );
  NAND U42348 ( .A(n33390), .B(n33391), .Z(n33388) );
  NAND U42349 ( .A(n33392), .B(n33393), .Z(n33391) );
  NANDN U42350 ( .A(n33394), .B(n33395), .Z(n33393) );
  NANDN U42351 ( .A(n33395), .B(n33394), .Z(n33390) );
  AND U42352 ( .A(n33396), .B(n33397), .Z(n33385) );
  NAND U42353 ( .A(n33398), .B(n33399), .Z(n33397) );
  NANDN U42354 ( .A(n33400), .B(n33401), .Z(n33399) );
  NANDN U42355 ( .A(n33401), .B(n33400), .Z(n33396) );
  IV U42356 ( .A(n33402), .Z(n33401) );
  AND U42357 ( .A(n33403), .B(n33404), .Z(n33387) );
  NAND U42358 ( .A(n33405), .B(n33406), .Z(n33404) );
  NANDN U42359 ( .A(n33407), .B(n33408), .Z(n33406) );
  NANDN U42360 ( .A(n33408), .B(n33407), .Z(n33403) );
  XOR U42361 ( .A(n33400), .B(n33409), .Z(N62414) );
  XNOR U42362 ( .A(n33398), .B(n33402), .Z(n33409) );
  XOR U42363 ( .A(n33395), .B(n33410), .Z(n33402) );
  XNOR U42364 ( .A(n33392), .B(n33394), .Z(n33410) );
  AND U42365 ( .A(n33411), .B(n33412), .Z(n33394) );
  NANDN U42366 ( .A(n33413), .B(n33414), .Z(n33412) );
  OR U42367 ( .A(n33415), .B(n33416), .Z(n33414) );
  IV U42368 ( .A(n33417), .Z(n33416) );
  NANDN U42369 ( .A(n33417), .B(n33415), .Z(n33411) );
  AND U42370 ( .A(n33418), .B(n33419), .Z(n33392) );
  NAND U42371 ( .A(n33420), .B(n33421), .Z(n33419) );
  NANDN U42372 ( .A(n33422), .B(n33423), .Z(n33421) );
  NANDN U42373 ( .A(n33423), .B(n33422), .Z(n33418) );
  IV U42374 ( .A(n33424), .Z(n33423) );
  NAND U42375 ( .A(n33425), .B(n33426), .Z(n33395) );
  NANDN U42376 ( .A(n33427), .B(n33428), .Z(n33426) );
  NANDN U42377 ( .A(n33429), .B(n33430), .Z(n33428) );
  NANDN U42378 ( .A(n33430), .B(n33429), .Z(n33425) );
  IV U42379 ( .A(n33431), .Z(n33429) );
  AND U42380 ( .A(n33432), .B(n33433), .Z(n33398) );
  NAND U42381 ( .A(n33434), .B(n33435), .Z(n33433) );
  NANDN U42382 ( .A(n33436), .B(n33437), .Z(n33435) );
  NANDN U42383 ( .A(n33437), .B(n33436), .Z(n33432) );
  XOR U42384 ( .A(n33408), .B(n33438), .Z(n33400) );
  XNOR U42385 ( .A(n33405), .B(n33407), .Z(n33438) );
  AND U42386 ( .A(n33439), .B(n33440), .Z(n33407) );
  NANDN U42387 ( .A(n33441), .B(n33442), .Z(n33440) );
  OR U42388 ( .A(n33443), .B(n33444), .Z(n33442) );
  IV U42389 ( .A(n33445), .Z(n33444) );
  NANDN U42390 ( .A(n33445), .B(n33443), .Z(n33439) );
  AND U42391 ( .A(n33446), .B(n33447), .Z(n33405) );
  NAND U42392 ( .A(n33448), .B(n33449), .Z(n33447) );
  NANDN U42393 ( .A(n33450), .B(n33451), .Z(n33449) );
  NANDN U42394 ( .A(n33451), .B(n33450), .Z(n33446) );
  IV U42395 ( .A(n33452), .Z(n33451) );
  NAND U42396 ( .A(n33453), .B(n33454), .Z(n33408) );
  NANDN U42397 ( .A(n33455), .B(n33456), .Z(n33454) );
  NANDN U42398 ( .A(n33457), .B(n33458), .Z(n33456) );
  NANDN U42399 ( .A(n33458), .B(n33457), .Z(n33453) );
  IV U42400 ( .A(n33459), .Z(n33457) );
  XOR U42401 ( .A(n33434), .B(n33460), .Z(N62413) );
  XNOR U42402 ( .A(n33437), .B(n33436), .Z(n33460) );
  XNOR U42403 ( .A(n33448), .B(n33461), .Z(n33436) );
  XNOR U42404 ( .A(n33452), .B(n33450), .Z(n33461) );
  XOR U42405 ( .A(n33458), .B(n33462), .Z(n33450) );
  XNOR U42406 ( .A(n33455), .B(n33459), .Z(n33462) );
  AND U42407 ( .A(n33463), .B(n33464), .Z(n33459) );
  NAND U42408 ( .A(n33465), .B(n33466), .Z(n33464) );
  NAND U42409 ( .A(n33467), .B(n33468), .Z(n33463) );
  AND U42410 ( .A(n33469), .B(n33470), .Z(n33455) );
  NAND U42411 ( .A(n33471), .B(n33472), .Z(n33470) );
  NAND U42412 ( .A(n33473), .B(n33474), .Z(n33469) );
  NANDN U42413 ( .A(n33475), .B(n33476), .Z(n33458) );
  ANDN U42414 ( .B(n33477), .A(n33478), .Z(n33452) );
  XNOR U42415 ( .A(n33443), .B(n33479), .Z(n33448) );
  XNOR U42416 ( .A(n33441), .B(n33445), .Z(n33479) );
  AND U42417 ( .A(n33480), .B(n33481), .Z(n33445) );
  NAND U42418 ( .A(n33482), .B(n33483), .Z(n33481) );
  NAND U42419 ( .A(n33484), .B(n33485), .Z(n33480) );
  AND U42420 ( .A(n33486), .B(n33487), .Z(n33441) );
  NAND U42421 ( .A(n33488), .B(n33489), .Z(n33487) );
  NAND U42422 ( .A(n33490), .B(n33491), .Z(n33486) );
  AND U42423 ( .A(n33492), .B(n33493), .Z(n33443) );
  NAND U42424 ( .A(n33494), .B(n33495), .Z(n33437) );
  XNOR U42425 ( .A(n33420), .B(n33496), .Z(n33434) );
  XNOR U42426 ( .A(n33424), .B(n33422), .Z(n33496) );
  XOR U42427 ( .A(n33430), .B(n33497), .Z(n33422) );
  XNOR U42428 ( .A(n33427), .B(n33431), .Z(n33497) );
  AND U42429 ( .A(n33498), .B(n33499), .Z(n33431) );
  NAND U42430 ( .A(n33500), .B(n33501), .Z(n33499) );
  NAND U42431 ( .A(n33502), .B(n33503), .Z(n33498) );
  AND U42432 ( .A(n33504), .B(n33505), .Z(n33427) );
  NAND U42433 ( .A(n33506), .B(n33507), .Z(n33505) );
  NAND U42434 ( .A(n33508), .B(n33509), .Z(n33504) );
  NANDN U42435 ( .A(n33510), .B(n33511), .Z(n33430) );
  ANDN U42436 ( .B(n33512), .A(n33513), .Z(n33424) );
  XNOR U42437 ( .A(n33415), .B(n33514), .Z(n33420) );
  XNOR U42438 ( .A(n33413), .B(n33417), .Z(n33514) );
  AND U42439 ( .A(n33515), .B(n33516), .Z(n33417) );
  NAND U42440 ( .A(n33517), .B(n33518), .Z(n33516) );
  NAND U42441 ( .A(n33519), .B(n33520), .Z(n33515) );
  AND U42442 ( .A(n33521), .B(n33522), .Z(n33413) );
  NAND U42443 ( .A(n33523), .B(n33524), .Z(n33522) );
  NAND U42444 ( .A(n33525), .B(n33526), .Z(n33521) );
  AND U42445 ( .A(n33527), .B(n33528), .Z(n33415) );
  XOR U42446 ( .A(n33495), .B(n33494), .Z(N62412) );
  XNOR U42447 ( .A(n33512), .B(n33513), .Z(n33494) );
  XNOR U42448 ( .A(n33527), .B(n33528), .Z(n33513) );
  XOR U42449 ( .A(n33524), .B(n33523), .Z(n33528) );
  XOR U42450 ( .A(y[3372]), .B(x[3372]), .Z(n33523) );
  XOR U42451 ( .A(n33526), .B(n33525), .Z(n33524) );
  XOR U42452 ( .A(y[3374]), .B(x[3374]), .Z(n33525) );
  XOR U42453 ( .A(y[3373]), .B(x[3373]), .Z(n33526) );
  XOR U42454 ( .A(n33518), .B(n33517), .Z(n33527) );
  XOR U42455 ( .A(n33520), .B(n33519), .Z(n33517) );
  XOR U42456 ( .A(y[3371]), .B(x[3371]), .Z(n33519) );
  XOR U42457 ( .A(y[3370]), .B(x[3370]), .Z(n33520) );
  XOR U42458 ( .A(y[3369]), .B(x[3369]), .Z(n33518) );
  XNOR U42459 ( .A(n33511), .B(n33510), .Z(n33512) );
  XNOR U42460 ( .A(n33507), .B(n33506), .Z(n33510) );
  XOR U42461 ( .A(n33509), .B(n33508), .Z(n33506) );
  XOR U42462 ( .A(y[3368]), .B(x[3368]), .Z(n33508) );
  XOR U42463 ( .A(y[3367]), .B(x[3367]), .Z(n33509) );
  XOR U42464 ( .A(y[3366]), .B(x[3366]), .Z(n33507) );
  XOR U42465 ( .A(n33501), .B(n33500), .Z(n33511) );
  XOR U42466 ( .A(n33503), .B(n33502), .Z(n33500) );
  XOR U42467 ( .A(y[3365]), .B(x[3365]), .Z(n33502) );
  XOR U42468 ( .A(y[3364]), .B(x[3364]), .Z(n33503) );
  XOR U42469 ( .A(y[3363]), .B(x[3363]), .Z(n33501) );
  XNOR U42470 ( .A(n33477), .B(n33478), .Z(n33495) );
  XNOR U42471 ( .A(n33492), .B(n33493), .Z(n33478) );
  XOR U42472 ( .A(n33489), .B(n33488), .Z(n33493) );
  XOR U42473 ( .A(y[3360]), .B(x[3360]), .Z(n33488) );
  XOR U42474 ( .A(n33491), .B(n33490), .Z(n33489) );
  XOR U42475 ( .A(y[3362]), .B(x[3362]), .Z(n33490) );
  XOR U42476 ( .A(y[3361]), .B(x[3361]), .Z(n33491) );
  XOR U42477 ( .A(n33483), .B(n33482), .Z(n33492) );
  XOR U42478 ( .A(n33485), .B(n33484), .Z(n33482) );
  XOR U42479 ( .A(y[3359]), .B(x[3359]), .Z(n33484) );
  XOR U42480 ( .A(y[3358]), .B(x[3358]), .Z(n33485) );
  XOR U42481 ( .A(y[3357]), .B(x[3357]), .Z(n33483) );
  XNOR U42482 ( .A(n33476), .B(n33475), .Z(n33477) );
  XNOR U42483 ( .A(n33472), .B(n33471), .Z(n33475) );
  XOR U42484 ( .A(n33474), .B(n33473), .Z(n33471) );
  XOR U42485 ( .A(y[3356]), .B(x[3356]), .Z(n33473) );
  XOR U42486 ( .A(y[3355]), .B(x[3355]), .Z(n33474) );
  XOR U42487 ( .A(y[3354]), .B(x[3354]), .Z(n33472) );
  XOR U42488 ( .A(n33466), .B(n33465), .Z(n33476) );
  XOR U42489 ( .A(n33468), .B(n33467), .Z(n33465) );
  XOR U42490 ( .A(y[3353]), .B(x[3353]), .Z(n33467) );
  XOR U42491 ( .A(y[3352]), .B(x[3352]), .Z(n33468) );
  XOR U42492 ( .A(y[3351]), .B(x[3351]), .Z(n33466) );
  NAND U42493 ( .A(n33529), .B(n33530), .Z(N62403) );
  NAND U42494 ( .A(n33531), .B(n33532), .Z(n33530) );
  NANDN U42495 ( .A(n33533), .B(n33534), .Z(n33532) );
  NANDN U42496 ( .A(n33534), .B(n33533), .Z(n33529) );
  XOR U42497 ( .A(n33533), .B(n33535), .Z(N62402) );
  XNOR U42498 ( .A(n33531), .B(n33534), .Z(n33535) );
  NAND U42499 ( .A(n33536), .B(n33537), .Z(n33534) );
  NAND U42500 ( .A(n33538), .B(n33539), .Z(n33537) );
  NANDN U42501 ( .A(n33540), .B(n33541), .Z(n33539) );
  NANDN U42502 ( .A(n33541), .B(n33540), .Z(n33536) );
  AND U42503 ( .A(n33542), .B(n33543), .Z(n33531) );
  NAND U42504 ( .A(n33544), .B(n33545), .Z(n33543) );
  NANDN U42505 ( .A(n33546), .B(n33547), .Z(n33545) );
  NANDN U42506 ( .A(n33547), .B(n33546), .Z(n33542) );
  IV U42507 ( .A(n33548), .Z(n33547) );
  AND U42508 ( .A(n33549), .B(n33550), .Z(n33533) );
  NAND U42509 ( .A(n33551), .B(n33552), .Z(n33550) );
  NANDN U42510 ( .A(n33553), .B(n33554), .Z(n33552) );
  NANDN U42511 ( .A(n33554), .B(n33553), .Z(n33549) );
  XOR U42512 ( .A(n33546), .B(n33555), .Z(N62401) );
  XNOR U42513 ( .A(n33544), .B(n33548), .Z(n33555) );
  XOR U42514 ( .A(n33541), .B(n33556), .Z(n33548) );
  XNOR U42515 ( .A(n33538), .B(n33540), .Z(n33556) );
  AND U42516 ( .A(n33557), .B(n33558), .Z(n33540) );
  NANDN U42517 ( .A(n33559), .B(n33560), .Z(n33558) );
  OR U42518 ( .A(n33561), .B(n33562), .Z(n33560) );
  IV U42519 ( .A(n33563), .Z(n33562) );
  NANDN U42520 ( .A(n33563), .B(n33561), .Z(n33557) );
  AND U42521 ( .A(n33564), .B(n33565), .Z(n33538) );
  NAND U42522 ( .A(n33566), .B(n33567), .Z(n33565) );
  NANDN U42523 ( .A(n33568), .B(n33569), .Z(n33567) );
  NANDN U42524 ( .A(n33569), .B(n33568), .Z(n33564) );
  IV U42525 ( .A(n33570), .Z(n33569) );
  NAND U42526 ( .A(n33571), .B(n33572), .Z(n33541) );
  NANDN U42527 ( .A(n33573), .B(n33574), .Z(n33572) );
  NANDN U42528 ( .A(n33575), .B(n33576), .Z(n33574) );
  NANDN U42529 ( .A(n33576), .B(n33575), .Z(n33571) );
  IV U42530 ( .A(n33577), .Z(n33575) );
  AND U42531 ( .A(n33578), .B(n33579), .Z(n33544) );
  NAND U42532 ( .A(n33580), .B(n33581), .Z(n33579) );
  NANDN U42533 ( .A(n33582), .B(n33583), .Z(n33581) );
  NANDN U42534 ( .A(n33583), .B(n33582), .Z(n33578) );
  XOR U42535 ( .A(n33554), .B(n33584), .Z(n33546) );
  XNOR U42536 ( .A(n33551), .B(n33553), .Z(n33584) );
  AND U42537 ( .A(n33585), .B(n33586), .Z(n33553) );
  NANDN U42538 ( .A(n33587), .B(n33588), .Z(n33586) );
  OR U42539 ( .A(n33589), .B(n33590), .Z(n33588) );
  IV U42540 ( .A(n33591), .Z(n33590) );
  NANDN U42541 ( .A(n33591), .B(n33589), .Z(n33585) );
  AND U42542 ( .A(n33592), .B(n33593), .Z(n33551) );
  NAND U42543 ( .A(n33594), .B(n33595), .Z(n33593) );
  NANDN U42544 ( .A(n33596), .B(n33597), .Z(n33595) );
  NANDN U42545 ( .A(n33597), .B(n33596), .Z(n33592) );
  IV U42546 ( .A(n33598), .Z(n33597) );
  NAND U42547 ( .A(n33599), .B(n33600), .Z(n33554) );
  NANDN U42548 ( .A(n33601), .B(n33602), .Z(n33600) );
  NANDN U42549 ( .A(n33603), .B(n33604), .Z(n33602) );
  NANDN U42550 ( .A(n33604), .B(n33603), .Z(n33599) );
  IV U42551 ( .A(n33605), .Z(n33603) );
  XOR U42552 ( .A(n33580), .B(n33606), .Z(N62400) );
  XNOR U42553 ( .A(n33583), .B(n33582), .Z(n33606) );
  XNOR U42554 ( .A(n33594), .B(n33607), .Z(n33582) );
  XNOR U42555 ( .A(n33598), .B(n33596), .Z(n33607) );
  XOR U42556 ( .A(n33604), .B(n33608), .Z(n33596) );
  XNOR U42557 ( .A(n33601), .B(n33605), .Z(n33608) );
  AND U42558 ( .A(n33609), .B(n33610), .Z(n33605) );
  NAND U42559 ( .A(n33611), .B(n33612), .Z(n33610) );
  NAND U42560 ( .A(n33613), .B(n33614), .Z(n33609) );
  AND U42561 ( .A(n33615), .B(n33616), .Z(n33601) );
  NAND U42562 ( .A(n33617), .B(n33618), .Z(n33616) );
  NAND U42563 ( .A(n33619), .B(n33620), .Z(n33615) );
  NANDN U42564 ( .A(n33621), .B(n33622), .Z(n33604) );
  ANDN U42565 ( .B(n33623), .A(n33624), .Z(n33598) );
  XNOR U42566 ( .A(n33589), .B(n33625), .Z(n33594) );
  XNOR U42567 ( .A(n33587), .B(n33591), .Z(n33625) );
  AND U42568 ( .A(n33626), .B(n33627), .Z(n33591) );
  NAND U42569 ( .A(n33628), .B(n33629), .Z(n33627) );
  NAND U42570 ( .A(n33630), .B(n33631), .Z(n33626) );
  AND U42571 ( .A(n33632), .B(n33633), .Z(n33587) );
  NAND U42572 ( .A(n33634), .B(n33635), .Z(n33633) );
  NAND U42573 ( .A(n33636), .B(n33637), .Z(n33632) );
  AND U42574 ( .A(n33638), .B(n33639), .Z(n33589) );
  NAND U42575 ( .A(n33640), .B(n33641), .Z(n33583) );
  XNOR U42576 ( .A(n33566), .B(n33642), .Z(n33580) );
  XNOR U42577 ( .A(n33570), .B(n33568), .Z(n33642) );
  XOR U42578 ( .A(n33576), .B(n33643), .Z(n33568) );
  XNOR U42579 ( .A(n33573), .B(n33577), .Z(n33643) );
  AND U42580 ( .A(n33644), .B(n33645), .Z(n33577) );
  NAND U42581 ( .A(n33646), .B(n33647), .Z(n33645) );
  NAND U42582 ( .A(n33648), .B(n33649), .Z(n33644) );
  AND U42583 ( .A(n33650), .B(n33651), .Z(n33573) );
  NAND U42584 ( .A(n33652), .B(n33653), .Z(n33651) );
  NAND U42585 ( .A(n33654), .B(n33655), .Z(n33650) );
  NANDN U42586 ( .A(n33656), .B(n33657), .Z(n33576) );
  ANDN U42587 ( .B(n33658), .A(n33659), .Z(n33570) );
  XNOR U42588 ( .A(n33561), .B(n33660), .Z(n33566) );
  XNOR U42589 ( .A(n33559), .B(n33563), .Z(n33660) );
  AND U42590 ( .A(n33661), .B(n33662), .Z(n33563) );
  NAND U42591 ( .A(n33663), .B(n33664), .Z(n33662) );
  NAND U42592 ( .A(n33665), .B(n33666), .Z(n33661) );
  AND U42593 ( .A(n33667), .B(n33668), .Z(n33559) );
  NAND U42594 ( .A(n33669), .B(n33670), .Z(n33668) );
  NAND U42595 ( .A(n33671), .B(n33672), .Z(n33667) );
  AND U42596 ( .A(n33673), .B(n33674), .Z(n33561) );
  XOR U42597 ( .A(n33641), .B(n33640), .Z(N62399) );
  XNOR U42598 ( .A(n33658), .B(n33659), .Z(n33640) );
  XNOR U42599 ( .A(n33673), .B(n33674), .Z(n33659) );
  XOR U42600 ( .A(n33670), .B(n33669), .Z(n33674) );
  XOR U42601 ( .A(y[3348]), .B(x[3348]), .Z(n33669) );
  XOR U42602 ( .A(n33672), .B(n33671), .Z(n33670) );
  XOR U42603 ( .A(y[3350]), .B(x[3350]), .Z(n33671) );
  XOR U42604 ( .A(y[3349]), .B(x[3349]), .Z(n33672) );
  XOR U42605 ( .A(n33664), .B(n33663), .Z(n33673) );
  XOR U42606 ( .A(n33666), .B(n33665), .Z(n33663) );
  XOR U42607 ( .A(y[3347]), .B(x[3347]), .Z(n33665) );
  XOR U42608 ( .A(y[3346]), .B(x[3346]), .Z(n33666) );
  XOR U42609 ( .A(y[3345]), .B(x[3345]), .Z(n33664) );
  XNOR U42610 ( .A(n33657), .B(n33656), .Z(n33658) );
  XNOR U42611 ( .A(n33653), .B(n33652), .Z(n33656) );
  XOR U42612 ( .A(n33655), .B(n33654), .Z(n33652) );
  XOR U42613 ( .A(y[3344]), .B(x[3344]), .Z(n33654) );
  XOR U42614 ( .A(y[3343]), .B(x[3343]), .Z(n33655) );
  XOR U42615 ( .A(y[3342]), .B(x[3342]), .Z(n33653) );
  XOR U42616 ( .A(n33647), .B(n33646), .Z(n33657) );
  XOR U42617 ( .A(n33649), .B(n33648), .Z(n33646) );
  XOR U42618 ( .A(y[3341]), .B(x[3341]), .Z(n33648) );
  XOR U42619 ( .A(y[3340]), .B(x[3340]), .Z(n33649) );
  XOR U42620 ( .A(y[3339]), .B(x[3339]), .Z(n33647) );
  XNOR U42621 ( .A(n33623), .B(n33624), .Z(n33641) );
  XNOR U42622 ( .A(n33638), .B(n33639), .Z(n33624) );
  XOR U42623 ( .A(n33635), .B(n33634), .Z(n33639) );
  XOR U42624 ( .A(y[3336]), .B(x[3336]), .Z(n33634) );
  XOR U42625 ( .A(n33637), .B(n33636), .Z(n33635) );
  XOR U42626 ( .A(y[3338]), .B(x[3338]), .Z(n33636) );
  XOR U42627 ( .A(y[3337]), .B(x[3337]), .Z(n33637) );
  XOR U42628 ( .A(n33629), .B(n33628), .Z(n33638) );
  XOR U42629 ( .A(n33631), .B(n33630), .Z(n33628) );
  XOR U42630 ( .A(y[3335]), .B(x[3335]), .Z(n33630) );
  XOR U42631 ( .A(y[3334]), .B(x[3334]), .Z(n33631) );
  XOR U42632 ( .A(y[3333]), .B(x[3333]), .Z(n33629) );
  XNOR U42633 ( .A(n33622), .B(n33621), .Z(n33623) );
  XNOR U42634 ( .A(n33618), .B(n33617), .Z(n33621) );
  XOR U42635 ( .A(n33620), .B(n33619), .Z(n33617) );
  XOR U42636 ( .A(y[3332]), .B(x[3332]), .Z(n33619) );
  XOR U42637 ( .A(y[3331]), .B(x[3331]), .Z(n33620) );
  XOR U42638 ( .A(y[3330]), .B(x[3330]), .Z(n33618) );
  XOR U42639 ( .A(n33612), .B(n33611), .Z(n33622) );
  XOR U42640 ( .A(n33614), .B(n33613), .Z(n33611) );
  XOR U42641 ( .A(y[3329]), .B(x[3329]), .Z(n33613) );
  XOR U42642 ( .A(y[3328]), .B(x[3328]), .Z(n33614) );
  XOR U42643 ( .A(y[3327]), .B(x[3327]), .Z(n33612) );
  NAND U42644 ( .A(n33675), .B(n33676), .Z(N62390) );
  NAND U42645 ( .A(n33677), .B(n33678), .Z(n33676) );
  NANDN U42646 ( .A(n33679), .B(n33680), .Z(n33678) );
  NANDN U42647 ( .A(n33680), .B(n33679), .Z(n33675) );
  XOR U42648 ( .A(n33679), .B(n33681), .Z(N62389) );
  XNOR U42649 ( .A(n33677), .B(n33680), .Z(n33681) );
  NAND U42650 ( .A(n33682), .B(n33683), .Z(n33680) );
  NAND U42651 ( .A(n33684), .B(n33685), .Z(n33683) );
  NANDN U42652 ( .A(n33686), .B(n33687), .Z(n33685) );
  NANDN U42653 ( .A(n33687), .B(n33686), .Z(n33682) );
  AND U42654 ( .A(n33688), .B(n33689), .Z(n33677) );
  NAND U42655 ( .A(n33690), .B(n33691), .Z(n33689) );
  NANDN U42656 ( .A(n33692), .B(n33693), .Z(n33691) );
  NANDN U42657 ( .A(n33693), .B(n33692), .Z(n33688) );
  IV U42658 ( .A(n33694), .Z(n33693) );
  AND U42659 ( .A(n33695), .B(n33696), .Z(n33679) );
  NAND U42660 ( .A(n33697), .B(n33698), .Z(n33696) );
  NANDN U42661 ( .A(n33699), .B(n33700), .Z(n33698) );
  NANDN U42662 ( .A(n33700), .B(n33699), .Z(n33695) );
  XOR U42663 ( .A(n33692), .B(n33701), .Z(N62388) );
  XNOR U42664 ( .A(n33690), .B(n33694), .Z(n33701) );
  XOR U42665 ( .A(n33687), .B(n33702), .Z(n33694) );
  XNOR U42666 ( .A(n33684), .B(n33686), .Z(n33702) );
  AND U42667 ( .A(n33703), .B(n33704), .Z(n33686) );
  NANDN U42668 ( .A(n33705), .B(n33706), .Z(n33704) );
  OR U42669 ( .A(n33707), .B(n33708), .Z(n33706) );
  IV U42670 ( .A(n33709), .Z(n33708) );
  NANDN U42671 ( .A(n33709), .B(n33707), .Z(n33703) );
  AND U42672 ( .A(n33710), .B(n33711), .Z(n33684) );
  NAND U42673 ( .A(n33712), .B(n33713), .Z(n33711) );
  NANDN U42674 ( .A(n33714), .B(n33715), .Z(n33713) );
  NANDN U42675 ( .A(n33715), .B(n33714), .Z(n33710) );
  IV U42676 ( .A(n33716), .Z(n33715) );
  NAND U42677 ( .A(n33717), .B(n33718), .Z(n33687) );
  NANDN U42678 ( .A(n33719), .B(n33720), .Z(n33718) );
  NANDN U42679 ( .A(n33721), .B(n33722), .Z(n33720) );
  NANDN U42680 ( .A(n33722), .B(n33721), .Z(n33717) );
  IV U42681 ( .A(n33723), .Z(n33721) );
  AND U42682 ( .A(n33724), .B(n33725), .Z(n33690) );
  NAND U42683 ( .A(n33726), .B(n33727), .Z(n33725) );
  NANDN U42684 ( .A(n33728), .B(n33729), .Z(n33727) );
  NANDN U42685 ( .A(n33729), .B(n33728), .Z(n33724) );
  XOR U42686 ( .A(n33700), .B(n33730), .Z(n33692) );
  XNOR U42687 ( .A(n33697), .B(n33699), .Z(n33730) );
  AND U42688 ( .A(n33731), .B(n33732), .Z(n33699) );
  NANDN U42689 ( .A(n33733), .B(n33734), .Z(n33732) );
  OR U42690 ( .A(n33735), .B(n33736), .Z(n33734) );
  IV U42691 ( .A(n33737), .Z(n33736) );
  NANDN U42692 ( .A(n33737), .B(n33735), .Z(n33731) );
  AND U42693 ( .A(n33738), .B(n33739), .Z(n33697) );
  NAND U42694 ( .A(n33740), .B(n33741), .Z(n33739) );
  NANDN U42695 ( .A(n33742), .B(n33743), .Z(n33741) );
  NANDN U42696 ( .A(n33743), .B(n33742), .Z(n33738) );
  IV U42697 ( .A(n33744), .Z(n33743) );
  NAND U42698 ( .A(n33745), .B(n33746), .Z(n33700) );
  NANDN U42699 ( .A(n33747), .B(n33748), .Z(n33746) );
  NANDN U42700 ( .A(n33749), .B(n33750), .Z(n33748) );
  NANDN U42701 ( .A(n33750), .B(n33749), .Z(n33745) );
  IV U42702 ( .A(n33751), .Z(n33749) );
  XOR U42703 ( .A(n33726), .B(n33752), .Z(N62387) );
  XNOR U42704 ( .A(n33729), .B(n33728), .Z(n33752) );
  XNOR U42705 ( .A(n33740), .B(n33753), .Z(n33728) );
  XNOR U42706 ( .A(n33744), .B(n33742), .Z(n33753) );
  XOR U42707 ( .A(n33750), .B(n33754), .Z(n33742) );
  XNOR U42708 ( .A(n33747), .B(n33751), .Z(n33754) );
  AND U42709 ( .A(n33755), .B(n33756), .Z(n33751) );
  NAND U42710 ( .A(n33757), .B(n33758), .Z(n33756) );
  NAND U42711 ( .A(n33759), .B(n33760), .Z(n33755) );
  AND U42712 ( .A(n33761), .B(n33762), .Z(n33747) );
  NAND U42713 ( .A(n33763), .B(n33764), .Z(n33762) );
  NAND U42714 ( .A(n33765), .B(n33766), .Z(n33761) );
  NANDN U42715 ( .A(n33767), .B(n33768), .Z(n33750) );
  ANDN U42716 ( .B(n33769), .A(n33770), .Z(n33744) );
  XNOR U42717 ( .A(n33735), .B(n33771), .Z(n33740) );
  XNOR U42718 ( .A(n33733), .B(n33737), .Z(n33771) );
  AND U42719 ( .A(n33772), .B(n33773), .Z(n33737) );
  NAND U42720 ( .A(n33774), .B(n33775), .Z(n33773) );
  NAND U42721 ( .A(n33776), .B(n33777), .Z(n33772) );
  AND U42722 ( .A(n33778), .B(n33779), .Z(n33733) );
  NAND U42723 ( .A(n33780), .B(n33781), .Z(n33779) );
  NAND U42724 ( .A(n33782), .B(n33783), .Z(n33778) );
  AND U42725 ( .A(n33784), .B(n33785), .Z(n33735) );
  NAND U42726 ( .A(n33786), .B(n33787), .Z(n33729) );
  XNOR U42727 ( .A(n33712), .B(n33788), .Z(n33726) );
  XNOR U42728 ( .A(n33716), .B(n33714), .Z(n33788) );
  XOR U42729 ( .A(n33722), .B(n33789), .Z(n33714) );
  XNOR U42730 ( .A(n33719), .B(n33723), .Z(n33789) );
  AND U42731 ( .A(n33790), .B(n33791), .Z(n33723) );
  NAND U42732 ( .A(n33792), .B(n33793), .Z(n33791) );
  NAND U42733 ( .A(n33794), .B(n33795), .Z(n33790) );
  AND U42734 ( .A(n33796), .B(n33797), .Z(n33719) );
  NAND U42735 ( .A(n33798), .B(n33799), .Z(n33797) );
  NAND U42736 ( .A(n33800), .B(n33801), .Z(n33796) );
  NANDN U42737 ( .A(n33802), .B(n33803), .Z(n33722) );
  ANDN U42738 ( .B(n33804), .A(n33805), .Z(n33716) );
  XNOR U42739 ( .A(n33707), .B(n33806), .Z(n33712) );
  XNOR U42740 ( .A(n33705), .B(n33709), .Z(n33806) );
  AND U42741 ( .A(n33807), .B(n33808), .Z(n33709) );
  NAND U42742 ( .A(n33809), .B(n33810), .Z(n33808) );
  NAND U42743 ( .A(n33811), .B(n33812), .Z(n33807) );
  AND U42744 ( .A(n33813), .B(n33814), .Z(n33705) );
  NAND U42745 ( .A(n33815), .B(n33816), .Z(n33814) );
  NAND U42746 ( .A(n33817), .B(n33818), .Z(n33813) );
  AND U42747 ( .A(n33819), .B(n33820), .Z(n33707) );
  XOR U42748 ( .A(n33787), .B(n33786), .Z(N62386) );
  XNOR U42749 ( .A(n33804), .B(n33805), .Z(n33786) );
  XNOR U42750 ( .A(n33819), .B(n33820), .Z(n33805) );
  XOR U42751 ( .A(n33816), .B(n33815), .Z(n33820) );
  XOR U42752 ( .A(y[3324]), .B(x[3324]), .Z(n33815) );
  XOR U42753 ( .A(n33818), .B(n33817), .Z(n33816) );
  XOR U42754 ( .A(y[3326]), .B(x[3326]), .Z(n33817) );
  XOR U42755 ( .A(y[3325]), .B(x[3325]), .Z(n33818) );
  XOR U42756 ( .A(n33810), .B(n33809), .Z(n33819) );
  XOR U42757 ( .A(n33812), .B(n33811), .Z(n33809) );
  XOR U42758 ( .A(y[3323]), .B(x[3323]), .Z(n33811) );
  XOR U42759 ( .A(y[3322]), .B(x[3322]), .Z(n33812) );
  XOR U42760 ( .A(y[3321]), .B(x[3321]), .Z(n33810) );
  XNOR U42761 ( .A(n33803), .B(n33802), .Z(n33804) );
  XNOR U42762 ( .A(n33799), .B(n33798), .Z(n33802) );
  XOR U42763 ( .A(n33801), .B(n33800), .Z(n33798) );
  XOR U42764 ( .A(y[3320]), .B(x[3320]), .Z(n33800) );
  XOR U42765 ( .A(y[3319]), .B(x[3319]), .Z(n33801) );
  XOR U42766 ( .A(y[3318]), .B(x[3318]), .Z(n33799) );
  XOR U42767 ( .A(n33793), .B(n33792), .Z(n33803) );
  XOR U42768 ( .A(n33795), .B(n33794), .Z(n33792) );
  XOR U42769 ( .A(y[3317]), .B(x[3317]), .Z(n33794) );
  XOR U42770 ( .A(y[3316]), .B(x[3316]), .Z(n33795) );
  XOR U42771 ( .A(y[3315]), .B(x[3315]), .Z(n33793) );
  XNOR U42772 ( .A(n33769), .B(n33770), .Z(n33787) );
  XNOR U42773 ( .A(n33784), .B(n33785), .Z(n33770) );
  XOR U42774 ( .A(n33781), .B(n33780), .Z(n33785) );
  XOR U42775 ( .A(y[3312]), .B(x[3312]), .Z(n33780) );
  XOR U42776 ( .A(n33783), .B(n33782), .Z(n33781) );
  XOR U42777 ( .A(y[3314]), .B(x[3314]), .Z(n33782) );
  XOR U42778 ( .A(y[3313]), .B(x[3313]), .Z(n33783) );
  XOR U42779 ( .A(n33775), .B(n33774), .Z(n33784) );
  XOR U42780 ( .A(n33777), .B(n33776), .Z(n33774) );
  XOR U42781 ( .A(y[3311]), .B(x[3311]), .Z(n33776) );
  XOR U42782 ( .A(y[3310]), .B(x[3310]), .Z(n33777) );
  XOR U42783 ( .A(y[3309]), .B(x[3309]), .Z(n33775) );
  XNOR U42784 ( .A(n33768), .B(n33767), .Z(n33769) );
  XNOR U42785 ( .A(n33764), .B(n33763), .Z(n33767) );
  XOR U42786 ( .A(n33766), .B(n33765), .Z(n33763) );
  XOR U42787 ( .A(y[3308]), .B(x[3308]), .Z(n33765) );
  XOR U42788 ( .A(y[3307]), .B(x[3307]), .Z(n33766) );
  XOR U42789 ( .A(y[3306]), .B(x[3306]), .Z(n33764) );
  XOR U42790 ( .A(n33758), .B(n33757), .Z(n33768) );
  XOR U42791 ( .A(n33760), .B(n33759), .Z(n33757) );
  XOR U42792 ( .A(y[3305]), .B(x[3305]), .Z(n33759) );
  XOR U42793 ( .A(y[3304]), .B(x[3304]), .Z(n33760) );
  XOR U42794 ( .A(y[3303]), .B(x[3303]), .Z(n33758) );
  NAND U42795 ( .A(n33821), .B(n33822), .Z(N62377) );
  NAND U42796 ( .A(n33823), .B(n33824), .Z(n33822) );
  NANDN U42797 ( .A(n33825), .B(n33826), .Z(n33824) );
  NANDN U42798 ( .A(n33826), .B(n33825), .Z(n33821) );
  XOR U42799 ( .A(n33825), .B(n33827), .Z(N62376) );
  XNOR U42800 ( .A(n33823), .B(n33826), .Z(n33827) );
  NAND U42801 ( .A(n33828), .B(n33829), .Z(n33826) );
  NAND U42802 ( .A(n33830), .B(n33831), .Z(n33829) );
  NANDN U42803 ( .A(n33832), .B(n33833), .Z(n33831) );
  NANDN U42804 ( .A(n33833), .B(n33832), .Z(n33828) );
  AND U42805 ( .A(n33834), .B(n33835), .Z(n33823) );
  NAND U42806 ( .A(n33836), .B(n33837), .Z(n33835) );
  NANDN U42807 ( .A(n33838), .B(n33839), .Z(n33837) );
  NANDN U42808 ( .A(n33839), .B(n33838), .Z(n33834) );
  IV U42809 ( .A(n33840), .Z(n33839) );
  AND U42810 ( .A(n33841), .B(n33842), .Z(n33825) );
  NAND U42811 ( .A(n33843), .B(n33844), .Z(n33842) );
  NANDN U42812 ( .A(n33845), .B(n33846), .Z(n33844) );
  NANDN U42813 ( .A(n33846), .B(n33845), .Z(n33841) );
  XOR U42814 ( .A(n33838), .B(n33847), .Z(N62375) );
  XNOR U42815 ( .A(n33836), .B(n33840), .Z(n33847) );
  XOR U42816 ( .A(n33833), .B(n33848), .Z(n33840) );
  XNOR U42817 ( .A(n33830), .B(n33832), .Z(n33848) );
  AND U42818 ( .A(n33849), .B(n33850), .Z(n33832) );
  NANDN U42819 ( .A(n33851), .B(n33852), .Z(n33850) );
  OR U42820 ( .A(n33853), .B(n33854), .Z(n33852) );
  IV U42821 ( .A(n33855), .Z(n33854) );
  NANDN U42822 ( .A(n33855), .B(n33853), .Z(n33849) );
  AND U42823 ( .A(n33856), .B(n33857), .Z(n33830) );
  NAND U42824 ( .A(n33858), .B(n33859), .Z(n33857) );
  NANDN U42825 ( .A(n33860), .B(n33861), .Z(n33859) );
  NANDN U42826 ( .A(n33861), .B(n33860), .Z(n33856) );
  IV U42827 ( .A(n33862), .Z(n33861) );
  NAND U42828 ( .A(n33863), .B(n33864), .Z(n33833) );
  NANDN U42829 ( .A(n33865), .B(n33866), .Z(n33864) );
  NANDN U42830 ( .A(n33867), .B(n33868), .Z(n33866) );
  NANDN U42831 ( .A(n33868), .B(n33867), .Z(n33863) );
  IV U42832 ( .A(n33869), .Z(n33867) );
  AND U42833 ( .A(n33870), .B(n33871), .Z(n33836) );
  NAND U42834 ( .A(n33872), .B(n33873), .Z(n33871) );
  NANDN U42835 ( .A(n33874), .B(n33875), .Z(n33873) );
  NANDN U42836 ( .A(n33875), .B(n33874), .Z(n33870) );
  XOR U42837 ( .A(n33846), .B(n33876), .Z(n33838) );
  XNOR U42838 ( .A(n33843), .B(n33845), .Z(n33876) );
  AND U42839 ( .A(n33877), .B(n33878), .Z(n33845) );
  NANDN U42840 ( .A(n33879), .B(n33880), .Z(n33878) );
  OR U42841 ( .A(n33881), .B(n33882), .Z(n33880) );
  IV U42842 ( .A(n33883), .Z(n33882) );
  NANDN U42843 ( .A(n33883), .B(n33881), .Z(n33877) );
  AND U42844 ( .A(n33884), .B(n33885), .Z(n33843) );
  NAND U42845 ( .A(n33886), .B(n33887), .Z(n33885) );
  NANDN U42846 ( .A(n33888), .B(n33889), .Z(n33887) );
  NANDN U42847 ( .A(n33889), .B(n33888), .Z(n33884) );
  IV U42848 ( .A(n33890), .Z(n33889) );
  NAND U42849 ( .A(n33891), .B(n33892), .Z(n33846) );
  NANDN U42850 ( .A(n33893), .B(n33894), .Z(n33892) );
  NANDN U42851 ( .A(n33895), .B(n33896), .Z(n33894) );
  NANDN U42852 ( .A(n33896), .B(n33895), .Z(n33891) );
  IV U42853 ( .A(n33897), .Z(n33895) );
  XOR U42854 ( .A(n33872), .B(n33898), .Z(N62374) );
  XNOR U42855 ( .A(n33875), .B(n33874), .Z(n33898) );
  XNOR U42856 ( .A(n33886), .B(n33899), .Z(n33874) );
  XNOR U42857 ( .A(n33890), .B(n33888), .Z(n33899) );
  XOR U42858 ( .A(n33896), .B(n33900), .Z(n33888) );
  XNOR U42859 ( .A(n33893), .B(n33897), .Z(n33900) );
  AND U42860 ( .A(n33901), .B(n33902), .Z(n33897) );
  NAND U42861 ( .A(n33903), .B(n33904), .Z(n33902) );
  NAND U42862 ( .A(n33905), .B(n33906), .Z(n33901) );
  AND U42863 ( .A(n33907), .B(n33908), .Z(n33893) );
  NAND U42864 ( .A(n33909), .B(n33910), .Z(n33908) );
  NAND U42865 ( .A(n33911), .B(n33912), .Z(n33907) );
  NANDN U42866 ( .A(n33913), .B(n33914), .Z(n33896) );
  ANDN U42867 ( .B(n33915), .A(n33916), .Z(n33890) );
  XNOR U42868 ( .A(n33881), .B(n33917), .Z(n33886) );
  XNOR U42869 ( .A(n33879), .B(n33883), .Z(n33917) );
  AND U42870 ( .A(n33918), .B(n33919), .Z(n33883) );
  NAND U42871 ( .A(n33920), .B(n33921), .Z(n33919) );
  NAND U42872 ( .A(n33922), .B(n33923), .Z(n33918) );
  AND U42873 ( .A(n33924), .B(n33925), .Z(n33879) );
  NAND U42874 ( .A(n33926), .B(n33927), .Z(n33925) );
  NAND U42875 ( .A(n33928), .B(n33929), .Z(n33924) );
  AND U42876 ( .A(n33930), .B(n33931), .Z(n33881) );
  NAND U42877 ( .A(n33932), .B(n33933), .Z(n33875) );
  XNOR U42878 ( .A(n33858), .B(n33934), .Z(n33872) );
  XNOR U42879 ( .A(n33862), .B(n33860), .Z(n33934) );
  XOR U42880 ( .A(n33868), .B(n33935), .Z(n33860) );
  XNOR U42881 ( .A(n33865), .B(n33869), .Z(n33935) );
  AND U42882 ( .A(n33936), .B(n33937), .Z(n33869) );
  NAND U42883 ( .A(n33938), .B(n33939), .Z(n33937) );
  NAND U42884 ( .A(n33940), .B(n33941), .Z(n33936) );
  AND U42885 ( .A(n33942), .B(n33943), .Z(n33865) );
  NAND U42886 ( .A(n33944), .B(n33945), .Z(n33943) );
  NAND U42887 ( .A(n33946), .B(n33947), .Z(n33942) );
  NANDN U42888 ( .A(n33948), .B(n33949), .Z(n33868) );
  ANDN U42889 ( .B(n33950), .A(n33951), .Z(n33862) );
  XNOR U42890 ( .A(n33853), .B(n33952), .Z(n33858) );
  XNOR U42891 ( .A(n33851), .B(n33855), .Z(n33952) );
  AND U42892 ( .A(n33953), .B(n33954), .Z(n33855) );
  NAND U42893 ( .A(n33955), .B(n33956), .Z(n33954) );
  NAND U42894 ( .A(n33957), .B(n33958), .Z(n33953) );
  AND U42895 ( .A(n33959), .B(n33960), .Z(n33851) );
  NAND U42896 ( .A(n33961), .B(n33962), .Z(n33960) );
  NAND U42897 ( .A(n33963), .B(n33964), .Z(n33959) );
  AND U42898 ( .A(n33965), .B(n33966), .Z(n33853) );
  XOR U42899 ( .A(n33933), .B(n33932), .Z(N62373) );
  XNOR U42900 ( .A(n33950), .B(n33951), .Z(n33932) );
  XNOR U42901 ( .A(n33965), .B(n33966), .Z(n33951) );
  XOR U42902 ( .A(n33962), .B(n33961), .Z(n33966) );
  XOR U42903 ( .A(y[3300]), .B(x[3300]), .Z(n33961) );
  XOR U42904 ( .A(n33964), .B(n33963), .Z(n33962) );
  XOR U42905 ( .A(y[3302]), .B(x[3302]), .Z(n33963) );
  XOR U42906 ( .A(y[3301]), .B(x[3301]), .Z(n33964) );
  XOR U42907 ( .A(n33956), .B(n33955), .Z(n33965) );
  XOR U42908 ( .A(n33958), .B(n33957), .Z(n33955) );
  XOR U42909 ( .A(y[3299]), .B(x[3299]), .Z(n33957) );
  XOR U42910 ( .A(y[3298]), .B(x[3298]), .Z(n33958) );
  XOR U42911 ( .A(y[3297]), .B(x[3297]), .Z(n33956) );
  XNOR U42912 ( .A(n33949), .B(n33948), .Z(n33950) );
  XNOR U42913 ( .A(n33945), .B(n33944), .Z(n33948) );
  XOR U42914 ( .A(n33947), .B(n33946), .Z(n33944) );
  XOR U42915 ( .A(y[3296]), .B(x[3296]), .Z(n33946) );
  XOR U42916 ( .A(y[3295]), .B(x[3295]), .Z(n33947) );
  XOR U42917 ( .A(y[3294]), .B(x[3294]), .Z(n33945) );
  XOR U42918 ( .A(n33939), .B(n33938), .Z(n33949) );
  XOR U42919 ( .A(n33941), .B(n33940), .Z(n33938) );
  XOR U42920 ( .A(y[3293]), .B(x[3293]), .Z(n33940) );
  XOR U42921 ( .A(y[3292]), .B(x[3292]), .Z(n33941) );
  XOR U42922 ( .A(y[3291]), .B(x[3291]), .Z(n33939) );
  XNOR U42923 ( .A(n33915), .B(n33916), .Z(n33933) );
  XNOR U42924 ( .A(n33930), .B(n33931), .Z(n33916) );
  XOR U42925 ( .A(n33927), .B(n33926), .Z(n33931) );
  XOR U42926 ( .A(y[3288]), .B(x[3288]), .Z(n33926) );
  XOR U42927 ( .A(n33929), .B(n33928), .Z(n33927) );
  XOR U42928 ( .A(y[3290]), .B(x[3290]), .Z(n33928) );
  XOR U42929 ( .A(y[3289]), .B(x[3289]), .Z(n33929) );
  XOR U42930 ( .A(n33921), .B(n33920), .Z(n33930) );
  XOR U42931 ( .A(n33923), .B(n33922), .Z(n33920) );
  XOR U42932 ( .A(y[3287]), .B(x[3287]), .Z(n33922) );
  XOR U42933 ( .A(y[3286]), .B(x[3286]), .Z(n33923) );
  XOR U42934 ( .A(y[3285]), .B(x[3285]), .Z(n33921) );
  XNOR U42935 ( .A(n33914), .B(n33913), .Z(n33915) );
  XNOR U42936 ( .A(n33910), .B(n33909), .Z(n33913) );
  XOR U42937 ( .A(n33912), .B(n33911), .Z(n33909) );
  XOR U42938 ( .A(y[3284]), .B(x[3284]), .Z(n33911) );
  XOR U42939 ( .A(y[3283]), .B(x[3283]), .Z(n33912) );
  XOR U42940 ( .A(y[3282]), .B(x[3282]), .Z(n33910) );
  XOR U42941 ( .A(n33904), .B(n33903), .Z(n33914) );
  XOR U42942 ( .A(n33906), .B(n33905), .Z(n33903) );
  XOR U42943 ( .A(y[3281]), .B(x[3281]), .Z(n33905) );
  XOR U42944 ( .A(y[3280]), .B(x[3280]), .Z(n33906) );
  XOR U42945 ( .A(y[3279]), .B(x[3279]), .Z(n33904) );
  NAND U42946 ( .A(n33967), .B(n33968), .Z(N62364) );
  NAND U42947 ( .A(n33969), .B(n33970), .Z(n33968) );
  NANDN U42948 ( .A(n33971), .B(n33972), .Z(n33970) );
  NANDN U42949 ( .A(n33972), .B(n33971), .Z(n33967) );
  XOR U42950 ( .A(n33971), .B(n33973), .Z(N62363) );
  XNOR U42951 ( .A(n33969), .B(n33972), .Z(n33973) );
  NAND U42952 ( .A(n33974), .B(n33975), .Z(n33972) );
  NAND U42953 ( .A(n33976), .B(n33977), .Z(n33975) );
  NANDN U42954 ( .A(n33978), .B(n33979), .Z(n33977) );
  NANDN U42955 ( .A(n33979), .B(n33978), .Z(n33974) );
  AND U42956 ( .A(n33980), .B(n33981), .Z(n33969) );
  NAND U42957 ( .A(n33982), .B(n33983), .Z(n33981) );
  NANDN U42958 ( .A(n33984), .B(n33985), .Z(n33983) );
  NANDN U42959 ( .A(n33985), .B(n33984), .Z(n33980) );
  IV U42960 ( .A(n33986), .Z(n33985) );
  AND U42961 ( .A(n33987), .B(n33988), .Z(n33971) );
  NAND U42962 ( .A(n33989), .B(n33990), .Z(n33988) );
  NANDN U42963 ( .A(n33991), .B(n33992), .Z(n33990) );
  NANDN U42964 ( .A(n33992), .B(n33991), .Z(n33987) );
  XOR U42965 ( .A(n33984), .B(n33993), .Z(N62362) );
  XNOR U42966 ( .A(n33982), .B(n33986), .Z(n33993) );
  XOR U42967 ( .A(n33979), .B(n33994), .Z(n33986) );
  XNOR U42968 ( .A(n33976), .B(n33978), .Z(n33994) );
  AND U42969 ( .A(n33995), .B(n33996), .Z(n33978) );
  NANDN U42970 ( .A(n33997), .B(n33998), .Z(n33996) );
  OR U42971 ( .A(n33999), .B(n34000), .Z(n33998) );
  IV U42972 ( .A(n34001), .Z(n34000) );
  NANDN U42973 ( .A(n34001), .B(n33999), .Z(n33995) );
  AND U42974 ( .A(n34002), .B(n34003), .Z(n33976) );
  NAND U42975 ( .A(n34004), .B(n34005), .Z(n34003) );
  NANDN U42976 ( .A(n34006), .B(n34007), .Z(n34005) );
  NANDN U42977 ( .A(n34007), .B(n34006), .Z(n34002) );
  IV U42978 ( .A(n34008), .Z(n34007) );
  NAND U42979 ( .A(n34009), .B(n34010), .Z(n33979) );
  NANDN U42980 ( .A(n34011), .B(n34012), .Z(n34010) );
  NANDN U42981 ( .A(n34013), .B(n34014), .Z(n34012) );
  NANDN U42982 ( .A(n34014), .B(n34013), .Z(n34009) );
  IV U42983 ( .A(n34015), .Z(n34013) );
  AND U42984 ( .A(n34016), .B(n34017), .Z(n33982) );
  NAND U42985 ( .A(n34018), .B(n34019), .Z(n34017) );
  NANDN U42986 ( .A(n34020), .B(n34021), .Z(n34019) );
  NANDN U42987 ( .A(n34021), .B(n34020), .Z(n34016) );
  XOR U42988 ( .A(n33992), .B(n34022), .Z(n33984) );
  XNOR U42989 ( .A(n33989), .B(n33991), .Z(n34022) );
  AND U42990 ( .A(n34023), .B(n34024), .Z(n33991) );
  NANDN U42991 ( .A(n34025), .B(n34026), .Z(n34024) );
  OR U42992 ( .A(n34027), .B(n34028), .Z(n34026) );
  IV U42993 ( .A(n34029), .Z(n34028) );
  NANDN U42994 ( .A(n34029), .B(n34027), .Z(n34023) );
  AND U42995 ( .A(n34030), .B(n34031), .Z(n33989) );
  NAND U42996 ( .A(n34032), .B(n34033), .Z(n34031) );
  NANDN U42997 ( .A(n34034), .B(n34035), .Z(n34033) );
  NANDN U42998 ( .A(n34035), .B(n34034), .Z(n34030) );
  IV U42999 ( .A(n34036), .Z(n34035) );
  NAND U43000 ( .A(n34037), .B(n34038), .Z(n33992) );
  NANDN U43001 ( .A(n34039), .B(n34040), .Z(n34038) );
  NANDN U43002 ( .A(n34041), .B(n34042), .Z(n34040) );
  NANDN U43003 ( .A(n34042), .B(n34041), .Z(n34037) );
  IV U43004 ( .A(n34043), .Z(n34041) );
  XOR U43005 ( .A(n34018), .B(n34044), .Z(N62361) );
  XNOR U43006 ( .A(n34021), .B(n34020), .Z(n34044) );
  XNOR U43007 ( .A(n34032), .B(n34045), .Z(n34020) );
  XNOR U43008 ( .A(n34036), .B(n34034), .Z(n34045) );
  XOR U43009 ( .A(n34042), .B(n34046), .Z(n34034) );
  XNOR U43010 ( .A(n34039), .B(n34043), .Z(n34046) );
  AND U43011 ( .A(n34047), .B(n34048), .Z(n34043) );
  NAND U43012 ( .A(n34049), .B(n34050), .Z(n34048) );
  NAND U43013 ( .A(n34051), .B(n34052), .Z(n34047) );
  AND U43014 ( .A(n34053), .B(n34054), .Z(n34039) );
  NAND U43015 ( .A(n34055), .B(n34056), .Z(n34054) );
  NAND U43016 ( .A(n34057), .B(n34058), .Z(n34053) );
  NANDN U43017 ( .A(n34059), .B(n34060), .Z(n34042) );
  ANDN U43018 ( .B(n34061), .A(n34062), .Z(n34036) );
  XNOR U43019 ( .A(n34027), .B(n34063), .Z(n34032) );
  XNOR U43020 ( .A(n34025), .B(n34029), .Z(n34063) );
  AND U43021 ( .A(n34064), .B(n34065), .Z(n34029) );
  NAND U43022 ( .A(n34066), .B(n34067), .Z(n34065) );
  NAND U43023 ( .A(n34068), .B(n34069), .Z(n34064) );
  AND U43024 ( .A(n34070), .B(n34071), .Z(n34025) );
  NAND U43025 ( .A(n34072), .B(n34073), .Z(n34071) );
  NAND U43026 ( .A(n34074), .B(n34075), .Z(n34070) );
  AND U43027 ( .A(n34076), .B(n34077), .Z(n34027) );
  NAND U43028 ( .A(n34078), .B(n34079), .Z(n34021) );
  XNOR U43029 ( .A(n34004), .B(n34080), .Z(n34018) );
  XNOR U43030 ( .A(n34008), .B(n34006), .Z(n34080) );
  XOR U43031 ( .A(n34014), .B(n34081), .Z(n34006) );
  XNOR U43032 ( .A(n34011), .B(n34015), .Z(n34081) );
  AND U43033 ( .A(n34082), .B(n34083), .Z(n34015) );
  NAND U43034 ( .A(n34084), .B(n34085), .Z(n34083) );
  NAND U43035 ( .A(n34086), .B(n34087), .Z(n34082) );
  AND U43036 ( .A(n34088), .B(n34089), .Z(n34011) );
  NAND U43037 ( .A(n34090), .B(n34091), .Z(n34089) );
  NAND U43038 ( .A(n34092), .B(n34093), .Z(n34088) );
  NANDN U43039 ( .A(n34094), .B(n34095), .Z(n34014) );
  ANDN U43040 ( .B(n34096), .A(n34097), .Z(n34008) );
  XNOR U43041 ( .A(n33999), .B(n34098), .Z(n34004) );
  XNOR U43042 ( .A(n33997), .B(n34001), .Z(n34098) );
  AND U43043 ( .A(n34099), .B(n34100), .Z(n34001) );
  NAND U43044 ( .A(n34101), .B(n34102), .Z(n34100) );
  NAND U43045 ( .A(n34103), .B(n34104), .Z(n34099) );
  AND U43046 ( .A(n34105), .B(n34106), .Z(n33997) );
  NAND U43047 ( .A(n34107), .B(n34108), .Z(n34106) );
  NAND U43048 ( .A(n34109), .B(n34110), .Z(n34105) );
  AND U43049 ( .A(n34111), .B(n34112), .Z(n33999) );
  XOR U43050 ( .A(n34079), .B(n34078), .Z(N62360) );
  XNOR U43051 ( .A(n34096), .B(n34097), .Z(n34078) );
  XNOR U43052 ( .A(n34111), .B(n34112), .Z(n34097) );
  XOR U43053 ( .A(n34108), .B(n34107), .Z(n34112) );
  XOR U43054 ( .A(y[3276]), .B(x[3276]), .Z(n34107) );
  XOR U43055 ( .A(n34110), .B(n34109), .Z(n34108) );
  XOR U43056 ( .A(y[3278]), .B(x[3278]), .Z(n34109) );
  XOR U43057 ( .A(y[3277]), .B(x[3277]), .Z(n34110) );
  XOR U43058 ( .A(n34102), .B(n34101), .Z(n34111) );
  XOR U43059 ( .A(n34104), .B(n34103), .Z(n34101) );
  XOR U43060 ( .A(y[3275]), .B(x[3275]), .Z(n34103) );
  XOR U43061 ( .A(y[3274]), .B(x[3274]), .Z(n34104) );
  XOR U43062 ( .A(y[3273]), .B(x[3273]), .Z(n34102) );
  XNOR U43063 ( .A(n34095), .B(n34094), .Z(n34096) );
  XNOR U43064 ( .A(n34091), .B(n34090), .Z(n34094) );
  XOR U43065 ( .A(n34093), .B(n34092), .Z(n34090) );
  XOR U43066 ( .A(y[3272]), .B(x[3272]), .Z(n34092) );
  XOR U43067 ( .A(y[3271]), .B(x[3271]), .Z(n34093) );
  XOR U43068 ( .A(y[3270]), .B(x[3270]), .Z(n34091) );
  XOR U43069 ( .A(n34085), .B(n34084), .Z(n34095) );
  XOR U43070 ( .A(n34087), .B(n34086), .Z(n34084) );
  XOR U43071 ( .A(y[3269]), .B(x[3269]), .Z(n34086) );
  XOR U43072 ( .A(y[3268]), .B(x[3268]), .Z(n34087) );
  XOR U43073 ( .A(y[3267]), .B(x[3267]), .Z(n34085) );
  XNOR U43074 ( .A(n34061), .B(n34062), .Z(n34079) );
  XNOR U43075 ( .A(n34076), .B(n34077), .Z(n34062) );
  XOR U43076 ( .A(n34073), .B(n34072), .Z(n34077) );
  XOR U43077 ( .A(y[3264]), .B(x[3264]), .Z(n34072) );
  XOR U43078 ( .A(n34075), .B(n34074), .Z(n34073) );
  XOR U43079 ( .A(y[3266]), .B(x[3266]), .Z(n34074) );
  XOR U43080 ( .A(y[3265]), .B(x[3265]), .Z(n34075) );
  XOR U43081 ( .A(n34067), .B(n34066), .Z(n34076) );
  XOR U43082 ( .A(n34069), .B(n34068), .Z(n34066) );
  XOR U43083 ( .A(y[3263]), .B(x[3263]), .Z(n34068) );
  XOR U43084 ( .A(y[3262]), .B(x[3262]), .Z(n34069) );
  XOR U43085 ( .A(y[3261]), .B(x[3261]), .Z(n34067) );
  XNOR U43086 ( .A(n34060), .B(n34059), .Z(n34061) );
  XNOR U43087 ( .A(n34056), .B(n34055), .Z(n34059) );
  XOR U43088 ( .A(n34058), .B(n34057), .Z(n34055) );
  XOR U43089 ( .A(y[3260]), .B(x[3260]), .Z(n34057) );
  XOR U43090 ( .A(y[3259]), .B(x[3259]), .Z(n34058) );
  XOR U43091 ( .A(y[3258]), .B(x[3258]), .Z(n34056) );
  XOR U43092 ( .A(n34050), .B(n34049), .Z(n34060) );
  XOR U43093 ( .A(n34052), .B(n34051), .Z(n34049) );
  XOR U43094 ( .A(y[3257]), .B(x[3257]), .Z(n34051) );
  XOR U43095 ( .A(y[3256]), .B(x[3256]), .Z(n34052) );
  XOR U43096 ( .A(y[3255]), .B(x[3255]), .Z(n34050) );
  NAND U43097 ( .A(n34113), .B(n34114), .Z(N62351) );
  NAND U43098 ( .A(n34115), .B(n34116), .Z(n34114) );
  NANDN U43099 ( .A(n34117), .B(n34118), .Z(n34116) );
  NANDN U43100 ( .A(n34118), .B(n34117), .Z(n34113) );
  XOR U43101 ( .A(n34117), .B(n34119), .Z(N62350) );
  XNOR U43102 ( .A(n34115), .B(n34118), .Z(n34119) );
  NAND U43103 ( .A(n34120), .B(n34121), .Z(n34118) );
  NAND U43104 ( .A(n34122), .B(n34123), .Z(n34121) );
  NANDN U43105 ( .A(n34124), .B(n34125), .Z(n34123) );
  NANDN U43106 ( .A(n34125), .B(n34124), .Z(n34120) );
  AND U43107 ( .A(n34126), .B(n34127), .Z(n34115) );
  NAND U43108 ( .A(n34128), .B(n34129), .Z(n34127) );
  NANDN U43109 ( .A(n34130), .B(n34131), .Z(n34129) );
  NANDN U43110 ( .A(n34131), .B(n34130), .Z(n34126) );
  IV U43111 ( .A(n34132), .Z(n34131) );
  AND U43112 ( .A(n34133), .B(n34134), .Z(n34117) );
  NAND U43113 ( .A(n34135), .B(n34136), .Z(n34134) );
  NANDN U43114 ( .A(n34137), .B(n34138), .Z(n34136) );
  NANDN U43115 ( .A(n34138), .B(n34137), .Z(n34133) );
  XOR U43116 ( .A(n34130), .B(n34139), .Z(N62349) );
  XNOR U43117 ( .A(n34128), .B(n34132), .Z(n34139) );
  XOR U43118 ( .A(n34125), .B(n34140), .Z(n34132) );
  XNOR U43119 ( .A(n34122), .B(n34124), .Z(n34140) );
  AND U43120 ( .A(n34141), .B(n34142), .Z(n34124) );
  NANDN U43121 ( .A(n34143), .B(n34144), .Z(n34142) );
  OR U43122 ( .A(n34145), .B(n34146), .Z(n34144) );
  IV U43123 ( .A(n34147), .Z(n34146) );
  NANDN U43124 ( .A(n34147), .B(n34145), .Z(n34141) );
  AND U43125 ( .A(n34148), .B(n34149), .Z(n34122) );
  NAND U43126 ( .A(n34150), .B(n34151), .Z(n34149) );
  NANDN U43127 ( .A(n34152), .B(n34153), .Z(n34151) );
  NANDN U43128 ( .A(n34153), .B(n34152), .Z(n34148) );
  IV U43129 ( .A(n34154), .Z(n34153) );
  NAND U43130 ( .A(n34155), .B(n34156), .Z(n34125) );
  NANDN U43131 ( .A(n34157), .B(n34158), .Z(n34156) );
  NANDN U43132 ( .A(n34159), .B(n34160), .Z(n34158) );
  NANDN U43133 ( .A(n34160), .B(n34159), .Z(n34155) );
  IV U43134 ( .A(n34161), .Z(n34159) );
  AND U43135 ( .A(n34162), .B(n34163), .Z(n34128) );
  NAND U43136 ( .A(n34164), .B(n34165), .Z(n34163) );
  NANDN U43137 ( .A(n34166), .B(n34167), .Z(n34165) );
  NANDN U43138 ( .A(n34167), .B(n34166), .Z(n34162) );
  XOR U43139 ( .A(n34138), .B(n34168), .Z(n34130) );
  XNOR U43140 ( .A(n34135), .B(n34137), .Z(n34168) );
  AND U43141 ( .A(n34169), .B(n34170), .Z(n34137) );
  NANDN U43142 ( .A(n34171), .B(n34172), .Z(n34170) );
  OR U43143 ( .A(n34173), .B(n34174), .Z(n34172) );
  IV U43144 ( .A(n34175), .Z(n34174) );
  NANDN U43145 ( .A(n34175), .B(n34173), .Z(n34169) );
  AND U43146 ( .A(n34176), .B(n34177), .Z(n34135) );
  NAND U43147 ( .A(n34178), .B(n34179), .Z(n34177) );
  NANDN U43148 ( .A(n34180), .B(n34181), .Z(n34179) );
  NANDN U43149 ( .A(n34181), .B(n34180), .Z(n34176) );
  IV U43150 ( .A(n34182), .Z(n34181) );
  NAND U43151 ( .A(n34183), .B(n34184), .Z(n34138) );
  NANDN U43152 ( .A(n34185), .B(n34186), .Z(n34184) );
  NANDN U43153 ( .A(n34187), .B(n34188), .Z(n34186) );
  NANDN U43154 ( .A(n34188), .B(n34187), .Z(n34183) );
  IV U43155 ( .A(n34189), .Z(n34187) );
  XOR U43156 ( .A(n34164), .B(n34190), .Z(N62348) );
  XNOR U43157 ( .A(n34167), .B(n34166), .Z(n34190) );
  XNOR U43158 ( .A(n34178), .B(n34191), .Z(n34166) );
  XNOR U43159 ( .A(n34182), .B(n34180), .Z(n34191) );
  XOR U43160 ( .A(n34188), .B(n34192), .Z(n34180) );
  XNOR U43161 ( .A(n34185), .B(n34189), .Z(n34192) );
  AND U43162 ( .A(n34193), .B(n34194), .Z(n34189) );
  NAND U43163 ( .A(n34195), .B(n34196), .Z(n34194) );
  NAND U43164 ( .A(n34197), .B(n34198), .Z(n34193) );
  AND U43165 ( .A(n34199), .B(n34200), .Z(n34185) );
  NAND U43166 ( .A(n34201), .B(n34202), .Z(n34200) );
  NAND U43167 ( .A(n34203), .B(n34204), .Z(n34199) );
  NANDN U43168 ( .A(n34205), .B(n34206), .Z(n34188) );
  ANDN U43169 ( .B(n34207), .A(n34208), .Z(n34182) );
  XNOR U43170 ( .A(n34173), .B(n34209), .Z(n34178) );
  XNOR U43171 ( .A(n34171), .B(n34175), .Z(n34209) );
  AND U43172 ( .A(n34210), .B(n34211), .Z(n34175) );
  NAND U43173 ( .A(n34212), .B(n34213), .Z(n34211) );
  NAND U43174 ( .A(n34214), .B(n34215), .Z(n34210) );
  AND U43175 ( .A(n34216), .B(n34217), .Z(n34171) );
  NAND U43176 ( .A(n34218), .B(n34219), .Z(n34217) );
  NAND U43177 ( .A(n34220), .B(n34221), .Z(n34216) );
  AND U43178 ( .A(n34222), .B(n34223), .Z(n34173) );
  NAND U43179 ( .A(n34224), .B(n34225), .Z(n34167) );
  XNOR U43180 ( .A(n34150), .B(n34226), .Z(n34164) );
  XNOR U43181 ( .A(n34154), .B(n34152), .Z(n34226) );
  XOR U43182 ( .A(n34160), .B(n34227), .Z(n34152) );
  XNOR U43183 ( .A(n34157), .B(n34161), .Z(n34227) );
  AND U43184 ( .A(n34228), .B(n34229), .Z(n34161) );
  NAND U43185 ( .A(n34230), .B(n34231), .Z(n34229) );
  NAND U43186 ( .A(n34232), .B(n34233), .Z(n34228) );
  AND U43187 ( .A(n34234), .B(n34235), .Z(n34157) );
  NAND U43188 ( .A(n34236), .B(n34237), .Z(n34235) );
  NAND U43189 ( .A(n34238), .B(n34239), .Z(n34234) );
  NANDN U43190 ( .A(n34240), .B(n34241), .Z(n34160) );
  ANDN U43191 ( .B(n34242), .A(n34243), .Z(n34154) );
  XNOR U43192 ( .A(n34145), .B(n34244), .Z(n34150) );
  XNOR U43193 ( .A(n34143), .B(n34147), .Z(n34244) );
  AND U43194 ( .A(n34245), .B(n34246), .Z(n34147) );
  NAND U43195 ( .A(n34247), .B(n34248), .Z(n34246) );
  NAND U43196 ( .A(n34249), .B(n34250), .Z(n34245) );
  AND U43197 ( .A(n34251), .B(n34252), .Z(n34143) );
  NAND U43198 ( .A(n34253), .B(n34254), .Z(n34252) );
  NAND U43199 ( .A(n34255), .B(n34256), .Z(n34251) );
  AND U43200 ( .A(n34257), .B(n34258), .Z(n34145) );
  XOR U43201 ( .A(n34225), .B(n34224), .Z(N62347) );
  XNOR U43202 ( .A(n34242), .B(n34243), .Z(n34224) );
  XNOR U43203 ( .A(n34257), .B(n34258), .Z(n34243) );
  XOR U43204 ( .A(n34254), .B(n34253), .Z(n34258) );
  XOR U43205 ( .A(y[3252]), .B(x[3252]), .Z(n34253) );
  XOR U43206 ( .A(n34256), .B(n34255), .Z(n34254) );
  XOR U43207 ( .A(y[3254]), .B(x[3254]), .Z(n34255) );
  XOR U43208 ( .A(y[3253]), .B(x[3253]), .Z(n34256) );
  XOR U43209 ( .A(n34248), .B(n34247), .Z(n34257) );
  XOR U43210 ( .A(n34250), .B(n34249), .Z(n34247) );
  XOR U43211 ( .A(y[3251]), .B(x[3251]), .Z(n34249) );
  XOR U43212 ( .A(y[3250]), .B(x[3250]), .Z(n34250) );
  XOR U43213 ( .A(y[3249]), .B(x[3249]), .Z(n34248) );
  XNOR U43214 ( .A(n34241), .B(n34240), .Z(n34242) );
  XNOR U43215 ( .A(n34237), .B(n34236), .Z(n34240) );
  XOR U43216 ( .A(n34239), .B(n34238), .Z(n34236) );
  XOR U43217 ( .A(y[3248]), .B(x[3248]), .Z(n34238) );
  XOR U43218 ( .A(y[3247]), .B(x[3247]), .Z(n34239) );
  XOR U43219 ( .A(y[3246]), .B(x[3246]), .Z(n34237) );
  XOR U43220 ( .A(n34231), .B(n34230), .Z(n34241) );
  XOR U43221 ( .A(n34233), .B(n34232), .Z(n34230) );
  XOR U43222 ( .A(y[3245]), .B(x[3245]), .Z(n34232) );
  XOR U43223 ( .A(y[3244]), .B(x[3244]), .Z(n34233) );
  XOR U43224 ( .A(y[3243]), .B(x[3243]), .Z(n34231) );
  XNOR U43225 ( .A(n34207), .B(n34208), .Z(n34225) );
  XNOR U43226 ( .A(n34222), .B(n34223), .Z(n34208) );
  XOR U43227 ( .A(n34219), .B(n34218), .Z(n34223) );
  XOR U43228 ( .A(y[3240]), .B(x[3240]), .Z(n34218) );
  XOR U43229 ( .A(n34221), .B(n34220), .Z(n34219) );
  XOR U43230 ( .A(y[3242]), .B(x[3242]), .Z(n34220) );
  XOR U43231 ( .A(y[3241]), .B(x[3241]), .Z(n34221) );
  XOR U43232 ( .A(n34213), .B(n34212), .Z(n34222) );
  XOR U43233 ( .A(n34215), .B(n34214), .Z(n34212) );
  XOR U43234 ( .A(y[3239]), .B(x[3239]), .Z(n34214) );
  XOR U43235 ( .A(y[3238]), .B(x[3238]), .Z(n34215) );
  XOR U43236 ( .A(y[3237]), .B(x[3237]), .Z(n34213) );
  XNOR U43237 ( .A(n34206), .B(n34205), .Z(n34207) );
  XNOR U43238 ( .A(n34202), .B(n34201), .Z(n34205) );
  XOR U43239 ( .A(n34204), .B(n34203), .Z(n34201) );
  XOR U43240 ( .A(y[3236]), .B(x[3236]), .Z(n34203) );
  XOR U43241 ( .A(y[3235]), .B(x[3235]), .Z(n34204) );
  XOR U43242 ( .A(y[3234]), .B(x[3234]), .Z(n34202) );
  XOR U43243 ( .A(n34196), .B(n34195), .Z(n34206) );
  XOR U43244 ( .A(n34198), .B(n34197), .Z(n34195) );
  XOR U43245 ( .A(y[3233]), .B(x[3233]), .Z(n34197) );
  XOR U43246 ( .A(y[3232]), .B(x[3232]), .Z(n34198) );
  XOR U43247 ( .A(y[3231]), .B(x[3231]), .Z(n34196) );
  NAND U43248 ( .A(n34259), .B(n34260), .Z(N62338) );
  NAND U43249 ( .A(n34261), .B(n34262), .Z(n34260) );
  NANDN U43250 ( .A(n34263), .B(n34264), .Z(n34262) );
  NANDN U43251 ( .A(n34264), .B(n34263), .Z(n34259) );
  XOR U43252 ( .A(n34263), .B(n34265), .Z(N62337) );
  XNOR U43253 ( .A(n34261), .B(n34264), .Z(n34265) );
  NAND U43254 ( .A(n34266), .B(n34267), .Z(n34264) );
  NAND U43255 ( .A(n34268), .B(n34269), .Z(n34267) );
  NANDN U43256 ( .A(n34270), .B(n34271), .Z(n34269) );
  NANDN U43257 ( .A(n34271), .B(n34270), .Z(n34266) );
  AND U43258 ( .A(n34272), .B(n34273), .Z(n34261) );
  NAND U43259 ( .A(n34274), .B(n34275), .Z(n34273) );
  NANDN U43260 ( .A(n34276), .B(n34277), .Z(n34275) );
  NANDN U43261 ( .A(n34277), .B(n34276), .Z(n34272) );
  IV U43262 ( .A(n34278), .Z(n34277) );
  AND U43263 ( .A(n34279), .B(n34280), .Z(n34263) );
  NAND U43264 ( .A(n34281), .B(n34282), .Z(n34280) );
  NANDN U43265 ( .A(n34283), .B(n34284), .Z(n34282) );
  NANDN U43266 ( .A(n34284), .B(n34283), .Z(n34279) );
  XOR U43267 ( .A(n34276), .B(n34285), .Z(N62336) );
  XNOR U43268 ( .A(n34274), .B(n34278), .Z(n34285) );
  XOR U43269 ( .A(n34271), .B(n34286), .Z(n34278) );
  XNOR U43270 ( .A(n34268), .B(n34270), .Z(n34286) );
  AND U43271 ( .A(n34287), .B(n34288), .Z(n34270) );
  NANDN U43272 ( .A(n34289), .B(n34290), .Z(n34288) );
  OR U43273 ( .A(n34291), .B(n34292), .Z(n34290) );
  IV U43274 ( .A(n34293), .Z(n34292) );
  NANDN U43275 ( .A(n34293), .B(n34291), .Z(n34287) );
  AND U43276 ( .A(n34294), .B(n34295), .Z(n34268) );
  NAND U43277 ( .A(n34296), .B(n34297), .Z(n34295) );
  NANDN U43278 ( .A(n34298), .B(n34299), .Z(n34297) );
  NANDN U43279 ( .A(n34299), .B(n34298), .Z(n34294) );
  IV U43280 ( .A(n34300), .Z(n34299) );
  NAND U43281 ( .A(n34301), .B(n34302), .Z(n34271) );
  NANDN U43282 ( .A(n34303), .B(n34304), .Z(n34302) );
  NANDN U43283 ( .A(n34305), .B(n34306), .Z(n34304) );
  NANDN U43284 ( .A(n34306), .B(n34305), .Z(n34301) );
  IV U43285 ( .A(n34307), .Z(n34305) );
  AND U43286 ( .A(n34308), .B(n34309), .Z(n34274) );
  NAND U43287 ( .A(n34310), .B(n34311), .Z(n34309) );
  NANDN U43288 ( .A(n34312), .B(n34313), .Z(n34311) );
  NANDN U43289 ( .A(n34313), .B(n34312), .Z(n34308) );
  XOR U43290 ( .A(n34284), .B(n34314), .Z(n34276) );
  XNOR U43291 ( .A(n34281), .B(n34283), .Z(n34314) );
  AND U43292 ( .A(n34315), .B(n34316), .Z(n34283) );
  NANDN U43293 ( .A(n34317), .B(n34318), .Z(n34316) );
  OR U43294 ( .A(n34319), .B(n34320), .Z(n34318) );
  IV U43295 ( .A(n34321), .Z(n34320) );
  NANDN U43296 ( .A(n34321), .B(n34319), .Z(n34315) );
  AND U43297 ( .A(n34322), .B(n34323), .Z(n34281) );
  NAND U43298 ( .A(n34324), .B(n34325), .Z(n34323) );
  NANDN U43299 ( .A(n34326), .B(n34327), .Z(n34325) );
  NANDN U43300 ( .A(n34327), .B(n34326), .Z(n34322) );
  IV U43301 ( .A(n34328), .Z(n34327) );
  NAND U43302 ( .A(n34329), .B(n34330), .Z(n34284) );
  NANDN U43303 ( .A(n34331), .B(n34332), .Z(n34330) );
  NANDN U43304 ( .A(n34333), .B(n34334), .Z(n34332) );
  NANDN U43305 ( .A(n34334), .B(n34333), .Z(n34329) );
  IV U43306 ( .A(n34335), .Z(n34333) );
  XOR U43307 ( .A(n34310), .B(n34336), .Z(N62335) );
  XNOR U43308 ( .A(n34313), .B(n34312), .Z(n34336) );
  XNOR U43309 ( .A(n34324), .B(n34337), .Z(n34312) );
  XNOR U43310 ( .A(n34328), .B(n34326), .Z(n34337) );
  XOR U43311 ( .A(n34334), .B(n34338), .Z(n34326) );
  XNOR U43312 ( .A(n34331), .B(n34335), .Z(n34338) );
  AND U43313 ( .A(n34339), .B(n34340), .Z(n34335) );
  NAND U43314 ( .A(n34341), .B(n34342), .Z(n34340) );
  NAND U43315 ( .A(n34343), .B(n34344), .Z(n34339) );
  AND U43316 ( .A(n34345), .B(n34346), .Z(n34331) );
  NAND U43317 ( .A(n34347), .B(n34348), .Z(n34346) );
  NAND U43318 ( .A(n34349), .B(n34350), .Z(n34345) );
  NANDN U43319 ( .A(n34351), .B(n34352), .Z(n34334) );
  ANDN U43320 ( .B(n34353), .A(n34354), .Z(n34328) );
  XNOR U43321 ( .A(n34319), .B(n34355), .Z(n34324) );
  XNOR U43322 ( .A(n34317), .B(n34321), .Z(n34355) );
  AND U43323 ( .A(n34356), .B(n34357), .Z(n34321) );
  NAND U43324 ( .A(n34358), .B(n34359), .Z(n34357) );
  NAND U43325 ( .A(n34360), .B(n34361), .Z(n34356) );
  AND U43326 ( .A(n34362), .B(n34363), .Z(n34317) );
  NAND U43327 ( .A(n34364), .B(n34365), .Z(n34363) );
  NAND U43328 ( .A(n34366), .B(n34367), .Z(n34362) );
  AND U43329 ( .A(n34368), .B(n34369), .Z(n34319) );
  NAND U43330 ( .A(n34370), .B(n34371), .Z(n34313) );
  XNOR U43331 ( .A(n34296), .B(n34372), .Z(n34310) );
  XNOR U43332 ( .A(n34300), .B(n34298), .Z(n34372) );
  XOR U43333 ( .A(n34306), .B(n34373), .Z(n34298) );
  XNOR U43334 ( .A(n34303), .B(n34307), .Z(n34373) );
  AND U43335 ( .A(n34374), .B(n34375), .Z(n34307) );
  NAND U43336 ( .A(n34376), .B(n34377), .Z(n34375) );
  NAND U43337 ( .A(n34378), .B(n34379), .Z(n34374) );
  AND U43338 ( .A(n34380), .B(n34381), .Z(n34303) );
  NAND U43339 ( .A(n34382), .B(n34383), .Z(n34381) );
  NAND U43340 ( .A(n34384), .B(n34385), .Z(n34380) );
  NANDN U43341 ( .A(n34386), .B(n34387), .Z(n34306) );
  ANDN U43342 ( .B(n34388), .A(n34389), .Z(n34300) );
  XNOR U43343 ( .A(n34291), .B(n34390), .Z(n34296) );
  XNOR U43344 ( .A(n34289), .B(n34293), .Z(n34390) );
  AND U43345 ( .A(n34391), .B(n34392), .Z(n34293) );
  NAND U43346 ( .A(n34393), .B(n34394), .Z(n34392) );
  NAND U43347 ( .A(n34395), .B(n34396), .Z(n34391) );
  AND U43348 ( .A(n34397), .B(n34398), .Z(n34289) );
  NAND U43349 ( .A(n34399), .B(n34400), .Z(n34398) );
  NAND U43350 ( .A(n34401), .B(n34402), .Z(n34397) );
  AND U43351 ( .A(n34403), .B(n34404), .Z(n34291) );
  XOR U43352 ( .A(n34371), .B(n34370), .Z(N62334) );
  XNOR U43353 ( .A(n34388), .B(n34389), .Z(n34370) );
  XNOR U43354 ( .A(n34403), .B(n34404), .Z(n34389) );
  XOR U43355 ( .A(n34400), .B(n34399), .Z(n34404) );
  XOR U43356 ( .A(y[3228]), .B(x[3228]), .Z(n34399) );
  XOR U43357 ( .A(n34402), .B(n34401), .Z(n34400) );
  XOR U43358 ( .A(y[3230]), .B(x[3230]), .Z(n34401) );
  XOR U43359 ( .A(y[3229]), .B(x[3229]), .Z(n34402) );
  XOR U43360 ( .A(n34394), .B(n34393), .Z(n34403) );
  XOR U43361 ( .A(n34396), .B(n34395), .Z(n34393) );
  XOR U43362 ( .A(y[3227]), .B(x[3227]), .Z(n34395) );
  XOR U43363 ( .A(y[3226]), .B(x[3226]), .Z(n34396) );
  XOR U43364 ( .A(y[3225]), .B(x[3225]), .Z(n34394) );
  XNOR U43365 ( .A(n34387), .B(n34386), .Z(n34388) );
  XNOR U43366 ( .A(n34383), .B(n34382), .Z(n34386) );
  XOR U43367 ( .A(n34385), .B(n34384), .Z(n34382) );
  XOR U43368 ( .A(y[3224]), .B(x[3224]), .Z(n34384) );
  XOR U43369 ( .A(y[3223]), .B(x[3223]), .Z(n34385) );
  XOR U43370 ( .A(y[3222]), .B(x[3222]), .Z(n34383) );
  XOR U43371 ( .A(n34377), .B(n34376), .Z(n34387) );
  XOR U43372 ( .A(n34379), .B(n34378), .Z(n34376) );
  XOR U43373 ( .A(y[3221]), .B(x[3221]), .Z(n34378) );
  XOR U43374 ( .A(y[3220]), .B(x[3220]), .Z(n34379) );
  XOR U43375 ( .A(y[3219]), .B(x[3219]), .Z(n34377) );
  XNOR U43376 ( .A(n34353), .B(n34354), .Z(n34371) );
  XNOR U43377 ( .A(n34368), .B(n34369), .Z(n34354) );
  XOR U43378 ( .A(n34365), .B(n34364), .Z(n34369) );
  XOR U43379 ( .A(y[3216]), .B(x[3216]), .Z(n34364) );
  XOR U43380 ( .A(n34367), .B(n34366), .Z(n34365) );
  XOR U43381 ( .A(y[3218]), .B(x[3218]), .Z(n34366) );
  XOR U43382 ( .A(y[3217]), .B(x[3217]), .Z(n34367) );
  XOR U43383 ( .A(n34359), .B(n34358), .Z(n34368) );
  XOR U43384 ( .A(n34361), .B(n34360), .Z(n34358) );
  XOR U43385 ( .A(y[3215]), .B(x[3215]), .Z(n34360) );
  XOR U43386 ( .A(y[3214]), .B(x[3214]), .Z(n34361) );
  XOR U43387 ( .A(y[3213]), .B(x[3213]), .Z(n34359) );
  XNOR U43388 ( .A(n34352), .B(n34351), .Z(n34353) );
  XNOR U43389 ( .A(n34348), .B(n34347), .Z(n34351) );
  XOR U43390 ( .A(n34350), .B(n34349), .Z(n34347) );
  XOR U43391 ( .A(y[3212]), .B(x[3212]), .Z(n34349) );
  XOR U43392 ( .A(y[3211]), .B(x[3211]), .Z(n34350) );
  XOR U43393 ( .A(y[3210]), .B(x[3210]), .Z(n34348) );
  XOR U43394 ( .A(n34342), .B(n34341), .Z(n34352) );
  XOR U43395 ( .A(n34344), .B(n34343), .Z(n34341) );
  XOR U43396 ( .A(y[3209]), .B(x[3209]), .Z(n34343) );
  XOR U43397 ( .A(y[3208]), .B(x[3208]), .Z(n34344) );
  XOR U43398 ( .A(y[3207]), .B(x[3207]), .Z(n34342) );
  NAND U43399 ( .A(n34405), .B(n34406), .Z(N62325) );
  NAND U43400 ( .A(n34407), .B(n34408), .Z(n34406) );
  NANDN U43401 ( .A(n34409), .B(n34410), .Z(n34408) );
  NANDN U43402 ( .A(n34410), .B(n34409), .Z(n34405) );
  XOR U43403 ( .A(n34409), .B(n34411), .Z(N62324) );
  XNOR U43404 ( .A(n34407), .B(n34410), .Z(n34411) );
  NAND U43405 ( .A(n34412), .B(n34413), .Z(n34410) );
  NAND U43406 ( .A(n34414), .B(n34415), .Z(n34413) );
  NANDN U43407 ( .A(n34416), .B(n34417), .Z(n34415) );
  NANDN U43408 ( .A(n34417), .B(n34416), .Z(n34412) );
  AND U43409 ( .A(n34418), .B(n34419), .Z(n34407) );
  NAND U43410 ( .A(n34420), .B(n34421), .Z(n34419) );
  NANDN U43411 ( .A(n34422), .B(n34423), .Z(n34421) );
  NANDN U43412 ( .A(n34423), .B(n34422), .Z(n34418) );
  IV U43413 ( .A(n34424), .Z(n34423) );
  AND U43414 ( .A(n34425), .B(n34426), .Z(n34409) );
  NAND U43415 ( .A(n34427), .B(n34428), .Z(n34426) );
  NANDN U43416 ( .A(n34429), .B(n34430), .Z(n34428) );
  NANDN U43417 ( .A(n34430), .B(n34429), .Z(n34425) );
  XOR U43418 ( .A(n34422), .B(n34431), .Z(N62323) );
  XNOR U43419 ( .A(n34420), .B(n34424), .Z(n34431) );
  XOR U43420 ( .A(n34417), .B(n34432), .Z(n34424) );
  XNOR U43421 ( .A(n34414), .B(n34416), .Z(n34432) );
  AND U43422 ( .A(n34433), .B(n34434), .Z(n34416) );
  NANDN U43423 ( .A(n34435), .B(n34436), .Z(n34434) );
  OR U43424 ( .A(n34437), .B(n34438), .Z(n34436) );
  IV U43425 ( .A(n34439), .Z(n34438) );
  NANDN U43426 ( .A(n34439), .B(n34437), .Z(n34433) );
  AND U43427 ( .A(n34440), .B(n34441), .Z(n34414) );
  NAND U43428 ( .A(n34442), .B(n34443), .Z(n34441) );
  NANDN U43429 ( .A(n34444), .B(n34445), .Z(n34443) );
  NANDN U43430 ( .A(n34445), .B(n34444), .Z(n34440) );
  IV U43431 ( .A(n34446), .Z(n34445) );
  NAND U43432 ( .A(n34447), .B(n34448), .Z(n34417) );
  NANDN U43433 ( .A(n34449), .B(n34450), .Z(n34448) );
  NANDN U43434 ( .A(n34451), .B(n34452), .Z(n34450) );
  NANDN U43435 ( .A(n34452), .B(n34451), .Z(n34447) );
  IV U43436 ( .A(n34453), .Z(n34451) );
  AND U43437 ( .A(n34454), .B(n34455), .Z(n34420) );
  NAND U43438 ( .A(n34456), .B(n34457), .Z(n34455) );
  NANDN U43439 ( .A(n34458), .B(n34459), .Z(n34457) );
  NANDN U43440 ( .A(n34459), .B(n34458), .Z(n34454) );
  XOR U43441 ( .A(n34430), .B(n34460), .Z(n34422) );
  XNOR U43442 ( .A(n34427), .B(n34429), .Z(n34460) );
  AND U43443 ( .A(n34461), .B(n34462), .Z(n34429) );
  NANDN U43444 ( .A(n34463), .B(n34464), .Z(n34462) );
  OR U43445 ( .A(n34465), .B(n34466), .Z(n34464) );
  IV U43446 ( .A(n34467), .Z(n34466) );
  NANDN U43447 ( .A(n34467), .B(n34465), .Z(n34461) );
  AND U43448 ( .A(n34468), .B(n34469), .Z(n34427) );
  NAND U43449 ( .A(n34470), .B(n34471), .Z(n34469) );
  NANDN U43450 ( .A(n34472), .B(n34473), .Z(n34471) );
  NANDN U43451 ( .A(n34473), .B(n34472), .Z(n34468) );
  IV U43452 ( .A(n34474), .Z(n34473) );
  NAND U43453 ( .A(n34475), .B(n34476), .Z(n34430) );
  NANDN U43454 ( .A(n34477), .B(n34478), .Z(n34476) );
  NANDN U43455 ( .A(n34479), .B(n34480), .Z(n34478) );
  NANDN U43456 ( .A(n34480), .B(n34479), .Z(n34475) );
  IV U43457 ( .A(n34481), .Z(n34479) );
  XOR U43458 ( .A(n34456), .B(n34482), .Z(N62322) );
  XNOR U43459 ( .A(n34459), .B(n34458), .Z(n34482) );
  XNOR U43460 ( .A(n34470), .B(n34483), .Z(n34458) );
  XNOR U43461 ( .A(n34474), .B(n34472), .Z(n34483) );
  XOR U43462 ( .A(n34480), .B(n34484), .Z(n34472) );
  XNOR U43463 ( .A(n34477), .B(n34481), .Z(n34484) );
  AND U43464 ( .A(n34485), .B(n34486), .Z(n34481) );
  NAND U43465 ( .A(n34487), .B(n34488), .Z(n34486) );
  NAND U43466 ( .A(n34489), .B(n34490), .Z(n34485) );
  AND U43467 ( .A(n34491), .B(n34492), .Z(n34477) );
  NAND U43468 ( .A(n34493), .B(n34494), .Z(n34492) );
  NAND U43469 ( .A(n34495), .B(n34496), .Z(n34491) );
  NANDN U43470 ( .A(n34497), .B(n34498), .Z(n34480) );
  ANDN U43471 ( .B(n34499), .A(n34500), .Z(n34474) );
  XNOR U43472 ( .A(n34465), .B(n34501), .Z(n34470) );
  XNOR U43473 ( .A(n34463), .B(n34467), .Z(n34501) );
  AND U43474 ( .A(n34502), .B(n34503), .Z(n34467) );
  NAND U43475 ( .A(n34504), .B(n34505), .Z(n34503) );
  NAND U43476 ( .A(n34506), .B(n34507), .Z(n34502) );
  AND U43477 ( .A(n34508), .B(n34509), .Z(n34463) );
  NAND U43478 ( .A(n34510), .B(n34511), .Z(n34509) );
  NAND U43479 ( .A(n34512), .B(n34513), .Z(n34508) );
  AND U43480 ( .A(n34514), .B(n34515), .Z(n34465) );
  NAND U43481 ( .A(n34516), .B(n34517), .Z(n34459) );
  XNOR U43482 ( .A(n34442), .B(n34518), .Z(n34456) );
  XNOR U43483 ( .A(n34446), .B(n34444), .Z(n34518) );
  XOR U43484 ( .A(n34452), .B(n34519), .Z(n34444) );
  XNOR U43485 ( .A(n34449), .B(n34453), .Z(n34519) );
  AND U43486 ( .A(n34520), .B(n34521), .Z(n34453) );
  NAND U43487 ( .A(n34522), .B(n34523), .Z(n34521) );
  NAND U43488 ( .A(n34524), .B(n34525), .Z(n34520) );
  AND U43489 ( .A(n34526), .B(n34527), .Z(n34449) );
  NAND U43490 ( .A(n34528), .B(n34529), .Z(n34527) );
  NAND U43491 ( .A(n34530), .B(n34531), .Z(n34526) );
  NANDN U43492 ( .A(n34532), .B(n34533), .Z(n34452) );
  ANDN U43493 ( .B(n34534), .A(n34535), .Z(n34446) );
  XNOR U43494 ( .A(n34437), .B(n34536), .Z(n34442) );
  XNOR U43495 ( .A(n34435), .B(n34439), .Z(n34536) );
  AND U43496 ( .A(n34537), .B(n34538), .Z(n34439) );
  NAND U43497 ( .A(n34539), .B(n34540), .Z(n34538) );
  NAND U43498 ( .A(n34541), .B(n34542), .Z(n34537) );
  AND U43499 ( .A(n34543), .B(n34544), .Z(n34435) );
  NAND U43500 ( .A(n34545), .B(n34546), .Z(n34544) );
  NAND U43501 ( .A(n34547), .B(n34548), .Z(n34543) );
  AND U43502 ( .A(n34549), .B(n34550), .Z(n34437) );
  XOR U43503 ( .A(n34517), .B(n34516), .Z(N62321) );
  XNOR U43504 ( .A(n34534), .B(n34535), .Z(n34516) );
  XNOR U43505 ( .A(n34549), .B(n34550), .Z(n34535) );
  XOR U43506 ( .A(n34546), .B(n34545), .Z(n34550) );
  XOR U43507 ( .A(y[3204]), .B(x[3204]), .Z(n34545) );
  XOR U43508 ( .A(n34548), .B(n34547), .Z(n34546) );
  XOR U43509 ( .A(y[3206]), .B(x[3206]), .Z(n34547) );
  XOR U43510 ( .A(y[3205]), .B(x[3205]), .Z(n34548) );
  XOR U43511 ( .A(n34540), .B(n34539), .Z(n34549) );
  XOR U43512 ( .A(n34542), .B(n34541), .Z(n34539) );
  XOR U43513 ( .A(y[3203]), .B(x[3203]), .Z(n34541) );
  XOR U43514 ( .A(y[3202]), .B(x[3202]), .Z(n34542) );
  XOR U43515 ( .A(y[3201]), .B(x[3201]), .Z(n34540) );
  XNOR U43516 ( .A(n34533), .B(n34532), .Z(n34534) );
  XNOR U43517 ( .A(n34529), .B(n34528), .Z(n34532) );
  XOR U43518 ( .A(n34531), .B(n34530), .Z(n34528) );
  XOR U43519 ( .A(y[3200]), .B(x[3200]), .Z(n34530) );
  XOR U43520 ( .A(y[3199]), .B(x[3199]), .Z(n34531) );
  XOR U43521 ( .A(y[3198]), .B(x[3198]), .Z(n34529) );
  XOR U43522 ( .A(n34523), .B(n34522), .Z(n34533) );
  XOR U43523 ( .A(n34525), .B(n34524), .Z(n34522) );
  XOR U43524 ( .A(y[3197]), .B(x[3197]), .Z(n34524) );
  XOR U43525 ( .A(y[3196]), .B(x[3196]), .Z(n34525) );
  XOR U43526 ( .A(y[3195]), .B(x[3195]), .Z(n34523) );
  XNOR U43527 ( .A(n34499), .B(n34500), .Z(n34517) );
  XNOR U43528 ( .A(n34514), .B(n34515), .Z(n34500) );
  XOR U43529 ( .A(n34511), .B(n34510), .Z(n34515) );
  XOR U43530 ( .A(y[3192]), .B(x[3192]), .Z(n34510) );
  XOR U43531 ( .A(n34513), .B(n34512), .Z(n34511) );
  XOR U43532 ( .A(y[3194]), .B(x[3194]), .Z(n34512) );
  XOR U43533 ( .A(y[3193]), .B(x[3193]), .Z(n34513) );
  XOR U43534 ( .A(n34505), .B(n34504), .Z(n34514) );
  XOR U43535 ( .A(n34507), .B(n34506), .Z(n34504) );
  XOR U43536 ( .A(y[3191]), .B(x[3191]), .Z(n34506) );
  XOR U43537 ( .A(y[3190]), .B(x[3190]), .Z(n34507) );
  XOR U43538 ( .A(y[3189]), .B(x[3189]), .Z(n34505) );
  XNOR U43539 ( .A(n34498), .B(n34497), .Z(n34499) );
  XNOR U43540 ( .A(n34494), .B(n34493), .Z(n34497) );
  XOR U43541 ( .A(n34496), .B(n34495), .Z(n34493) );
  XOR U43542 ( .A(y[3188]), .B(x[3188]), .Z(n34495) );
  XOR U43543 ( .A(y[3187]), .B(x[3187]), .Z(n34496) );
  XOR U43544 ( .A(y[3186]), .B(x[3186]), .Z(n34494) );
  XOR U43545 ( .A(n34488), .B(n34487), .Z(n34498) );
  XOR U43546 ( .A(n34490), .B(n34489), .Z(n34487) );
  XOR U43547 ( .A(y[3185]), .B(x[3185]), .Z(n34489) );
  XOR U43548 ( .A(y[3184]), .B(x[3184]), .Z(n34490) );
  XOR U43549 ( .A(y[3183]), .B(x[3183]), .Z(n34488) );
  NAND U43550 ( .A(n34551), .B(n34552), .Z(N62312) );
  NAND U43551 ( .A(n34553), .B(n34554), .Z(n34552) );
  NANDN U43552 ( .A(n34555), .B(n34556), .Z(n34554) );
  NANDN U43553 ( .A(n34556), .B(n34555), .Z(n34551) );
  XOR U43554 ( .A(n34555), .B(n34557), .Z(N62311) );
  XNOR U43555 ( .A(n34553), .B(n34556), .Z(n34557) );
  NAND U43556 ( .A(n34558), .B(n34559), .Z(n34556) );
  NAND U43557 ( .A(n34560), .B(n34561), .Z(n34559) );
  NANDN U43558 ( .A(n34562), .B(n34563), .Z(n34561) );
  NANDN U43559 ( .A(n34563), .B(n34562), .Z(n34558) );
  AND U43560 ( .A(n34564), .B(n34565), .Z(n34553) );
  NAND U43561 ( .A(n34566), .B(n34567), .Z(n34565) );
  NANDN U43562 ( .A(n34568), .B(n34569), .Z(n34567) );
  NANDN U43563 ( .A(n34569), .B(n34568), .Z(n34564) );
  IV U43564 ( .A(n34570), .Z(n34569) );
  AND U43565 ( .A(n34571), .B(n34572), .Z(n34555) );
  NAND U43566 ( .A(n34573), .B(n34574), .Z(n34572) );
  NANDN U43567 ( .A(n34575), .B(n34576), .Z(n34574) );
  NANDN U43568 ( .A(n34576), .B(n34575), .Z(n34571) );
  XOR U43569 ( .A(n34568), .B(n34577), .Z(N62310) );
  XNOR U43570 ( .A(n34566), .B(n34570), .Z(n34577) );
  XOR U43571 ( .A(n34563), .B(n34578), .Z(n34570) );
  XNOR U43572 ( .A(n34560), .B(n34562), .Z(n34578) );
  AND U43573 ( .A(n34579), .B(n34580), .Z(n34562) );
  NANDN U43574 ( .A(n34581), .B(n34582), .Z(n34580) );
  OR U43575 ( .A(n34583), .B(n34584), .Z(n34582) );
  IV U43576 ( .A(n34585), .Z(n34584) );
  NANDN U43577 ( .A(n34585), .B(n34583), .Z(n34579) );
  AND U43578 ( .A(n34586), .B(n34587), .Z(n34560) );
  NAND U43579 ( .A(n34588), .B(n34589), .Z(n34587) );
  NANDN U43580 ( .A(n34590), .B(n34591), .Z(n34589) );
  NANDN U43581 ( .A(n34591), .B(n34590), .Z(n34586) );
  IV U43582 ( .A(n34592), .Z(n34591) );
  NAND U43583 ( .A(n34593), .B(n34594), .Z(n34563) );
  NANDN U43584 ( .A(n34595), .B(n34596), .Z(n34594) );
  NANDN U43585 ( .A(n34597), .B(n34598), .Z(n34596) );
  NANDN U43586 ( .A(n34598), .B(n34597), .Z(n34593) );
  IV U43587 ( .A(n34599), .Z(n34597) );
  AND U43588 ( .A(n34600), .B(n34601), .Z(n34566) );
  NAND U43589 ( .A(n34602), .B(n34603), .Z(n34601) );
  NANDN U43590 ( .A(n34604), .B(n34605), .Z(n34603) );
  NANDN U43591 ( .A(n34605), .B(n34604), .Z(n34600) );
  XOR U43592 ( .A(n34576), .B(n34606), .Z(n34568) );
  XNOR U43593 ( .A(n34573), .B(n34575), .Z(n34606) );
  AND U43594 ( .A(n34607), .B(n34608), .Z(n34575) );
  NANDN U43595 ( .A(n34609), .B(n34610), .Z(n34608) );
  OR U43596 ( .A(n34611), .B(n34612), .Z(n34610) );
  IV U43597 ( .A(n34613), .Z(n34612) );
  NANDN U43598 ( .A(n34613), .B(n34611), .Z(n34607) );
  AND U43599 ( .A(n34614), .B(n34615), .Z(n34573) );
  NAND U43600 ( .A(n34616), .B(n34617), .Z(n34615) );
  NANDN U43601 ( .A(n34618), .B(n34619), .Z(n34617) );
  NANDN U43602 ( .A(n34619), .B(n34618), .Z(n34614) );
  IV U43603 ( .A(n34620), .Z(n34619) );
  NAND U43604 ( .A(n34621), .B(n34622), .Z(n34576) );
  NANDN U43605 ( .A(n34623), .B(n34624), .Z(n34622) );
  NANDN U43606 ( .A(n34625), .B(n34626), .Z(n34624) );
  NANDN U43607 ( .A(n34626), .B(n34625), .Z(n34621) );
  IV U43608 ( .A(n34627), .Z(n34625) );
  XOR U43609 ( .A(n34602), .B(n34628), .Z(N62309) );
  XNOR U43610 ( .A(n34605), .B(n34604), .Z(n34628) );
  XNOR U43611 ( .A(n34616), .B(n34629), .Z(n34604) );
  XNOR U43612 ( .A(n34620), .B(n34618), .Z(n34629) );
  XOR U43613 ( .A(n34626), .B(n34630), .Z(n34618) );
  XNOR U43614 ( .A(n34623), .B(n34627), .Z(n34630) );
  AND U43615 ( .A(n34631), .B(n34632), .Z(n34627) );
  NAND U43616 ( .A(n34633), .B(n34634), .Z(n34632) );
  NAND U43617 ( .A(n34635), .B(n34636), .Z(n34631) );
  AND U43618 ( .A(n34637), .B(n34638), .Z(n34623) );
  NAND U43619 ( .A(n34639), .B(n34640), .Z(n34638) );
  NAND U43620 ( .A(n34641), .B(n34642), .Z(n34637) );
  NANDN U43621 ( .A(n34643), .B(n34644), .Z(n34626) );
  ANDN U43622 ( .B(n34645), .A(n34646), .Z(n34620) );
  XNOR U43623 ( .A(n34611), .B(n34647), .Z(n34616) );
  XNOR U43624 ( .A(n34609), .B(n34613), .Z(n34647) );
  AND U43625 ( .A(n34648), .B(n34649), .Z(n34613) );
  NAND U43626 ( .A(n34650), .B(n34651), .Z(n34649) );
  NAND U43627 ( .A(n34652), .B(n34653), .Z(n34648) );
  AND U43628 ( .A(n34654), .B(n34655), .Z(n34609) );
  NAND U43629 ( .A(n34656), .B(n34657), .Z(n34655) );
  NAND U43630 ( .A(n34658), .B(n34659), .Z(n34654) );
  AND U43631 ( .A(n34660), .B(n34661), .Z(n34611) );
  NAND U43632 ( .A(n34662), .B(n34663), .Z(n34605) );
  XNOR U43633 ( .A(n34588), .B(n34664), .Z(n34602) );
  XNOR U43634 ( .A(n34592), .B(n34590), .Z(n34664) );
  XOR U43635 ( .A(n34598), .B(n34665), .Z(n34590) );
  XNOR U43636 ( .A(n34595), .B(n34599), .Z(n34665) );
  AND U43637 ( .A(n34666), .B(n34667), .Z(n34599) );
  NAND U43638 ( .A(n34668), .B(n34669), .Z(n34667) );
  NAND U43639 ( .A(n34670), .B(n34671), .Z(n34666) );
  AND U43640 ( .A(n34672), .B(n34673), .Z(n34595) );
  NAND U43641 ( .A(n34674), .B(n34675), .Z(n34673) );
  NAND U43642 ( .A(n34676), .B(n34677), .Z(n34672) );
  NANDN U43643 ( .A(n34678), .B(n34679), .Z(n34598) );
  ANDN U43644 ( .B(n34680), .A(n34681), .Z(n34592) );
  XNOR U43645 ( .A(n34583), .B(n34682), .Z(n34588) );
  XNOR U43646 ( .A(n34581), .B(n34585), .Z(n34682) );
  AND U43647 ( .A(n34683), .B(n34684), .Z(n34585) );
  NAND U43648 ( .A(n34685), .B(n34686), .Z(n34684) );
  NAND U43649 ( .A(n34687), .B(n34688), .Z(n34683) );
  AND U43650 ( .A(n34689), .B(n34690), .Z(n34581) );
  NAND U43651 ( .A(n34691), .B(n34692), .Z(n34690) );
  NAND U43652 ( .A(n34693), .B(n34694), .Z(n34689) );
  AND U43653 ( .A(n34695), .B(n34696), .Z(n34583) );
  XOR U43654 ( .A(n34663), .B(n34662), .Z(N62308) );
  XNOR U43655 ( .A(n34680), .B(n34681), .Z(n34662) );
  XNOR U43656 ( .A(n34695), .B(n34696), .Z(n34681) );
  XOR U43657 ( .A(n34692), .B(n34691), .Z(n34696) );
  XOR U43658 ( .A(y[3180]), .B(x[3180]), .Z(n34691) );
  XOR U43659 ( .A(n34694), .B(n34693), .Z(n34692) );
  XOR U43660 ( .A(y[3182]), .B(x[3182]), .Z(n34693) );
  XOR U43661 ( .A(y[3181]), .B(x[3181]), .Z(n34694) );
  XOR U43662 ( .A(n34686), .B(n34685), .Z(n34695) );
  XOR U43663 ( .A(n34688), .B(n34687), .Z(n34685) );
  XOR U43664 ( .A(y[3179]), .B(x[3179]), .Z(n34687) );
  XOR U43665 ( .A(y[3178]), .B(x[3178]), .Z(n34688) );
  XOR U43666 ( .A(y[3177]), .B(x[3177]), .Z(n34686) );
  XNOR U43667 ( .A(n34679), .B(n34678), .Z(n34680) );
  XNOR U43668 ( .A(n34675), .B(n34674), .Z(n34678) );
  XOR U43669 ( .A(n34677), .B(n34676), .Z(n34674) );
  XOR U43670 ( .A(y[3176]), .B(x[3176]), .Z(n34676) );
  XOR U43671 ( .A(y[3175]), .B(x[3175]), .Z(n34677) );
  XOR U43672 ( .A(y[3174]), .B(x[3174]), .Z(n34675) );
  XOR U43673 ( .A(n34669), .B(n34668), .Z(n34679) );
  XOR U43674 ( .A(n34671), .B(n34670), .Z(n34668) );
  XOR U43675 ( .A(y[3173]), .B(x[3173]), .Z(n34670) );
  XOR U43676 ( .A(y[3172]), .B(x[3172]), .Z(n34671) );
  XOR U43677 ( .A(y[3171]), .B(x[3171]), .Z(n34669) );
  XNOR U43678 ( .A(n34645), .B(n34646), .Z(n34663) );
  XNOR U43679 ( .A(n34660), .B(n34661), .Z(n34646) );
  XOR U43680 ( .A(n34657), .B(n34656), .Z(n34661) );
  XOR U43681 ( .A(y[3168]), .B(x[3168]), .Z(n34656) );
  XOR U43682 ( .A(n34659), .B(n34658), .Z(n34657) );
  XOR U43683 ( .A(y[3170]), .B(x[3170]), .Z(n34658) );
  XOR U43684 ( .A(y[3169]), .B(x[3169]), .Z(n34659) );
  XOR U43685 ( .A(n34651), .B(n34650), .Z(n34660) );
  XOR U43686 ( .A(n34653), .B(n34652), .Z(n34650) );
  XOR U43687 ( .A(y[3167]), .B(x[3167]), .Z(n34652) );
  XOR U43688 ( .A(y[3166]), .B(x[3166]), .Z(n34653) );
  XOR U43689 ( .A(y[3165]), .B(x[3165]), .Z(n34651) );
  XNOR U43690 ( .A(n34644), .B(n34643), .Z(n34645) );
  XNOR U43691 ( .A(n34640), .B(n34639), .Z(n34643) );
  XOR U43692 ( .A(n34642), .B(n34641), .Z(n34639) );
  XOR U43693 ( .A(y[3164]), .B(x[3164]), .Z(n34641) );
  XOR U43694 ( .A(y[3163]), .B(x[3163]), .Z(n34642) );
  XOR U43695 ( .A(y[3162]), .B(x[3162]), .Z(n34640) );
  XOR U43696 ( .A(n34634), .B(n34633), .Z(n34644) );
  XOR U43697 ( .A(n34636), .B(n34635), .Z(n34633) );
  XOR U43698 ( .A(y[3161]), .B(x[3161]), .Z(n34635) );
  XOR U43699 ( .A(y[3160]), .B(x[3160]), .Z(n34636) );
  XOR U43700 ( .A(y[3159]), .B(x[3159]), .Z(n34634) );
  NAND U43701 ( .A(n34697), .B(n34698), .Z(N62299) );
  NAND U43702 ( .A(n34699), .B(n34700), .Z(n34698) );
  NANDN U43703 ( .A(n34701), .B(n34702), .Z(n34700) );
  NANDN U43704 ( .A(n34702), .B(n34701), .Z(n34697) );
  XOR U43705 ( .A(n34701), .B(n34703), .Z(N62298) );
  XNOR U43706 ( .A(n34699), .B(n34702), .Z(n34703) );
  NAND U43707 ( .A(n34704), .B(n34705), .Z(n34702) );
  NAND U43708 ( .A(n34706), .B(n34707), .Z(n34705) );
  NANDN U43709 ( .A(n34708), .B(n34709), .Z(n34707) );
  NANDN U43710 ( .A(n34709), .B(n34708), .Z(n34704) );
  AND U43711 ( .A(n34710), .B(n34711), .Z(n34699) );
  NAND U43712 ( .A(n34712), .B(n34713), .Z(n34711) );
  NANDN U43713 ( .A(n34714), .B(n34715), .Z(n34713) );
  NANDN U43714 ( .A(n34715), .B(n34714), .Z(n34710) );
  IV U43715 ( .A(n34716), .Z(n34715) );
  AND U43716 ( .A(n34717), .B(n34718), .Z(n34701) );
  NAND U43717 ( .A(n34719), .B(n34720), .Z(n34718) );
  NANDN U43718 ( .A(n34721), .B(n34722), .Z(n34720) );
  NANDN U43719 ( .A(n34722), .B(n34721), .Z(n34717) );
  XOR U43720 ( .A(n34714), .B(n34723), .Z(N62297) );
  XNOR U43721 ( .A(n34712), .B(n34716), .Z(n34723) );
  XOR U43722 ( .A(n34709), .B(n34724), .Z(n34716) );
  XNOR U43723 ( .A(n34706), .B(n34708), .Z(n34724) );
  AND U43724 ( .A(n34725), .B(n34726), .Z(n34708) );
  NANDN U43725 ( .A(n34727), .B(n34728), .Z(n34726) );
  OR U43726 ( .A(n34729), .B(n34730), .Z(n34728) );
  IV U43727 ( .A(n34731), .Z(n34730) );
  NANDN U43728 ( .A(n34731), .B(n34729), .Z(n34725) );
  AND U43729 ( .A(n34732), .B(n34733), .Z(n34706) );
  NAND U43730 ( .A(n34734), .B(n34735), .Z(n34733) );
  NANDN U43731 ( .A(n34736), .B(n34737), .Z(n34735) );
  NANDN U43732 ( .A(n34737), .B(n34736), .Z(n34732) );
  IV U43733 ( .A(n34738), .Z(n34737) );
  NAND U43734 ( .A(n34739), .B(n34740), .Z(n34709) );
  NANDN U43735 ( .A(n34741), .B(n34742), .Z(n34740) );
  NANDN U43736 ( .A(n34743), .B(n34744), .Z(n34742) );
  NANDN U43737 ( .A(n34744), .B(n34743), .Z(n34739) );
  IV U43738 ( .A(n34745), .Z(n34743) );
  AND U43739 ( .A(n34746), .B(n34747), .Z(n34712) );
  NAND U43740 ( .A(n34748), .B(n34749), .Z(n34747) );
  NANDN U43741 ( .A(n34750), .B(n34751), .Z(n34749) );
  NANDN U43742 ( .A(n34751), .B(n34750), .Z(n34746) );
  XOR U43743 ( .A(n34722), .B(n34752), .Z(n34714) );
  XNOR U43744 ( .A(n34719), .B(n34721), .Z(n34752) );
  AND U43745 ( .A(n34753), .B(n34754), .Z(n34721) );
  NANDN U43746 ( .A(n34755), .B(n34756), .Z(n34754) );
  OR U43747 ( .A(n34757), .B(n34758), .Z(n34756) );
  IV U43748 ( .A(n34759), .Z(n34758) );
  NANDN U43749 ( .A(n34759), .B(n34757), .Z(n34753) );
  AND U43750 ( .A(n34760), .B(n34761), .Z(n34719) );
  NAND U43751 ( .A(n34762), .B(n34763), .Z(n34761) );
  NANDN U43752 ( .A(n34764), .B(n34765), .Z(n34763) );
  NANDN U43753 ( .A(n34765), .B(n34764), .Z(n34760) );
  IV U43754 ( .A(n34766), .Z(n34765) );
  NAND U43755 ( .A(n34767), .B(n34768), .Z(n34722) );
  NANDN U43756 ( .A(n34769), .B(n34770), .Z(n34768) );
  NANDN U43757 ( .A(n34771), .B(n34772), .Z(n34770) );
  NANDN U43758 ( .A(n34772), .B(n34771), .Z(n34767) );
  IV U43759 ( .A(n34773), .Z(n34771) );
  XOR U43760 ( .A(n34748), .B(n34774), .Z(N62296) );
  XNOR U43761 ( .A(n34751), .B(n34750), .Z(n34774) );
  XNOR U43762 ( .A(n34762), .B(n34775), .Z(n34750) );
  XNOR U43763 ( .A(n34766), .B(n34764), .Z(n34775) );
  XOR U43764 ( .A(n34772), .B(n34776), .Z(n34764) );
  XNOR U43765 ( .A(n34769), .B(n34773), .Z(n34776) );
  AND U43766 ( .A(n34777), .B(n34778), .Z(n34773) );
  NAND U43767 ( .A(n34779), .B(n34780), .Z(n34778) );
  NAND U43768 ( .A(n34781), .B(n34782), .Z(n34777) );
  AND U43769 ( .A(n34783), .B(n34784), .Z(n34769) );
  NAND U43770 ( .A(n34785), .B(n34786), .Z(n34784) );
  NAND U43771 ( .A(n34787), .B(n34788), .Z(n34783) );
  NANDN U43772 ( .A(n34789), .B(n34790), .Z(n34772) );
  ANDN U43773 ( .B(n34791), .A(n34792), .Z(n34766) );
  XNOR U43774 ( .A(n34757), .B(n34793), .Z(n34762) );
  XNOR U43775 ( .A(n34755), .B(n34759), .Z(n34793) );
  AND U43776 ( .A(n34794), .B(n34795), .Z(n34759) );
  NAND U43777 ( .A(n34796), .B(n34797), .Z(n34795) );
  NAND U43778 ( .A(n34798), .B(n34799), .Z(n34794) );
  AND U43779 ( .A(n34800), .B(n34801), .Z(n34755) );
  NAND U43780 ( .A(n34802), .B(n34803), .Z(n34801) );
  NAND U43781 ( .A(n34804), .B(n34805), .Z(n34800) );
  AND U43782 ( .A(n34806), .B(n34807), .Z(n34757) );
  NAND U43783 ( .A(n34808), .B(n34809), .Z(n34751) );
  XNOR U43784 ( .A(n34734), .B(n34810), .Z(n34748) );
  XNOR U43785 ( .A(n34738), .B(n34736), .Z(n34810) );
  XOR U43786 ( .A(n34744), .B(n34811), .Z(n34736) );
  XNOR U43787 ( .A(n34741), .B(n34745), .Z(n34811) );
  AND U43788 ( .A(n34812), .B(n34813), .Z(n34745) );
  NAND U43789 ( .A(n34814), .B(n34815), .Z(n34813) );
  NAND U43790 ( .A(n34816), .B(n34817), .Z(n34812) );
  AND U43791 ( .A(n34818), .B(n34819), .Z(n34741) );
  NAND U43792 ( .A(n34820), .B(n34821), .Z(n34819) );
  NAND U43793 ( .A(n34822), .B(n34823), .Z(n34818) );
  NANDN U43794 ( .A(n34824), .B(n34825), .Z(n34744) );
  ANDN U43795 ( .B(n34826), .A(n34827), .Z(n34738) );
  XNOR U43796 ( .A(n34729), .B(n34828), .Z(n34734) );
  XNOR U43797 ( .A(n34727), .B(n34731), .Z(n34828) );
  AND U43798 ( .A(n34829), .B(n34830), .Z(n34731) );
  NAND U43799 ( .A(n34831), .B(n34832), .Z(n34830) );
  NAND U43800 ( .A(n34833), .B(n34834), .Z(n34829) );
  AND U43801 ( .A(n34835), .B(n34836), .Z(n34727) );
  NAND U43802 ( .A(n34837), .B(n34838), .Z(n34836) );
  NAND U43803 ( .A(n34839), .B(n34840), .Z(n34835) );
  AND U43804 ( .A(n34841), .B(n34842), .Z(n34729) );
  XOR U43805 ( .A(n34809), .B(n34808), .Z(N62295) );
  XNOR U43806 ( .A(n34826), .B(n34827), .Z(n34808) );
  XNOR U43807 ( .A(n34841), .B(n34842), .Z(n34827) );
  XOR U43808 ( .A(n34838), .B(n34837), .Z(n34842) );
  XOR U43809 ( .A(y[3156]), .B(x[3156]), .Z(n34837) );
  XOR U43810 ( .A(n34840), .B(n34839), .Z(n34838) );
  XOR U43811 ( .A(y[3158]), .B(x[3158]), .Z(n34839) );
  XOR U43812 ( .A(y[3157]), .B(x[3157]), .Z(n34840) );
  XOR U43813 ( .A(n34832), .B(n34831), .Z(n34841) );
  XOR U43814 ( .A(n34834), .B(n34833), .Z(n34831) );
  XOR U43815 ( .A(y[3155]), .B(x[3155]), .Z(n34833) );
  XOR U43816 ( .A(y[3154]), .B(x[3154]), .Z(n34834) );
  XOR U43817 ( .A(y[3153]), .B(x[3153]), .Z(n34832) );
  XNOR U43818 ( .A(n34825), .B(n34824), .Z(n34826) );
  XNOR U43819 ( .A(n34821), .B(n34820), .Z(n34824) );
  XOR U43820 ( .A(n34823), .B(n34822), .Z(n34820) );
  XOR U43821 ( .A(y[3152]), .B(x[3152]), .Z(n34822) );
  XOR U43822 ( .A(y[3151]), .B(x[3151]), .Z(n34823) );
  XOR U43823 ( .A(y[3150]), .B(x[3150]), .Z(n34821) );
  XOR U43824 ( .A(n34815), .B(n34814), .Z(n34825) );
  XOR U43825 ( .A(n34817), .B(n34816), .Z(n34814) );
  XOR U43826 ( .A(y[3149]), .B(x[3149]), .Z(n34816) );
  XOR U43827 ( .A(y[3148]), .B(x[3148]), .Z(n34817) );
  XOR U43828 ( .A(y[3147]), .B(x[3147]), .Z(n34815) );
  XNOR U43829 ( .A(n34791), .B(n34792), .Z(n34809) );
  XNOR U43830 ( .A(n34806), .B(n34807), .Z(n34792) );
  XOR U43831 ( .A(n34803), .B(n34802), .Z(n34807) );
  XOR U43832 ( .A(y[3144]), .B(x[3144]), .Z(n34802) );
  XOR U43833 ( .A(n34805), .B(n34804), .Z(n34803) );
  XOR U43834 ( .A(y[3146]), .B(x[3146]), .Z(n34804) );
  XOR U43835 ( .A(y[3145]), .B(x[3145]), .Z(n34805) );
  XOR U43836 ( .A(n34797), .B(n34796), .Z(n34806) );
  XOR U43837 ( .A(n34799), .B(n34798), .Z(n34796) );
  XOR U43838 ( .A(y[3143]), .B(x[3143]), .Z(n34798) );
  XOR U43839 ( .A(y[3142]), .B(x[3142]), .Z(n34799) );
  XOR U43840 ( .A(y[3141]), .B(x[3141]), .Z(n34797) );
  XNOR U43841 ( .A(n34790), .B(n34789), .Z(n34791) );
  XNOR U43842 ( .A(n34786), .B(n34785), .Z(n34789) );
  XOR U43843 ( .A(n34788), .B(n34787), .Z(n34785) );
  XOR U43844 ( .A(y[3140]), .B(x[3140]), .Z(n34787) );
  XOR U43845 ( .A(y[3139]), .B(x[3139]), .Z(n34788) );
  XOR U43846 ( .A(y[3138]), .B(x[3138]), .Z(n34786) );
  XOR U43847 ( .A(n34780), .B(n34779), .Z(n34790) );
  XOR U43848 ( .A(n34782), .B(n34781), .Z(n34779) );
  XOR U43849 ( .A(y[3137]), .B(x[3137]), .Z(n34781) );
  XOR U43850 ( .A(y[3136]), .B(x[3136]), .Z(n34782) );
  XOR U43851 ( .A(y[3135]), .B(x[3135]), .Z(n34780) );
  NAND U43852 ( .A(n34843), .B(n34844), .Z(N62286) );
  NAND U43853 ( .A(n34845), .B(n34846), .Z(n34844) );
  NANDN U43854 ( .A(n34847), .B(n34848), .Z(n34846) );
  NANDN U43855 ( .A(n34848), .B(n34847), .Z(n34843) );
  XOR U43856 ( .A(n34847), .B(n34849), .Z(N62285) );
  XNOR U43857 ( .A(n34845), .B(n34848), .Z(n34849) );
  NAND U43858 ( .A(n34850), .B(n34851), .Z(n34848) );
  NAND U43859 ( .A(n34852), .B(n34853), .Z(n34851) );
  NANDN U43860 ( .A(n34854), .B(n34855), .Z(n34853) );
  NANDN U43861 ( .A(n34855), .B(n34854), .Z(n34850) );
  AND U43862 ( .A(n34856), .B(n34857), .Z(n34845) );
  NAND U43863 ( .A(n34858), .B(n34859), .Z(n34857) );
  NANDN U43864 ( .A(n34860), .B(n34861), .Z(n34859) );
  NANDN U43865 ( .A(n34861), .B(n34860), .Z(n34856) );
  IV U43866 ( .A(n34862), .Z(n34861) );
  AND U43867 ( .A(n34863), .B(n34864), .Z(n34847) );
  NAND U43868 ( .A(n34865), .B(n34866), .Z(n34864) );
  NANDN U43869 ( .A(n34867), .B(n34868), .Z(n34866) );
  NANDN U43870 ( .A(n34868), .B(n34867), .Z(n34863) );
  XOR U43871 ( .A(n34860), .B(n34869), .Z(N62284) );
  XNOR U43872 ( .A(n34858), .B(n34862), .Z(n34869) );
  XOR U43873 ( .A(n34855), .B(n34870), .Z(n34862) );
  XNOR U43874 ( .A(n34852), .B(n34854), .Z(n34870) );
  AND U43875 ( .A(n34871), .B(n34872), .Z(n34854) );
  NANDN U43876 ( .A(n34873), .B(n34874), .Z(n34872) );
  OR U43877 ( .A(n34875), .B(n34876), .Z(n34874) );
  IV U43878 ( .A(n34877), .Z(n34876) );
  NANDN U43879 ( .A(n34877), .B(n34875), .Z(n34871) );
  AND U43880 ( .A(n34878), .B(n34879), .Z(n34852) );
  NAND U43881 ( .A(n34880), .B(n34881), .Z(n34879) );
  NANDN U43882 ( .A(n34882), .B(n34883), .Z(n34881) );
  NANDN U43883 ( .A(n34883), .B(n34882), .Z(n34878) );
  IV U43884 ( .A(n34884), .Z(n34883) );
  NAND U43885 ( .A(n34885), .B(n34886), .Z(n34855) );
  NANDN U43886 ( .A(n34887), .B(n34888), .Z(n34886) );
  NANDN U43887 ( .A(n34889), .B(n34890), .Z(n34888) );
  NANDN U43888 ( .A(n34890), .B(n34889), .Z(n34885) );
  IV U43889 ( .A(n34891), .Z(n34889) );
  AND U43890 ( .A(n34892), .B(n34893), .Z(n34858) );
  NAND U43891 ( .A(n34894), .B(n34895), .Z(n34893) );
  NANDN U43892 ( .A(n34896), .B(n34897), .Z(n34895) );
  NANDN U43893 ( .A(n34897), .B(n34896), .Z(n34892) );
  XOR U43894 ( .A(n34868), .B(n34898), .Z(n34860) );
  XNOR U43895 ( .A(n34865), .B(n34867), .Z(n34898) );
  AND U43896 ( .A(n34899), .B(n34900), .Z(n34867) );
  NANDN U43897 ( .A(n34901), .B(n34902), .Z(n34900) );
  OR U43898 ( .A(n34903), .B(n34904), .Z(n34902) );
  IV U43899 ( .A(n34905), .Z(n34904) );
  NANDN U43900 ( .A(n34905), .B(n34903), .Z(n34899) );
  AND U43901 ( .A(n34906), .B(n34907), .Z(n34865) );
  NAND U43902 ( .A(n34908), .B(n34909), .Z(n34907) );
  NANDN U43903 ( .A(n34910), .B(n34911), .Z(n34909) );
  NANDN U43904 ( .A(n34911), .B(n34910), .Z(n34906) );
  IV U43905 ( .A(n34912), .Z(n34911) );
  NAND U43906 ( .A(n34913), .B(n34914), .Z(n34868) );
  NANDN U43907 ( .A(n34915), .B(n34916), .Z(n34914) );
  NANDN U43908 ( .A(n34917), .B(n34918), .Z(n34916) );
  NANDN U43909 ( .A(n34918), .B(n34917), .Z(n34913) );
  IV U43910 ( .A(n34919), .Z(n34917) );
  XOR U43911 ( .A(n34894), .B(n34920), .Z(N62283) );
  XNOR U43912 ( .A(n34897), .B(n34896), .Z(n34920) );
  XNOR U43913 ( .A(n34908), .B(n34921), .Z(n34896) );
  XNOR U43914 ( .A(n34912), .B(n34910), .Z(n34921) );
  XOR U43915 ( .A(n34918), .B(n34922), .Z(n34910) );
  XNOR U43916 ( .A(n34915), .B(n34919), .Z(n34922) );
  AND U43917 ( .A(n34923), .B(n34924), .Z(n34919) );
  NAND U43918 ( .A(n34925), .B(n34926), .Z(n34924) );
  NAND U43919 ( .A(n34927), .B(n34928), .Z(n34923) );
  AND U43920 ( .A(n34929), .B(n34930), .Z(n34915) );
  NAND U43921 ( .A(n34931), .B(n34932), .Z(n34930) );
  NAND U43922 ( .A(n34933), .B(n34934), .Z(n34929) );
  NANDN U43923 ( .A(n34935), .B(n34936), .Z(n34918) );
  ANDN U43924 ( .B(n34937), .A(n34938), .Z(n34912) );
  XNOR U43925 ( .A(n34903), .B(n34939), .Z(n34908) );
  XNOR U43926 ( .A(n34901), .B(n34905), .Z(n34939) );
  AND U43927 ( .A(n34940), .B(n34941), .Z(n34905) );
  NAND U43928 ( .A(n34942), .B(n34943), .Z(n34941) );
  NAND U43929 ( .A(n34944), .B(n34945), .Z(n34940) );
  AND U43930 ( .A(n34946), .B(n34947), .Z(n34901) );
  NAND U43931 ( .A(n34948), .B(n34949), .Z(n34947) );
  NAND U43932 ( .A(n34950), .B(n34951), .Z(n34946) );
  AND U43933 ( .A(n34952), .B(n34953), .Z(n34903) );
  NAND U43934 ( .A(n34954), .B(n34955), .Z(n34897) );
  XNOR U43935 ( .A(n34880), .B(n34956), .Z(n34894) );
  XNOR U43936 ( .A(n34884), .B(n34882), .Z(n34956) );
  XOR U43937 ( .A(n34890), .B(n34957), .Z(n34882) );
  XNOR U43938 ( .A(n34887), .B(n34891), .Z(n34957) );
  AND U43939 ( .A(n34958), .B(n34959), .Z(n34891) );
  NAND U43940 ( .A(n34960), .B(n34961), .Z(n34959) );
  NAND U43941 ( .A(n34962), .B(n34963), .Z(n34958) );
  AND U43942 ( .A(n34964), .B(n34965), .Z(n34887) );
  NAND U43943 ( .A(n34966), .B(n34967), .Z(n34965) );
  NAND U43944 ( .A(n34968), .B(n34969), .Z(n34964) );
  NANDN U43945 ( .A(n34970), .B(n34971), .Z(n34890) );
  ANDN U43946 ( .B(n34972), .A(n34973), .Z(n34884) );
  XNOR U43947 ( .A(n34875), .B(n34974), .Z(n34880) );
  XNOR U43948 ( .A(n34873), .B(n34877), .Z(n34974) );
  AND U43949 ( .A(n34975), .B(n34976), .Z(n34877) );
  NAND U43950 ( .A(n34977), .B(n34978), .Z(n34976) );
  NAND U43951 ( .A(n34979), .B(n34980), .Z(n34975) );
  AND U43952 ( .A(n34981), .B(n34982), .Z(n34873) );
  NAND U43953 ( .A(n34983), .B(n34984), .Z(n34982) );
  NAND U43954 ( .A(n34985), .B(n34986), .Z(n34981) );
  AND U43955 ( .A(n34987), .B(n34988), .Z(n34875) );
  XOR U43956 ( .A(n34955), .B(n34954), .Z(N62282) );
  XNOR U43957 ( .A(n34972), .B(n34973), .Z(n34954) );
  XNOR U43958 ( .A(n34987), .B(n34988), .Z(n34973) );
  XOR U43959 ( .A(n34984), .B(n34983), .Z(n34988) );
  XOR U43960 ( .A(y[3132]), .B(x[3132]), .Z(n34983) );
  XOR U43961 ( .A(n34986), .B(n34985), .Z(n34984) );
  XOR U43962 ( .A(y[3134]), .B(x[3134]), .Z(n34985) );
  XOR U43963 ( .A(y[3133]), .B(x[3133]), .Z(n34986) );
  XOR U43964 ( .A(n34978), .B(n34977), .Z(n34987) );
  XOR U43965 ( .A(n34980), .B(n34979), .Z(n34977) );
  XOR U43966 ( .A(y[3131]), .B(x[3131]), .Z(n34979) );
  XOR U43967 ( .A(y[3130]), .B(x[3130]), .Z(n34980) );
  XOR U43968 ( .A(y[3129]), .B(x[3129]), .Z(n34978) );
  XNOR U43969 ( .A(n34971), .B(n34970), .Z(n34972) );
  XNOR U43970 ( .A(n34967), .B(n34966), .Z(n34970) );
  XOR U43971 ( .A(n34969), .B(n34968), .Z(n34966) );
  XOR U43972 ( .A(y[3128]), .B(x[3128]), .Z(n34968) );
  XOR U43973 ( .A(y[3127]), .B(x[3127]), .Z(n34969) );
  XOR U43974 ( .A(y[3126]), .B(x[3126]), .Z(n34967) );
  XOR U43975 ( .A(n34961), .B(n34960), .Z(n34971) );
  XOR U43976 ( .A(n34963), .B(n34962), .Z(n34960) );
  XOR U43977 ( .A(y[3125]), .B(x[3125]), .Z(n34962) );
  XOR U43978 ( .A(y[3124]), .B(x[3124]), .Z(n34963) );
  XOR U43979 ( .A(y[3123]), .B(x[3123]), .Z(n34961) );
  XNOR U43980 ( .A(n34937), .B(n34938), .Z(n34955) );
  XNOR U43981 ( .A(n34952), .B(n34953), .Z(n34938) );
  XOR U43982 ( .A(n34949), .B(n34948), .Z(n34953) );
  XOR U43983 ( .A(y[3120]), .B(x[3120]), .Z(n34948) );
  XOR U43984 ( .A(n34951), .B(n34950), .Z(n34949) );
  XOR U43985 ( .A(y[3122]), .B(x[3122]), .Z(n34950) );
  XOR U43986 ( .A(y[3121]), .B(x[3121]), .Z(n34951) );
  XOR U43987 ( .A(n34943), .B(n34942), .Z(n34952) );
  XOR U43988 ( .A(n34945), .B(n34944), .Z(n34942) );
  XOR U43989 ( .A(y[3119]), .B(x[3119]), .Z(n34944) );
  XOR U43990 ( .A(y[3118]), .B(x[3118]), .Z(n34945) );
  XOR U43991 ( .A(y[3117]), .B(x[3117]), .Z(n34943) );
  XNOR U43992 ( .A(n34936), .B(n34935), .Z(n34937) );
  XNOR U43993 ( .A(n34932), .B(n34931), .Z(n34935) );
  XOR U43994 ( .A(n34934), .B(n34933), .Z(n34931) );
  XOR U43995 ( .A(y[3116]), .B(x[3116]), .Z(n34933) );
  XOR U43996 ( .A(y[3115]), .B(x[3115]), .Z(n34934) );
  XOR U43997 ( .A(y[3114]), .B(x[3114]), .Z(n34932) );
  XOR U43998 ( .A(n34926), .B(n34925), .Z(n34936) );
  XOR U43999 ( .A(n34928), .B(n34927), .Z(n34925) );
  XOR U44000 ( .A(y[3113]), .B(x[3113]), .Z(n34927) );
  XOR U44001 ( .A(y[3112]), .B(x[3112]), .Z(n34928) );
  XOR U44002 ( .A(y[3111]), .B(x[3111]), .Z(n34926) );
  NAND U44003 ( .A(n34989), .B(n34990), .Z(N62273) );
  NAND U44004 ( .A(n34991), .B(n34992), .Z(n34990) );
  NANDN U44005 ( .A(n34993), .B(n34994), .Z(n34992) );
  NANDN U44006 ( .A(n34994), .B(n34993), .Z(n34989) );
  XOR U44007 ( .A(n34993), .B(n34995), .Z(N62272) );
  XNOR U44008 ( .A(n34991), .B(n34994), .Z(n34995) );
  NAND U44009 ( .A(n34996), .B(n34997), .Z(n34994) );
  NAND U44010 ( .A(n34998), .B(n34999), .Z(n34997) );
  NANDN U44011 ( .A(n35000), .B(n35001), .Z(n34999) );
  NANDN U44012 ( .A(n35001), .B(n35000), .Z(n34996) );
  AND U44013 ( .A(n35002), .B(n35003), .Z(n34991) );
  NAND U44014 ( .A(n35004), .B(n35005), .Z(n35003) );
  NANDN U44015 ( .A(n35006), .B(n35007), .Z(n35005) );
  NANDN U44016 ( .A(n35007), .B(n35006), .Z(n35002) );
  IV U44017 ( .A(n35008), .Z(n35007) );
  AND U44018 ( .A(n35009), .B(n35010), .Z(n34993) );
  NAND U44019 ( .A(n35011), .B(n35012), .Z(n35010) );
  NANDN U44020 ( .A(n35013), .B(n35014), .Z(n35012) );
  NANDN U44021 ( .A(n35014), .B(n35013), .Z(n35009) );
  XOR U44022 ( .A(n35006), .B(n35015), .Z(N62271) );
  XNOR U44023 ( .A(n35004), .B(n35008), .Z(n35015) );
  XOR U44024 ( .A(n35001), .B(n35016), .Z(n35008) );
  XNOR U44025 ( .A(n34998), .B(n35000), .Z(n35016) );
  AND U44026 ( .A(n35017), .B(n35018), .Z(n35000) );
  NANDN U44027 ( .A(n35019), .B(n35020), .Z(n35018) );
  OR U44028 ( .A(n35021), .B(n35022), .Z(n35020) );
  IV U44029 ( .A(n35023), .Z(n35022) );
  NANDN U44030 ( .A(n35023), .B(n35021), .Z(n35017) );
  AND U44031 ( .A(n35024), .B(n35025), .Z(n34998) );
  NAND U44032 ( .A(n35026), .B(n35027), .Z(n35025) );
  NANDN U44033 ( .A(n35028), .B(n35029), .Z(n35027) );
  NANDN U44034 ( .A(n35029), .B(n35028), .Z(n35024) );
  IV U44035 ( .A(n35030), .Z(n35029) );
  NAND U44036 ( .A(n35031), .B(n35032), .Z(n35001) );
  NANDN U44037 ( .A(n35033), .B(n35034), .Z(n35032) );
  NANDN U44038 ( .A(n35035), .B(n35036), .Z(n35034) );
  NANDN U44039 ( .A(n35036), .B(n35035), .Z(n35031) );
  IV U44040 ( .A(n35037), .Z(n35035) );
  AND U44041 ( .A(n35038), .B(n35039), .Z(n35004) );
  NAND U44042 ( .A(n35040), .B(n35041), .Z(n35039) );
  NANDN U44043 ( .A(n35042), .B(n35043), .Z(n35041) );
  NANDN U44044 ( .A(n35043), .B(n35042), .Z(n35038) );
  XOR U44045 ( .A(n35014), .B(n35044), .Z(n35006) );
  XNOR U44046 ( .A(n35011), .B(n35013), .Z(n35044) );
  AND U44047 ( .A(n35045), .B(n35046), .Z(n35013) );
  NANDN U44048 ( .A(n35047), .B(n35048), .Z(n35046) );
  OR U44049 ( .A(n35049), .B(n35050), .Z(n35048) );
  IV U44050 ( .A(n35051), .Z(n35050) );
  NANDN U44051 ( .A(n35051), .B(n35049), .Z(n35045) );
  AND U44052 ( .A(n35052), .B(n35053), .Z(n35011) );
  NAND U44053 ( .A(n35054), .B(n35055), .Z(n35053) );
  NANDN U44054 ( .A(n35056), .B(n35057), .Z(n35055) );
  NANDN U44055 ( .A(n35057), .B(n35056), .Z(n35052) );
  IV U44056 ( .A(n35058), .Z(n35057) );
  NAND U44057 ( .A(n35059), .B(n35060), .Z(n35014) );
  NANDN U44058 ( .A(n35061), .B(n35062), .Z(n35060) );
  NANDN U44059 ( .A(n35063), .B(n35064), .Z(n35062) );
  NANDN U44060 ( .A(n35064), .B(n35063), .Z(n35059) );
  IV U44061 ( .A(n35065), .Z(n35063) );
  XOR U44062 ( .A(n35040), .B(n35066), .Z(N62270) );
  XNOR U44063 ( .A(n35043), .B(n35042), .Z(n35066) );
  XNOR U44064 ( .A(n35054), .B(n35067), .Z(n35042) );
  XNOR U44065 ( .A(n35058), .B(n35056), .Z(n35067) );
  XOR U44066 ( .A(n35064), .B(n35068), .Z(n35056) );
  XNOR U44067 ( .A(n35061), .B(n35065), .Z(n35068) );
  AND U44068 ( .A(n35069), .B(n35070), .Z(n35065) );
  NAND U44069 ( .A(n35071), .B(n35072), .Z(n35070) );
  NAND U44070 ( .A(n35073), .B(n35074), .Z(n35069) );
  AND U44071 ( .A(n35075), .B(n35076), .Z(n35061) );
  NAND U44072 ( .A(n35077), .B(n35078), .Z(n35076) );
  NAND U44073 ( .A(n35079), .B(n35080), .Z(n35075) );
  NANDN U44074 ( .A(n35081), .B(n35082), .Z(n35064) );
  ANDN U44075 ( .B(n35083), .A(n35084), .Z(n35058) );
  XNOR U44076 ( .A(n35049), .B(n35085), .Z(n35054) );
  XNOR U44077 ( .A(n35047), .B(n35051), .Z(n35085) );
  AND U44078 ( .A(n35086), .B(n35087), .Z(n35051) );
  NAND U44079 ( .A(n35088), .B(n35089), .Z(n35087) );
  NAND U44080 ( .A(n35090), .B(n35091), .Z(n35086) );
  AND U44081 ( .A(n35092), .B(n35093), .Z(n35047) );
  NAND U44082 ( .A(n35094), .B(n35095), .Z(n35093) );
  NAND U44083 ( .A(n35096), .B(n35097), .Z(n35092) );
  AND U44084 ( .A(n35098), .B(n35099), .Z(n35049) );
  NAND U44085 ( .A(n35100), .B(n35101), .Z(n35043) );
  XNOR U44086 ( .A(n35026), .B(n35102), .Z(n35040) );
  XNOR U44087 ( .A(n35030), .B(n35028), .Z(n35102) );
  XOR U44088 ( .A(n35036), .B(n35103), .Z(n35028) );
  XNOR U44089 ( .A(n35033), .B(n35037), .Z(n35103) );
  AND U44090 ( .A(n35104), .B(n35105), .Z(n35037) );
  NAND U44091 ( .A(n35106), .B(n35107), .Z(n35105) );
  NAND U44092 ( .A(n35108), .B(n35109), .Z(n35104) );
  AND U44093 ( .A(n35110), .B(n35111), .Z(n35033) );
  NAND U44094 ( .A(n35112), .B(n35113), .Z(n35111) );
  NAND U44095 ( .A(n35114), .B(n35115), .Z(n35110) );
  NANDN U44096 ( .A(n35116), .B(n35117), .Z(n35036) );
  ANDN U44097 ( .B(n35118), .A(n35119), .Z(n35030) );
  XNOR U44098 ( .A(n35021), .B(n35120), .Z(n35026) );
  XNOR U44099 ( .A(n35019), .B(n35023), .Z(n35120) );
  AND U44100 ( .A(n35121), .B(n35122), .Z(n35023) );
  NAND U44101 ( .A(n35123), .B(n35124), .Z(n35122) );
  NAND U44102 ( .A(n35125), .B(n35126), .Z(n35121) );
  AND U44103 ( .A(n35127), .B(n35128), .Z(n35019) );
  NAND U44104 ( .A(n35129), .B(n35130), .Z(n35128) );
  NAND U44105 ( .A(n35131), .B(n35132), .Z(n35127) );
  AND U44106 ( .A(n35133), .B(n35134), .Z(n35021) );
  XOR U44107 ( .A(n35101), .B(n35100), .Z(N62269) );
  XNOR U44108 ( .A(n35118), .B(n35119), .Z(n35100) );
  XNOR U44109 ( .A(n35133), .B(n35134), .Z(n35119) );
  XOR U44110 ( .A(n35130), .B(n35129), .Z(n35134) );
  XOR U44111 ( .A(y[3108]), .B(x[3108]), .Z(n35129) );
  XOR U44112 ( .A(n35132), .B(n35131), .Z(n35130) );
  XOR U44113 ( .A(y[3110]), .B(x[3110]), .Z(n35131) );
  XOR U44114 ( .A(y[3109]), .B(x[3109]), .Z(n35132) );
  XOR U44115 ( .A(n35124), .B(n35123), .Z(n35133) );
  XOR U44116 ( .A(n35126), .B(n35125), .Z(n35123) );
  XOR U44117 ( .A(y[3107]), .B(x[3107]), .Z(n35125) );
  XOR U44118 ( .A(y[3106]), .B(x[3106]), .Z(n35126) );
  XOR U44119 ( .A(y[3105]), .B(x[3105]), .Z(n35124) );
  XNOR U44120 ( .A(n35117), .B(n35116), .Z(n35118) );
  XNOR U44121 ( .A(n35113), .B(n35112), .Z(n35116) );
  XOR U44122 ( .A(n35115), .B(n35114), .Z(n35112) );
  XOR U44123 ( .A(y[3104]), .B(x[3104]), .Z(n35114) );
  XOR U44124 ( .A(y[3103]), .B(x[3103]), .Z(n35115) );
  XOR U44125 ( .A(y[3102]), .B(x[3102]), .Z(n35113) );
  XOR U44126 ( .A(n35107), .B(n35106), .Z(n35117) );
  XOR U44127 ( .A(n35109), .B(n35108), .Z(n35106) );
  XOR U44128 ( .A(y[3101]), .B(x[3101]), .Z(n35108) );
  XOR U44129 ( .A(y[3100]), .B(x[3100]), .Z(n35109) );
  XOR U44130 ( .A(y[3099]), .B(x[3099]), .Z(n35107) );
  XNOR U44131 ( .A(n35083), .B(n35084), .Z(n35101) );
  XNOR U44132 ( .A(n35098), .B(n35099), .Z(n35084) );
  XOR U44133 ( .A(n35095), .B(n35094), .Z(n35099) );
  XOR U44134 ( .A(y[3096]), .B(x[3096]), .Z(n35094) );
  XOR U44135 ( .A(n35097), .B(n35096), .Z(n35095) );
  XOR U44136 ( .A(y[3098]), .B(x[3098]), .Z(n35096) );
  XOR U44137 ( .A(y[3097]), .B(x[3097]), .Z(n35097) );
  XOR U44138 ( .A(n35089), .B(n35088), .Z(n35098) );
  XOR U44139 ( .A(n35091), .B(n35090), .Z(n35088) );
  XOR U44140 ( .A(y[3095]), .B(x[3095]), .Z(n35090) );
  XOR U44141 ( .A(y[3094]), .B(x[3094]), .Z(n35091) );
  XOR U44142 ( .A(y[3093]), .B(x[3093]), .Z(n35089) );
  XNOR U44143 ( .A(n35082), .B(n35081), .Z(n35083) );
  XNOR U44144 ( .A(n35078), .B(n35077), .Z(n35081) );
  XOR U44145 ( .A(n35080), .B(n35079), .Z(n35077) );
  XOR U44146 ( .A(y[3092]), .B(x[3092]), .Z(n35079) );
  XOR U44147 ( .A(y[3091]), .B(x[3091]), .Z(n35080) );
  XOR U44148 ( .A(y[3090]), .B(x[3090]), .Z(n35078) );
  XOR U44149 ( .A(n35072), .B(n35071), .Z(n35082) );
  XOR U44150 ( .A(n35074), .B(n35073), .Z(n35071) );
  XOR U44151 ( .A(y[3089]), .B(x[3089]), .Z(n35073) );
  XOR U44152 ( .A(y[3088]), .B(x[3088]), .Z(n35074) );
  XOR U44153 ( .A(y[3087]), .B(x[3087]), .Z(n35072) );
  NAND U44154 ( .A(n35135), .B(n35136), .Z(N62260) );
  NAND U44155 ( .A(n35137), .B(n35138), .Z(n35136) );
  NANDN U44156 ( .A(n35139), .B(n35140), .Z(n35138) );
  NANDN U44157 ( .A(n35140), .B(n35139), .Z(n35135) );
  XOR U44158 ( .A(n35139), .B(n35141), .Z(N62259) );
  XNOR U44159 ( .A(n35137), .B(n35140), .Z(n35141) );
  NAND U44160 ( .A(n35142), .B(n35143), .Z(n35140) );
  NAND U44161 ( .A(n35144), .B(n35145), .Z(n35143) );
  NANDN U44162 ( .A(n35146), .B(n35147), .Z(n35145) );
  NANDN U44163 ( .A(n35147), .B(n35146), .Z(n35142) );
  AND U44164 ( .A(n35148), .B(n35149), .Z(n35137) );
  NAND U44165 ( .A(n35150), .B(n35151), .Z(n35149) );
  NANDN U44166 ( .A(n35152), .B(n35153), .Z(n35151) );
  NANDN U44167 ( .A(n35153), .B(n35152), .Z(n35148) );
  IV U44168 ( .A(n35154), .Z(n35153) );
  AND U44169 ( .A(n35155), .B(n35156), .Z(n35139) );
  NAND U44170 ( .A(n35157), .B(n35158), .Z(n35156) );
  NANDN U44171 ( .A(n35159), .B(n35160), .Z(n35158) );
  NANDN U44172 ( .A(n35160), .B(n35159), .Z(n35155) );
  XOR U44173 ( .A(n35152), .B(n35161), .Z(N62258) );
  XNOR U44174 ( .A(n35150), .B(n35154), .Z(n35161) );
  XOR U44175 ( .A(n35147), .B(n35162), .Z(n35154) );
  XNOR U44176 ( .A(n35144), .B(n35146), .Z(n35162) );
  AND U44177 ( .A(n35163), .B(n35164), .Z(n35146) );
  NANDN U44178 ( .A(n35165), .B(n35166), .Z(n35164) );
  OR U44179 ( .A(n35167), .B(n35168), .Z(n35166) );
  IV U44180 ( .A(n35169), .Z(n35168) );
  NANDN U44181 ( .A(n35169), .B(n35167), .Z(n35163) );
  AND U44182 ( .A(n35170), .B(n35171), .Z(n35144) );
  NAND U44183 ( .A(n35172), .B(n35173), .Z(n35171) );
  NANDN U44184 ( .A(n35174), .B(n35175), .Z(n35173) );
  NANDN U44185 ( .A(n35175), .B(n35174), .Z(n35170) );
  IV U44186 ( .A(n35176), .Z(n35175) );
  NAND U44187 ( .A(n35177), .B(n35178), .Z(n35147) );
  NANDN U44188 ( .A(n35179), .B(n35180), .Z(n35178) );
  NANDN U44189 ( .A(n35181), .B(n35182), .Z(n35180) );
  NANDN U44190 ( .A(n35182), .B(n35181), .Z(n35177) );
  IV U44191 ( .A(n35183), .Z(n35181) );
  AND U44192 ( .A(n35184), .B(n35185), .Z(n35150) );
  NAND U44193 ( .A(n35186), .B(n35187), .Z(n35185) );
  NANDN U44194 ( .A(n35188), .B(n35189), .Z(n35187) );
  NANDN U44195 ( .A(n35189), .B(n35188), .Z(n35184) );
  XOR U44196 ( .A(n35160), .B(n35190), .Z(n35152) );
  XNOR U44197 ( .A(n35157), .B(n35159), .Z(n35190) );
  AND U44198 ( .A(n35191), .B(n35192), .Z(n35159) );
  NANDN U44199 ( .A(n35193), .B(n35194), .Z(n35192) );
  OR U44200 ( .A(n35195), .B(n35196), .Z(n35194) );
  IV U44201 ( .A(n35197), .Z(n35196) );
  NANDN U44202 ( .A(n35197), .B(n35195), .Z(n35191) );
  AND U44203 ( .A(n35198), .B(n35199), .Z(n35157) );
  NAND U44204 ( .A(n35200), .B(n35201), .Z(n35199) );
  NANDN U44205 ( .A(n35202), .B(n35203), .Z(n35201) );
  NANDN U44206 ( .A(n35203), .B(n35202), .Z(n35198) );
  IV U44207 ( .A(n35204), .Z(n35203) );
  NAND U44208 ( .A(n35205), .B(n35206), .Z(n35160) );
  NANDN U44209 ( .A(n35207), .B(n35208), .Z(n35206) );
  NANDN U44210 ( .A(n35209), .B(n35210), .Z(n35208) );
  NANDN U44211 ( .A(n35210), .B(n35209), .Z(n35205) );
  IV U44212 ( .A(n35211), .Z(n35209) );
  XOR U44213 ( .A(n35186), .B(n35212), .Z(N62257) );
  XNOR U44214 ( .A(n35189), .B(n35188), .Z(n35212) );
  XNOR U44215 ( .A(n35200), .B(n35213), .Z(n35188) );
  XNOR U44216 ( .A(n35204), .B(n35202), .Z(n35213) );
  XOR U44217 ( .A(n35210), .B(n35214), .Z(n35202) );
  XNOR U44218 ( .A(n35207), .B(n35211), .Z(n35214) );
  AND U44219 ( .A(n35215), .B(n35216), .Z(n35211) );
  NAND U44220 ( .A(n35217), .B(n35218), .Z(n35216) );
  NAND U44221 ( .A(n35219), .B(n35220), .Z(n35215) );
  AND U44222 ( .A(n35221), .B(n35222), .Z(n35207) );
  NAND U44223 ( .A(n35223), .B(n35224), .Z(n35222) );
  NAND U44224 ( .A(n35225), .B(n35226), .Z(n35221) );
  NANDN U44225 ( .A(n35227), .B(n35228), .Z(n35210) );
  ANDN U44226 ( .B(n35229), .A(n35230), .Z(n35204) );
  XNOR U44227 ( .A(n35195), .B(n35231), .Z(n35200) );
  XNOR U44228 ( .A(n35193), .B(n35197), .Z(n35231) );
  AND U44229 ( .A(n35232), .B(n35233), .Z(n35197) );
  NAND U44230 ( .A(n35234), .B(n35235), .Z(n35233) );
  NAND U44231 ( .A(n35236), .B(n35237), .Z(n35232) );
  AND U44232 ( .A(n35238), .B(n35239), .Z(n35193) );
  NAND U44233 ( .A(n35240), .B(n35241), .Z(n35239) );
  NAND U44234 ( .A(n35242), .B(n35243), .Z(n35238) );
  AND U44235 ( .A(n35244), .B(n35245), .Z(n35195) );
  NAND U44236 ( .A(n35246), .B(n35247), .Z(n35189) );
  XNOR U44237 ( .A(n35172), .B(n35248), .Z(n35186) );
  XNOR U44238 ( .A(n35176), .B(n35174), .Z(n35248) );
  XOR U44239 ( .A(n35182), .B(n35249), .Z(n35174) );
  XNOR U44240 ( .A(n35179), .B(n35183), .Z(n35249) );
  AND U44241 ( .A(n35250), .B(n35251), .Z(n35183) );
  NAND U44242 ( .A(n35252), .B(n35253), .Z(n35251) );
  NAND U44243 ( .A(n35254), .B(n35255), .Z(n35250) );
  AND U44244 ( .A(n35256), .B(n35257), .Z(n35179) );
  NAND U44245 ( .A(n35258), .B(n35259), .Z(n35257) );
  NAND U44246 ( .A(n35260), .B(n35261), .Z(n35256) );
  NANDN U44247 ( .A(n35262), .B(n35263), .Z(n35182) );
  ANDN U44248 ( .B(n35264), .A(n35265), .Z(n35176) );
  XNOR U44249 ( .A(n35167), .B(n35266), .Z(n35172) );
  XNOR U44250 ( .A(n35165), .B(n35169), .Z(n35266) );
  AND U44251 ( .A(n35267), .B(n35268), .Z(n35169) );
  NAND U44252 ( .A(n35269), .B(n35270), .Z(n35268) );
  NAND U44253 ( .A(n35271), .B(n35272), .Z(n35267) );
  AND U44254 ( .A(n35273), .B(n35274), .Z(n35165) );
  NAND U44255 ( .A(n35275), .B(n35276), .Z(n35274) );
  NAND U44256 ( .A(n35277), .B(n35278), .Z(n35273) );
  AND U44257 ( .A(n35279), .B(n35280), .Z(n35167) );
  XOR U44258 ( .A(n35247), .B(n35246), .Z(N62256) );
  XNOR U44259 ( .A(n35264), .B(n35265), .Z(n35246) );
  XNOR U44260 ( .A(n35279), .B(n35280), .Z(n35265) );
  XOR U44261 ( .A(n35276), .B(n35275), .Z(n35280) );
  XOR U44262 ( .A(y[3084]), .B(x[3084]), .Z(n35275) );
  XOR U44263 ( .A(n35278), .B(n35277), .Z(n35276) );
  XOR U44264 ( .A(y[3086]), .B(x[3086]), .Z(n35277) );
  XOR U44265 ( .A(y[3085]), .B(x[3085]), .Z(n35278) );
  XOR U44266 ( .A(n35270), .B(n35269), .Z(n35279) );
  XOR U44267 ( .A(n35272), .B(n35271), .Z(n35269) );
  XOR U44268 ( .A(y[3083]), .B(x[3083]), .Z(n35271) );
  XOR U44269 ( .A(y[3082]), .B(x[3082]), .Z(n35272) );
  XOR U44270 ( .A(y[3081]), .B(x[3081]), .Z(n35270) );
  XNOR U44271 ( .A(n35263), .B(n35262), .Z(n35264) );
  XNOR U44272 ( .A(n35259), .B(n35258), .Z(n35262) );
  XOR U44273 ( .A(n35261), .B(n35260), .Z(n35258) );
  XOR U44274 ( .A(y[3080]), .B(x[3080]), .Z(n35260) );
  XOR U44275 ( .A(y[3079]), .B(x[3079]), .Z(n35261) );
  XOR U44276 ( .A(y[3078]), .B(x[3078]), .Z(n35259) );
  XOR U44277 ( .A(n35253), .B(n35252), .Z(n35263) );
  XOR U44278 ( .A(n35255), .B(n35254), .Z(n35252) );
  XOR U44279 ( .A(y[3077]), .B(x[3077]), .Z(n35254) );
  XOR U44280 ( .A(y[3076]), .B(x[3076]), .Z(n35255) );
  XOR U44281 ( .A(y[3075]), .B(x[3075]), .Z(n35253) );
  XNOR U44282 ( .A(n35229), .B(n35230), .Z(n35247) );
  XNOR U44283 ( .A(n35244), .B(n35245), .Z(n35230) );
  XOR U44284 ( .A(n35241), .B(n35240), .Z(n35245) );
  XOR U44285 ( .A(y[3072]), .B(x[3072]), .Z(n35240) );
  XOR U44286 ( .A(n35243), .B(n35242), .Z(n35241) );
  XOR U44287 ( .A(y[3074]), .B(x[3074]), .Z(n35242) );
  XOR U44288 ( .A(y[3073]), .B(x[3073]), .Z(n35243) );
  XOR U44289 ( .A(n35235), .B(n35234), .Z(n35244) );
  XOR U44290 ( .A(n35237), .B(n35236), .Z(n35234) );
  XOR U44291 ( .A(y[3071]), .B(x[3071]), .Z(n35236) );
  XOR U44292 ( .A(y[3070]), .B(x[3070]), .Z(n35237) );
  XOR U44293 ( .A(y[3069]), .B(x[3069]), .Z(n35235) );
  XNOR U44294 ( .A(n35228), .B(n35227), .Z(n35229) );
  XNOR U44295 ( .A(n35224), .B(n35223), .Z(n35227) );
  XOR U44296 ( .A(n35226), .B(n35225), .Z(n35223) );
  XOR U44297 ( .A(y[3068]), .B(x[3068]), .Z(n35225) );
  XOR U44298 ( .A(y[3067]), .B(x[3067]), .Z(n35226) );
  XOR U44299 ( .A(y[3066]), .B(x[3066]), .Z(n35224) );
  XOR U44300 ( .A(n35218), .B(n35217), .Z(n35228) );
  XOR U44301 ( .A(n35220), .B(n35219), .Z(n35217) );
  XOR U44302 ( .A(y[3065]), .B(x[3065]), .Z(n35219) );
  XOR U44303 ( .A(y[3064]), .B(x[3064]), .Z(n35220) );
  XOR U44304 ( .A(y[3063]), .B(x[3063]), .Z(n35218) );
  NAND U44305 ( .A(n35281), .B(n35282), .Z(N62247) );
  NAND U44306 ( .A(n35283), .B(n35284), .Z(n35282) );
  NANDN U44307 ( .A(n35285), .B(n35286), .Z(n35284) );
  NANDN U44308 ( .A(n35286), .B(n35285), .Z(n35281) );
  XOR U44309 ( .A(n35285), .B(n35287), .Z(N62246) );
  XNOR U44310 ( .A(n35283), .B(n35286), .Z(n35287) );
  NAND U44311 ( .A(n35288), .B(n35289), .Z(n35286) );
  NAND U44312 ( .A(n35290), .B(n35291), .Z(n35289) );
  NANDN U44313 ( .A(n35292), .B(n35293), .Z(n35291) );
  NANDN U44314 ( .A(n35293), .B(n35292), .Z(n35288) );
  AND U44315 ( .A(n35294), .B(n35295), .Z(n35283) );
  NAND U44316 ( .A(n35296), .B(n35297), .Z(n35295) );
  NANDN U44317 ( .A(n35298), .B(n35299), .Z(n35297) );
  NANDN U44318 ( .A(n35299), .B(n35298), .Z(n35294) );
  IV U44319 ( .A(n35300), .Z(n35299) );
  AND U44320 ( .A(n35301), .B(n35302), .Z(n35285) );
  NAND U44321 ( .A(n35303), .B(n35304), .Z(n35302) );
  NANDN U44322 ( .A(n35305), .B(n35306), .Z(n35304) );
  NANDN U44323 ( .A(n35306), .B(n35305), .Z(n35301) );
  XOR U44324 ( .A(n35298), .B(n35307), .Z(N62245) );
  XNOR U44325 ( .A(n35296), .B(n35300), .Z(n35307) );
  XOR U44326 ( .A(n35293), .B(n35308), .Z(n35300) );
  XNOR U44327 ( .A(n35290), .B(n35292), .Z(n35308) );
  AND U44328 ( .A(n35309), .B(n35310), .Z(n35292) );
  NANDN U44329 ( .A(n35311), .B(n35312), .Z(n35310) );
  OR U44330 ( .A(n35313), .B(n35314), .Z(n35312) );
  IV U44331 ( .A(n35315), .Z(n35314) );
  NANDN U44332 ( .A(n35315), .B(n35313), .Z(n35309) );
  AND U44333 ( .A(n35316), .B(n35317), .Z(n35290) );
  NAND U44334 ( .A(n35318), .B(n35319), .Z(n35317) );
  NANDN U44335 ( .A(n35320), .B(n35321), .Z(n35319) );
  NANDN U44336 ( .A(n35321), .B(n35320), .Z(n35316) );
  IV U44337 ( .A(n35322), .Z(n35321) );
  NAND U44338 ( .A(n35323), .B(n35324), .Z(n35293) );
  NANDN U44339 ( .A(n35325), .B(n35326), .Z(n35324) );
  NANDN U44340 ( .A(n35327), .B(n35328), .Z(n35326) );
  NANDN U44341 ( .A(n35328), .B(n35327), .Z(n35323) );
  IV U44342 ( .A(n35329), .Z(n35327) );
  AND U44343 ( .A(n35330), .B(n35331), .Z(n35296) );
  NAND U44344 ( .A(n35332), .B(n35333), .Z(n35331) );
  NANDN U44345 ( .A(n35334), .B(n35335), .Z(n35333) );
  NANDN U44346 ( .A(n35335), .B(n35334), .Z(n35330) );
  XOR U44347 ( .A(n35306), .B(n35336), .Z(n35298) );
  XNOR U44348 ( .A(n35303), .B(n35305), .Z(n35336) );
  AND U44349 ( .A(n35337), .B(n35338), .Z(n35305) );
  NANDN U44350 ( .A(n35339), .B(n35340), .Z(n35338) );
  OR U44351 ( .A(n35341), .B(n35342), .Z(n35340) );
  IV U44352 ( .A(n35343), .Z(n35342) );
  NANDN U44353 ( .A(n35343), .B(n35341), .Z(n35337) );
  AND U44354 ( .A(n35344), .B(n35345), .Z(n35303) );
  NAND U44355 ( .A(n35346), .B(n35347), .Z(n35345) );
  NANDN U44356 ( .A(n35348), .B(n35349), .Z(n35347) );
  NANDN U44357 ( .A(n35349), .B(n35348), .Z(n35344) );
  IV U44358 ( .A(n35350), .Z(n35349) );
  NAND U44359 ( .A(n35351), .B(n35352), .Z(n35306) );
  NANDN U44360 ( .A(n35353), .B(n35354), .Z(n35352) );
  NANDN U44361 ( .A(n35355), .B(n35356), .Z(n35354) );
  NANDN U44362 ( .A(n35356), .B(n35355), .Z(n35351) );
  IV U44363 ( .A(n35357), .Z(n35355) );
  XOR U44364 ( .A(n35332), .B(n35358), .Z(N62244) );
  XNOR U44365 ( .A(n35335), .B(n35334), .Z(n35358) );
  XNOR U44366 ( .A(n35346), .B(n35359), .Z(n35334) );
  XNOR U44367 ( .A(n35350), .B(n35348), .Z(n35359) );
  XOR U44368 ( .A(n35356), .B(n35360), .Z(n35348) );
  XNOR U44369 ( .A(n35353), .B(n35357), .Z(n35360) );
  AND U44370 ( .A(n35361), .B(n35362), .Z(n35357) );
  NAND U44371 ( .A(n35363), .B(n35364), .Z(n35362) );
  NAND U44372 ( .A(n35365), .B(n35366), .Z(n35361) );
  AND U44373 ( .A(n35367), .B(n35368), .Z(n35353) );
  NAND U44374 ( .A(n35369), .B(n35370), .Z(n35368) );
  NAND U44375 ( .A(n35371), .B(n35372), .Z(n35367) );
  NANDN U44376 ( .A(n35373), .B(n35374), .Z(n35356) );
  ANDN U44377 ( .B(n35375), .A(n35376), .Z(n35350) );
  XNOR U44378 ( .A(n35341), .B(n35377), .Z(n35346) );
  XNOR U44379 ( .A(n35339), .B(n35343), .Z(n35377) );
  AND U44380 ( .A(n35378), .B(n35379), .Z(n35343) );
  NAND U44381 ( .A(n35380), .B(n35381), .Z(n35379) );
  NAND U44382 ( .A(n35382), .B(n35383), .Z(n35378) );
  AND U44383 ( .A(n35384), .B(n35385), .Z(n35339) );
  NAND U44384 ( .A(n35386), .B(n35387), .Z(n35385) );
  NAND U44385 ( .A(n35388), .B(n35389), .Z(n35384) );
  AND U44386 ( .A(n35390), .B(n35391), .Z(n35341) );
  NAND U44387 ( .A(n35392), .B(n35393), .Z(n35335) );
  XNOR U44388 ( .A(n35318), .B(n35394), .Z(n35332) );
  XNOR U44389 ( .A(n35322), .B(n35320), .Z(n35394) );
  XOR U44390 ( .A(n35328), .B(n35395), .Z(n35320) );
  XNOR U44391 ( .A(n35325), .B(n35329), .Z(n35395) );
  AND U44392 ( .A(n35396), .B(n35397), .Z(n35329) );
  NAND U44393 ( .A(n35398), .B(n35399), .Z(n35397) );
  NAND U44394 ( .A(n35400), .B(n35401), .Z(n35396) );
  AND U44395 ( .A(n35402), .B(n35403), .Z(n35325) );
  NAND U44396 ( .A(n35404), .B(n35405), .Z(n35403) );
  NAND U44397 ( .A(n35406), .B(n35407), .Z(n35402) );
  NANDN U44398 ( .A(n35408), .B(n35409), .Z(n35328) );
  ANDN U44399 ( .B(n35410), .A(n35411), .Z(n35322) );
  XNOR U44400 ( .A(n35313), .B(n35412), .Z(n35318) );
  XNOR U44401 ( .A(n35311), .B(n35315), .Z(n35412) );
  AND U44402 ( .A(n35413), .B(n35414), .Z(n35315) );
  NAND U44403 ( .A(n35415), .B(n35416), .Z(n35414) );
  NAND U44404 ( .A(n35417), .B(n35418), .Z(n35413) );
  AND U44405 ( .A(n35419), .B(n35420), .Z(n35311) );
  NAND U44406 ( .A(n35421), .B(n35422), .Z(n35420) );
  NAND U44407 ( .A(n35423), .B(n35424), .Z(n35419) );
  AND U44408 ( .A(n35425), .B(n35426), .Z(n35313) );
  XOR U44409 ( .A(n35393), .B(n35392), .Z(N62243) );
  XNOR U44410 ( .A(n35410), .B(n35411), .Z(n35392) );
  XNOR U44411 ( .A(n35425), .B(n35426), .Z(n35411) );
  XOR U44412 ( .A(n35422), .B(n35421), .Z(n35426) );
  XOR U44413 ( .A(y[3060]), .B(x[3060]), .Z(n35421) );
  XOR U44414 ( .A(n35424), .B(n35423), .Z(n35422) );
  XOR U44415 ( .A(y[3062]), .B(x[3062]), .Z(n35423) );
  XOR U44416 ( .A(y[3061]), .B(x[3061]), .Z(n35424) );
  XOR U44417 ( .A(n35416), .B(n35415), .Z(n35425) );
  XOR U44418 ( .A(n35418), .B(n35417), .Z(n35415) );
  XOR U44419 ( .A(y[3059]), .B(x[3059]), .Z(n35417) );
  XOR U44420 ( .A(y[3058]), .B(x[3058]), .Z(n35418) );
  XOR U44421 ( .A(y[3057]), .B(x[3057]), .Z(n35416) );
  XNOR U44422 ( .A(n35409), .B(n35408), .Z(n35410) );
  XNOR U44423 ( .A(n35405), .B(n35404), .Z(n35408) );
  XOR U44424 ( .A(n35407), .B(n35406), .Z(n35404) );
  XOR U44425 ( .A(y[3056]), .B(x[3056]), .Z(n35406) );
  XOR U44426 ( .A(y[3055]), .B(x[3055]), .Z(n35407) );
  XOR U44427 ( .A(y[3054]), .B(x[3054]), .Z(n35405) );
  XOR U44428 ( .A(n35399), .B(n35398), .Z(n35409) );
  XOR U44429 ( .A(n35401), .B(n35400), .Z(n35398) );
  XOR U44430 ( .A(y[3053]), .B(x[3053]), .Z(n35400) );
  XOR U44431 ( .A(y[3052]), .B(x[3052]), .Z(n35401) );
  XOR U44432 ( .A(y[3051]), .B(x[3051]), .Z(n35399) );
  XNOR U44433 ( .A(n35375), .B(n35376), .Z(n35393) );
  XNOR U44434 ( .A(n35390), .B(n35391), .Z(n35376) );
  XOR U44435 ( .A(n35387), .B(n35386), .Z(n35391) );
  XOR U44436 ( .A(y[3048]), .B(x[3048]), .Z(n35386) );
  XOR U44437 ( .A(n35389), .B(n35388), .Z(n35387) );
  XOR U44438 ( .A(y[3050]), .B(x[3050]), .Z(n35388) );
  XOR U44439 ( .A(y[3049]), .B(x[3049]), .Z(n35389) );
  XOR U44440 ( .A(n35381), .B(n35380), .Z(n35390) );
  XOR U44441 ( .A(n35383), .B(n35382), .Z(n35380) );
  XOR U44442 ( .A(y[3047]), .B(x[3047]), .Z(n35382) );
  XOR U44443 ( .A(y[3046]), .B(x[3046]), .Z(n35383) );
  XOR U44444 ( .A(y[3045]), .B(x[3045]), .Z(n35381) );
  XNOR U44445 ( .A(n35374), .B(n35373), .Z(n35375) );
  XNOR U44446 ( .A(n35370), .B(n35369), .Z(n35373) );
  XOR U44447 ( .A(n35372), .B(n35371), .Z(n35369) );
  XOR U44448 ( .A(y[3044]), .B(x[3044]), .Z(n35371) );
  XOR U44449 ( .A(y[3043]), .B(x[3043]), .Z(n35372) );
  XOR U44450 ( .A(y[3042]), .B(x[3042]), .Z(n35370) );
  XOR U44451 ( .A(n35364), .B(n35363), .Z(n35374) );
  XOR U44452 ( .A(n35366), .B(n35365), .Z(n35363) );
  XOR U44453 ( .A(y[3041]), .B(x[3041]), .Z(n35365) );
  XOR U44454 ( .A(y[3040]), .B(x[3040]), .Z(n35366) );
  XOR U44455 ( .A(y[3039]), .B(x[3039]), .Z(n35364) );
  NAND U44456 ( .A(n35427), .B(n35428), .Z(N62234) );
  NAND U44457 ( .A(n35429), .B(n35430), .Z(n35428) );
  NANDN U44458 ( .A(n35431), .B(n35432), .Z(n35430) );
  NANDN U44459 ( .A(n35432), .B(n35431), .Z(n35427) );
  XOR U44460 ( .A(n35431), .B(n35433), .Z(N62233) );
  XNOR U44461 ( .A(n35429), .B(n35432), .Z(n35433) );
  NAND U44462 ( .A(n35434), .B(n35435), .Z(n35432) );
  NAND U44463 ( .A(n35436), .B(n35437), .Z(n35435) );
  NANDN U44464 ( .A(n35438), .B(n35439), .Z(n35437) );
  NANDN U44465 ( .A(n35439), .B(n35438), .Z(n35434) );
  AND U44466 ( .A(n35440), .B(n35441), .Z(n35429) );
  NAND U44467 ( .A(n35442), .B(n35443), .Z(n35441) );
  NANDN U44468 ( .A(n35444), .B(n35445), .Z(n35443) );
  NANDN U44469 ( .A(n35445), .B(n35444), .Z(n35440) );
  IV U44470 ( .A(n35446), .Z(n35445) );
  AND U44471 ( .A(n35447), .B(n35448), .Z(n35431) );
  NAND U44472 ( .A(n35449), .B(n35450), .Z(n35448) );
  NANDN U44473 ( .A(n35451), .B(n35452), .Z(n35450) );
  NANDN U44474 ( .A(n35452), .B(n35451), .Z(n35447) );
  XOR U44475 ( .A(n35444), .B(n35453), .Z(N62232) );
  XNOR U44476 ( .A(n35442), .B(n35446), .Z(n35453) );
  XOR U44477 ( .A(n35439), .B(n35454), .Z(n35446) );
  XNOR U44478 ( .A(n35436), .B(n35438), .Z(n35454) );
  AND U44479 ( .A(n35455), .B(n35456), .Z(n35438) );
  NANDN U44480 ( .A(n35457), .B(n35458), .Z(n35456) );
  OR U44481 ( .A(n35459), .B(n35460), .Z(n35458) );
  IV U44482 ( .A(n35461), .Z(n35460) );
  NANDN U44483 ( .A(n35461), .B(n35459), .Z(n35455) );
  AND U44484 ( .A(n35462), .B(n35463), .Z(n35436) );
  NAND U44485 ( .A(n35464), .B(n35465), .Z(n35463) );
  NANDN U44486 ( .A(n35466), .B(n35467), .Z(n35465) );
  NANDN U44487 ( .A(n35467), .B(n35466), .Z(n35462) );
  IV U44488 ( .A(n35468), .Z(n35467) );
  NAND U44489 ( .A(n35469), .B(n35470), .Z(n35439) );
  NANDN U44490 ( .A(n35471), .B(n35472), .Z(n35470) );
  NANDN U44491 ( .A(n35473), .B(n35474), .Z(n35472) );
  NANDN U44492 ( .A(n35474), .B(n35473), .Z(n35469) );
  IV U44493 ( .A(n35475), .Z(n35473) );
  AND U44494 ( .A(n35476), .B(n35477), .Z(n35442) );
  NAND U44495 ( .A(n35478), .B(n35479), .Z(n35477) );
  NANDN U44496 ( .A(n35480), .B(n35481), .Z(n35479) );
  NANDN U44497 ( .A(n35481), .B(n35480), .Z(n35476) );
  XOR U44498 ( .A(n35452), .B(n35482), .Z(n35444) );
  XNOR U44499 ( .A(n35449), .B(n35451), .Z(n35482) );
  AND U44500 ( .A(n35483), .B(n35484), .Z(n35451) );
  NANDN U44501 ( .A(n35485), .B(n35486), .Z(n35484) );
  OR U44502 ( .A(n35487), .B(n35488), .Z(n35486) );
  IV U44503 ( .A(n35489), .Z(n35488) );
  NANDN U44504 ( .A(n35489), .B(n35487), .Z(n35483) );
  AND U44505 ( .A(n35490), .B(n35491), .Z(n35449) );
  NAND U44506 ( .A(n35492), .B(n35493), .Z(n35491) );
  NANDN U44507 ( .A(n35494), .B(n35495), .Z(n35493) );
  NANDN U44508 ( .A(n35495), .B(n35494), .Z(n35490) );
  IV U44509 ( .A(n35496), .Z(n35495) );
  NAND U44510 ( .A(n35497), .B(n35498), .Z(n35452) );
  NANDN U44511 ( .A(n35499), .B(n35500), .Z(n35498) );
  NANDN U44512 ( .A(n35501), .B(n35502), .Z(n35500) );
  NANDN U44513 ( .A(n35502), .B(n35501), .Z(n35497) );
  IV U44514 ( .A(n35503), .Z(n35501) );
  XOR U44515 ( .A(n35478), .B(n35504), .Z(N62231) );
  XNOR U44516 ( .A(n35481), .B(n35480), .Z(n35504) );
  XNOR U44517 ( .A(n35492), .B(n35505), .Z(n35480) );
  XNOR U44518 ( .A(n35496), .B(n35494), .Z(n35505) );
  XOR U44519 ( .A(n35502), .B(n35506), .Z(n35494) );
  XNOR U44520 ( .A(n35499), .B(n35503), .Z(n35506) );
  AND U44521 ( .A(n35507), .B(n35508), .Z(n35503) );
  NAND U44522 ( .A(n35509), .B(n35510), .Z(n35508) );
  NAND U44523 ( .A(n35511), .B(n35512), .Z(n35507) );
  AND U44524 ( .A(n35513), .B(n35514), .Z(n35499) );
  NAND U44525 ( .A(n35515), .B(n35516), .Z(n35514) );
  NAND U44526 ( .A(n35517), .B(n35518), .Z(n35513) );
  NANDN U44527 ( .A(n35519), .B(n35520), .Z(n35502) );
  ANDN U44528 ( .B(n35521), .A(n35522), .Z(n35496) );
  XNOR U44529 ( .A(n35487), .B(n35523), .Z(n35492) );
  XNOR U44530 ( .A(n35485), .B(n35489), .Z(n35523) );
  AND U44531 ( .A(n35524), .B(n35525), .Z(n35489) );
  NAND U44532 ( .A(n35526), .B(n35527), .Z(n35525) );
  NAND U44533 ( .A(n35528), .B(n35529), .Z(n35524) );
  AND U44534 ( .A(n35530), .B(n35531), .Z(n35485) );
  NAND U44535 ( .A(n35532), .B(n35533), .Z(n35531) );
  NAND U44536 ( .A(n35534), .B(n35535), .Z(n35530) );
  AND U44537 ( .A(n35536), .B(n35537), .Z(n35487) );
  NAND U44538 ( .A(n35538), .B(n35539), .Z(n35481) );
  XNOR U44539 ( .A(n35464), .B(n35540), .Z(n35478) );
  XNOR U44540 ( .A(n35468), .B(n35466), .Z(n35540) );
  XOR U44541 ( .A(n35474), .B(n35541), .Z(n35466) );
  XNOR U44542 ( .A(n35471), .B(n35475), .Z(n35541) );
  AND U44543 ( .A(n35542), .B(n35543), .Z(n35475) );
  NAND U44544 ( .A(n35544), .B(n35545), .Z(n35543) );
  NAND U44545 ( .A(n35546), .B(n35547), .Z(n35542) );
  AND U44546 ( .A(n35548), .B(n35549), .Z(n35471) );
  NAND U44547 ( .A(n35550), .B(n35551), .Z(n35549) );
  NAND U44548 ( .A(n35552), .B(n35553), .Z(n35548) );
  NANDN U44549 ( .A(n35554), .B(n35555), .Z(n35474) );
  ANDN U44550 ( .B(n35556), .A(n35557), .Z(n35468) );
  XNOR U44551 ( .A(n35459), .B(n35558), .Z(n35464) );
  XNOR U44552 ( .A(n35457), .B(n35461), .Z(n35558) );
  AND U44553 ( .A(n35559), .B(n35560), .Z(n35461) );
  NAND U44554 ( .A(n35561), .B(n35562), .Z(n35560) );
  NAND U44555 ( .A(n35563), .B(n35564), .Z(n35559) );
  AND U44556 ( .A(n35565), .B(n35566), .Z(n35457) );
  NAND U44557 ( .A(n35567), .B(n35568), .Z(n35566) );
  NAND U44558 ( .A(n35569), .B(n35570), .Z(n35565) );
  AND U44559 ( .A(n35571), .B(n35572), .Z(n35459) );
  XOR U44560 ( .A(n35539), .B(n35538), .Z(N62230) );
  XNOR U44561 ( .A(n35556), .B(n35557), .Z(n35538) );
  XNOR U44562 ( .A(n35571), .B(n35572), .Z(n35557) );
  XOR U44563 ( .A(n35568), .B(n35567), .Z(n35572) );
  XOR U44564 ( .A(y[3036]), .B(x[3036]), .Z(n35567) );
  XOR U44565 ( .A(n35570), .B(n35569), .Z(n35568) );
  XOR U44566 ( .A(y[3038]), .B(x[3038]), .Z(n35569) );
  XOR U44567 ( .A(y[3037]), .B(x[3037]), .Z(n35570) );
  XOR U44568 ( .A(n35562), .B(n35561), .Z(n35571) );
  XOR U44569 ( .A(n35564), .B(n35563), .Z(n35561) );
  XOR U44570 ( .A(y[3035]), .B(x[3035]), .Z(n35563) );
  XOR U44571 ( .A(y[3034]), .B(x[3034]), .Z(n35564) );
  XOR U44572 ( .A(y[3033]), .B(x[3033]), .Z(n35562) );
  XNOR U44573 ( .A(n35555), .B(n35554), .Z(n35556) );
  XNOR U44574 ( .A(n35551), .B(n35550), .Z(n35554) );
  XOR U44575 ( .A(n35553), .B(n35552), .Z(n35550) );
  XOR U44576 ( .A(y[3032]), .B(x[3032]), .Z(n35552) );
  XOR U44577 ( .A(y[3031]), .B(x[3031]), .Z(n35553) );
  XOR U44578 ( .A(y[3030]), .B(x[3030]), .Z(n35551) );
  XOR U44579 ( .A(n35545), .B(n35544), .Z(n35555) );
  XOR U44580 ( .A(n35547), .B(n35546), .Z(n35544) );
  XOR U44581 ( .A(y[3029]), .B(x[3029]), .Z(n35546) );
  XOR U44582 ( .A(y[3028]), .B(x[3028]), .Z(n35547) );
  XOR U44583 ( .A(y[3027]), .B(x[3027]), .Z(n35545) );
  XNOR U44584 ( .A(n35521), .B(n35522), .Z(n35539) );
  XNOR U44585 ( .A(n35536), .B(n35537), .Z(n35522) );
  XOR U44586 ( .A(n35533), .B(n35532), .Z(n35537) );
  XOR U44587 ( .A(y[3024]), .B(x[3024]), .Z(n35532) );
  XOR U44588 ( .A(n35535), .B(n35534), .Z(n35533) );
  XOR U44589 ( .A(y[3026]), .B(x[3026]), .Z(n35534) );
  XOR U44590 ( .A(y[3025]), .B(x[3025]), .Z(n35535) );
  XOR U44591 ( .A(n35527), .B(n35526), .Z(n35536) );
  XOR U44592 ( .A(n35529), .B(n35528), .Z(n35526) );
  XOR U44593 ( .A(y[3023]), .B(x[3023]), .Z(n35528) );
  XOR U44594 ( .A(y[3022]), .B(x[3022]), .Z(n35529) );
  XOR U44595 ( .A(y[3021]), .B(x[3021]), .Z(n35527) );
  XNOR U44596 ( .A(n35520), .B(n35519), .Z(n35521) );
  XNOR U44597 ( .A(n35516), .B(n35515), .Z(n35519) );
  XOR U44598 ( .A(n35518), .B(n35517), .Z(n35515) );
  XOR U44599 ( .A(y[3020]), .B(x[3020]), .Z(n35517) );
  XOR U44600 ( .A(y[3019]), .B(x[3019]), .Z(n35518) );
  XOR U44601 ( .A(y[3018]), .B(x[3018]), .Z(n35516) );
  XOR U44602 ( .A(n35510), .B(n35509), .Z(n35520) );
  XOR U44603 ( .A(n35512), .B(n35511), .Z(n35509) );
  XOR U44604 ( .A(y[3017]), .B(x[3017]), .Z(n35511) );
  XOR U44605 ( .A(y[3016]), .B(x[3016]), .Z(n35512) );
  XOR U44606 ( .A(y[3015]), .B(x[3015]), .Z(n35510) );
  NAND U44607 ( .A(n35573), .B(n35574), .Z(N62221) );
  NAND U44608 ( .A(n35575), .B(n35576), .Z(n35574) );
  NANDN U44609 ( .A(n35577), .B(n35578), .Z(n35576) );
  NANDN U44610 ( .A(n35578), .B(n35577), .Z(n35573) );
  XOR U44611 ( .A(n35577), .B(n35579), .Z(N62220) );
  XNOR U44612 ( .A(n35575), .B(n35578), .Z(n35579) );
  NAND U44613 ( .A(n35580), .B(n35581), .Z(n35578) );
  NAND U44614 ( .A(n35582), .B(n35583), .Z(n35581) );
  NANDN U44615 ( .A(n35584), .B(n35585), .Z(n35583) );
  NANDN U44616 ( .A(n35585), .B(n35584), .Z(n35580) );
  AND U44617 ( .A(n35586), .B(n35587), .Z(n35575) );
  NAND U44618 ( .A(n35588), .B(n35589), .Z(n35587) );
  NANDN U44619 ( .A(n35590), .B(n35591), .Z(n35589) );
  NANDN U44620 ( .A(n35591), .B(n35590), .Z(n35586) );
  IV U44621 ( .A(n35592), .Z(n35591) );
  AND U44622 ( .A(n35593), .B(n35594), .Z(n35577) );
  NAND U44623 ( .A(n35595), .B(n35596), .Z(n35594) );
  NANDN U44624 ( .A(n35597), .B(n35598), .Z(n35596) );
  NANDN U44625 ( .A(n35598), .B(n35597), .Z(n35593) );
  XOR U44626 ( .A(n35590), .B(n35599), .Z(N62219) );
  XNOR U44627 ( .A(n35588), .B(n35592), .Z(n35599) );
  XOR U44628 ( .A(n35585), .B(n35600), .Z(n35592) );
  XNOR U44629 ( .A(n35582), .B(n35584), .Z(n35600) );
  AND U44630 ( .A(n35601), .B(n35602), .Z(n35584) );
  NANDN U44631 ( .A(n35603), .B(n35604), .Z(n35602) );
  OR U44632 ( .A(n35605), .B(n35606), .Z(n35604) );
  IV U44633 ( .A(n35607), .Z(n35606) );
  NANDN U44634 ( .A(n35607), .B(n35605), .Z(n35601) );
  AND U44635 ( .A(n35608), .B(n35609), .Z(n35582) );
  NAND U44636 ( .A(n35610), .B(n35611), .Z(n35609) );
  NANDN U44637 ( .A(n35612), .B(n35613), .Z(n35611) );
  NANDN U44638 ( .A(n35613), .B(n35612), .Z(n35608) );
  IV U44639 ( .A(n35614), .Z(n35613) );
  NAND U44640 ( .A(n35615), .B(n35616), .Z(n35585) );
  NANDN U44641 ( .A(n35617), .B(n35618), .Z(n35616) );
  NANDN U44642 ( .A(n35619), .B(n35620), .Z(n35618) );
  NANDN U44643 ( .A(n35620), .B(n35619), .Z(n35615) );
  IV U44644 ( .A(n35621), .Z(n35619) );
  AND U44645 ( .A(n35622), .B(n35623), .Z(n35588) );
  NAND U44646 ( .A(n35624), .B(n35625), .Z(n35623) );
  NANDN U44647 ( .A(n35626), .B(n35627), .Z(n35625) );
  NANDN U44648 ( .A(n35627), .B(n35626), .Z(n35622) );
  XOR U44649 ( .A(n35598), .B(n35628), .Z(n35590) );
  XNOR U44650 ( .A(n35595), .B(n35597), .Z(n35628) );
  AND U44651 ( .A(n35629), .B(n35630), .Z(n35597) );
  NANDN U44652 ( .A(n35631), .B(n35632), .Z(n35630) );
  OR U44653 ( .A(n35633), .B(n35634), .Z(n35632) );
  IV U44654 ( .A(n35635), .Z(n35634) );
  NANDN U44655 ( .A(n35635), .B(n35633), .Z(n35629) );
  AND U44656 ( .A(n35636), .B(n35637), .Z(n35595) );
  NAND U44657 ( .A(n35638), .B(n35639), .Z(n35637) );
  NANDN U44658 ( .A(n35640), .B(n35641), .Z(n35639) );
  NANDN U44659 ( .A(n35641), .B(n35640), .Z(n35636) );
  IV U44660 ( .A(n35642), .Z(n35641) );
  NAND U44661 ( .A(n35643), .B(n35644), .Z(n35598) );
  NANDN U44662 ( .A(n35645), .B(n35646), .Z(n35644) );
  NANDN U44663 ( .A(n35647), .B(n35648), .Z(n35646) );
  NANDN U44664 ( .A(n35648), .B(n35647), .Z(n35643) );
  IV U44665 ( .A(n35649), .Z(n35647) );
  XOR U44666 ( .A(n35624), .B(n35650), .Z(N62218) );
  XNOR U44667 ( .A(n35627), .B(n35626), .Z(n35650) );
  XNOR U44668 ( .A(n35638), .B(n35651), .Z(n35626) );
  XNOR U44669 ( .A(n35642), .B(n35640), .Z(n35651) );
  XOR U44670 ( .A(n35648), .B(n35652), .Z(n35640) );
  XNOR U44671 ( .A(n35645), .B(n35649), .Z(n35652) );
  AND U44672 ( .A(n35653), .B(n35654), .Z(n35649) );
  NAND U44673 ( .A(n35655), .B(n35656), .Z(n35654) );
  NAND U44674 ( .A(n35657), .B(n35658), .Z(n35653) );
  AND U44675 ( .A(n35659), .B(n35660), .Z(n35645) );
  NAND U44676 ( .A(n35661), .B(n35662), .Z(n35660) );
  NAND U44677 ( .A(n35663), .B(n35664), .Z(n35659) );
  NANDN U44678 ( .A(n35665), .B(n35666), .Z(n35648) );
  ANDN U44679 ( .B(n35667), .A(n35668), .Z(n35642) );
  XNOR U44680 ( .A(n35633), .B(n35669), .Z(n35638) );
  XNOR U44681 ( .A(n35631), .B(n35635), .Z(n35669) );
  AND U44682 ( .A(n35670), .B(n35671), .Z(n35635) );
  NAND U44683 ( .A(n35672), .B(n35673), .Z(n35671) );
  NAND U44684 ( .A(n35674), .B(n35675), .Z(n35670) );
  AND U44685 ( .A(n35676), .B(n35677), .Z(n35631) );
  NAND U44686 ( .A(n35678), .B(n35679), .Z(n35677) );
  NAND U44687 ( .A(n35680), .B(n35681), .Z(n35676) );
  AND U44688 ( .A(n35682), .B(n35683), .Z(n35633) );
  NAND U44689 ( .A(n35684), .B(n35685), .Z(n35627) );
  XNOR U44690 ( .A(n35610), .B(n35686), .Z(n35624) );
  XNOR U44691 ( .A(n35614), .B(n35612), .Z(n35686) );
  XOR U44692 ( .A(n35620), .B(n35687), .Z(n35612) );
  XNOR U44693 ( .A(n35617), .B(n35621), .Z(n35687) );
  AND U44694 ( .A(n35688), .B(n35689), .Z(n35621) );
  NAND U44695 ( .A(n35690), .B(n35691), .Z(n35689) );
  NAND U44696 ( .A(n35692), .B(n35693), .Z(n35688) );
  AND U44697 ( .A(n35694), .B(n35695), .Z(n35617) );
  NAND U44698 ( .A(n35696), .B(n35697), .Z(n35695) );
  NAND U44699 ( .A(n35698), .B(n35699), .Z(n35694) );
  NANDN U44700 ( .A(n35700), .B(n35701), .Z(n35620) );
  ANDN U44701 ( .B(n35702), .A(n35703), .Z(n35614) );
  XNOR U44702 ( .A(n35605), .B(n35704), .Z(n35610) );
  XNOR U44703 ( .A(n35603), .B(n35607), .Z(n35704) );
  AND U44704 ( .A(n35705), .B(n35706), .Z(n35607) );
  NAND U44705 ( .A(n35707), .B(n35708), .Z(n35706) );
  NAND U44706 ( .A(n35709), .B(n35710), .Z(n35705) );
  AND U44707 ( .A(n35711), .B(n35712), .Z(n35603) );
  NAND U44708 ( .A(n35713), .B(n35714), .Z(n35712) );
  NAND U44709 ( .A(n35715), .B(n35716), .Z(n35711) );
  AND U44710 ( .A(n35717), .B(n35718), .Z(n35605) );
  XOR U44711 ( .A(n35685), .B(n35684), .Z(N62217) );
  XNOR U44712 ( .A(n35702), .B(n35703), .Z(n35684) );
  XNOR U44713 ( .A(n35717), .B(n35718), .Z(n35703) );
  XOR U44714 ( .A(n35714), .B(n35713), .Z(n35718) );
  XOR U44715 ( .A(y[3012]), .B(x[3012]), .Z(n35713) );
  XOR U44716 ( .A(n35716), .B(n35715), .Z(n35714) );
  XOR U44717 ( .A(y[3014]), .B(x[3014]), .Z(n35715) );
  XOR U44718 ( .A(y[3013]), .B(x[3013]), .Z(n35716) );
  XOR U44719 ( .A(n35708), .B(n35707), .Z(n35717) );
  XOR U44720 ( .A(n35710), .B(n35709), .Z(n35707) );
  XOR U44721 ( .A(y[3011]), .B(x[3011]), .Z(n35709) );
  XOR U44722 ( .A(y[3010]), .B(x[3010]), .Z(n35710) );
  XOR U44723 ( .A(y[3009]), .B(x[3009]), .Z(n35708) );
  XNOR U44724 ( .A(n35701), .B(n35700), .Z(n35702) );
  XNOR U44725 ( .A(n35697), .B(n35696), .Z(n35700) );
  XOR U44726 ( .A(n35699), .B(n35698), .Z(n35696) );
  XOR U44727 ( .A(y[3008]), .B(x[3008]), .Z(n35698) );
  XOR U44728 ( .A(y[3007]), .B(x[3007]), .Z(n35699) );
  XOR U44729 ( .A(y[3006]), .B(x[3006]), .Z(n35697) );
  XOR U44730 ( .A(n35691), .B(n35690), .Z(n35701) );
  XOR U44731 ( .A(n35693), .B(n35692), .Z(n35690) );
  XOR U44732 ( .A(y[3005]), .B(x[3005]), .Z(n35692) );
  XOR U44733 ( .A(y[3004]), .B(x[3004]), .Z(n35693) );
  XOR U44734 ( .A(y[3003]), .B(x[3003]), .Z(n35691) );
  XNOR U44735 ( .A(n35667), .B(n35668), .Z(n35685) );
  XNOR U44736 ( .A(n35682), .B(n35683), .Z(n35668) );
  XOR U44737 ( .A(n35679), .B(n35678), .Z(n35683) );
  XOR U44738 ( .A(y[3000]), .B(x[3000]), .Z(n35678) );
  XOR U44739 ( .A(n35681), .B(n35680), .Z(n35679) );
  XOR U44740 ( .A(y[3002]), .B(x[3002]), .Z(n35680) );
  XOR U44741 ( .A(y[3001]), .B(x[3001]), .Z(n35681) );
  XOR U44742 ( .A(n35673), .B(n35672), .Z(n35682) );
  XOR U44743 ( .A(n35675), .B(n35674), .Z(n35672) );
  XOR U44744 ( .A(y[2999]), .B(x[2999]), .Z(n35674) );
  XOR U44745 ( .A(y[2998]), .B(x[2998]), .Z(n35675) );
  XOR U44746 ( .A(y[2997]), .B(x[2997]), .Z(n35673) );
  XNOR U44747 ( .A(n35666), .B(n35665), .Z(n35667) );
  XNOR U44748 ( .A(n35662), .B(n35661), .Z(n35665) );
  XOR U44749 ( .A(n35664), .B(n35663), .Z(n35661) );
  XOR U44750 ( .A(y[2996]), .B(x[2996]), .Z(n35663) );
  XOR U44751 ( .A(y[2995]), .B(x[2995]), .Z(n35664) );
  XOR U44752 ( .A(y[2994]), .B(x[2994]), .Z(n35662) );
  XOR U44753 ( .A(n35656), .B(n35655), .Z(n35666) );
  XOR U44754 ( .A(n35658), .B(n35657), .Z(n35655) );
  XOR U44755 ( .A(y[2993]), .B(x[2993]), .Z(n35657) );
  XOR U44756 ( .A(y[2992]), .B(x[2992]), .Z(n35658) );
  XOR U44757 ( .A(y[2991]), .B(x[2991]), .Z(n35656) );
  NAND U44758 ( .A(n35719), .B(n35720), .Z(N62208) );
  NAND U44759 ( .A(n35721), .B(n35722), .Z(n35720) );
  NANDN U44760 ( .A(n35723), .B(n35724), .Z(n35722) );
  NANDN U44761 ( .A(n35724), .B(n35723), .Z(n35719) );
  XOR U44762 ( .A(n35723), .B(n35725), .Z(N62207) );
  XNOR U44763 ( .A(n35721), .B(n35724), .Z(n35725) );
  NAND U44764 ( .A(n35726), .B(n35727), .Z(n35724) );
  NAND U44765 ( .A(n35728), .B(n35729), .Z(n35727) );
  NANDN U44766 ( .A(n35730), .B(n35731), .Z(n35729) );
  NANDN U44767 ( .A(n35731), .B(n35730), .Z(n35726) );
  AND U44768 ( .A(n35732), .B(n35733), .Z(n35721) );
  NAND U44769 ( .A(n35734), .B(n35735), .Z(n35733) );
  NANDN U44770 ( .A(n35736), .B(n35737), .Z(n35735) );
  NANDN U44771 ( .A(n35737), .B(n35736), .Z(n35732) );
  IV U44772 ( .A(n35738), .Z(n35737) );
  AND U44773 ( .A(n35739), .B(n35740), .Z(n35723) );
  NAND U44774 ( .A(n35741), .B(n35742), .Z(n35740) );
  NANDN U44775 ( .A(n35743), .B(n35744), .Z(n35742) );
  NANDN U44776 ( .A(n35744), .B(n35743), .Z(n35739) );
  XOR U44777 ( .A(n35736), .B(n35745), .Z(N62206) );
  XNOR U44778 ( .A(n35734), .B(n35738), .Z(n35745) );
  XOR U44779 ( .A(n35731), .B(n35746), .Z(n35738) );
  XNOR U44780 ( .A(n35728), .B(n35730), .Z(n35746) );
  AND U44781 ( .A(n35747), .B(n35748), .Z(n35730) );
  NANDN U44782 ( .A(n35749), .B(n35750), .Z(n35748) );
  OR U44783 ( .A(n35751), .B(n35752), .Z(n35750) );
  IV U44784 ( .A(n35753), .Z(n35752) );
  NANDN U44785 ( .A(n35753), .B(n35751), .Z(n35747) );
  AND U44786 ( .A(n35754), .B(n35755), .Z(n35728) );
  NAND U44787 ( .A(n35756), .B(n35757), .Z(n35755) );
  NANDN U44788 ( .A(n35758), .B(n35759), .Z(n35757) );
  NANDN U44789 ( .A(n35759), .B(n35758), .Z(n35754) );
  IV U44790 ( .A(n35760), .Z(n35759) );
  NAND U44791 ( .A(n35761), .B(n35762), .Z(n35731) );
  NANDN U44792 ( .A(n35763), .B(n35764), .Z(n35762) );
  NANDN U44793 ( .A(n35765), .B(n35766), .Z(n35764) );
  NANDN U44794 ( .A(n35766), .B(n35765), .Z(n35761) );
  IV U44795 ( .A(n35767), .Z(n35765) );
  AND U44796 ( .A(n35768), .B(n35769), .Z(n35734) );
  NAND U44797 ( .A(n35770), .B(n35771), .Z(n35769) );
  NANDN U44798 ( .A(n35772), .B(n35773), .Z(n35771) );
  NANDN U44799 ( .A(n35773), .B(n35772), .Z(n35768) );
  XOR U44800 ( .A(n35744), .B(n35774), .Z(n35736) );
  XNOR U44801 ( .A(n35741), .B(n35743), .Z(n35774) );
  AND U44802 ( .A(n35775), .B(n35776), .Z(n35743) );
  NANDN U44803 ( .A(n35777), .B(n35778), .Z(n35776) );
  OR U44804 ( .A(n35779), .B(n35780), .Z(n35778) );
  IV U44805 ( .A(n35781), .Z(n35780) );
  NANDN U44806 ( .A(n35781), .B(n35779), .Z(n35775) );
  AND U44807 ( .A(n35782), .B(n35783), .Z(n35741) );
  NAND U44808 ( .A(n35784), .B(n35785), .Z(n35783) );
  NANDN U44809 ( .A(n35786), .B(n35787), .Z(n35785) );
  NANDN U44810 ( .A(n35787), .B(n35786), .Z(n35782) );
  IV U44811 ( .A(n35788), .Z(n35787) );
  NAND U44812 ( .A(n35789), .B(n35790), .Z(n35744) );
  NANDN U44813 ( .A(n35791), .B(n35792), .Z(n35790) );
  NANDN U44814 ( .A(n35793), .B(n35794), .Z(n35792) );
  NANDN U44815 ( .A(n35794), .B(n35793), .Z(n35789) );
  IV U44816 ( .A(n35795), .Z(n35793) );
  XOR U44817 ( .A(n35770), .B(n35796), .Z(N62205) );
  XNOR U44818 ( .A(n35773), .B(n35772), .Z(n35796) );
  XNOR U44819 ( .A(n35784), .B(n35797), .Z(n35772) );
  XNOR U44820 ( .A(n35788), .B(n35786), .Z(n35797) );
  XOR U44821 ( .A(n35794), .B(n35798), .Z(n35786) );
  XNOR U44822 ( .A(n35791), .B(n35795), .Z(n35798) );
  AND U44823 ( .A(n35799), .B(n35800), .Z(n35795) );
  NAND U44824 ( .A(n35801), .B(n35802), .Z(n35800) );
  NAND U44825 ( .A(n35803), .B(n35804), .Z(n35799) );
  AND U44826 ( .A(n35805), .B(n35806), .Z(n35791) );
  NAND U44827 ( .A(n35807), .B(n35808), .Z(n35806) );
  NAND U44828 ( .A(n35809), .B(n35810), .Z(n35805) );
  NANDN U44829 ( .A(n35811), .B(n35812), .Z(n35794) );
  ANDN U44830 ( .B(n35813), .A(n35814), .Z(n35788) );
  XNOR U44831 ( .A(n35779), .B(n35815), .Z(n35784) );
  XNOR U44832 ( .A(n35777), .B(n35781), .Z(n35815) );
  AND U44833 ( .A(n35816), .B(n35817), .Z(n35781) );
  NAND U44834 ( .A(n35818), .B(n35819), .Z(n35817) );
  NAND U44835 ( .A(n35820), .B(n35821), .Z(n35816) );
  AND U44836 ( .A(n35822), .B(n35823), .Z(n35777) );
  NAND U44837 ( .A(n35824), .B(n35825), .Z(n35823) );
  NAND U44838 ( .A(n35826), .B(n35827), .Z(n35822) );
  AND U44839 ( .A(n35828), .B(n35829), .Z(n35779) );
  NAND U44840 ( .A(n35830), .B(n35831), .Z(n35773) );
  XNOR U44841 ( .A(n35756), .B(n35832), .Z(n35770) );
  XNOR U44842 ( .A(n35760), .B(n35758), .Z(n35832) );
  XOR U44843 ( .A(n35766), .B(n35833), .Z(n35758) );
  XNOR U44844 ( .A(n35763), .B(n35767), .Z(n35833) );
  AND U44845 ( .A(n35834), .B(n35835), .Z(n35767) );
  NAND U44846 ( .A(n35836), .B(n35837), .Z(n35835) );
  NAND U44847 ( .A(n35838), .B(n35839), .Z(n35834) );
  AND U44848 ( .A(n35840), .B(n35841), .Z(n35763) );
  NAND U44849 ( .A(n35842), .B(n35843), .Z(n35841) );
  NAND U44850 ( .A(n35844), .B(n35845), .Z(n35840) );
  NANDN U44851 ( .A(n35846), .B(n35847), .Z(n35766) );
  ANDN U44852 ( .B(n35848), .A(n35849), .Z(n35760) );
  XNOR U44853 ( .A(n35751), .B(n35850), .Z(n35756) );
  XNOR U44854 ( .A(n35749), .B(n35753), .Z(n35850) );
  AND U44855 ( .A(n35851), .B(n35852), .Z(n35753) );
  NAND U44856 ( .A(n35853), .B(n35854), .Z(n35852) );
  NAND U44857 ( .A(n35855), .B(n35856), .Z(n35851) );
  AND U44858 ( .A(n35857), .B(n35858), .Z(n35749) );
  NAND U44859 ( .A(n35859), .B(n35860), .Z(n35858) );
  NAND U44860 ( .A(n35861), .B(n35862), .Z(n35857) );
  AND U44861 ( .A(n35863), .B(n35864), .Z(n35751) );
  XOR U44862 ( .A(n35831), .B(n35830), .Z(N62204) );
  XNOR U44863 ( .A(n35848), .B(n35849), .Z(n35830) );
  XNOR U44864 ( .A(n35863), .B(n35864), .Z(n35849) );
  XOR U44865 ( .A(n35860), .B(n35859), .Z(n35864) );
  XOR U44866 ( .A(y[2988]), .B(x[2988]), .Z(n35859) );
  XOR U44867 ( .A(n35862), .B(n35861), .Z(n35860) );
  XOR U44868 ( .A(y[2990]), .B(x[2990]), .Z(n35861) );
  XOR U44869 ( .A(y[2989]), .B(x[2989]), .Z(n35862) );
  XOR U44870 ( .A(n35854), .B(n35853), .Z(n35863) );
  XOR U44871 ( .A(n35856), .B(n35855), .Z(n35853) );
  XOR U44872 ( .A(y[2987]), .B(x[2987]), .Z(n35855) );
  XOR U44873 ( .A(y[2986]), .B(x[2986]), .Z(n35856) );
  XOR U44874 ( .A(y[2985]), .B(x[2985]), .Z(n35854) );
  XNOR U44875 ( .A(n35847), .B(n35846), .Z(n35848) );
  XNOR U44876 ( .A(n35843), .B(n35842), .Z(n35846) );
  XOR U44877 ( .A(n35845), .B(n35844), .Z(n35842) );
  XOR U44878 ( .A(y[2984]), .B(x[2984]), .Z(n35844) );
  XOR U44879 ( .A(y[2983]), .B(x[2983]), .Z(n35845) );
  XOR U44880 ( .A(y[2982]), .B(x[2982]), .Z(n35843) );
  XOR U44881 ( .A(n35837), .B(n35836), .Z(n35847) );
  XOR U44882 ( .A(n35839), .B(n35838), .Z(n35836) );
  XOR U44883 ( .A(y[2981]), .B(x[2981]), .Z(n35838) );
  XOR U44884 ( .A(y[2980]), .B(x[2980]), .Z(n35839) );
  XOR U44885 ( .A(y[2979]), .B(x[2979]), .Z(n35837) );
  XNOR U44886 ( .A(n35813), .B(n35814), .Z(n35831) );
  XNOR U44887 ( .A(n35828), .B(n35829), .Z(n35814) );
  XOR U44888 ( .A(n35825), .B(n35824), .Z(n35829) );
  XOR U44889 ( .A(y[2976]), .B(x[2976]), .Z(n35824) );
  XOR U44890 ( .A(n35827), .B(n35826), .Z(n35825) );
  XOR U44891 ( .A(y[2978]), .B(x[2978]), .Z(n35826) );
  XOR U44892 ( .A(y[2977]), .B(x[2977]), .Z(n35827) );
  XOR U44893 ( .A(n35819), .B(n35818), .Z(n35828) );
  XOR U44894 ( .A(n35821), .B(n35820), .Z(n35818) );
  XOR U44895 ( .A(y[2975]), .B(x[2975]), .Z(n35820) );
  XOR U44896 ( .A(y[2974]), .B(x[2974]), .Z(n35821) );
  XOR U44897 ( .A(y[2973]), .B(x[2973]), .Z(n35819) );
  XNOR U44898 ( .A(n35812), .B(n35811), .Z(n35813) );
  XNOR U44899 ( .A(n35808), .B(n35807), .Z(n35811) );
  XOR U44900 ( .A(n35810), .B(n35809), .Z(n35807) );
  XOR U44901 ( .A(y[2972]), .B(x[2972]), .Z(n35809) );
  XOR U44902 ( .A(y[2971]), .B(x[2971]), .Z(n35810) );
  XOR U44903 ( .A(y[2970]), .B(x[2970]), .Z(n35808) );
  XOR U44904 ( .A(n35802), .B(n35801), .Z(n35812) );
  XOR U44905 ( .A(n35804), .B(n35803), .Z(n35801) );
  XOR U44906 ( .A(y[2969]), .B(x[2969]), .Z(n35803) );
  XOR U44907 ( .A(y[2968]), .B(x[2968]), .Z(n35804) );
  XOR U44908 ( .A(y[2967]), .B(x[2967]), .Z(n35802) );
  NAND U44909 ( .A(n35865), .B(n35866), .Z(N62195) );
  NAND U44910 ( .A(n35867), .B(n35868), .Z(n35866) );
  NANDN U44911 ( .A(n35869), .B(n35870), .Z(n35868) );
  NANDN U44912 ( .A(n35870), .B(n35869), .Z(n35865) );
  XOR U44913 ( .A(n35869), .B(n35871), .Z(N62194) );
  XNOR U44914 ( .A(n35867), .B(n35870), .Z(n35871) );
  NAND U44915 ( .A(n35872), .B(n35873), .Z(n35870) );
  NAND U44916 ( .A(n35874), .B(n35875), .Z(n35873) );
  NANDN U44917 ( .A(n35876), .B(n35877), .Z(n35875) );
  NANDN U44918 ( .A(n35877), .B(n35876), .Z(n35872) );
  AND U44919 ( .A(n35878), .B(n35879), .Z(n35867) );
  NAND U44920 ( .A(n35880), .B(n35881), .Z(n35879) );
  NANDN U44921 ( .A(n35882), .B(n35883), .Z(n35881) );
  NANDN U44922 ( .A(n35883), .B(n35882), .Z(n35878) );
  IV U44923 ( .A(n35884), .Z(n35883) );
  AND U44924 ( .A(n35885), .B(n35886), .Z(n35869) );
  NAND U44925 ( .A(n35887), .B(n35888), .Z(n35886) );
  NANDN U44926 ( .A(n35889), .B(n35890), .Z(n35888) );
  NANDN U44927 ( .A(n35890), .B(n35889), .Z(n35885) );
  XOR U44928 ( .A(n35882), .B(n35891), .Z(N62193) );
  XNOR U44929 ( .A(n35880), .B(n35884), .Z(n35891) );
  XOR U44930 ( .A(n35877), .B(n35892), .Z(n35884) );
  XNOR U44931 ( .A(n35874), .B(n35876), .Z(n35892) );
  AND U44932 ( .A(n35893), .B(n35894), .Z(n35876) );
  NANDN U44933 ( .A(n35895), .B(n35896), .Z(n35894) );
  OR U44934 ( .A(n35897), .B(n35898), .Z(n35896) );
  IV U44935 ( .A(n35899), .Z(n35898) );
  NANDN U44936 ( .A(n35899), .B(n35897), .Z(n35893) );
  AND U44937 ( .A(n35900), .B(n35901), .Z(n35874) );
  NAND U44938 ( .A(n35902), .B(n35903), .Z(n35901) );
  NANDN U44939 ( .A(n35904), .B(n35905), .Z(n35903) );
  NANDN U44940 ( .A(n35905), .B(n35904), .Z(n35900) );
  IV U44941 ( .A(n35906), .Z(n35905) );
  NAND U44942 ( .A(n35907), .B(n35908), .Z(n35877) );
  NANDN U44943 ( .A(n35909), .B(n35910), .Z(n35908) );
  NANDN U44944 ( .A(n35911), .B(n35912), .Z(n35910) );
  NANDN U44945 ( .A(n35912), .B(n35911), .Z(n35907) );
  IV U44946 ( .A(n35913), .Z(n35911) );
  AND U44947 ( .A(n35914), .B(n35915), .Z(n35880) );
  NAND U44948 ( .A(n35916), .B(n35917), .Z(n35915) );
  NANDN U44949 ( .A(n35918), .B(n35919), .Z(n35917) );
  NANDN U44950 ( .A(n35919), .B(n35918), .Z(n35914) );
  XOR U44951 ( .A(n35890), .B(n35920), .Z(n35882) );
  XNOR U44952 ( .A(n35887), .B(n35889), .Z(n35920) );
  AND U44953 ( .A(n35921), .B(n35922), .Z(n35889) );
  NANDN U44954 ( .A(n35923), .B(n35924), .Z(n35922) );
  OR U44955 ( .A(n35925), .B(n35926), .Z(n35924) );
  IV U44956 ( .A(n35927), .Z(n35926) );
  NANDN U44957 ( .A(n35927), .B(n35925), .Z(n35921) );
  AND U44958 ( .A(n35928), .B(n35929), .Z(n35887) );
  NAND U44959 ( .A(n35930), .B(n35931), .Z(n35929) );
  NANDN U44960 ( .A(n35932), .B(n35933), .Z(n35931) );
  NANDN U44961 ( .A(n35933), .B(n35932), .Z(n35928) );
  IV U44962 ( .A(n35934), .Z(n35933) );
  NAND U44963 ( .A(n35935), .B(n35936), .Z(n35890) );
  NANDN U44964 ( .A(n35937), .B(n35938), .Z(n35936) );
  NANDN U44965 ( .A(n35939), .B(n35940), .Z(n35938) );
  NANDN U44966 ( .A(n35940), .B(n35939), .Z(n35935) );
  IV U44967 ( .A(n35941), .Z(n35939) );
  XOR U44968 ( .A(n35916), .B(n35942), .Z(N62192) );
  XNOR U44969 ( .A(n35919), .B(n35918), .Z(n35942) );
  XNOR U44970 ( .A(n35930), .B(n35943), .Z(n35918) );
  XNOR U44971 ( .A(n35934), .B(n35932), .Z(n35943) );
  XOR U44972 ( .A(n35940), .B(n35944), .Z(n35932) );
  XNOR U44973 ( .A(n35937), .B(n35941), .Z(n35944) );
  AND U44974 ( .A(n35945), .B(n35946), .Z(n35941) );
  NAND U44975 ( .A(n35947), .B(n35948), .Z(n35946) );
  NAND U44976 ( .A(n35949), .B(n35950), .Z(n35945) );
  AND U44977 ( .A(n35951), .B(n35952), .Z(n35937) );
  NAND U44978 ( .A(n35953), .B(n35954), .Z(n35952) );
  NAND U44979 ( .A(n35955), .B(n35956), .Z(n35951) );
  NANDN U44980 ( .A(n35957), .B(n35958), .Z(n35940) );
  ANDN U44981 ( .B(n35959), .A(n35960), .Z(n35934) );
  XNOR U44982 ( .A(n35925), .B(n35961), .Z(n35930) );
  XNOR U44983 ( .A(n35923), .B(n35927), .Z(n35961) );
  AND U44984 ( .A(n35962), .B(n35963), .Z(n35927) );
  NAND U44985 ( .A(n35964), .B(n35965), .Z(n35963) );
  NAND U44986 ( .A(n35966), .B(n35967), .Z(n35962) );
  AND U44987 ( .A(n35968), .B(n35969), .Z(n35923) );
  NAND U44988 ( .A(n35970), .B(n35971), .Z(n35969) );
  NAND U44989 ( .A(n35972), .B(n35973), .Z(n35968) );
  AND U44990 ( .A(n35974), .B(n35975), .Z(n35925) );
  NAND U44991 ( .A(n35976), .B(n35977), .Z(n35919) );
  XNOR U44992 ( .A(n35902), .B(n35978), .Z(n35916) );
  XNOR U44993 ( .A(n35906), .B(n35904), .Z(n35978) );
  XOR U44994 ( .A(n35912), .B(n35979), .Z(n35904) );
  XNOR U44995 ( .A(n35909), .B(n35913), .Z(n35979) );
  AND U44996 ( .A(n35980), .B(n35981), .Z(n35913) );
  NAND U44997 ( .A(n35982), .B(n35983), .Z(n35981) );
  NAND U44998 ( .A(n35984), .B(n35985), .Z(n35980) );
  AND U44999 ( .A(n35986), .B(n35987), .Z(n35909) );
  NAND U45000 ( .A(n35988), .B(n35989), .Z(n35987) );
  NAND U45001 ( .A(n35990), .B(n35991), .Z(n35986) );
  NANDN U45002 ( .A(n35992), .B(n35993), .Z(n35912) );
  ANDN U45003 ( .B(n35994), .A(n35995), .Z(n35906) );
  XNOR U45004 ( .A(n35897), .B(n35996), .Z(n35902) );
  XNOR U45005 ( .A(n35895), .B(n35899), .Z(n35996) );
  AND U45006 ( .A(n35997), .B(n35998), .Z(n35899) );
  NAND U45007 ( .A(n35999), .B(n36000), .Z(n35998) );
  NAND U45008 ( .A(n36001), .B(n36002), .Z(n35997) );
  AND U45009 ( .A(n36003), .B(n36004), .Z(n35895) );
  NAND U45010 ( .A(n36005), .B(n36006), .Z(n36004) );
  NAND U45011 ( .A(n36007), .B(n36008), .Z(n36003) );
  AND U45012 ( .A(n36009), .B(n36010), .Z(n35897) );
  XOR U45013 ( .A(n35977), .B(n35976), .Z(N62191) );
  XNOR U45014 ( .A(n35994), .B(n35995), .Z(n35976) );
  XNOR U45015 ( .A(n36009), .B(n36010), .Z(n35995) );
  XOR U45016 ( .A(n36006), .B(n36005), .Z(n36010) );
  XOR U45017 ( .A(y[2964]), .B(x[2964]), .Z(n36005) );
  XOR U45018 ( .A(n36008), .B(n36007), .Z(n36006) );
  XOR U45019 ( .A(y[2966]), .B(x[2966]), .Z(n36007) );
  XOR U45020 ( .A(y[2965]), .B(x[2965]), .Z(n36008) );
  XOR U45021 ( .A(n36000), .B(n35999), .Z(n36009) );
  XOR U45022 ( .A(n36002), .B(n36001), .Z(n35999) );
  XOR U45023 ( .A(y[2963]), .B(x[2963]), .Z(n36001) );
  XOR U45024 ( .A(y[2962]), .B(x[2962]), .Z(n36002) );
  XOR U45025 ( .A(y[2961]), .B(x[2961]), .Z(n36000) );
  XNOR U45026 ( .A(n35993), .B(n35992), .Z(n35994) );
  XNOR U45027 ( .A(n35989), .B(n35988), .Z(n35992) );
  XOR U45028 ( .A(n35991), .B(n35990), .Z(n35988) );
  XOR U45029 ( .A(y[2960]), .B(x[2960]), .Z(n35990) );
  XOR U45030 ( .A(y[2959]), .B(x[2959]), .Z(n35991) );
  XOR U45031 ( .A(y[2958]), .B(x[2958]), .Z(n35989) );
  XOR U45032 ( .A(n35983), .B(n35982), .Z(n35993) );
  XOR U45033 ( .A(n35985), .B(n35984), .Z(n35982) );
  XOR U45034 ( .A(y[2957]), .B(x[2957]), .Z(n35984) );
  XOR U45035 ( .A(y[2956]), .B(x[2956]), .Z(n35985) );
  XOR U45036 ( .A(y[2955]), .B(x[2955]), .Z(n35983) );
  XNOR U45037 ( .A(n35959), .B(n35960), .Z(n35977) );
  XNOR U45038 ( .A(n35974), .B(n35975), .Z(n35960) );
  XOR U45039 ( .A(n35971), .B(n35970), .Z(n35975) );
  XOR U45040 ( .A(y[2952]), .B(x[2952]), .Z(n35970) );
  XOR U45041 ( .A(n35973), .B(n35972), .Z(n35971) );
  XOR U45042 ( .A(y[2954]), .B(x[2954]), .Z(n35972) );
  XOR U45043 ( .A(y[2953]), .B(x[2953]), .Z(n35973) );
  XOR U45044 ( .A(n35965), .B(n35964), .Z(n35974) );
  XOR U45045 ( .A(n35967), .B(n35966), .Z(n35964) );
  XOR U45046 ( .A(y[2951]), .B(x[2951]), .Z(n35966) );
  XOR U45047 ( .A(y[2950]), .B(x[2950]), .Z(n35967) );
  XOR U45048 ( .A(y[2949]), .B(x[2949]), .Z(n35965) );
  XNOR U45049 ( .A(n35958), .B(n35957), .Z(n35959) );
  XNOR U45050 ( .A(n35954), .B(n35953), .Z(n35957) );
  XOR U45051 ( .A(n35956), .B(n35955), .Z(n35953) );
  XOR U45052 ( .A(y[2948]), .B(x[2948]), .Z(n35955) );
  XOR U45053 ( .A(y[2947]), .B(x[2947]), .Z(n35956) );
  XOR U45054 ( .A(y[2946]), .B(x[2946]), .Z(n35954) );
  XOR U45055 ( .A(n35948), .B(n35947), .Z(n35958) );
  XOR U45056 ( .A(n35950), .B(n35949), .Z(n35947) );
  XOR U45057 ( .A(y[2945]), .B(x[2945]), .Z(n35949) );
  XOR U45058 ( .A(y[2944]), .B(x[2944]), .Z(n35950) );
  XOR U45059 ( .A(y[2943]), .B(x[2943]), .Z(n35948) );
  NAND U45060 ( .A(n36011), .B(n36012), .Z(N62182) );
  NAND U45061 ( .A(n36013), .B(n36014), .Z(n36012) );
  NANDN U45062 ( .A(n36015), .B(n36016), .Z(n36014) );
  NANDN U45063 ( .A(n36016), .B(n36015), .Z(n36011) );
  XOR U45064 ( .A(n36015), .B(n36017), .Z(N62181) );
  XNOR U45065 ( .A(n36013), .B(n36016), .Z(n36017) );
  NAND U45066 ( .A(n36018), .B(n36019), .Z(n36016) );
  NAND U45067 ( .A(n36020), .B(n36021), .Z(n36019) );
  NANDN U45068 ( .A(n36022), .B(n36023), .Z(n36021) );
  NANDN U45069 ( .A(n36023), .B(n36022), .Z(n36018) );
  AND U45070 ( .A(n36024), .B(n36025), .Z(n36013) );
  NAND U45071 ( .A(n36026), .B(n36027), .Z(n36025) );
  NANDN U45072 ( .A(n36028), .B(n36029), .Z(n36027) );
  NANDN U45073 ( .A(n36029), .B(n36028), .Z(n36024) );
  IV U45074 ( .A(n36030), .Z(n36029) );
  AND U45075 ( .A(n36031), .B(n36032), .Z(n36015) );
  NAND U45076 ( .A(n36033), .B(n36034), .Z(n36032) );
  NANDN U45077 ( .A(n36035), .B(n36036), .Z(n36034) );
  NANDN U45078 ( .A(n36036), .B(n36035), .Z(n36031) );
  XOR U45079 ( .A(n36028), .B(n36037), .Z(N62180) );
  XNOR U45080 ( .A(n36026), .B(n36030), .Z(n36037) );
  XOR U45081 ( .A(n36023), .B(n36038), .Z(n36030) );
  XNOR U45082 ( .A(n36020), .B(n36022), .Z(n36038) );
  AND U45083 ( .A(n36039), .B(n36040), .Z(n36022) );
  NANDN U45084 ( .A(n36041), .B(n36042), .Z(n36040) );
  OR U45085 ( .A(n36043), .B(n36044), .Z(n36042) );
  IV U45086 ( .A(n36045), .Z(n36044) );
  NANDN U45087 ( .A(n36045), .B(n36043), .Z(n36039) );
  AND U45088 ( .A(n36046), .B(n36047), .Z(n36020) );
  NAND U45089 ( .A(n36048), .B(n36049), .Z(n36047) );
  NANDN U45090 ( .A(n36050), .B(n36051), .Z(n36049) );
  NANDN U45091 ( .A(n36051), .B(n36050), .Z(n36046) );
  IV U45092 ( .A(n36052), .Z(n36051) );
  NAND U45093 ( .A(n36053), .B(n36054), .Z(n36023) );
  NANDN U45094 ( .A(n36055), .B(n36056), .Z(n36054) );
  NANDN U45095 ( .A(n36057), .B(n36058), .Z(n36056) );
  NANDN U45096 ( .A(n36058), .B(n36057), .Z(n36053) );
  IV U45097 ( .A(n36059), .Z(n36057) );
  AND U45098 ( .A(n36060), .B(n36061), .Z(n36026) );
  NAND U45099 ( .A(n36062), .B(n36063), .Z(n36061) );
  NANDN U45100 ( .A(n36064), .B(n36065), .Z(n36063) );
  NANDN U45101 ( .A(n36065), .B(n36064), .Z(n36060) );
  XOR U45102 ( .A(n36036), .B(n36066), .Z(n36028) );
  XNOR U45103 ( .A(n36033), .B(n36035), .Z(n36066) );
  AND U45104 ( .A(n36067), .B(n36068), .Z(n36035) );
  NANDN U45105 ( .A(n36069), .B(n36070), .Z(n36068) );
  OR U45106 ( .A(n36071), .B(n36072), .Z(n36070) );
  IV U45107 ( .A(n36073), .Z(n36072) );
  NANDN U45108 ( .A(n36073), .B(n36071), .Z(n36067) );
  AND U45109 ( .A(n36074), .B(n36075), .Z(n36033) );
  NAND U45110 ( .A(n36076), .B(n36077), .Z(n36075) );
  NANDN U45111 ( .A(n36078), .B(n36079), .Z(n36077) );
  NANDN U45112 ( .A(n36079), .B(n36078), .Z(n36074) );
  IV U45113 ( .A(n36080), .Z(n36079) );
  NAND U45114 ( .A(n36081), .B(n36082), .Z(n36036) );
  NANDN U45115 ( .A(n36083), .B(n36084), .Z(n36082) );
  NANDN U45116 ( .A(n36085), .B(n36086), .Z(n36084) );
  NANDN U45117 ( .A(n36086), .B(n36085), .Z(n36081) );
  IV U45118 ( .A(n36087), .Z(n36085) );
  XOR U45119 ( .A(n36062), .B(n36088), .Z(N62179) );
  XNOR U45120 ( .A(n36065), .B(n36064), .Z(n36088) );
  XNOR U45121 ( .A(n36076), .B(n36089), .Z(n36064) );
  XNOR U45122 ( .A(n36080), .B(n36078), .Z(n36089) );
  XOR U45123 ( .A(n36086), .B(n36090), .Z(n36078) );
  XNOR U45124 ( .A(n36083), .B(n36087), .Z(n36090) );
  AND U45125 ( .A(n36091), .B(n36092), .Z(n36087) );
  NAND U45126 ( .A(n36093), .B(n36094), .Z(n36092) );
  NAND U45127 ( .A(n36095), .B(n36096), .Z(n36091) );
  AND U45128 ( .A(n36097), .B(n36098), .Z(n36083) );
  NAND U45129 ( .A(n36099), .B(n36100), .Z(n36098) );
  NAND U45130 ( .A(n36101), .B(n36102), .Z(n36097) );
  NANDN U45131 ( .A(n36103), .B(n36104), .Z(n36086) );
  ANDN U45132 ( .B(n36105), .A(n36106), .Z(n36080) );
  XNOR U45133 ( .A(n36071), .B(n36107), .Z(n36076) );
  XNOR U45134 ( .A(n36069), .B(n36073), .Z(n36107) );
  AND U45135 ( .A(n36108), .B(n36109), .Z(n36073) );
  NAND U45136 ( .A(n36110), .B(n36111), .Z(n36109) );
  NAND U45137 ( .A(n36112), .B(n36113), .Z(n36108) );
  AND U45138 ( .A(n36114), .B(n36115), .Z(n36069) );
  NAND U45139 ( .A(n36116), .B(n36117), .Z(n36115) );
  NAND U45140 ( .A(n36118), .B(n36119), .Z(n36114) );
  AND U45141 ( .A(n36120), .B(n36121), .Z(n36071) );
  NAND U45142 ( .A(n36122), .B(n36123), .Z(n36065) );
  XNOR U45143 ( .A(n36048), .B(n36124), .Z(n36062) );
  XNOR U45144 ( .A(n36052), .B(n36050), .Z(n36124) );
  XOR U45145 ( .A(n36058), .B(n36125), .Z(n36050) );
  XNOR U45146 ( .A(n36055), .B(n36059), .Z(n36125) );
  AND U45147 ( .A(n36126), .B(n36127), .Z(n36059) );
  NAND U45148 ( .A(n36128), .B(n36129), .Z(n36127) );
  NAND U45149 ( .A(n36130), .B(n36131), .Z(n36126) );
  AND U45150 ( .A(n36132), .B(n36133), .Z(n36055) );
  NAND U45151 ( .A(n36134), .B(n36135), .Z(n36133) );
  NAND U45152 ( .A(n36136), .B(n36137), .Z(n36132) );
  NANDN U45153 ( .A(n36138), .B(n36139), .Z(n36058) );
  ANDN U45154 ( .B(n36140), .A(n36141), .Z(n36052) );
  XNOR U45155 ( .A(n36043), .B(n36142), .Z(n36048) );
  XNOR U45156 ( .A(n36041), .B(n36045), .Z(n36142) );
  AND U45157 ( .A(n36143), .B(n36144), .Z(n36045) );
  NAND U45158 ( .A(n36145), .B(n36146), .Z(n36144) );
  NAND U45159 ( .A(n36147), .B(n36148), .Z(n36143) );
  AND U45160 ( .A(n36149), .B(n36150), .Z(n36041) );
  NAND U45161 ( .A(n36151), .B(n36152), .Z(n36150) );
  NAND U45162 ( .A(n36153), .B(n36154), .Z(n36149) );
  AND U45163 ( .A(n36155), .B(n36156), .Z(n36043) );
  XOR U45164 ( .A(n36123), .B(n36122), .Z(N62178) );
  XNOR U45165 ( .A(n36140), .B(n36141), .Z(n36122) );
  XNOR U45166 ( .A(n36155), .B(n36156), .Z(n36141) );
  XOR U45167 ( .A(n36152), .B(n36151), .Z(n36156) );
  XOR U45168 ( .A(y[2940]), .B(x[2940]), .Z(n36151) );
  XOR U45169 ( .A(n36154), .B(n36153), .Z(n36152) );
  XOR U45170 ( .A(y[2942]), .B(x[2942]), .Z(n36153) );
  XOR U45171 ( .A(y[2941]), .B(x[2941]), .Z(n36154) );
  XOR U45172 ( .A(n36146), .B(n36145), .Z(n36155) );
  XOR U45173 ( .A(n36148), .B(n36147), .Z(n36145) );
  XOR U45174 ( .A(y[2939]), .B(x[2939]), .Z(n36147) );
  XOR U45175 ( .A(y[2938]), .B(x[2938]), .Z(n36148) );
  XOR U45176 ( .A(y[2937]), .B(x[2937]), .Z(n36146) );
  XNOR U45177 ( .A(n36139), .B(n36138), .Z(n36140) );
  XNOR U45178 ( .A(n36135), .B(n36134), .Z(n36138) );
  XOR U45179 ( .A(n36137), .B(n36136), .Z(n36134) );
  XOR U45180 ( .A(y[2936]), .B(x[2936]), .Z(n36136) );
  XOR U45181 ( .A(y[2935]), .B(x[2935]), .Z(n36137) );
  XOR U45182 ( .A(y[2934]), .B(x[2934]), .Z(n36135) );
  XOR U45183 ( .A(n36129), .B(n36128), .Z(n36139) );
  XOR U45184 ( .A(n36131), .B(n36130), .Z(n36128) );
  XOR U45185 ( .A(y[2933]), .B(x[2933]), .Z(n36130) );
  XOR U45186 ( .A(y[2932]), .B(x[2932]), .Z(n36131) );
  XOR U45187 ( .A(y[2931]), .B(x[2931]), .Z(n36129) );
  XNOR U45188 ( .A(n36105), .B(n36106), .Z(n36123) );
  XNOR U45189 ( .A(n36120), .B(n36121), .Z(n36106) );
  XOR U45190 ( .A(n36117), .B(n36116), .Z(n36121) );
  XOR U45191 ( .A(y[2928]), .B(x[2928]), .Z(n36116) );
  XOR U45192 ( .A(n36119), .B(n36118), .Z(n36117) );
  XOR U45193 ( .A(y[2930]), .B(x[2930]), .Z(n36118) );
  XOR U45194 ( .A(y[2929]), .B(x[2929]), .Z(n36119) );
  XOR U45195 ( .A(n36111), .B(n36110), .Z(n36120) );
  XOR U45196 ( .A(n36113), .B(n36112), .Z(n36110) );
  XOR U45197 ( .A(y[2927]), .B(x[2927]), .Z(n36112) );
  XOR U45198 ( .A(y[2926]), .B(x[2926]), .Z(n36113) );
  XOR U45199 ( .A(y[2925]), .B(x[2925]), .Z(n36111) );
  XNOR U45200 ( .A(n36104), .B(n36103), .Z(n36105) );
  XNOR U45201 ( .A(n36100), .B(n36099), .Z(n36103) );
  XOR U45202 ( .A(n36102), .B(n36101), .Z(n36099) );
  XOR U45203 ( .A(y[2924]), .B(x[2924]), .Z(n36101) );
  XOR U45204 ( .A(y[2923]), .B(x[2923]), .Z(n36102) );
  XOR U45205 ( .A(y[2922]), .B(x[2922]), .Z(n36100) );
  XOR U45206 ( .A(n36094), .B(n36093), .Z(n36104) );
  XOR U45207 ( .A(n36096), .B(n36095), .Z(n36093) );
  XOR U45208 ( .A(y[2921]), .B(x[2921]), .Z(n36095) );
  XOR U45209 ( .A(y[2920]), .B(x[2920]), .Z(n36096) );
  XOR U45210 ( .A(y[2919]), .B(x[2919]), .Z(n36094) );
  NAND U45211 ( .A(n36157), .B(n36158), .Z(N62169) );
  NAND U45212 ( .A(n36159), .B(n36160), .Z(n36158) );
  NANDN U45213 ( .A(n36161), .B(n36162), .Z(n36160) );
  NANDN U45214 ( .A(n36162), .B(n36161), .Z(n36157) );
  XOR U45215 ( .A(n36161), .B(n36163), .Z(N62168) );
  XNOR U45216 ( .A(n36159), .B(n36162), .Z(n36163) );
  NAND U45217 ( .A(n36164), .B(n36165), .Z(n36162) );
  NAND U45218 ( .A(n36166), .B(n36167), .Z(n36165) );
  NANDN U45219 ( .A(n36168), .B(n36169), .Z(n36167) );
  NANDN U45220 ( .A(n36169), .B(n36168), .Z(n36164) );
  AND U45221 ( .A(n36170), .B(n36171), .Z(n36159) );
  NAND U45222 ( .A(n36172), .B(n36173), .Z(n36171) );
  NANDN U45223 ( .A(n36174), .B(n36175), .Z(n36173) );
  NANDN U45224 ( .A(n36175), .B(n36174), .Z(n36170) );
  IV U45225 ( .A(n36176), .Z(n36175) );
  AND U45226 ( .A(n36177), .B(n36178), .Z(n36161) );
  NAND U45227 ( .A(n36179), .B(n36180), .Z(n36178) );
  NANDN U45228 ( .A(n36181), .B(n36182), .Z(n36180) );
  NANDN U45229 ( .A(n36182), .B(n36181), .Z(n36177) );
  XOR U45230 ( .A(n36174), .B(n36183), .Z(N62167) );
  XNOR U45231 ( .A(n36172), .B(n36176), .Z(n36183) );
  XOR U45232 ( .A(n36169), .B(n36184), .Z(n36176) );
  XNOR U45233 ( .A(n36166), .B(n36168), .Z(n36184) );
  AND U45234 ( .A(n36185), .B(n36186), .Z(n36168) );
  NANDN U45235 ( .A(n36187), .B(n36188), .Z(n36186) );
  OR U45236 ( .A(n36189), .B(n36190), .Z(n36188) );
  IV U45237 ( .A(n36191), .Z(n36190) );
  NANDN U45238 ( .A(n36191), .B(n36189), .Z(n36185) );
  AND U45239 ( .A(n36192), .B(n36193), .Z(n36166) );
  NAND U45240 ( .A(n36194), .B(n36195), .Z(n36193) );
  NANDN U45241 ( .A(n36196), .B(n36197), .Z(n36195) );
  NANDN U45242 ( .A(n36197), .B(n36196), .Z(n36192) );
  IV U45243 ( .A(n36198), .Z(n36197) );
  NAND U45244 ( .A(n36199), .B(n36200), .Z(n36169) );
  NANDN U45245 ( .A(n36201), .B(n36202), .Z(n36200) );
  NANDN U45246 ( .A(n36203), .B(n36204), .Z(n36202) );
  NANDN U45247 ( .A(n36204), .B(n36203), .Z(n36199) );
  IV U45248 ( .A(n36205), .Z(n36203) );
  AND U45249 ( .A(n36206), .B(n36207), .Z(n36172) );
  NAND U45250 ( .A(n36208), .B(n36209), .Z(n36207) );
  NANDN U45251 ( .A(n36210), .B(n36211), .Z(n36209) );
  NANDN U45252 ( .A(n36211), .B(n36210), .Z(n36206) );
  XOR U45253 ( .A(n36182), .B(n36212), .Z(n36174) );
  XNOR U45254 ( .A(n36179), .B(n36181), .Z(n36212) );
  AND U45255 ( .A(n36213), .B(n36214), .Z(n36181) );
  NANDN U45256 ( .A(n36215), .B(n36216), .Z(n36214) );
  OR U45257 ( .A(n36217), .B(n36218), .Z(n36216) );
  IV U45258 ( .A(n36219), .Z(n36218) );
  NANDN U45259 ( .A(n36219), .B(n36217), .Z(n36213) );
  AND U45260 ( .A(n36220), .B(n36221), .Z(n36179) );
  NAND U45261 ( .A(n36222), .B(n36223), .Z(n36221) );
  NANDN U45262 ( .A(n36224), .B(n36225), .Z(n36223) );
  NANDN U45263 ( .A(n36225), .B(n36224), .Z(n36220) );
  IV U45264 ( .A(n36226), .Z(n36225) );
  NAND U45265 ( .A(n36227), .B(n36228), .Z(n36182) );
  NANDN U45266 ( .A(n36229), .B(n36230), .Z(n36228) );
  NANDN U45267 ( .A(n36231), .B(n36232), .Z(n36230) );
  NANDN U45268 ( .A(n36232), .B(n36231), .Z(n36227) );
  IV U45269 ( .A(n36233), .Z(n36231) );
  XOR U45270 ( .A(n36208), .B(n36234), .Z(N62166) );
  XNOR U45271 ( .A(n36211), .B(n36210), .Z(n36234) );
  XNOR U45272 ( .A(n36222), .B(n36235), .Z(n36210) );
  XNOR U45273 ( .A(n36226), .B(n36224), .Z(n36235) );
  XOR U45274 ( .A(n36232), .B(n36236), .Z(n36224) );
  XNOR U45275 ( .A(n36229), .B(n36233), .Z(n36236) );
  AND U45276 ( .A(n36237), .B(n36238), .Z(n36233) );
  NAND U45277 ( .A(n36239), .B(n36240), .Z(n36238) );
  NAND U45278 ( .A(n36241), .B(n36242), .Z(n36237) );
  AND U45279 ( .A(n36243), .B(n36244), .Z(n36229) );
  NAND U45280 ( .A(n36245), .B(n36246), .Z(n36244) );
  NAND U45281 ( .A(n36247), .B(n36248), .Z(n36243) );
  NANDN U45282 ( .A(n36249), .B(n36250), .Z(n36232) );
  ANDN U45283 ( .B(n36251), .A(n36252), .Z(n36226) );
  XNOR U45284 ( .A(n36217), .B(n36253), .Z(n36222) );
  XNOR U45285 ( .A(n36215), .B(n36219), .Z(n36253) );
  AND U45286 ( .A(n36254), .B(n36255), .Z(n36219) );
  NAND U45287 ( .A(n36256), .B(n36257), .Z(n36255) );
  NAND U45288 ( .A(n36258), .B(n36259), .Z(n36254) );
  AND U45289 ( .A(n36260), .B(n36261), .Z(n36215) );
  NAND U45290 ( .A(n36262), .B(n36263), .Z(n36261) );
  NAND U45291 ( .A(n36264), .B(n36265), .Z(n36260) );
  AND U45292 ( .A(n36266), .B(n36267), .Z(n36217) );
  NAND U45293 ( .A(n36268), .B(n36269), .Z(n36211) );
  XNOR U45294 ( .A(n36194), .B(n36270), .Z(n36208) );
  XNOR U45295 ( .A(n36198), .B(n36196), .Z(n36270) );
  XOR U45296 ( .A(n36204), .B(n36271), .Z(n36196) );
  XNOR U45297 ( .A(n36201), .B(n36205), .Z(n36271) );
  AND U45298 ( .A(n36272), .B(n36273), .Z(n36205) );
  NAND U45299 ( .A(n36274), .B(n36275), .Z(n36273) );
  NAND U45300 ( .A(n36276), .B(n36277), .Z(n36272) );
  AND U45301 ( .A(n36278), .B(n36279), .Z(n36201) );
  NAND U45302 ( .A(n36280), .B(n36281), .Z(n36279) );
  NAND U45303 ( .A(n36282), .B(n36283), .Z(n36278) );
  NANDN U45304 ( .A(n36284), .B(n36285), .Z(n36204) );
  ANDN U45305 ( .B(n36286), .A(n36287), .Z(n36198) );
  XNOR U45306 ( .A(n36189), .B(n36288), .Z(n36194) );
  XNOR U45307 ( .A(n36187), .B(n36191), .Z(n36288) );
  AND U45308 ( .A(n36289), .B(n36290), .Z(n36191) );
  NAND U45309 ( .A(n36291), .B(n36292), .Z(n36290) );
  NAND U45310 ( .A(n36293), .B(n36294), .Z(n36289) );
  AND U45311 ( .A(n36295), .B(n36296), .Z(n36187) );
  NAND U45312 ( .A(n36297), .B(n36298), .Z(n36296) );
  NAND U45313 ( .A(n36299), .B(n36300), .Z(n36295) );
  AND U45314 ( .A(n36301), .B(n36302), .Z(n36189) );
  XOR U45315 ( .A(n36269), .B(n36268), .Z(N62165) );
  XNOR U45316 ( .A(n36286), .B(n36287), .Z(n36268) );
  XNOR U45317 ( .A(n36301), .B(n36302), .Z(n36287) );
  XOR U45318 ( .A(n36298), .B(n36297), .Z(n36302) );
  XOR U45319 ( .A(y[2916]), .B(x[2916]), .Z(n36297) );
  XOR U45320 ( .A(n36300), .B(n36299), .Z(n36298) );
  XOR U45321 ( .A(y[2918]), .B(x[2918]), .Z(n36299) );
  XOR U45322 ( .A(y[2917]), .B(x[2917]), .Z(n36300) );
  XOR U45323 ( .A(n36292), .B(n36291), .Z(n36301) );
  XOR U45324 ( .A(n36294), .B(n36293), .Z(n36291) );
  XOR U45325 ( .A(y[2915]), .B(x[2915]), .Z(n36293) );
  XOR U45326 ( .A(y[2914]), .B(x[2914]), .Z(n36294) );
  XOR U45327 ( .A(y[2913]), .B(x[2913]), .Z(n36292) );
  XNOR U45328 ( .A(n36285), .B(n36284), .Z(n36286) );
  XNOR U45329 ( .A(n36281), .B(n36280), .Z(n36284) );
  XOR U45330 ( .A(n36283), .B(n36282), .Z(n36280) );
  XOR U45331 ( .A(y[2912]), .B(x[2912]), .Z(n36282) );
  XOR U45332 ( .A(y[2911]), .B(x[2911]), .Z(n36283) );
  XOR U45333 ( .A(y[2910]), .B(x[2910]), .Z(n36281) );
  XOR U45334 ( .A(n36275), .B(n36274), .Z(n36285) );
  XOR U45335 ( .A(n36277), .B(n36276), .Z(n36274) );
  XOR U45336 ( .A(y[2909]), .B(x[2909]), .Z(n36276) );
  XOR U45337 ( .A(y[2908]), .B(x[2908]), .Z(n36277) );
  XOR U45338 ( .A(y[2907]), .B(x[2907]), .Z(n36275) );
  XNOR U45339 ( .A(n36251), .B(n36252), .Z(n36269) );
  XNOR U45340 ( .A(n36266), .B(n36267), .Z(n36252) );
  XOR U45341 ( .A(n36263), .B(n36262), .Z(n36267) );
  XOR U45342 ( .A(y[2904]), .B(x[2904]), .Z(n36262) );
  XOR U45343 ( .A(n36265), .B(n36264), .Z(n36263) );
  XOR U45344 ( .A(y[2906]), .B(x[2906]), .Z(n36264) );
  XOR U45345 ( .A(y[2905]), .B(x[2905]), .Z(n36265) );
  XOR U45346 ( .A(n36257), .B(n36256), .Z(n36266) );
  XOR U45347 ( .A(n36259), .B(n36258), .Z(n36256) );
  XOR U45348 ( .A(y[2903]), .B(x[2903]), .Z(n36258) );
  XOR U45349 ( .A(y[2902]), .B(x[2902]), .Z(n36259) );
  XOR U45350 ( .A(y[2901]), .B(x[2901]), .Z(n36257) );
  XNOR U45351 ( .A(n36250), .B(n36249), .Z(n36251) );
  XNOR U45352 ( .A(n36246), .B(n36245), .Z(n36249) );
  XOR U45353 ( .A(n36248), .B(n36247), .Z(n36245) );
  XOR U45354 ( .A(y[2900]), .B(x[2900]), .Z(n36247) );
  XOR U45355 ( .A(y[2899]), .B(x[2899]), .Z(n36248) );
  XOR U45356 ( .A(y[2898]), .B(x[2898]), .Z(n36246) );
  XOR U45357 ( .A(n36240), .B(n36239), .Z(n36250) );
  XOR U45358 ( .A(n36242), .B(n36241), .Z(n36239) );
  XOR U45359 ( .A(y[2897]), .B(x[2897]), .Z(n36241) );
  XOR U45360 ( .A(y[2896]), .B(x[2896]), .Z(n36242) );
  XOR U45361 ( .A(y[2895]), .B(x[2895]), .Z(n36240) );
  NAND U45362 ( .A(n36303), .B(n36304), .Z(N62156) );
  NAND U45363 ( .A(n36305), .B(n36306), .Z(n36304) );
  NANDN U45364 ( .A(n36307), .B(n36308), .Z(n36306) );
  NANDN U45365 ( .A(n36308), .B(n36307), .Z(n36303) );
  XOR U45366 ( .A(n36307), .B(n36309), .Z(N62155) );
  XNOR U45367 ( .A(n36305), .B(n36308), .Z(n36309) );
  NAND U45368 ( .A(n36310), .B(n36311), .Z(n36308) );
  NAND U45369 ( .A(n36312), .B(n36313), .Z(n36311) );
  NANDN U45370 ( .A(n36314), .B(n36315), .Z(n36313) );
  NANDN U45371 ( .A(n36315), .B(n36314), .Z(n36310) );
  AND U45372 ( .A(n36316), .B(n36317), .Z(n36305) );
  NAND U45373 ( .A(n36318), .B(n36319), .Z(n36317) );
  NANDN U45374 ( .A(n36320), .B(n36321), .Z(n36319) );
  NANDN U45375 ( .A(n36321), .B(n36320), .Z(n36316) );
  IV U45376 ( .A(n36322), .Z(n36321) );
  AND U45377 ( .A(n36323), .B(n36324), .Z(n36307) );
  NAND U45378 ( .A(n36325), .B(n36326), .Z(n36324) );
  NANDN U45379 ( .A(n36327), .B(n36328), .Z(n36326) );
  NANDN U45380 ( .A(n36328), .B(n36327), .Z(n36323) );
  XOR U45381 ( .A(n36320), .B(n36329), .Z(N62154) );
  XNOR U45382 ( .A(n36318), .B(n36322), .Z(n36329) );
  XOR U45383 ( .A(n36315), .B(n36330), .Z(n36322) );
  XNOR U45384 ( .A(n36312), .B(n36314), .Z(n36330) );
  AND U45385 ( .A(n36331), .B(n36332), .Z(n36314) );
  NANDN U45386 ( .A(n36333), .B(n36334), .Z(n36332) );
  OR U45387 ( .A(n36335), .B(n36336), .Z(n36334) );
  IV U45388 ( .A(n36337), .Z(n36336) );
  NANDN U45389 ( .A(n36337), .B(n36335), .Z(n36331) );
  AND U45390 ( .A(n36338), .B(n36339), .Z(n36312) );
  NAND U45391 ( .A(n36340), .B(n36341), .Z(n36339) );
  NANDN U45392 ( .A(n36342), .B(n36343), .Z(n36341) );
  NANDN U45393 ( .A(n36343), .B(n36342), .Z(n36338) );
  IV U45394 ( .A(n36344), .Z(n36343) );
  NAND U45395 ( .A(n36345), .B(n36346), .Z(n36315) );
  NANDN U45396 ( .A(n36347), .B(n36348), .Z(n36346) );
  NANDN U45397 ( .A(n36349), .B(n36350), .Z(n36348) );
  NANDN U45398 ( .A(n36350), .B(n36349), .Z(n36345) );
  IV U45399 ( .A(n36351), .Z(n36349) );
  AND U45400 ( .A(n36352), .B(n36353), .Z(n36318) );
  NAND U45401 ( .A(n36354), .B(n36355), .Z(n36353) );
  NANDN U45402 ( .A(n36356), .B(n36357), .Z(n36355) );
  NANDN U45403 ( .A(n36357), .B(n36356), .Z(n36352) );
  XOR U45404 ( .A(n36328), .B(n36358), .Z(n36320) );
  XNOR U45405 ( .A(n36325), .B(n36327), .Z(n36358) );
  AND U45406 ( .A(n36359), .B(n36360), .Z(n36327) );
  NANDN U45407 ( .A(n36361), .B(n36362), .Z(n36360) );
  OR U45408 ( .A(n36363), .B(n36364), .Z(n36362) );
  IV U45409 ( .A(n36365), .Z(n36364) );
  NANDN U45410 ( .A(n36365), .B(n36363), .Z(n36359) );
  AND U45411 ( .A(n36366), .B(n36367), .Z(n36325) );
  NAND U45412 ( .A(n36368), .B(n36369), .Z(n36367) );
  NANDN U45413 ( .A(n36370), .B(n36371), .Z(n36369) );
  NANDN U45414 ( .A(n36371), .B(n36370), .Z(n36366) );
  IV U45415 ( .A(n36372), .Z(n36371) );
  NAND U45416 ( .A(n36373), .B(n36374), .Z(n36328) );
  NANDN U45417 ( .A(n36375), .B(n36376), .Z(n36374) );
  NANDN U45418 ( .A(n36377), .B(n36378), .Z(n36376) );
  NANDN U45419 ( .A(n36378), .B(n36377), .Z(n36373) );
  IV U45420 ( .A(n36379), .Z(n36377) );
  XOR U45421 ( .A(n36354), .B(n36380), .Z(N62153) );
  XNOR U45422 ( .A(n36357), .B(n36356), .Z(n36380) );
  XNOR U45423 ( .A(n36368), .B(n36381), .Z(n36356) );
  XNOR U45424 ( .A(n36372), .B(n36370), .Z(n36381) );
  XOR U45425 ( .A(n36378), .B(n36382), .Z(n36370) );
  XNOR U45426 ( .A(n36375), .B(n36379), .Z(n36382) );
  AND U45427 ( .A(n36383), .B(n36384), .Z(n36379) );
  NAND U45428 ( .A(n36385), .B(n36386), .Z(n36384) );
  NAND U45429 ( .A(n36387), .B(n36388), .Z(n36383) );
  AND U45430 ( .A(n36389), .B(n36390), .Z(n36375) );
  NAND U45431 ( .A(n36391), .B(n36392), .Z(n36390) );
  NAND U45432 ( .A(n36393), .B(n36394), .Z(n36389) );
  NANDN U45433 ( .A(n36395), .B(n36396), .Z(n36378) );
  ANDN U45434 ( .B(n36397), .A(n36398), .Z(n36372) );
  XNOR U45435 ( .A(n36363), .B(n36399), .Z(n36368) );
  XNOR U45436 ( .A(n36361), .B(n36365), .Z(n36399) );
  AND U45437 ( .A(n36400), .B(n36401), .Z(n36365) );
  NAND U45438 ( .A(n36402), .B(n36403), .Z(n36401) );
  NAND U45439 ( .A(n36404), .B(n36405), .Z(n36400) );
  AND U45440 ( .A(n36406), .B(n36407), .Z(n36361) );
  NAND U45441 ( .A(n36408), .B(n36409), .Z(n36407) );
  NAND U45442 ( .A(n36410), .B(n36411), .Z(n36406) );
  AND U45443 ( .A(n36412), .B(n36413), .Z(n36363) );
  NAND U45444 ( .A(n36414), .B(n36415), .Z(n36357) );
  XNOR U45445 ( .A(n36340), .B(n36416), .Z(n36354) );
  XNOR U45446 ( .A(n36344), .B(n36342), .Z(n36416) );
  XOR U45447 ( .A(n36350), .B(n36417), .Z(n36342) );
  XNOR U45448 ( .A(n36347), .B(n36351), .Z(n36417) );
  AND U45449 ( .A(n36418), .B(n36419), .Z(n36351) );
  NAND U45450 ( .A(n36420), .B(n36421), .Z(n36419) );
  NAND U45451 ( .A(n36422), .B(n36423), .Z(n36418) );
  AND U45452 ( .A(n36424), .B(n36425), .Z(n36347) );
  NAND U45453 ( .A(n36426), .B(n36427), .Z(n36425) );
  NAND U45454 ( .A(n36428), .B(n36429), .Z(n36424) );
  NANDN U45455 ( .A(n36430), .B(n36431), .Z(n36350) );
  ANDN U45456 ( .B(n36432), .A(n36433), .Z(n36344) );
  XNOR U45457 ( .A(n36335), .B(n36434), .Z(n36340) );
  XNOR U45458 ( .A(n36333), .B(n36337), .Z(n36434) );
  AND U45459 ( .A(n36435), .B(n36436), .Z(n36337) );
  NAND U45460 ( .A(n36437), .B(n36438), .Z(n36436) );
  NAND U45461 ( .A(n36439), .B(n36440), .Z(n36435) );
  AND U45462 ( .A(n36441), .B(n36442), .Z(n36333) );
  NAND U45463 ( .A(n36443), .B(n36444), .Z(n36442) );
  NAND U45464 ( .A(n36445), .B(n36446), .Z(n36441) );
  AND U45465 ( .A(n36447), .B(n36448), .Z(n36335) );
  XOR U45466 ( .A(n36415), .B(n36414), .Z(N62152) );
  XNOR U45467 ( .A(n36432), .B(n36433), .Z(n36414) );
  XNOR U45468 ( .A(n36447), .B(n36448), .Z(n36433) );
  XOR U45469 ( .A(n36444), .B(n36443), .Z(n36448) );
  XOR U45470 ( .A(y[2892]), .B(x[2892]), .Z(n36443) );
  XOR U45471 ( .A(n36446), .B(n36445), .Z(n36444) );
  XOR U45472 ( .A(y[2894]), .B(x[2894]), .Z(n36445) );
  XOR U45473 ( .A(y[2893]), .B(x[2893]), .Z(n36446) );
  XOR U45474 ( .A(n36438), .B(n36437), .Z(n36447) );
  XOR U45475 ( .A(n36440), .B(n36439), .Z(n36437) );
  XOR U45476 ( .A(y[2891]), .B(x[2891]), .Z(n36439) );
  XOR U45477 ( .A(y[2890]), .B(x[2890]), .Z(n36440) );
  XOR U45478 ( .A(y[2889]), .B(x[2889]), .Z(n36438) );
  XNOR U45479 ( .A(n36431), .B(n36430), .Z(n36432) );
  XNOR U45480 ( .A(n36427), .B(n36426), .Z(n36430) );
  XOR U45481 ( .A(n36429), .B(n36428), .Z(n36426) );
  XOR U45482 ( .A(y[2888]), .B(x[2888]), .Z(n36428) );
  XOR U45483 ( .A(y[2887]), .B(x[2887]), .Z(n36429) );
  XOR U45484 ( .A(y[2886]), .B(x[2886]), .Z(n36427) );
  XOR U45485 ( .A(n36421), .B(n36420), .Z(n36431) );
  XOR U45486 ( .A(n36423), .B(n36422), .Z(n36420) );
  XOR U45487 ( .A(y[2885]), .B(x[2885]), .Z(n36422) );
  XOR U45488 ( .A(y[2884]), .B(x[2884]), .Z(n36423) );
  XOR U45489 ( .A(y[2883]), .B(x[2883]), .Z(n36421) );
  XNOR U45490 ( .A(n36397), .B(n36398), .Z(n36415) );
  XNOR U45491 ( .A(n36412), .B(n36413), .Z(n36398) );
  XOR U45492 ( .A(n36409), .B(n36408), .Z(n36413) );
  XOR U45493 ( .A(y[2880]), .B(x[2880]), .Z(n36408) );
  XOR U45494 ( .A(n36411), .B(n36410), .Z(n36409) );
  XOR U45495 ( .A(y[2882]), .B(x[2882]), .Z(n36410) );
  XOR U45496 ( .A(y[2881]), .B(x[2881]), .Z(n36411) );
  XOR U45497 ( .A(n36403), .B(n36402), .Z(n36412) );
  XOR U45498 ( .A(n36405), .B(n36404), .Z(n36402) );
  XOR U45499 ( .A(y[2879]), .B(x[2879]), .Z(n36404) );
  XOR U45500 ( .A(y[2878]), .B(x[2878]), .Z(n36405) );
  XOR U45501 ( .A(y[2877]), .B(x[2877]), .Z(n36403) );
  XNOR U45502 ( .A(n36396), .B(n36395), .Z(n36397) );
  XNOR U45503 ( .A(n36392), .B(n36391), .Z(n36395) );
  XOR U45504 ( .A(n36394), .B(n36393), .Z(n36391) );
  XOR U45505 ( .A(y[2876]), .B(x[2876]), .Z(n36393) );
  XOR U45506 ( .A(y[2875]), .B(x[2875]), .Z(n36394) );
  XOR U45507 ( .A(y[2874]), .B(x[2874]), .Z(n36392) );
  XOR U45508 ( .A(n36386), .B(n36385), .Z(n36396) );
  XOR U45509 ( .A(n36388), .B(n36387), .Z(n36385) );
  XOR U45510 ( .A(y[2873]), .B(x[2873]), .Z(n36387) );
  XOR U45511 ( .A(y[2872]), .B(x[2872]), .Z(n36388) );
  XOR U45512 ( .A(y[2871]), .B(x[2871]), .Z(n36386) );
  NAND U45513 ( .A(n36449), .B(n36450), .Z(N62143) );
  NAND U45514 ( .A(n36451), .B(n36452), .Z(n36450) );
  NANDN U45515 ( .A(n36453), .B(n36454), .Z(n36452) );
  NANDN U45516 ( .A(n36454), .B(n36453), .Z(n36449) );
  XOR U45517 ( .A(n36453), .B(n36455), .Z(N62142) );
  XNOR U45518 ( .A(n36451), .B(n36454), .Z(n36455) );
  NAND U45519 ( .A(n36456), .B(n36457), .Z(n36454) );
  NAND U45520 ( .A(n36458), .B(n36459), .Z(n36457) );
  NANDN U45521 ( .A(n36460), .B(n36461), .Z(n36459) );
  NANDN U45522 ( .A(n36461), .B(n36460), .Z(n36456) );
  AND U45523 ( .A(n36462), .B(n36463), .Z(n36451) );
  NAND U45524 ( .A(n36464), .B(n36465), .Z(n36463) );
  NANDN U45525 ( .A(n36466), .B(n36467), .Z(n36465) );
  NANDN U45526 ( .A(n36467), .B(n36466), .Z(n36462) );
  IV U45527 ( .A(n36468), .Z(n36467) );
  AND U45528 ( .A(n36469), .B(n36470), .Z(n36453) );
  NAND U45529 ( .A(n36471), .B(n36472), .Z(n36470) );
  NANDN U45530 ( .A(n36473), .B(n36474), .Z(n36472) );
  NANDN U45531 ( .A(n36474), .B(n36473), .Z(n36469) );
  XOR U45532 ( .A(n36466), .B(n36475), .Z(N62141) );
  XNOR U45533 ( .A(n36464), .B(n36468), .Z(n36475) );
  XOR U45534 ( .A(n36461), .B(n36476), .Z(n36468) );
  XNOR U45535 ( .A(n36458), .B(n36460), .Z(n36476) );
  AND U45536 ( .A(n36477), .B(n36478), .Z(n36460) );
  NANDN U45537 ( .A(n36479), .B(n36480), .Z(n36478) );
  OR U45538 ( .A(n36481), .B(n36482), .Z(n36480) );
  IV U45539 ( .A(n36483), .Z(n36482) );
  NANDN U45540 ( .A(n36483), .B(n36481), .Z(n36477) );
  AND U45541 ( .A(n36484), .B(n36485), .Z(n36458) );
  NAND U45542 ( .A(n36486), .B(n36487), .Z(n36485) );
  NANDN U45543 ( .A(n36488), .B(n36489), .Z(n36487) );
  NANDN U45544 ( .A(n36489), .B(n36488), .Z(n36484) );
  IV U45545 ( .A(n36490), .Z(n36489) );
  NAND U45546 ( .A(n36491), .B(n36492), .Z(n36461) );
  NANDN U45547 ( .A(n36493), .B(n36494), .Z(n36492) );
  NANDN U45548 ( .A(n36495), .B(n36496), .Z(n36494) );
  NANDN U45549 ( .A(n36496), .B(n36495), .Z(n36491) );
  IV U45550 ( .A(n36497), .Z(n36495) );
  AND U45551 ( .A(n36498), .B(n36499), .Z(n36464) );
  NAND U45552 ( .A(n36500), .B(n36501), .Z(n36499) );
  NANDN U45553 ( .A(n36502), .B(n36503), .Z(n36501) );
  NANDN U45554 ( .A(n36503), .B(n36502), .Z(n36498) );
  XOR U45555 ( .A(n36474), .B(n36504), .Z(n36466) );
  XNOR U45556 ( .A(n36471), .B(n36473), .Z(n36504) );
  AND U45557 ( .A(n36505), .B(n36506), .Z(n36473) );
  NANDN U45558 ( .A(n36507), .B(n36508), .Z(n36506) );
  OR U45559 ( .A(n36509), .B(n36510), .Z(n36508) );
  IV U45560 ( .A(n36511), .Z(n36510) );
  NANDN U45561 ( .A(n36511), .B(n36509), .Z(n36505) );
  AND U45562 ( .A(n36512), .B(n36513), .Z(n36471) );
  NAND U45563 ( .A(n36514), .B(n36515), .Z(n36513) );
  NANDN U45564 ( .A(n36516), .B(n36517), .Z(n36515) );
  NANDN U45565 ( .A(n36517), .B(n36516), .Z(n36512) );
  IV U45566 ( .A(n36518), .Z(n36517) );
  NAND U45567 ( .A(n36519), .B(n36520), .Z(n36474) );
  NANDN U45568 ( .A(n36521), .B(n36522), .Z(n36520) );
  NANDN U45569 ( .A(n36523), .B(n36524), .Z(n36522) );
  NANDN U45570 ( .A(n36524), .B(n36523), .Z(n36519) );
  IV U45571 ( .A(n36525), .Z(n36523) );
  XOR U45572 ( .A(n36500), .B(n36526), .Z(N62140) );
  XNOR U45573 ( .A(n36503), .B(n36502), .Z(n36526) );
  XNOR U45574 ( .A(n36514), .B(n36527), .Z(n36502) );
  XNOR U45575 ( .A(n36518), .B(n36516), .Z(n36527) );
  XOR U45576 ( .A(n36524), .B(n36528), .Z(n36516) );
  XNOR U45577 ( .A(n36521), .B(n36525), .Z(n36528) );
  AND U45578 ( .A(n36529), .B(n36530), .Z(n36525) );
  NAND U45579 ( .A(n36531), .B(n36532), .Z(n36530) );
  NAND U45580 ( .A(n36533), .B(n36534), .Z(n36529) );
  AND U45581 ( .A(n36535), .B(n36536), .Z(n36521) );
  NAND U45582 ( .A(n36537), .B(n36538), .Z(n36536) );
  NAND U45583 ( .A(n36539), .B(n36540), .Z(n36535) );
  NANDN U45584 ( .A(n36541), .B(n36542), .Z(n36524) );
  ANDN U45585 ( .B(n36543), .A(n36544), .Z(n36518) );
  XNOR U45586 ( .A(n36509), .B(n36545), .Z(n36514) );
  XNOR U45587 ( .A(n36507), .B(n36511), .Z(n36545) );
  AND U45588 ( .A(n36546), .B(n36547), .Z(n36511) );
  NAND U45589 ( .A(n36548), .B(n36549), .Z(n36547) );
  NAND U45590 ( .A(n36550), .B(n36551), .Z(n36546) );
  AND U45591 ( .A(n36552), .B(n36553), .Z(n36507) );
  NAND U45592 ( .A(n36554), .B(n36555), .Z(n36553) );
  NAND U45593 ( .A(n36556), .B(n36557), .Z(n36552) );
  AND U45594 ( .A(n36558), .B(n36559), .Z(n36509) );
  NAND U45595 ( .A(n36560), .B(n36561), .Z(n36503) );
  XNOR U45596 ( .A(n36486), .B(n36562), .Z(n36500) );
  XNOR U45597 ( .A(n36490), .B(n36488), .Z(n36562) );
  XOR U45598 ( .A(n36496), .B(n36563), .Z(n36488) );
  XNOR U45599 ( .A(n36493), .B(n36497), .Z(n36563) );
  AND U45600 ( .A(n36564), .B(n36565), .Z(n36497) );
  NAND U45601 ( .A(n36566), .B(n36567), .Z(n36565) );
  NAND U45602 ( .A(n36568), .B(n36569), .Z(n36564) );
  AND U45603 ( .A(n36570), .B(n36571), .Z(n36493) );
  NAND U45604 ( .A(n36572), .B(n36573), .Z(n36571) );
  NAND U45605 ( .A(n36574), .B(n36575), .Z(n36570) );
  NANDN U45606 ( .A(n36576), .B(n36577), .Z(n36496) );
  ANDN U45607 ( .B(n36578), .A(n36579), .Z(n36490) );
  XNOR U45608 ( .A(n36481), .B(n36580), .Z(n36486) );
  XNOR U45609 ( .A(n36479), .B(n36483), .Z(n36580) );
  AND U45610 ( .A(n36581), .B(n36582), .Z(n36483) );
  NAND U45611 ( .A(n36583), .B(n36584), .Z(n36582) );
  NAND U45612 ( .A(n36585), .B(n36586), .Z(n36581) );
  AND U45613 ( .A(n36587), .B(n36588), .Z(n36479) );
  NAND U45614 ( .A(n36589), .B(n36590), .Z(n36588) );
  NAND U45615 ( .A(n36591), .B(n36592), .Z(n36587) );
  AND U45616 ( .A(n36593), .B(n36594), .Z(n36481) );
  XOR U45617 ( .A(n36561), .B(n36560), .Z(N62139) );
  XNOR U45618 ( .A(n36578), .B(n36579), .Z(n36560) );
  XNOR U45619 ( .A(n36593), .B(n36594), .Z(n36579) );
  XOR U45620 ( .A(n36590), .B(n36589), .Z(n36594) );
  XOR U45621 ( .A(y[2868]), .B(x[2868]), .Z(n36589) );
  XOR U45622 ( .A(n36592), .B(n36591), .Z(n36590) );
  XOR U45623 ( .A(y[2870]), .B(x[2870]), .Z(n36591) );
  XOR U45624 ( .A(y[2869]), .B(x[2869]), .Z(n36592) );
  XOR U45625 ( .A(n36584), .B(n36583), .Z(n36593) );
  XOR U45626 ( .A(n36586), .B(n36585), .Z(n36583) );
  XOR U45627 ( .A(y[2867]), .B(x[2867]), .Z(n36585) );
  XOR U45628 ( .A(y[2866]), .B(x[2866]), .Z(n36586) );
  XOR U45629 ( .A(y[2865]), .B(x[2865]), .Z(n36584) );
  XNOR U45630 ( .A(n36577), .B(n36576), .Z(n36578) );
  XNOR U45631 ( .A(n36573), .B(n36572), .Z(n36576) );
  XOR U45632 ( .A(n36575), .B(n36574), .Z(n36572) );
  XOR U45633 ( .A(y[2864]), .B(x[2864]), .Z(n36574) );
  XOR U45634 ( .A(y[2863]), .B(x[2863]), .Z(n36575) );
  XOR U45635 ( .A(y[2862]), .B(x[2862]), .Z(n36573) );
  XOR U45636 ( .A(n36567), .B(n36566), .Z(n36577) );
  XOR U45637 ( .A(n36569), .B(n36568), .Z(n36566) );
  XOR U45638 ( .A(y[2861]), .B(x[2861]), .Z(n36568) );
  XOR U45639 ( .A(y[2860]), .B(x[2860]), .Z(n36569) );
  XOR U45640 ( .A(y[2859]), .B(x[2859]), .Z(n36567) );
  XNOR U45641 ( .A(n36543), .B(n36544), .Z(n36561) );
  XNOR U45642 ( .A(n36558), .B(n36559), .Z(n36544) );
  XOR U45643 ( .A(n36555), .B(n36554), .Z(n36559) );
  XOR U45644 ( .A(y[2856]), .B(x[2856]), .Z(n36554) );
  XOR U45645 ( .A(n36557), .B(n36556), .Z(n36555) );
  XOR U45646 ( .A(y[2858]), .B(x[2858]), .Z(n36556) );
  XOR U45647 ( .A(y[2857]), .B(x[2857]), .Z(n36557) );
  XOR U45648 ( .A(n36549), .B(n36548), .Z(n36558) );
  XOR U45649 ( .A(n36551), .B(n36550), .Z(n36548) );
  XOR U45650 ( .A(y[2855]), .B(x[2855]), .Z(n36550) );
  XOR U45651 ( .A(y[2854]), .B(x[2854]), .Z(n36551) );
  XOR U45652 ( .A(y[2853]), .B(x[2853]), .Z(n36549) );
  XNOR U45653 ( .A(n36542), .B(n36541), .Z(n36543) );
  XNOR U45654 ( .A(n36538), .B(n36537), .Z(n36541) );
  XOR U45655 ( .A(n36540), .B(n36539), .Z(n36537) );
  XOR U45656 ( .A(y[2852]), .B(x[2852]), .Z(n36539) );
  XOR U45657 ( .A(y[2851]), .B(x[2851]), .Z(n36540) );
  XOR U45658 ( .A(y[2850]), .B(x[2850]), .Z(n36538) );
  XOR U45659 ( .A(n36532), .B(n36531), .Z(n36542) );
  XOR U45660 ( .A(n36534), .B(n36533), .Z(n36531) );
  XOR U45661 ( .A(y[2849]), .B(x[2849]), .Z(n36533) );
  XOR U45662 ( .A(y[2848]), .B(x[2848]), .Z(n36534) );
  XOR U45663 ( .A(y[2847]), .B(x[2847]), .Z(n36532) );
  NAND U45664 ( .A(n36595), .B(n36596), .Z(N62130) );
  NAND U45665 ( .A(n36597), .B(n36598), .Z(n36596) );
  NANDN U45666 ( .A(n36599), .B(n36600), .Z(n36598) );
  NANDN U45667 ( .A(n36600), .B(n36599), .Z(n36595) );
  XOR U45668 ( .A(n36599), .B(n36601), .Z(N62129) );
  XNOR U45669 ( .A(n36597), .B(n36600), .Z(n36601) );
  NAND U45670 ( .A(n36602), .B(n36603), .Z(n36600) );
  NAND U45671 ( .A(n36604), .B(n36605), .Z(n36603) );
  NANDN U45672 ( .A(n36606), .B(n36607), .Z(n36605) );
  NANDN U45673 ( .A(n36607), .B(n36606), .Z(n36602) );
  AND U45674 ( .A(n36608), .B(n36609), .Z(n36597) );
  NAND U45675 ( .A(n36610), .B(n36611), .Z(n36609) );
  NANDN U45676 ( .A(n36612), .B(n36613), .Z(n36611) );
  NANDN U45677 ( .A(n36613), .B(n36612), .Z(n36608) );
  IV U45678 ( .A(n36614), .Z(n36613) );
  AND U45679 ( .A(n36615), .B(n36616), .Z(n36599) );
  NAND U45680 ( .A(n36617), .B(n36618), .Z(n36616) );
  NANDN U45681 ( .A(n36619), .B(n36620), .Z(n36618) );
  NANDN U45682 ( .A(n36620), .B(n36619), .Z(n36615) );
  XOR U45683 ( .A(n36612), .B(n36621), .Z(N62128) );
  XNOR U45684 ( .A(n36610), .B(n36614), .Z(n36621) );
  XOR U45685 ( .A(n36607), .B(n36622), .Z(n36614) );
  XNOR U45686 ( .A(n36604), .B(n36606), .Z(n36622) );
  AND U45687 ( .A(n36623), .B(n36624), .Z(n36606) );
  NANDN U45688 ( .A(n36625), .B(n36626), .Z(n36624) );
  OR U45689 ( .A(n36627), .B(n36628), .Z(n36626) );
  IV U45690 ( .A(n36629), .Z(n36628) );
  NANDN U45691 ( .A(n36629), .B(n36627), .Z(n36623) );
  AND U45692 ( .A(n36630), .B(n36631), .Z(n36604) );
  NAND U45693 ( .A(n36632), .B(n36633), .Z(n36631) );
  NANDN U45694 ( .A(n36634), .B(n36635), .Z(n36633) );
  NANDN U45695 ( .A(n36635), .B(n36634), .Z(n36630) );
  IV U45696 ( .A(n36636), .Z(n36635) );
  NAND U45697 ( .A(n36637), .B(n36638), .Z(n36607) );
  NANDN U45698 ( .A(n36639), .B(n36640), .Z(n36638) );
  NANDN U45699 ( .A(n36641), .B(n36642), .Z(n36640) );
  NANDN U45700 ( .A(n36642), .B(n36641), .Z(n36637) );
  IV U45701 ( .A(n36643), .Z(n36641) );
  AND U45702 ( .A(n36644), .B(n36645), .Z(n36610) );
  NAND U45703 ( .A(n36646), .B(n36647), .Z(n36645) );
  NANDN U45704 ( .A(n36648), .B(n36649), .Z(n36647) );
  NANDN U45705 ( .A(n36649), .B(n36648), .Z(n36644) );
  XOR U45706 ( .A(n36620), .B(n36650), .Z(n36612) );
  XNOR U45707 ( .A(n36617), .B(n36619), .Z(n36650) );
  AND U45708 ( .A(n36651), .B(n36652), .Z(n36619) );
  NANDN U45709 ( .A(n36653), .B(n36654), .Z(n36652) );
  OR U45710 ( .A(n36655), .B(n36656), .Z(n36654) );
  IV U45711 ( .A(n36657), .Z(n36656) );
  NANDN U45712 ( .A(n36657), .B(n36655), .Z(n36651) );
  AND U45713 ( .A(n36658), .B(n36659), .Z(n36617) );
  NAND U45714 ( .A(n36660), .B(n36661), .Z(n36659) );
  NANDN U45715 ( .A(n36662), .B(n36663), .Z(n36661) );
  NANDN U45716 ( .A(n36663), .B(n36662), .Z(n36658) );
  IV U45717 ( .A(n36664), .Z(n36663) );
  NAND U45718 ( .A(n36665), .B(n36666), .Z(n36620) );
  NANDN U45719 ( .A(n36667), .B(n36668), .Z(n36666) );
  NANDN U45720 ( .A(n36669), .B(n36670), .Z(n36668) );
  NANDN U45721 ( .A(n36670), .B(n36669), .Z(n36665) );
  IV U45722 ( .A(n36671), .Z(n36669) );
  XOR U45723 ( .A(n36646), .B(n36672), .Z(N62127) );
  XNOR U45724 ( .A(n36649), .B(n36648), .Z(n36672) );
  XNOR U45725 ( .A(n36660), .B(n36673), .Z(n36648) );
  XNOR U45726 ( .A(n36664), .B(n36662), .Z(n36673) );
  XOR U45727 ( .A(n36670), .B(n36674), .Z(n36662) );
  XNOR U45728 ( .A(n36667), .B(n36671), .Z(n36674) );
  AND U45729 ( .A(n36675), .B(n36676), .Z(n36671) );
  NAND U45730 ( .A(n36677), .B(n36678), .Z(n36676) );
  NAND U45731 ( .A(n36679), .B(n36680), .Z(n36675) );
  AND U45732 ( .A(n36681), .B(n36682), .Z(n36667) );
  NAND U45733 ( .A(n36683), .B(n36684), .Z(n36682) );
  NAND U45734 ( .A(n36685), .B(n36686), .Z(n36681) );
  NANDN U45735 ( .A(n36687), .B(n36688), .Z(n36670) );
  ANDN U45736 ( .B(n36689), .A(n36690), .Z(n36664) );
  XNOR U45737 ( .A(n36655), .B(n36691), .Z(n36660) );
  XNOR U45738 ( .A(n36653), .B(n36657), .Z(n36691) );
  AND U45739 ( .A(n36692), .B(n36693), .Z(n36657) );
  NAND U45740 ( .A(n36694), .B(n36695), .Z(n36693) );
  NAND U45741 ( .A(n36696), .B(n36697), .Z(n36692) );
  AND U45742 ( .A(n36698), .B(n36699), .Z(n36653) );
  NAND U45743 ( .A(n36700), .B(n36701), .Z(n36699) );
  NAND U45744 ( .A(n36702), .B(n36703), .Z(n36698) );
  AND U45745 ( .A(n36704), .B(n36705), .Z(n36655) );
  NAND U45746 ( .A(n36706), .B(n36707), .Z(n36649) );
  XNOR U45747 ( .A(n36632), .B(n36708), .Z(n36646) );
  XNOR U45748 ( .A(n36636), .B(n36634), .Z(n36708) );
  XOR U45749 ( .A(n36642), .B(n36709), .Z(n36634) );
  XNOR U45750 ( .A(n36639), .B(n36643), .Z(n36709) );
  AND U45751 ( .A(n36710), .B(n36711), .Z(n36643) );
  NAND U45752 ( .A(n36712), .B(n36713), .Z(n36711) );
  NAND U45753 ( .A(n36714), .B(n36715), .Z(n36710) );
  AND U45754 ( .A(n36716), .B(n36717), .Z(n36639) );
  NAND U45755 ( .A(n36718), .B(n36719), .Z(n36717) );
  NAND U45756 ( .A(n36720), .B(n36721), .Z(n36716) );
  NANDN U45757 ( .A(n36722), .B(n36723), .Z(n36642) );
  ANDN U45758 ( .B(n36724), .A(n36725), .Z(n36636) );
  XNOR U45759 ( .A(n36627), .B(n36726), .Z(n36632) );
  XNOR U45760 ( .A(n36625), .B(n36629), .Z(n36726) );
  AND U45761 ( .A(n36727), .B(n36728), .Z(n36629) );
  NAND U45762 ( .A(n36729), .B(n36730), .Z(n36728) );
  NAND U45763 ( .A(n36731), .B(n36732), .Z(n36727) );
  AND U45764 ( .A(n36733), .B(n36734), .Z(n36625) );
  NAND U45765 ( .A(n36735), .B(n36736), .Z(n36734) );
  NAND U45766 ( .A(n36737), .B(n36738), .Z(n36733) );
  AND U45767 ( .A(n36739), .B(n36740), .Z(n36627) );
  XOR U45768 ( .A(n36707), .B(n36706), .Z(N62126) );
  XNOR U45769 ( .A(n36724), .B(n36725), .Z(n36706) );
  XNOR U45770 ( .A(n36739), .B(n36740), .Z(n36725) );
  XOR U45771 ( .A(n36736), .B(n36735), .Z(n36740) );
  XOR U45772 ( .A(y[2844]), .B(x[2844]), .Z(n36735) );
  XOR U45773 ( .A(n36738), .B(n36737), .Z(n36736) );
  XOR U45774 ( .A(y[2846]), .B(x[2846]), .Z(n36737) );
  XOR U45775 ( .A(y[2845]), .B(x[2845]), .Z(n36738) );
  XOR U45776 ( .A(n36730), .B(n36729), .Z(n36739) );
  XOR U45777 ( .A(n36732), .B(n36731), .Z(n36729) );
  XOR U45778 ( .A(y[2843]), .B(x[2843]), .Z(n36731) );
  XOR U45779 ( .A(y[2842]), .B(x[2842]), .Z(n36732) );
  XOR U45780 ( .A(y[2841]), .B(x[2841]), .Z(n36730) );
  XNOR U45781 ( .A(n36723), .B(n36722), .Z(n36724) );
  XNOR U45782 ( .A(n36719), .B(n36718), .Z(n36722) );
  XOR U45783 ( .A(n36721), .B(n36720), .Z(n36718) );
  XOR U45784 ( .A(y[2840]), .B(x[2840]), .Z(n36720) );
  XOR U45785 ( .A(y[2839]), .B(x[2839]), .Z(n36721) );
  XOR U45786 ( .A(y[2838]), .B(x[2838]), .Z(n36719) );
  XOR U45787 ( .A(n36713), .B(n36712), .Z(n36723) );
  XOR U45788 ( .A(n36715), .B(n36714), .Z(n36712) );
  XOR U45789 ( .A(y[2837]), .B(x[2837]), .Z(n36714) );
  XOR U45790 ( .A(y[2836]), .B(x[2836]), .Z(n36715) );
  XOR U45791 ( .A(y[2835]), .B(x[2835]), .Z(n36713) );
  XNOR U45792 ( .A(n36689), .B(n36690), .Z(n36707) );
  XNOR U45793 ( .A(n36704), .B(n36705), .Z(n36690) );
  XOR U45794 ( .A(n36701), .B(n36700), .Z(n36705) );
  XOR U45795 ( .A(y[2832]), .B(x[2832]), .Z(n36700) );
  XOR U45796 ( .A(n36703), .B(n36702), .Z(n36701) );
  XOR U45797 ( .A(y[2834]), .B(x[2834]), .Z(n36702) );
  XOR U45798 ( .A(y[2833]), .B(x[2833]), .Z(n36703) );
  XOR U45799 ( .A(n36695), .B(n36694), .Z(n36704) );
  XOR U45800 ( .A(n36697), .B(n36696), .Z(n36694) );
  XOR U45801 ( .A(y[2831]), .B(x[2831]), .Z(n36696) );
  XOR U45802 ( .A(y[2830]), .B(x[2830]), .Z(n36697) );
  XOR U45803 ( .A(y[2829]), .B(x[2829]), .Z(n36695) );
  XNOR U45804 ( .A(n36688), .B(n36687), .Z(n36689) );
  XNOR U45805 ( .A(n36684), .B(n36683), .Z(n36687) );
  XOR U45806 ( .A(n36686), .B(n36685), .Z(n36683) );
  XOR U45807 ( .A(y[2828]), .B(x[2828]), .Z(n36685) );
  XOR U45808 ( .A(y[2827]), .B(x[2827]), .Z(n36686) );
  XOR U45809 ( .A(y[2826]), .B(x[2826]), .Z(n36684) );
  XOR U45810 ( .A(n36678), .B(n36677), .Z(n36688) );
  XOR U45811 ( .A(n36680), .B(n36679), .Z(n36677) );
  XOR U45812 ( .A(y[2825]), .B(x[2825]), .Z(n36679) );
  XOR U45813 ( .A(y[2824]), .B(x[2824]), .Z(n36680) );
  XOR U45814 ( .A(y[2823]), .B(x[2823]), .Z(n36678) );
  NAND U45815 ( .A(n36741), .B(n36742), .Z(N62117) );
  NAND U45816 ( .A(n36743), .B(n36744), .Z(n36742) );
  NANDN U45817 ( .A(n36745), .B(n36746), .Z(n36744) );
  NANDN U45818 ( .A(n36746), .B(n36745), .Z(n36741) );
  XOR U45819 ( .A(n36745), .B(n36747), .Z(N62116) );
  XNOR U45820 ( .A(n36743), .B(n36746), .Z(n36747) );
  NAND U45821 ( .A(n36748), .B(n36749), .Z(n36746) );
  NAND U45822 ( .A(n36750), .B(n36751), .Z(n36749) );
  NANDN U45823 ( .A(n36752), .B(n36753), .Z(n36751) );
  NANDN U45824 ( .A(n36753), .B(n36752), .Z(n36748) );
  AND U45825 ( .A(n36754), .B(n36755), .Z(n36743) );
  NAND U45826 ( .A(n36756), .B(n36757), .Z(n36755) );
  NANDN U45827 ( .A(n36758), .B(n36759), .Z(n36757) );
  NANDN U45828 ( .A(n36759), .B(n36758), .Z(n36754) );
  IV U45829 ( .A(n36760), .Z(n36759) );
  AND U45830 ( .A(n36761), .B(n36762), .Z(n36745) );
  NAND U45831 ( .A(n36763), .B(n36764), .Z(n36762) );
  NANDN U45832 ( .A(n36765), .B(n36766), .Z(n36764) );
  NANDN U45833 ( .A(n36766), .B(n36765), .Z(n36761) );
  XOR U45834 ( .A(n36758), .B(n36767), .Z(N62115) );
  XNOR U45835 ( .A(n36756), .B(n36760), .Z(n36767) );
  XOR U45836 ( .A(n36753), .B(n36768), .Z(n36760) );
  XNOR U45837 ( .A(n36750), .B(n36752), .Z(n36768) );
  AND U45838 ( .A(n36769), .B(n36770), .Z(n36752) );
  NANDN U45839 ( .A(n36771), .B(n36772), .Z(n36770) );
  OR U45840 ( .A(n36773), .B(n36774), .Z(n36772) );
  IV U45841 ( .A(n36775), .Z(n36774) );
  NANDN U45842 ( .A(n36775), .B(n36773), .Z(n36769) );
  AND U45843 ( .A(n36776), .B(n36777), .Z(n36750) );
  NAND U45844 ( .A(n36778), .B(n36779), .Z(n36777) );
  NANDN U45845 ( .A(n36780), .B(n36781), .Z(n36779) );
  NANDN U45846 ( .A(n36781), .B(n36780), .Z(n36776) );
  IV U45847 ( .A(n36782), .Z(n36781) );
  NAND U45848 ( .A(n36783), .B(n36784), .Z(n36753) );
  NANDN U45849 ( .A(n36785), .B(n36786), .Z(n36784) );
  NANDN U45850 ( .A(n36787), .B(n36788), .Z(n36786) );
  NANDN U45851 ( .A(n36788), .B(n36787), .Z(n36783) );
  IV U45852 ( .A(n36789), .Z(n36787) );
  AND U45853 ( .A(n36790), .B(n36791), .Z(n36756) );
  NAND U45854 ( .A(n36792), .B(n36793), .Z(n36791) );
  NANDN U45855 ( .A(n36794), .B(n36795), .Z(n36793) );
  NANDN U45856 ( .A(n36795), .B(n36794), .Z(n36790) );
  XOR U45857 ( .A(n36766), .B(n36796), .Z(n36758) );
  XNOR U45858 ( .A(n36763), .B(n36765), .Z(n36796) );
  AND U45859 ( .A(n36797), .B(n36798), .Z(n36765) );
  NANDN U45860 ( .A(n36799), .B(n36800), .Z(n36798) );
  OR U45861 ( .A(n36801), .B(n36802), .Z(n36800) );
  IV U45862 ( .A(n36803), .Z(n36802) );
  NANDN U45863 ( .A(n36803), .B(n36801), .Z(n36797) );
  AND U45864 ( .A(n36804), .B(n36805), .Z(n36763) );
  NAND U45865 ( .A(n36806), .B(n36807), .Z(n36805) );
  NANDN U45866 ( .A(n36808), .B(n36809), .Z(n36807) );
  NANDN U45867 ( .A(n36809), .B(n36808), .Z(n36804) );
  IV U45868 ( .A(n36810), .Z(n36809) );
  NAND U45869 ( .A(n36811), .B(n36812), .Z(n36766) );
  NANDN U45870 ( .A(n36813), .B(n36814), .Z(n36812) );
  NANDN U45871 ( .A(n36815), .B(n36816), .Z(n36814) );
  NANDN U45872 ( .A(n36816), .B(n36815), .Z(n36811) );
  IV U45873 ( .A(n36817), .Z(n36815) );
  XOR U45874 ( .A(n36792), .B(n36818), .Z(N62114) );
  XNOR U45875 ( .A(n36795), .B(n36794), .Z(n36818) );
  XNOR U45876 ( .A(n36806), .B(n36819), .Z(n36794) );
  XNOR U45877 ( .A(n36810), .B(n36808), .Z(n36819) );
  XOR U45878 ( .A(n36816), .B(n36820), .Z(n36808) );
  XNOR U45879 ( .A(n36813), .B(n36817), .Z(n36820) );
  AND U45880 ( .A(n36821), .B(n36822), .Z(n36817) );
  NAND U45881 ( .A(n36823), .B(n36824), .Z(n36822) );
  NAND U45882 ( .A(n36825), .B(n36826), .Z(n36821) );
  AND U45883 ( .A(n36827), .B(n36828), .Z(n36813) );
  NAND U45884 ( .A(n36829), .B(n36830), .Z(n36828) );
  NAND U45885 ( .A(n36831), .B(n36832), .Z(n36827) );
  NANDN U45886 ( .A(n36833), .B(n36834), .Z(n36816) );
  ANDN U45887 ( .B(n36835), .A(n36836), .Z(n36810) );
  XNOR U45888 ( .A(n36801), .B(n36837), .Z(n36806) );
  XNOR U45889 ( .A(n36799), .B(n36803), .Z(n36837) );
  AND U45890 ( .A(n36838), .B(n36839), .Z(n36803) );
  NAND U45891 ( .A(n36840), .B(n36841), .Z(n36839) );
  NAND U45892 ( .A(n36842), .B(n36843), .Z(n36838) );
  AND U45893 ( .A(n36844), .B(n36845), .Z(n36799) );
  NAND U45894 ( .A(n36846), .B(n36847), .Z(n36845) );
  NAND U45895 ( .A(n36848), .B(n36849), .Z(n36844) );
  AND U45896 ( .A(n36850), .B(n36851), .Z(n36801) );
  NAND U45897 ( .A(n36852), .B(n36853), .Z(n36795) );
  XNOR U45898 ( .A(n36778), .B(n36854), .Z(n36792) );
  XNOR U45899 ( .A(n36782), .B(n36780), .Z(n36854) );
  XOR U45900 ( .A(n36788), .B(n36855), .Z(n36780) );
  XNOR U45901 ( .A(n36785), .B(n36789), .Z(n36855) );
  AND U45902 ( .A(n36856), .B(n36857), .Z(n36789) );
  NAND U45903 ( .A(n36858), .B(n36859), .Z(n36857) );
  NAND U45904 ( .A(n36860), .B(n36861), .Z(n36856) );
  AND U45905 ( .A(n36862), .B(n36863), .Z(n36785) );
  NAND U45906 ( .A(n36864), .B(n36865), .Z(n36863) );
  NAND U45907 ( .A(n36866), .B(n36867), .Z(n36862) );
  NANDN U45908 ( .A(n36868), .B(n36869), .Z(n36788) );
  ANDN U45909 ( .B(n36870), .A(n36871), .Z(n36782) );
  XNOR U45910 ( .A(n36773), .B(n36872), .Z(n36778) );
  XNOR U45911 ( .A(n36771), .B(n36775), .Z(n36872) );
  AND U45912 ( .A(n36873), .B(n36874), .Z(n36775) );
  NAND U45913 ( .A(n36875), .B(n36876), .Z(n36874) );
  NAND U45914 ( .A(n36877), .B(n36878), .Z(n36873) );
  AND U45915 ( .A(n36879), .B(n36880), .Z(n36771) );
  NAND U45916 ( .A(n36881), .B(n36882), .Z(n36880) );
  NAND U45917 ( .A(n36883), .B(n36884), .Z(n36879) );
  AND U45918 ( .A(n36885), .B(n36886), .Z(n36773) );
  XOR U45919 ( .A(n36853), .B(n36852), .Z(N62113) );
  XNOR U45920 ( .A(n36870), .B(n36871), .Z(n36852) );
  XNOR U45921 ( .A(n36885), .B(n36886), .Z(n36871) );
  XOR U45922 ( .A(n36882), .B(n36881), .Z(n36886) );
  XOR U45923 ( .A(y[2820]), .B(x[2820]), .Z(n36881) );
  XOR U45924 ( .A(n36884), .B(n36883), .Z(n36882) );
  XOR U45925 ( .A(y[2822]), .B(x[2822]), .Z(n36883) );
  XOR U45926 ( .A(y[2821]), .B(x[2821]), .Z(n36884) );
  XOR U45927 ( .A(n36876), .B(n36875), .Z(n36885) );
  XOR U45928 ( .A(n36878), .B(n36877), .Z(n36875) );
  XOR U45929 ( .A(y[2819]), .B(x[2819]), .Z(n36877) );
  XOR U45930 ( .A(y[2818]), .B(x[2818]), .Z(n36878) );
  XOR U45931 ( .A(y[2817]), .B(x[2817]), .Z(n36876) );
  XNOR U45932 ( .A(n36869), .B(n36868), .Z(n36870) );
  XNOR U45933 ( .A(n36865), .B(n36864), .Z(n36868) );
  XOR U45934 ( .A(n36867), .B(n36866), .Z(n36864) );
  XOR U45935 ( .A(y[2816]), .B(x[2816]), .Z(n36866) );
  XOR U45936 ( .A(y[2815]), .B(x[2815]), .Z(n36867) );
  XOR U45937 ( .A(y[2814]), .B(x[2814]), .Z(n36865) );
  XOR U45938 ( .A(n36859), .B(n36858), .Z(n36869) );
  XOR U45939 ( .A(n36861), .B(n36860), .Z(n36858) );
  XOR U45940 ( .A(y[2813]), .B(x[2813]), .Z(n36860) );
  XOR U45941 ( .A(y[2812]), .B(x[2812]), .Z(n36861) );
  XOR U45942 ( .A(y[2811]), .B(x[2811]), .Z(n36859) );
  XNOR U45943 ( .A(n36835), .B(n36836), .Z(n36853) );
  XNOR U45944 ( .A(n36850), .B(n36851), .Z(n36836) );
  XOR U45945 ( .A(n36847), .B(n36846), .Z(n36851) );
  XOR U45946 ( .A(y[2808]), .B(x[2808]), .Z(n36846) );
  XOR U45947 ( .A(n36849), .B(n36848), .Z(n36847) );
  XOR U45948 ( .A(y[2810]), .B(x[2810]), .Z(n36848) );
  XOR U45949 ( .A(y[2809]), .B(x[2809]), .Z(n36849) );
  XOR U45950 ( .A(n36841), .B(n36840), .Z(n36850) );
  XOR U45951 ( .A(n36843), .B(n36842), .Z(n36840) );
  XOR U45952 ( .A(y[2807]), .B(x[2807]), .Z(n36842) );
  XOR U45953 ( .A(y[2806]), .B(x[2806]), .Z(n36843) );
  XOR U45954 ( .A(y[2805]), .B(x[2805]), .Z(n36841) );
  XNOR U45955 ( .A(n36834), .B(n36833), .Z(n36835) );
  XNOR U45956 ( .A(n36830), .B(n36829), .Z(n36833) );
  XOR U45957 ( .A(n36832), .B(n36831), .Z(n36829) );
  XOR U45958 ( .A(y[2804]), .B(x[2804]), .Z(n36831) );
  XOR U45959 ( .A(y[2803]), .B(x[2803]), .Z(n36832) );
  XOR U45960 ( .A(y[2802]), .B(x[2802]), .Z(n36830) );
  XOR U45961 ( .A(n36824), .B(n36823), .Z(n36834) );
  XOR U45962 ( .A(n36826), .B(n36825), .Z(n36823) );
  XOR U45963 ( .A(y[2801]), .B(x[2801]), .Z(n36825) );
  XOR U45964 ( .A(y[2800]), .B(x[2800]), .Z(n36826) );
  XOR U45965 ( .A(y[2799]), .B(x[2799]), .Z(n36824) );
  NAND U45966 ( .A(n36887), .B(n36888), .Z(N62104) );
  NAND U45967 ( .A(n36889), .B(n36890), .Z(n36888) );
  NANDN U45968 ( .A(n36891), .B(n36892), .Z(n36890) );
  NANDN U45969 ( .A(n36892), .B(n36891), .Z(n36887) );
  XOR U45970 ( .A(n36891), .B(n36893), .Z(N62103) );
  XNOR U45971 ( .A(n36889), .B(n36892), .Z(n36893) );
  NAND U45972 ( .A(n36894), .B(n36895), .Z(n36892) );
  NAND U45973 ( .A(n36896), .B(n36897), .Z(n36895) );
  NANDN U45974 ( .A(n36898), .B(n36899), .Z(n36897) );
  NANDN U45975 ( .A(n36899), .B(n36898), .Z(n36894) );
  AND U45976 ( .A(n36900), .B(n36901), .Z(n36889) );
  NAND U45977 ( .A(n36902), .B(n36903), .Z(n36901) );
  NANDN U45978 ( .A(n36904), .B(n36905), .Z(n36903) );
  NANDN U45979 ( .A(n36905), .B(n36904), .Z(n36900) );
  IV U45980 ( .A(n36906), .Z(n36905) );
  AND U45981 ( .A(n36907), .B(n36908), .Z(n36891) );
  NAND U45982 ( .A(n36909), .B(n36910), .Z(n36908) );
  NANDN U45983 ( .A(n36911), .B(n36912), .Z(n36910) );
  NANDN U45984 ( .A(n36912), .B(n36911), .Z(n36907) );
  XOR U45985 ( .A(n36904), .B(n36913), .Z(N62102) );
  XNOR U45986 ( .A(n36902), .B(n36906), .Z(n36913) );
  XOR U45987 ( .A(n36899), .B(n36914), .Z(n36906) );
  XNOR U45988 ( .A(n36896), .B(n36898), .Z(n36914) );
  AND U45989 ( .A(n36915), .B(n36916), .Z(n36898) );
  NANDN U45990 ( .A(n36917), .B(n36918), .Z(n36916) );
  OR U45991 ( .A(n36919), .B(n36920), .Z(n36918) );
  IV U45992 ( .A(n36921), .Z(n36920) );
  NANDN U45993 ( .A(n36921), .B(n36919), .Z(n36915) );
  AND U45994 ( .A(n36922), .B(n36923), .Z(n36896) );
  NAND U45995 ( .A(n36924), .B(n36925), .Z(n36923) );
  NANDN U45996 ( .A(n36926), .B(n36927), .Z(n36925) );
  NANDN U45997 ( .A(n36927), .B(n36926), .Z(n36922) );
  IV U45998 ( .A(n36928), .Z(n36927) );
  NAND U45999 ( .A(n36929), .B(n36930), .Z(n36899) );
  NANDN U46000 ( .A(n36931), .B(n36932), .Z(n36930) );
  NANDN U46001 ( .A(n36933), .B(n36934), .Z(n36932) );
  NANDN U46002 ( .A(n36934), .B(n36933), .Z(n36929) );
  IV U46003 ( .A(n36935), .Z(n36933) );
  AND U46004 ( .A(n36936), .B(n36937), .Z(n36902) );
  NAND U46005 ( .A(n36938), .B(n36939), .Z(n36937) );
  NANDN U46006 ( .A(n36940), .B(n36941), .Z(n36939) );
  NANDN U46007 ( .A(n36941), .B(n36940), .Z(n36936) );
  XOR U46008 ( .A(n36912), .B(n36942), .Z(n36904) );
  XNOR U46009 ( .A(n36909), .B(n36911), .Z(n36942) );
  AND U46010 ( .A(n36943), .B(n36944), .Z(n36911) );
  NANDN U46011 ( .A(n36945), .B(n36946), .Z(n36944) );
  OR U46012 ( .A(n36947), .B(n36948), .Z(n36946) );
  IV U46013 ( .A(n36949), .Z(n36948) );
  NANDN U46014 ( .A(n36949), .B(n36947), .Z(n36943) );
  AND U46015 ( .A(n36950), .B(n36951), .Z(n36909) );
  NAND U46016 ( .A(n36952), .B(n36953), .Z(n36951) );
  NANDN U46017 ( .A(n36954), .B(n36955), .Z(n36953) );
  NANDN U46018 ( .A(n36955), .B(n36954), .Z(n36950) );
  IV U46019 ( .A(n36956), .Z(n36955) );
  NAND U46020 ( .A(n36957), .B(n36958), .Z(n36912) );
  NANDN U46021 ( .A(n36959), .B(n36960), .Z(n36958) );
  NANDN U46022 ( .A(n36961), .B(n36962), .Z(n36960) );
  NANDN U46023 ( .A(n36962), .B(n36961), .Z(n36957) );
  IV U46024 ( .A(n36963), .Z(n36961) );
  XOR U46025 ( .A(n36938), .B(n36964), .Z(N62101) );
  XNOR U46026 ( .A(n36941), .B(n36940), .Z(n36964) );
  XNOR U46027 ( .A(n36952), .B(n36965), .Z(n36940) );
  XNOR U46028 ( .A(n36956), .B(n36954), .Z(n36965) );
  XOR U46029 ( .A(n36962), .B(n36966), .Z(n36954) );
  XNOR U46030 ( .A(n36959), .B(n36963), .Z(n36966) );
  AND U46031 ( .A(n36967), .B(n36968), .Z(n36963) );
  NAND U46032 ( .A(n36969), .B(n36970), .Z(n36968) );
  NAND U46033 ( .A(n36971), .B(n36972), .Z(n36967) );
  AND U46034 ( .A(n36973), .B(n36974), .Z(n36959) );
  NAND U46035 ( .A(n36975), .B(n36976), .Z(n36974) );
  NAND U46036 ( .A(n36977), .B(n36978), .Z(n36973) );
  NANDN U46037 ( .A(n36979), .B(n36980), .Z(n36962) );
  ANDN U46038 ( .B(n36981), .A(n36982), .Z(n36956) );
  XNOR U46039 ( .A(n36947), .B(n36983), .Z(n36952) );
  XNOR U46040 ( .A(n36945), .B(n36949), .Z(n36983) );
  AND U46041 ( .A(n36984), .B(n36985), .Z(n36949) );
  NAND U46042 ( .A(n36986), .B(n36987), .Z(n36985) );
  NAND U46043 ( .A(n36988), .B(n36989), .Z(n36984) );
  AND U46044 ( .A(n36990), .B(n36991), .Z(n36945) );
  NAND U46045 ( .A(n36992), .B(n36993), .Z(n36991) );
  NAND U46046 ( .A(n36994), .B(n36995), .Z(n36990) );
  AND U46047 ( .A(n36996), .B(n36997), .Z(n36947) );
  NAND U46048 ( .A(n36998), .B(n36999), .Z(n36941) );
  XNOR U46049 ( .A(n36924), .B(n37000), .Z(n36938) );
  XNOR U46050 ( .A(n36928), .B(n36926), .Z(n37000) );
  XOR U46051 ( .A(n36934), .B(n37001), .Z(n36926) );
  XNOR U46052 ( .A(n36931), .B(n36935), .Z(n37001) );
  AND U46053 ( .A(n37002), .B(n37003), .Z(n36935) );
  NAND U46054 ( .A(n37004), .B(n37005), .Z(n37003) );
  NAND U46055 ( .A(n37006), .B(n37007), .Z(n37002) );
  AND U46056 ( .A(n37008), .B(n37009), .Z(n36931) );
  NAND U46057 ( .A(n37010), .B(n37011), .Z(n37009) );
  NAND U46058 ( .A(n37012), .B(n37013), .Z(n37008) );
  NANDN U46059 ( .A(n37014), .B(n37015), .Z(n36934) );
  ANDN U46060 ( .B(n37016), .A(n37017), .Z(n36928) );
  XNOR U46061 ( .A(n36919), .B(n37018), .Z(n36924) );
  XNOR U46062 ( .A(n36917), .B(n36921), .Z(n37018) );
  AND U46063 ( .A(n37019), .B(n37020), .Z(n36921) );
  NAND U46064 ( .A(n37021), .B(n37022), .Z(n37020) );
  NAND U46065 ( .A(n37023), .B(n37024), .Z(n37019) );
  AND U46066 ( .A(n37025), .B(n37026), .Z(n36917) );
  NAND U46067 ( .A(n37027), .B(n37028), .Z(n37026) );
  NAND U46068 ( .A(n37029), .B(n37030), .Z(n37025) );
  AND U46069 ( .A(n37031), .B(n37032), .Z(n36919) );
  XOR U46070 ( .A(n36999), .B(n36998), .Z(N62100) );
  XNOR U46071 ( .A(n37016), .B(n37017), .Z(n36998) );
  XNOR U46072 ( .A(n37031), .B(n37032), .Z(n37017) );
  XOR U46073 ( .A(n37028), .B(n37027), .Z(n37032) );
  XOR U46074 ( .A(y[2796]), .B(x[2796]), .Z(n37027) );
  XOR U46075 ( .A(n37030), .B(n37029), .Z(n37028) );
  XOR U46076 ( .A(y[2798]), .B(x[2798]), .Z(n37029) );
  XOR U46077 ( .A(y[2797]), .B(x[2797]), .Z(n37030) );
  XOR U46078 ( .A(n37022), .B(n37021), .Z(n37031) );
  XOR U46079 ( .A(n37024), .B(n37023), .Z(n37021) );
  XOR U46080 ( .A(y[2795]), .B(x[2795]), .Z(n37023) );
  XOR U46081 ( .A(y[2794]), .B(x[2794]), .Z(n37024) );
  XOR U46082 ( .A(y[2793]), .B(x[2793]), .Z(n37022) );
  XNOR U46083 ( .A(n37015), .B(n37014), .Z(n37016) );
  XNOR U46084 ( .A(n37011), .B(n37010), .Z(n37014) );
  XOR U46085 ( .A(n37013), .B(n37012), .Z(n37010) );
  XOR U46086 ( .A(y[2792]), .B(x[2792]), .Z(n37012) );
  XOR U46087 ( .A(y[2791]), .B(x[2791]), .Z(n37013) );
  XOR U46088 ( .A(y[2790]), .B(x[2790]), .Z(n37011) );
  XOR U46089 ( .A(n37005), .B(n37004), .Z(n37015) );
  XOR U46090 ( .A(n37007), .B(n37006), .Z(n37004) );
  XOR U46091 ( .A(y[2789]), .B(x[2789]), .Z(n37006) );
  XOR U46092 ( .A(y[2788]), .B(x[2788]), .Z(n37007) );
  XOR U46093 ( .A(y[2787]), .B(x[2787]), .Z(n37005) );
  XNOR U46094 ( .A(n36981), .B(n36982), .Z(n36999) );
  XNOR U46095 ( .A(n36996), .B(n36997), .Z(n36982) );
  XOR U46096 ( .A(n36993), .B(n36992), .Z(n36997) );
  XOR U46097 ( .A(y[2784]), .B(x[2784]), .Z(n36992) );
  XOR U46098 ( .A(n36995), .B(n36994), .Z(n36993) );
  XOR U46099 ( .A(y[2786]), .B(x[2786]), .Z(n36994) );
  XOR U46100 ( .A(y[2785]), .B(x[2785]), .Z(n36995) );
  XOR U46101 ( .A(n36987), .B(n36986), .Z(n36996) );
  XOR U46102 ( .A(n36989), .B(n36988), .Z(n36986) );
  XOR U46103 ( .A(y[2783]), .B(x[2783]), .Z(n36988) );
  XOR U46104 ( .A(y[2782]), .B(x[2782]), .Z(n36989) );
  XOR U46105 ( .A(y[2781]), .B(x[2781]), .Z(n36987) );
  XNOR U46106 ( .A(n36980), .B(n36979), .Z(n36981) );
  XNOR U46107 ( .A(n36976), .B(n36975), .Z(n36979) );
  XOR U46108 ( .A(n36978), .B(n36977), .Z(n36975) );
  XOR U46109 ( .A(y[2780]), .B(x[2780]), .Z(n36977) );
  XOR U46110 ( .A(y[2779]), .B(x[2779]), .Z(n36978) );
  XOR U46111 ( .A(y[2778]), .B(x[2778]), .Z(n36976) );
  XOR U46112 ( .A(n36970), .B(n36969), .Z(n36980) );
  XOR U46113 ( .A(n36972), .B(n36971), .Z(n36969) );
  XOR U46114 ( .A(y[2777]), .B(x[2777]), .Z(n36971) );
  XOR U46115 ( .A(y[2776]), .B(x[2776]), .Z(n36972) );
  XOR U46116 ( .A(y[2775]), .B(x[2775]), .Z(n36970) );
  NAND U46117 ( .A(n37033), .B(n37034), .Z(N62091) );
  NAND U46118 ( .A(n37035), .B(n37036), .Z(n37034) );
  NANDN U46119 ( .A(n37037), .B(n37038), .Z(n37036) );
  NANDN U46120 ( .A(n37038), .B(n37037), .Z(n37033) );
  XOR U46121 ( .A(n37037), .B(n37039), .Z(N62090) );
  XNOR U46122 ( .A(n37035), .B(n37038), .Z(n37039) );
  NAND U46123 ( .A(n37040), .B(n37041), .Z(n37038) );
  NAND U46124 ( .A(n37042), .B(n37043), .Z(n37041) );
  NANDN U46125 ( .A(n37044), .B(n37045), .Z(n37043) );
  NANDN U46126 ( .A(n37045), .B(n37044), .Z(n37040) );
  AND U46127 ( .A(n37046), .B(n37047), .Z(n37035) );
  NAND U46128 ( .A(n37048), .B(n37049), .Z(n37047) );
  NANDN U46129 ( .A(n37050), .B(n37051), .Z(n37049) );
  NANDN U46130 ( .A(n37051), .B(n37050), .Z(n37046) );
  IV U46131 ( .A(n37052), .Z(n37051) );
  AND U46132 ( .A(n37053), .B(n37054), .Z(n37037) );
  NAND U46133 ( .A(n37055), .B(n37056), .Z(n37054) );
  NANDN U46134 ( .A(n37057), .B(n37058), .Z(n37056) );
  NANDN U46135 ( .A(n37058), .B(n37057), .Z(n37053) );
  XOR U46136 ( .A(n37050), .B(n37059), .Z(N62089) );
  XNOR U46137 ( .A(n37048), .B(n37052), .Z(n37059) );
  XOR U46138 ( .A(n37045), .B(n37060), .Z(n37052) );
  XNOR U46139 ( .A(n37042), .B(n37044), .Z(n37060) );
  AND U46140 ( .A(n37061), .B(n37062), .Z(n37044) );
  NANDN U46141 ( .A(n37063), .B(n37064), .Z(n37062) );
  OR U46142 ( .A(n37065), .B(n37066), .Z(n37064) );
  IV U46143 ( .A(n37067), .Z(n37066) );
  NANDN U46144 ( .A(n37067), .B(n37065), .Z(n37061) );
  AND U46145 ( .A(n37068), .B(n37069), .Z(n37042) );
  NAND U46146 ( .A(n37070), .B(n37071), .Z(n37069) );
  NANDN U46147 ( .A(n37072), .B(n37073), .Z(n37071) );
  NANDN U46148 ( .A(n37073), .B(n37072), .Z(n37068) );
  IV U46149 ( .A(n37074), .Z(n37073) );
  NAND U46150 ( .A(n37075), .B(n37076), .Z(n37045) );
  NANDN U46151 ( .A(n37077), .B(n37078), .Z(n37076) );
  NANDN U46152 ( .A(n37079), .B(n37080), .Z(n37078) );
  NANDN U46153 ( .A(n37080), .B(n37079), .Z(n37075) );
  IV U46154 ( .A(n37081), .Z(n37079) );
  AND U46155 ( .A(n37082), .B(n37083), .Z(n37048) );
  NAND U46156 ( .A(n37084), .B(n37085), .Z(n37083) );
  NANDN U46157 ( .A(n37086), .B(n37087), .Z(n37085) );
  NANDN U46158 ( .A(n37087), .B(n37086), .Z(n37082) );
  XOR U46159 ( .A(n37058), .B(n37088), .Z(n37050) );
  XNOR U46160 ( .A(n37055), .B(n37057), .Z(n37088) );
  AND U46161 ( .A(n37089), .B(n37090), .Z(n37057) );
  NANDN U46162 ( .A(n37091), .B(n37092), .Z(n37090) );
  OR U46163 ( .A(n37093), .B(n37094), .Z(n37092) );
  IV U46164 ( .A(n37095), .Z(n37094) );
  NANDN U46165 ( .A(n37095), .B(n37093), .Z(n37089) );
  AND U46166 ( .A(n37096), .B(n37097), .Z(n37055) );
  NAND U46167 ( .A(n37098), .B(n37099), .Z(n37097) );
  NANDN U46168 ( .A(n37100), .B(n37101), .Z(n37099) );
  NANDN U46169 ( .A(n37101), .B(n37100), .Z(n37096) );
  IV U46170 ( .A(n37102), .Z(n37101) );
  NAND U46171 ( .A(n37103), .B(n37104), .Z(n37058) );
  NANDN U46172 ( .A(n37105), .B(n37106), .Z(n37104) );
  NANDN U46173 ( .A(n37107), .B(n37108), .Z(n37106) );
  NANDN U46174 ( .A(n37108), .B(n37107), .Z(n37103) );
  IV U46175 ( .A(n37109), .Z(n37107) );
  XOR U46176 ( .A(n37084), .B(n37110), .Z(N62088) );
  XNOR U46177 ( .A(n37087), .B(n37086), .Z(n37110) );
  XNOR U46178 ( .A(n37098), .B(n37111), .Z(n37086) );
  XNOR U46179 ( .A(n37102), .B(n37100), .Z(n37111) );
  XOR U46180 ( .A(n37108), .B(n37112), .Z(n37100) );
  XNOR U46181 ( .A(n37105), .B(n37109), .Z(n37112) );
  AND U46182 ( .A(n37113), .B(n37114), .Z(n37109) );
  NAND U46183 ( .A(n37115), .B(n37116), .Z(n37114) );
  NAND U46184 ( .A(n37117), .B(n37118), .Z(n37113) );
  AND U46185 ( .A(n37119), .B(n37120), .Z(n37105) );
  NAND U46186 ( .A(n37121), .B(n37122), .Z(n37120) );
  NAND U46187 ( .A(n37123), .B(n37124), .Z(n37119) );
  NANDN U46188 ( .A(n37125), .B(n37126), .Z(n37108) );
  ANDN U46189 ( .B(n37127), .A(n37128), .Z(n37102) );
  XNOR U46190 ( .A(n37093), .B(n37129), .Z(n37098) );
  XNOR U46191 ( .A(n37091), .B(n37095), .Z(n37129) );
  AND U46192 ( .A(n37130), .B(n37131), .Z(n37095) );
  NAND U46193 ( .A(n37132), .B(n37133), .Z(n37131) );
  NAND U46194 ( .A(n37134), .B(n37135), .Z(n37130) );
  AND U46195 ( .A(n37136), .B(n37137), .Z(n37091) );
  NAND U46196 ( .A(n37138), .B(n37139), .Z(n37137) );
  NAND U46197 ( .A(n37140), .B(n37141), .Z(n37136) );
  AND U46198 ( .A(n37142), .B(n37143), .Z(n37093) );
  NAND U46199 ( .A(n37144), .B(n37145), .Z(n37087) );
  XNOR U46200 ( .A(n37070), .B(n37146), .Z(n37084) );
  XNOR U46201 ( .A(n37074), .B(n37072), .Z(n37146) );
  XOR U46202 ( .A(n37080), .B(n37147), .Z(n37072) );
  XNOR U46203 ( .A(n37077), .B(n37081), .Z(n37147) );
  AND U46204 ( .A(n37148), .B(n37149), .Z(n37081) );
  NAND U46205 ( .A(n37150), .B(n37151), .Z(n37149) );
  NAND U46206 ( .A(n37152), .B(n37153), .Z(n37148) );
  AND U46207 ( .A(n37154), .B(n37155), .Z(n37077) );
  NAND U46208 ( .A(n37156), .B(n37157), .Z(n37155) );
  NAND U46209 ( .A(n37158), .B(n37159), .Z(n37154) );
  NANDN U46210 ( .A(n37160), .B(n37161), .Z(n37080) );
  ANDN U46211 ( .B(n37162), .A(n37163), .Z(n37074) );
  XNOR U46212 ( .A(n37065), .B(n37164), .Z(n37070) );
  XNOR U46213 ( .A(n37063), .B(n37067), .Z(n37164) );
  AND U46214 ( .A(n37165), .B(n37166), .Z(n37067) );
  NAND U46215 ( .A(n37167), .B(n37168), .Z(n37166) );
  NAND U46216 ( .A(n37169), .B(n37170), .Z(n37165) );
  AND U46217 ( .A(n37171), .B(n37172), .Z(n37063) );
  NAND U46218 ( .A(n37173), .B(n37174), .Z(n37172) );
  NAND U46219 ( .A(n37175), .B(n37176), .Z(n37171) );
  AND U46220 ( .A(n37177), .B(n37178), .Z(n37065) );
  XOR U46221 ( .A(n37145), .B(n37144), .Z(N62087) );
  XNOR U46222 ( .A(n37162), .B(n37163), .Z(n37144) );
  XNOR U46223 ( .A(n37177), .B(n37178), .Z(n37163) );
  XOR U46224 ( .A(n37174), .B(n37173), .Z(n37178) );
  XOR U46225 ( .A(y[2772]), .B(x[2772]), .Z(n37173) );
  XOR U46226 ( .A(n37176), .B(n37175), .Z(n37174) );
  XOR U46227 ( .A(y[2774]), .B(x[2774]), .Z(n37175) );
  XOR U46228 ( .A(y[2773]), .B(x[2773]), .Z(n37176) );
  XOR U46229 ( .A(n37168), .B(n37167), .Z(n37177) );
  XOR U46230 ( .A(n37170), .B(n37169), .Z(n37167) );
  XOR U46231 ( .A(y[2771]), .B(x[2771]), .Z(n37169) );
  XOR U46232 ( .A(y[2770]), .B(x[2770]), .Z(n37170) );
  XOR U46233 ( .A(y[2769]), .B(x[2769]), .Z(n37168) );
  XNOR U46234 ( .A(n37161), .B(n37160), .Z(n37162) );
  XNOR U46235 ( .A(n37157), .B(n37156), .Z(n37160) );
  XOR U46236 ( .A(n37159), .B(n37158), .Z(n37156) );
  XOR U46237 ( .A(y[2768]), .B(x[2768]), .Z(n37158) );
  XOR U46238 ( .A(y[2767]), .B(x[2767]), .Z(n37159) );
  XOR U46239 ( .A(y[2766]), .B(x[2766]), .Z(n37157) );
  XOR U46240 ( .A(n37151), .B(n37150), .Z(n37161) );
  XOR U46241 ( .A(n37153), .B(n37152), .Z(n37150) );
  XOR U46242 ( .A(y[2765]), .B(x[2765]), .Z(n37152) );
  XOR U46243 ( .A(y[2764]), .B(x[2764]), .Z(n37153) );
  XOR U46244 ( .A(y[2763]), .B(x[2763]), .Z(n37151) );
  XNOR U46245 ( .A(n37127), .B(n37128), .Z(n37145) );
  XNOR U46246 ( .A(n37142), .B(n37143), .Z(n37128) );
  XOR U46247 ( .A(n37139), .B(n37138), .Z(n37143) );
  XOR U46248 ( .A(y[2760]), .B(x[2760]), .Z(n37138) );
  XOR U46249 ( .A(n37141), .B(n37140), .Z(n37139) );
  XOR U46250 ( .A(y[2762]), .B(x[2762]), .Z(n37140) );
  XOR U46251 ( .A(y[2761]), .B(x[2761]), .Z(n37141) );
  XOR U46252 ( .A(n37133), .B(n37132), .Z(n37142) );
  XOR U46253 ( .A(n37135), .B(n37134), .Z(n37132) );
  XOR U46254 ( .A(y[2759]), .B(x[2759]), .Z(n37134) );
  XOR U46255 ( .A(y[2758]), .B(x[2758]), .Z(n37135) );
  XOR U46256 ( .A(y[2757]), .B(x[2757]), .Z(n37133) );
  XNOR U46257 ( .A(n37126), .B(n37125), .Z(n37127) );
  XNOR U46258 ( .A(n37122), .B(n37121), .Z(n37125) );
  XOR U46259 ( .A(n37124), .B(n37123), .Z(n37121) );
  XOR U46260 ( .A(y[2756]), .B(x[2756]), .Z(n37123) );
  XOR U46261 ( .A(y[2755]), .B(x[2755]), .Z(n37124) );
  XOR U46262 ( .A(y[2754]), .B(x[2754]), .Z(n37122) );
  XOR U46263 ( .A(n37116), .B(n37115), .Z(n37126) );
  XOR U46264 ( .A(n37118), .B(n37117), .Z(n37115) );
  XOR U46265 ( .A(y[2753]), .B(x[2753]), .Z(n37117) );
  XOR U46266 ( .A(y[2752]), .B(x[2752]), .Z(n37118) );
  XOR U46267 ( .A(y[2751]), .B(x[2751]), .Z(n37116) );
  NAND U46268 ( .A(n37179), .B(n37180), .Z(N62078) );
  NAND U46269 ( .A(n37181), .B(n37182), .Z(n37180) );
  NANDN U46270 ( .A(n37183), .B(n37184), .Z(n37182) );
  NANDN U46271 ( .A(n37184), .B(n37183), .Z(n37179) );
  XOR U46272 ( .A(n37183), .B(n37185), .Z(N62077) );
  XNOR U46273 ( .A(n37181), .B(n37184), .Z(n37185) );
  NAND U46274 ( .A(n37186), .B(n37187), .Z(n37184) );
  NAND U46275 ( .A(n37188), .B(n37189), .Z(n37187) );
  NANDN U46276 ( .A(n37190), .B(n37191), .Z(n37189) );
  NANDN U46277 ( .A(n37191), .B(n37190), .Z(n37186) );
  AND U46278 ( .A(n37192), .B(n37193), .Z(n37181) );
  NAND U46279 ( .A(n37194), .B(n37195), .Z(n37193) );
  NANDN U46280 ( .A(n37196), .B(n37197), .Z(n37195) );
  NANDN U46281 ( .A(n37197), .B(n37196), .Z(n37192) );
  IV U46282 ( .A(n37198), .Z(n37197) );
  AND U46283 ( .A(n37199), .B(n37200), .Z(n37183) );
  NAND U46284 ( .A(n37201), .B(n37202), .Z(n37200) );
  NANDN U46285 ( .A(n37203), .B(n37204), .Z(n37202) );
  NANDN U46286 ( .A(n37204), .B(n37203), .Z(n37199) );
  XOR U46287 ( .A(n37196), .B(n37205), .Z(N62076) );
  XNOR U46288 ( .A(n37194), .B(n37198), .Z(n37205) );
  XOR U46289 ( .A(n37191), .B(n37206), .Z(n37198) );
  XNOR U46290 ( .A(n37188), .B(n37190), .Z(n37206) );
  AND U46291 ( .A(n37207), .B(n37208), .Z(n37190) );
  NANDN U46292 ( .A(n37209), .B(n37210), .Z(n37208) );
  OR U46293 ( .A(n37211), .B(n37212), .Z(n37210) );
  IV U46294 ( .A(n37213), .Z(n37212) );
  NANDN U46295 ( .A(n37213), .B(n37211), .Z(n37207) );
  AND U46296 ( .A(n37214), .B(n37215), .Z(n37188) );
  NAND U46297 ( .A(n37216), .B(n37217), .Z(n37215) );
  NANDN U46298 ( .A(n37218), .B(n37219), .Z(n37217) );
  NANDN U46299 ( .A(n37219), .B(n37218), .Z(n37214) );
  IV U46300 ( .A(n37220), .Z(n37219) );
  NAND U46301 ( .A(n37221), .B(n37222), .Z(n37191) );
  NANDN U46302 ( .A(n37223), .B(n37224), .Z(n37222) );
  NANDN U46303 ( .A(n37225), .B(n37226), .Z(n37224) );
  NANDN U46304 ( .A(n37226), .B(n37225), .Z(n37221) );
  IV U46305 ( .A(n37227), .Z(n37225) );
  AND U46306 ( .A(n37228), .B(n37229), .Z(n37194) );
  NAND U46307 ( .A(n37230), .B(n37231), .Z(n37229) );
  NANDN U46308 ( .A(n37232), .B(n37233), .Z(n37231) );
  NANDN U46309 ( .A(n37233), .B(n37232), .Z(n37228) );
  XOR U46310 ( .A(n37204), .B(n37234), .Z(n37196) );
  XNOR U46311 ( .A(n37201), .B(n37203), .Z(n37234) );
  AND U46312 ( .A(n37235), .B(n37236), .Z(n37203) );
  NANDN U46313 ( .A(n37237), .B(n37238), .Z(n37236) );
  OR U46314 ( .A(n37239), .B(n37240), .Z(n37238) );
  IV U46315 ( .A(n37241), .Z(n37240) );
  NANDN U46316 ( .A(n37241), .B(n37239), .Z(n37235) );
  AND U46317 ( .A(n37242), .B(n37243), .Z(n37201) );
  NAND U46318 ( .A(n37244), .B(n37245), .Z(n37243) );
  NANDN U46319 ( .A(n37246), .B(n37247), .Z(n37245) );
  NANDN U46320 ( .A(n37247), .B(n37246), .Z(n37242) );
  IV U46321 ( .A(n37248), .Z(n37247) );
  NAND U46322 ( .A(n37249), .B(n37250), .Z(n37204) );
  NANDN U46323 ( .A(n37251), .B(n37252), .Z(n37250) );
  NANDN U46324 ( .A(n37253), .B(n37254), .Z(n37252) );
  NANDN U46325 ( .A(n37254), .B(n37253), .Z(n37249) );
  IV U46326 ( .A(n37255), .Z(n37253) );
  XOR U46327 ( .A(n37230), .B(n37256), .Z(N62075) );
  XNOR U46328 ( .A(n37233), .B(n37232), .Z(n37256) );
  XNOR U46329 ( .A(n37244), .B(n37257), .Z(n37232) );
  XNOR U46330 ( .A(n37248), .B(n37246), .Z(n37257) );
  XOR U46331 ( .A(n37254), .B(n37258), .Z(n37246) );
  XNOR U46332 ( .A(n37251), .B(n37255), .Z(n37258) );
  AND U46333 ( .A(n37259), .B(n37260), .Z(n37255) );
  NAND U46334 ( .A(n37261), .B(n37262), .Z(n37260) );
  NAND U46335 ( .A(n37263), .B(n37264), .Z(n37259) );
  AND U46336 ( .A(n37265), .B(n37266), .Z(n37251) );
  NAND U46337 ( .A(n37267), .B(n37268), .Z(n37266) );
  NAND U46338 ( .A(n37269), .B(n37270), .Z(n37265) );
  NANDN U46339 ( .A(n37271), .B(n37272), .Z(n37254) );
  ANDN U46340 ( .B(n37273), .A(n37274), .Z(n37248) );
  XNOR U46341 ( .A(n37239), .B(n37275), .Z(n37244) );
  XNOR U46342 ( .A(n37237), .B(n37241), .Z(n37275) );
  AND U46343 ( .A(n37276), .B(n37277), .Z(n37241) );
  NAND U46344 ( .A(n37278), .B(n37279), .Z(n37277) );
  NAND U46345 ( .A(n37280), .B(n37281), .Z(n37276) );
  AND U46346 ( .A(n37282), .B(n37283), .Z(n37237) );
  NAND U46347 ( .A(n37284), .B(n37285), .Z(n37283) );
  NAND U46348 ( .A(n37286), .B(n37287), .Z(n37282) );
  AND U46349 ( .A(n37288), .B(n37289), .Z(n37239) );
  NAND U46350 ( .A(n37290), .B(n37291), .Z(n37233) );
  XNOR U46351 ( .A(n37216), .B(n37292), .Z(n37230) );
  XNOR U46352 ( .A(n37220), .B(n37218), .Z(n37292) );
  XOR U46353 ( .A(n37226), .B(n37293), .Z(n37218) );
  XNOR U46354 ( .A(n37223), .B(n37227), .Z(n37293) );
  AND U46355 ( .A(n37294), .B(n37295), .Z(n37227) );
  NAND U46356 ( .A(n37296), .B(n37297), .Z(n37295) );
  NAND U46357 ( .A(n37298), .B(n37299), .Z(n37294) );
  AND U46358 ( .A(n37300), .B(n37301), .Z(n37223) );
  NAND U46359 ( .A(n37302), .B(n37303), .Z(n37301) );
  NAND U46360 ( .A(n37304), .B(n37305), .Z(n37300) );
  NANDN U46361 ( .A(n37306), .B(n37307), .Z(n37226) );
  ANDN U46362 ( .B(n37308), .A(n37309), .Z(n37220) );
  XNOR U46363 ( .A(n37211), .B(n37310), .Z(n37216) );
  XNOR U46364 ( .A(n37209), .B(n37213), .Z(n37310) );
  AND U46365 ( .A(n37311), .B(n37312), .Z(n37213) );
  NAND U46366 ( .A(n37313), .B(n37314), .Z(n37312) );
  NAND U46367 ( .A(n37315), .B(n37316), .Z(n37311) );
  AND U46368 ( .A(n37317), .B(n37318), .Z(n37209) );
  NAND U46369 ( .A(n37319), .B(n37320), .Z(n37318) );
  NAND U46370 ( .A(n37321), .B(n37322), .Z(n37317) );
  AND U46371 ( .A(n37323), .B(n37324), .Z(n37211) );
  XOR U46372 ( .A(n37291), .B(n37290), .Z(N62074) );
  XNOR U46373 ( .A(n37308), .B(n37309), .Z(n37290) );
  XNOR U46374 ( .A(n37323), .B(n37324), .Z(n37309) );
  XOR U46375 ( .A(n37320), .B(n37319), .Z(n37324) );
  XOR U46376 ( .A(y[2748]), .B(x[2748]), .Z(n37319) );
  XOR U46377 ( .A(n37322), .B(n37321), .Z(n37320) );
  XOR U46378 ( .A(y[2750]), .B(x[2750]), .Z(n37321) );
  XOR U46379 ( .A(y[2749]), .B(x[2749]), .Z(n37322) );
  XOR U46380 ( .A(n37314), .B(n37313), .Z(n37323) );
  XOR U46381 ( .A(n37316), .B(n37315), .Z(n37313) );
  XOR U46382 ( .A(y[2747]), .B(x[2747]), .Z(n37315) );
  XOR U46383 ( .A(y[2746]), .B(x[2746]), .Z(n37316) );
  XOR U46384 ( .A(y[2745]), .B(x[2745]), .Z(n37314) );
  XNOR U46385 ( .A(n37307), .B(n37306), .Z(n37308) );
  XNOR U46386 ( .A(n37303), .B(n37302), .Z(n37306) );
  XOR U46387 ( .A(n37305), .B(n37304), .Z(n37302) );
  XOR U46388 ( .A(y[2744]), .B(x[2744]), .Z(n37304) );
  XOR U46389 ( .A(y[2743]), .B(x[2743]), .Z(n37305) );
  XOR U46390 ( .A(y[2742]), .B(x[2742]), .Z(n37303) );
  XOR U46391 ( .A(n37297), .B(n37296), .Z(n37307) );
  XOR U46392 ( .A(n37299), .B(n37298), .Z(n37296) );
  XOR U46393 ( .A(y[2741]), .B(x[2741]), .Z(n37298) );
  XOR U46394 ( .A(y[2740]), .B(x[2740]), .Z(n37299) );
  XOR U46395 ( .A(y[2739]), .B(x[2739]), .Z(n37297) );
  XNOR U46396 ( .A(n37273), .B(n37274), .Z(n37291) );
  XNOR U46397 ( .A(n37288), .B(n37289), .Z(n37274) );
  XOR U46398 ( .A(n37285), .B(n37284), .Z(n37289) );
  XOR U46399 ( .A(y[2736]), .B(x[2736]), .Z(n37284) );
  XOR U46400 ( .A(n37287), .B(n37286), .Z(n37285) );
  XOR U46401 ( .A(y[2738]), .B(x[2738]), .Z(n37286) );
  XOR U46402 ( .A(y[2737]), .B(x[2737]), .Z(n37287) );
  XOR U46403 ( .A(n37279), .B(n37278), .Z(n37288) );
  XOR U46404 ( .A(n37281), .B(n37280), .Z(n37278) );
  XOR U46405 ( .A(y[2735]), .B(x[2735]), .Z(n37280) );
  XOR U46406 ( .A(y[2734]), .B(x[2734]), .Z(n37281) );
  XOR U46407 ( .A(y[2733]), .B(x[2733]), .Z(n37279) );
  XNOR U46408 ( .A(n37272), .B(n37271), .Z(n37273) );
  XNOR U46409 ( .A(n37268), .B(n37267), .Z(n37271) );
  XOR U46410 ( .A(n37270), .B(n37269), .Z(n37267) );
  XOR U46411 ( .A(y[2732]), .B(x[2732]), .Z(n37269) );
  XOR U46412 ( .A(y[2731]), .B(x[2731]), .Z(n37270) );
  XOR U46413 ( .A(y[2730]), .B(x[2730]), .Z(n37268) );
  XOR U46414 ( .A(n37262), .B(n37261), .Z(n37272) );
  XOR U46415 ( .A(n37264), .B(n37263), .Z(n37261) );
  XOR U46416 ( .A(y[2729]), .B(x[2729]), .Z(n37263) );
  XOR U46417 ( .A(y[2728]), .B(x[2728]), .Z(n37264) );
  XOR U46418 ( .A(y[2727]), .B(x[2727]), .Z(n37262) );
  NAND U46419 ( .A(n37325), .B(n37326), .Z(N62065) );
  NAND U46420 ( .A(n37327), .B(n37328), .Z(n37326) );
  NANDN U46421 ( .A(n37329), .B(n37330), .Z(n37328) );
  NANDN U46422 ( .A(n37330), .B(n37329), .Z(n37325) );
  XOR U46423 ( .A(n37329), .B(n37331), .Z(N62064) );
  XNOR U46424 ( .A(n37327), .B(n37330), .Z(n37331) );
  NAND U46425 ( .A(n37332), .B(n37333), .Z(n37330) );
  NAND U46426 ( .A(n37334), .B(n37335), .Z(n37333) );
  NANDN U46427 ( .A(n37336), .B(n37337), .Z(n37335) );
  NANDN U46428 ( .A(n37337), .B(n37336), .Z(n37332) );
  AND U46429 ( .A(n37338), .B(n37339), .Z(n37327) );
  NAND U46430 ( .A(n37340), .B(n37341), .Z(n37339) );
  NANDN U46431 ( .A(n37342), .B(n37343), .Z(n37341) );
  NANDN U46432 ( .A(n37343), .B(n37342), .Z(n37338) );
  IV U46433 ( .A(n37344), .Z(n37343) );
  AND U46434 ( .A(n37345), .B(n37346), .Z(n37329) );
  NAND U46435 ( .A(n37347), .B(n37348), .Z(n37346) );
  NANDN U46436 ( .A(n37349), .B(n37350), .Z(n37348) );
  NANDN U46437 ( .A(n37350), .B(n37349), .Z(n37345) );
  XOR U46438 ( .A(n37342), .B(n37351), .Z(N62063) );
  XNOR U46439 ( .A(n37340), .B(n37344), .Z(n37351) );
  XOR U46440 ( .A(n37337), .B(n37352), .Z(n37344) );
  XNOR U46441 ( .A(n37334), .B(n37336), .Z(n37352) );
  AND U46442 ( .A(n37353), .B(n37354), .Z(n37336) );
  NANDN U46443 ( .A(n37355), .B(n37356), .Z(n37354) );
  OR U46444 ( .A(n37357), .B(n37358), .Z(n37356) );
  IV U46445 ( .A(n37359), .Z(n37358) );
  NANDN U46446 ( .A(n37359), .B(n37357), .Z(n37353) );
  AND U46447 ( .A(n37360), .B(n37361), .Z(n37334) );
  NAND U46448 ( .A(n37362), .B(n37363), .Z(n37361) );
  NANDN U46449 ( .A(n37364), .B(n37365), .Z(n37363) );
  NANDN U46450 ( .A(n37365), .B(n37364), .Z(n37360) );
  IV U46451 ( .A(n37366), .Z(n37365) );
  NAND U46452 ( .A(n37367), .B(n37368), .Z(n37337) );
  NANDN U46453 ( .A(n37369), .B(n37370), .Z(n37368) );
  NANDN U46454 ( .A(n37371), .B(n37372), .Z(n37370) );
  NANDN U46455 ( .A(n37372), .B(n37371), .Z(n37367) );
  IV U46456 ( .A(n37373), .Z(n37371) );
  AND U46457 ( .A(n37374), .B(n37375), .Z(n37340) );
  NAND U46458 ( .A(n37376), .B(n37377), .Z(n37375) );
  NANDN U46459 ( .A(n37378), .B(n37379), .Z(n37377) );
  NANDN U46460 ( .A(n37379), .B(n37378), .Z(n37374) );
  XOR U46461 ( .A(n37350), .B(n37380), .Z(n37342) );
  XNOR U46462 ( .A(n37347), .B(n37349), .Z(n37380) );
  AND U46463 ( .A(n37381), .B(n37382), .Z(n37349) );
  NANDN U46464 ( .A(n37383), .B(n37384), .Z(n37382) );
  OR U46465 ( .A(n37385), .B(n37386), .Z(n37384) );
  IV U46466 ( .A(n37387), .Z(n37386) );
  NANDN U46467 ( .A(n37387), .B(n37385), .Z(n37381) );
  AND U46468 ( .A(n37388), .B(n37389), .Z(n37347) );
  NAND U46469 ( .A(n37390), .B(n37391), .Z(n37389) );
  NANDN U46470 ( .A(n37392), .B(n37393), .Z(n37391) );
  NANDN U46471 ( .A(n37393), .B(n37392), .Z(n37388) );
  IV U46472 ( .A(n37394), .Z(n37393) );
  NAND U46473 ( .A(n37395), .B(n37396), .Z(n37350) );
  NANDN U46474 ( .A(n37397), .B(n37398), .Z(n37396) );
  NANDN U46475 ( .A(n37399), .B(n37400), .Z(n37398) );
  NANDN U46476 ( .A(n37400), .B(n37399), .Z(n37395) );
  IV U46477 ( .A(n37401), .Z(n37399) );
  XOR U46478 ( .A(n37376), .B(n37402), .Z(N62062) );
  XNOR U46479 ( .A(n37379), .B(n37378), .Z(n37402) );
  XNOR U46480 ( .A(n37390), .B(n37403), .Z(n37378) );
  XNOR U46481 ( .A(n37394), .B(n37392), .Z(n37403) );
  XOR U46482 ( .A(n37400), .B(n37404), .Z(n37392) );
  XNOR U46483 ( .A(n37397), .B(n37401), .Z(n37404) );
  AND U46484 ( .A(n37405), .B(n37406), .Z(n37401) );
  NAND U46485 ( .A(n37407), .B(n37408), .Z(n37406) );
  NAND U46486 ( .A(n37409), .B(n37410), .Z(n37405) );
  AND U46487 ( .A(n37411), .B(n37412), .Z(n37397) );
  NAND U46488 ( .A(n37413), .B(n37414), .Z(n37412) );
  NAND U46489 ( .A(n37415), .B(n37416), .Z(n37411) );
  NANDN U46490 ( .A(n37417), .B(n37418), .Z(n37400) );
  ANDN U46491 ( .B(n37419), .A(n37420), .Z(n37394) );
  XNOR U46492 ( .A(n37385), .B(n37421), .Z(n37390) );
  XNOR U46493 ( .A(n37383), .B(n37387), .Z(n37421) );
  AND U46494 ( .A(n37422), .B(n37423), .Z(n37387) );
  NAND U46495 ( .A(n37424), .B(n37425), .Z(n37423) );
  NAND U46496 ( .A(n37426), .B(n37427), .Z(n37422) );
  AND U46497 ( .A(n37428), .B(n37429), .Z(n37383) );
  NAND U46498 ( .A(n37430), .B(n37431), .Z(n37429) );
  NAND U46499 ( .A(n37432), .B(n37433), .Z(n37428) );
  AND U46500 ( .A(n37434), .B(n37435), .Z(n37385) );
  NAND U46501 ( .A(n37436), .B(n37437), .Z(n37379) );
  XNOR U46502 ( .A(n37362), .B(n37438), .Z(n37376) );
  XNOR U46503 ( .A(n37366), .B(n37364), .Z(n37438) );
  XOR U46504 ( .A(n37372), .B(n37439), .Z(n37364) );
  XNOR U46505 ( .A(n37369), .B(n37373), .Z(n37439) );
  AND U46506 ( .A(n37440), .B(n37441), .Z(n37373) );
  NAND U46507 ( .A(n37442), .B(n37443), .Z(n37441) );
  NAND U46508 ( .A(n37444), .B(n37445), .Z(n37440) );
  AND U46509 ( .A(n37446), .B(n37447), .Z(n37369) );
  NAND U46510 ( .A(n37448), .B(n37449), .Z(n37447) );
  NAND U46511 ( .A(n37450), .B(n37451), .Z(n37446) );
  NANDN U46512 ( .A(n37452), .B(n37453), .Z(n37372) );
  ANDN U46513 ( .B(n37454), .A(n37455), .Z(n37366) );
  XNOR U46514 ( .A(n37357), .B(n37456), .Z(n37362) );
  XNOR U46515 ( .A(n37355), .B(n37359), .Z(n37456) );
  AND U46516 ( .A(n37457), .B(n37458), .Z(n37359) );
  NAND U46517 ( .A(n37459), .B(n37460), .Z(n37458) );
  NAND U46518 ( .A(n37461), .B(n37462), .Z(n37457) );
  AND U46519 ( .A(n37463), .B(n37464), .Z(n37355) );
  NAND U46520 ( .A(n37465), .B(n37466), .Z(n37464) );
  NAND U46521 ( .A(n37467), .B(n37468), .Z(n37463) );
  AND U46522 ( .A(n37469), .B(n37470), .Z(n37357) );
  XOR U46523 ( .A(n37437), .B(n37436), .Z(N62061) );
  XNOR U46524 ( .A(n37454), .B(n37455), .Z(n37436) );
  XNOR U46525 ( .A(n37469), .B(n37470), .Z(n37455) );
  XOR U46526 ( .A(n37466), .B(n37465), .Z(n37470) );
  XOR U46527 ( .A(y[2724]), .B(x[2724]), .Z(n37465) );
  XOR U46528 ( .A(n37468), .B(n37467), .Z(n37466) );
  XOR U46529 ( .A(y[2726]), .B(x[2726]), .Z(n37467) );
  XOR U46530 ( .A(y[2725]), .B(x[2725]), .Z(n37468) );
  XOR U46531 ( .A(n37460), .B(n37459), .Z(n37469) );
  XOR U46532 ( .A(n37462), .B(n37461), .Z(n37459) );
  XOR U46533 ( .A(y[2723]), .B(x[2723]), .Z(n37461) );
  XOR U46534 ( .A(y[2722]), .B(x[2722]), .Z(n37462) );
  XOR U46535 ( .A(y[2721]), .B(x[2721]), .Z(n37460) );
  XNOR U46536 ( .A(n37453), .B(n37452), .Z(n37454) );
  XNOR U46537 ( .A(n37449), .B(n37448), .Z(n37452) );
  XOR U46538 ( .A(n37451), .B(n37450), .Z(n37448) );
  XOR U46539 ( .A(y[2720]), .B(x[2720]), .Z(n37450) );
  XOR U46540 ( .A(y[2719]), .B(x[2719]), .Z(n37451) );
  XOR U46541 ( .A(y[2718]), .B(x[2718]), .Z(n37449) );
  XOR U46542 ( .A(n37443), .B(n37442), .Z(n37453) );
  XOR U46543 ( .A(n37445), .B(n37444), .Z(n37442) );
  XOR U46544 ( .A(y[2717]), .B(x[2717]), .Z(n37444) );
  XOR U46545 ( .A(y[2716]), .B(x[2716]), .Z(n37445) );
  XOR U46546 ( .A(y[2715]), .B(x[2715]), .Z(n37443) );
  XNOR U46547 ( .A(n37419), .B(n37420), .Z(n37437) );
  XNOR U46548 ( .A(n37434), .B(n37435), .Z(n37420) );
  XOR U46549 ( .A(n37431), .B(n37430), .Z(n37435) );
  XOR U46550 ( .A(y[2712]), .B(x[2712]), .Z(n37430) );
  XOR U46551 ( .A(n37433), .B(n37432), .Z(n37431) );
  XOR U46552 ( .A(y[2714]), .B(x[2714]), .Z(n37432) );
  XOR U46553 ( .A(y[2713]), .B(x[2713]), .Z(n37433) );
  XOR U46554 ( .A(n37425), .B(n37424), .Z(n37434) );
  XOR U46555 ( .A(n37427), .B(n37426), .Z(n37424) );
  XOR U46556 ( .A(y[2711]), .B(x[2711]), .Z(n37426) );
  XOR U46557 ( .A(y[2710]), .B(x[2710]), .Z(n37427) );
  XOR U46558 ( .A(y[2709]), .B(x[2709]), .Z(n37425) );
  XNOR U46559 ( .A(n37418), .B(n37417), .Z(n37419) );
  XNOR U46560 ( .A(n37414), .B(n37413), .Z(n37417) );
  XOR U46561 ( .A(n37416), .B(n37415), .Z(n37413) );
  XOR U46562 ( .A(y[2708]), .B(x[2708]), .Z(n37415) );
  XOR U46563 ( .A(y[2707]), .B(x[2707]), .Z(n37416) );
  XOR U46564 ( .A(y[2706]), .B(x[2706]), .Z(n37414) );
  XOR U46565 ( .A(n37408), .B(n37407), .Z(n37418) );
  XOR U46566 ( .A(n37410), .B(n37409), .Z(n37407) );
  XOR U46567 ( .A(y[2705]), .B(x[2705]), .Z(n37409) );
  XOR U46568 ( .A(y[2704]), .B(x[2704]), .Z(n37410) );
  XOR U46569 ( .A(y[2703]), .B(x[2703]), .Z(n37408) );
  NAND U46570 ( .A(n37471), .B(n37472), .Z(N62052) );
  NAND U46571 ( .A(n37473), .B(n37474), .Z(n37472) );
  NANDN U46572 ( .A(n37475), .B(n37476), .Z(n37474) );
  NANDN U46573 ( .A(n37476), .B(n37475), .Z(n37471) );
  XOR U46574 ( .A(n37475), .B(n37477), .Z(N62051) );
  XNOR U46575 ( .A(n37473), .B(n37476), .Z(n37477) );
  NAND U46576 ( .A(n37478), .B(n37479), .Z(n37476) );
  NAND U46577 ( .A(n37480), .B(n37481), .Z(n37479) );
  NANDN U46578 ( .A(n37482), .B(n37483), .Z(n37481) );
  NANDN U46579 ( .A(n37483), .B(n37482), .Z(n37478) );
  AND U46580 ( .A(n37484), .B(n37485), .Z(n37473) );
  NAND U46581 ( .A(n37486), .B(n37487), .Z(n37485) );
  NANDN U46582 ( .A(n37488), .B(n37489), .Z(n37487) );
  NANDN U46583 ( .A(n37489), .B(n37488), .Z(n37484) );
  IV U46584 ( .A(n37490), .Z(n37489) );
  AND U46585 ( .A(n37491), .B(n37492), .Z(n37475) );
  NAND U46586 ( .A(n37493), .B(n37494), .Z(n37492) );
  NANDN U46587 ( .A(n37495), .B(n37496), .Z(n37494) );
  NANDN U46588 ( .A(n37496), .B(n37495), .Z(n37491) );
  XOR U46589 ( .A(n37488), .B(n37497), .Z(N62050) );
  XNOR U46590 ( .A(n37486), .B(n37490), .Z(n37497) );
  XOR U46591 ( .A(n37483), .B(n37498), .Z(n37490) );
  XNOR U46592 ( .A(n37480), .B(n37482), .Z(n37498) );
  AND U46593 ( .A(n37499), .B(n37500), .Z(n37482) );
  NANDN U46594 ( .A(n37501), .B(n37502), .Z(n37500) );
  OR U46595 ( .A(n37503), .B(n37504), .Z(n37502) );
  IV U46596 ( .A(n37505), .Z(n37504) );
  NANDN U46597 ( .A(n37505), .B(n37503), .Z(n37499) );
  AND U46598 ( .A(n37506), .B(n37507), .Z(n37480) );
  NAND U46599 ( .A(n37508), .B(n37509), .Z(n37507) );
  NANDN U46600 ( .A(n37510), .B(n37511), .Z(n37509) );
  NANDN U46601 ( .A(n37511), .B(n37510), .Z(n37506) );
  IV U46602 ( .A(n37512), .Z(n37511) );
  NAND U46603 ( .A(n37513), .B(n37514), .Z(n37483) );
  NANDN U46604 ( .A(n37515), .B(n37516), .Z(n37514) );
  NANDN U46605 ( .A(n37517), .B(n37518), .Z(n37516) );
  NANDN U46606 ( .A(n37518), .B(n37517), .Z(n37513) );
  IV U46607 ( .A(n37519), .Z(n37517) );
  AND U46608 ( .A(n37520), .B(n37521), .Z(n37486) );
  NAND U46609 ( .A(n37522), .B(n37523), .Z(n37521) );
  NANDN U46610 ( .A(n37524), .B(n37525), .Z(n37523) );
  NANDN U46611 ( .A(n37525), .B(n37524), .Z(n37520) );
  XOR U46612 ( .A(n37496), .B(n37526), .Z(n37488) );
  XNOR U46613 ( .A(n37493), .B(n37495), .Z(n37526) );
  AND U46614 ( .A(n37527), .B(n37528), .Z(n37495) );
  NANDN U46615 ( .A(n37529), .B(n37530), .Z(n37528) );
  OR U46616 ( .A(n37531), .B(n37532), .Z(n37530) );
  IV U46617 ( .A(n37533), .Z(n37532) );
  NANDN U46618 ( .A(n37533), .B(n37531), .Z(n37527) );
  AND U46619 ( .A(n37534), .B(n37535), .Z(n37493) );
  NAND U46620 ( .A(n37536), .B(n37537), .Z(n37535) );
  NANDN U46621 ( .A(n37538), .B(n37539), .Z(n37537) );
  NANDN U46622 ( .A(n37539), .B(n37538), .Z(n37534) );
  IV U46623 ( .A(n37540), .Z(n37539) );
  NAND U46624 ( .A(n37541), .B(n37542), .Z(n37496) );
  NANDN U46625 ( .A(n37543), .B(n37544), .Z(n37542) );
  NANDN U46626 ( .A(n37545), .B(n37546), .Z(n37544) );
  NANDN U46627 ( .A(n37546), .B(n37545), .Z(n37541) );
  IV U46628 ( .A(n37547), .Z(n37545) );
  XOR U46629 ( .A(n37522), .B(n37548), .Z(N62049) );
  XNOR U46630 ( .A(n37525), .B(n37524), .Z(n37548) );
  XNOR U46631 ( .A(n37536), .B(n37549), .Z(n37524) );
  XNOR U46632 ( .A(n37540), .B(n37538), .Z(n37549) );
  XOR U46633 ( .A(n37546), .B(n37550), .Z(n37538) );
  XNOR U46634 ( .A(n37543), .B(n37547), .Z(n37550) );
  AND U46635 ( .A(n37551), .B(n37552), .Z(n37547) );
  NAND U46636 ( .A(n37553), .B(n37554), .Z(n37552) );
  NAND U46637 ( .A(n37555), .B(n37556), .Z(n37551) );
  AND U46638 ( .A(n37557), .B(n37558), .Z(n37543) );
  NAND U46639 ( .A(n37559), .B(n37560), .Z(n37558) );
  NAND U46640 ( .A(n37561), .B(n37562), .Z(n37557) );
  NANDN U46641 ( .A(n37563), .B(n37564), .Z(n37546) );
  ANDN U46642 ( .B(n37565), .A(n37566), .Z(n37540) );
  XNOR U46643 ( .A(n37531), .B(n37567), .Z(n37536) );
  XNOR U46644 ( .A(n37529), .B(n37533), .Z(n37567) );
  AND U46645 ( .A(n37568), .B(n37569), .Z(n37533) );
  NAND U46646 ( .A(n37570), .B(n37571), .Z(n37569) );
  NAND U46647 ( .A(n37572), .B(n37573), .Z(n37568) );
  AND U46648 ( .A(n37574), .B(n37575), .Z(n37529) );
  NAND U46649 ( .A(n37576), .B(n37577), .Z(n37575) );
  NAND U46650 ( .A(n37578), .B(n37579), .Z(n37574) );
  AND U46651 ( .A(n37580), .B(n37581), .Z(n37531) );
  NAND U46652 ( .A(n37582), .B(n37583), .Z(n37525) );
  XNOR U46653 ( .A(n37508), .B(n37584), .Z(n37522) );
  XNOR U46654 ( .A(n37512), .B(n37510), .Z(n37584) );
  XOR U46655 ( .A(n37518), .B(n37585), .Z(n37510) );
  XNOR U46656 ( .A(n37515), .B(n37519), .Z(n37585) );
  AND U46657 ( .A(n37586), .B(n37587), .Z(n37519) );
  NAND U46658 ( .A(n37588), .B(n37589), .Z(n37587) );
  NAND U46659 ( .A(n37590), .B(n37591), .Z(n37586) );
  AND U46660 ( .A(n37592), .B(n37593), .Z(n37515) );
  NAND U46661 ( .A(n37594), .B(n37595), .Z(n37593) );
  NAND U46662 ( .A(n37596), .B(n37597), .Z(n37592) );
  NANDN U46663 ( .A(n37598), .B(n37599), .Z(n37518) );
  ANDN U46664 ( .B(n37600), .A(n37601), .Z(n37512) );
  XNOR U46665 ( .A(n37503), .B(n37602), .Z(n37508) );
  XNOR U46666 ( .A(n37501), .B(n37505), .Z(n37602) );
  AND U46667 ( .A(n37603), .B(n37604), .Z(n37505) );
  NAND U46668 ( .A(n37605), .B(n37606), .Z(n37604) );
  NAND U46669 ( .A(n37607), .B(n37608), .Z(n37603) );
  AND U46670 ( .A(n37609), .B(n37610), .Z(n37501) );
  NAND U46671 ( .A(n37611), .B(n37612), .Z(n37610) );
  NAND U46672 ( .A(n37613), .B(n37614), .Z(n37609) );
  AND U46673 ( .A(n37615), .B(n37616), .Z(n37503) );
  XOR U46674 ( .A(n37583), .B(n37582), .Z(N62048) );
  XNOR U46675 ( .A(n37600), .B(n37601), .Z(n37582) );
  XNOR U46676 ( .A(n37615), .B(n37616), .Z(n37601) );
  XOR U46677 ( .A(n37612), .B(n37611), .Z(n37616) );
  XOR U46678 ( .A(y[2700]), .B(x[2700]), .Z(n37611) );
  XOR U46679 ( .A(n37614), .B(n37613), .Z(n37612) );
  XOR U46680 ( .A(y[2702]), .B(x[2702]), .Z(n37613) );
  XOR U46681 ( .A(y[2701]), .B(x[2701]), .Z(n37614) );
  XOR U46682 ( .A(n37606), .B(n37605), .Z(n37615) );
  XOR U46683 ( .A(n37608), .B(n37607), .Z(n37605) );
  XOR U46684 ( .A(y[2699]), .B(x[2699]), .Z(n37607) );
  XOR U46685 ( .A(y[2698]), .B(x[2698]), .Z(n37608) );
  XOR U46686 ( .A(y[2697]), .B(x[2697]), .Z(n37606) );
  XNOR U46687 ( .A(n37599), .B(n37598), .Z(n37600) );
  XNOR U46688 ( .A(n37595), .B(n37594), .Z(n37598) );
  XOR U46689 ( .A(n37597), .B(n37596), .Z(n37594) );
  XOR U46690 ( .A(y[2696]), .B(x[2696]), .Z(n37596) );
  XOR U46691 ( .A(y[2695]), .B(x[2695]), .Z(n37597) );
  XOR U46692 ( .A(y[2694]), .B(x[2694]), .Z(n37595) );
  XOR U46693 ( .A(n37589), .B(n37588), .Z(n37599) );
  XOR U46694 ( .A(n37591), .B(n37590), .Z(n37588) );
  XOR U46695 ( .A(y[2693]), .B(x[2693]), .Z(n37590) );
  XOR U46696 ( .A(y[2692]), .B(x[2692]), .Z(n37591) );
  XOR U46697 ( .A(y[2691]), .B(x[2691]), .Z(n37589) );
  XNOR U46698 ( .A(n37565), .B(n37566), .Z(n37583) );
  XNOR U46699 ( .A(n37580), .B(n37581), .Z(n37566) );
  XOR U46700 ( .A(n37577), .B(n37576), .Z(n37581) );
  XOR U46701 ( .A(y[2688]), .B(x[2688]), .Z(n37576) );
  XOR U46702 ( .A(n37579), .B(n37578), .Z(n37577) );
  XOR U46703 ( .A(y[2690]), .B(x[2690]), .Z(n37578) );
  XOR U46704 ( .A(y[2689]), .B(x[2689]), .Z(n37579) );
  XOR U46705 ( .A(n37571), .B(n37570), .Z(n37580) );
  XOR U46706 ( .A(n37573), .B(n37572), .Z(n37570) );
  XOR U46707 ( .A(y[2687]), .B(x[2687]), .Z(n37572) );
  XOR U46708 ( .A(y[2686]), .B(x[2686]), .Z(n37573) );
  XOR U46709 ( .A(y[2685]), .B(x[2685]), .Z(n37571) );
  XNOR U46710 ( .A(n37564), .B(n37563), .Z(n37565) );
  XNOR U46711 ( .A(n37560), .B(n37559), .Z(n37563) );
  XOR U46712 ( .A(n37562), .B(n37561), .Z(n37559) );
  XOR U46713 ( .A(y[2684]), .B(x[2684]), .Z(n37561) );
  XOR U46714 ( .A(y[2683]), .B(x[2683]), .Z(n37562) );
  XOR U46715 ( .A(y[2682]), .B(x[2682]), .Z(n37560) );
  XOR U46716 ( .A(n37554), .B(n37553), .Z(n37564) );
  XOR U46717 ( .A(n37556), .B(n37555), .Z(n37553) );
  XOR U46718 ( .A(y[2681]), .B(x[2681]), .Z(n37555) );
  XOR U46719 ( .A(y[2680]), .B(x[2680]), .Z(n37556) );
  XOR U46720 ( .A(y[2679]), .B(x[2679]), .Z(n37554) );
  NAND U46721 ( .A(n37617), .B(n37618), .Z(N62039) );
  NAND U46722 ( .A(n37619), .B(n37620), .Z(n37618) );
  NANDN U46723 ( .A(n37621), .B(n37622), .Z(n37620) );
  NANDN U46724 ( .A(n37622), .B(n37621), .Z(n37617) );
  XOR U46725 ( .A(n37621), .B(n37623), .Z(N62038) );
  XNOR U46726 ( .A(n37619), .B(n37622), .Z(n37623) );
  NAND U46727 ( .A(n37624), .B(n37625), .Z(n37622) );
  NAND U46728 ( .A(n37626), .B(n37627), .Z(n37625) );
  NANDN U46729 ( .A(n37628), .B(n37629), .Z(n37627) );
  NANDN U46730 ( .A(n37629), .B(n37628), .Z(n37624) );
  AND U46731 ( .A(n37630), .B(n37631), .Z(n37619) );
  NAND U46732 ( .A(n37632), .B(n37633), .Z(n37631) );
  NANDN U46733 ( .A(n37634), .B(n37635), .Z(n37633) );
  NANDN U46734 ( .A(n37635), .B(n37634), .Z(n37630) );
  IV U46735 ( .A(n37636), .Z(n37635) );
  AND U46736 ( .A(n37637), .B(n37638), .Z(n37621) );
  NAND U46737 ( .A(n37639), .B(n37640), .Z(n37638) );
  NANDN U46738 ( .A(n37641), .B(n37642), .Z(n37640) );
  NANDN U46739 ( .A(n37642), .B(n37641), .Z(n37637) );
  XOR U46740 ( .A(n37634), .B(n37643), .Z(N62037) );
  XNOR U46741 ( .A(n37632), .B(n37636), .Z(n37643) );
  XOR U46742 ( .A(n37629), .B(n37644), .Z(n37636) );
  XNOR U46743 ( .A(n37626), .B(n37628), .Z(n37644) );
  AND U46744 ( .A(n37645), .B(n37646), .Z(n37628) );
  NANDN U46745 ( .A(n37647), .B(n37648), .Z(n37646) );
  OR U46746 ( .A(n37649), .B(n37650), .Z(n37648) );
  IV U46747 ( .A(n37651), .Z(n37650) );
  NANDN U46748 ( .A(n37651), .B(n37649), .Z(n37645) );
  AND U46749 ( .A(n37652), .B(n37653), .Z(n37626) );
  NAND U46750 ( .A(n37654), .B(n37655), .Z(n37653) );
  NANDN U46751 ( .A(n37656), .B(n37657), .Z(n37655) );
  NANDN U46752 ( .A(n37657), .B(n37656), .Z(n37652) );
  IV U46753 ( .A(n37658), .Z(n37657) );
  NAND U46754 ( .A(n37659), .B(n37660), .Z(n37629) );
  NANDN U46755 ( .A(n37661), .B(n37662), .Z(n37660) );
  NANDN U46756 ( .A(n37663), .B(n37664), .Z(n37662) );
  NANDN U46757 ( .A(n37664), .B(n37663), .Z(n37659) );
  IV U46758 ( .A(n37665), .Z(n37663) );
  AND U46759 ( .A(n37666), .B(n37667), .Z(n37632) );
  NAND U46760 ( .A(n37668), .B(n37669), .Z(n37667) );
  NANDN U46761 ( .A(n37670), .B(n37671), .Z(n37669) );
  NANDN U46762 ( .A(n37671), .B(n37670), .Z(n37666) );
  XOR U46763 ( .A(n37642), .B(n37672), .Z(n37634) );
  XNOR U46764 ( .A(n37639), .B(n37641), .Z(n37672) );
  AND U46765 ( .A(n37673), .B(n37674), .Z(n37641) );
  NANDN U46766 ( .A(n37675), .B(n37676), .Z(n37674) );
  OR U46767 ( .A(n37677), .B(n37678), .Z(n37676) );
  IV U46768 ( .A(n37679), .Z(n37678) );
  NANDN U46769 ( .A(n37679), .B(n37677), .Z(n37673) );
  AND U46770 ( .A(n37680), .B(n37681), .Z(n37639) );
  NAND U46771 ( .A(n37682), .B(n37683), .Z(n37681) );
  NANDN U46772 ( .A(n37684), .B(n37685), .Z(n37683) );
  NANDN U46773 ( .A(n37685), .B(n37684), .Z(n37680) );
  IV U46774 ( .A(n37686), .Z(n37685) );
  NAND U46775 ( .A(n37687), .B(n37688), .Z(n37642) );
  NANDN U46776 ( .A(n37689), .B(n37690), .Z(n37688) );
  NANDN U46777 ( .A(n37691), .B(n37692), .Z(n37690) );
  NANDN U46778 ( .A(n37692), .B(n37691), .Z(n37687) );
  IV U46779 ( .A(n37693), .Z(n37691) );
  XOR U46780 ( .A(n37668), .B(n37694), .Z(N62036) );
  XNOR U46781 ( .A(n37671), .B(n37670), .Z(n37694) );
  XNOR U46782 ( .A(n37682), .B(n37695), .Z(n37670) );
  XNOR U46783 ( .A(n37686), .B(n37684), .Z(n37695) );
  XOR U46784 ( .A(n37692), .B(n37696), .Z(n37684) );
  XNOR U46785 ( .A(n37689), .B(n37693), .Z(n37696) );
  AND U46786 ( .A(n37697), .B(n37698), .Z(n37693) );
  NAND U46787 ( .A(n37699), .B(n37700), .Z(n37698) );
  NAND U46788 ( .A(n37701), .B(n37702), .Z(n37697) );
  AND U46789 ( .A(n37703), .B(n37704), .Z(n37689) );
  NAND U46790 ( .A(n37705), .B(n37706), .Z(n37704) );
  NAND U46791 ( .A(n37707), .B(n37708), .Z(n37703) );
  NANDN U46792 ( .A(n37709), .B(n37710), .Z(n37692) );
  ANDN U46793 ( .B(n37711), .A(n37712), .Z(n37686) );
  XNOR U46794 ( .A(n37677), .B(n37713), .Z(n37682) );
  XNOR U46795 ( .A(n37675), .B(n37679), .Z(n37713) );
  AND U46796 ( .A(n37714), .B(n37715), .Z(n37679) );
  NAND U46797 ( .A(n37716), .B(n37717), .Z(n37715) );
  NAND U46798 ( .A(n37718), .B(n37719), .Z(n37714) );
  AND U46799 ( .A(n37720), .B(n37721), .Z(n37675) );
  NAND U46800 ( .A(n37722), .B(n37723), .Z(n37721) );
  NAND U46801 ( .A(n37724), .B(n37725), .Z(n37720) );
  AND U46802 ( .A(n37726), .B(n37727), .Z(n37677) );
  NAND U46803 ( .A(n37728), .B(n37729), .Z(n37671) );
  XNOR U46804 ( .A(n37654), .B(n37730), .Z(n37668) );
  XNOR U46805 ( .A(n37658), .B(n37656), .Z(n37730) );
  XOR U46806 ( .A(n37664), .B(n37731), .Z(n37656) );
  XNOR U46807 ( .A(n37661), .B(n37665), .Z(n37731) );
  AND U46808 ( .A(n37732), .B(n37733), .Z(n37665) );
  NAND U46809 ( .A(n37734), .B(n37735), .Z(n37733) );
  NAND U46810 ( .A(n37736), .B(n37737), .Z(n37732) );
  AND U46811 ( .A(n37738), .B(n37739), .Z(n37661) );
  NAND U46812 ( .A(n37740), .B(n37741), .Z(n37739) );
  NAND U46813 ( .A(n37742), .B(n37743), .Z(n37738) );
  NANDN U46814 ( .A(n37744), .B(n37745), .Z(n37664) );
  ANDN U46815 ( .B(n37746), .A(n37747), .Z(n37658) );
  XNOR U46816 ( .A(n37649), .B(n37748), .Z(n37654) );
  XNOR U46817 ( .A(n37647), .B(n37651), .Z(n37748) );
  AND U46818 ( .A(n37749), .B(n37750), .Z(n37651) );
  NAND U46819 ( .A(n37751), .B(n37752), .Z(n37750) );
  NAND U46820 ( .A(n37753), .B(n37754), .Z(n37749) );
  AND U46821 ( .A(n37755), .B(n37756), .Z(n37647) );
  NAND U46822 ( .A(n37757), .B(n37758), .Z(n37756) );
  NAND U46823 ( .A(n37759), .B(n37760), .Z(n37755) );
  AND U46824 ( .A(n37761), .B(n37762), .Z(n37649) );
  XOR U46825 ( .A(n37729), .B(n37728), .Z(N62035) );
  XNOR U46826 ( .A(n37746), .B(n37747), .Z(n37728) );
  XNOR U46827 ( .A(n37761), .B(n37762), .Z(n37747) );
  XOR U46828 ( .A(n37758), .B(n37757), .Z(n37762) );
  XOR U46829 ( .A(y[2676]), .B(x[2676]), .Z(n37757) );
  XOR U46830 ( .A(n37760), .B(n37759), .Z(n37758) );
  XOR U46831 ( .A(y[2678]), .B(x[2678]), .Z(n37759) );
  XOR U46832 ( .A(y[2677]), .B(x[2677]), .Z(n37760) );
  XOR U46833 ( .A(n37752), .B(n37751), .Z(n37761) );
  XOR U46834 ( .A(n37754), .B(n37753), .Z(n37751) );
  XOR U46835 ( .A(y[2675]), .B(x[2675]), .Z(n37753) );
  XOR U46836 ( .A(y[2674]), .B(x[2674]), .Z(n37754) );
  XOR U46837 ( .A(y[2673]), .B(x[2673]), .Z(n37752) );
  XNOR U46838 ( .A(n37745), .B(n37744), .Z(n37746) );
  XNOR U46839 ( .A(n37741), .B(n37740), .Z(n37744) );
  XOR U46840 ( .A(n37743), .B(n37742), .Z(n37740) );
  XOR U46841 ( .A(y[2672]), .B(x[2672]), .Z(n37742) );
  XOR U46842 ( .A(y[2671]), .B(x[2671]), .Z(n37743) );
  XOR U46843 ( .A(y[2670]), .B(x[2670]), .Z(n37741) );
  XOR U46844 ( .A(n37735), .B(n37734), .Z(n37745) );
  XOR U46845 ( .A(n37737), .B(n37736), .Z(n37734) );
  XOR U46846 ( .A(y[2669]), .B(x[2669]), .Z(n37736) );
  XOR U46847 ( .A(y[2668]), .B(x[2668]), .Z(n37737) );
  XOR U46848 ( .A(y[2667]), .B(x[2667]), .Z(n37735) );
  XNOR U46849 ( .A(n37711), .B(n37712), .Z(n37729) );
  XNOR U46850 ( .A(n37726), .B(n37727), .Z(n37712) );
  XOR U46851 ( .A(n37723), .B(n37722), .Z(n37727) );
  XOR U46852 ( .A(y[2664]), .B(x[2664]), .Z(n37722) );
  XOR U46853 ( .A(n37725), .B(n37724), .Z(n37723) );
  XOR U46854 ( .A(y[2666]), .B(x[2666]), .Z(n37724) );
  XOR U46855 ( .A(y[2665]), .B(x[2665]), .Z(n37725) );
  XOR U46856 ( .A(n37717), .B(n37716), .Z(n37726) );
  XOR U46857 ( .A(n37719), .B(n37718), .Z(n37716) );
  XOR U46858 ( .A(y[2663]), .B(x[2663]), .Z(n37718) );
  XOR U46859 ( .A(y[2662]), .B(x[2662]), .Z(n37719) );
  XOR U46860 ( .A(y[2661]), .B(x[2661]), .Z(n37717) );
  XNOR U46861 ( .A(n37710), .B(n37709), .Z(n37711) );
  XNOR U46862 ( .A(n37706), .B(n37705), .Z(n37709) );
  XOR U46863 ( .A(n37708), .B(n37707), .Z(n37705) );
  XOR U46864 ( .A(y[2660]), .B(x[2660]), .Z(n37707) );
  XOR U46865 ( .A(y[2659]), .B(x[2659]), .Z(n37708) );
  XOR U46866 ( .A(y[2658]), .B(x[2658]), .Z(n37706) );
  XOR U46867 ( .A(n37700), .B(n37699), .Z(n37710) );
  XOR U46868 ( .A(n37702), .B(n37701), .Z(n37699) );
  XOR U46869 ( .A(y[2657]), .B(x[2657]), .Z(n37701) );
  XOR U46870 ( .A(y[2656]), .B(x[2656]), .Z(n37702) );
  XOR U46871 ( .A(y[2655]), .B(x[2655]), .Z(n37700) );
  NAND U46872 ( .A(n37763), .B(n37764), .Z(N62026) );
  NAND U46873 ( .A(n37765), .B(n37766), .Z(n37764) );
  NANDN U46874 ( .A(n37767), .B(n37768), .Z(n37766) );
  NANDN U46875 ( .A(n37768), .B(n37767), .Z(n37763) );
  XOR U46876 ( .A(n37767), .B(n37769), .Z(N62025) );
  XNOR U46877 ( .A(n37765), .B(n37768), .Z(n37769) );
  NAND U46878 ( .A(n37770), .B(n37771), .Z(n37768) );
  NAND U46879 ( .A(n37772), .B(n37773), .Z(n37771) );
  NANDN U46880 ( .A(n37774), .B(n37775), .Z(n37773) );
  NANDN U46881 ( .A(n37775), .B(n37774), .Z(n37770) );
  AND U46882 ( .A(n37776), .B(n37777), .Z(n37765) );
  NAND U46883 ( .A(n37778), .B(n37779), .Z(n37777) );
  NANDN U46884 ( .A(n37780), .B(n37781), .Z(n37779) );
  NANDN U46885 ( .A(n37781), .B(n37780), .Z(n37776) );
  IV U46886 ( .A(n37782), .Z(n37781) );
  AND U46887 ( .A(n37783), .B(n37784), .Z(n37767) );
  NAND U46888 ( .A(n37785), .B(n37786), .Z(n37784) );
  NANDN U46889 ( .A(n37787), .B(n37788), .Z(n37786) );
  NANDN U46890 ( .A(n37788), .B(n37787), .Z(n37783) );
  XOR U46891 ( .A(n37780), .B(n37789), .Z(N62024) );
  XNOR U46892 ( .A(n37778), .B(n37782), .Z(n37789) );
  XOR U46893 ( .A(n37775), .B(n37790), .Z(n37782) );
  XNOR U46894 ( .A(n37772), .B(n37774), .Z(n37790) );
  AND U46895 ( .A(n37791), .B(n37792), .Z(n37774) );
  NANDN U46896 ( .A(n37793), .B(n37794), .Z(n37792) );
  OR U46897 ( .A(n37795), .B(n37796), .Z(n37794) );
  IV U46898 ( .A(n37797), .Z(n37796) );
  NANDN U46899 ( .A(n37797), .B(n37795), .Z(n37791) );
  AND U46900 ( .A(n37798), .B(n37799), .Z(n37772) );
  NAND U46901 ( .A(n37800), .B(n37801), .Z(n37799) );
  NANDN U46902 ( .A(n37802), .B(n37803), .Z(n37801) );
  NANDN U46903 ( .A(n37803), .B(n37802), .Z(n37798) );
  IV U46904 ( .A(n37804), .Z(n37803) );
  NAND U46905 ( .A(n37805), .B(n37806), .Z(n37775) );
  NANDN U46906 ( .A(n37807), .B(n37808), .Z(n37806) );
  NANDN U46907 ( .A(n37809), .B(n37810), .Z(n37808) );
  NANDN U46908 ( .A(n37810), .B(n37809), .Z(n37805) );
  IV U46909 ( .A(n37811), .Z(n37809) );
  AND U46910 ( .A(n37812), .B(n37813), .Z(n37778) );
  NAND U46911 ( .A(n37814), .B(n37815), .Z(n37813) );
  NANDN U46912 ( .A(n37816), .B(n37817), .Z(n37815) );
  NANDN U46913 ( .A(n37817), .B(n37816), .Z(n37812) );
  XOR U46914 ( .A(n37788), .B(n37818), .Z(n37780) );
  XNOR U46915 ( .A(n37785), .B(n37787), .Z(n37818) );
  AND U46916 ( .A(n37819), .B(n37820), .Z(n37787) );
  NANDN U46917 ( .A(n37821), .B(n37822), .Z(n37820) );
  OR U46918 ( .A(n37823), .B(n37824), .Z(n37822) );
  IV U46919 ( .A(n37825), .Z(n37824) );
  NANDN U46920 ( .A(n37825), .B(n37823), .Z(n37819) );
  AND U46921 ( .A(n37826), .B(n37827), .Z(n37785) );
  NAND U46922 ( .A(n37828), .B(n37829), .Z(n37827) );
  NANDN U46923 ( .A(n37830), .B(n37831), .Z(n37829) );
  NANDN U46924 ( .A(n37831), .B(n37830), .Z(n37826) );
  IV U46925 ( .A(n37832), .Z(n37831) );
  NAND U46926 ( .A(n37833), .B(n37834), .Z(n37788) );
  NANDN U46927 ( .A(n37835), .B(n37836), .Z(n37834) );
  NANDN U46928 ( .A(n37837), .B(n37838), .Z(n37836) );
  NANDN U46929 ( .A(n37838), .B(n37837), .Z(n37833) );
  IV U46930 ( .A(n37839), .Z(n37837) );
  XOR U46931 ( .A(n37814), .B(n37840), .Z(N62023) );
  XNOR U46932 ( .A(n37817), .B(n37816), .Z(n37840) );
  XNOR U46933 ( .A(n37828), .B(n37841), .Z(n37816) );
  XNOR U46934 ( .A(n37832), .B(n37830), .Z(n37841) );
  XOR U46935 ( .A(n37838), .B(n37842), .Z(n37830) );
  XNOR U46936 ( .A(n37835), .B(n37839), .Z(n37842) );
  AND U46937 ( .A(n37843), .B(n37844), .Z(n37839) );
  NAND U46938 ( .A(n37845), .B(n37846), .Z(n37844) );
  NAND U46939 ( .A(n37847), .B(n37848), .Z(n37843) );
  AND U46940 ( .A(n37849), .B(n37850), .Z(n37835) );
  NAND U46941 ( .A(n37851), .B(n37852), .Z(n37850) );
  NAND U46942 ( .A(n37853), .B(n37854), .Z(n37849) );
  NANDN U46943 ( .A(n37855), .B(n37856), .Z(n37838) );
  ANDN U46944 ( .B(n37857), .A(n37858), .Z(n37832) );
  XNOR U46945 ( .A(n37823), .B(n37859), .Z(n37828) );
  XNOR U46946 ( .A(n37821), .B(n37825), .Z(n37859) );
  AND U46947 ( .A(n37860), .B(n37861), .Z(n37825) );
  NAND U46948 ( .A(n37862), .B(n37863), .Z(n37861) );
  NAND U46949 ( .A(n37864), .B(n37865), .Z(n37860) );
  AND U46950 ( .A(n37866), .B(n37867), .Z(n37821) );
  NAND U46951 ( .A(n37868), .B(n37869), .Z(n37867) );
  NAND U46952 ( .A(n37870), .B(n37871), .Z(n37866) );
  AND U46953 ( .A(n37872), .B(n37873), .Z(n37823) );
  NAND U46954 ( .A(n37874), .B(n37875), .Z(n37817) );
  XNOR U46955 ( .A(n37800), .B(n37876), .Z(n37814) );
  XNOR U46956 ( .A(n37804), .B(n37802), .Z(n37876) );
  XOR U46957 ( .A(n37810), .B(n37877), .Z(n37802) );
  XNOR U46958 ( .A(n37807), .B(n37811), .Z(n37877) );
  AND U46959 ( .A(n37878), .B(n37879), .Z(n37811) );
  NAND U46960 ( .A(n37880), .B(n37881), .Z(n37879) );
  NAND U46961 ( .A(n37882), .B(n37883), .Z(n37878) );
  AND U46962 ( .A(n37884), .B(n37885), .Z(n37807) );
  NAND U46963 ( .A(n37886), .B(n37887), .Z(n37885) );
  NAND U46964 ( .A(n37888), .B(n37889), .Z(n37884) );
  NANDN U46965 ( .A(n37890), .B(n37891), .Z(n37810) );
  ANDN U46966 ( .B(n37892), .A(n37893), .Z(n37804) );
  XNOR U46967 ( .A(n37795), .B(n37894), .Z(n37800) );
  XNOR U46968 ( .A(n37793), .B(n37797), .Z(n37894) );
  AND U46969 ( .A(n37895), .B(n37896), .Z(n37797) );
  NAND U46970 ( .A(n37897), .B(n37898), .Z(n37896) );
  NAND U46971 ( .A(n37899), .B(n37900), .Z(n37895) );
  AND U46972 ( .A(n37901), .B(n37902), .Z(n37793) );
  NAND U46973 ( .A(n37903), .B(n37904), .Z(n37902) );
  NAND U46974 ( .A(n37905), .B(n37906), .Z(n37901) );
  AND U46975 ( .A(n37907), .B(n37908), .Z(n37795) );
  XOR U46976 ( .A(n37875), .B(n37874), .Z(N62022) );
  XNOR U46977 ( .A(n37892), .B(n37893), .Z(n37874) );
  XNOR U46978 ( .A(n37907), .B(n37908), .Z(n37893) );
  XOR U46979 ( .A(n37904), .B(n37903), .Z(n37908) );
  XOR U46980 ( .A(y[2652]), .B(x[2652]), .Z(n37903) );
  XOR U46981 ( .A(n37906), .B(n37905), .Z(n37904) );
  XOR U46982 ( .A(y[2654]), .B(x[2654]), .Z(n37905) );
  XOR U46983 ( .A(y[2653]), .B(x[2653]), .Z(n37906) );
  XOR U46984 ( .A(n37898), .B(n37897), .Z(n37907) );
  XOR U46985 ( .A(n37900), .B(n37899), .Z(n37897) );
  XOR U46986 ( .A(y[2651]), .B(x[2651]), .Z(n37899) );
  XOR U46987 ( .A(y[2650]), .B(x[2650]), .Z(n37900) );
  XOR U46988 ( .A(y[2649]), .B(x[2649]), .Z(n37898) );
  XNOR U46989 ( .A(n37891), .B(n37890), .Z(n37892) );
  XNOR U46990 ( .A(n37887), .B(n37886), .Z(n37890) );
  XOR U46991 ( .A(n37889), .B(n37888), .Z(n37886) );
  XOR U46992 ( .A(y[2648]), .B(x[2648]), .Z(n37888) );
  XOR U46993 ( .A(y[2647]), .B(x[2647]), .Z(n37889) );
  XOR U46994 ( .A(y[2646]), .B(x[2646]), .Z(n37887) );
  XOR U46995 ( .A(n37881), .B(n37880), .Z(n37891) );
  XOR U46996 ( .A(n37883), .B(n37882), .Z(n37880) );
  XOR U46997 ( .A(y[2645]), .B(x[2645]), .Z(n37882) );
  XOR U46998 ( .A(y[2644]), .B(x[2644]), .Z(n37883) );
  XOR U46999 ( .A(y[2643]), .B(x[2643]), .Z(n37881) );
  XNOR U47000 ( .A(n37857), .B(n37858), .Z(n37875) );
  XNOR U47001 ( .A(n37872), .B(n37873), .Z(n37858) );
  XOR U47002 ( .A(n37869), .B(n37868), .Z(n37873) );
  XOR U47003 ( .A(y[2640]), .B(x[2640]), .Z(n37868) );
  XOR U47004 ( .A(n37871), .B(n37870), .Z(n37869) );
  XOR U47005 ( .A(y[2642]), .B(x[2642]), .Z(n37870) );
  XOR U47006 ( .A(y[2641]), .B(x[2641]), .Z(n37871) );
  XOR U47007 ( .A(n37863), .B(n37862), .Z(n37872) );
  XOR U47008 ( .A(n37865), .B(n37864), .Z(n37862) );
  XOR U47009 ( .A(y[2639]), .B(x[2639]), .Z(n37864) );
  XOR U47010 ( .A(y[2638]), .B(x[2638]), .Z(n37865) );
  XOR U47011 ( .A(y[2637]), .B(x[2637]), .Z(n37863) );
  XNOR U47012 ( .A(n37856), .B(n37855), .Z(n37857) );
  XNOR U47013 ( .A(n37852), .B(n37851), .Z(n37855) );
  XOR U47014 ( .A(n37854), .B(n37853), .Z(n37851) );
  XOR U47015 ( .A(y[2636]), .B(x[2636]), .Z(n37853) );
  XOR U47016 ( .A(y[2635]), .B(x[2635]), .Z(n37854) );
  XOR U47017 ( .A(y[2634]), .B(x[2634]), .Z(n37852) );
  XOR U47018 ( .A(n37846), .B(n37845), .Z(n37856) );
  XOR U47019 ( .A(n37848), .B(n37847), .Z(n37845) );
  XOR U47020 ( .A(y[2633]), .B(x[2633]), .Z(n37847) );
  XOR U47021 ( .A(y[2632]), .B(x[2632]), .Z(n37848) );
  XOR U47022 ( .A(y[2631]), .B(x[2631]), .Z(n37846) );
  NAND U47023 ( .A(n37909), .B(n37910), .Z(N62013) );
  NAND U47024 ( .A(n37911), .B(n37912), .Z(n37910) );
  NANDN U47025 ( .A(n37913), .B(n37914), .Z(n37912) );
  NANDN U47026 ( .A(n37914), .B(n37913), .Z(n37909) );
  XOR U47027 ( .A(n37913), .B(n37915), .Z(N62012) );
  XNOR U47028 ( .A(n37911), .B(n37914), .Z(n37915) );
  NAND U47029 ( .A(n37916), .B(n37917), .Z(n37914) );
  NAND U47030 ( .A(n37918), .B(n37919), .Z(n37917) );
  NANDN U47031 ( .A(n37920), .B(n37921), .Z(n37919) );
  NANDN U47032 ( .A(n37921), .B(n37920), .Z(n37916) );
  AND U47033 ( .A(n37922), .B(n37923), .Z(n37911) );
  NAND U47034 ( .A(n37924), .B(n37925), .Z(n37923) );
  NANDN U47035 ( .A(n37926), .B(n37927), .Z(n37925) );
  NANDN U47036 ( .A(n37927), .B(n37926), .Z(n37922) );
  IV U47037 ( .A(n37928), .Z(n37927) );
  AND U47038 ( .A(n37929), .B(n37930), .Z(n37913) );
  NAND U47039 ( .A(n37931), .B(n37932), .Z(n37930) );
  NANDN U47040 ( .A(n37933), .B(n37934), .Z(n37932) );
  NANDN U47041 ( .A(n37934), .B(n37933), .Z(n37929) );
  XOR U47042 ( .A(n37926), .B(n37935), .Z(N62011) );
  XNOR U47043 ( .A(n37924), .B(n37928), .Z(n37935) );
  XOR U47044 ( .A(n37921), .B(n37936), .Z(n37928) );
  XNOR U47045 ( .A(n37918), .B(n37920), .Z(n37936) );
  AND U47046 ( .A(n37937), .B(n37938), .Z(n37920) );
  NANDN U47047 ( .A(n37939), .B(n37940), .Z(n37938) );
  OR U47048 ( .A(n37941), .B(n37942), .Z(n37940) );
  IV U47049 ( .A(n37943), .Z(n37942) );
  NANDN U47050 ( .A(n37943), .B(n37941), .Z(n37937) );
  AND U47051 ( .A(n37944), .B(n37945), .Z(n37918) );
  NAND U47052 ( .A(n37946), .B(n37947), .Z(n37945) );
  NANDN U47053 ( .A(n37948), .B(n37949), .Z(n37947) );
  NANDN U47054 ( .A(n37949), .B(n37948), .Z(n37944) );
  IV U47055 ( .A(n37950), .Z(n37949) );
  NAND U47056 ( .A(n37951), .B(n37952), .Z(n37921) );
  NANDN U47057 ( .A(n37953), .B(n37954), .Z(n37952) );
  NANDN U47058 ( .A(n37955), .B(n37956), .Z(n37954) );
  NANDN U47059 ( .A(n37956), .B(n37955), .Z(n37951) );
  IV U47060 ( .A(n37957), .Z(n37955) );
  AND U47061 ( .A(n37958), .B(n37959), .Z(n37924) );
  NAND U47062 ( .A(n37960), .B(n37961), .Z(n37959) );
  NANDN U47063 ( .A(n37962), .B(n37963), .Z(n37961) );
  NANDN U47064 ( .A(n37963), .B(n37962), .Z(n37958) );
  XOR U47065 ( .A(n37934), .B(n37964), .Z(n37926) );
  XNOR U47066 ( .A(n37931), .B(n37933), .Z(n37964) );
  AND U47067 ( .A(n37965), .B(n37966), .Z(n37933) );
  NANDN U47068 ( .A(n37967), .B(n37968), .Z(n37966) );
  OR U47069 ( .A(n37969), .B(n37970), .Z(n37968) );
  IV U47070 ( .A(n37971), .Z(n37970) );
  NANDN U47071 ( .A(n37971), .B(n37969), .Z(n37965) );
  AND U47072 ( .A(n37972), .B(n37973), .Z(n37931) );
  NAND U47073 ( .A(n37974), .B(n37975), .Z(n37973) );
  NANDN U47074 ( .A(n37976), .B(n37977), .Z(n37975) );
  NANDN U47075 ( .A(n37977), .B(n37976), .Z(n37972) );
  IV U47076 ( .A(n37978), .Z(n37977) );
  NAND U47077 ( .A(n37979), .B(n37980), .Z(n37934) );
  NANDN U47078 ( .A(n37981), .B(n37982), .Z(n37980) );
  NANDN U47079 ( .A(n37983), .B(n37984), .Z(n37982) );
  NANDN U47080 ( .A(n37984), .B(n37983), .Z(n37979) );
  IV U47081 ( .A(n37985), .Z(n37983) );
  XOR U47082 ( .A(n37960), .B(n37986), .Z(N62010) );
  XNOR U47083 ( .A(n37963), .B(n37962), .Z(n37986) );
  XNOR U47084 ( .A(n37974), .B(n37987), .Z(n37962) );
  XNOR U47085 ( .A(n37978), .B(n37976), .Z(n37987) );
  XOR U47086 ( .A(n37984), .B(n37988), .Z(n37976) );
  XNOR U47087 ( .A(n37981), .B(n37985), .Z(n37988) );
  AND U47088 ( .A(n37989), .B(n37990), .Z(n37985) );
  NAND U47089 ( .A(n37991), .B(n37992), .Z(n37990) );
  NAND U47090 ( .A(n37993), .B(n37994), .Z(n37989) );
  AND U47091 ( .A(n37995), .B(n37996), .Z(n37981) );
  NAND U47092 ( .A(n37997), .B(n37998), .Z(n37996) );
  NAND U47093 ( .A(n37999), .B(n38000), .Z(n37995) );
  NANDN U47094 ( .A(n38001), .B(n38002), .Z(n37984) );
  ANDN U47095 ( .B(n38003), .A(n38004), .Z(n37978) );
  XNOR U47096 ( .A(n37969), .B(n38005), .Z(n37974) );
  XNOR U47097 ( .A(n37967), .B(n37971), .Z(n38005) );
  AND U47098 ( .A(n38006), .B(n38007), .Z(n37971) );
  NAND U47099 ( .A(n38008), .B(n38009), .Z(n38007) );
  NAND U47100 ( .A(n38010), .B(n38011), .Z(n38006) );
  AND U47101 ( .A(n38012), .B(n38013), .Z(n37967) );
  NAND U47102 ( .A(n38014), .B(n38015), .Z(n38013) );
  NAND U47103 ( .A(n38016), .B(n38017), .Z(n38012) );
  AND U47104 ( .A(n38018), .B(n38019), .Z(n37969) );
  NAND U47105 ( .A(n38020), .B(n38021), .Z(n37963) );
  XNOR U47106 ( .A(n37946), .B(n38022), .Z(n37960) );
  XNOR U47107 ( .A(n37950), .B(n37948), .Z(n38022) );
  XOR U47108 ( .A(n37956), .B(n38023), .Z(n37948) );
  XNOR U47109 ( .A(n37953), .B(n37957), .Z(n38023) );
  AND U47110 ( .A(n38024), .B(n38025), .Z(n37957) );
  NAND U47111 ( .A(n38026), .B(n38027), .Z(n38025) );
  NAND U47112 ( .A(n38028), .B(n38029), .Z(n38024) );
  AND U47113 ( .A(n38030), .B(n38031), .Z(n37953) );
  NAND U47114 ( .A(n38032), .B(n38033), .Z(n38031) );
  NAND U47115 ( .A(n38034), .B(n38035), .Z(n38030) );
  NANDN U47116 ( .A(n38036), .B(n38037), .Z(n37956) );
  ANDN U47117 ( .B(n38038), .A(n38039), .Z(n37950) );
  XNOR U47118 ( .A(n37941), .B(n38040), .Z(n37946) );
  XNOR U47119 ( .A(n37939), .B(n37943), .Z(n38040) );
  AND U47120 ( .A(n38041), .B(n38042), .Z(n37943) );
  NAND U47121 ( .A(n38043), .B(n38044), .Z(n38042) );
  NAND U47122 ( .A(n38045), .B(n38046), .Z(n38041) );
  AND U47123 ( .A(n38047), .B(n38048), .Z(n37939) );
  NAND U47124 ( .A(n38049), .B(n38050), .Z(n38048) );
  NAND U47125 ( .A(n38051), .B(n38052), .Z(n38047) );
  AND U47126 ( .A(n38053), .B(n38054), .Z(n37941) );
  XOR U47127 ( .A(n38021), .B(n38020), .Z(N62009) );
  XNOR U47128 ( .A(n38038), .B(n38039), .Z(n38020) );
  XNOR U47129 ( .A(n38053), .B(n38054), .Z(n38039) );
  XOR U47130 ( .A(n38050), .B(n38049), .Z(n38054) );
  XOR U47131 ( .A(y[2628]), .B(x[2628]), .Z(n38049) );
  XOR U47132 ( .A(n38052), .B(n38051), .Z(n38050) );
  XOR U47133 ( .A(y[2630]), .B(x[2630]), .Z(n38051) );
  XOR U47134 ( .A(y[2629]), .B(x[2629]), .Z(n38052) );
  XOR U47135 ( .A(n38044), .B(n38043), .Z(n38053) );
  XOR U47136 ( .A(n38046), .B(n38045), .Z(n38043) );
  XOR U47137 ( .A(y[2627]), .B(x[2627]), .Z(n38045) );
  XOR U47138 ( .A(y[2626]), .B(x[2626]), .Z(n38046) );
  XOR U47139 ( .A(y[2625]), .B(x[2625]), .Z(n38044) );
  XNOR U47140 ( .A(n38037), .B(n38036), .Z(n38038) );
  XNOR U47141 ( .A(n38033), .B(n38032), .Z(n38036) );
  XOR U47142 ( .A(n38035), .B(n38034), .Z(n38032) );
  XOR U47143 ( .A(y[2624]), .B(x[2624]), .Z(n38034) );
  XOR U47144 ( .A(y[2623]), .B(x[2623]), .Z(n38035) );
  XOR U47145 ( .A(y[2622]), .B(x[2622]), .Z(n38033) );
  XOR U47146 ( .A(n38027), .B(n38026), .Z(n38037) );
  XOR U47147 ( .A(n38029), .B(n38028), .Z(n38026) );
  XOR U47148 ( .A(y[2621]), .B(x[2621]), .Z(n38028) );
  XOR U47149 ( .A(y[2620]), .B(x[2620]), .Z(n38029) );
  XOR U47150 ( .A(y[2619]), .B(x[2619]), .Z(n38027) );
  XNOR U47151 ( .A(n38003), .B(n38004), .Z(n38021) );
  XNOR U47152 ( .A(n38018), .B(n38019), .Z(n38004) );
  XOR U47153 ( .A(n38015), .B(n38014), .Z(n38019) );
  XOR U47154 ( .A(y[2616]), .B(x[2616]), .Z(n38014) );
  XOR U47155 ( .A(n38017), .B(n38016), .Z(n38015) );
  XOR U47156 ( .A(y[2618]), .B(x[2618]), .Z(n38016) );
  XOR U47157 ( .A(y[2617]), .B(x[2617]), .Z(n38017) );
  XOR U47158 ( .A(n38009), .B(n38008), .Z(n38018) );
  XOR U47159 ( .A(n38011), .B(n38010), .Z(n38008) );
  XOR U47160 ( .A(y[2615]), .B(x[2615]), .Z(n38010) );
  XOR U47161 ( .A(y[2614]), .B(x[2614]), .Z(n38011) );
  XOR U47162 ( .A(y[2613]), .B(x[2613]), .Z(n38009) );
  XNOR U47163 ( .A(n38002), .B(n38001), .Z(n38003) );
  XNOR U47164 ( .A(n37998), .B(n37997), .Z(n38001) );
  XOR U47165 ( .A(n38000), .B(n37999), .Z(n37997) );
  XOR U47166 ( .A(y[2612]), .B(x[2612]), .Z(n37999) );
  XOR U47167 ( .A(y[2611]), .B(x[2611]), .Z(n38000) );
  XOR U47168 ( .A(y[2610]), .B(x[2610]), .Z(n37998) );
  XOR U47169 ( .A(n37992), .B(n37991), .Z(n38002) );
  XOR U47170 ( .A(n37994), .B(n37993), .Z(n37991) );
  XOR U47171 ( .A(y[2609]), .B(x[2609]), .Z(n37993) );
  XOR U47172 ( .A(y[2608]), .B(x[2608]), .Z(n37994) );
  XOR U47173 ( .A(y[2607]), .B(x[2607]), .Z(n37992) );
  NAND U47174 ( .A(n38055), .B(n38056), .Z(N62000) );
  NAND U47175 ( .A(n38057), .B(n38058), .Z(n38056) );
  NANDN U47176 ( .A(n38059), .B(n38060), .Z(n38058) );
  NANDN U47177 ( .A(n38060), .B(n38059), .Z(n38055) );
  XOR U47178 ( .A(n38059), .B(n38061), .Z(N61999) );
  XNOR U47179 ( .A(n38057), .B(n38060), .Z(n38061) );
  NAND U47180 ( .A(n38062), .B(n38063), .Z(n38060) );
  NAND U47181 ( .A(n38064), .B(n38065), .Z(n38063) );
  NANDN U47182 ( .A(n38066), .B(n38067), .Z(n38065) );
  NANDN U47183 ( .A(n38067), .B(n38066), .Z(n38062) );
  AND U47184 ( .A(n38068), .B(n38069), .Z(n38057) );
  NAND U47185 ( .A(n38070), .B(n38071), .Z(n38069) );
  NANDN U47186 ( .A(n38072), .B(n38073), .Z(n38071) );
  NANDN U47187 ( .A(n38073), .B(n38072), .Z(n38068) );
  IV U47188 ( .A(n38074), .Z(n38073) );
  AND U47189 ( .A(n38075), .B(n38076), .Z(n38059) );
  NAND U47190 ( .A(n38077), .B(n38078), .Z(n38076) );
  NANDN U47191 ( .A(n38079), .B(n38080), .Z(n38078) );
  NANDN U47192 ( .A(n38080), .B(n38079), .Z(n38075) );
  XOR U47193 ( .A(n38072), .B(n38081), .Z(N61998) );
  XNOR U47194 ( .A(n38070), .B(n38074), .Z(n38081) );
  XOR U47195 ( .A(n38067), .B(n38082), .Z(n38074) );
  XNOR U47196 ( .A(n38064), .B(n38066), .Z(n38082) );
  AND U47197 ( .A(n38083), .B(n38084), .Z(n38066) );
  NANDN U47198 ( .A(n38085), .B(n38086), .Z(n38084) );
  OR U47199 ( .A(n38087), .B(n38088), .Z(n38086) );
  IV U47200 ( .A(n38089), .Z(n38088) );
  NANDN U47201 ( .A(n38089), .B(n38087), .Z(n38083) );
  AND U47202 ( .A(n38090), .B(n38091), .Z(n38064) );
  NAND U47203 ( .A(n38092), .B(n38093), .Z(n38091) );
  NANDN U47204 ( .A(n38094), .B(n38095), .Z(n38093) );
  NANDN U47205 ( .A(n38095), .B(n38094), .Z(n38090) );
  IV U47206 ( .A(n38096), .Z(n38095) );
  NAND U47207 ( .A(n38097), .B(n38098), .Z(n38067) );
  NANDN U47208 ( .A(n38099), .B(n38100), .Z(n38098) );
  NANDN U47209 ( .A(n38101), .B(n38102), .Z(n38100) );
  NANDN U47210 ( .A(n38102), .B(n38101), .Z(n38097) );
  IV U47211 ( .A(n38103), .Z(n38101) );
  AND U47212 ( .A(n38104), .B(n38105), .Z(n38070) );
  NAND U47213 ( .A(n38106), .B(n38107), .Z(n38105) );
  NANDN U47214 ( .A(n38108), .B(n38109), .Z(n38107) );
  NANDN U47215 ( .A(n38109), .B(n38108), .Z(n38104) );
  XOR U47216 ( .A(n38080), .B(n38110), .Z(n38072) );
  XNOR U47217 ( .A(n38077), .B(n38079), .Z(n38110) );
  AND U47218 ( .A(n38111), .B(n38112), .Z(n38079) );
  NANDN U47219 ( .A(n38113), .B(n38114), .Z(n38112) );
  OR U47220 ( .A(n38115), .B(n38116), .Z(n38114) );
  IV U47221 ( .A(n38117), .Z(n38116) );
  NANDN U47222 ( .A(n38117), .B(n38115), .Z(n38111) );
  AND U47223 ( .A(n38118), .B(n38119), .Z(n38077) );
  NAND U47224 ( .A(n38120), .B(n38121), .Z(n38119) );
  NANDN U47225 ( .A(n38122), .B(n38123), .Z(n38121) );
  NANDN U47226 ( .A(n38123), .B(n38122), .Z(n38118) );
  IV U47227 ( .A(n38124), .Z(n38123) );
  NAND U47228 ( .A(n38125), .B(n38126), .Z(n38080) );
  NANDN U47229 ( .A(n38127), .B(n38128), .Z(n38126) );
  NANDN U47230 ( .A(n38129), .B(n38130), .Z(n38128) );
  NANDN U47231 ( .A(n38130), .B(n38129), .Z(n38125) );
  IV U47232 ( .A(n38131), .Z(n38129) );
  XOR U47233 ( .A(n38106), .B(n38132), .Z(N61997) );
  XNOR U47234 ( .A(n38109), .B(n38108), .Z(n38132) );
  XNOR U47235 ( .A(n38120), .B(n38133), .Z(n38108) );
  XNOR U47236 ( .A(n38124), .B(n38122), .Z(n38133) );
  XOR U47237 ( .A(n38130), .B(n38134), .Z(n38122) );
  XNOR U47238 ( .A(n38127), .B(n38131), .Z(n38134) );
  AND U47239 ( .A(n38135), .B(n38136), .Z(n38131) );
  NAND U47240 ( .A(n38137), .B(n38138), .Z(n38136) );
  NAND U47241 ( .A(n38139), .B(n38140), .Z(n38135) );
  AND U47242 ( .A(n38141), .B(n38142), .Z(n38127) );
  NAND U47243 ( .A(n38143), .B(n38144), .Z(n38142) );
  NAND U47244 ( .A(n38145), .B(n38146), .Z(n38141) );
  NANDN U47245 ( .A(n38147), .B(n38148), .Z(n38130) );
  ANDN U47246 ( .B(n38149), .A(n38150), .Z(n38124) );
  XNOR U47247 ( .A(n38115), .B(n38151), .Z(n38120) );
  XNOR U47248 ( .A(n38113), .B(n38117), .Z(n38151) );
  AND U47249 ( .A(n38152), .B(n38153), .Z(n38117) );
  NAND U47250 ( .A(n38154), .B(n38155), .Z(n38153) );
  NAND U47251 ( .A(n38156), .B(n38157), .Z(n38152) );
  AND U47252 ( .A(n38158), .B(n38159), .Z(n38113) );
  NAND U47253 ( .A(n38160), .B(n38161), .Z(n38159) );
  NAND U47254 ( .A(n38162), .B(n38163), .Z(n38158) );
  AND U47255 ( .A(n38164), .B(n38165), .Z(n38115) );
  NAND U47256 ( .A(n38166), .B(n38167), .Z(n38109) );
  XNOR U47257 ( .A(n38092), .B(n38168), .Z(n38106) );
  XNOR U47258 ( .A(n38096), .B(n38094), .Z(n38168) );
  XOR U47259 ( .A(n38102), .B(n38169), .Z(n38094) );
  XNOR U47260 ( .A(n38099), .B(n38103), .Z(n38169) );
  AND U47261 ( .A(n38170), .B(n38171), .Z(n38103) );
  NAND U47262 ( .A(n38172), .B(n38173), .Z(n38171) );
  NAND U47263 ( .A(n38174), .B(n38175), .Z(n38170) );
  AND U47264 ( .A(n38176), .B(n38177), .Z(n38099) );
  NAND U47265 ( .A(n38178), .B(n38179), .Z(n38177) );
  NAND U47266 ( .A(n38180), .B(n38181), .Z(n38176) );
  NANDN U47267 ( .A(n38182), .B(n38183), .Z(n38102) );
  ANDN U47268 ( .B(n38184), .A(n38185), .Z(n38096) );
  XNOR U47269 ( .A(n38087), .B(n38186), .Z(n38092) );
  XNOR U47270 ( .A(n38085), .B(n38089), .Z(n38186) );
  AND U47271 ( .A(n38187), .B(n38188), .Z(n38089) );
  NAND U47272 ( .A(n38189), .B(n38190), .Z(n38188) );
  NAND U47273 ( .A(n38191), .B(n38192), .Z(n38187) );
  AND U47274 ( .A(n38193), .B(n38194), .Z(n38085) );
  NAND U47275 ( .A(n38195), .B(n38196), .Z(n38194) );
  NAND U47276 ( .A(n38197), .B(n38198), .Z(n38193) );
  AND U47277 ( .A(n38199), .B(n38200), .Z(n38087) );
  XOR U47278 ( .A(n38167), .B(n38166), .Z(N61996) );
  XNOR U47279 ( .A(n38184), .B(n38185), .Z(n38166) );
  XNOR U47280 ( .A(n38199), .B(n38200), .Z(n38185) );
  XOR U47281 ( .A(n38196), .B(n38195), .Z(n38200) );
  XOR U47282 ( .A(y[2604]), .B(x[2604]), .Z(n38195) );
  XOR U47283 ( .A(n38198), .B(n38197), .Z(n38196) );
  XOR U47284 ( .A(y[2606]), .B(x[2606]), .Z(n38197) );
  XOR U47285 ( .A(y[2605]), .B(x[2605]), .Z(n38198) );
  XOR U47286 ( .A(n38190), .B(n38189), .Z(n38199) );
  XOR U47287 ( .A(n38192), .B(n38191), .Z(n38189) );
  XOR U47288 ( .A(y[2603]), .B(x[2603]), .Z(n38191) );
  XOR U47289 ( .A(y[2602]), .B(x[2602]), .Z(n38192) );
  XOR U47290 ( .A(y[2601]), .B(x[2601]), .Z(n38190) );
  XNOR U47291 ( .A(n38183), .B(n38182), .Z(n38184) );
  XNOR U47292 ( .A(n38179), .B(n38178), .Z(n38182) );
  XOR U47293 ( .A(n38181), .B(n38180), .Z(n38178) );
  XOR U47294 ( .A(y[2600]), .B(x[2600]), .Z(n38180) );
  XOR U47295 ( .A(y[2599]), .B(x[2599]), .Z(n38181) );
  XOR U47296 ( .A(y[2598]), .B(x[2598]), .Z(n38179) );
  XOR U47297 ( .A(n38173), .B(n38172), .Z(n38183) );
  XOR U47298 ( .A(n38175), .B(n38174), .Z(n38172) );
  XOR U47299 ( .A(y[2597]), .B(x[2597]), .Z(n38174) );
  XOR U47300 ( .A(y[2596]), .B(x[2596]), .Z(n38175) );
  XOR U47301 ( .A(y[2595]), .B(x[2595]), .Z(n38173) );
  XNOR U47302 ( .A(n38149), .B(n38150), .Z(n38167) );
  XNOR U47303 ( .A(n38164), .B(n38165), .Z(n38150) );
  XOR U47304 ( .A(n38161), .B(n38160), .Z(n38165) );
  XOR U47305 ( .A(y[2592]), .B(x[2592]), .Z(n38160) );
  XOR U47306 ( .A(n38163), .B(n38162), .Z(n38161) );
  XOR U47307 ( .A(y[2594]), .B(x[2594]), .Z(n38162) );
  XOR U47308 ( .A(y[2593]), .B(x[2593]), .Z(n38163) );
  XOR U47309 ( .A(n38155), .B(n38154), .Z(n38164) );
  XOR U47310 ( .A(n38157), .B(n38156), .Z(n38154) );
  XOR U47311 ( .A(y[2591]), .B(x[2591]), .Z(n38156) );
  XOR U47312 ( .A(y[2590]), .B(x[2590]), .Z(n38157) );
  XOR U47313 ( .A(y[2589]), .B(x[2589]), .Z(n38155) );
  XNOR U47314 ( .A(n38148), .B(n38147), .Z(n38149) );
  XNOR U47315 ( .A(n38144), .B(n38143), .Z(n38147) );
  XOR U47316 ( .A(n38146), .B(n38145), .Z(n38143) );
  XOR U47317 ( .A(y[2588]), .B(x[2588]), .Z(n38145) );
  XOR U47318 ( .A(y[2587]), .B(x[2587]), .Z(n38146) );
  XOR U47319 ( .A(y[2586]), .B(x[2586]), .Z(n38144) );
  XOR U47320 ( .A(n38138), .B(n38137), .Z(n38148) );
  XOR U47321 ( .A(n38140), .B(n38139), .Z(n38137) );
  XOR U47322 ( .A(y[2585]), .B(x[2585]), .Z(n38139) );
  XOR U47323 ( .A(y[2584]), .B(x[2584]), .Z(n38140) );
  XOR U47324 ( .A(y[2583]), .B(x[2583]), .Z(n38138) );
  NAND U47325 ( .A(n38201), .B(n38202), .Z(N61987) );
  NAND U47326 ( .A(n38203), .B(n38204), .Z(n38202) );
  NANDN U47327 ( .A(n38205), .B(n38206), .Z(n38204) );
  NANDN U47328 ( .A(n38206), .B(n38205), .Z(n38201) );
  XOR U47329 ( .A(n38205), .B(n38207), .Z(N61986) );
  XNOR U47330 ( .A(n38203), .B(n38206), .Z(n38207) );
  NAND U47331 ( .A(n38208), .B(n38209), .Z(n38206) );
  NAND U47332 ( .A(n38210), .B(n38211), .Z(n38209) );
  NANDN U47333 ( .A(n38212), .B(n38213), .Z(n38211) );
  NANDN U47334 ( .A(n38213), .B(n38212), .Z(n38208) );
  AND U47335 ( .A(n38214), .B(n38215), .Z(n38203) );
  NAND U47336 ( .A(n38216), .B(n38217), .Z(n38215) );
  NANDN U47337 ( .A(n38218), .B(n38219), .Z(n38217) );
  NANDN U47338 ( .A(n38219), .B(n38218), .Z(n38214) );
  IV U47339 ( .A(n38220), .Z(n38219) );
  AND U47340 ( .A(n38221), .B(n38222), .Z(n38205) );
  NAND U47341 ( .A(n38223), .B(n38224), .Z(n38222) );
  NANDN U47342 ( .A(n38225), .B(n38226), .Z(n38224) );
  NANDN U47343 ( .A(n38226), .B(n38225), .Z(n38221) );
  XOR U47344 ( .A(n38218), .B(n38227), .Z(N61985) );
  XNOR U47345 ( .A(n38216), .B(n38220), .Z(n38227) );
  XOR U47346 ( .A(n38213), .B(n38228), .Z(n38220) );
  XNOR U47347 ( .A(n38210), .B(n38212), .Z(n38228) );
  AND U47348 ( .A(n38229), .B(n38230), .Z(n38212) );
  NANDN U47349 ( .A(n38231), .B(n38232), .Z(n38230) );
  OR U47350 ( .A(n38233), .B(n38234), .Z(n38232) );
  IV U47351 ( .A(n38235), .Z(n38234) );
  NANDN U47352 ( .A(n38235), .B(n38233), .Z(n38229) );
  AND U47353 ( .A(n38236), .B(n38237), .Z(n38210) );
  NAND U47354 ( .A(n38238), .B(n38239), .Z(n38237) );
  NANDN U47355 ( .A(n38240), .B(n38241), .Z(n38239) );
  NANDN U47356 ( .A(n38241), .B(n38240), .Z(n38236) );
  IV U47357 ( .A(n38242), .Z(n38241) );
  NAND U47358 ( .A(n38243), .B(n38244), .Z(n38213) );
  NANDN U47359 ( .A(n38245), .B(n38246), .Z(n38244) );
  NANDN U47360 ( .A(n38247), .B(n38248), .Z(n38246) );
  NANDN U47361 ( .A(n38248), .B(n38247), .Z(n38243) );
  IV U47362 ( .A(n38249), .Z(n38247) );
  AND U47363 ( .A(n38250), .B(n38251), .Z(n38216) );
  NAND U47364 ( .A(n38252), .B(n38253), .Z(n38251) );
  NANDN U47365 ( .A(n38254), .B(n38255), .Z(n38253) );
  NANDN U47366 ( .A(n38255), .B(n38254), .Z(n38250) );
  XOR U47367 ( .A(n38226), .B(n38256), .Z(n38218) );
  XNOR U47368 ( .A(n38223), .B(n38225), .Z(n38256) );
  AND U47369 ( .A(n38257), .B(n38258), .Z(n38225) );
  NANDN U47370 ( .A(n38259), .B(n38260), .Z(n38258) );
  OR U47371 ( .A(n38261), .B(n38262), .Z(n38260) );
  IV U47372 ( .A(n38263), .Z(n38262) );
  NANDN U47373 ( .A(n38263), .B(n38261), .Z(n38257) );
  AND U47374 ( .A(n38264), .B(n38265), .Z(n38223) );
  NAND U47375 ( .A(n38266), .B(n38267), .Z(n38265) );
  NANDN U47376 ( .A(n38268), .B(n38269), .Z(n38267) );
  NANDN U47377 ( .A(n38269), .B(n38268), .Z(n38264) );
  IV U47378 ( .A(n38270), .Z(n38269) );
  NAND U47379 ( .A(n38271), .B(n38272), .Z(n38226) );
  NANDN U47380 ( .A(n38273), .B(n38274), .Z(n38272) );
  NANDN U47381 ( .A(n38275), .B(n38276), .Z(n38274) );
  NANDN U47382 ( .A(n38276), .B(n38275), .Z(n38271) );
  IV U47383 ( .A(n38277), .Z(n38275) );
  XOR U47384 ( .A(n38252), .B(n38278), .Z(N61984) );
  XNOR U47385 ( .A(n38255), .B(n38254), .Z(n38278) );
  XNOR U47386 ( .A(n38266), .B(n38279), .Z(n38254) );
  XNOR U47387 ( .A(n38270), .B(n38268), .Z(n38279) );
  XOR U47388 ( .A(n38276), .B(n38280), .Z(n38268) );
  XNOR U47389 ( .A(n38273), .B(n38277), .Z(n38280) );
  AND U47390 ( .A(n38281), .B(n38282), .Z(n38277) );
  NAND U47391 ( .A(n38283), .B(n38284), .Z(n38282) );
  NAND U47392 ( .A(n38285), .B(n38286), .Z(n38281) );
  AND U47393 ( .A(n38287), .B(n38288), .Z(n38273) );
  NAND U47394 ( .A(n38289), .B(n38290), .Z(n38288) );
  NAND U47395 ( .A(n38291), .B(n38292), .Z(n38287) );
  NANDN U47396 ( .A(n38293), .B(n38294), .Z(n38276) );
  ANDN U47397 ( .B(n38295), .A(n38296), .Z(n38270) );
  XNOR U47398 ( .A(n38261), .B(n38297), .Z(n38266) );
  XNOR U47399 ( .A(n38259), .B(n38263), .Z(n38297) );
  AND U47400 ( .A(n38298), .B(n38299), .Z(n38263) );
  NAND U47401 ( .A(n38300), .B(n38301), .Z(n38299) );
  NAND U47402 ( .A(n38302), .B(n38303), .Z(n38298) );
  AND U47403 ( .A(n38304), .B(n38305), .Z(n38259) );
  NAND U47404 ( .A(n38306), .B(n38307), .Z(n38305) );
  NAND U47405 ( .A(n38308), .B(n38309), .Z(n38304) );
  AND U47406 ( .A(n38310), .B(n38311), .Z(n38261) );
  NAND U47407 ( .A(n38312), .B(n38313), .Z(n38255) );
  XNOR U47408 ( .A(n38238), .B(n38314), .Z(n38252) );
  XNOR U47409 ( .A(n38242), .B(n38240), .Z(n38314) );
  XOR U47410 ( .A(n38248), .B(n38315), .Z(n38240) );
  XNOR U47411 ( .A(n38245), .B(n38249), .Z(n38315) );
  AND U47412 ( .A(n38316), .B(n38317), .Z(n38249) );
  NAND U47413 ( .A(n38318), .B(n38319), .Z(n38317) );
  NAND U47414 ( .A(n38320), .B(n38321), .Z(n38316) );
  AND U47415 ( .A(n38322), .B(n38323), .Z(n38245) );
  NAND U47416 ( .A(n38324), .B(n38325), .Z(n38323) );
  NAND U47417 ( .A(n38326), .B(n38327), .Z(n38322) );
  NANDN U47418 ( .A(n38328), .B(n38329), .Z(n38248) );
  ANDN U47419 ( .B(n38330), .A(n38331), .Z(n38242) );
  XNOR U47420 ( .A(n38233), .B(n38332), .Z(n38238) );
  XNOR U47421 ( .A(n38231), .B(n38235), .Z(n38332) );
  AND U47422 ( .A(n38333), .B(n38334), .Z(n38235) );
  NAND U47423 ( .A(n38335), .B(n38336), .Z(n38334) );
  NAND U47424 ( .A(n38337), .B(n38338), .Z(n38333) );
  AND U47425 ( .A(n38339), .B(n38340), .Z(n38231) );
  NAND U47426 ( .A(n38341), .B(n38342), .Z(n38340) );
  NAND U47427 ( .A(n38343), .B(n38344), .Z(n38339) );
  AND U47428 ( .A(n38345), .B(n38346), .Z(n38233) );
  XOR U47429 ( .A(n38313), .B(n38312), .Z(N61983) );
  XNOR U47430 ( .A(n38330), .B(n38331), .Z(n38312) );
  XNOR U47431 ( .A(n38345), .B(n38346), .Z(n38331) );
  XOR U47432 ( .A(n38342), .B(n38341), .Z(n38346) );
  XOR U47433 ( .A(y[2580]), .B(x[2580]), .Z(n38341) );
  XOR U47434 ( .A(n38344), .B(n38343), .Z(n38342) );
  XOR U47435 ( .A(y[2582]), .B(x[2582]), .Z(n38343) );
  XOR U47436 ( .A(y[2581]), .B(x[2581]), .Z(n38344) );
  XOR U47437 ( .A(n38336), .B(n38335), .Z(n38345) );
  XOR U47438 ( .A(n38338), .B(n38337), .Z(n38335) );
  XOR U47439 ( .A(y[2579]), .B(x[2579]), .Z(n38337) );
  XOR U47440 ( .A(y[2578]), .B(x[2578]), .Z(n38338) );
  XOR U47441 ( .A(y[2577]), .B(x[2577]), .Z(n38336) );
  XNOR U47442 ( .A(n38329), .B(n38328), .Z(n38330) );
  XNOR U47443 ( .A(n38325), .B(n38324), .Z(n38328) );
  XOR U47444 ( .A(n38327), .B(n38326), .Z(n38324) );
  XOR U47445 ( .A(y[2576]), .B(x[2576]), .Z(n38326) );
  XOR U47446 ( .A(y[2575]), .B(x[2575]), .Z(n38327) );
  XOR U47447 ( .A(y[2574]), .B(x[2574]), .Z(n38325) );
  XOR U47448 ( .A(n38319), .B(n38318), .Z(n38329) );
  XOR U47449 ( .A(n38321), .B(n38320), .Z(n38318) );
  XOR U47450 ( .A(y[2573]), .B(x[2573]), .Z(n38320) );
  XOR U47451 ( .A(y[2572]), .B(x[2572]), .Z(n38321) );
  XOR U47452 ( .A(y[2571]), .B(x[2571]), .Z(n38319) );
  XNOR U47453 ( .A(n38295), .B(n38296), .Z(n38313) );
  XNOR U47454 ( .A(n38310), .B(n38311), .Z(n38296) );
  XOR U47455 ( .A(n38307), .B(n38306), .Z(n38311) );
  XOR U47456 ( .A(y[2568]), .B(x[2568]), .Z(n38306) );
  XOR U47457 ( .A(n38309), .B(n38308), .Z(n38307) );
  XOR U47458 ( .A(y[2570]), .B(x[2570]), .Z(n38308) );
  XOR U47459 ( .A(y[2569]), .B(x[2569]), .Z(n38309) );
  XOR U47460 ( .A(n38301), .B(n38300), .Z(n38310) );
  XOR U47461 ( .A(n38303), .B(n38302), .Z(n38300) );
  XOR U47462 ( .A(y[2567]), .B(x[2567]), .Z(n38302) );
  XOR U47463 ( .A(y[2566]), .B(x[2566]), .Z(n38303) );
  XOR U47464 ( .A(y[2565]), .B(x[2565]), .Z(n38301) );
  XNOR U47465 ( .A(n38294), .B(n38293), .Z(n38295) );
  XNOR U47466 ( .A(n38290), .B(n38289), .Z(n38293) );
  XOR U47467 ( .A(n38292), .B(n38291), .Z(n38289) );
  XOR U47468 ( .A(y[2564]), .B(x[2564]), .Z(n38291) );
  XOR U47469 ( .A(y[2563]), .B(x[2563]), .Z(n38292) );
  XOR U47470 ( .A(y[2562]), .B(x[2562]), .Z(n38290) );
  XOR U47471 ( .A(n38284), .B(n38283), .Z(n38294) );
  XOR U47472 ( .A(n38286), .B(n38285), .Z(n38283) );
  XOR U47473 ( .A(y[2561]), .B(x[2561]), .Z(n38285) );
  XOR U47474 ( .A(y[2560]), .B(x[2560]), .Z(n38286) );
  XOR U47475 ( .A(y[2559]), .B(x[2559]), .Z(n38284) );
  NAND U47476 ( .A(n38347), .B(n38348), .Z(N61974) );
  NAND U47477 ( .A(n38349), .B(n38350), .Z(n38348) );
  NANDN U47478 ( .A(n38351), .B(n38352), .Z(n38350) );
  NANDN U47479 ( .A(n38352), .B(n38351), .Z(n38347) );
  XOR U47480 ( .A(n38351), .B(n38353), .Z(N61973) );
  XNOR U47481 ( .A(n38349), .B(n38352), .Z(n38353) );
  NAND U47482 ( .A(n38354), .B(n38355), .Z(n38352) );
  NAND U47483 ( .A(n38356), .B(n38357), .Z(n38355) );
  NANDN U47484 ( .A(n38358), .B(n38359), .Z(n38357) );
  NANDN U47485 ( .A(n38359), .B(n38358), .Z(n38354) );
  AND U47486 ( .A(n38360), .B(n38361), .Z(n38349) );
  NAND U47487 ( .A(n38362), .B(n38363), .Z(n38361) );
  NANDN U47488 ( .A(n38364), .B(n38365), .Z(n38363) );
  NANDN U47489 ( .A(n38365), .B(n38364), .Z(n38360) );
  IV U47490 ( .A(n38366), .Z(n38365) );
  AND U47491 ( .A(n38367), .B(n38368), .Z(n38351) );
  NAND U47492 ( .A(n38369), .B(n38370), .Z(n38368) );
  NANDN U47493 ( .A(n38371), .B(n38372), .Z(n38370) );
  NANDN U47494 ( .A(n38372), .B(n38371), .Z(n38367) );
  XOR U47495 ( .A(n38364), .B(n38373), .Z(N61972) );
  XNOR U47496 ( .A(n38362), .B(n38366), .Z(n38373) );
  XOR U47497 ( .A(n38359), .B(n38374), .Z(n38366) );
  XNOR U47498 ( .A(n38356), .B(n38358), .Z(n38374) );
  AND U47499 ( .A(n38375), .B(n38376), .Z(n38358) );
  NANDN U47500 ( .A(n38377), .B(n38378), .Z(n38376) );
  OR U47501 ( .A(n38379), .B(n38380), .Z(n38378) );
  IV U47502 ( .A(n38381), .Z(n38380) );
  NANDN U47503 ( .A(n38381), .B(n38379), .Z(n38375) );
  AND U47504 ( .A(n38382), .B(n38383), .Z(n38356) );
  NAND U47505 ( .A(n38384), .B(n38385), .Z(n38383) );
  NANDN U47506 ( .A(n38386), .B(n38387), .Z(n38385) );
  NANDN U47507 ( .A(n38387), .B(n38386), .Z(n38382) );
  IV U47508 ( .A(n38388), .Z(n38387) );
  NAND U47509 ( .A(n38389), .B(n38390), .Z(n38359) );
  NANDN U47510 ( .A(n38391), .B(n38392), .Z(n38390) );
  NANDN U47511 ( .A(n38393), .B(n38394), .Z(n38392) );
  NANDN U47512 ( .A(n38394), .B(n38393), .Z(n38389) );
  IV U47513 ( .A(n38395), .Z(n38393) );
  AND U47514 ( .A(n38396), .B(n38397), .Z(n38362) );
  NAND U47515 ( .A(n38398), .B(n38399), .Z(n38397) );
  NANDN U47516 ( .A(n38400), .B(n38401), .Z(n38399) );
  NANDN U47517 ( .A(n38401), .B(n38400), .Z(n38396) );
  XOR U47518 ( .A(n38372), .B(n38402), .Z(n38364) );
  XNOR U47519 ( .A(n38369), .B(n38371), .Z(n38402) );
  AND U47520 ( .A(n38403), .B(n38404), .Z(n38371) );
  NANDN U47521 ( .A(n38405), .B(n38406), .Z(n38404) );
  OR U47522 ( .A(n38407), .B(n38408), .Z(n38406) );
  IV U47523 ( .A(n38409), .Z(n38408) );
  NANDN U47524 ( .A(n38409), .B(n38407), .Z(n38403) );
  AND U47525 ( .A(n38410), .B(n38411), .Z(n38369) );
  NAND U47526 ( .A(n38412), .B(n38413), .Z(n38411) );
  NANDN U47527 ( .A(n38414), .B(n38415), .Z(n38413) );
  NANDN U47528 ( .A(n38415), .B(n38414), .Z(n38410) );
  IV U47529 ( .A(n38416), .Z(n38415) );
  NAND U47530 ( .A(n38417), .B(n38418), .Z(n38372) );
  NANDN U47531 ( .A(n38419), .B(n38420), .Z(n38418) );
  NANDN U47532 ( .A(n38421), .B(n38422), .Z(n38420) );
  NANDN U47533 ( .A(n38422), .B(n38421), .Z(n38417) );
  IV U47534 ( .A(n38423), .Z(n38421) );
  XOR U47535 ( .A(n38398), .B(n38424), .Z(N61971) );
  XNOR U47536 ( .A(n38401), .B(n38400), .Z(n38424) );
  XNOR U47537 ( .A(n38412), .B(n38425), .Z(n38400) );
  XNOR U47538 ( .A(n38416), .B(n38414), .Z(n38425) );
  XOR U47539 ( .A(n38422), .B(n38426), .Z(n38414) );
  XNOR U47540 ( .A(n38419), .B(n38423), .Z(n38426) );
  AND U47541 ( .A(n38427), .B(n38428), .Z(n38423) );
  NAND U47542 ( .A(n38429), .B(n38430), .Z(n38428) );
  NAND U47543 ( .A(n38431), .B(n38432), .Z(n38427) );
  AND U47544 ( .A(n38433), .B(n38434), .Z(n38419) );
  NAND U47545 ( .A(n38435), .B(n38436), .Z(n38434) );
  NAND U47546 ( .A(n38437), .B(n38438), .Z(n38433) );
  NANDN U47547 ( .A(n38439), .B(n38440), .Z(n38422) );
  ANDN U47548 ( .B(n38441), .A(n38442), .Z(n38416) );
  XNOR U47549 ( .A(n38407), .B(n38443), .Z(n38412) );
  XNOR U47550 ( .A(n38405), .B(n38409), .Z(n38443) );
  AND U47551 ( .A(n38444), .B(n38445), .Z(n38409) );
  NAND U47552 ( .A(n38446), .B(n38447), .Z(n38445) );
  NAND U47553 ( .A(n38448), .B(n38449), .Z(n38444) );
  AND U47554 ( .A(n38450), .B(n38451), .Z(n38405) );
  NAND U47555 ( .A(n38452), .B(n38453), .Z(n38451) );
  NAND U47556 ( .A(n38454), .B(n38455), .Z(n38450) );
  AND U47557 ( .A(n38456), .B(n38457), .Z(n38407) );
  NAND U47558 ( .A(n38458), .B(n38459), .Z(n38401) );
  XNOR U47559 ( .A(n38384), .B(n38460), .Z(n38398) );
  XNOR U47560 ( .A(n38388), .B(n38386), .Z(n38460) );
  XOR U47561 ( .A(n38394), .B(n38461), .Z(n38386) );
  XNOR U47562 ( .A(n38391), .B(n38395), .Z(n38461) );
  AND U47563 ( .A(n38462), .B(n38463), .Z(n38395) );
  NAND U47564 ( .A(n38464), .B(n38465), .Z(n38463) );
  NAND U47565 ( .A(n38466), .B(n38467), .Z(n38462) );
  AND U47566 ( .A(n38468), .B(n38469), .Z(n38391) );
  NAND U47567 ( .A(n38470), .B(n38471), .Z(n38469) );
  NAND U47568 ( .A(n38472), .B(n38473), .Z(n38468) );
  NANDN U47569 ( .A(n38474), .B(n38475), .Z(n38394) );
  ANDN U47570 ( .B(n38476), .A(n38477), .Z(n38388) );
  XNOR U47571 ( .A(n38379), .B(n38478), .Z(n38384) );
  XNOR U47572 ( .A(n38377), .B(n38381), .Z(n38478) );
  AND U47573 ( .A(n38479), .B(n38480), .Z(n38381) );
  NAND U47574 ( .A(n38481), .B(n38482), .Z(n38480) );
  NAND U47575 ( .A(n38483), .B(n38484), .Z(n38479) );
  AND U47576 ( .A(n38485), .B(n38486), .Z(n38377) );
  NAND U47577 ( .A(n38487), .B(n38488), .Z(n38486) );
  NAND U47578 ( .A(n38489), .B(n38490), .Z(n38485) );
  AND U47579 ( .A(n38491), .B(n38492), .Z(n38379) );
  XOR U47580 ( .A(n38459), .B(n38458), .Z(N61970) );
  XNOR U47581 ( .A(n38476), .B(n38477), .Z(n38458) );
  XNOR U47582 ( .A(n38491), .B(n38492), .Z(n38477) );
  XOR U47583 ( .A(n38488), .B(n38487), .Z(n38492) );
  XOR U47584 ( .A(y[2556]), .B(x[2556]), .Z(n38487) );
  XOR U47585 ( .A(n38490), .B(n38489), .Z(n38488) );
  XOR U47586 ( .A(y[2558]), .B(x[2558]), .Z(n38489) );
  XOR U47587 ( .A(y[2557]), .B(x[2557]), .Z(n38490) );
  XOR U47588 ( .A(n38482), .B(n38481), .Z(n38491) );
  XOR U47589 ( .A(n38484), .B(n38483), .Z(n38481) );
  XOR U47590 ( .A(y[2555]), .B(x[2555]), .Z(n38483) );
  XOR U47591 ( .A(y[2554]), .B(x[2554]), .Z(n38484) );
  XOR U47592 ( .A(y[2553]), .B(x[2553]), .Z(n38482) );
  XNOR U47593 ( .A(n38475), .B(n38474), .Z(n38476) );
  XNOR U47594 ( .A(n38471), .B(n38470), .Z(n38474) );
  XOR U47595 ( .A(n38473), .B(n38472), .Z(n38470) );
  XOR U47596 ( .A(y[2552]), .B(x[2552]), .Z(n38472) );
  XOR U47597 ( .A(y[2551]), .B(x[2551]), .Z(n38473) );
  XOR U47598 ( .A(y[2550]), .B(x[2550]), .Z(n38471) );
  XOR U47599 ( .A(n38465), .B(n38464), .Z(n38475) );
  XOR U47600 ( .A(n38467), .B(n38466), .Z(n38464) );
  XOR U47601 ( .A(y[2549]), .B(x[2549]), .Z(n38466) );
  XOR U47602 ( .A(y[2548]), .B(x[2548]), .Z(n38467) );
  XOR U47603 ( .A(y[2547]), .B(x[2547]), .Z(n38465) );
  XNOR U47604 ( .A(n38441), .B(n38442), .Z(n38459) );
  XNOR U47605 ( .A(n38456), .B(n38457), .Z(n38442) );
  XOR U47606 ( .A(n38453), .B(n38452), .Z(n38457) );
  XOR U47607 ( .A(y[2544]), .B(x[2544]), .Z(n38452) );
  XOR U47608 ( .A(n38455), .B(n38454), .Z(n38453) );
  XOR U47609 ( .A(y[2546]), .B(x[2546]), .Z(n38454) );
  XOR U47610 ( .A(y[2545]), .B(x[2545]), .Z(n38455) );
  XOR U47611 ( .A(n38447), .B(n38446), .Z(n38456) );
  XOR U47612 ( .A(n38449), .B(n38448), .Z(n38446) );
  XOR U47613 ( .A(y[2543]), .B(x[2543]), .Z(n38448) );
  XOR U47614 ( .A(y[2542]), .B(x[2542]), .Z(n38449) );
  XOR U47615 ( .A(y[2541]), .B(x[2541]), .Z(n38447) );
  XNOR U47616 ( .A(n38440), .B(n38439), .Z(n38441) );
  XNOR U47617 ( .A(n38436), .B(n38435), .Z(n38439) );
  XOR U47618 ( .A(n38438), .B(n38437), .Z(n38435) );
  XOR U47619 ( .A(y[2540]), .B(x[2540]), .Z(n38437) );
  XOR U47620 ( .A(y[2539]), .B(x[2539]), .Z(n38438) );
  XOR U47621 ( .A(y[2538]), .B(x[2538]), .Z(n38436) );
  XOR U47622 ( .A(n38430), .B(n38429), .Z(n38440) );
  XOR U47623 ( .A(n38432), .B(n38431), .Z(n38429) );
  XOR U47624 ( .A(y[2537]), .B(x[2537]), .Z(n38431) );
  XOR U47625 ( .A(y[2536]), .B(x[2536]), .Z(n38432) );
  XOR U47626 ( .A(y[2535]), .B(x[2535]), .Z(n38430) );
  NAND U47627 ( .A(n38493), .B(n38494), .Z(N61961) );
  NAND U47628 ( .A(n38495), .B(n38496), .Z(n38494) );
  NANDN U47629 ( .A(n38497), .B(n38498), .Z(n38496) );
  NANDN U47630 ( .A(n38498), .B(n38497), .Z(n38493) );
  XOR U47631 ( .A(n38497), .B(n38499), .Z(N61960) );
  XNOR U47632 ( .A(n38495), .B(n38498), .Z(n38499) );
  NAND U47633 ( .A(n38500), .B(n38501), .Z(n38498) );
  NAND U47634 ( .A(n38502), .B(n38503), .Z(n38501) );
  NANDN U47635 ( .A(n38504), .B(n38505), .Z(n38503) );
  NANDN U47636 ( .A(n38505), .B(n38504), .Z(n38500) );
  AND U47637 ( .A(n38506), .B(n38507), .Z(n38495) );
  NAND U47638 ( .A(n38508), .B(n38509), .Z(n38507) );
  NANDN U47639 ( .A(n38510), .B(n38511), .Z(n38509) );
  NANDN U47640 ( .A(n38511), .B(n38510), .Z(n38506) );
  IV U47641 ( .A(n38512), .Z(n38511) );
  AND U47642 ( .A(n38513), .B(n38514), .Z(n38497) );
  NAND U47643 ( .A(n38515), .B(n38516), .Z(n38514) );
  NANDN U47644 ( .A(n38517), .B(n38518), .Z(n38516) );
  NANDN U47645 ( .A(n38518), .B(n38517), .Z(n38513) );
  XOR U47646 ( .A(n38510), .B(n38519), .Z(N61959) );
  XNOR U47647 ( .A(n38508), .B(n38512), .Z(n38519) );
  XOR U47648 ( .A(n38505), .B(n38520), .Z(n38512) );
  XNOR U47649 ( .A(n38502), .B(n38504), .Z(n38520) );
  AND U47650 ( .A(n38521), .B(n38522), .Z(n38504) );
  NANDN U47651 ( .A(n38523), .B(n38524), .Z(n38522) );
  OR U47652 ( .A(n38525), .B(n38526), .Z(n38524) );
  IV U47653 ( .A(n38527), .Z(n38526) );
  NANDN U47654 ( .A(n38527), .B(n38525), .Z(n38521) );
  AND U47655 ( .A(n38528), .B(n38529), .Z(n38502) );
  NAND U47656 ( .A(n38530), .B(n38531), .Z(n38529) );
  NANDN U47657 ( .A(n38532), .B(n38533), .Z(n38531) );
  NANDN U47658 ( .A(n38533), .B(n38532), .Z(n38528) );
  IV U47659 ( .A(n38534), .Z(n38533) );
  NAND U47660 ( .A(n38535), .B(n38536), .Z(n38505) );
  NANDN U47661 ( .A(n38537), .B(n38538), .Z(n38536) );
  NANDN U47662 ( .A(n38539), .B(n38540), .Z(n38538) );
  NANDN U47663 ( .A(n38540), .B(n38539), .Z(n38535) );
  IV U47664 ( .A(n38541), .Z(n38539) );
  AND U47665 ( .A(n38542), .B(n38543), .Z(n38508) );
  NAND U47666 ( .A(n38544), .B(n38545), .Z(n38543) );
  NANDN U47667 ( .A(n38546), .B(n38547), .Z(n38545) );
  NANDN U47668 ( .A(n38547), .B(n38546), .Z(n38542) );
  XOR U47669 ( .A(n38518), .B(n38548), .Z(n38510) );
  XNOR U47670 ( .A(n38515), .B(n38517), .Z(n38548) );
  AND U47671 ( .A(n38549), .B(n38550), .Z(n38517) );
  NANDN U47672 ( .A(n38551), .B(n38552), .Z(n38550) );
  OR U47673 ( .A(n38553), .B(n38554), .Z(n38552) );
  IV U47674 ( .A(n38555), .Z(n38554) );
  NANDN U47675 ( .A(n38555), .B(n38553), .Z(n38549) );
  AND U47676 ( .A(n38556), .B(n38557), .Z(n38515) );
  NAND U47677 ( .A(n38558), .B(n38559), .Z(n38557) );
  NANDN U47678 ( .A(n38560), .B(n38561), .Z(n38559) );
  NANDN U47679 ( .A(n38561), .B(n38560), .Z(n38556) );
  IV U47680 ( .A(n38562), .Z(n38561) );
  NAND U47681 ( .A(n38563), .B(n38564), .Z(n38518) );
  NANDN U47682 ( .A(n38565), .B(n38566), .Z(n38564) );
  NANDN U47683 ( .A(n38567), .B(n38568), .Z(n38566) );
  NANDN U47684 ( .A(n38568), .B(n38567), .Z(n38563) );
  IV U47685 ( .A(n38569), .Z(n38567) );
  XOR U47686 ( .A(n38544), .B(n38570), .Z(N61958) );
  XNOR U47687 ( .A(n38547), .B(n38546), .Z(n38570) );
  XNOR U47688 ( .A(n38558), .B(n38571), .Z(n38546) );
  XNOR U47689 ( .A(n38562), .B(n38560), .Z(n38571) );
  XOR U47690 ( .A(n38568), .B(n38572), .Z(n38560) );
  XNOR U47691 ( .A(n38565), .B(n38569), .Z(n38572) );
  AND U47692 ( .A(n38573), .B(n38574), .Z(n38569) );
  NAND U47693 ( .A(n38575), .B(n38576), .Z(n38574) );
  NAND U47694 ( .A(n38577), .B(n38578), .Z(n38573) );
  AND U47695 ( .A(n38579), .B(n38580), .Z(n38565) );
  NAND U47696 ( .A(n38581), .B(n38582), .Z(n38580) );
  NAND U47697 ( .A(n38583), .B(n38584), .Z(n38579) );
  NANDN U47698 ( .A(n38585), .B(n38586), .Z(n38568) );
  ANDN U47699 ( .B(n38587), .A(n38588), .Z(n38562) );
  XNOR U47700 ( .A(n38553), .B(n38589), .Z(n38558) );
  XNOR U47701 ( .A(n38551), .B(n38555), .Z(n38589) );
  AND U47702 ( .A(n38590), .B(n38591), .Z(n38555) );
  NAND U47703 ( .A(n38592), .B(n38593), .Z(n38591) );
  NAND U47704 ( .A(n38594), .B(n38595), .Z(n38590) );
  AND U47705 ( .A(n38596), .B(n38597), .Z(n38551) );
  NAND U47706 ( .A(n38598), .B(n38599), .Z(n38597) );
  NAND U47707 ( .A(n38600), .B(n38601), .Z(n38596) );
  AND U47708 ( .A(n38602), .B(n38603), .Z(n38553) );
  NAND U47709 ( .A(n38604), .B(n38605), .Z(n38547) );
  XNOR U47710 ( .A(n38530), .B(n38606), .Z(n38544) );
  XNOR U47711 ( .A(n38534), .B(n38532), .Z(n38606) );
  XOR U47712 ( .A(n38540), .B(n38607), .Z(n38532) );
  XNOR U47713 ( .A(n38537), .B(n38541), .Z(n38607) );
  AND U47714 ( .A(n38608), .B(n38609), .Z(n38541) );
  NAND U47715 ( .A(n38610), .B(n38611), .Z(n38609) );
  NAND U47716 ( .A(n38612), .B(n38613), .Z(n38608) );
  AND U47717 ( .A(n38614), .B(n38615), .Z(n38537) );
  NAND U47718 ( .A(n38616), .B(n38617), .Z(n38615) );
  NAND U47719 ( .A(n38618), .B(n38619), .Z(n38614) );
  NANDN U47720 ( .A(n38620), .B(n38621), .Z(n38540) );
  ANDN U47721 ( .B(n38622), .A(n38623), .Z(n38534) );
  XNOR U47722 ( .A(n38525), .B(n38624), .Z(n38530) );
  XNOR U47723 ( .A(n38523), .B(n38527), .Z(n38624) );
  AND U47724 ( .A(n38625), .B(n38626), .Z(n38527) );
  NAND U47725 ( .A(n38627), .B(n38628), .Z(n38626) );
  NAND U47726 ( .A(n38629), .B(n38630), .Z(n38625) );
  AND U47727 ( .A(n38631), .B(n38632), .Z(n38523) );
  NAND U47728 ( .A(n38633), .B(n38634), .Z(n38632) );
  NAND U47729 ( .A(n38635), .B(n38636), .Z(n38631) );
  AND U47730 ( .A(n38637), .B(n38638), .Z(n38525) );
  XOR U47731 ( .A(n38605), .B(n38604), .Z(N61957) );
  XNOR U47732 ( .A(n38622), .B(n38623), .Z(n38604) );
  XNOR U47733 ( .A(n38637), .B(n38638), .Z(n38623) );
  XOR U47734 ( .A(n38634), .B(n38633), .Z(n38638) );
  XOR U47735 ( .A(y[2532]), .B(x[2532]), .Z(n38633) );
  XOR U47736 ( .A(n38636), .B(n38635), .Z(n38634) );
  XOR U47737 ( .A(y[2534]), .B(x[2534]), .Z(n38635) );
  XOR U47738 ( .A(y[2533]), .B(x[2533]), .Z(n38636) );
  XOR U47739 ( .A(n38628), .B(n38627), .Z(n38637) );
  XOR U47740 ( .A(n38630), .B(n38629), .Z(n38627) );
  XOR U47741 ( .A(y[2531]), .B(x[2531]), .Z(n38629) );
  XOR U47742 ( .A(y[2530]), .B(x[2530]), .Z(n38630) );
  XOR U47743 ( .A(y[2529]), .B(x[2529]), .Z(n38628) );
  XNOR U47744 ( .A(n38621), .B(n38620), .Z(n38622) );
  XNOR U47745 ( .A(n38617), .B(n38616), .Z(n38620) );
  XOR U47746 ( .A(n38619), .B(n38618), .Z(n38616) );
  XOR U47747 ( .A(y[2528]), .B(x[2528]), .Z(n38618) );
  XOR U47748 ( .A(y[2527]), .B(x[2527]), .Z(n38619) );
  XOR U47749 ( .A(y[2526]), .B(x[2526]), .Z(n38617) );
  XOR U47750 ( .A(n38611), .B(n38610), .Z(n38621) );
  XOR U47751 ( .A(n38613), .B(n38612), .Z(n38610) );
  XOR U47752 ( .A(y[2525]), .B(x[2525]), .Z(n38612) );
  XOR U47753 ( .A(y[2524]), .B(x[2524]), .Z(n38613) );
  XOR U47754 ( .A(y[2523]), .B(x[2523]), .Z(n38611) );
  XNOR U47755 ( .A(n38587), .B(n38588), .Z(n38605) );
  XNOR U47756 ( .A(n38602), .B(n38603), .Z(n38588) );
  XOR U47757 ( .A(n38599), .B(n38598), .Z(n38603) );
  XOR U47758 ( .A(y[2520]), .B(x[2520]), .Z(n38598) );
  XOR U47759 ( .A(n38601), .B(n38600), .Z(n38599) );
  XOR U47760 ( .A(y[2522]), .B(x[2522]), .Z(n38600) );
  XOR U47761 ( .A(y[2521]), .B(x[2521]), .Z(n38601) );
  XOR U47762 ( .A(n38593), .B(n38592), .Z(n38602) );
  XOR U47763 ( .A(n38595), .B(n38594), .Z(n38592) );
  XOR U47764 ( .A(y[2519]), .B(x[2519]), .Z(n38594) );
  XOR U47765 ( .A(y[2518]), .B(x[2518]), .Z(n38595) );
  XOR U47766 ( .A(y[2517]), .B(x[2517]), .Z(n38593) );
  XNOR U47767 ( .A(n38586), .B(n38585), .Z(n38587) );
  XNOR U47768 ( .A(n38582), .B(n38581), .Z(n38585) );
  XOR U47769 ( .A(n38584), .B(n38583), .Z(n38581) );
  XOR U47770 ( .A(y[2516]), .B(x[2516]), .Z(n38583) );
  XOR U47771 ( .A(y[2515]), .B(x[2515]), .Z(n38584) );
  XOR U47772 ( .A(y[2514]), .B(x[2514]), .Z(n38582) );
  XOR U47773 ( .A(n38576), .B(n38575), .Z(n38586) );
  XOR U47774 ( .A(n38578), .B(n38577), .Z(n38575) );
  XOR U47775 ( .A(y[2513]), .B(x[2513]), .Z(n38577) );
  XOR U47776 ( .A(y[2512]), .B(x[2512]), .Z(n38578) );
  XOR U47777 ( .A(y[2511]), .B(x[2511]), .Z(n38576) );
  NAND U47778 ( .A(n38639), .B(n38640), .Z(N61948) );
  NAND U47779 ( .A(n38641), .B(n38642), .Z(n38640) );
  NANDN U47780 ( .A(n38643), .B(n38644), .Z(n38642) );
  NANDN U47781 ( .A(n38644), .B(n38643), .Z(n38639) );
  XOR U47782 ( .A(n38643), .B(n38645), .Z(N61947) );
  XNOR U47783 ( .A(n38641), .B(n38644), .Z(n38645) );
  NAND U47784 ( .A(n38646), .B(n38647), .Z(n38644) );
  NAND U47785 ( .A(n38648), .B(n38649), .Z(n38647) );
  NANDN U47786 ( .A(n38650), .B(n38651), .Z(n38649) );
  NANDN U47787 ( .A(n38651), .B(n38650), .Z(n38646) );
  AND U47788 ( .A(n38652), .B(n38653), .Z(n38641) );
  NAND U47789 ( .A(n38654), .B(n38655), .Z(n38653) );
  NANDN U47790 ( .A(n38656), .B(n38657), .Z(n38655) );
  NANDN U47791 ( .A(n38657), .B(n38656), .Z(n38652) );
  IV U47792 ( .A(n38658), .Z(n38657) );
  AND U47793 ( .A(n38659), .B(n38660), .Z(n38643) );
  NAND U47794 ( .A(n38661), .B(n38662), .Z(n38660) );
  NANDN U47795 ( .A(n38663), .B(n38664), .Z(n38662) );
  NANDN U47796 ( .A(n38664), .B(n38663), .Z(n38659) );
  XOR U47797 ( .A(n38656), .B(n38665), .Z(N61946) );
  XNOR U47798 ( .A(n38654), .B(n38658), .Z(n38665) );
  XOR U47799 ( .A(n38651), .B(n38666), .Z(n38658) );
  XNOR U47800 ( .A(n38648), .B(n38650), .Z(n38666) );
  AND U47801 ( .A(n38667), .B(n38668), .Z(n38650) );
  NANDN U47802 ( .A(n38669), .B(n38670), .Z(n38668) );
  OR U47803 ( .A(n38671), .B(n38672), .Z(n38670) );
  IV U47804 ( .A(n38673), .Z(n38672) );
  NANDN U47805 ( .A(n38673), .B(n38671), .Z(n38667) );
  AND U47806 ( .A(n38674), .B(n38675), .Z(n38648) );
  NAND U47807 ( .A(n38676), .B(n38677), .Z(n38675) );
  NANDN U47808 ( .A(n38678), .B(n38679), .Z(n38677) );
  NANDN U47809 ( .A(n38679), .B(n38678), .Z(n38674) );
  IV U47810 ( .A(n38680), .Z(n38679) );
  NAND U47811 ( .A(n38681), .B(n38682), .Z(n38651) );
  NANDN U47812 ( .A(n38683), .B(n38684), .Z(n38682) );
  NANDN U47813 ( .A(n38685), .B(n38686), .Z(n38684) );
  NANDN U47814 ( .A(n38686), .B(n38685), .Z(n38681) );
  IV U47815 ( .A(n38687), .Z(n38685) );
  AND U47816 ( .A(n38688), .B(n38689), .Z(n38654) );
  NAND U47817 ( .A(n38690), .B(n38691), .Z(n38689) );
  NANDN U47818 ( .A(n38692), .B(n38693), .Z(n38691) );
  NANDN U47819 ( .A(n38693), .B(n38692), .Z(n38688) );
  XOR U47820 ( .A(n38664), .B(n38694), .Z(n38656) );
  XNOR U47821 ( .A(n38661), .B(n38663), .Z(n38694) );
  AND U47822 ( .A(n38695), .B(n38696), .Z(n38663) );
  NANDN U47823 ( .A(n38697), .B(n38698), .Z(n38696) );
  OR U47824 ( .A(n38699), .B(n38700), .Z(n38698) );
  IV U47825 ( .A(n38701), .Z(n38700) );
  NANDN U47826 ( .A(n38701), .B(n38699), .Z(n38695) );
  AND U47827 ( .A(n38702), .B(n38703), .Z(n38661) );
  NAND U47828 ( .A(n38704), .B(n38705), .Z(n38703) );
  NANDN U47829 ( .A(n38706), .B(n38707), .Z(n38705) );
  NANDN U47830 ( .A(n38707), .B(n38706), .Z(n38702) );
  IV U47831 ( .A(n38708), .Z(n38707) );
  NAND U47832 ( .A(n38709), .B(n38710), .Z(n38664) );
  NANDN U47833 ( .A(n38711), .B(n38712), .Z(n38710) );
  NANDN U47834 ( .A(n38713), .B(n38714), .Z(n38712) );
  NANDN U47835 ( .A(n38714), .B(n38713), .Z(n38709) );
  IV U47836 ( .A(n38715), .Z(n38713) );
  XOR U47837 ( .A(n38690), .B(n38716), .Z(N61945) );
  XNOR U47838 ( .A(n38693), .B(n38692), .Z(n38716) );
  XNOR U47839 ( .A(n38704), .B(n38717), .Z(n38692) );
  XNOR U47840 ( .A(n38708), .B(n38706), .Z(n38717) );
  XOR U47841 ( .A(n38714), .B(n38718), .Z(n38706) );
  XNOR U47842 ( .A(n38711), .B(n38715), .Z(n38718) );
  AND U47843 ( .A(n38719), .B(n38720), .Z(n38715) );
  NAND U47844 ( .A(n38721), .B(n38722), .Z(n38720) );
  NAND U47845 ( .A(n38723), .B(n38724), .Z(n38719) );
  AND U47846 ( .A(n38725), .B(n38726), .Z(n38711) );
  NAND U47847 ( .A(n38727), .B(n38728), .Z(n38726) );
  NAND U47848 ( .A(n38729), .B(n38730), .Z(n38725) );
  NANDN U47849 ( .A(n38731), .B(n38732), .Z(n38714) );
  ANDN U47850 ( .B(n38733), .A(n38734), .Z(n38708) );
  XNOR U47851 ( .A(n38699), .B(n38735), .Z(n38704) );
  XNOR U47852 ( .A(n38697), .B(n38701), .Z(n38735) );
  AND U47853 ( .A(n38736), .B(n38737), .Z(n38701) );
  NAND U47854 ( .A(n38738), .B(n38739), .Z(n38737) );
  NAND U47855 ( .A(n38740), .B(n38741), .Z(n38736) );
  AND U47856 ( .A(n38742), .B(n38743), .Z(n38697) );
  NAND U47857 ( .A(n38744), .B(n38745), .Z(n38743) );
  NAND U47858 ( .A(n38746), .B(n38747), .Z(n38742) );
  AND U47859 ( .A(n38748), .B(n38749), .Z(n38699) );
  NAND U47860 ( .A(n38750), .B(n38751), .Z(n38693) );
  XNOR U47861 ( .A(n38676), .B(n38752), .Z(n38690) );
  XNOR U47862 ( .A(n38680), .B(n38678), .Z(n38752) );
  XOR U47863 ( .A(n38686), .B(n38753), .Z(n38678) );
  XNOR U47864 ( .A(n38683), .B(n38687), .Z(n38753) );
  AND U47865 ( .A(n38754), .B(n38755), .Z(n38687) );
  NAND U47866 ( .A(n38756), .B(n38757), .Z(n38755) );
  NAND U47867 ( .A(n38758), .B(n38759), .Z(n38754) );
  AND U47868 ( .A(n38760), .B(n38761), .Z(n38683) );
  NAND U47869 ( .A(n38762), .B(n38763), .Z(n38761) );
  NAND U47870 ( .A(n38764), .B(n38765), .Z(n38760) );
  NANDN U47871 ( .A(n38766), .B(n38767), .Z(n38686) );
  ANDN U47872 ( .B(n38768), .A(n38769), .Z(n38680) );
  XNOR U47873 ( .A(n38671), .B(n38770), .Z(n38676) );
  XNOR U47874 ( .A(n38669), .B(n38673), .Z(n38770) );
  AND U47875 ( .A(n38771), .B(n38772), .Z(n38673) );
  NAND U47876 ( .A(n38773), .B(n38774), .Z(n38772) );
  NAND U47877 ( .A(n38775), .B(n38776), .Z(n38771) );
  AND U47878 ( .A(n38777), .B(n38778), .Z(n38669) );
  NAND U47879 ( .A(n38779), .B(n38780), .Z(n38778) );
  NAND U47880 ( .A(n38781), .B(n38782), .Z(n38777) );
  AND U47881 ( .A(n38783), .B(n38784), .Z(n38671) );
  XOR U47882 ( .A(n38751), .B(n38750), .Z(N61944) );
  XNOR U47883 ( .A(n38768), .B(n38769), .Z(n38750) );
  XNOR U47884 ( .A(n38783), .B(n38784), .Z(n38769) );
  XOR U47885 ( .A(n38780), .B(n38779), .Z(n38784) );
  XOR U47886 ( .A(y[2508]), .B(x[2508]), .Z(n38779) );
  XOR U47887 ( .A(n38782), .B(n38781), .Z(n38780) );
  XOR U47888 ( .A(y[2510]), .B(x[2510]), .Z(n38781) );
  XOR U47889 ( .A(y[2509]), .B(x[2509]), .Z(n38782) );
  XOR U47890 ( .A(n38774), .B(n38773), .Z(n38783) );
  XOR U47891 ( .A(n38776), .B(n38775), .Z(n38773) );
  XOR U47892 ( .A(y[2507]), .B(x[2507]), .Z(n38775) );
  XOR U47893 ( .A(y[2506]), .B(x[2506]), .Z(n38776) );
  XOR U47894 ( .A(y[2505]), .B(x[2505]), .Z(n38774) );
  XNOR U47895 ( .A(n38767), .B(n38766), .Z(n38768) );
  XNOR U47896 ( .A(n38763), .B(n38762), .Z(n38766) );
  XOR U47897 ( .A(n38765), .B(n38764), .Z(n38762) );
  XOR U47898 ( .A(y[2504]), .B(x[2504]), .Z(n38764) );
  XOR U47899 ( .A(y[2503]), .B(x[2503]), .Z(n38765) );
  XOR U47900 ( .A(y[2502]), .B(x[2502]), .Z(n38763) );
  XOR U47901 ( .A(n38757), .B(n38756), .Z(n38767) );
  XOR U47902 ( .A(n38759), .B(n38758), .Z(n38756) );
  XOR U47903 ( .A(y[2501]), .B(x[2501]), .Z(n38758) );
  XOR U47904 ( .A(y[2500]), .B(x[2500]), .Z(n38759) );
  XOR U47905 ( .A(y[2499]), .B(x[2499]), .Z(n38757) );
  XNOR U47906 ( .A(n38733), .B(n38734), .Z(n38751) );
  XNOR U47907 ( .A(n38748), .B(n38749), .Z(n38734) );
  XOR U47908 ( .A(n38745), .B(n38744), .Z(n38749) );
  XOR U47909 ( .A(y[2496]), .B(x[2496]), .Z(n38744) );
  XOR U47910 ( .A(n38747), .B(n38746), .Z(n38745) );
  XOR U47911 ( .A(y[2498]), .B(x[2498]), .Z(n38746) );
  XOR U47912 ( .A(y[2497]), .B(x[2497]), .Z(n38747) );
  XOR U47913 ( .A(n38739), .B(n38738), .Z(n38748) );
  XOR U47914 ( .A(n38741), .B(n38740), .Z(n38738) );
  XOR U47915 ( .A(y[2495]), .B(x[2495]), .Z(n38740) );
  XOR U47916 ( .A(y[2494]), .B(x[2494]), .Z(n38741) );
  XOR U47917 ( .A(y[2493]), .B(x[2493]), .Z(n38739) );
  XNOR U47918 ( .A(n38732), .B(n38731), .Z(n38733) );
  XNOR U47919 ( .A(n38728), .B(n38727), .Z(n38731) );
  XOR U47920 ( .A(n38730), .B(n38729), .Z(n38727) );
  XOR U47921 ( .A(y[2492]), .B(x[2492]), .Z(n38729) );
  XOR U47922 ( .A(y[2491]), .B(x[2491]), .Z(n38730) );
  XOR U47923 ( .A(y[2490]), .B(x[2490]), .Z(n38728) );
  XOR U47924 ( .A(n38722), .B(n38721), .Z(n38732) );
  XOR U47925 ( .A(n38724), .B(n38723), .Z(n38721) );
  XOR U47926 ( .A(y[2489]), .B(x[2489]), .Z(n38723) );
  XOR U47927 ( .A(y[2488]), .B(x[2488]), .Z(n38724) );
  XOR U47928 ( .A(y[2487]), .B(x[2487]), .Z(n38722) );
  NAND U47929 ( .A(n38785), .B(n38786), .Z(N61935) );
  NAND U47930 ( .A(n38787), .B(n38788), .Z(n38786) );
  NANDN U47931 ( .A(n38789), .B(n38790), .Z(n38788) );
  NANDN U47932 ( .A(n38790), .B(n38789), .Z(n38785) );
  XOR U47933 ( .A(n38789), .B(n38791), .Z(N61934) );
  XNOR U47934 ( .A(n38787), .B(n38790), .Z(n38791) );
  NAND U47935 ( .A(n38792), .B(n38793), .Z(n38790) );
  NAND U47936 ( .A(n38794), .B(n38795), .Z(n38793) );
  NANDN U47937 ( .A(n38796), .B(n38797), .Z(n38795) );
  NANDN U47938 ( .A(n38797), .B(n38796), .Z(n38792) );
  AND U47939 ( .A(n38798), .B(n38799), .Z(n38787) );
  NAND U47940 ( .A(n38800), .B(n38801), .Z(n38799) );
  NANDN U47941 ( .A(n38802), .B(n38803), .Z(n38801) );
  NANDN U47942 ( .A(n38803), .B(n38802), .Z(n38798) );
  IV U47943 ( .A(n38804), .Z(n38803) );
  AND U47944 ( .A(n38805), .B(n38806), .Z(n38789) );
  NAND U47945 ( .A(n38807), .B(n38808), .Z(n38806) );
  NANDN U47946 ( .A(n38809), .B(n38810), .Z(n38808) );
  NANDN U47947 ( .A(n38810), .B(n38809), .Z(n38805) );
  XOR U47948 ( .A(n38802), .B(n38811), .Z(N61933) );
  XNOR U47949 ( .A(n38800), .B(n38804), .Z(n38811) );
  XOR U47950 ( .A(n38797), .B(n38812), .Z(n38804) );
  XNOR U47951 ( .A(n38794), .B(n38796), .Z(n38812) );
  AND U47952 ( .A(n38813), .B(n38814), .Z(n38796) );
  NANDN U47953 ( .A(n38815), .B(n38816), .Z(n38814) );
  OR U47954 ( .A(n38817), .B(n38818), .Z(n38816) );
  IV U47955 ( .A(n38819), .Z(n38818) );
  NANDN U47956 ( .A(n38819), .B(n38817), .Z(n38813) );
  AND U47957 ( .A(n38820), .B(n38821), .Z(n38794) );
  NAND U47958 ( .A(n38822), .B(n38823), .Z(n38821) );
  NANDN U47959 ( .A(n38824), .B(n38825), .Z(n38823) );
  NANDN U47960 ( .A(n38825), .B(n38824), .Z(n38820) );
  IV U47961 ( .A(n38826), .Z(n38825) );
  NAND U47962 ( .A(n38827), .B(n38828), .Z(n38797) );
  NANDN U47963 ( .A(n38829), .B(n38830), .Z(n38828) );
  NANDN U47964 ( .A(n38831), .B(n38832), .Z(n38830) );
  NANDN U47965 ( .A(n38832), .B(n38831), .Z(n38827) );
  IV U47966 ( .A(n38833), .Z(n38831) );
  AND U47967 ( .A(n38834), .B(n38835), .Z(n38800) );
  NAND U47968 ( .A(n38836), .B(n38837), .Z(n38835) );
  NANDN U47969 ( .A(n38838), .B(n38839), .Z(n38837) );
  NANDN U47970 ( .A(n38839), .B(n38838), .Z(n38834) );
  XOR U47971 ( .A(n38810), .B(n38840), .Z(n38802) );
  XNOR U47972 ( .A(n38807), .B(n38809), .Z(n38840) );
  AND U47973 ( .A(n38841), .B(n38842), .Z(n38809) );
  NANDN U47974 ( .A(n38843), .B(n38844), .Z(n38842) );
  OR U47975 ( .A(n38845), .B(n38846), .Z(n38844) );
  IV U47976 ( .A(n38847), .Z(n38846) );
  NANDN U47977 ( .A(n38847), .B(n38845), .Z(n38841) );
  AND U47978 ( .A(n38848), .B(n38849), .Z(n38807) );
  NAND U47979 ( .A(n38850), .B(n38851), .Z(n38849) );
  NANDN U47980 ( .A(n38852), .B(n38853), .Z(n38851) );
  NANDN U47981 ( .A(n38853), .B(n38852), .Z(n38848) );
  IV U47982 ( .A(n38854), .Z(n38853) );
  NAND U47983 ( .A(n38855), .B(n38856), .Z(n38810) );
  NANDN U47984 ( .A(n38857), .B(n38858), .Z(n38856) );
  NANDN U47985 ( .A(n38859), .B(n38860), .Z(n38858) );
  NANDN U47986 ( .A(n38860), .B(n38859), .Z(n38855) );
  IV U47987 ( .A(n38861), .Z(n38859) );
  XOR U47988 ( .A(n38836), .B(n38862), .Z(N61932) );
  XNOR U47989 ( .A(n38839), .B(n38838), .Z(n38862) );
  XNOR U47990 ( .A(n38850), .B(n38863), .Z(n38838) );
  XNOR U47991 ( .A(n38854), .B(n38852), .Z(n38863) );
  XOR U47992 ( .A(n38860), .B(n38864), .Z(n38852) );
  XNOR U47993 ( .A(n38857), .B(n38861), .Z(n38864) );
  AND U47994 ( .A(n38865), .B(n38866), .Z(n38861) );
  NAND U47995 ( .A(n38867), .B(n38868), .Z(n38866) );
  NAND U47996 ( .A(n38869), .B(n38870), .Z(n38865) );
  AND U47997 ( .A(n38871), .B(n38872), .Z(n38857) );
  NAND U47998 ( .A(n38873), .B(n38874), .Z(n38872) );
  NAND U47999 ( .A(n38875), .B(n38876), .Z(n38871) );
  NANDN U48000 ( .A(n38877), .B(n38878), .Z(n38860) );
  ANDN U48001 ( .B(n38879), .A(n38880), .Z(n38854) );
  XNOR U48002 ( .A(n38845), .B(n38881), .Z(n38850) );
  XNOR U48003 ( .A(n38843), .B(n38847), .Z(n38881) );
  AND U48004 ( .A(n38882), .B(n38883), .Z(n38847) );
  NAND U48005 ( .A(n38884), .B(n38885), .Z(n38883) );
  NAND U48006 ( .A(n38886), .B(n38887), .Z(n38882) );
  AND U48007 ( .A(n38888), .B(n38889), .Z(n38843) );
  NAND U48008 ( .A(n38890), .B(n38891), .Z(n38889) );
  NAND U48009 ( .A(n38892), .B(n38893), .Z(n38888) );
  AND U48010 ( .A(n38894), .B(n38895), .Z(n38845) );
  NAND U48011 ( .A(n38896), .B(n38897), .Z(n38839) );
  XNOR U48012 ( .A(n38822), .B(n38898), .Z(n38836) );
  XNOR U48013 ( .A(n38826), .B(n38824), .Z(n38898) );
  XOR U48014 ( .A(n38832), .B(n38899), .Z(n38824) );
  XNOR U48015 ( .A(n38829), .B(n38833), .Z(n38899) );
  AND U48016 ( .A(n38900), .B(n38901), .Z(n38833) );
  NAND U48017 ( .A(n38902), .B(n38903), .Z(n38901) );
  NAND U48018 ( .A(n38904), .B(n38905), .Z(n38900) );
  AND U48019 ( .A(n38906), .B(n38907), .Z(n38829) );
  NAND U48020 ( .A(n38908), .B(n38909), .Z(n38907) );
  NAND U48021 ( .A(n38910), .B(n38911), .Z(n38906) );
  NANDN U48022 ( .A(n38912), .B(n38913), .Z(n38832) );
  ANDN U48023 ( .B(n38914), .A(n38915), .Z(n38826) );
  XNOR U48024 ( .A(n38817), .B(n38916), .Z(n38822) );
  XNOR U48025 ( .A(n38815), .B(n38819), .Z(n38916) );
  AND U48026 ( .A(n38917), .B(n38918), .Z(n38819) );
  NAND U48027 ( .A(n38919), .B(n38920), .Z(n38918) );
  NAND U48028 ( .A(n38921), .B(n38922), .Z(n38917) );
  AND U48029 ( .A(n38923), .B(n38924), .Z(n38815) );
  NAND U48030 ( .A(n38925), .B(n38926), .Z(n38924) );
  NAND U48031 ( .A(n38927), .B(n38928), .Z(n38923) );
  AND U48032 ( .A(n38929), .B(n38930), .Z(n38817) );
  XOR U48033 ( .A(n38897), .B(n38896), .Z(N61931) );
  XNOR U48034 ( .A(n38914), .B(n38915), .Z(n38896) );
  XNOR U48035 ( .A(n38929), .B(n38930), .Z(n38915) );
  XOR U48036 ( .A(n38926), .B(n38925), .Z(n38930) );
  XOR U48037 ( .A(y[2484]), .B(x[2484]), .Z(n38925) );
  XOR U48038 ( .A(n38928), .B(n38927), .Z(n38926) );
  XOR U48039 ( .A(y[2486]), .B(x[2486]), .Z(n38927) );
  XOR U48040 ( .A(y[2485]), .B(x[2485]), .Z(n38928) );
  XOR U48041 ( .A(n38920), .B(n38919), .Z(n38929) );
  XOR U48042 ( .A(n38922), .B(n38921), .Z(n38919) );
  XOR U48043 ( .A(y[2483]), .B(x[2483]), .Z(n38921) );
  XOR U48044 ( .A(y[2482]), .B(x[2482]), .Z(n38922) );
  XOR U48045 ( .A(y[2481]), .B(x[2481]), .Z(n38920) );
  XNOR U48046 ( .A(n38913), .B(n38912), .Z(n38914) );
  XNOR U48047 ( .A(n38909), .B(n38908), .Z(n38912) );
  XOR U48048 ( .A(n38911), .B(n38910), .Z(n38908) );
  XOR U48049 ( .A(y[2480]), .B(x[2480]), .Z(n38910) );
  XOR U48050 ( .A(y[2479]), .B(x[2479]), .Z(n38911) );
  XOR U48051 ( .A(y[2478]), .B(x[2478]), .Z(n38909) );
  XOR U48052 ( .A(n38903), .B(n38902), .Z(n38913) );
  XOR U48053 ( .A(n38905), .B(n38904), .Z(n38902) );
  XOR U48054 ( .A(y[2477]), .B(x[2477]), .Z(n38904) );
  XOR U48055 ( .A(y[2476]), .B(x[2476]), .Z(n38905) );
  XOR U48056 ( .A(y[2475]), .B(x[2475]), .Z(n38903) );
  XNOR U48057 ( .A(n38879), .B(n38880), .Z(n38897) );
  XNOR U48058 ( .A(n38894), .B(n38895), .Z(n38880) );
  XOR U48059 ( .A(n38891), .B(n38890), .Z(n38895) );
  XOR U48060 ( .A(y[2472]), .B(x[2472]), .Z(n38890) );
  XOR U48061 ( .A(n38893), .B(n38892), .Z(n38891) );
  XOR U48062 ( .A(y[2474]), .B(x[2474]), .Z(n38892) );
  XOR U48063 ( .A(y[2473]), .B(x[2473]), .Z(n38893) );
  XOR U48064 ( .A(n38885), .B(n38884), .Z(n38894) );
  XOR U48065 ( .A(n38887), .B(n38886), .Z(n38884) );
  XOR U48066 ( .A(y[2471]), .B(x[2471]), .Z(n38886) );
  XOR U48067 ( .A(y[2470]), .B(x[2470]), .Z(n38887) );
  XOR U48068 ( .A(y[2469]), .B(x[2469]), .Z(n38885) );
  XNOR U48069 ( .A(n38878), .B(n38877), .Z(n38879) );
  XNOR U48070 ( .A(n38874), .B(n38873), .Z(n38877) );
  XOR U48071 ( .A(n38876), .B(n38875), .Z(n38873) );
  XOR U48072 ( .A(y[2468]), .B(x[2468]), .Z(n38875) );
  XOR U48073 ( .A(y[2467]), .B(x[2467]), .Z(n38876) );
  XOR U48074 ( .A(y[2466]), .B(x[2466]), .Z(n38874) );
  XOR U48075 ( .A(n38868), .B(n38867), .Z(n38878) );
  XOR U48076 ( .A(n38870), .B(n38869), .Z(n38867) );
  XOR U48077 ( .A(y[2465]), .B(x[2465]), .Z(n38869) );
  XOR U48078 ( .A(y[2464]), .B(x[2464]), .Z(n38870) );
  XOR U48079 ( .A(y[2463]), .B(x[2463]), .Z(n38868) );
  NAND U48080 ( .A(n38931), .B(n38932), .Z(N61922) );
  NAND U48081 ( .A(n38933), .B(n38934), .Z(n38932) );
  NANDN U48082 ( .A(n38935), .B(n38936), .Z(n38934) );
  NANDN U48083 ( .A(n38936), .B(n38935), .Z(n38931) );
  XOR U48084 ( .A(n38935), .B(n38937), .Z(N61921) );
  XNOR U48085 ( .A(n38933), .B(n38936), .Z(n38937) );
  NAND U48086 ( .A(n38938), .B(n38939), .Z(n38936) );
  NAND U48087 ( .A(n38940), .B(n38941), .Z(n38939) );
  NANDN U48088 ( .A(n38942), .B(n38943), .Z(n38941) );
  NANDN U48089 ( .A(n38943), .B(n38942), .Z(n38938) );
  AND U48090 ( .A(n38944), .B(n38945), .Z(n38933) );
  NAND U48091 ( .A(n38946), .B(n38947), .Z(n38945) );
  NANDN U48092 ( .A(n38948), .B(n38949), .Z(n38947) );
  NANDN U48093 ( .A(n38949), .B(n38948), .Z(n38944) );
  IV U48094 ( .A(n38950), .Z(n38949) );
  AND U48095 ( .A(n38951), .B(n38952), .Z(n38935) );
  NAND U48096 ( .A(n38953), .B(n38954), .Z(n38952) );
  NANDN U48097 ( .A(n38955), .B(n38956), .Z(n38954) );
  NANDN U48098 ( .A(n38956), .B(n38955), .Z(n38951) );
  XOR U48099 ( .A(n38948), .B(n38957), .Z(N61920) );
  XNOR U48100 ( .A(n38946), .B(n38950), .Z(n38957) );
  XOR U48101 ( .A(n38943), .B(n38958), .Z(n38950) );
  XNOR U48102 ( .A(n38940), .B(n38942), .Z(n38958) );
  AND U48103 ( .A(n38959), .B(n38960), .Z(n38942) );
  NANDN U48104 ( .A(n38961), .B(n38962), .Z(n38960) );
  OR U48105 ( .A(n38963), .B(n38964), .Z(n38962) );
  IV U48106 ( .A(n38965), .Z(n38964) );
  NANDN U48107 ( .A(n38965), .B(n38963), .Z(n38959) );
  AND U48108 ( .A(n38966), .B(n38967), .Z(n38940) );
  NAND U48109 ( .A(n38968), .B(n38969), .Z(n38967) );
  NANDN U48110 ( .A(n38970), .B(n38971), .Z(n38969) );
  NANDN U48111 ( .A(n38971), .B(n38970), .Z(n38966) );
  IV U48112 ( .A(n38972), .Z(n38971) );
  NAND U48113 ( .A(n38973), .B(n38974), .Z(n38943) );
  NANDN U48114 ( .A(n38975), .B(n38976), .Z(n38974) );
  NANDN U48115 ( .A(n38977), .B(n38978), .Z(n38976) );
  NANDN U48116 ( .A(n38978), .B(n38977), .Z(n38973) );
  IV U48117 ( .A(n38979), .Z(n38977) );
  AND U48118 ( .A(n38980), .B(n38981), .Z(n38946) );
  NAND U48119 ( .A(n38982), .B(n38983), .Z(n38981) );
  NANDN U48120 ( .A(n38984), .B(n38985), .Z(n38983) );
  NANDN U48121 ( .A(n38985), .B(n38984), .Z(n38980) );
  XOR U48122 ( .A(n38956), .B(n38986), .Z(n38948) );
  XNOR U48123 ( .A(n38953), .B(n38955), .Z(n38986) );
  AND U48124 ( .A(n38987), .B(n38988), .Z(n38955) );
  NANDN U48125 ( .A(n38989), .B(n38990), .Z(n38988) );
  OR U48126 ( .A(n38991), .B(n38992), .Z(n38990) );
  IV U48127 ( .A(n38993), .Z(n38992) );
  NANDN U48128 ( .A(n38993), .B(n38991), .Z(n38987) );
  AND U48129 ( .A(n38994), .B(n38995), .Z(n38953) );
  NAND U48130 ( .A(n38996), .B(n38997), .Z(n38995) );
  NANDN U48131 ( .A(n38998), .B(n38999), .Z(n38997) );
  NANDN U48132 ( .A(n38999), .B(n38998), .Z(n38994) );
  IV U48133 ( .A(n39000), .Z(n38999) );
  NAND U48134 ( .A(n39001), .B(n39002), .Z(n38956) );
  NANDN U48135 ( .A(n39003), .B(n39004), .Z(n39002) );
  NANDN U48136 ( .A(n39005), .B(n39006), .Z(n39004) );
  NANDN U48137 ( .A(n39006), .B(n39005), .Z(n39001) );
  IV U48138 ( .A(n39007), .Z(n39005) );
  XOR U48139 ( .A(n38982), .B(n39008), .Z(N61919) );
  XNOR U48140 ( .A(n38985), .B(n38984), .Z(n39008) );
  XNOR U48141 ( .A(n38996), .B(n39009), .Z(n38984) );
  XNOR U48142 ( .A(n39000), .B(n38998), .Z(n39009) );
  XOR U48143 ( .A(n39006), .B(n39010), .Z(n38998) );
  XNOR U48144 ( .A(n39003), .B(n39007), .Z(n39010) );
  AND U48145 ( .A(n39011), .B(n39012), .Z(n39007) );
  NAND U48146 ( .A(n39013), .B(n39014), .Z(n39012) );
  NAND U48147 ( .A(n39015), .B(n39016), .Z(n39011) );
  AND U48148 ( .A(n39017), .B(n39018), .Z(n39003) );
  NAND U48149 ( .A(n39019), .B(n39020), .Z(n39018) );
  NAND U48150 ( .A(n39021), .B(n39022), .Z(n39017) );
  NANDN U48151 ( .A(n39023), .B(n39024), .Z(n39006) );
  ANDN U48152 ( .B(n39025), .A(n39026), .Z(n39000) );
  XNOR U48153 ( .A(n38991), .B(n39027), .Z(n38996) );
  XNOR U48154 ( .A(n38989), .B(n38993), .Z(n39027) );
  AND U48155 ( .A(n39028), .B(n39029), .Z(n38993) );
  NAND U48156 ( .A(n39030), .B(n39031), .Z(n39029) );
  NAND U48157 ( .A(n39032), .B(n39033), .Z(n39028) );
  AND U48158 ( .A(n39034), .B(n39035), .Z(n38989) );
  NAND U48159 ( .A(n39036), .B(n39037), .Z(n39035) );
  NAND U48160 ( .A(n39038), .B(n39039), .Z(n39034) );
  AND U48161 ( .A(n39040), .B(n39041), .Z(n38991) );
  NAND U48162 ( .A(n39042), .B(n39043), .Z(n38985) );
  XNOR U48163 ( .A(n38968), .B(n39044), .Z(n38982) );
  XNOR U48164 ( .A(n38972), .B(n38970), .Z(n39044) );
  XOR U48165 ( .A(n38978), .B(n39045), .Z(n38970) );
  XNOR U48166 ( .A(n38975), .B(n38979), .Z(n39045) );
  AND U48167 ( .A(n39046), .B(n39047), .Z(n38979) );
  NAND U48168 ( .A(n39048), .B(n39049), .Z(n39047) );
  NAND U48169 ( .A(n39050), .B(n39051), .Z(n39046) );
  AND U48170 ( .A(n39052), .B(n39053), .Z(n38975) );
  NAND U48171 ( .A(n39054), .B(n39055), .Z(n39053) );
  NAND U48172 ( .A(n39056), .B(n39057), .Z(n39052) );
  NANDN U48173 ( .A(n39058), .B(n39059), .Z(n38978) );
  ANDN U48174 ( .B(n39060), .A(n39061), .Z(n38972) );
  XNOR U48175 ( .A(n38963), .B(n39062), .Z(n38968) );
  XNOR U48176 ( .A(n38961), .B(n38965), .Z(n39062) );
  AND U48177 ( .A(n39063), .B(n39064), .Z(n38965) );
  NAND U48178 ( .A(n39065), .B(n39066), .Z(n39064) );
  NAND U48179 ( .A(n39067), .B(n39068), .Z(n39063) );
  AND U48180 ( .A(n39069), .B(n39070), .Z(n38961) );
  NAND U48181 ( .A(n39071), .B(n39072), .Z(n39070) );
  NAND U48182 ( .A(n39073), .B(n39074), .Z(n39069) );
  AND U48183 ( .A(n39075), .B(n39076), .Z(n38963) );
  XOR U48184 ( .A(n39043), .B(n39042), .Z(N61918) );
  XNOR U48185 ( .A(n39060), .B(n39061), .Z(n39042) );
  XNOR U48186 ( .A(n39075), .B(n39076), .Z(n39061) );
  XOR U48187 ( .A(n39072), .B(n39071), .Z(n39076) );
  XOR U48188 ( .A(y[2460]), .B(x[2460]), .Z(n39071) );
  XOR U48189 ( .A(n39074), .B(n39073), .Z(n39072) );
  XOR U48190 ( .A(y[2462]), .B(x[2462]), .Z(n39073) );
  XOR U48191 ( .A(y[2461]), .B(x[2461]), .Z(n39074) );
  XOR U48192 ( .A(n39066), .B(n39065), .Z(n39075) );
  XOR U48193 ( .A(n39068), .B(n39067), .Z(n39065) );
  XOR U48194 ( .A(y[2459]), .B(x[2459]), .Z(n39067) );
  XOR U48195 ( .A(y[2458]), .B(x[2458]), .Z(n39068) );
  XOR U48196 ( .A(y[2457]), .B(x[2457]), .Z(n39066) );
  XNOR U48197 ( .A(n39059), .B(n39058), .Z(n39060) );
  XNOR U48198 ( .A(n39055), .B(n39054), .Z(n39058) );
  XOR U48199 ( .A(n39057), .B(n39056), .Z(n39054) );
  XOR U48200 ( .A(y[2456]), .B(x[2456]), .Z(n39056) );
  XOR U48201 ( .A(y[2455]), .B(x[2455]), .Z(n39057) );
  XOR U48202 ( .A(y[2454]), .B(x[2454]), .Z(n39055) );
  XOR U48203 ( .A(n39049), .B(n39048), .Z(n39059) );
  XOR U48204 ( .A(n39051), .B(n39050), .Z(n39048) );
  XOR U48205 ( .A(y[2453]), .B(x[2453]), .Z(n39050) );
  XOR U48206 ( .A(y[2452]), .B(x[2452]), .Z(n39051) );
  XOR U48207 ( .A(y[2451]), .B(x[2451]), .Z(n39049) );
  XNOR U48208 ( .A(n39025), .B(n39026), .Z(n39043) );
  XNOR U48209 ( .A(n39040), .B(n39041), .Z(n39026) );
  XOR U48210 ( .A(n39037), .B(n39036), .Z(n39041) );
  XOR U48211 ( .A(y[2448]), .B(x[2448]), .Z(n39036) );
  XOR U48212 ( .A(n39039), .B(n39038), .Z(n39037) );
  XOR U48213 ( .A(y[2450]), .B(x[2450]), .Z(n39038) );
  XOR U48214 ( .A(y[2449]), .B(x[2449]), .Z(n39039) );
  XOR U48215 ( .A(n39031), .B(n39030), .Z(n39040) );
  XOR U48216 ( .A(n39033), .B(n39032), .Z(n39030) );
  XOR U48217 ( .A(y[2447]), .B(x[2447]), .Z(n39032) );
  XOR U48218 ( .A(y[2446]), .B(x[2446]), .Z(n39033) );
  XOR U48219 ( .A(y[2445]), .B(x[2445]), .Z(n39031) );
  XNOR U48220 ( .A(n39024), .B(n39023), .Z(n39025) );
  XNOR U48221 ( .A(n39020), .B(n39019), .Z(n39023) );
  XOR U48222 ( .A(n39022), .B(n39021), .Z(n39019) );
  XOR U48223 ( .A(y[2444]), .B(x[2444]), .Z(n39021) );
  XOR U48224 ( .A(y[2443]), .B(x[2443]), .Z(n39022) );
  XOR U48225 ( .A(y[2442]), .B(x[2442]), .Z(n39020) );
  XOR U48226 ( .A(n39014), .B(n39013), .Z(n39024) );
  XOR U48227 ( .A(n39016), .B(n39015), .Z(n39013) );
  XOR U48228 ( .A(y[2441]), .B(x[2441]), .Z(n39015) );
  XOR U48229 ( .A(y[2440]), .B(x[2440]), .Z(n39016) );
  XOR U48230 ( .A(y[2439]), .B(x[2439]), .Z(n39014) );
  NAND U48231 ( .A(n39077), .B(n39078), .Z(N61909) );
  NAND U48232 ( .A(n39079), .B(n39080), .Z(n39078) );
  NANDN U48233 ( .A(n39081), .B(n39082), .Z(n39080) );
  NANDN U48234 ( .A(n39082), .B(n39081), .Z(n39077) );
  XOR U48235 ( .A(n39081), .B(n39083), .Z(N61908) );
  XNOR U48236 ( .A(n39079), .B(n39082), .Z(n39083) );
  NAND U48237 ( .A(n39084), .B(n39085), .Z(n39082) );
  NAND U48238 ( .A(n39086), .B(n39087), .Z(n39085) );
  NANDN U48239 ( .A(n39088), .B(n39089), .Z(n39087) );
  NANDN U48240 ( .A(n39089), .B(n39088), .Z(n39084) );
  AND U48241 ( .A(n39090), .B(n39091), .Z(n39079) );
  NAND U48242 ( .A(n39092), .B(n39093), .Z(n39091) );
  NANDN U48243 ( .A(n39094), .B(n39095), .Z(n39093) );
  NANDN U48244 ( .A(n39095), .B(n39094), .Z(n39090) );
  IV U48245 ( .A(n39096), .Z(n39095) );
  AND U48246 ( .A(n39097), .B(n39098), .Z(n39081) );
  NAND U48247 ( .A(n39099), .B(n39100), .Z(n39098) );
  NANDN U48248 ( .A(n39101), .B(n39102), .Z(n39100) );
  NANDN U48249 ( .A(n39102), .B(n39101), .Z(n39097) );
  XOR U48250 ( .A(n39094), .B(n39103), .Z(N61907) );
  XNOR U48251 ( .A(n39092), .B(n39096), .Z(n39103) );
  XOR U48252 ( .A(n39089), .B(n39104), .Z(n39096) );
  XNOR U48253 ( .A(n39086), .B(n39088), .Z(n39104) );
  AND U48254 ( .A(n39105), .B(n39106), .Z(n39088) );
  NANDN U48255 ( .A(n39107), .B(n39108), .Z(n39106) );
  OR U48256 ( .A(n39109), .B(n39110), .Z(n39108) );
  IV U48257 ( .A(n39111), .Z(n39110) );
  NANDN U48258 ( .A(n39111), .B(n39109), .Z(n39105) );
  AND U48259 ( .A(n39112), .B(n39113), .Z(n39086) );
  NAND U48260 ( .A(n39114), .B(n39115), .Z(n39113) );
  NANDN U48261 ( .A(n39116), .B(n39117), .Z(n39115) );
  NANDN U48262 ( .A(n39117), .B(n39116), .Z(n39112) );
  IV U48263 ( .A(n39118), .Z(n39117) );
  NAND U48264 ( .A(n39119), .B(n39120), .Z(n39089) );
  NANDN U48265 ( .A(n39121), .B(n39122), .Z(n39120) );
  NANDN U48266 ( .A(n39123), .B(n39124), .Z(n39122) );
  NANDN U48267 ( .A(n39124), .B(n39123), .Z(n39119) );
  IV U48268 ( .A(n39125), .Z(n39123) );
  AND U48269 ( .A(n39126), .B(n39127), .Z(n39092) );
  NAND U48270 ( .A(n39128), .B(n39129), .Z(n39127) );
  NANDN U48271 ( .A(n39130), .B(n39131), .Z(n39129) );
  NANDN U48272 ( .A(n39131), .B(n39130), .Z(n39126) );
  XOR U48273 ( .A(n39102), .B(n39132), .Z(n39094) );
  XNOR U48274 ( .A(n39099), .B(n39101), .Z(n39132) );
  AND U48275 ( .A(n39133), .B(n39134), .Z(n39101) );
  NANDN U48276 ( .A(n39135), .B(n39136), .Z(n39134) );
  OR U48277 ( .A(n39137), .B(n39138), .Z(n39136) );
  IV U48278 ( .A(n39139), .Z(n39138) );
  NANDN U48279 ( .A(n39139), .B(n39137), .Z(n39133) );
  AND U48280 ( .A(n39140), .B(n39141), .Z(n39099) );
  NAND U48281 ( .A(n39142), .B(n39143), .Z(n39141) );
  NANDN U48282 ( .A(n39144), .B(n39145), .Z(n39143) );
  NANDN U48283 ( .A(n39145), .B(n39144), .Z(n39140) );
  IV U48284 ( .A(n39146), .Z(n39145) );
  NAND U48285 ( .A(n39147), .B(n39148), .Z(n39102) );
  NANDN U48286 ( .A(n39149), .B(n39150), .Z(n39148) );
  NANDN U48287 ( .A(n39151), .B(n39152), .Z(n39150) );
  NANDN U48288 ( .A(n39152), .B(n39151), .Z(n39147) );
  IV U48289 ( .A(n39153), .Z(n39151) );
  XOR U48290 ( .A(n39128), .B(n39154), .Z(N61906) );
  XNOR U48291 ( .A(n39131), .B(n39130), .Z(n39154) );
  XNOR U48292 ( .A(n39142), .B(n39155), .Z(n39130) );
  XNOR U48293 ( .A(n39146), .B(n39144), .Z(n39155) );
  XOR U48294 ( .A(n39152), .B(n39156), .Z(n39144) );
  XNOR U48295 ( .A(n39149), .B(n39153), .Z(n39156) );
  AND U48296 ( .A(n39157), .B(n39158), .Z(n39153) );
  NAND U48297 ( .A(n39159), .B(n39160), .Z(n39158) );
  NAND U48298 ( .A(n39161), .B(n39162), .Z(n39157) );
  AND U48299 ( .A(n39163), .B(n39164), .Z(n39149) );
  NAND U48300 ( .A(n39165), .B(n39166), .Z(n39164) );
  NAND U48301 ( .A(n39167), .B(n39168), .Z(n39163) );
  NANDN U48302 ( .A(n39169), .B(n39170), .Z(n39152) );
  ANDN U48303 ( .B(n39171), .A(n39172), .Z(n39146) );
  XNOR U48304 ( .A(n39137), .B(n39173), .Z(n39142) );
  XNOR U48305 ( .A(n39135), .B(n39139), .Z(n39173) );
  AND U48306 ( .A(n39174), .B(n39175), .Z(n39139) );
  NAND U48307 ( .A(n39176), .B(n39177), .Z(n39175) );
  NAND U48308 ( .A(n39178), .B(n39179), .Z(n39174) );
  AND U48309 ( .A(n39180), .B(n39181), .Z(n39135) );
  NAND U48310 ( .A(n39182), .B(n39183), .Z(n39181) );
  NAND U48311 ( .A(n39184), .B(n39185), .Z(n39180) );
  AND U48312 ( .A(n39186), .B(n39187), .Z(n39137) );
  NAND U48313 ( .A(n39188), .B(n39189), .Z(n39131) );
  XNOR U48314 ( .A(n39114), .B(n39190), .Z(n39128) );
  XNOR U48315 ( .A(n39118), .B(n39116), .Z(n39190) );
  XOR U48316 ( .A(n39124), .B(n39191), .Z(n39116) );
  XNOR U48317 ( .A(n39121), .B(n39125), .Z(n39191) );
  AND U48318 ( .A(n39192), .B(n39193), .Z(n39125) );
  NAND U48319 ( .A(n39194), .B(n39195), .Z(n39193) );
  NAND U48320 ( .A(n39196), .B(n39197), .Z(n39192) );
  AND U48321 ( .A(n39198), .B(n39199), .Z(n39121) );
  NAND U48322 ( .A(n39200), .B(n39201), .Z(n39199) );
  NAND U48323 ( .A(n39202), .B(n39203), .Z(n39198) );
  NANDN U48324 ( .A(n39204), .B(n39205), .Z(n39124) );
  ANDN U48325 ( .B(n39206), .A(n39207), .Z(n39118) );
  XNOR U48326 ( .A(n39109), .B(n39208), .Z(n39114) );
  XNOR U48327 ( .A(n39107), .B(n39111), .Z(n39208) );
  AND U48328 ( .A(n39209), .B(n39210), .Z(n39111) );
  NAND U48329 ( .A(n39211), .B(n39212), .Z(n39210) );
  NAND U48330 ( .A(n39213), .B(n39214), .Z(n39209) );
  AND U48331 ( .A(n39215), .B(n39216), .Z(n39107) );
  NAND U48332 ( .A(n39217), .B(n39218), .Z(n39216) );
  NAND U48333 ( .A(n39219), .B(n39220), .Z(n39215) );
  AND U48334 ( .A(n39221), .B(n39222), .Z(n39109) );
  XOR U48335 ( .A(n39189), .B(n39188), .Z(N61905) );
  XNOR U48336 ( .A(n39206), .B(n39207), .Z(n39188) );
  XNOR U48337 ( .A(n39221), .B(n39222), .Z(n39207) );
  XOR U48338 ( .A(n39218), .B(n39217), .Z(n39222) );
  XOR U48339 ( .A(y[2436]), .B(x[2436]), .Z(n39217) );
  XOR U48340 ( .A(n39220), .B(n39219), .Z(n39218) );
  XOR U48341 ( .A(y[2438]), .B(x[2438]), .Z(n39219) );
  XOR U48342 ( .A(y[2437]), .B(x[2437]), .Z(n39220) );
  XOR U48343 ( .A(n39212), .B(n39211), .Z(n39221) );
  XOR U48344 ( .A(n39214), .B(n39213), .Z(n39211) );
  XOR U48345 ( .A(y[2435]), .B(x[2435]), .Z(n39213) );
  XOR U48346 ( .A(y[2434]), .B(x[2434]), .Z(n39214) );
  XOR U48347 ( .A(y[2433]), .B(x[2433]), .Z(n39212) );
  XNOR U48348 ( .A(n39205), .B(n39204), .Z(n39206) );
  XNOR U48349 ( .A(n39201), .B(n39200), .Z(n39204) );
  XOR U48350 ( .A(n39203), .B(n39202), .Z(n39200) );
  XOR U48351 ( .A(y[2432]), .B(x[2432]), .Z(n39202) );
  XOR U48352 ( .A(y[2431]), .B(x[2431]), .Z(n39203) );
  XOR U48353 ( .A(y[2430]), .B(x[2430]), .Z(n39201) );
  XOR U48354 ( .A(n39195), .B(n39194), .Z(n39205) );
  XOR U48355 ( .A(n39197), .B(n39196), .Z(n39194) );
  XOR U48356 ( .A(y[2429]), .B(x[2429]), .Z(n39196) );
  XOR U48357 ( .A(y[2428]), .B(x[2428]), .Z(n39197) );
  XOR U48358 ( .A(y[2427]), .B(x[2427]), .Z(n39195) );
  XNOR U48359 ( .A(n39171), .B(n39172), .Z(n39189) );
  XNOR U48360 ( .A(n39186), .B(n39187), .Z(n39172) );
  XOR U48361 ( .A(n39183), .B(n39182), .Z(n39187) );
  XOR U48362 ( .A(y[2424]), .B(x[2424]), .Z(n39182) );
  XOR U48363 ( .A(n39185), .B(n39184), .Z(n39183) );
  XOR U48364 ( .A(y[2426]), .B(x[2426]), .Z(n39184) );
  XOR U48365 ( .A(y[2425]), .B(x[2425]), .Z(n39185) );
  XOR U48366 ( .A(n39177), .B(n39176), .Z(n39186) );
  XOR U48367 ( .A(n39179), .B(n39178), .Z(n39176) );
  XOR U48368 ( .A(y[2423]), .B(x[2423]), .Z(n39178) );
  XOR U48369 ( .A(y[2422]), .B(x[2422]), .Z(n39179) );
  XOR U48370 ( .A(y[2421]), .B(x[2421]), .Z(n39177) );
  XNOR U48371 ( .A(n39170), .B(n39169), .Z(n39171) );
  XNOR U48372 ( .A(n39166), .B(n39165), .Z(n39169) );
  XOR U48373 ( .A(n39168), .B(n39167), .Z(n39165) );
  XOR U48374 ( .A(y[2420]), .B(x[2420]), .Z(n39167) );
  XOR U48375 ( .A(y[2419]), .B(x[2419]), .Z(n39168) );
  XOR U48376 ( .A(y[2418]), .B(x[2418]), .Z(n39166) );
  XOR U48377 ( .A(n39160), .B(n39159), .Z(n39170) );
  XOR U48378 ( .A(n39162), .B(n39161), .Z(n39159) );
  XOR U48379 ( .A(y[2417]), .B(x[2417]), .Z(n39161) );
  XOR U48380 ( .A(y[2416]), .B(x[2416]), .Z(n39162) );
  XOR U48381 ( .A(y[2415]), .B(x[2415]), .Z(n39160) );
  NAND U48382 ( .A(n39223), .B(n39224), .Z(N61896) );
  NAND U48383 ( .A(n39225), .B(n39226), .Z(n39224) );
  NANDN U48384 ( .A(n39227), .B(n39228), .Z(n39226) );
  NANDN U48385 ( .A(n39228), .B(n39227), .Z(n39223) );
  XOR U48386 ( .A(n39227), .B(n39229), .Z(N61895) );
  XNOR U48387 ( .A(n39225), .B(n39228), .Z(n39229) );
  NAND U48388 ( .A(n39230), .B(n39231), .Z(n39228) );
  NAND U48389 ( .A(n39232), .B(n39233), .Z(n39231) );
  NANDN U48390 ( .A(n39234), .B(n39235), .Z(n39233) );
  NANDN U48391 ( .A(n39235), .B(n39234), .Z(n39230) );
  AND U48392 ( .A(n39236), .B(n39237), .Z(n39225) );
  NAND U48393 ( .A(n39238), .B(n39239), .Z(n39237) );
  NANDN U48394 ( .A(n39240), .B(n39241), .Z(n39239) );
  NANDN U48395 ( .A(n39241), .B(n39240), .Z(n39236) );
  IV U48396 ( .A(n39242), .Z(n39241) );
  AND U48397 ( .A(n39243), .B(n39244), .Z(n39227) );
  NAND U48398 ( .A(n39245), .B(n39246), .Z(n39244) );
  NANDN U48399 ( .A(n39247), .B(n39248), .Z(n39246) );
  NANDN U48400 ( .A(n39248), .B(n39247), .Z(n39243) );
  XOR U48401 ( .A(n39240), .B(n39249), .Z(N61894) );
  XNOR U48402 ( .A(n39238), .B(n39242), .Z(n39249) );
  XOR U48403 ( .A(n39235), .B(n39250), .Z(n39242) );
  XNOR U48404 ( .A(n39232), .B(n39234), .Z(n39250) );
  AND U48405 ( .A(n39251), .B(n39252), .Z(n39234) );
  NANDN U48406 ( .A(n39253), .B(n39254), .Z(n39252) );
  OR U48407 ( .A(n39255), .B(n39256), .Z(n39254) );
  IV U48408 ( .A(n39257), .Z(n39256) );
  NANDN U48409 ( .A(n39257), .B(n39255), .Z(n39251) );
  AND U48410 ( .A(n39258), .B(n39259), .Z(n39232) );
  NAND U48411 ( .A(n39260), .B(n39261), .Z(n39259) );
  NANDN U48412 ( .A(n39262), .B(n39263), .Z(n39261) );
  NANDN U48413 ( .A(n39263), .B(n39262), .Z(n39258) );
  IV U48414 ( .A(n39264), .Z(n39263) );
  NAND U48415 ( .A(n39265), .B(n39266), .Z(n39235) );
  NANDN U48416 ( .A(n39267), .B(n39268), .Z(n39266) );
  NANDN U48417 ( .A(n39269), .B(n39270), .Z(n39268) );
  NANDN U48418 ( .A(n39270), .B(n39269), .Z(n39265) );
  IV U48419 ( .A(n39271), .Z(n39269) );
  AND U48420 ( .A(n39272), .B(n39273), .Z(n39238) );
  NAND U48421 ( .A(n39274), .B(n39275), .Z(n39273) );
  NANDN U48422 ( .A(n39276), .B(n39277), .Z(n39275) );
  NANDN U48423 ( .A(n39277), .B(n39276), .Z(n39272) );
  XOR U48424 ( .A(n39248), .B(n39278), .Z(n39240) );
  XNOR U48425 ( .A(n39245), .B(n39247), .Z(n39278) );
  AND U48426 ( .A(n39279), .B(n39280), .Z(n39247) );
  NANDN U48427 ( .A(n39281), .B(n39282), .Z(n39280) );
  OR U48428 ( .A(n39283), .B(n39284), .Z(n39282) );
  IV U48429 ( .A(n39285), .Z(n39284) );
  NANDN U48430 ( .A(n39285), .B(n39283), .Z(n39279) );
  AND U48431 ( .A(n39286), .B(n39287), .Z(n39245) );
  NAND U48432 ( .A(n39288), .B(n39289), .Z(n39287) );
  NANDN U48433 ( .A(n39290), .B(n39291), .Z(n39289) );
  NANDN U48434 ( .A(n39291), .B(n39290), .Z(n39286) );
  IV U48435 ( .A(n39292), .Z(n39291) );
  NAND U48436 ( .A(n39293), .B(n39294), .Z(n39248) );
  NANDN U48437 ( .A(n39295), .B(n39296), .Z(n39294) );
  NANDN U48438 ( .A(n39297), .B(n39298), .Z(n39296) );
  NANDN U48439 ( .A(n39298), .B(n39297), .Z(n39293) );
  IV U48440 ( .A(n39299), .Z(n39297) );
  XOR U48441 ( .A(n39274), .B(n39300), .Z(N61893) );
  XNOR U48442 ( .A(n39277), .B(n39276), .Z(n39300) );
  XNOR U48443 ( .A(n39288), .B(n39301), .Z(n39276) );
  XNOR U48444 ( .A(n39292), .B(n39290), .Z(n39301) );
  XOR U48445 ( .A(n39298), .B(n39302), .Z(n39290) );
  XNOR U48446 ( .A(n39295), .B(n39299), .Z(n39302) );
  AND U48447 ( .A(n39303), .B(n39304), .Z(n39299) );
  NAND U48448 ( .A(n39305), .B(n39306), .Z(n39304) );
  NAND U48449 ( .A(n39307), .B(n39308), .Z(n39303) );
  AND U48450 ( .A(n39309), .B(n39310), .Z(n39295) );
  NAND U48451 ( .A(n39311), .B(n39312), .Z(n39310) );
  NAND U48452 ( .A(n39313), .B(n39314), .Z(n39309) );
  NANDN U48453 ( .A(n39315), .B(n39316), .Z(n39298) );
  ANDN U48454 ( .B(n39317), .A(n39318), .Z(n39292) );
  XNOR U48455 ( .A(n39283), .B(n39319), .Z(n39288) );
  XNOR U48456 ( .A(n39281), .B(n39285), .Z(n39319) );
  AND U48457 ( .A(n39320), .B(n39321), .Z(n39285) );
  NAND U48458 ( .A(n39322), .B(n39323), .Z(n39321) );
  NAND U48459 ( .A(n39324), .B(n39325), .Z(n39320) );
  AND U48460 ( .A(n39326), .B(n39327), .Z(n39281) );
  NAND U48461 ( .A(n39328), .B(n39329), .Z(n39327) );
  NAND U48462 ( .A(n39330), .B(n39331), .Z(n39326) );
  AND U48463 ( .A(n39332), .B(n39333), .Z(n39283) );
  NAND U48464 ( .A(n39334), .B(n39335), .Z(n39277) );
  XNOR U48465 ( .A(n39260), .B(n39336), .Z(n39274) );
  XNOR U48466 ( .A(n39264), .B(n39262), .Z(n39336) );
  XOR U48467 ( .A(n39270), .B(n39337), .Z(n39262) );
  XNOR U48468 ( .A(n39267), .B(n39271), .Z(n39337) );
  AND U48469 ( .A(n39338), .B(n39339), .Z(n39271) );
  NAND U48470 ( .A(n39340), .B(n39341), .Z(n39339) );
  NAND U48471 ( .A(n39342), .B(n39343), .Z(n39338) );
  AND U48472 ( .A(n39344), .B(n39345), .Z(n39267) );
  NAND U48473 ( .A(n39346), .B(n39347), .Z(n39345) );
  NAND U48474 ( .A(n39348), .B(n39349), .Z(n39344) );
  NANDN U48475 ( .A(n39350), .B(n39351), .Z(n39270) );
  ANDN U48476 ( .B(n39352), .A(n39353), .Z(n39264) );
  XNOR U48477 ( .A(n39255), .B(n39354), .Z(n39260) );
  XNOR U48478 ( .A(n39253), .B(n39257), .Z(n39354) );
  AND U48479 ( .A(n39355), .B(n39356), .Z(n39257) );
  NAND U48480 ( .A(n39357), .B(n39358), .Z(n39356) );
  NAND U48481 ( .A(n39359), .B(n39360), .Z(n39355) );
  AND U48482 ( .A(n39361), .B(n39362), .Z(n39253) );
  NAND U48483 ( .A(n39363), .B(n39364), .Z(n39362) );
  NAND U48484 ( .A(n39365), .B(n39366), .Z(n39361) );
  AND U48485 ( .A(n39367), .B(n39368), .Z(n39255) );
  XOR U48486 ( .A(n39335), .B(n39334), .Z(N61892) );
  XNOR U48487 ( .A(n39352), .B(n39353), .Z(n39334) );
  XNOR U48488 ( .A(n39367), .B(n39368), .Z(n39353) );
  XOR U48489 ( .A(n39364), .B(n39363), .Z(n39368) );
  XOR U48490 ( .A(y[2412]), .B(x[2412]), .Z(n39363) );
  XOR U48491 ( .A(n39366), .B(n39365), .Z(n39364) );
  XOR U48492 ( .A(y[2414]), .B(x[2414]), .Z(n39365) );
  XOR U48493 ( .A(y[2413]), .B(x[2413]), .Z(n39366) );
  XOR U48494 ( .A(n39358), .B(n39357), .Z(n39367) );
  XOR U48495 ( .A(n39360), .B(n39359), .Z(n39357) );
  XOR U48496 ( .A(y[2411]), .B(x[2411]), .Z(n39359) );
  XOR U48497 ( .A(y[2410]), .B(x[2410]), .Z(n39360) );
  XOR U48498 ( .A(y[2409]), .B(x[2409]), .Z(n39358) );
  XNOR U48499 ( .A(n39351), .B(n39350), .Z(n39352) );
  XNOR U48500 ( .A(n39347), .B(n39346), .Z(n39350) );
  XOR U48501 ( .A(n39349), .B(n39348), .Z(n39346) );
  XOR U48502 ( .A(y[2408]), .B(x[2408]), .Z(n39348) );
  XOR U48503 ( .A(y[2407]), .B(x[2407]), .Z(n39349) );
  XOR U48504 ( .A(y[2406]), .B(x[2406]), .Z(n39347) );
  XOR U48505 ( .A(n39341), .B(n39340), .Z(n39351) );
  XOR U48506 ( .A(n39343), .B(n39342), .Z(n39340) );
  XOR U48507 ( .A(y[2405]), .B(x[2405]), .Z(n39342) );
  XOR U48508 ( .A(y[2404]), .B(x[2404]), .Z(n39343) );
  XOR U48509 ( .A(y[2403]), .B(x[2403]), .Z(n39341) );
  XNOR U48510 ( .A(n39317), .B(n39318), .Z(n39335) );
  XNOR U48511 ( .A(n39332), .B(n39333), .Z(n39318) );
  XOR U48512 ( .A(n39329), .B(n39328), .Z(n39333) );
  XOR U48513 ( .A(y[2400]), .B(x[2400]), .Z(n39328) );
  XOR U48514 ( .A(n39331), .B(n39330), .Z(n39329) );
  XOR U48515 ( .A(y[2402]), .B(x[2402]), .Z(n39330) );
  XOR U48516 ( .A(y[2401]), .B(x[2401]), .Z(n39331) );
  XOR U48517 ( .A(n39323), .B(n39322), .Z(n39332) );
  XOR U48518 ( .A(n39325), .B(n39324), .Z(n39322) );
  XOR U48519 ( .A(y[2399]), .B(x[2399]), .Z(n39324) );
  XOR U48520 ( .A(y[2398]), .B(x[2398]), .Z(n39325) );
  XOR U48521 ( .A(y[2397]), .B(x[2397]), .Z(n39323) );
  XNOR U48522 ( .A(n39316), .B(n39315), .Z(n39317) );
  XNOR U48523 ( .A(n39312), .B(n39311), .Z(n39315) );
  XOR U48524 ( .A(n39314), .B(n39313), .Z(n39311) );
  XOR U48525 ( .A(y[2396]), .B(x[2396]), .Z(n39313) );
  XOR U48526 ( .A(y[2395]), .B(x[2395]), .Z(n39314) );
  XOR U48527 ( .A(y[2394]), .B(x[2394]), .Z(n39312) );
  XOR U48528 ( .A(n39306), .B(n39305), .Z(n39316) );
  XOR U48529 ( .A(n39308), .B(n39307), .Z(n39305) );
  XOR U48530 ( .A(y[2393]), .B(x[2393]), .Z(n39307) );
  XOR U48531 ( .A(y[2392]), .B(x[2392]), .Z(n39308) );
  XOR U48532 ( .A(y[2391]), .B(x[2391]), .Z(n39306) );
  NAND U48533 ( .A(n39369), .B(n39370), .Z(N61883) );
  NAND U48534 ( .A(n39371), .B(n39372), .Z(n39370) );
  NANDN U48535 ( .A(n39373), .B(n39374), .Z(n39372) );
  NANDN U48536 ( .A(n39374), .B(n39373), .Z(n39369) );
  XOR U48537 ( .A(n39373), .B(n39375), .Z(N61882) );
  XNOR U48538 ( .A(n39371), .B(n39374), .Z(n39375) );
  NAND U48539 ( .A(n39376), .B(n39377), .Z(n39374) );
  NAND U48540 ( .A(n39378), .B(n39379), .Z(n39377) );
  NANDN U48541 ( .A(n39380), .B(n39381), .Z(n39379) );
  NANDN U48542 ( .A(n39381), .B(n39380), .Z(n39376) );
  AND U48543 ( .A(n39382), .B(n39383), .Z(n39371) );
  NAND U48544 ( .A(n39384), .B(n39385), .Z(n39383) );
  NANDN U48545 ( .A(n39386), .B(n39387), .Z(n39385) );
  NANDN U48546 ( .A(n39387), .B(n39386), .Z(n39382) );
  IV U48547 ( .A(n39388), .Z(n39387) );
  AND U48548 ( .A(n39389), .B(n39390), .Z(n39373) );
  NAND U48549 ( .A(n39391), .B(n39392), .Z(n39390) );
  NANDN U48550 ( .A(n39393), .B(n39394), .Z(n39392) );
  NANDN U48551 ( .A(n39394), .B(n39393), .Z(n39389) );
  XOR U48552 ( .A(n39386), .B(n39395), .Z(N61881) );
  XNOR U48553 ( .A(n39384), .B(n39388), .Z(n39395) );
  XOR U48554 ( .A(n39381), .B(n39396), .Z(n39388) );
  XNOR U48555 ( .A(n39378), .B(n39380), .Z(n39396) );
  AND U48556 ( .A(n39397), .B(n39398), .Z(n39380) );
  NANDN U48557 ( .A(n39399), .B(n39400), .Z(n39398) );
  OR U48558 ( .A(n39401), .B(n39402), .Z(n39400) );
  IV U48559 ( .A(n39403), .Z(n39402) );
  NANDN U48560 ( .A(n39403), .B(n39401), .Z(n39397) );
  AND U48561 ( .A(n39404), .B(n39405), .Z(n39378) );
  NAND U48562 ( .A(n39406), .B(n39407), .Z(n39405) );
  NANDN U48563 ( .A(n39408), .B(n39409), .Z(n39407) );
  NANDN U48564 ( .A(n39409), .B(n39408), .Z(n39404) );
  IV U48565 ( .A(n39410), .Z(n39409) );
  NAND U48566 ( .A(n39411), .B(n39412), .Z(n39381) );
  NANDN U48567 ( .A(n39413), .B(n39414), .Z(n39412) );
  NANDN U48568 ( .A(n39415), .B(n39416), .Z(n39414) );
  NANDN U48569 ( .A(n39416), .B(n39415), .Z(n39411) );
  IV U48570 ( .A(n39417), .Z(n39415) );
  AND U48571 ( .A(n39418), .B(n39419), .Z(n39384) );
  NAND U48572 ( .A(n39420), .B(n39421), .Z(n39419) );
  NANDN U48573 ( .A(n39422), .B(n39423), .Z(n39421) );
  NANDN U48574 ( .A(n39423), .B(n39422), .Z(n39418) );
  XOR U48575 ( .A(n39394), .B(n39424), .Z(n39386) );
  XNOR U48576 ( .A(n39391), .B(n39393), .Z(n39424) );
  AND U48577 ( .A(n39425), .B(n39426), .Z(n39393) );
  NANDN U48578 ( .A(n39427), .B(n39428), .Z(n39426) );
  OR U48579 ( .A(n39429), .B(n39430), .Z(n39428) );
  IV U48580 ( .A(n39431), .Z(n39430) );
  NANDN U48581 ( .A(n39431), .B(n39429), .Z(n39425) );
  AND U48582 ( .A(n39432), .B(n39433), .Z(n39391) );
  NAND U48583 ( .A(n39434), .B(n39435), .Z(n39433) );
  NANDN U48584 ( .A(n39436), .B(n39437), .Z(n39435) );
  NANDN U48585 ( .A(n39437), .B(n39436), .Z(n39432) );
  IV U48586 ( .A(n39438), .Z(n39437) );
  NAND U48587 ( .A(n39439), .B(n39440), .Z(n39394) );
  NANDN U48588 ( .A(n39441), .B(n39442), .Z(n39440) );
  NANDN U48589 ( .A(n39443), .B(n39444), .Z(n39442) );
  NANDN U48590 ( .A(n39444), .B(n39443), .Z(n39439) );
  IV U48591 ( .A(n39445), .Z(n39443) );
  XOR U48592 ( .A(n39420), .B(n39446), .Z(N61880) );
  XNOR U48593 ( .A(n39423), .B(n39422), .Z(n39446) );
  XNOR U48594 ( .A(n39434), .B(n39447), .Z(n39422) );
  XNOR U48595 ( .A(n39438), .B(n39436), .Z(n39447) );
  XOR U48596 ( .A(n39444), .B(n39448), .Z(n39436) );
  XNOR U48597 ( .A(n39441), .B(n39445), .Z(n39448) );
  AND U48598 ( .A(n39449), .B(n39450), .Z(n39445) );
  NAND U48599 ( .A(n39451), .B(n39452), .Z(n39450) );
  NAND U48600 ( .A(n39453), .B(n39454), .Z(n39449) );
  AND U48601 ( .A(n39455), .B(n39456), .Z(n39441) );
  NAND U48602 ( .A(n39457), .B(n39458), .Z(n39456) );
  NAND U48603 ( .A(n39459), .B(n39460), .Z(n39455) );
  NANDN U48604 ( .A(n39461), .B(n39462), .Z(n39444) );
  ANDN U48605 ( .B(n39463), .A(n39464), .Z(n39438) );
  XNOR U48606 ( .A(n39429), .B(n39465), .Z(n39434) );
  XNOR U48607 ( .A(n39427), .B(n39431), .Z(n39465) );
  AND U48608 ( .A(n39466), .B(n39467), .Z(n39431) );
  NAND U48609 ( .A(n39468), .B(n39469), .Z(n39467) );
  NAND U48610 ( .A(n39470), .B(n39471), .Z(n39466) );
  AND U48611 ( .A(n39472), .B(n39473), .Z(n39427) );
  NAND U48612 ( .A(n39474), .B(n39475), .Z(n39473) );
  NAND U48613 ( .A(n39476), .B(n39477), .Z(n39472) );
  AND U48614 ( .A(n39478), .B(n39479), .Z(n39429) );
  NAND U48615 ( .A(n39480), .B(n39481), .Z(n39423) );
  XNOR U48616 ( .A(n39406), .B(n39482), .Z(n39420) );
  XNOR U48617 ( .A(n39410), .B(n39408), .Z(n39482) );
  XOR U48618 ( .A(n39416), .B(n39483), .Z(n39408) );
  XNOR U48619 ( .A(n39413), .B(n39417), .Z(n39483) );
  AND U48620 ( .A(n39484), .B(n39485), .Z(n39417) );
  NAND U48621 ( .A(n39486), .B(n39487), .Z(n39485) );
  NAND U48622 ( .A(n39488), .B(n39489), .Z(n39484) );
  AND U48623 ( .A(n39490), .B(n39491), .Z(n39413) );
  NAND U48624 ( .A(n39492), .B(n39493), .Z(n39491) );
  NAND U48625 ( .A(n39494), .B(n39495), .Z(n39490) );
  NANDN U48626 ( .A(n39496), .B(n39497), .Z(n39416) );
  ANDN U48627 ( .B(n39498), .A(n39499), .Z(n39410) );
  XNOR U48628 ( .A(n39401), .B(n39500), .Z(n39406) );
  XNOR U48629 ( .A(n39399), .B(n39403), .Z(n39500) );
  AND U48630 ( .A(n39501), .B(n39502), .Z(n39403) );
  NAND U48631 ( .A(n39503), .B(n39504), .Z(n39502) );
  NAND U48632 ( .A(n39505), .B(n39506), .Z(n39501) );
  AND U48633 ( .A(n39507), .B(n39508), .Z(n39399) );
  NAND U48634 ( .A(n39509), .B(n39510), .Z(n39508) );
  NAND U48635 ( .A(n39511), .B(n39512), .Z(n39507) );
  AND U48636 ( .A(n39513), .B(n39514), .Z(n39401) );
  XOR U48637 ( .A(n39481), .B(n39480), .Z(N61879) );
  XNOR U48638 ( .A(n39498), .B(n39499), .Z(n39480) );
  XNOR U48639 ( .A(n39513), .B(n39514), .Z(n39499) );
  XOR U48640 ( .A(n39510), .B(n39509), .Z(n39514) );
  XOR U48641 ( .A(y[2388]), .B(x[2388]), .Z(n39509) );
  XOR U48642 ( .A(n39512), .B(n39511), .Z(n39510) );
  XOR U48643 ( .A(y[2390]), .B(x[2390]), .Z(n39511) );
  XOR U48644 ( .A(y[2389]), .B(x[2389]), .Z(n39512) );
  XOR U48645 ( .A(n39504), .B(n39503), .Z(n39513) );
  XOR U48646 ( .A(n39506), .B(n39505), .Z(n39503) );
  XOR U48647 ( .A(y[2387]), .B(x[2387]), .Z(n39505) );
  XOR U48648 ( .A(y[2386]), .B(x[2386]), .Z(n39506) );
  XOR U48649 ( .A(y[2385]), .B(x[2385]), .Z(n39504) );
  XNOR U48650 ( .A(n39497), .B(n39496), .Z(n39498) );
  XNOR U48651 ( .A(n39493), .B(n39492), .Z(n39496) );
  XOR U48652 ( .A(n39495), .B(n39494), .Z(n39492) );
  XOR U48653 ( .A(y[2384]), .B(x[2384]), .Z(n39494) );
  XOR U48654 ( .A(y[2383]), .B(x[2383]), .Z(n39495) );
  XOR U48655 ( .A(y[2382]), .B(x[2382]), .Z(n39493) );
  XOR U48656 ( .A(n39487), .B(n39486), .Z(n39497) );
  XOR U48657 ( .A(n39489), .B(n39488), .Z(n39486) );
  XOR U48658 ( .A(y[2381]), .B(x[2381]), .Z(n39488) );
  XOR U48659 ( .A(y[2380]), .B(x[2380]), .Z(n39489) );
  XOR U48660 ( .A(y[2379]), .B(x[2379]), .Z(n39487) );
  XNOR U48661 ( .A(n39463), .B(n39464), .Z(n39481) );
  XNOR U48662 ( .A(n39478), .B(n39479), .Z(n39464) );
  XOR U48663 ( .A(n39475), .B(n39474), .Z(n39479) );
  XOR U48664 ( .A(y[2376]), .B(x[2376]), .Z(n39474) );
  XOR U48665 ( .A(n39477), .B(n39476), .Z(n39475) );
  XOR U48666 ( .A(y[2378]), .B(x[2378]), .Z(n39476) );
  XOR U48667 ( .A(y[2377]), .B(x[2377]), .Z(n39477) );
  XOR U48668 ( .A(n39469), .B(n39468), .Z(n39478) );
  XOR U48669 ( .A(n39471), .B(n39470), .Z(n39468) );
  XOR U48670 ( .A(y[2375]), .B(x[2375]), .Z(n39470) );
  XOR U48671 ( .A(y[2374]), .B(x[2374]), .Z(n39471) );
  XOR U48672 ( .A(y[2373]), .B(x[2373]), .Z(n39469) );
  XNOR U48673 ( .A(n39462), .B(n39461), .Z(n39463) );
  XNOR U48674 ( .A(n39458), .B(n39457), .Z(n39461) );
  XOR U48675 ( .A(n39460), .B(n39459), .Z(n39457) );
  XOR U48676 ( .A(y[2372]), .B(x[2372]), .Z(n39459) );
  XOR U48677 ( .A(y[2371]), .B(x[2371]), .Z(n39460) );
  XOR U48678 ( .A(y[2370]), .B(x[2370]), .Z(n39458) );
  XOR U48679 ( .A(n39452), .B(n39451), .Z(n39462) );
  XOR U48680 ( .A(n39454), .B(n39453), .Z(n39451) );
  XOR U48681 ( .A(y[2369]), .B(x[2369]), .Z(n39453) );
  XOR U48682 ( .A(y[2368]), .B(x[2368]), .Z(n39454) );
  XOR U48683 ( .A(y[2367]), .B(x[2367]), .Z(n39452) );
  NAND U48684 ( .A(n39515), .B(n39516), .Z(N61870) );
  NAND U48685 ( .A(n39517), .B(n39518), .Z(n39516) );
  NANDN U48686 ( .A(n39519), .B(n39520), .Z(n39518) );
  NANDN U48687 ( .A(n39520), .B(n39519), .Z(n39515) );
  XOR U48688 ( .A(n39519), .B(n39521), .Z(N61869) );
  XNOR U48689 ( .A(n39517), .B(n39520), .Z(n39521) );
  NAND U48690 ( .A(n39522), .B(n39523), .Z(n39520) );
  NAND U48691 ( .A(n39524), .B(n39525), .Z(n39523) );
  NANDN U48692 ( .A(n39526), .B(n39527), .Z(n39525) );
  NANDN U48693 ( .A(n39527), .B(n39526), .Z(n39522) );
  AND U48694 ( .A(n39528), .B(n39529), .Z(n39517) );
  NAND U48695 ( .A(n39530), .B(n39531), .Z(n39529) );
  NANDN U48696 ( .A(n39532), .B(n39533), .Z(n39531) );
  NANDN U48697 ( .A(n39533), .B(n39532), .Z(n39528) );
  IV U48698 ( .A(n39534), .Z(n39533) );
  AND U48699 ( .A(n39535), .B(n39536), .Z(n39519) );
  NAND U48700 ( .A(n39537), .B(n39538), .Z(n39536) );
  NANDN U48701 ( .A(n39539), .B(n39540), .Z(n39538) );
  NANDN U48702 ( .A(n39540), .B(n39539), .Z(n39535) );
  XOR U48703 ( .A(n39532), .B(n39541), .Z(N61868) );
  XNOR U48704 ( .A(n39530), .B(n39534), .Z(n39541) );
  XOR U48705 ( .A(n39527), .B(n39542), .Z(n39534) );
  XNOR U48706 ( .A(n39524), .B(n39526), .Z(n39542) );
  AND U48707 ( .A(n39543), .B(n39544), .Z(n39526) );
  NANDN U48708 ( .A(n39545), .B(n39546), .Z(n39544) );
  OR U48709 ( .A(n39547), .B(n39548), .Z(n39546) );
  IV U48710 ( .A(n39549), .Z(n39548) );
  NANDN U48711 ( .A(n39549), .B(n39547), .Z(n39543) );
  AND U48712 ( .A(n39550), .B(n39551), .Z(n39524) );
  NAND U48713 ( .A(n39552), .B(n39553), .Z(n39551) );
  NANDN U48714 ( .A(n39554), .B(n39555), .Z(n39553) );
  NANDN U48715 ( .A(n39555), .B(n39554), .Z(n39550) );
  IV U48716 ( .A(n39556), .Z(n39555) );
  NAND U48717 ( .A(n39557), .B(n39558), .Z(n39527) );
  NANDN U48718 ( .A(n39559), .B(n39560), .Z(n39558) );
  NANDN U48719 ( .A(n39561), .B(n39562), .Z(n39560) );
  NANDN U48720 ( .A(n39562), .B(n39561), .Z(n39557) );
  IV U48721 ( .A(n39563), .Z(n39561) );
  AND U48722 ( .A(n39564), .B(n39565), .Z(n39530) );
  NAND U48723 ( .A(n39566), .B(n39567), .Z(n39565) );
  NANDN U48724 ( .A(n39568), .B(n39569), .Z(n39567) );
  NANDN U48725 ( .A(n39569), .B(n39568), .Z(n39564) );
  XOR U48726 ( .A(n39540), .B(n39570), .Z(n39532) );
  XNOR U48727 ( .A(n39537), .B(n39539), .Z(n39570) );
  AND U48728 ( .A(n39571), .B(n39572), .Z(n39539) );
  NANDN U48729 ( .A(n39573), .B(n39574), .Z(n39572) );
  OR U48730 ( .A(n39575), .B(n39576), .Z(n39574) );
  IV U48731 ( .A(n39577), .Z(n39576) );
  NANDN U48732 ( .A(n39577), .B(n39575), .Z(n39571) );
  AND U48733 ( .A(n39578), .B(n39579), .Z(n39537) );
  NAND U48734 ( .A(n39580), .B(n39581), .Z(n39579) );
  NANDN U48735 ( .A(n39582), .B(n39583), .Z(n39581) );
  NANDN U48736 ( .A(n39583), .B(n39582), .Z(n39578) );
  IV U48737 ( .A(n39584), .Z(n39583) );
  NAND U48738 ( .A(n39585), .B(n39586), .Z(n39540) );
  NANDN U48739 ( .A(n39587), .B(n39588), .Z(n39586) );
  NANDN U48740 ( .A(n39589), .B(n39590), .Z(n39588) );
  NANDN U48741 ( .A(n39590), .B(n39589), .Z(n39585) );
  IV U48742 ( .A(n39591), .Z(n39589) );
  XOR U48743 ( .A(n39566), .B(n39592), .Z(N61867) );
  XNOR U48744 ( .A(n39569), .B(n39568), .Z(n39592) );
  XNOR U48745 ( .A(n39580), .B(n39593), .Z(n39568) );
  XNOR U48746 ( .A(n39584), .B(n39582), .Z(n39593) );
  XOR U48747 ( .A(n39590), .B(n39594), .Z(n39582) );
  XNOR U48748 ( .A(n39587), .B(n39591), .Z(n39594) );
  AND U48749 ( .A(n39595), .B(n39596), .Z(n39591) );
  NAND U48750 ( .A(n39597), .B(n39598), .Z(n39596) );
  NAND U48751 ( .A(n39599), .B(n39600), .Z(n39595) );
  AND U48752 ( .A(n39601), .B(n39602), .Z(n39587) );
  NAND U48753 ( .A(n39603), .B(n39604), .Z(n39602) );
  NAND U48754 ( .A(n39605), .B(n39606), .Z(n39601) );
  NANDN U48755 ( .A(n39607), .B(n39608), .Z(n39590) );
  ANDN U48756 ( .B(n39609), .A(n39610), .Z(n39584) );
  XNOR U48757 ( .A(n39575), .B(n39611), .Z(n39580) );
  XNOR U48758 ( .A(n39573), .B(n39577), .Z(n39611) );
  AND U48759 ( .A(n39612), .B(n39613), .Z(n39577) );
  NAND U48760 ( .A(n39614), .B(n39615), .Z(n39613) );
  NAND U48761 ( .A(n39616), .B(n39617), .Z(n39612) );
  AND U48762 ( .A(n39618), .B(n39619), .Z(n39573) );
  NAND U48763 ( .A(n39620), .B(n39621), .Z(n39619) );
  NAND U48764 ( .A(n39622), .B(n39623), .Z(n39618) );
  AND U48765 ( .A(n39624), .B(n39625), .Z(n39575) );
  NAND U48766 ( .A(n39626), .B(n39627), .Z(n39569) );
  XNOR U48767 ( .A(n39552), .B(n39628), .Z(n39566) );
  XNOR U48768 ( .A(n39556), .B(n39554), .Z(n39628) );
  XOR U48769 ( .A(n39562), .B(n39629), .Z(n39554) );
  XNOR U48770 ( .A(n39559), .B(n39563), .Z(n39629) );
  AND U48771 ( .A(n39630), .B(n39631), .Z(n39563) );
  NAND U48772 ( .A(n39632), .B(n39633), .Z(n39631) );
  NAND U48773 ( .A(n39634), .B(n39635), .Z(n39630) );
  AND U48774 ( .A(n39636), .B(n39637), .Z(n39559) );
  NAND U48775 ( .A(n39638), .B(n39639), .Z(n39637) );
  NAND U48776 ( .A(n39640), .B(n39641), .Z(n39636) );
  NANDN U48777 ( .A(n39642), .B(n39643), .Z(n39562) );
  ANDN U48778 ( .B(n39644), .A(n39645), .Z(n39556) );
  XNOR U48779 ( .A(n39547), .B(n39646), .Z(n39552) );
  XNOR U48780 ( .A(n39545), .B(n39549), .Z(n39646) );
  AND U48781 ( .A(n39647), .B(n39648), .Z(n39549) );
  NAND U48782 ( .A(n39649), .B(n39650), .Z(n39648) );
  NAND U48783 ( .A(n39651), .B(n39652), .Z(n39647) );
  AND U48784 ( .A(n39653), .B(n39654), .Z(n39545) );
  NAND U48785 ( .A(n39655), .B(n39656), .Z(n39654) );
  NAND U48786 ( .A(n39657), .B(n39658), .Z(n39653) );
  AND U48787 ( .A(n39659), .B(n39660), .Z(n39547) );
  XOR U48788 ( .A(n39627), .B(n39626), .Z(N61866) );
  XNOR U48789 ( .A(n39644), .B(n39645), .Z(n39626) );
  XNOR U48790 ( .A(n39659), .B(n39660), .Z(n39645) );
  XOR U48791 ( .A(n39656), .B(n39655), .Z(n39660) );
  XOR U48792 ( .A(y[2364]), .B(x[2364]), .Z(n39655) );
  XOR U48793 ( .A(n39658), .B(n39657), .Z(n39656) );
  XOR U48794 ( .A(y[2366]), .B(x[2366]), .Z(n39657) );
  XOR U48795 ( .A(y[2365]), .B(x[2365]), .Z(n39658) );
  XOR U48796 ( .A(n39650), .B(n39649), .Z(n39659) );
  XOR U48797 ( .A(n39652), .B(n39651), .Z(n39649) );
  XOR U48798 ( .A(y[2363]), .B(x[2363]), .Z(n39651) );
  XOR U48799 ( .A(y[2362]), .B(x[2362]), .Z(n39652) );
  XOR U48800 ( .A(y[2361]), .B(x[2361]), .Z(n39650) );
  XNOR U48801 ( .A(n39643), .B(n39642), .Z(n39644) );
  XNOR U48802 ( .A(n39639), .B(n39638), .Z(n39642) );
  XOR U48803 ( .A(n39641), .B(n39640), .Z(n39638) );
  XOR U48804 ( .A(y[2360]), .B(x[2360]), .Z(n39640) );
  XOR U48805 ( .A(y[2359]), .B(x[2359]), .Z(n39641) );
  XOR U48806 ( .A(y[2358]), .B(x[2358]), .Z(n39639) );
  XOR U48807 ( .A(n39633), .B(n39632), .Z(n39643) );
  XOR U48808 ( .A(n39635), .B(n39634), .Z(n39632) );
  XOR U48809 ( .A(y[2357]), .B(x[2357]), .Z(n39634) );
  XOR U48810 ( .A(y[2356]), .B(x[2356]), .Z(n39635) );
  XOR U48811 ( .A(y[2355]), .B(x[2355]), .Z(n39633) );
  XNOR U48812 ( .A(n39609), .B(n39610), .Z(n39627) );
  XNOR U48813 ( .A(n39624), .B(n39625), .Z(n39610) );
  XOR U48814 ( .A(n39621), .B(n39620), .Z(n39625) );
  XOR U48815 ( .A(y[2352]), .B(x[2352]), .Z(n39620) );
  XOR U48816 ( .A(n39623), .B(n39622), .Z(n39621) );
  XOR U48817 ( .A(y[2354]), .B(x[2354]), .Z(n39622) );
  XOR U48818 ( .A(y[2353]), .B(x[2353]), .Z(n39623) );
  XOR U48819 ( .A(n39615), .B(n39614), .Z(n39624) );
  XOR U48820 ( .A(n39617), .B(n39616), .Z(n39614) );
  XOR U48821 ( .A(y[2351]), .B(x[2351]), .Z(n39616) );
  XOR U48822 ( .A(y[2350]), .B(x[2350]), .Z(n39617) );
  XOR U48823 ( .A(y[2349]), .B(x[2349]), .Z(n39615) );
  XNOR U48824 ( .A(n39608), .B(n39607), .Z(n39609) );
  XNOR U48825 ( .A(n39604), .B(n39603), .Z(n39607) );
  XOR U48826 ( .A(n39606), .B(n39605), .Z(n39603) );
  XOR U48827 ( .A(y[2348]), .B(x[2348]), .Z(n39605) );
  XOR U48828 ( .A(y[2347]), .B(x[2347]), .Z(n39606) );
  XOR U48829 ( .A(y[2346]), .B(x[2346]), .Z(n39604) );
  XOR U48830 ( .A(n39598), .B(n39597), .Z(n39608) );
  XOR U48831 ( .A(n39600), .B(n39599), .Z(n39597) );
  XOR U48832 ( .A(y[2345]), .B(x[2345]), .Z(n39599) );
  XOR U48833 ( .A(y[2344]), .B(x[2344]), .Z(n39600) );
  XOR U48834 ( .A(y[2343]), .B(x[2343]), .Z(n39598) );
  NAND U48835 ( .A(n39661), .B(n39662), .Z(N61857) );
  NAND U48836 ( .A(n39663), .B(n39664), .Z(n39662) );
  NANDN U48837 ( .A(n39665), .B(n39666), .Z(n39664) );
  NANDN U48838 ( .A(n39666), .B(n39665), .Z(n39661) );
  XOR U48839 ( .A(n39665), .B(n39667), .Z(N61856) );
  XNOR U48840 ( .A(n39663), .B(n39666), .Z(n39667) );
  NAND U48841 ( .A(n39668), .B(n39669), .Z(n39666) );
  NAND U48842 ( .A(n39670), .B(n39671), .Z(n39669) );
  NANDN U48843 ( .A(n39672), .B(n39673), .Z(n39671) );
  NANDN U48844 ( .A(n39673), .B(n39672), .Z(n39668) );
  AND U48845 ( .A(n39674), .B(n39675), .Z(n39663) );
  NAND U48846 ( .A(n39676), .B(n39677), .Z(n39675) );
  NANDN U48847 ( .A(n39678), .B(n39679), .Z(n39677) );
  NANDN U48848 ( .A(n39679), .B(n39678), .Z(n39674) );
  IV U48849 ( .A(n39680), .Z(n39679) );
  AND U48850 ( .A(n39681), .B(n39682), .Z(n39665) );
  NAND U48851 ( .A(n39683), .B(n39684), .Z(n39682) );
  NANDN U48852 ( .A(n39685), .B(n39686), .Z(n39684) );
  NANDN U48853 ( .A(n39686), .B(n39685), .Z(n39681) );
  XOR U48854 ( .A(n39678), .B(n39687), .Z(N61855) );
  XNOR U48855 ( .A(n39676), .B(n39680), .Z(n39687) );
  XOR U48856 ( .A(n39673), .B(n39688), .Z(n39680) );
  XNOR U48857 ( .A(n39670), .B(n39672), .Z(n39688) );
  AND U48858 ( .A(n39689), .B(n39690), .Z(n39672) );
  NANDN U48859 ( .A(n39691), .B(n39692), .Z(n39690) );
  OR U48860 ( .A(n39693), .B(n39694), .Z(n39692) );
  IV U48861 ( .A(n39695), .Z(n39694) );
  NANDN U48862 ( .A(n39695), .B(n39693), .Z(n39689) );
  AND U48863 ( .A(n39696), .B(n39697), .Z(n39670) );
  NAND U48864 ( .A(n39698), .B(n39699), .Z(n39697) );
  NANDN U48865 ( .A(n39700), .B(n39701), .Z(n39699) );
  NANDN U48866 ( .A(n39701), .B(n39700), .Z(n39696) );
  IV U48867 ( .A(n39702), .Z(n39701) );
  NAND U48868 ( .A(n39703), .B(n39704), .Z(n39673) );
  NANDN U48869 ( .A(n39705), .B(n39706), .Z(n39704) );
  NANDN U48870 ( .A(n39707), .B(n39708), .Z(n39706) );
  NANDN U48871 ( .A(n39708), .B(n39707), .Z(n39703) );
  IV U48872 ( .A(n39709), .Z(n39707) );
  AND U48873 ( .A(n39710), .B(n39711), .Z(n39676) );
  NAND U48874 ( .A(n39712), .B(n39713), .Z(n39711) );
  NANDN U48875 ( .A(n39714), .B(n39715), .Z(n39713) );
  NANDN U48876 ( .A(n39715), .B(n39714), .Z(n39710) );
  XOR U48877 ( .A(n39686), .B(n39716), .Z(n39678) );
  XNOR U48878 ( .A(n39683), .B(n39685), .Z(n39716) );
  AND U48879 ( .A(n39717), .B(n39718), .Z(n39685) );
  NANDN U48880 ( .A(n39719), .B(n39720), .Z(n39718) );
  OR U48881 ( .A(n39721), .B(n39722), .Z(n39720) );
  IV U48882 ( .A(n39723), .Z(n39722) );
  NANDN U48883 ( .A(n39723), .B(n39721), .Z(n39717) );
  AND U48884 ( .A(n39724), .B(n39725), .Z(n39683) );
  NAND U48885 ( .A(n39726), .B(n39727), .Z(n39725) );
  NANDN U48886 ( .A(n39728), .B(n39729), .Z(n39727) );
  NANDN U48887 ( .A(n39729), .B(n39728), .Z(n39724) );
  IV U48888 ( .A(n39730), .Z(n39729) );
  NAND U48889 ( .A(n39731), .B(n39732), .Z(n39686) );
  NANDN U48890 ( .A(n39733), .B(n39734), .Z(n39732) );
  NANDN U48891 ( .A(n39735), .B(n39736), .Z(n39734) );
  NANDN U48892 ( .A(n39736), .B(n39735), .Z(n39731) );
  IV U48893 ( .A(n39737), .Z(n39735) );
  XOR U48894 ( .A(n39712), .B(n39738), .Z(N61854) );
  XNOR U48895 ( .A(n39715), .B(n39714), .Z(n39738) );
  XNOR U48896 ( .A(n39726), .B(n39739), .Z(n39714) );
  XNOR U48897 ( .A(n39730), .B(n39728), .Z(n39739) );
  XOR U48898 ( .A(n39736), .B(n39740), .Z(n39728) );
  XNOR U48899 ( .A(n39733), .B(n39737), .Z(n39740) );
  AND U48900 ( .A(n39741), .B(n39742), .Z(n39737) );
  NAND U48901 ( .A(n39743), .B(n39744), .Z(n39742) );
  NAND U48902 ( .A(n39745), .B(n39746), .Z(n39741) );
  AND U48903 ( .A(n39747), .B(n39748), .Z(n39733) );
  NAND U48904 ( .A(n39749), .B(n39750), .Z(n39748) );
  NAND U48905 ( .A(n39751), .B(n39752), .Z(n39747) );
  NANDN U48906 ( .A(n39753), .B(n39754), .Z(n39736) );
  ANDN U48907 ( .B(n39755), .A(n39756), .Z(n39730) );
  XNOR U48908 ( .A(n39721), .B(n39757), .Z(n39726) );
  XNOR U48909 ( .A(n39719), .B(n39723), .Z(n39757) );
  AND U48910 ( .A(n39758), .B(n39759), .Z(n39723) );
  NAND U48911 ( .A(n39760), .B(n39761), .Z(n39759) );
  NAND U48912 ( .A(n39762), .B(n39763), .Z(n39758) );
  AND U48913 ( .A(n39764), .B(n39765), .Z(n39719) );
  NAND U48914 ( .A(n39766), .B(n39767), .Z(n39765) );
  NAND U48915 ( .A(n39768), .B(n39769), .Z(n39764) );
  AND U48916 ( .A(n39770), .B(n39771), .Z(n39721) );
  NAND U48917 ( .A(n39772), .B(n39773), .Z(n39715) );
  XNOR U48918 ( .A(n39698), .B(n39774), .Z(n39712) );
  XNOR U48919 ( .A(n39702), .B(n39700), .Z(n39774) );
  XOR U48920 ( .A(n39708), .B(n39775), .Z(n39700) );
  XNOR U48921 ( .A(n39705), .B(n39709), .Z(n39775) );
  AND U48922 ( .A(n39776), .B(n39777), .Z(n39709) );
  NAND U48923 ( .A(n39778), .B(n39779), .Z(n39777) );
  NAND U48924 ( .A(n39780), .B(n39781), .Z(n39776) );
  AND U48925 ( .A(n39782), .B(n39783), .Z(n39705) );
  NAND U48926 ( .A(n39784), .B(n39785), .Z(n39783) );
  NAND U48927 ( .A(n39786), .B(n39787), .Z(n39782) );
  NANDN U48928 ( .A(n39788), .B(n39789), .Z(n39708) );
  ANDN U48929 ( .B(n39790), .A(n39791), .Z(n39702) );
  XNOR U48930 ( .A(n39693), .B(n39792), .Z(n39698) );
  XNOR U48931 ( .A(n39691), .B(n39695), .Z(n39792) );
  AND U48932 ( .A(n39793), .B(n39794), .Z(n39695) );
  NAND U48933 ( .A(n39795), .B(n39796), .Z(n39794) );
  NAND U48934 ( .A(n39797), .B(n39798), .Z(n39793) );
  AND U48935 ( .A(n39799), .B(n39800), .Z(n39691) );
  NAND U48936 ( .A(n39801), .B(n39802), .Z(n39800) );
  NAND U48937 ( .A(n39803), .B(n39804), .Z(n39799) );
  AND U48938 ( .A(n39805), .B(n39806), .Z(n39693) );
  XOR U48939 ( .A(n39773), .B(n39772), .Z(N61853) );
  XNOR U48940 ( .A(n39790), .B(n39791), .Z(n39772) );
  XNOR U48941 ( .A(n39805), .B(n39806), .Z(n39791) );
  XOR U48942 ( .A(n39802), .B(n39801), .Z(n39806) );
  XOR U48943 ( .A(y[2340]), .B(x[2340]), .Z(n39801) );
  XOR U48944 ( .A(n39804), .B(n39803), .Z(n39802) );
  XOR U48945 ( .A(y[2342]), .B(x[2342]), .Z(n39803) );
  XOR U48946 ( .A(y[2341]), .B(x[2341]), .Z(n39804) );
  XOR U48947 ( .A(n39796), .B(n39795), .Z(n39805) );
  XOR U48948 ( .A(n39798), .B(n39797), .Z(n39795) );
  XOR U48949 ( .A(y[2339]), .B(x[2339]), .Z(n39797) );
  XOR U48950 ( .A(y[2338]), .B(x[2338]), .Z(n39798) );
  XOR U48951 ( .A(y[2337]), .B(x[2337]), .Z(n39796) );
  XNOR U48952 ( .A(n39789), .B(n39788), .Z(n39790) );
  XNOR U48953 ( .A(n39785), .B(n39784), .Z(n39788) );
  XOR U48954 ( .A(n39787), .B(n39786), .Z(n39784) );
  XOR U48955 ( .A(y[2336]), .B(x[2336]), .Z(n39786) );
  XOR U48956 ( .A(y[2335]), .B(x[2335]), .Z(n39787) );
  XOR U48957 ( .A(y[2334]), .B(x[2334]), .Z(n39785) );
  XOR U48958 ( .A(n39779), .B(n39778), .Z(n39789) );
  XOR U48959 ( .A(n39781), .B(n39780), .Z(n39778) );
  XOR U48960 ( .A(y[2333]), .B(x[2333]), .Z(n39780) );
  XOR U48961 ( .A(y[2332]), .B(x[2332]), .Z(n39781) );
  XOR U48962 ( .A(y[2331]), .B(x[2331]), .Z(n39779) );
  XNOR U48963 ( .A(n39755), .B(n39756), .Z(n39773) );
  XNOR U48964 ( .A(n39770), .B(n39771), .Z(n39756) );
  XOR U48965 ( .A(n39767), .B(n39766), .Z(n39771) );
  XOR U48966 ( .A(y[2328]), .B(x[2328]), .Z(n39766) );
  XOR U48967 ( .A(n39769), .B(n39768), .Z(n39767) );
  XOR U48968 ( .A(y[2330]), .B(x[2330]), .Z(n39768) );
  XOR U48969 ( .A(y[2329]), .B(x[2329]), .Z(n39769) );
  XOR U48970 ( .A(n39761), .B(n39760), .Z(n39770) );
  XOR U48971 ( .A(n39763), .B(n39762), .Z(n39760) );
  XOR U48972 ( .A(y[2327]), .B(x[2327]), .Z(n39762) );
  XOR U48973 ( .A(y[2326]), .B(x[2326]), .Z(n39763) );
  XOR U48974 ( .A(y[2325]), .B(x[2325]), .Z(n39761) );
  XNOR U48975 ( .A(n39754), .B(n39753), .Z(n39755) );
  XNOR U48976 ( .A(n39750), .B(n39749), .Z(n39753) );
  XOR U48977 ( .A(n39752), .B(n39751), .Z(n39749) );
  XOR U48978 ( .A(y[2324]), .B(x[2324]), .Z(n39751) );
  XOR U48979 ( .A(y[2323]), .B(x[2323]), .Z(n39752) );
  XOR U48980 ( .A(y[2322]), .B(x[2322]), .Z(n39750) );
  XOR U48981 ( .A(n39744), .B(n39743), .Z(n39754) );
  XOR U48982 ( .A(n39746), .B(n39745), .Z(n39743) );
  XOR U48983 ( .A(y[2321]), .B(x[2321]), .Z(n39745) );
  XOR U48984 ( .A(y[2320]), .B(x[2320]), .Z(n39746) );
  XOR U48985 ( .A(y[2319]), .B(x[2319]), .Z(n39744) );
  NAND U48986 ( .A(n39807), .B(n39808), .Z(N61844) );
  NAND U48987 ( .A(n39809), .B(n39810), .Z(n39808) );
  NANDN U48988 ( .A(n39811), .B(n39812), .Z(n39810) );
  NANDN U48989 ( .A(n39812), .B(n39811), .Z(n39807) );
  XOR U48990 ( .A(n39811), .B(n39813), .Z(N61843) );
  XNOR U48991 ( .A(n39809), .B(n39812), .Z(n39813) );
  NAND U48992 ( .A(n39814), .B(n39815), .Z(n39812) );
  NAND U48993 ( .A(n39816), .B(n39817), .Z(n39815) );
  NANDN U48994 ( .A(n39818), .B(n39819), .Z(n39817) );
  NANDN U48995 ( .A(n39819), .B(n39818), .Z(n39814) );
  AND U48996 ( .A(n39820), .B(n39821), .Z(n39809) );
  NAND U48997 ( .A(n39822), .B(n39823), .Z(n39821) );
  NANDN U48998 ( .A(n39824), .B(n39825), .Z(n39823) );
  NANDN U48999 ( .A(n39825), .B(n39824), .Z(n39820) );
  IV U49000 ( .A(n39826), .Z(n39825) );
  AND U49001 ( .A(n39827), .B(n39828), .Z(n39811) );
  NAND U49002 ( .A(n39829), .B(n39830), .Z(n39828) );
  NANDN U49003 ( .A(n39831), .B(n39832), .Z(n39830) );
  NANDN U49004 ( .A(n39832), .B(n39831), .Z(n39827) );
  XOR U49005 ( .A(n39824), .B(n39833), .Z(N61842) );
  XNOR U49006 ( .A(n39822), .B(n39826), .Z(n39833) );
  XOR U49007 ( .A(n39819), .B(n39834), .Z(n39826) );
  XNOR U49008 ( .A(n39816), .B(n39818), .Z(n39834) );
  AND U49009 ( .A(n39835), .B(n39836), .Z(n39818) );
  NANDN U49010 ( .A(n39837), .B(n39838), .Z(n39836) );
  OR U49011 ( .A(n39839), .B(n39840), .Z(n39838) );
  IV U49012 ( .A(n39841), .Z(n39840) );
  NANDN U49013 ( .A(n39841), .B(n39839), .Z(n39835) );
  AND U49014 ( .A(n39842), .B(n39843), .Z(n39816) );
  NAND U49015 ( .A(n39844), .B(n39845), .Z(n39843) );
  NANDN U49016 ( .A(n39846), .B(n39847), .Z(n39845) );
  NANDN U49017 ( .A(n39847), .B(n39846), .Z(n39842) );
  IV U49018 ( .A(n39848), .Z(n39847) );
  NAND U49019 ( .A(n39849), .B(n39850), .Z(n39819) );
  NANDN U49020 ( .A(n39851), .B(n39852), .Z(n39850) );
  NANDN U49021 ( .A(n39853), .B(n39854), .Z(n39852) );
  NANDN U49022 ( .A(n39854), .B(n39853), .Z(n39849) );
  IV U49023 ( .A(n39855), .Z(n39853) );
  AND U49024 ( .A(n39856), .B(n39857), .Z(n39822) );
  NAND U49025 ( .A(n39858), .B(n39859), .Z(n39857) );
  NANDN U49026 ( .A(n39860), .B(n39861), .Z(n39859) );
  NANDN U49027 ( .A(n39861), .B(n39860), .Z(n39856) );
  XOR U49028 ( .A(n39832), .B(n39862), .Z(n39824) );
  XNOR U49029 ( .A(n39829), .B(n39831), .Z(n39862) );
  AND U49030 ( .A(n39863), .B(n39864), .Z(n39831) );
  NANDN U49031 ( .A(n39865), .B(n39866), .Z(n39864) );
  OR U49032 ( .A(n39867), .B(n39868), .Z(n39866) );
  IV U49033 ( .A(n39869), .Z(n39868) );
  NANDN U49034 ( .A(n39869), .B(n39867), .Z(n39863) );
  AND U49035 ( .A(n39870), .B(n39871), .Z(n39829) );
  NAND U49036 ( .A(n39872), .B(n39873), .Z(n39871) );
  NANDN U49037 ( .A(n39874), .B(n39875), .Z(n39873) );
  NANDN U49038 ( .A(n39875), .B(n39874), .Z(n39870) );
  IV U49039 ( .A(n39876), .Z(n39875) );
  NAND U49040 ( .A(n39877), .B(n39878), .Z(n39832) );
  NANDN U49041 ( .A(n39879), .B(n39880), .Z(n39878) );
  NANDN U49042 ( .A(n39881), .B(n39882), .Z(n39880) );
  NANDN U49043 ( .A(n39882), .B(n39881), .Z(n39877) );
  IV U49044 ( .A(n39883), .Z(n39881) );
  XOR U49045 ( .A(n39858), .B(n39884), .Z(N61841) );
  XNOR U49046 ( .A(n39861), .B(n39860), .Z(n39884) );
  XNOR U49047 ( .A(n39872), .B(n39885), .Z(n39860) );
  XNOR U49048 ( .A(n39876), .B(n39874), .Z(n39885) );
  XOR U49049 ( .A(n39882), .B(n39886), .Z(n39874) );
  XNOR U49050 ( .A(n39879), .B(n39883), .Z(n39886) );
  AND U49051 ( .A(n39887), .B(n39888), .Z(n39883) );
  NAND U49052 ( .A(n39889), .B(n39890), .Z(n39888) );
  NAND U49053 ( .A(n39891), .B(n39892), .Z(n39887) );
  AND U49054 ( .A(n39893), .B(n39894), .Z(n39879) );
  NAND U49055 ( .A(n39895), .B(n39896), .Z(n39894) );
  NAND U49056 ( .A(n39897), .B(n39898), .Z(n39893) );
  NANDN U49057 ( .A(n39899), .B(n39900), .Z(n39882) );
  ANDN U49058 ( .B(n39901), .A(n39902), .Z(n39876) );
  XNOR U49059 ( .A(n39867), .B(n39903), .Z(n39872) );
  XNOR U49060 ( .A(n39865), .B(n39869), .Z(n39903) );
  AND U49061 ( .A(n39904), .B(n39905), .Z(n39869) );
  NAND U49062 ( .A(n39906), .B(n39907), .Z(n39905) );
  NAND U49063 ( .A(n39908), .B(n39909), .Z(n39904) );
  AND U49064 ( .A(n39910), .B(n39911), .Z(n39865) );
  NAND U49065 ( .A(n39912), .B(n39913), .Z(n39911) );
  NAND U49066 ( .A(n39914), .B(n39915), .Z(n39910) );
  AND U49067 ( .A(n39916), .B(n39917), .Z(n39867) );
  NAND U49068 ( .A(n39918), .B(n39919), .Z(n39861) );
  XNOR U49069 ( .A(n39844), .B(n39920), .Z(n39858) );
  XNOR U49070 ( .A(n39848), .B(n39846), .Z(n39920) );
  XOR U49071 ( .A(n39854), .B(n39921), .Z(n39846) );
  XNOR U49072 ( .A(n39851), .B(n39855), .Z(n39921) );
  AND U49073 ( .A(n39922), .B(n39923), .Z(n39855) );
  NAND U49074 ( .A(n39924), .B(n39925), .Z(n39923) );
  NAND U49075 ( .A(n39926), .B(n39927), .Z(n39922) );
  AND U49076 ( .A(n39928), .B(n39929), .Z(n39851) );
  NAND U49077 ( .A(n39930), .B(n39931), .Z(n39929) );
  NAND U49078 ( .A(n39932), .B(n39933), .Z(n39928) );
  NANDN U49079 ( .A(n39934), .B(n39935), .Z(n39854) );
  ANDN U49080 ( .B(n39936), .A(n39937), .Z(n39848) );
  XNOR U49081 ( .A(n39839), .B(n39938), .Z(n39844) );
  XNOR U49082 ( .A(n39837), .B(n39841), .Z(n39938) );
  AND U49083 ( .A(n39939), .B(n39940), .Z(n39841) );
  NAND U49084 ( .A(n39941), .B(n39942), .Z(n39940) );
  NAND U49085 ( .A(n39943), .B(n39944), .Z(n39939) );
  AND U49086 ( .A(n39945), .B(n39946), .Z(n39837) );
  NAND U49087 ( .A(n39947), .B(n39948), .Z(n39946) );
  NAND U49088 ( .A(n39949), .B(n39950), .Z(n39945) );
  AND U49089 ( .A(n39951), .B(n39952), .Z(n39839) );
  XOR U49090 ( .A(n39919), .B(n39918), .Z(N61840) );
  XNOR U49091 ( .A(n39936), .B(n39937), .Z(n39918) );
  XNOR U49092 ( .A(n39951), .B(n39952), .Z(n39937) );
  XOR U49093 ( .A(n39948), .B(n39947), .Z(n39952) );
  XOR U49094 ( .A(y[2316]), .B(x[2316]), .Z(n39947) );
  XOR U49095 ( .A(n39950), .B(n39949), .Z(n39948) );
  XOR U49096 ( .A(y[2318]), .B(x[2318]), .Z(n39949) );
  XOR U49097 ( .A(y[2317]), .B(x[2317]), .Z(n39950) );
  XOR U49098 ( .A(n39942), .B(n39941), .Z(n39951) );
  XOR U49099 ( .A(n39944), .B(n39943), .Z(n39941) );
  XOR U49100 ( .A(y[2315]), .B(x[2315]), .Z(n39943) );
  XOR U49101 ( .A(y[2314]), .B(x[2314]), .Z(n39944) );
  XOR U49102 ( .A(y[2313]), .B(x[2313]), .Z(n39942) );
  XNOR U49103 ( .A(n39935), .B(n39934), .Z(n39936) );
  XNOR U49104 ( .A(n39931), .B(n39930), .Z(n39934) );
  XOR U49105 ( .A(n39933), .B(n39932), .Z(n39930) );
  XOR U49106 ( .A(y[2312]), .B(x[2312]), .Z(n39932) );
  XOR U49107 ( .A(y[2311]), .B(x[2311]), .Z(n39933) );
  XOR U49108 ( .A(y[2310]), .B(x[2310]), .Z(n39931) );
  XOR U49109 ( .A(n39925), .B(n39924), .Z(n39935) );
  XOR U49110 ( .A(n39927), .B(n39926), .Z(n39924) );
  XOR U49111 ( .A(y[2309]), .B(x[2309]), .Z(n39926) );
  XOR U49112 ( .A(y[2308]), .B(x[2308]), .Z(n39927) );
  XOR U49113 ( .A(y[2307]), .B(x[2307]), .Z(n39925) );
  XNOR U49114 ( .A(n39901), .B(n39902), .Z(n39919) );
  XNOR U49115 ( .A(n39916), .B(n39917), .Z(n39902) );
  XOR U49116 ( .A(n39913), .B(n39912), .Z(n39917) );
  XOR U49117 ( .A(y[2304]), .B(x[2304]), .Z(n39912) );
  XOR U49118 ( .A(n39915), .B(n39914), .Z(n39913) );
  XOR U49119 ( .A(y[2306]), .B(x[2306]), .Z(n39914) );
  XOR U49120 ( .A(y[2305]), .B(x[2305]), .Z(n39915) );
  XOR U49121 ( .A(n39907), .B(n39906), .Z(n39916) );
  XOR U49122 ( .A(n39909), .B(n39908), .Z(n39906) );
  XOR U49123 ( .A(y[2303]), .B(x[2303]), .Z(n39908) );
  XOR U49124 ( .A(y[2302]), .B(x[2302]), .Z(n39909) );
  XOR U49125 ( .A(y[2301]), .B(x[2301]), .Z(n39907) );
  XNOR U49126 ( .A(n39900), .B(n39899), .Z(n39901) );
  XNOR U49127 ( .A(n39896), .B(n39895), .Z(n39899) );
  XOR U49128 ( .A(n39898), .B(n39897), .Z(n39895) );
  XOR U49129 ( .A(y[2300]), .B(x[2300]), .Z(n39897) );
  XOR U49130 ( .A(y[2299]), .B(x[2299]), .Z(n39898) );
  XOR U49131 ( .A(y[2298]), .B(x[2298]), .Z(n39896) );
  XOR U49132 ( .A(n39890), .B(n39889), .Z(n39900) );
  XOR U49133 ( .A(n39892), .B(n39891), .Z(n39889) );
  XOR U49134 ( .A(y[2297]), .B(x[2297]), .Z(n39891) );
  XOR U49135 ( .A(y[2296]), .B(x[2296]), .Z(n39892) );
  XOR U49136 ( .A(y[2295]), .B(x[2295]), .Z(n39890) );
  NAND U49137 ( .A(n39953), .B(n39954), .Z(N61831) );
  NAND U49138 ( .A(n39955), .B(n39956), .Z(n39954) );
  NANDN U49139 ( .A(n39957), .B(n39958), .Z(n39956) );
  NANDN U49140 ( .A(n39958), .B(n39957), .Z(n39953) );
  XOR U49141 ( .A(n39957), .B(n39959), .Z(N61830) );
  XNOR U49142 ( .A(n39955), .B(n39958), .Z(n39959) );
  NAND U49143 ( .A(n39960), .B(n39961), .Z(n39958) );
  NAND U49144 ( .A(n39962), .B(n39963), .Z(n39961) );
  NANDN U49145 ( .A(n39964), .B(n39965), .Z(n39963) );
  NANDN U49146 ( .A(n39965), .B(n39964), .Z(n39960) );
  AND U49147 ( .A(n39966), .B(n39967), .Z(n39955) );
  NAND U49148 ( .A(n39968), .B(n39969), .Z(n39967) );
  NANDN U49149 ( .A(n39970), .B(n39971), .Z(n39969) );
  NANDN U49150 ( .A(n39971), .B(n39970), .Z(n39966) );
  IV U49151 ( .A(n39972), .Z(n39971) );
  AND U49152 ( .A(n39973), .B(n39974), .Z(n39957) );
  NAND U49153 ( .A(n39975), .B(n39976), .Z(n39974) );
  NANDN U49154 ( .A(n39977), .B(n39978), .Z(n39976) );
  NANDN U49155 ( .A(n39978), .B(n39977), .Z(n39973) );
  XOR U49156 ( .A(n39970), .B(n39979), .Z(N61829) );
  XNOR U49157 ( .A(n39968), .B(n39972), .Z(n39979) );
  XOR U49158 ( .A(n39965), .B(n39980), .Z(n39972) );
  XNOR U49159 ( .A(n39962), .B(n39964), .Z(n39980) );
  AND U49160 ( .A(n39981), .B(n39982), .Z(n39964) );
  NANDN U49161 ( .A(n39983), .B(n39984), .Z(n39982) );
  OR U49162 ( .A(n39985), .B(n39986), .Z(n39984) );
  IV U49163 ( .A(n39987), .Z(n39986) );
  NANDN U49164 ( .A(n39987), .B(n39985), .Z(n39981) );
  AND U49165 ( .A(n39988), .B(n39989), .Z(n39962) );
  NAND U49166 ( .A(n39990), .B(n39991), .Z(n39989) );
  NANDN U49167 ( .A(n39992), .B(n39993), .Z(n39991) );
  NANDN U49168 ( .A(n39993), .B(n39992), .Z(n39988) );
  IV U49169 ( .A(n39994), .Z(n39993) );
  NAND U49170 ( .A(n39995), .B(n39996), .Z(n39965) );
  NANDN U49171 ( .A(n39997), .B(n39998), .Z(n39996) );
  NANDN U49172 ( .A(n39999), .B(n40000), .Z(n39998) );
  NANDN U49173 ( .A(n40000), .B(n39999), .Z(n39995) );
  IV U49174 ( .A(n40001), .Z(n39999) );
  AND U49175 ( .A(n40002), .B(n40003), .Z(n39968) );
  NAND U49176 ( .A(n40004), .B(n40005), .Z(n40003) );
  NANDN U49177 ( .A(n40006), .B(n40007), .Z(n40005) );
  NANDN U49178 ( .A(n40007), .B(n40006), .Z(n40002) );
  XOR U49179 ( .A(n39978), .B(n40008), .Z(n39970) );
  XNOR U49180 ( .A(n39975), .B(n39977), .Z(n40008) );
  AND U49181 ( .A(n40009), .B(n40010), .Z(n39977) );
  NANDN U49182 ( .A(n40011), .B(n40012), .Z(n40010) );
  OR U49183 ( .A(n40013), .B(n40014), .Z(n40012) );
  IV U49184 ( .A(n40015), .Z(n40014) );
  NANDN U49185 ( .A(n40015), .B(n40013), .Z(n40009) );
  AND U49186 ( .A(n40016), .B(n40017), .Z(n39975) );
  NAND U49187 ( .A(n40018), .B(n40019), .Z(n40017) );
  NANDN U49188 ( .A(n40020), .B(n40021), .Z(n40019) );
  NANDN U49189 ( .A(n40021), .B(n40020), .Z(n40016) );
  IV U49190 ( .A(n40022), .Z(n40021) );
  NAND U49191 ( .A(n40023), .B(n40024), .Z(n39978) );
  NANDN U49192 ( .A(n40025), .B(n40026), .Z(n40024) );
  NANDN U49193 ( .A(n40027), .B(n40028), .Z(n40026) );
  NANDN U49194 ( .A(n40028), .B(n40027), .Z(n40023) );
  IV U49195 ( .A(n40029), .Z(n40027) );
  XOR U49196 ( .A(n40004), .B(n40030), .Z(N61828) );
  XNOR U49197 ( .A(n40007), .B(n40006), .Z(n40030) );
  XNOR U49198 ( .A(n40018), .B(n40031), .Z(n40006) );
  XNOR U49199 ( .A(n40022), .B(n40020), .Z(n40031) );
  XOR U49200 ( .A(n40028), .B(n40032), .Z(n40020) );
  XNOR U49201 ( .A(n40025), .B(n40029), .Z(n40032) );
  AND U49202 ( .A(n40033), .B(n40034), .Z(n40029) );
  NAND U49203 ( .A(n40035), .B(n40036), .Z(n40034) );
  NAND U49204 ( .A(n40037), .B(n40038), .Z(n40033) );
  AND U49205 ( .A(n40039), .B(n40040), .Z(n40025) );
  NAND U49206 ( .A(n40041), .B(n40042), .Z(n40040) );
  NAND U49207 ( .A(n40043), .B(n40044), .Z(n40039) );
  NANDN U49208 ( .A(n40045), .B(n40046), .Z(n40028) );
  ANDN U49209 ( .B(n40047), .A(n40048), .Z(n40022) );
  XNOR U49210 ( .A(n40013), .B(n40049), .Z(n40018) );
  XNOR U49211 ( .A(n40011), .B(n40015), .Z(n40049) );
  AND U49212 ( .A(n40050), .B(n40051), .Z(n40015) );
  NAND U49213 ( .A(n40052), .B(n40053), .Z(n40051) );
  NAND U49214 ( .A(n40054), .B(n40055), .Z(n40050) );
  AND U49215 ( .A(n40056), .B(n40057), .Z(n40011) );
  NAND U49216 ( .A(n40058), .B(n40059), .Z(n40057) );
  NAND U49217 ( .A(n40060), .B(n40061), .Z(n40056) );
  AND U49218 ( .A(n40062), .B(n40063), .Z(n40013) );
  NAND U49219 ( .A(n40064), .B(n40065), .Z(n40007) );
  XNOR U49220 ( .A(n39990), .B(n40066), .Z(n40004) );
  XNOR U49221 ( .A(n39994), .B(n39992), .Z(n40066) );
  XOR U49222 ( .A(n40000), .B(n40067), .Z(n39992) );
  XNOR U49223 ( .A(n39997), .B(n40001), .Z(n40067) );
  AND U49224 ( .A(n40068), .B(n40069), .Z(n40001) );
  NAND U49225 ( .A(n40070), .B(n40071), .Z(n40069) );
  NAND U49226 ( .A(n40072), .B(n40073), .Z(n40068) );
  AND U49227 ( .A(n40074), .B(n40075), .Z(n39997) );
  NAND U49228 ( .A(n40076), .B(n40077), .Z(n40075) );
  NAND U49229 ( .A(n40078), .B(n40079), .Z(n40074) );
  NANDN U49230 ( .A(n40080), .B(n40081), .Z(n40000) );
  ANDN U49231 ( .B(n40082), .A(n40083), .Z(n39994) );
  XNOR U49232 ( .A(n39985), .B(n40084), .Z(n39990) );
  XNOR U49233 ( .A(n39983), .B(n39987), .Z(n40084) );
  AND U49234 ( .A(n40085), .B(n40086), .Z(n39987) );
  NAND U49235 ( .A(n40087), .B(n40088), .Z(n40086) );
  NAND U49236 ( .A(n40089), .B(n40090), .Z(n40085) );
  AND U49237 ( .A(n40091), .B(n40092), .Z(n39983) );
  NAND U49238 ( .A(n40093), .B(n40094), .Z(n40092) );
  NAND U49239 ( .A(n40095), .B(n40096), .Z(n40091) );
  AND U49240 ( .A(n40097), .B(n40098), .Z(n39985) );
  XOR U49241 ( .A(n40065), .B(n40064), .Z(N61827) );
  XNOR U49242 ( .A(n40082), .B(n40083), .Z(n40064) );
  XNOR U49243 ( .A(n40097), .B(n40098), .Z(n40083) );
  XOR U49244 ( .A(n40094), .B(n40093), .Z(n40098) );
  XOR U49245 ( .A(y[2292]), .B(x[2292]), .Z(n40093) );
  XOR U49246 ( .A(n40096), .B(n40095), .Z(n40094) );
  XOR U49247 ( .A(y[2294]), .B(x[2294]), .Z(n40095) );
  XOR U49248 ( .A(y[2293]), .B(x[2293]), .Z(n40096) );
  XOR U49249 ( .A(n40088), .B(n40087), .Z(n40097) );
  XOR U49250 ( .A(n40090), .B(n40089), .Z(n40087) );
  XOR U49251 ( .A(y[2291]), .B(x[2291]), .Z(n40089) );
  XOR U49252 ( .A(y[2290]), .B(x[2290]), .Z(n40090) );
  XOR U49253 ( .A(y[2289]), .B(x[2289]), .Z(n40088) );
  XNOR U49254 ( .A(n40081), .B(n40080), .Z(n40082) );
  XNOR U49255 ( .A(n40077), .B(n40076), .Z(n40080) );
  XOR U49256 ( .A(n40079), .B(n40078), .Z(n40076) );
  XOR U49257 ( .A(y[2288]), .B(x[2288]), .Z(n40078) );
  XOR U49258 ( .A(y[2287]), .B(x[2287]), .Z(n40079) );
  XOR U49259 ( .A(y[2286]), .B(x[2286]), .Z(n40077) );
  XOR U49260 ( .A(n40071), .B(n40070), .Z(n40081) );
  XOR U49261 ( .A(n40073), .B(n40072), .Z(n40070) );
  XOR U49262 ( .A(y[2285]), .B(x[2285]), .Z(n40072) );
  XOR U49263 ( .A(y[2284]), .B(x[2284]), .Z(n40073) );
  XOR U49264 ( .A(y[2283]), .B(x[2283]), .Z(n40071) );
  XNOR U49265 ( .A(n40047), .B(n40048), .Z(n40065) );
  XNOR U49266 ( .A(n40062), .B(n40063), .Z(n40048) );
  XOR U49267 ( .A(n40059), .B(n40058), .Z(n40063) );
  XOR U49268 ( .A(y[2280]), .B(x[2280]), .Z(n40058) );
  XOR U49269 ( .A(n40061), .B(n40060), .Z(n40059) );
  XOR U49270 ( .A(y[2282]), .B(x[2282]), .Z(n40060) );
  XOR U49271 ( .A(y[2281]), .B(x[2281]), .Z(n40061) );
  XOR U49272 ( .A(n40053), .B(n40052), .Z(n40062) );
  XOR U49273 ( .A(n40055), .B(n40054), .Z(n40052) );
  XOR U49274 ( .A(y[2279]), .B(x[2279]), .Z(n40054) );
  XOR U49275 ( .A(y[2278]), .B(x[2278]), .Z(n40055) );
  XOR U49276 ( .A(y[2277]), .B(x[2277]), .Z(n40053) );
  XNOR U49277 ( .A(n40046), .B(n40045), .Z(n40047) );
  XNOR U49278 ( .A(n40042), .B(n40041), .Z(n40045) );
  XOR U49279 ( .A(n40044), .B(n40043), .Z(n40041) );
  XOR U49280 ( .A(y[2276]), .B(x[2276]), .Z(n40043) );
  XOR U49281 ( .A(y[2275]), .B(x[2275]), .Z(n40044) );
  XOR U49282 ( .A(y[2274]), .B(x[2274]), .Z(n40042) );
  XOR U49283 ( .A(n40036), .B(n40035), .Z(n40046) );
  XOR U49284 ( .A(n40038), .B(n40037), .Z(n40035) );
  XOR U49285 ( .A(y[2273]), .B(x[2273]), .Z(n40037) );
  XOR U49286 ( .A(y[2272]), .B(x[2272]), .Z(n40038) );
  XOR U49287 ( .A(y[2271]), .B(x[2271]), .Z(n40036) );
  NAND U49288 ( .A(n40099), .B(n40100), .Z(N61818) );
  NAND U49289 ( .A(n40101), .B(n40102), .Z(n40100) );
  NANDN U49290 ( .A(n40103), .B(n40104), .Z(n40102) );
  NANDN U49291 ( .A(n40104), .B(n40103), .Z(n40099) );
  XOR U49292 ( .A(n40103), .B(n40105), .Z(N61817) );
  XNOR U49293 ( .A(n40101), .B(n40104), .Z(n40105) );
  NAND U49294 ( .A(n40106), .B(n40107), .Z(n40104) );
  NAND U49295 ( .A(n40108), .B(n40109), .Z(n40107) );
  NANDN U49296 ( .A(n40110), .B(n40111), .Z(n40109) );
  NANDN U49297 ( .A(n40111), .B(n40110), .Z(n40106) );
  AND U49298 ( .A(n40112), .B(n40113), .Z(n40101) );
  NAND U49299 ( .A(n40114), .B(n40115), .Z(n40113) );
  NANDN U49300 ( .A(n40116), .B(n40117), .Z(n40115) );
  NANDN U49301 ( .A(n40117), .B(n40116), .Z(n40112) );
  IV U49302 ( .A(n40118), .Z(n40117) );
  AND U49303 ( .A(n40119), .B(n40120), .Z(n40103) );
  NAND U49304 ( .A(n40121), .B(n40122), .Z(n40120) );
  NANDN U49305 ( .A(n40123), .B(n40124), .Z(n40122) );
  NANDN U49306 ( .A(n40124), .B(n40123), .Z(n40119) );
  XOR U49307 ( .A(n40116), .B(n40125), .Z(N61816) );
  XNOR U49308 ( .A(n40114), .B(n40118), .Z(n40125) );
  XOR U49309 ( .A(n40111), .B(n40126), .Z(n40118) );
  XNOR U49310 ( .A(n40108), .B(n40110), .Z(n40126) );
  AND U49311 ( .A(n40127), .B(n40128), .Z(n40110) );
  NANDN U49312 ( .A(n40129), .B(n40130), .Z(n40128) );
  OR U49313 ( .A(n40131), .B(n40132), .Z(n40130) );
  IV U49314 ( .A(n40133), .Z(n40132) );
  NANDN U49315 ( .A(n40133), .B(n40131), .Z(n40127) );
  AND U49316 ( .A(n40134), .B(n40135), .Z(n40108) );
  NAND U49317 ( .A(n40136), .B(n40137), .Z(n40135) );
  NANDN U49318 ( .A(n40138), .B(n40139), .Z(n40137) );
  NANDN U49319 ( .A(n40139), .B(n40138), .Z(n40134) );
  IV U49320 ( .A(n40140), .Z(n40139) );
  NAND U49321 ( .A(n40141), .B(n40142), .Z(n40111) );
  NANDN U49322 ( .A(n40143), .B(n40144), .Z(n40142) );
  NANDN U49323 ( .A(n40145), .B(n40146), .Z(n40144) );
  NANDN U49324 ( .A(n40146), .B(n40145), .Z(n40141) );
  IV U49325 ( .A(n40147), .Z(n40145) );
  AND U49326 ( .A(n40148), .B(n40149), .Z(n40114) );
  NAND U49327 ( .A(n40150), .B(n40151), .Z(n40149) );
  NANDN U49328 ( .A(n40152), .B(n40153), .Z(n40151) );
  NANDN U49329 ( .A(n40153), .B(n40152), .Z(n40148) );
  XOR U49330 ( .A(n40124), .B(n40154), .Z(n40116) );
  XNOR U49331 ( .A(n40121), .B(n40123), .Z(n40154) );
  AND U49332 ( .A(n40155), .B(n40156), .Z(n40123) );
  NANDN U49333 ( .A(n40157), .B(n40158), .Z(n40156) );
  OR U49334 ( .A(n40159), .B(n40160), .Z(n40158) );
  IV U49335 ( .A(n40161), .Z(n40160) );
  NANDN U49336 ( .A(n40161), .B(n40159), .Z(n40155) );
  AND U49337 ( .A(n40162), .B(n40163), .Z(n40121) );
  NAND U49338 ( .A(n40164), .B(n40165), .Z(n40163) );
  NANDN U49339 ( .A(n40166), .B(n40167), .Z(n40165) );
  NANDN U49340 ( .A(n40167), .B(n40166), .Z(n40162) );
  IV U49341 ( .A(n40168), .Z(n40167) );
  NAND U49342 ( .A(n40169), .B(n40170), .Z(n40124) );
  NANDN U49343 ( .A(n40171), .B(n40172), .Z(n40170) );
  NANDN U49344 ( .A(n40173), .B(n40174), .Z(n40172) );
  NANDN U49345 ( .A(n40174), .B(n40173), .Z(n40169) );
  IV U49346 ( .A(n40175), .Z(n40173) );
  XOR U49347 ( .A(n40150), .B(n40176), .Z(N61815) );
  XNOR U49348 ( .A(n40153), .B(n40152), .Z(n40176) );
  XNOR U49349 ( .A(n40164), .B(n40177), .Z(n40152) );
  XNOR U49350 ( .A(n40168), .B(n40166), .Z(n40177) );
  XOR U49351 ( .A(n40174), .B(n40178), .Z(n40166) );
  XNOR U49352 ( .A(n40171), .B(n40175), .Z(n40178) );
  AND U49353 ( .A(n40179), .B(n40180), .Z(n40175) );
  NAND U49354 ( .A(n40181), .B(n40182), .Z(n40180) );
  NAND U49355 ( .A(n40183), .B(n40184), .Z(n40179) );
  AND U49356 ( .A(n40185), .B(n40186), .Z(n40171) );
  NAND U49357 ( .A(n40187), .B(n40188), .Z(n40186) );
  NAND U49358 ( .A(n40189), .B(n40190), .Z(n40185) );
  NANDN U49359 ( .A(n40191), .B(n40192), .Z(n40174) );
  ANDN U49360 ( .B(n40193), .A(n40194), .Z(n40168) );
  XNOR U49361 ( .A(n40159), .B(n40195), .Z(n40164) );
  XNOR U49362 ( .A(n40157), .B(n40161), .Z(n40195) );
  AND U49363 ( .A(n40196), .B(n40197), .Z(n40161) );
  NAND U49364 ( .A(n40198), .B(n40199), .Z(n40197) );
  NAND U49365 ( .A(n40200), .B(n40201), .Z(n40196) );
  AND U49366 ( .A(n40202), .B(n40203), .Z(n40157) );
  NAND U49367 ( .A(n40204), .B(n40205), .Z(n40203) );
  NAND U49368 ( .A(n40206), .B(n40207), .Z(n40202) );
  AND U49369 ( .A(n40208), .B(n40209), .Z(n40159) );
  NAND U49370 ( .A(n40210), .B(n40211), .Z(n40153) );
  XNOR U49371 ( .A(n40136), .B(n40212), .Z(n40150) );
  XNOR U49372 ( .A(n40140), .B(n40138), .Z(n40212) );
  XOR U49373 ( .A(n40146), .B(n40213), .Z(n40138) );
  XNOR U49374 ( .A(n40143), .B(n40147), .Z(n40213) );
  AND U49375 ( .A(n40214), .B(n40215), .Z(n40147) );
  NAND U49376 ( .A(n40216), .B(n40217), .Z(n40215) );
  NAND U49377 ( .A(n40218), .B(n40219), .Z(n40214) );
  AND U49378 ( .A(n40220), .B(n40221), .Z(n40143) );
  NAND U49379 ( .A(n40222), .B(n40223), .Z(n40221) );
  NAND U49380 ( .A(n40224), .B(n40225), .Z(n40220) );
  NANDN U49381 ( .A(n40226), .B(n40227), .Z(n40146) );
  ANDN U49382 ( .B(n40228), .A(n40229), .Z(n40140) );
  XNOR U49383 ( .A(n40131), .B(n40230), .Z(n40136) );
  XNOR U49384 ( .A(n40129), .B(n40133), .Z(n40230) );
  AND U49385 ( .A(n40231), .B(n40232), .Z(n40133) );
  NAND U49386 ( .A(n40233), .B(n40234), .Z(n40232) );
  NAND U49387 ( .A(n40235), .B(n40236), .Z(n40231) );
  AND U49388 ( .A(n40237), .B(n40238), .Z(n40129) );
  NAND U49389 ( .A(n40239), .B(n40240), .Z(n40238) );
  NAND U49390 ( .A(n40241), .B(n40242), .Z(n40237) );
  AND U49391 ( .A(n40243), .B(n40244), .Z(n40131) );
  XOR U49392 ( .A(n40211), .B(n40210), .Z(N61814) );
  XNOR U49393 ( .A(n40228), .B(n40229), .Z(n40210) );
  XNOR U49394 ( .A(n40243), .B(n40244), .Z(n40229) );
  XOR U49395 ( .A(n40240), .B(n40239), .Z(n40244) );
  XOR U49396 ( .A(y[2268]), .B(x[2268]), .Z(n40239) );
  XOR U49397 ( .A(n40242), .B(n40241), .Z(n40240) );
  XOR U49398 ( .A(y[2270]), .B(x[2270]), .Z(n40241) );
  XOR U49399 ( .A(y[2269]), .B(x[2269]), .Z(n40242) );
  XOR U49400 ( .A(n40234), .B(n40233), .Z(n40243) );
  XOR U49401 ( .A(n40236), .B(n40235), .Z(n40233) );
  XOR U49402 ( .A(y[2267]), .B(x[2267]), .Z(n40235) );
  XOR U49403 ( .A(y[2266]), .B(x[2266]), .Z(n40236) );
  XOR U49404 ( .A(y[2265]), .B(x[2265]), .Z(n40234) );
  XNOR U49405 ( .A(n40227), .B(n40226), .Z(n40228) );
  XNOR U49406 ( .A(n40223), .B(n40222), .Z(n40226) );
  XOR U49407 ( .A(n40225), .B(n40224), .Z(n40222) );
  XOR U49408 ( .A(y[2264]), .B(x[2264]), .Z(n40224) );
  XOR U49409 ( .A(y[2263]), .B(x[2263]), .Z(n40225) );
  XOR U49410 ( .A(y[2262]), .B(x[2262]), .Z(n40223) );
  XOR U49411 ( .A(n40217), .B(n40216), .Z(n40227) );
  XOR U49412 ( .A(n40219), .B(n40218), .Z(n40216) );
  XOR U49413 ( .A(y[2261]), .B(x[2261]), .Z(n40218) );
  XOR U49414 ( .A(y[2260]), .B(x[2260]), .Z(n40219) );
  XOR U49415 ( .A(y[2259]), .B(x[2259]), .Z(n40217) );
  XNOR U49416 ( .A(n40193), .B(n40194), .Z(n40211) );
  XNOR U49417 ( .A(n40208), .B(n40209), .Z(n40194) );
  XOR U49418 ( .A(n40205), .B(n40204), .Z(n40209) );
  XOR U49419 ( .A(y[2256]), .B(x[2256]), .Z(n40204) );
  XOR U49420 ( .A(n40207), .B(n40206), .Z(n40205) );
  XOR U49421 ( .A(y[2258]), .B(x[2258]), .Z(n40206) );
  XOR U49422 ( .A(y[2257]), .B(x[2257]), .Z(n40207) );
  XOR U49423 ( .A(n40199), .B(n40198), .Z(n40208) );
  XOR U49424 ( .A(n40201), .B(n40200), .Z(n40198) );
  XOR U49425 ( .A(y[2255]), .B(x[2255]), .Z(n40200) );
  XOR U49426 ( .A(y[2254]), .B(x[2254]), .Z(n40201) );
  XOR U49427 ( .A(y[2253]), .B(x[2253]), .Z(n40199) );
  XNOR U49428 ( .A(n40192), .B(n40191), .Z(n40193) );
  XNOR U49429 ( .A(n40188), .B(n40187), .Z(n40191) );
  XOR U49430 ( .A(n40190), .B(n40189), .Z(n40187) );
  XOR U49431 ( .A(y[2252]), .B(x[2252]), .Z(n40189) );
  XOR U49432 ( .A(y[2251]), .B(x[2251]), .Z(n40190) );
  XOR U49433 ( .A(y[2250]), .B(x[2250]), .Z(n40188) );
  XOR U49434 ( .A(n40182), .B(n40181), .Z(n40192) );
  XOR U49435 ( .A(n40184), .B(n40183), .Z(n40181) );
  XOR U49436 ( .A(y[2249]), .B(x[2249]), .Z(n40183) );
  XOR U49437 ( .A(y[2248]), .B(x[2248]), .Z(n40184) );
  XOR U49438 ( .A(y[2247]), .B(x[2247]), .Z(n40182) );
  NAND U49439 ( .A(n40245), .B(n40246), .Z(N61805) );
  NAND U49440 ( .A(n40247), .B(n40248), .Z(n40246) );
  NANDN U49441 ( .A(n40249), .B(n40250), .Z(n40248) );
  NANDN U49442 ( .A(n40250), .B(n40249), .Z(n40245) );
  XOR U49443 ( .A(n40249), .B(n40251), .Z(N61804) );
  XNOR U49444 ( .A(n40247), .B(n40250), .Z(n40251) );
  NAND U49445 ( .A(n40252), .B(n40253), .Z(n40250) );
  NAND U49446 ( .A(n40254), .B(n40255), .Z(n40253) );
  NANDN U49447 ( .A(n40256), .B(n40257), .Z(n40255) );
  NANDN U49448 ( .A(n40257), .B(n40256), .Z(n40252) );
  AND U49449 ( .A(n40258), .B(n40259), .Z(n40247) );
  NAND U49450 ( .A(n40260), .B(n40261), .Z(n40259) );
  NANDN U49451 ( .A(n40262), .B(n40263), .Z(n40261) );
  NANDN U49452 ( .A(n40263), .B(n40262), .Z(n40258) );
  IV U49453 ( .A(n40264), .Z(n40263) );
  AND U49454 ( .A(n40265), .B(n40266), .Z(n40249) );
  NAND U49455 ( .A(n40267), .B(n40268), .Z(n40266) );
  NANDN U49456 ( .A(n40269), .B(n40270), .Z(n40268) );
  NANDN U49457 ( .A(n40270), .B(n40269), .Z(n40265) );
  XOR U49458 ( .A(n40262), .B(n40271), .Z(N61803) );
  XNOR U49459 ( .A(n40260), .B(n40264), .Z(n40271) );
  XOR U49460 ( .A(n40257), .B(n40272), .Z(n40264) );
  XNOR U49461 ( .A(n40254), .B(n40256), .Z(n40272) );
  AND U49462 ( .A(n40273), .B(n40274), .Z(n40256) );
  NANDN U49463 ( .A(n40275), .B(n40276), .Z(n40274) );
  OR U49464 ( .A(n40277), .B(n40278), .Z(n40276) );
  IV U49465 ( .A(n40279), .Z(n40278) );
  NANDN U49466 ( .A(n40279), .B(n40277), .Z(n40273) );
  AND U49467 ( .A(n40280), .B(n40281), .Z(n40254) );
  NAND U49468 ( .A(n40282), .B(n40283), .Z(n40281) );
  NANDN U49469 ( .A(n40284), .B(n40285), .Z(n40283) );
  NANDN U49470 ( .A(n40285), .B(n40284), .Z(n40280) );
  IV U49471 ( .A(n40286), .Z(n40285) );
  NAND U49472 ( .A(n40287), .B(n40288), .Z(n40257) );
  NANDN U49473 ( .A(n40289), .B(n40290), .Z(n40288) );
  NANDN U49474 ( .A(n40291), .B(n40292), .Z(n40290) );
  NANDN U49475 ( .A(n40292), .B(n40291), .Z(n40287) );
  IV U49476 ( .A(n40293), .Z(n40291) );
  AND U49477 ( .A(n40294), .B(n40295), .Z(n40260) );
  NAND U49478 ( .A(n40296), .B(n40297), .Z(n40295) );
  NANDN U49479 ( .A(n40298), .B(n40299), .Z(n40297) );
  NANDN U49480 ( .A(n40299), .B(n40298), .Z(n40294) );
  XOR U49481 ( .A(n40270), .B(n40300), .Z(n40262) );
  XNOR U49482 ( .A(n40267), .B(n40269), .Z(n40300) );
  AND U49483 ( .A(n40301), .B(n40302), .Z(n40269) );
  NANDN U49484 ( .A(n40303), .B(n40304), .Z(n40302) );
  OR U49485 ( .A(n40305), .B(n40306), .Z(n40304) );
  IV U49486 ( .A(n40307), .Z(n40306) );
  NANDN U49487 ( .A(n40307), .B(n40305), .Z(n40301) );
  AND U49488 ( .A(n40308), .B(n40309), .Z(n40267) );
  NAND U49489 ( .A(n40310), .B(n40311), .Z(n40309) );
  NANDN U49490 ( .A(n40312), .B(n40313), .Z(n40311) );
  NANDN U49491 ( .A(n40313), .B(n40312), .Z(n40308) );
  IV U49492 ( .A(n40314), .Z(n40313) );
  NAND U49493 ( .A(n40315), .B(n40316), .Z(n40270) );
  NANDN U49494 ( .A(n40317), .B(n40318), .Z(n40316) );
  NANDN U49495 ( .A(n40319), .B(n40320), .Z(n40318) );
  NANDN U49496 ( .A(n40320), .B(n40319), .Z(n40315) );
  IV U49497 ( .A(n40321), .Z(n40319) );
  XOR U49498 ( .A(n40296), .B(n40322), .Z(N61802) );
  XNOR U49499 ( .A(n40299), .B(n40298), .Z(n40322) );
  XNOR U49500 ( .A(n40310), .B(n40323), .Z(n40298) );
  XNOR U49501 ( .A(n40314), .B(n40312), .Z(n40323) );
  XOR U49502 ( .A(n40320), .B(n40324), .Z(n40312) );
  XNOR U49503 ( .A(n40317), .B(n40321), .Z(n40324) );
  AND U49504 ( .A(n40325), .B(n40326), .Z(n40321) );
  NAND U49505 ( .A(n40327), .B(n40328), .Z(n40326) );
  NAND U49506 ( .A(n40329), .B(n40330), .Z(n40325) );
  AND U49507 ( .A(n40331), .B(n40332), .Z(n40317) );
  NAND U49508 ( .A(n40333), .B(n40334), .Z(n40332) );
  NAND U49509 ( .A(n40335), .B(n40336), .Z(n40331) );
  NANDN U49510 ( .A(n40337), .B(n40338), .Z(n40320) );
  ANDN U49511 ( .B(n40339), .A(n40340), .Z(n40314) );
  XNOR U49512 ( .A(n40305), .B(n40341), .Z(n40310) );
  XNOR U49513 ( .A(n40303), .B(n40307), .Z(n40341) );
  AND U49514 ( .A(n40342), .B(n40343), .Z(n40307) );
  NAND U49515 ( .A(n40344), .B(n40345), .Z(n40343) );
  NAND U49516 ( .A(n40346), .B(n40347), .Z(n40342) );
  AND U49517 ( .A(n40348), .B(n40349), .Z(n40303) );
  NAND U49518 ( .A(n40350), .B(n40351), .Z(n40349) );
  NAND U49519 ( .A(n40352), .B(n40353), .Z(n40348) );
  AND U49520 ( .A(n40354), .B(n40355), .Z(n40305) );
  NAND U49521 ( .A(n40356), .B(n40357), .Z(n40299) );
  XNOR U49522 ( .A(n40282), .B(n40358), .Z(n40296) );
  XNOR U49523 ( .A(n40286), .B(n40284), .Z(n40358) );
  XOR U49524 ( .A(n40292), .B(n40359), .Z(n40284) );
  XNOR U49525 ( .A(n40289), .B(n40293), .Z(n40359) );
  AND U49526 ( .A(n40360), .B(n40361), .Z(n40293) );
  NAND U49527 ( .A(n40362), .B(n40363), .Z(n40361) );
  NAND U49528 ( .A(n40364), .B(n40365), .Z(n40360) );
  AND U49529 ( .A(n40366), .B(n40367), .Z(n40289) );
  NAND U49530 ( .A(n40368), .B(n40369), .Z(n40367) );
  NAND U49531 ( .A(n40370), .B(n40371), .Z(n40366) );
  NANDN U49532 ( .A(n40372), .B(n40373), .Z(n40292) );
  ANDN U49533 ( .B(n40374), .A(n40375), .Z(n40286) );
  XNOR U49534 ( .A(n40277), .B(n40376), .Z(n40282) );
  XNOR U49535 ( .A(n40275), .B(n40279), .Z(n40376) );
  AND U49536 ( .A(n40377), .B(n40378), .Z(n40279) );
  NAND U49537 ( .A(n40379), .B(n40380), .Z(n40378) );
  NAND U49538 ( .A(n40381), .B(n40382), .Z(n40377) );
  AND U49539 ( .A(n40383), .B(n40384), .Z(n40275) );
  NAND U49540 ( .A(n40385), .B(n40386), .Z(n40384) );
  NAND U49541 ( .A(n40387), .B(n40388), .Z(n40383) );
  AND U49542 ( .A(n40389), .B(n40390), .Z(n40277) );
  XOR U49543 ( .A(n40357), .B(n40356), .Z(N61801) );
  XNOR U49544 ( .A(n40374), .B(n40375), .Z(n40356) );
  XNOR U49545 ( .A(n40389), .B(n40390), .Z(n40375) );
  XOR U49546 ( .A(n40386), .B(n40385), .Z(n40390) );
  XOR U49547 ( .A(y[2244]), .B(x[2244]), .Z(n40385) );
  XOR U49548 ( .A(n40388), .B(n40387), .Z(n40386) );
  XOR U49549 ( .A(y[2246]), .B(x[2246]), .Z(n40387) );
  XOR U49550 ( .A(y[2245]), .B(x[2245]), .Z(n40388) );
  XOR U49551 ( .A(n40380), .B(n40379), .Z(n40389) );
  XOR U49552 ( .A(n40382), .B(n40381), .Z(n40379) );
  XOR U49553 ( .A(y[2243]), .B(x[2243]), .Z(n40381) );
  XOR U49554 ( .A(y[2242]), .B(x[2242]), .Z(n40382) );
  XOR U49555 ( .A(y[2241]), .B(x[2241]), .Z(n40380) );
  XNOR U49556 ( .A(n40373), .B(n40372), .Z(n40374) );
  XNOR U49557 ( .A(n40369), .B(n40368), .Z(n40372) );
  XOR U49558 ( .A(n40371), .B(n40370), .Z(n40368) );
  XOR U49559 ( .A(y[2240]), .B(x[2240]), .Z(n40370) );
  XOR U49560 ( .A(y[2239]), .B(x[2239]), .Z(n40371) );
  XOR U49561 ( .A(y[2238]), .B(x[2238]), .Z(n40369) );
  XOR U49562 ( .A(n40363), .B(n40362), .Z(n40373) );
  XOR U49563 ( .A(n40365), .B(n40364), .Z(n40362) );
  XOR U49564 ( .A(y[2237]), .B(x[2237]), .Z(n40364) );
  XOR U49565 ( .A(y[2236]), .B(x[2236]), .Z(n40365) );
  XOR U49566 ( .A(y[2235]), .B(x[2235]), .Z(n40363) );
  XNOR U49567 ( .A(n40339), .B(n40340), .Z(n40357) );
  XNOR U49568 ( .A(n40354), .B(n40355), .Z(n40340) );
  XOR U49569 ( .A(n40351), .B(n40350), .Z(n40355) );
  XOR U49570 ( .A(y[2232]), .B(x[2232]), .Z(n40350) );
  XOR U49571 ( .A(n40353), .B(n40352), .Z(n40351) );
  XOR U49572 ( .A(y[2234]), .B(x[2234]), .Z(n40352) );
  XOR U49573 ( .A(y[2233]), .B(x[2233]), .Z(n40353) );
  XOR U49574 ( .A(n40345), .B(n40344), .Z(n40354) );
  XOR U49575 ( .A(n40347), .B(n40346), .Z(n40344) );
  XOR U49576 ( .A(y[2231]), .B(x[2231]), .Z(n40346) );
  XOR U49577 ( .A(y[2230]), .B(x[2230]), .Z(n40347) );
  XOR U49578 ( .A(y[2229]), .B(x[2229]), .Z(n40345) );
  XNOR U49579 ( .A(n40338), .B(n40337), .Z(n40339) );
  XNOR U49580 ( .A(n40334), .B(n40333), .Z(n40337) );
  XOR U49581 ( .A(n40336), .B(n40335), .Z(n40333) );
  XOR U49582 ( .A(y[2228]), .B(x[2228]), .Z(n40335) );
  XOR U49583 ( .A(y[2227]), .B(x[2227]), .Z(n40336) );
  XOR U49584 ( .A(y[2226]), .B(x[2226]), .Z(n40334) );
  XOR U49585 ( .A(n40328), .B(n40327), .Z(n40338) );
  XOR U49586 ( .A(n40330), .B(n40329), .Z(n40327) );
  XOR U49587 ( .A(y[2225]), .B(x[2225]), .Z(n40329) );
  XOR U49588 ( .A(y[2224]), .B(x[2224]), .Z(n40330) );
  XOR U49589 ( .A(y[2223]), .B(x[2223]), .Z(n40328) );
  NAND U49590 ( .A(n40391), .B(n40392), .Z(N61792) );
  NAND U49591 ( .A(n40393), .B(n40394), .Z(n40392) );
  NANDN U49592 ( .A(n40395), .B(n40396), .Z(n40394) );
  NANDN U49593 ( .A(n40396), .B(n40395), .Z(n40391) );
  XOR U49594 ( .A(n40395), .B(n40397), .Z(N61791) );
  XNOR U49595 ( .A(n40393), .B(n40396), .Z(n40397) );
  NAND U49596 ( .A(n40398), .B(n40399), .Z(n40396) );
  NAND U49597 ( .A(n40400), .B(n40401), .Z(n40399) );
  NANDN U49598 ( .A(n40402), .B(n40403), .Z(n40401) );
  NANDN U49599 ( .A(n40403), .B(n40402), .Z(n40398) );
  AND U49600 ( .A(n40404), .B(n40405), .Z(n40393) );
  NAND U49601 ( .A(n40406), .B(n40407), .Z(n40405) );
  NANDN U49602 ( .A(n40408), .B(n40409), .Z(n40407) );
  NANDN U49603 ( .A(n40409), .B(n40408), .Z(n40404) );
  IV U49604 ( .A(n40410), .Z(n40409) );
  AND U49605 ( .A(n40411), .B(n40412), .Z(n40395) );
  NAND U49606 ( .A(n40413), .B(n40414), .Z(n40412) );
  NANDN U49607 ( .A(n40415), .B(n40416), .Z(n40414) );
  NANDN U49608 ( .A(n40416), .B(n40415), .Z(n40411) );
  XOR U49609 ( .A(n40408), .B(n40417), .Z(N61790) );
  XNOR U49610 ( .A(n40406), .B(n40410), .Z(n40417) );
  XOR U49611 ( .A(n40403), .B(n40418), .Z(n40410) );
  XNOR U49612 ( .A(n40400), .B(n40402), .Z(n40418) );
  AND U49613 ( .A(n40419), .B(n40420), .Z(n40402) );
  NANDN U49614 ( .A(n40421), .B(n40422), .Z(n40420) );
  OR U49615 ( .A(n40423), .B(n40424), .Z(n40422) );
  IV U49616 ( .A(n40425), .Z(n40424) );
  NANDN U49617 ( .A(n40425), .B(n40423), .Z(n40419) );
  AND U49618 ( .A(n40426), .B(n40427), .Z(n40400) );
  NAND U49619 ( .A(n40428), .B(n40429), .Z(n40427) );
  NANDN U49620 ( .A(n40430), .B(n40431), .Z(n40429) );
  NANDN U49621 ( .A(n40431), .B(n40430), .Z(n40426) );
  IV U49622 ( .A(n40432), .Z(n40431) );
  NAND U49623 ( .A(n40433), .B(n40434), .Z(n40403) );
  NANDN U49624 ( .A(n40435), .B(n40436), .Z(n40434) );
  NANDN U49625 ( .A(n40437), .B(n40438), .Z(n40436) );
  NANDN U49626 ( .A(n40438), .B(n40437), .Z(n40433) );
  IV U49627 ( .A(n40439), .Z(n40437) );
  AND U49628 ( .A(n40440), .B(n40441), .Z(n40406) );
  NAND U49629 ( .A(n40442), .B(n40443), .Z(n40441) );
  NANDN U49630 ( .A(n40444), .B(n40445), .Z(n40443) );
  NANDN U49631 ( .A(n40445), .B(n40444), .Z(n40440) );
  XOR U49632 ( .A(n40416), .B(n40446), .Z(n40408) );
  XNOR U49633 ( .A(n40413), .B(n40415), .Z(n40446) );
  AND U49634 ( .A(n40447), .B(n40448), .Z(n40415) );
  NANDN U49635 ( .A(n40449), .B(n40450), .Z(n40448) );
  OR U49636 ( .A(n40451), .B(n40452), .Z(n40450) );
  IV U49637 ( .A(n40453), .Z(n40452) );
  NANDN U49638 ( .A(n40453), .B(n40451), .Z(n40447) );
  AND U49639 ( .A(n40454), .B(n40455), .Z(n40413) );
  NAND U49640 ( .A(n40456), .B(n40457), .Z(n40455) );
  NANDN U49641 ( .A(n40458), .B(n40459), .Z(n40457) );
  NANDN U49642 ( .A(n40459), .B(n40458), .Z(n40454) );
  IV U49643 ( .A(n40460), .Z(n40459) );
  NAND U49644 ( .A(n40461), .B(n40462), .Z(n40416) );
  NANDN U49645 ( .A(n40463), .B(n40464), .Z(n40462) );
  NANDN U49646 ( .A(n40465), .B(n40466), .Z(n40464) );
  NANDN U49647 ( .A(n40466), .B(n40465), .Z(n40461) );
  IV U49648 ( .A(n40467), .Z(n40465) );
  XOR U49649 ( .A(n40442), .B(n40468), .Z(N61789) );
  XNOR U49650 ( .A(n40445), .B(n40444), .Z(n40468) );
  XNOR U49651 ( .A(n40456), .B(n40469), .Z(n40444) );
  XNOR U49652 ( .A(n40460), .B(n40458), .Z(n40469) );
  XOR U49653 ( .A(n40466), .B(n40470), .Z(n40458) );
  XNOR U49654 ( .A(n40463), .B(n40467), .Z(n40470) );
  AND U49655 ( .A(n40471), .B(n40472), .Z(n40467) );
  NAND U49656 ( .A(n40473), .B(n40474), .Z(n40472) );
  NAND U49657 ( .A(n40475), .B(n40476), .Z(n40471) );
  AND U49658 ( .A(n40477), .B(n40478), .Z(n40463) );
  NAND U49659 ( .A(n40479), .B(n40480), .Z(n40478) );
  NAND U49660 ( .A(n40481), .B(n40482), .Z(n40477) );
  NANDN U49661 ( .A(n40483), .B(n40484), .Z(n40466) );
  ANDN U49662 ( .B(n40485), .A(n40486), .Z(n40460) );
  XNOR U49663 ( .A(n40451), .B(n40487), .Z(n40456) );
  XNOR U49664 ( .A(n40449), .B(n40453), .Z(n40487) );
  AND U49665 ( .A(n40488), .B(n40489), .Z(n40453) );
  NAND U49666 ( .A(n40490), .B(n40491), .Z(n40489) );
  NAND U49667 ( .A(n40492), .B(n40493), .Z(n40488) );
  AND U49668 ( .A(n40494), .B(n40495), .Z(n40449) );
  NAND U49669 ( .A(n40496), .B(n40497), .Z(n40495) );
  NAND U49670 ( .A(n40498), .B(n40499), .Z(n40494) );
  AND U49671 ( .A(n40500), .B(n40501), .Z(n40451) );
  NAND U49672 ( .A(n40502), .B(n40503), .Z(n40445) );
  XNOR U49673 ( .A(n40428), .B(n40504), .Z(n40442) );
  XNOR U49674 ( .A(n40432), .B(n40430), .Z(n40504) );
  XOR U49675 ( .A(n40438), .B(n40505), .Z(n40430) );
  XNOR U49676 ( .A(n40435), .B(n40439), .Z(n40505) );
  AND U49677 ( .A(n40506), .B(n40507), .Z(n40439) );
  NAND U49678 ( .A(n40508), .B(n40509), .Z(n40507) );
  NAND U49679 ( .A(n40510), .B(n40511), .Z(n40506) );
  AND U49680 ( .A(n40512), .B(n40513), .Z(n40435) );
  NAND U49681 ( .A(n40514), .B(n40515), .Z(n40513) );
  NAND U49682 ( .A(n40516), .B(n40517), .Z(n40512) );
  NANDN U49683 ( .A(n40518), .B(n40519), .Z(n40438) );
  ANDN U49684 ( .B(n40520), .A(n40521), .Z(n40432) );
  XNOR U49685 ( .A(n40423), .B(n40522), .Z(n40428) );
  XNOR U49686 ( .A(n40421), .B(n40425), .Z(n40522) );
  AND U49687 ( .A(n40523), .B(n40524), .Z(n40425) );
  NAND U49688 ( .A(n40525), .B(n40526), .Z(n40524) );
  NAND U49689 ( .A(n40527), .B(n40528), .Z(n40523) );
  AND U49690 ( .A(n40529), .B(n40530), .Z(n40421) );
  NAND U49691 ( .A(n40531), .B(n40532), .Z(n40530) );
  NAND U49692 ( .A(n40533), .B(n40534), .Z(n40529) );
  AND U49693 ( .A(n40535), .B(n40536), .Z(n40423) );
  XOR U49694 ( .A(n40503), .B(n40502), .Z(N61788) );
  XNOR U49695 ( .A(n40520), .B(n40521), .Z(n40502) );
  XNOR U49696 ( .A(n40535), .B(n40536), .Z(n40521) );
  XOR U49697 ( .A(n40532), .B(n40531), .Z(n40536) );
  XOR U49698 ( .A(y[2220]), .B(x[2220]), .Z(n40531) );
  XOR U49699 ( .A(n40534), .B(n40533), .Z(n40532) );
  XOR U49700 ( .A(y[2222]), .B(x[2222]), .Z(n40533) );
  XOR U49701 ( .A(y[2221]), .B(x[2221]), .Z(n40534) );
  XOR U49702 ( .A(n40526), .B(n40525), .Z(n40535) );
  XOR U49703 ( .A(n40528), .B(n40527), .Z(n40525) );
  XOR U49704 ( .A(y[2219]), .B(x[2219]), .Z(n40527) );
  XOR U49705 ( .A(y[2218]), .B(x[2218]), .Z(n40528) );
  XOR U49706 ( .A(y[2217]), .B(x[2217]), .Z(n40526) );
  XNOR U49707 ( .A(n40519), .B(n40518), .Z(n40520) );
  XNOR U49708 ( .A(n40515), .B(n40514), .Z(n40518) );
  XOR U49709 ( .A(n40517), .B(n40516), .Z(n40514) );
  XOR U49710 ( .A(y[2216]), .B(x[2216]), .Z(n40516) );
  XOR U49711 ( .A(y[2215]), .B(x[2215]), .Z(n40517) );
  XOR U49712 ( .A(y[2214]), .B(x[2214]), .Z(n40515) );
  XOR U49713 ( .A(n40509), .B(n40508), .Z(n40519) );
  XOR U49714 ( .A(n40511), .B(n40510), .Z(n40508) );
  XOR U49715 ( .A(y[2213]), .B(x[2213]), .Z(n40510) );
  XOR U49716 ( .A(y[2212]), .B(x[2212]), .Z(n40511) );
  XOR U49717 ( .A(y[2211]), .B(x[2211]), .Z(n40509) );
  XNOR U49718 ( .A(n40485), .B(n40486), .Z(n40503) );
  XNOR U49719 ( .A(n40500), .B(n40501), .Z(n40486) );
  XOR U49720 ( .A(n40497), .B(n40496), .Z(n40501) );
  XOR U49721 ( .A(y[2208]), .B(x[2208]), .Z(n40496) );
  XOR U49722 ( .A(n40499), .B(n40498), .Z(n40497) );
  XOR U49723 ( .A(y[2210]), .B(x[2210]), .Z(n40498) );
  XOR U49724 ( .A(y[2209]), .B(x[2209]), .Z(n40499) );
  XOR U49725 ( .A(n40491), .B(n40490), .Z(n40500) );
  XOR U49726 ( .A(n40493), .B(n40492), .Z(n40490) );
  XOR U49727 ( .A(y[2207]), .B(x[2207]), .Z(n40492) );
  XOR U49728 ( .A(y[2206]), .B(x[2206]), .Z(n40493) );
  XOR U49729 ( .A(y[2205]), .B(x[2205]), .Z(n40491) );
  XNOR U49730 ( .A(n40484), .B(n40483), .Z(n40485) );
  XNOR U49731 ( .A(n40480), .B(n40479), .Z(n40483) );
  XOR U49732 ( .A(n40482), .B(n40481), .Z(n40479) );
  XOR U49733 ( .A(y[2204]), .B(x[2204]), .Z(n40481) );
  XOR U49734 ( .A(y[2203]), .B(x[2203]), .Z(n40482) );
  XOR U49735 ( .A(y[2202]), .B(x[2202]), .Z(n40480) );
  XOR U49736 ( .A(n40474), .B(n40473), .Z(n40484) );
  XOR U49737 ( .A(n40476), .B(n40475), .Z(n40473) );
  XOR U49738 ( .A(y[2201]), .B(x[2201]), .Z(n40475) );
  XOR U49739 ( .A(y[2200]), .B(x[2200]), .Z(n40476) );
  XOR U49740 ( .A(y[2199]), .B(x[2199]), .Z(n40474) );
  NAND U49741 ( .A(n40537), .B(n40538), .Z(N61779) );
  NAND U49742 ( .A(n40539), .B(n40540), .Z(n40538) );
  NANDN U49743 ( .A(n40541), .B(n40542), .Z(n40540) );
  NANDN U49744 ( .A(n40542), .B(n40541), .Z(n40537) );
  XOR U49745 ( .A(n40541), .B(n40543), .Z(N61778) );
  XNOR U49746 ( .A(n40539), .B(n40542), .Z(n40543) );
  NAND U49747 ( .A(n40544), .B(n40545), .Z(n40542) );
  NAND U49748 ( .A(n40546), .B(n40547), .Z(n40545) );
  NANDN U49749 ( .A(n40548), .B(n40549), .Z(n40547) );
  NANDN U49750 ( .A(n40549), .B(n40548), .Z(n40544) );
  AND U49751 ( .A(n40550), .B(n40551), .Z(n40539) );
  NAND U49752 ( .A(n40552), .B(n40553), .Z(n40551) );
  NANDN U49753 ( .A(n40554), .B(n40555), .Z(n40553) );
  NANDN U49754 ( .A(n40555), .B(n40554), .Z(n40550) );
  IV U49755 ( .A(n40556), .Z(n40555) );
  AND U49756 ( .A(n40557), .B(n40558), .Z(n40541) );
  NAND U49757 ( .A(n40559), .B(n40560), .Z(n40558) );
  NANDN U49758 ( .A(n40561), .B(n40562), .Z(n40560) );
  NANDN U49759 ( .A(n40562), .B(n40561), .Z(n40557) );
  XOR U49760 ( .A(n40554), .B(n40563), .Z(N61777) );
  XNOR U49761 ( .A(n40552), .B(n40556), .Z(n40563) );
  XOR U49762 ( .A(n40549), .B(n40564), .Z(n40556) );
  XNOR U49763 ( .A(n40546), .B(n40548), .Z(n40564) );
  AND U49764 ( .A(n40565), .B(n40566), .Z(n40548) );
  NANDN U49765 ( .A(n40567), .B(n40568), .Z(n40566) );
  OR U49766 ( .A(n40569), .B(n40570), .Z(n40568) );
  IV U49767 ( .A(n40571), .Z(n40570) );
  NANDN U49768 ( .A(n40571), .B(n40569), .Z(n40565) );
  AND U49769 ( .A(n40572), .B(n40573), .Z(n40546) );
  NAND U49770 ( .A(n40574), .B(n40575), .Z(n40573) );
  NANDN U49771 ( .A(n40576), .B(n40577), .Z(n40575) );
  NANDN U49772 ( .A(n40577), .B(n40576), .Z(n40572) );
  IV U49773 ( .A(n40578), .Z(n40577) );
  NAND U49774 ( .A(n40579), .B(n40580), .Z(n40549) );
  NANDN U49775 ( .A(n40581), .B(n40582), .Z(n40580) );
  NANDN U49776 ( .A(n40583), .B(n40584), .Z(n40582) );
  NANDN U49777 ( .A(n40584), .B(n40583), .Z(n40579) );
  IV U49778 ( .A(n40585), .Z(n40583) );
  AND U49779 ( .A(n40586), .B(n40587), .Z(n40552) );
  NAND U49780 ( .A(n40588), .B(n40589), .Z(n40587) );
  NANDN U49781 ( .A(n40590), .B(n40591), .Z(n40589) );
  NANDN U49782 ( .A(n40591), .B(n40590), .Z(n40586) );
  XOR U49783 ( .A(n40562), .B(n40592), .Z(n40554) );
  XNOR U49784 ( .A(n40559), .B(n40561), .Z(n40592) );
  AND U49785 ( .A(n40593), .B(n40594), .Z(n40561) );
  NANDN U49786 ( .A(n40595), .B(n40596), .Z(n40594) );
  OR U49787 ( .A(n40597), .B(n40598), .Z(n40596) );
  IV U49788 ( .A(n40599), .Z(n40598) );
  NANDN U49789 ( .A(n40599), .B(n40597), .Z(n40593) );
  AND U49790 ( .A(n40600), .B(n40601), .Z(n40559) );
  NAND U49791 ( .A(n40602), .B(n40603), .Z(n40601) );
  NANDN U49792 ( .A(n40604), .B(n40605), .Z(n40603) );
  NANDN U49793 ( .A(n40605), .B(n40604), .Z(n40600) );
  IV U49794 ( .A(n40606), .Z(n40605) );
  NAND U49795 ( .A(n40607), .B(n40608), .Z(n40562) );
  NANDN U49796 ( .A(n40609), .B(n40610), .Z(n40608) );
  NANDN U49797 ( .A(n40611), .B(n40612), .Z(n40610) );
  NANDN U49798 ( .A(n40612), .B(n40611), .Z(n40607) );
  IV U49799 ( .A(n40613), .Z(n40611) );
  XOR U49800 ( .A(n40588), .B(n40614), .Z(N61776) );
  XNOR U49801 ( .A(n40591), .B(n40590), .Z(n40614) );
  XNOR U49802 ( .A(n40602), .B(n40615), .Z(n40590) );
  XNOR U49803 ( .A(n40606), .B(n40604), .Z(n40615) );
  XOR U49804 ( .A(n40612), .B(n40616), .Z(n40604) );
  XNOR U49805 ( .A(n40609), .B(n40613), .Z(n40616) );
  AND U49806 ( .A(n40617), .B(n40618), .Z(n40613) );
  NAND U49807 ( .A(n40619), .B(n40620), .Z(n40618) );
  NAND U49808 ( .A(n40621), .B(n40622), .Z(n40617) );
  AND U49809 ( .A(n40623), .B(n40624), .Z(n40609) );
  NAND U49810 ( .A(n40625), .B(n40626), .Z(n40624) );
  NAND U49811 ( .A(n40627), .B(n40628), .Z(n40623) );
  NANDN U49812 ( .A(n40629), .B(n40630), .Z(n40612) );
  ANDN U49813 ( .B(n40631), .A(n40632), .Z(n40606) );
  XNOR U49814 ( .A(n40597), .B(n40633), .Z(n40602) );
  XNOR U49815 ( .A(n40595), .B(n40599), .Z(n40633) );
  AND U49816 ( .A(n40634), .B(n40635), .Z(n40599) );
  NAND U49817 ( .A(n40636), .B(n40637), .Z(n40635) );
  NAND U49818 ( .A(n40638), .B(n40639), .Z(n40634) );
  AND U49819 ( .A(n40640), .B(n40641), .Z(n40595) );
  NAND U49820 ( .A(n40642), .B(n40643), .Z(n40641) );
  NAND U49821 ( .A(n40644), .B(n40645), .Z(n40640) );
  AND U49822 ( .A(n40646), .B(n40647), .Z(n40597) );
  NAND U49823 ( .A(n40648), .B(n40649), .Z(n40591) );
  XNOR U49824 ( .A(n40574), .B(n40650), .Z(n40588) );
  XNOR U49825 ( .A(n40578), .B(n40576), .Z(n40650) );
  XOR U49826 ( .A(n40584), .B(n40651), .Z(n40576) );
  XNOR U49827 ( .A(n40581), .B(n40585), .Z(n40651) );
  AND U49828 ( .A(n40652), .B(n40653), .Z(n40585) );
  NAND U49829 ( .A(n40654), .B(n40655), .Z(n40653) );
  NAND U49830 ( .A(n40656), .B(n40657), .Z(n40652) );
  AND U49831 ( .A(n40658), .B(n40659), .Z(n40581) );
  NAND U49832 ( .A(n40660), .B(n40661), .Z(n40659) );
  NAND U49833 ( .A(n40662), .B(n40663), .Z(n40658) );
  NANDN U49834 ( .A(n40664), .B(n40665), .Z(n40584) );
  ANDN U49835 ( .B(n40666), .A(n40667), .Z(n40578) );
  XNOR U49836 ( .A(n40569), .B(n40668), .Z(n40574) );
  XNOR U49837 ( .A(n40567), .B(n40571), .Z(n40668) );
  AND U49838 ( .A(n40669), .B(n40670), .Z(n40571) );
  NAND U49839 ( .A(n40671), .B(n40672), .Z(n40670) );
  NAND U49840 ( .A(n40673), .B(n40674), .Z(n40669) );
  AND U49841 ( .A(n40675), .B(n40676), .Z(n40567) );
  NAND U49842 ( .A(n40677), .B(n40678), .Z(n40676) );
  NAND U49843 ( .A(n40679), .B(n40680), .Z(n40675) );
  AND U49844 ( .A(n40681), .B(n40682), .Z(n40569) );
  XOR U49845 ( .A(n40649), .B(n40648), .Z(N61775) );
  XNOR U49846 ( .A(n40666), .B(n40667), .Z(n40648) );
  XNOR U49847 ( .A(n40681), .B(n40682), .Z(n40667) );
  XOR U49848 ( .A(n40678), .B(n40677), .Z(n40682) );
  XOR U49849 ( .A(y[2196]), .B(x[2196]), .Z(n40677) );
  XOR U49850 ( .A(n40680), .B(n40679), .Z(n40678) );
  XOR U49851 ( .A(y[2198]), .B(x[2198]), .Z(n40679) );
  XOR U49852 ( .A(y[2197]), .B(x[2197]), .Z(n40680) );
  XOR U49853 ( .A(n40672), .B(n40671), .Z(n40681) );
  XOR U49854 ( .A(n40674), .B(n40673), .Z(n40671) );
  XOR U49855 ( .A(y[2195]), .B(x[2195]), .Z(n40673) );
  XOR U49856 ( .A(y[2194]), .B(x[2194]), .Z(n40674) );
  XOR U49857 ( .A(y[2193]), .B(x[2193]), .Z(n40672) );
  XNOR U49858 ( .A(n40665), .B(n40664), .Z(n40666) );
  XNOR U49859 ( .A(n40661), .B(n40660), .Z(n40664) );
  XOR U49860 ( .A(n40663), .B(n40662), .Z(n40660) );
  XOR U49861 ( .A(y[2192]), .B(x[2192]), .Z(n40662) );
  XOR U49862 ( .A(y[2191]), .B(x[2191]), .Z(n40663) );
  XOR U49863 ( .A(y[2190]), .B(x[2190]), .Z(n40661) );
  XOR U49864 ( .A(n40655), .B(n40654), .Z(n40665) );
  XOR U49865 ( .A(n40657), .B(n40656), .Z(n40654) );
  XOR U49866 ( .A(y[2189]), .B(x[2189]), .Z(n40656) );
  XOR U49867 ( .A(y[2188]), .B(x[2188]), .Z(n40657) );
  XOR U49868 ( .A(y[2187]), .B(x[2187]), .Z(n40655) );
  XNOR U49869 ( .A(n40631), .B(n40632), .Z(n40649) );
  XNOR U49870 ( .A(n40646), .B(n40647), .Z(n40632) );
  XOR U49871 ( .A(n40643), .B(n40642), .Z(n40647) );
  XOR U49872 ( .A(y[2184]), .B(x[2184]), .Z(n40642) );
  XOR U49873 ( .A(n40645), .B(n40644), .Z(n40643) );
  XOR U49874 ( .A(y[2186]), .B(x[2186]), .Z(n40644) );
  XOR U49875 ( .A(y[2185]), .B(x[2185]), .Z(n40645) );
  XOR U49876 ( .A(n40637), .B(n40636), .Z(n40646) );
  XOR U49877 ( .A(n40639), .B(n40638), .Z(n40636) );
  XOR U49878 ( .A(y[2183]), .B(x[2183]), .Z(n40638) );
  XOR U49879 ( .A(y[2182]), .B(x[2182]), .Z(n40639) );
  XOR U49880 ( .A(y[2181]), .B(x[2181]), .Z(n40637) );
  XNOR U49881 ( .A(n40630), .B(n40629), .Z(n40631) );
  XNOR U49882 ( .A(n40626), .B(n40625), .Z(n40629) );
  XOR U49883 ( .A(n40628), .B(n40627), .Z(n40625) );
  XOR U49884 ( .A(y[2180]), .B(x[2180]), .Z(n40627) );
  XOR U49885 ( .A(y[2179]), .B(x[2179]), .Z(n40628) );
  XOR U49886 ( .A(y[2178]), .B(x[2178]), .Z(n40626) );
  XOR U49887 ( .A(n40620), .B(n40619), .Z(n40630) );
  XOR U49888 ( .A(n40622), .B(n40621), .Z(n40619) );
  XOR U49889 ( .A(y[2177]), .B(x[2177]), .Z(n40621) );
  XOR U49890 ( .A(y[2176]), .B(x[2176]), .Z(n40622) );
  XOR U49891 ( .A(y[2175]), .B(x[2175]), .Z(n40620) );
  NAND U49892 ( .A(n40683), .B(n40684), .Z(N61766) );
  NAND U49893 ( .A(n40685), .B(n40686), .Z(n40684) );
  NANDN U49894 ( .A(n40687), .B(n40688), .Z(n40686) );
  NANDN U49895 ( .A(n40688), .B(n40687), .Z(n40683) );
  XOR U49896 ( .A(n40687), .B(n40689), .Z(N61765) );
  XNOR U49897 ( .A(n40685), .B(n40688), .Z(n40689) );
  NAND U49898 ( .A(n40690), .B(n40691), .Z(n40688) );
  NAND U49899 ( .A(n40692), .B(n40693), .Z(n40691) );
  NANDN U49900 ( .A(n40694), .B(n40695), .Z(n40693) );
  NANDN U49901 ( .A(n40695), .B(n40694), .Z(n40690) );
  AND U49902 ( .A(n40696), .B(n40697), .Z(n40685) );
  NAND U49903 ( .A(n40698), .B(n40699), .Z(n40697) );
  NANDN U49904 ( .A(n40700), .B(n40701), .Z(n40699) );
  NANDN U49905 ( .A(n40701), .B(n40700), .Z(n40696) );
  IV U49906 ( .A(n40702), .Z(n40701) );
  AND U49907 ( .A(n40703), .B(n40704), .Z(n40687) );
  NAND U49908 ( .A(n40705), .B(n40706), .Z(n40704) );
  NANDN U49909 ( .A(n40707), .B(n40708), .Z(n40706) );
  NANDN U49910 ( .A(n40708), .B(n40707), .Z(n40703) );
  XOR U49911 ( .A(n40700), .B(n40709), .Z(N61764) );
  XNOR U49912 ( .A(n40698), .B(n40702), .Z(n40709) );
  XOR U49913 ( .A(n40695), .B(n40710), .Z(n40702) );
  XNOR U49914 ( .A(n40692), .B(n40694), .Z(n40710) );
  AND U49915 ( .A(n40711), .B(n40712), .Z(n40694) );
  NANDN U49916 ( .A(n40713), .B(n40714), .Z(n40712) );
  OR U49917 ( .A(n40715), .B(n40716), .Z(n40714) );
  IV U49918 ( .A(n40717), .Z(n40716) );
  NANDN U49919 ( .A(n40717), .B(n40715), .Z(n40711) );
  AND U49920 ( .A(n40718), .B(n40719), .Z(n40692) );
  NAND U49921 ( .A(n40720), .B(n40721), .Z(n40719) );
  NANDN U49922 ( .A(n40722), .B(n40723), .Z(n40721) );
  NANDN U49923 ( .A(n40723), .B(n40722), .Z(n40718) );
  IV U49924 ( .A(n40724), .Z(n40723) );
  NAND U49925 ( .A(n40725), .B(n40726), .Z(n40695) );
  NANDN U49926 ( .A(n40727), .B(n40728), .Z(n40726) );
  NANDN U49927 ( .A(n40729), .B(n40730), .Z(n40728) );
  NANDN U49928 ( .A(n40730), .B(n40729), .Z(n40725) );
  IV U49929 ( .A(n40731), .Z(n40729) );
  AND U49930 ( .A(n40732), .B(n40733), .Z(n40698) );
  NAND U49931 ( .A(n40734), .B(n40735), .Z(n40733) );
  NANDN U49932 ( .A(n40736), .B(n40737), .Z(n40735) );
  NANDN U49933 ( .A(n40737), .B(n40736), .Z(n40732) );
  XOR U49934 ( .A(n40708), .B(n40738), .Z(n40700) );
  XNOR U49935 ( .A(n40705), .B(n40707), .Z(n40738) );
  AND U49936 ( .A(n40739), .B(n40740), .Z(n40707) );
  NANDN U49937 ( .A(n40741), .B(n40742), .Z(n40740) );
  OR U49938 ( .A(n40743), .B(n40744), .Z(n40742) );
  IV U49939 ( .A(n40745), .Z(n40744) );
  NANDN U49940 ( .A(n40745), .B(n40743), .Z(n40739) );
  AND U49941 ( .A(n40746), .B(n40747), .Z(n40705) );
  NAND U49942 ( .A(n40748), .B(n40749), .Z(n40747) );
  NANDN U49943 ( .A(n40750), .B(n40751), .Z(n40749) );
  NANDN U49944 ( .A(n40751), .B(n40750), .Z(n40746) );
  IV U49945 ( .A(n40752), .Z(n40751) );
  NAND U49946 ( .A(n40753), .B(n40754), .Z(n40708) );
  NANDN U49947 ( .A(n40755), .B(n40756), .Z(n40754) );
  NANDN U49948 ( .A(n40757), .B(n40758), .Z(n40756) );
  NANDN U49949 ( .A(n40758), .B(n40757), .Z(n40753) );
  IV U49950 ( .A(n40759), .Z(n40757) );
  XOR U49951 ( .A(n40734), .B(n40760), .Z(N61763) );
  XNOR U49952 ( .A(n40737), .B(n40736), .Z(n40760) );
  XNOR U49953 ( .A(n40748), .B(n40761), .Z(n40736) );
  XNOR U49954 ( .A(n40752), .B(n40750), .Z(n40761) );
  XOR U49955 ( .A(n40758), .B(n40762), .Z(n40750) );
  XNOR U49956 ( .A(n40755), .B(n40759), .Z(n40762) );
  AND U49957 ( .A(n40763), .B(n40764), .Z(n40759) );
  NAND U49958 ( .A(n40765), .B(n40766), .Z(n40764) );
  NAND U49959 ( .A(n40767), .B(n40768), .Z(n40763) );
  AND U49960 ( .A(n40769), .B(n40770), .Z(n40755) );
  NAND U49961 ( .A(n40771), .B(n40772), .Z(n40770) );
  NAND U49962 ( .A(n40773), .B(n40774), .Z(n40769) );
  NANDN U49963 ( .A(n40775), .B(n40776), .Z(n40758) );
  ANDN U49964 ( .B(n40777), .A(n40778), .Z(n40752) );
  XNOR U49965 ( .A(n40743), .B(n40779), .Z(n40748) );
  XNOR U49966 ( .A(n40741), .B(n40745), .Z(n40779) );
  AND U49967 ( .A(n40780), .B(n40781), .Z(n40745) );
  NAND U49968 ( .A(n40782), .B(n40783), .Z(n40781) );
  NAND U49969 ( .A(n40784), .B(n40785), .Z(n40780) );
  AND U49970 ( .A(n40786), .B(n40787), .Z(n40741) );
  NAND U49971 ( .A(n40788), .B(n40789), .Z(n40787) );
  NAND U49972 ( .A(n40790), .B(n40791), .Z(n40786) );
  AND U49973 ( .A(n40792), .B(n40793), .Z(n40743) );
  NAND U49974 ( .A(n40794), .B(n40795), .Z(n40737) );
  XNOR U49975 ( .A(n40720), .B(n40796), .Z(n40734) );
  XNOR U49976 ( .A(n40724), .B(n40722), .Z(n40796) );
  XOR U49977 ( .A(n40730), .B(n40797), .Z(n40722) );
  XNOR U49978 ( .A(n40727), .B(n40731), .Z(n40797) );
  AND U49979 ( .A(n40798), .B(n40799), .Z(n40731) );
  NAND U49980 ( .A(n40800), .B(n40801), .Z(n40799) );
  NAND U49981 ( .A(n40802), .B(n40803), .Z(n40798) );
  AND U49982 ( .A(n40804), .B(n40805), .Z(n40727) );
  NAND U49983 ( .A(n40806), .B(n40807), .Z(n40805) );
  NAND U49984 ( .A(n40808), .B(n40809), .Z(n40804) );
  NANDN U49985 ( .A(n40810), .B(n40811), .Z(n40730) );
  ANDN U49986 ( .B(n40812), .A(n40813), .Z(n40724) );
  XNOR U49987 ( .A(n40715), .B(n40814), .Z(n40720) );
  XNOR U49988 ( .A(n40713), .B(n40717), .Z(n40814) );
  AND U49989 ( .A(n40815), .B(n40816), .Z(n40717) );
  NAND U49990 ( .A(n40817), .B(n40818), .Z(n40816) );
  NAND U49991 ( .A(n40819), .B(n40820), .Z(n40815) );
  AND U49992 ( .A(n40821), .B(n40822), .Z(n40713) );
  NAND U49993 ( .A(n40823), .B(n40824), .Z(n40822) );
  NAND U49994 ( .A(n40825), .B(n40826), .Z(n40821) );
  AND U49995 ( .A(n40827), .B(n40828), .Z(n40715) );
  XOR U49996 ( .A(n40795), .B(n40794), .Z(N61762) );
  XNOR U49997 ( .A(n40812), .B(n40813), .Z(n40794) );
  XNOR U49998 ( .A(n40827), .B(n40828), .Z(n40813) );
  XOR U49999 ( .A(n40824), .B(n40823), .Z(n40828) );
  XOR U50000 ( .A(y[2172]), .B(x[2172]), .Z(n40823) );
  XOR U50001 ( .A(n40826), .B(n40825), .Z(n40824) );
  XOR U50002 ( .A(y[2174]), .B(x[2174]), .Z(n40825) );
  XOR U50003 ( .A(y[2173]), .B(x[2173]), .Z(n40826) );
  XOR U50004 ( .A(n40818), .B(n40817), .Z(n40827) );
  XOR U50005 ( .A(n40820), .B(n40819), .Z(n40817) );
  XOR U50006 ( .A(y[2171]), .B(x[2171]), .Z(n40819) );
  XOR U50007 ( .A(y[2170]), .B(x[2170]), .Z(n40820) );
  XOR U50008 ( .A(y[2169]), .B(x[2169]), .Z(n40818) );
  XNOR U50009 ( .A(n40811), .B(n40810), .Z(n40812) );
  XNOR U50010 ( .A(n40807), .B(n40806), .Z(n40810) );
  XOR U50011 ( .A(n40809), .B(n40808), .Z(n40806) );
  XOR U50012 ( .A(y[2168]), .B(x[2168]), .Z(n40808) );
  XOR U50013 ( .A(y[2167]), .B(x[2167]), .Z(n40809) );
  XOR U50014 ( .A(y[2166]), .B(x[2166]), .Z(n40807) );
  XOR U50015 ( .A(n40801), .B(n40800), .Z(n40811) );
  XOR U50016 ( .A(n40803), .B(n40802), .Z(n40800) );
  XOR U50017 ( .A(y[2165]), .B(x[2165]), .Z(n40802) );
  XOR U50018 ( .A(y[2164]), .B(x[2164]), .Z(n40803) );
  XOR U50019 ( .A(y[2163]), .B(x[2163]), .Z(n40801) );
  XNOR U50020 ( .A(n40777), .B(n40778), .Z(n40795) );
  XNOR U50021 ( .A(n40792), .B(n40793), .Z(n40778) );
  XOR U50022 ( .A(n40789), .B(n40788), .Z(n40793) );
  XOR U50023 ( .A(y[2160]), .B(x[2160]), .Z(n40788) );
  XOR U50024 ( .A(n40791), .B(n40790), .Z(n40789) );
  XOR U50025 ( .A(y[2162]), .B(x[2162]), .Z(n40790) );
  XOR U50026 ( .A(y[2161]), .B(x[2161]), .Z(n40791) );
  XOR U50027 ( .A(n40783), .B(n40782), .Z(n40792) );
  XOR U50028 ( .A(n40785), .B(n40784), .Z(n40782) );
  XOR U50029 ( .A(y[2159]), .B(x[2159]), .Z(n40784) );
  XOR U50030 ( .A(y[2158]), .B(x[2158]), .Z(n40785) );
  XOR U50031 ( .A(y[2157]), .B(x[2157]), .Z(n40783) );
  XNOR U50032 ( .A(n40776), .B(n40775), .Z(n40777) );
  XNOR U50033 ( .A(n40772), .B(n40771), .Z(n40775) );
  XOR U50034 ( .A(n40774), .B(n40773), .Z(n40771) );
  XOR U50035 ( .A(y[2156]), .B(x[2156]), .Z(n40773) );
  XOR U50036 ( .A(y[2155]), .B(x[2155]), .Z(n40774) );
  XOR U50037 ( .A(y[2154]), .B(x[2154]), .Z(n40772) );
  XOR U50038 ( .A(n40766), .B(n40765), .Z(n40776) );
  XOR U50039 ( .A(n40768), .B(n40767), .Z(n40765) );
  XOR U50040 ( .A(y[2153]), .B(x[2153]), .Z(n40767) );
  XOR U50041 ( .A(y[2152]), .B(x[2152]), .Z(n40768) );
  XOR U50042 ( .A(y[2151]), .B(x[2151]), .Z(n40766) );
  NAND U50043 ( .A(n40829), .B(n40830), .Z(N61753) );
  NAND U50044 ( .A(n40831), .B(n40832), .Z(n40830) );
  NANDN U50045 ( .A(n40833), .B(n40834), .Z(n40832) );
  NANDN U50046 ( .A(n40834), .B(n40833), .Z(n40829) );
  XOR U50047 ( .A(n40833), .B(n40835), .Z(N61752) );
  XNOR U50048 ( .A(n40831), .B(n40834), .Z(n40835) );
  NAND U50049 ( .A(n40836), .B(n40837), .Z(n40834) );
  NAND U50050 ( .A(n40838), .B(n40839), .Z(n40837) );
  NANDN U50051 ( .A(n40840), .B(n40841), .Z(n40839) );
  NANDN U50052 ( .A(n40841), .B(n40840), .Z(n40836) );
  AND U50053 ( .A(n40842), .B(n40843), .Z(n40831) );
  NAND U50054 ( .A(n40844), .B(n40845), .Z(n40843) );
  NANDN U50055 ( .A(n40846), .B(n40847), .Z(n40845) );
  NANDN U50056 ( .A(n40847), .B(n40846), .Z(n40842) );
  IV U50057 ( .A(n40848), .Z(n40847) );
  AND U50058 ( .A(n40849), .B(n40850), .Z(n40833) );
  NAND U50059 ( .A(n40851), .B(n40852), .Z(n40850) );
  NANDN U50060 ( .A(n40853), .B(n40854), .Z(n40852) );
  NANDN U50061 ( .A(n40854), .B(n40853), .Z(n40849) );
  XOR U50062 ( .A(n40846), .B(n40855), .Z(N61751) );
  XNOR U50063 ( .A(n40844), .B(n40848), .Z(n40855) );
  XOR U50064 ( .A(n40841), .B(n40856), .Z(n40848) );
  XNOR U50065 ( .A(n40838), .B(n40840), .Z(n40856) );
  AND U50066 ( .A(n40857), .B(n40858), .Z(n40840) );
  NANDN U50067 ( .A(n40859), .B(n40860), .Z(n40858) );
  OR U50068 ( .A(n40861), .B(n40862), .Z(n40860) );
  IV U50069 ( .A(n40863), .Z(n40862) );
  NANDN U50070 ( .A(n40863), .B(n40861), .Z(n40857) );
  AND U50071 ( .A(n40864), .B(n40865), .Z(n40838) );
  NAND U50072 ( .A(n40866), .B(n40867), .Z(n40865) );
  NANDN U50073 ( .A(n40868), .B(n40869), .Z(n40867) );
  NANDN U50074 ( .A(n40869), .B(n40868), .Z(n40864) );
  IV U50075 ( .A(n40870), .Z(n40869) );
  NAND U50076 ( .A(n40871), .B(n40872), .Z(n40841) );
  NANDN U50077 ( .A(n40873), .B(n40874), .Z(n40872) );
  NANDN U50078 ( .A(n40875), .B(n40876), .Z(n40874) );
  NANDN U50079 ( .A(n40876), .B(n40875), .Z(n40871) );
  IV U50080 ( .A(n40877), .Z(n40875) );
  AND U50081 ( .A(n40878), .B(n40879), .Z(n40844) );
  NAND U50082 ( .A(n40880), .B(n40881), .Z(n40879) );
  NANDN U50083 ( .A(n40882), .B(n40883), .Z(n40881) );
  NANDN U50084 ( .A(n40883), .B(n40882), .Z(n40878) );
  XOR U50085 ( .A(n40854), .B(n40884), .Z(n40846) );
  XNOR U50086 ( .A(n40851), .B(n40853), .Z(n40884) );
  AND U50087 ( .A(n40885), .B(n40886), .Z(n40853) );
  NANDN U50088 ( .A(n40887), .B(n40888), .Z(n40886) );
  OR U50089 ( .A(n40889), .B(n40890), .Z(n40888) );
  IV U50090 ( .A(n40891), .Z(n40890) );
  NANDN U50091 ( .A(n40891), .B(n40889), .Z(n40885) );
  AND U50092 ( .A(n40892), .B(n40893), .Z(n40851) );
  NAND U50093 ( .A(n40894), .B(n40895), .Z(n40893) );
  NANDN U50094 ( .A(n40896), .B(n40897), .Z(n40895) );
  NANDN U50095 ( .A(n40897), .B(n40896), .Z(n40892) );
  IV U50096 ( .A(n40898), .Z(n40897) );
  NAND U50097 ( .A(n40899), .B(n40900), .Z(n40854) );
  NANDN U50098 ( .A(n40901), .B(n40902), .Z(n40900) );
  NANDN U50099 ( .A(n40903), .B(n40904), .Z(n40902) );
  NANDN U50100 ( .A(n40904), .B(n40903), .Z(n40899) );
  IV U50101 ( .A(n40905), .Z(n40903) );
  XOR U50102 ( .A(n40880), .B(n40906), .Z(N61750) );
  XNOR U50103 ( .A(n40883), .B(n40882), .Z(n40906) );
  XNOR U50104 ( .A(n40894), .B(n40907), .Z(n40882) );
  XNOR U50105 ( .A(n40898), .B(n40896), .Z(n40907) );
  XOR U50106 ( .A(n40904), .B(n40908), .Z(n40896) );
  XNOR U50107 ( .A(n40901), .B(n40905), .Z(n40908) );
  AND U50108 ( .A(n40909), .B(n40910), .Z(n40905) );
  NAND U50109 ( .A(n40911), .B(n40912), .Z(n40910) );
  NAND U50110 ( .A(n40913), .B(n40914), .Z(n40909) );
  AND U50111 ( .A(n40915), .B(n40916), .Z(n40901) );
  NAND U50112 ( .A(n40917), .B(n40918), .Z(n40916) );
  NAND U50113 ( .A(n40919), .B(n40920), .Z(n40915) );
  NANDN U50114 ( .A(n40921), .B(n40922), .Z(n40904) );
  ANDN U50115 ( .B(n40923), .A(n40924), .Z(n40898) );
  XNOR U50116 ( .A(n40889), .B(n40925), .Z(n40894) );
  XNOR U50117 ( .A(n40887), .B(n40891), .Z(n40925) );
  AND U50118 ( .A(n40926), .B(n40927), .Z(n40891) );
  NAND U50119 ( .A(n40928), .B(n40929), .Z(n40927) );
  NAND U50120 ( .A(n40930), .B(n40931), .Z(n40926) );
  AND U50121 ( .A(n40932), .B(n40933), .Z(n40887) );
  NAND U50122 ( .A(n40934), .B(n40935), .Z(n40933) );
  NAND U50123 ( .A(n40936), .B(n40937), .Z(n40932) );
  AND U50124 ( .A(n40938), .B(n40939), .Z(n40889) );
  NAND U50125 ( .A(n40940), .B(n40941), .Z(n40883) );
  XNOR U50126 ( .A(n40866), .B(n40942), .Z(n40880) );
  XNOR U50127 ( .A(n40870), .B(n40868), .Z(n40942) );
  XOR U50128 ( .A(n40876), .B(n40943), .Z(n40868) );
  XNOR U50129 ( .A(n40873), .B(n40877), .Z(n40943) );
  AND U50130 ( .A(n40944), .B(n40945), .Z(n40877) );
  NAND U50131 ( .A(n40946), .B(n40947), .Z(n40945) );
  NAND U50132 ( .A(n40948), .B(n40949), .Z(n40944) );
  AND U50133 ( .A(n40950), .B(n40951), .Z(n40873) );
  NAND U50134 ( .A(n40952), .B(n40953), .Z(n40951) );
  NAND U50135 ( .A(n40954), .B(n40955), .Z(n40950) );
  NANDN U50136 ( .A(n40956), .B(n40957), .Z(n40876) );
  ANDN U50137 ( .B(n40958), .A(n40959), .Z(n40870) );
  XNOR U50138 ( .A(n40861), .B(n40960), .Z(n40866) );
  XNOR U50139 ( .A(n40859), .B(n40863), .Z(n40960) );
  AND U50140 ( .A(n40961), .B(n40962), .Z(n40863) );
  NAND U50141 ( .A(n40963), .B(n40964), .Z(n40962) );
  NAND U50142 ( .A(n40965), .B(n40966), .Z(n40961) );
  AND U50143 ( .A(n40967), .B(n40968), .Z(n40859) );
  NAND U50144 ( .A(n40969), .B(n40970), .Z(n40968) );
  NAND U50145 ( .A(n40971), .B(n40972), .Z(n40967) );
  AND U50146 ( .A(n40973), .B(n40974), .Z(n40861) );
  XOR U50147 ( .A(n40941), .B(n40940), .Z(N61749) );
  XNOR U50148 ( .A(n40958), .B(n40959), .Z(n40940) );
  XNOR U50149 ( .A(n40973), .B(n40974), .Z(n40959) );
  XOR U50150 ( .A(n40970), .B(n40969), .Z(n40974) );
  XOR U50151 ( .A(y[2148]), .B(x[2148]), .Z(n40969) );
  XOR U50152 ( .A(n40972), .B(n40971), .Z(n40970) );
  XOR U50153 ( .A(y[2150]), .B(x[2150]), .Z(n40971) );
  XOR U50154 ( .A(y[2149]), .B(x[2149]), .Z(n40972) );
  XOR U50155 ( .A(n40964), .B(n40963), .Z(n40973) );
  XOR U50156 ( .A(n40966), .B(n40965), .Z(n40963) );
  XOR U50157 ( .A(y[2147]), .B(x[2147]), .Z(n40965) );
  XOR U50158 ( .A(y[2146]), .B(x[2146]), .Z(n40966) );
  XOR U50159 ( .A(y[2145]), .B(x[2145]), .Z(n40964) );
  XNOR U50160 ( .A(n40957), .B(n40956), .Z(n40958) );
  XNOR U50161 ( .A(n40953), .B(n40952), .Z(n40956) );
  XOR U50162 ( .A(n40955), .B(n40954), .Z(n40952) );
  XOR U50163 ( .A(y[2144]), .B(x[2144]), .Z(n40954) );
  XOR U50164 ( .A(y[2143]), .B(x[2143]), .Z(n40955) );
  XOR U50165 ( .A(y[2142]), .B(x[2142]), .Z(n40953) );
  XOR U50166 ( .A(n40947), .B(n40946), .Z(n40957) );
  XOR U50167 ( .A(n40949), .B(n40948), .Z(n40946) );
  XOR U50168 ( .A(y[2141]), .B(x[2141]), .Z(n40948) );
  XOR U50169 ( .A(y[2140]), .B(x[2140]), .Z(n40949) );
  XOR U50170 ( .A(y[2139]), .B(x[2139]), .Z(n40947) );
  XNOR U50171 ( .A(n40923), .B(n40924), .Z(n40941) );
  XNOR U50172 ( .A(n40938), .B(n40939), .Z(n40924) );
  XOR U50173 ( .A(n40935), .B(n40934), .Z(n40939) );
  XOR U50174 ( .A(y[2136]), .B(x[2136]), .Z(n40934) );
  XOR U50175 ( .A(n40937), .B(n40936), .Z(n40935) );
  XOR U50176 ( .A(y[2138]), .B(x[2138]), .Z(n40936) );
  XOR U50177 ( .A(y[2137]), .B(x[2137]), .Z(n40937) );
  XOR U50178 ( .A(n40929), .B(n40928), .Z(n40938) );
  XOR U50179 ( .A(n40931), .B(n40930), .Z(n40928) );
  XOR U50180 ( .A(y[2135]), .B(x[2135]), .Z(n40930) );
  XOR U50181 ( .A(y[2134]), .B(x[2134]), .Z(n40931) );
  XOR U50182 ( .A(y[2133]), .B(x[2133]), .Z(n40929) );
  XNOR U50183 ( .A(n40922), .B(n40921), .Z(n40923) );
  XNOR U50184 ( .A(n40918), .B(n40917), .Z(n40921) );
  XOR U50185 ( .A(n40920), .B(n40919), .Z(n40917) );
  XOR U50186 ( .A(y[2132]), .B(x[2132]), .Z(n40919) );
  XOR U50187 ( .A(y[2131]), .B(x[2131]), .Z(n40920) );
  XOR U50188 ( .A(y[2130]), .B(x[2130]), .Z(n40918) );
  XOR U50189 ( .A(n40912), .B(n40911), .Z(n40922) );
  XOR U50190 ( .A(n40914), .B(n40913), .Z(n40911) );
  XOR U50191 ( .A(y[2129]), .B(x[2129]), .Z(n40913) );
  XOR U50192 ( .A(y[2128]), .B(x[2128]), .Z(n40914) );
  XOR U50193 ( .A(y[2127]), .B(x[2127]), .Z(n40912) );
  NAND U50194 ( .A(n40975), .B(n40976), .Z(N61740) );
  NAND U50195 ( .A(n40977), .B(n40978), .Z(n40976) );
  NANDN U50196 ( .A(n40979), .B(n40980), .Z(n40978) );
  NANDN U50197 ( .A(n40980), .B(n40979), .Z(n40975) );
  XOR U50198 ( .A(n40979), .B(n40981), .Z(N61739) );
  XNOR U50199 ( .A(n40977), .B(n40980), .Z(n40981) );
  NAND U50200 ( .A(n40982), .B(n40983), .Z(n40980) );
  NAND U50201 ( .A(n40984), .B(n40985), .Z(n40983) );
  NANDN U50202 ( .A(n40986), .B(n40987), .Z(n40985) );
  NANDN U50203 ( .A(n40987), .B(n40986), .Z(n40982) );
  AND U50204 ( .A(n40988), .B(n40989), .Z(n40977) );
  NAND U50205 ( .A(n40990), .B(n40991), .Z(n40989) );
  NANDN U50206 ( .A(n40992), .B(n40993), .Z(n40991) );
  NANDN U50207 ( .A(n40993), .B(n40992), .Z(n40988) );
  IV U50208 ( .A(n40994), .Z(n40993) );
  AND U50209 ( .A(n40995), .B(n40996), .Z(n40979) );
  NAND U50210 ( .A(n40997), .B(n40998), .Z(n40996) );
  NANDN U50211 ( .A(n40999), .B(n41000), .Z(n40998) );
  NANDN U50212 ( .A(n41000), .B(n40999), .Z(n40995) );
  XOR U50213 ( .A(n40992), .B(n41001), .Z(N61738) );
  XNOR U50214 ( .A(n40990), .B(n40994), .Z(n41001) );
  XOR U50215 ( .A(n40987), .B(n41002), .Z(n40994) );
  XNOR U50216 ( .A(n40984), .B(n40986), .Z(n41002) );
  AND U50217 ( .A(n41003), .B(n41004), .Z(n40986) );
  NANDN U50218 ( .A(n41005), .B(n41006), .Z(n41004) );
  OR U50219 ( .A(n41007), .B(n41008), .Z(n41006) );
  IV U50220 ( .A(n41009), .Z(n41008) );
  NANDN U50221 ( .A(n41009), .B(n41007), .Z(n41003) );
  AND U50222 ( .A(n41010), .B(n41011), .Z(n40984) );
  NAND U50223 ( .A(n41012), .B(n41013), .Z(n41011) );
  NANDN U50224 ( .A(n41014), .B(n41015), .Z(n41013) );
  NANDN U50225 ( .A(n41015), .B(n41014), .Z(n41010) );
  IV U50226 ( .A(n41016), .Z(n41015) );
  NAND U50227 ( .A(n41017), .B(n41018), .Z(n40987) );
  NANDN U50228 ( .A(n41019), .B(n41020), .Z(n41018) );
  NANDN U50229 ( .A(n41021), .B(n41022), .Z(n41020) );
  NANDN U50230 ( .A(n41022), .B(n41021), .Z(n41017) );
  IV U50231 ( .A(n41023), .Z(n41021) );
  AND U50232 ( .A(n41024), .B(n41025), .Z(n40990) );
  NAND U50233 ( .A(n41026), .B(n41027), .Z(n41025) );
  NANDN U50234 ( .A(n41028), .B(n41029), .Z(n41027) );
  NANDN U50235 ( .A(n41029), .B(n41028), .Z(n41024) );
  XOR U50236 ( .A(n41000), .B(n41030), .Z(n40992) );
  XNOR U50237 ( .A(n40997), .B(n40999), .Z(n41030) );
  AND U50238 ( .A(n41031), .B(n41032), .Z(n40999) );
  NANDN U50239 ( .A(n41033), .B(n41034), .Z(n41032) );
  OR U50240 ( .A(n41035), .B(n41036), .Z(n41034) );
  IV U50241 ( .A(n41037), .Z(n41036) );
  NANDN U50242 ( .A(n41037), .B(n41035), .Z(n41031) );
  AND U50243 ( .A(n41038), .B(n41039), .Z(n40997) );
  NAND U50244 ( .A(n41040), .B(n41041), .Z(n41039) );
  NANDN U50245 ( .A(n41042), .B(n41043), .Z(n41041) );
  NANDN U50246 ( .A(n41043), .B(n41042), .Z(n41038) );
  IV U50247 ( .A(n41044), .Z(n41043) );
  NAND U50248 ( .A(n41045), .B(n41046), .Z(n41000) );
  NANDN U50249 ( .A(n41047), .B(n41048), .Z(n41046) );
  NANDN U50250 ( .A(n41049), .B(n41050), .Z(n41048) );
  NANDN U50251 ( .A(n41050), .B(n41049), .Z(n41045) );
  IV U50252 ( .A(n41051), .Z(n41049) );
  XOR U50253 ( .A(n41026), .B(n41052), .Z(N61737) );
  XNOR U50254 ( .A(n41029), .B(n41028), .Z(n41052) );
  XNOR U50255 ( .A(n41040), .B(n41053), .Z(n41028) );
  XNOR U50256 ( .A(n41044), .B(n41042), .Z(n41053) );
  XOR U50257 ( .A(n41050), .B(n41054), .Z(n41042) );
  XNOR U50258 ( .A(n41047), .B(n41051), .Z(n41054) );
  AND U50259 ( .A(n41055), .B(n41056), .Z(n41051) );
  NAND U50260 ( .A(n41057), .B(n41058), .Z(n41056) );
  NAND U50261 ( .A(n41059), .B(n41060), .Z(n41055) );
  AND U50262 ( .A(n41061), .B(n41062), .Z(n41047) );
  NAND U50263 ( .A(n41063), .B(n41064), .Z(n41062) );
  NAND U50264 ( .A(n41065), .B(n41066), .Z(n41061) );
  NANDN U50265 ( .A(n41067), .B(n41068), .Z(n41050) );
  ANDN U50266 ( .B(n41069), .A(n41070), .Z(n41044) );
  XNOR U50267 ( .A(n41035), .B(n41071), .Z(n41040) );
  XNOR U50268 ( .A(n41033), .B(n41037), .Z(n41071) );
  AND U50269 ( .A(n41072), .B(n41073), .Z(n41037) );
  NAND U50270 ( .A(n41074), .B(n41075), .Z(n41073) );
  NAND U50271 ( .A(n41076), .B(n41077), .Z(n41072) );
  AND U50272 ( .A(n41078), .B(n41079), .Z(n41033) );
  NAND U50273 ( .A(n41080), .B(n41081), .Z(n41079) );
  NAND U50274 ( .A(n41082), .B(n41083), .Z(n41078) );
  AND U50275 ( .A(n41084), .B(n41085), .Z(n41035) );
  NAND U50276 ( .A(n41086), .B(n41087), .Z(n41029) );
  XNOR U50277 ( .A(n41012), .B(n41088), .Z(n41026) );
  XNOR U50278 ( .A(n41016), .B(n41014), .Z(n41088) );
  XOR U50279 ( .A(n41022), .B(n41089), .Z(n41014) );
  XNOR U50280 ( .A(n41019), .B(n41023), .Z(n41089) );
  AND U50281 ( .A(n41090), .B(n41091), .Z(n41023) );
  NAND U50282 ( .A(n41092), .B(n41093), .Z(n41091) );
  NAND U50283 ( .A(n41094), .B(n41095), .Z(n41090) );
  AND U50284 ( .A(n41096), .B(n41097), .Z(n41019) );
  NAND U50285 ( .A(n41098), .B(n41099), .Z(n41097) );
  NAND U50286 ( .A(n41100), .B(n41101), .Z(n41096) );
  NANDN U50287 ( .A(n41102), .B(n41103), .Z(n41022) );
  ANDN U50288 ( .B(n41104), .A(n41105), .Z(n41016) );
  XNOR U50289 ( .A(n41007), .B(n41106), .Z(n41012) );
  XNOR U50290 ( .A(n41005), .B(n41009), .Z(n41106) );
  AND U50291 ( .A(n41107), .B(n41108), .Z(n41009) );
  NAND U50292 ( .A(n41109), .B(n41110), .Z(n41108) );
  NAND U50293 ( .A(n41111), .B(n41112), .Z(n41107) );
  AND U50294 ( .A(n41113), .B(n41114), .Z(n41005) );
  NAND U50295 ( .A(n41115), .B(n41116), .Z(n41114) );
  NAND U50296 ( .A(n41117), .B(n41118), .Z(n41113) );
  AND U50297 ( .A(n41119), .B(n41120), .Z(n41007) );
  XOR U50298 ( .A(n41087), .B(n41086), .Z(N61736) );
  XNOR U50299 ( .A(n41104), .B(n41105), .Z(n41086) );
  XNOR U50300 ( .A(n41119), .B(n41120), .Z(n41105) );
  XOR U50301 ( .A(n41116), .B(n41115), .Z(n41120) );
  XOR U50302 ( .A(y[2124]), .B(x[2124]), .Z(n41115) );
  XOR U50303 ( .A(n41118), .B(n41117), .Z(n41116) );
  XOR U50304 ( .A(y[2126]), .B(x[2126]), .Z(n41117) );
  XOR U50305 ( .A(y[2125]), .B(x[2125]), .Z(n41118) );
  XOR U50306 ( .A(n41110), .B(n41109), .Z(n41119) );
  XOR U50307 ( .A(n41112), .B(n41111), .Z(n41109) );
  XOR U50308 ( .A(y[2123]), .B(x[2123]), .Z(n41111) );
  XOR U50309 ( .A(y[2122]), .B(x[2122]), .Z(n41112) );
  XOR U50310 ( .A(y[2121]), .B(x[2121]), .Z(n41110) );
  XNOR U50311 ( .A(n41103), .B(n41102), .Z(n41104) );
  XNOR U50312 ( .A(n41099), .B(n41098), .Z(n41102) );
  XOR U50313 ( .A(n41101), .B(n41100), .Z(n41098) );
  XOR U50314 ( .A(y[2120]), .B(x[2120]), .Z(n41100) );
  XOR U50315 ( .A(y[2119]), .B(x[2119]), .Z(n41101) );
  XOR U50316 ( .A(y[2118]), .B(x[2118]), .Z(n41099) );
  XOR U50317 ( .A(n41093), .B(n41092), .Z(n41103) );
  XOR U50318 ( .A(n41095), .B(n41094), .Z(n41092) );
  XOR U50319 ( .A(y[2117]), .B(x[2117]), .Z(n41094) );
  XOR U50320 ( .A(y[2116]), .B(x[2116]), .Z(n41095) );
  XOR U50321 ( .A(y[2115]), .B(x[2115]), .Z(n41093) );
  XNOR U50322 ( .A(n41069), .B(n41070), .Z(n41087) );
  XNOR U50323 ( .A(n41084), .B(n41085), .Z(n41070) );
  XOR U50324 ( .A(n41081), .B(n41080), .Z(n41085) );
  XOR U50325 ( .A(y[2112]), .B(x[2112]), .Z(n41080) );
  XOR U50326 ( .A(n41083), .B(n41082), .Z(n41081) );
  XOR U50327 ( .A(y[2114]), .B(x[2114]), .Z(n41082) );
  XOR U50328 ( .A(y[2113]), .B(x[2113]), .Z(n41083) );
  XOR U50329 ( .A(n41075), .B(n41074), .Z(n41084) );
  XOR U50330 ( .A(n41077), .B(n41076), .Z(n41074) );
  XOR U50331 ( .A(y[2111]), .B(x[2111]), .Z(n41076) );
  XOR U50332 ( .A(y[2110]), .B(x[2110]), .Z(n41077) );
  XOR U50333 ( .A(y[2109]), .B(x[2109]), .Z(n41075) );
  XNOR U50334 ( .A(n41068), .B(n41067), .Z(n41069) );
  XNOR U50335 ( .A(n41064), .B(n41063), .Z(n41067) );
  XOR U50336 ( .A(n41066), .B(n41065), .Z(n41063) );
  XOR U50337 ( .A(y[2108]), .B(x[2108]), .Z(n41065) );
  XOR U50338 ( .A(y[2107]), .B(x[2107]), .Z(n41066) );
  XOR U50339 ( .A(y[2106]), .B(x[2106]), .Z(n41064) );
  XOR U50340 ( .A(n41058), .B(n41057), .Z(n41068) );
  XOR U50341 ( .A(n41060), .B(n41059), .Z(n41057) );
  XOR U50342 ( .A(y[2105]), .B(x[2105]), .Z(n41059) );
  XOR U50343 ( .A(y[2104]), .B(x[2104]), .Z(n41060) );
  XOR U50344 ( .A(y[2103]), .B(x[2103]), .Z(n41058) );
  NAND U50345 ( .A(n41121), .B(n41122), .Z(N61727) );
  NAND U50346 ( .A(n41123), .B(n41124), .Z(n41122) );
  NANDN U50347 ( .A(n41125), .B(n41126), .Z(n41124) );
  NANDN U50348 ( .A(n41126), .B(n41125), .Z(n41121) );
  XOR U50349 ( .A(n41125), .B(n41127), .Z(N61726) );
  XNOR U50350 ( .A(n41123), .B(n41126), .Z(n41127) );
  NAND U50351 ( .A(n41128), .B(n41129), .Z(n41126) );
  NAND U50352 ( .A(n41130), .B(n41131), .Z(n41129) );
  NANDN U50353 ( .A(n41132), .B(n41133), .Z(n41131) );
  NANDN U50354 ( .A(n41133), .B(n41132), .Z(n41128) );
  AND U50355 ( .A(n41134), .B(n41135), .Z(n41123) );
  NAND U50356 ( .A(n41136), .B(n41137), .Z(n41135) );
  NANDN U50357 ( .A(n41138), .B(n41139), .Z(n41137) );
  NANDN U50358 ( .A(n41139), .B(n41138), .Z(n41134) );
  IV U50359 ( .A(n41140), .Z(n41139) );
  AND U50360 ( .A(n41141), .B(n41142), .Z(n41125) );
  NAND U50361 ( .A(n41143), .B(n41144), .Z(n41142) );
  NANDN U50362 ( .A(n41145), .B(n41146), .Z(n41144) );
  NANDN U50363 ( .A(n41146), .B(n41145), .Z(n41141) );
  XOR U50364 ( .A(n41138), .B(n41147), .Z(N61725) );
  XNOR U50365 ( .A(n41136), .B(n41140), .Z(n41147) );
  XOR U50366 ( .A(n41133), .B(n41148), .Z(n41140) );
  XNOR U50367 ( .A(n41130), .B(n41132), .Z(n41148) );
  AND U50368 ( .A(n41149), .B(n41150), .Z(n41132) );
  NANDN U50369 ( .A(n41151), .B(n41152), .Z(n41150) );
  OR U50370 ( .A(n41153), .B(n41154), .Z(n41152) );
  IV U50371 ( .A(n41155), .Z(n41154) );
  NANDN U50372 ( .A(n41155), .B(n41153), .Z(n41149) );
  AND U50373 ( .A(n41156), .B(n41157), .Z(n41130) );
  NAND U50374 ( .A(n41158), .B(n41159), .Z(n41157) );
  NANDN U50375 ( .A(n41160), .B(n41161), .Z(n41159) );
  NANDN U50376 ( .A(n41161), .B(n41160), .Z(n41156) );
  IV U50377 ( .A(n41162), .Z(n41161) );
  NAND U50378 ( .A(n41163), .B(n41164), .Z(n41133) );
  NANDN U50379 ( .A(n41165), .B(n41166), .Z(n41164) );
  NANDN U50380 ( .A(n41167), .B(n41168), .Z(n41166) );
  NANDN U50381 ( .A(n41168), .B(n41167), .Z(n41163) );
  IV U50382 ( .A(n41169), .Z(n41167) );
  AND U50383 ( .A(n41170), .B(n41171), .Z(n41136) );
  NAND U50384 ( .A(n41172), .B(n41173), .Z(n41171) );
  NANDN U50385 ( .A(n41174), .B(n41175), .Z(n41173) );
  NANDN U50386 ( .A(n41175), .B(n41174), .Z(n41170) );
  XOR U50387 ( .A(n41146), .B(n41176), .Z(n41138) );
  XNOR U50388 ( .A(n41143), .B(n41145), .Z(n41176) );
  AND U50389 ( .A(n41177), .B(n41178), .Z(n41145) );
  NANDN U50390 ( .A(n41179), .B(n41180), .Z(n41178) );
  OR U50391 ( .A(n41181), .B(n41182), .Z(n41180) );
  IV U50392 ( .A(n41183), .Z(n41182) );
  NANDN U50393 ( .A(n41183), .B(n41181), .Z(n41177) );
  AND U50394 ( .A(n41184), .B(n41185), .Z(n41143) );
  NAND U50395 ( .A(n41186), .B(n41187), .Z(n41185) );
  NANDN U50396 ( .A(n41188), .B(n41189), .Z(n41187) );
  NANDN U50397 ( .A(n41189), .B(n41188), .Z(n41184) );
  IV U50398 ( .A(n41190), .Z(n41189) );
  NAND U50399 ( .A(n41191), .B(n41192), .Z(n41146) );
  NANDN U50400 ( .A(n41193), .B(n41194), .Z(n41192) );
  NANDN U50401 ( .A(n41195), .B(n41196), .Z(n41194) );
  NANDN U50402 ( .A(n41196), .B(n41195), .Z(n41191) );
  IV U50403 ( .A(n41197), .Z(n41195) );
  XOR U50404 ( .A(n41172), .B(n41198), .Z(N61724) );
  XNOR U50405 ( .A(n41175), .B(n41174), .Z(n41198) );
  XNOR U50406 ( .A(n41186), .B(n41199), .Z(n41174) );
  XNOR U50407 ( .A(n41190), .B(n41188), .Z(n41199) );
  XOR U50408 ( .A(n41196), .B(n41200), .Z(n41188) );
  XNOR U50409 ( .A(n41193), .B(n41197), .Z(n41200) );
  AND U50410 ( .A(n41201), .B(n41202), .Z(n41197) );
  NAND U50411 ( .A(n41203), .B(n41204), .Z(n41202) );
  NAND U50412 ( .A(n41205), .B(n41206), .Z(n41201) );
  AND U50413 ( .A(n41207), .B(n41208), .Z(n41193) );
  NAND U50414 ( .A(n41209), .B(n41210), .Z(n41208) );
  NAND U50415 ( .A(n41211), .B(n41212), .Z(n41207) );
  NANDN U50416 ( .A(n41213), .B(n41214), .Z(n41196) );
  ANDN U50417 ( .B(n41215), .A(n41216), .Z(n41190) );
  XNOR U50418 ( .A(n41181), .B(n41217), .Z(n41186) );
  XNOR U50419 ( .A(n41179), .B(n41183), .Z(n41217) );
  AND U50420 ( .A(n41218), .B(n41219), .Z(n41183) );
  NAND U50421 ( .A(n41220), .B(n41221), .Z(n41219) );
  NAND U50422 ( .A(n41222), .B(n41223), .Z(n41218) );
  AND U50423 ( .A(n41224), .B(n41225), .Z(n41179) );
  NAND U50424 ( .A(n41226), .B(n41227), .Z(n41225) );
  NAND U50425 ( .A(n41228), .B(n41229), .Z(n41224) );
  AND U50426 ( .A(n41230), .B(n41231), .Z(n41181) );
  NAND U50427 ( .A(n41232), .B(n41233), .Z(n41175) );
  XNOR U50428 ( .A(n41158), .B(n41234), .Z(n41172) );
  XNOR U50429 ( .A(n41162), .B(n41160), .Z(n41234) );
  XOR U50430 ( .A(n41168), .B(n41235), .Z(n41160) );
  XNOR U50431 ( .A(n41165), .B(n41169), .Z(n41235) );
  AND U50432 ( .A(n41236), .B(n41237), .Z(n41169) );
  NAND U50433 ( .A(n41238), .B(n41239), .Z(n41237) );
  NAND U50434 ( .A(n41240), .B(n41241), .Z(n41236) );
  AND U50435 ( .A(n41242), .B(n41243), .Z(n41165) );
  NAND U50436 ( .A(n41244), .B(n41245), .Z(n41243) );
  NAND U50437 ( .A(n41246), .B(n41247), .Z(n41242) );
  NANDN U50438 ( .A(n41248), .B(n41249), .Z(n41168) );
  ANDN U50439 ( .B(n41250), .A(n41251), .Z(n41162) );
  XNOR U50440 ( .A(n41153), .B(n41252), .Z(n41158) );
  XNOR U50441 ( .A(n41151), .B(n41155), .Z(n41252) );
  AND U50442 ( .A(n41253), .B(n41254), .Z(n41155) );
  NAND U50443 ( .A(n41255), .B(n41256), .Z(n41254) );
  NAND U50444 ( .A(n41257), .B(n41258), .Z(n41253) );
  AND U50445 ( .A(n41259), .B(n41260), .Z(n41151) );
  NAND U50446 ( .A(n41261), .B(n41262), .Z(n41260) );
  NAND U50447 ( .A(n41263), .B(n41264), .Z(n41259) );
  AND U50448 ( .A(n41265), .B(n41266), .Z(n41153) );
  XOR U50449 ( .A(n41233), .B(n41232), .Z(N61723) );
  XNOR U50450 ( .A(n41250), .B(n41251), .Z(n41232) );
  XNOR U50451 ( .A(n41265), .B(n41266), .Z(n41251) );
  XOR U50452 ( .A(n41262), .B(n41261), .Z(n41266) );
  XOR U50453 ( .A(y[2100]), .B(x[2100]), .Z(n41261) );
  XOR U50454 ( .A(n41264), .B(n41263), .Z(n41262) );
  XOR U50455 ( .A(y[2102]), .B(x[2102]), .Z(n41263) );
  XOR U50456 ( .A(y[2101]), .B(x[2101]), .Z(n41264) );
  XOR U50457 ( .A(n41256), .B(n41255), .Z(n41265) );
  XOR U50458 ( .A(n41258), .B(n41257), .Z(n41255) );
  XOR U50459 ( .A(y[2099]), .B(x[2099]), .Z(n41257) );
  XOR U50460 ( .A(y[2098]), .B(x[2098]), .Z(n41258) );
  XOR U50461 ( .A(y[2097]), .B(x[2097]), .Z(n41256) );
  XNOR U50462 ( .A(n41249), .B(n41248), .Z(n41250) );
  XNOR U50463 ( .A(n41245), .B(n41244), .Z(n41248) );
  XOR U50464 ( .A(n41247), .B(n41246), .Z(n41244) );
  XOR U50465 ( .A(y[2096]), .B(x[2096]), .Z(n41246) );
  XOR U50466 ( .A(y[2095]), .B(x[2095]), .Z(n41247) );
  XOR U50467 ( .A(y[2094]), .B(x[2094]), .Z(n41245) );
  XOR U50468 ( .A(n41239), .B(n41238), .Z(n41249) );
  XOR U50469 ( .A(n41241), .B(n41240), .Z(n41238) );
  XOR U50470 ( .A(y[2093]), .B(x[2093]), .Z(n41240) );
  XOR U50471 ( .A(y[2092]), .B(x[2092]), .Z(n41241) );
  XOR U50472 ( .A(y[2091]), .B(x[2091]), .Z(n41239) );
  XNOR U50473 ( .A(n41215), .B(n41216), .Z(n41233) );
  XNOR U50474 ( .A(n41230), .B(n41231), .Z(n41216) );
  XOR U50475 ( .A(n41227), .B(n41226), .Z(n41231) );
  XOR U50476 ( .A(y[2088]), .B(x[2088]), .Z(n41226) );
  XOR U50477 ( .A(n41229), .B(n41228), .Z(n41227) );
  XOR U50478 ( .A(y[2090]), .B(x[2090]), .Z(n41228) );
  XOR U50479 ( .A(y[2089]), .B(x[2089]), .Z(n41229) );
  XOR U50480 ( .A(n41221), .B(n41220), .Z(n41230) );
  XOR U50481 ( .A(n41223), .B(n41222), .Z(n41220) );
  XOR U50482 ( .A(y[2087]), .B(x[2087]), .Z(n41222) );
  XOR U50483 ( .A(y[2086]), .B(x[2086]), .Z(n41223) );
  XOR U50484 ( .A(y[2085]), .B(x[2085]), .Z(n41221) );
  XNOR U50485 ( .A(n41214), .B(n41213), .Z(n41215) );
  XNOR U50486 ( .A(n41210), .B(n41209), .Z(n41213) );
  XOR U50487 ( .A(n41212), .B(n41211), .Z(n41209) );
  XOR U50488 ( .A(y[2084]), .B(x[2084]), .Z(n41211) );
  XOR U50489 ( .A(y[2083]), .B(x[2083]), .Z(n41212) );
  XOR U50490 ( .A(y[2082]), .B(x[2082]), .Z(n41210) );
  XOR U50491 ( .A(n41204), .B(n41203), .Z(n41214) );
  XOR U50492 ( .A(n41206), .B(n41205), .Z(n41203) );
  XOR U50493 ( .A(y[2081]), .B(x[2081]), .Z(n41205) );
  XOR U50494 ( .A(y[2080]), .B(x[2080]), .Z(n41206) );
  XOR U50495 ( .A(y[2079]), .B(x[2079]), .Z(n41204) );
  NAND U50496 ( .A(n41267), .B(n41268), .Z(N61714) );
  NAND U50497 ( .A(n41269), .B(n41270), .Z(n41268) );
  NANDN U50498 ( .A(n41271), .B(n41272), .Z(n41270) );
  NANDN U50499 ( .A(n41272), .B(n41271), .Z(n41267) );
  XOR U50500 ( .A(n41271), .B(n41273), .Z(N61713) );
  XNOR U50501 ( .A(n41269), .B(n41272), .Z(n41273) );
  NAND U50502 ( .A(n41274), .B(n41275), .Z(n41272) );
  NAND U50503 ( .A(n41276), .B(n41277), .Z(n41275) );
  NANDN U50504 ( .A(n41278), .B(n41279), .Z(n41277) );
  NANDN U50505 ( .A(n41279), .B(n41278), .Z(n41274) );
  AND U50506 ( .A(n41280), .B(n41281), .Z(n41269) );
  NAND U50507 ( .A(n41282), .B(n41283), .Z(n41281) );
  NANDN U50508 ( .A(n41284), .B(n41285), .Z(n41283) );
  NANDN U50509 ( .A(n41285), .B(n41284), .Z(n41280) );
  IV U50510 ( .A(n41286), .Z(n41285) );
  AND U50511 ( .A(n41287), .B(n41288), .Z(n41271) );
  NAND U50512 ( .A(n41289), .B(n41290), .Z(n41288) );
  NANDN U50513 ( .A(n41291), .B(n41292), .Z(n41290) );
  NANDN U50514 ( .A(n41292), .B(n41291), .Z(n41287) );
  XOR U50515 ( .A(n41284), .B(n41293), .Z(N61712) );
  XNOR U50516 ( .A(n41282), .B(n41286), .Z(n41293) );
  XOR U50517 ( .A(n41279), .B(n41294), .Z(n41286) );
  XNOR U50518 ( .A(n41276), .B(n41278), .Z(n41294) );
  AND U50519 ( .A(n41295), .B(n41296), .Z(n41278) );
  NANDN U50520 ( .A(n41297), .B(n41298), .Z(n41296) );
  OR U50521 ( .A(n41299), .B(n41300), .Z(n41298) );
  IV U50522 ( .A(n41301), .Z(n41300) );
  NANDN U50523 ( .A(n41301), .B(n41299), .Z(n41295) );
  AND U50524 ( .A(n41302), .B(n41303), .Z(n41276) );
  NAND U50525 ( .A(n41304), .B(n41305), .Z(n41303) );
  NANDN U50526 ( .A(n41306), .B(n41307), .Z(n41305) );
  NANDN U50527 ( .A(n41307), .B(n41306), .Z(n41302) );
  IV U50528 ( .A(n41308), .Z(n41307) );
  NAND U50529 ( .A(n41309), .B(n41310), .Z(n41279) );
  NANDN U50530 ( .A(n41311), .B(n41312), .Z(n41310) );
  NANDN U50531 ( .A(n41313), .B(n41314), .Z(n41312) );
  NANDN U50532 ( .A(n41314), .B(n41313), .Z(n41309) );
  IV U50533 ( .A(n41315), .Z(n41313) );
  AND U50534 ( .A(n41316), .B(n41317), .Z(n41282) );
  NAND U50535 ( .A(n41318), .B(n41319), .Z(n41317) );
  NANDN U50536 ( .A(n41320), .B(n41321), .Z(n41319) );
  NANDN U50537 ( .A(n41321), .B(n41320), .Z(n41316) );
  XOR U50538 ( .A(n41292), .B(n41322), .Z(n41284) );
  XNOR U50539 ( .A(n41289), .B(n41291), .Z(n41322) );
  AND U50540 ( .A(n41323), .B(n41324), .Z(n41291) );
  NANDN U50541 ( .A(n41325), .B(n41326), .Z(n41324) );
  OR U50542 ( .A(n41327), .B(n41328), .Z(n41326) );
  IV U50543 ( .A(n41329), .Z(n41328) );
  NANDN U50544 ( .A(n41329), .B(n41327), .Z(n41323) );
  AND U50545 ( .A(n41330), .B(n41331), .Z(n41289) );
  NAND U50546 ( .A(n41332), .B(n41333), .Z(n41331) );
  NANDN U50547 ( .A(n41334), .B(n41335), .Z(n41333) );
  NANDN U50548 ( .A(n41335), .B(n41334), .Z(n41330) );
  IV U50549 ( .A(n41336), .Z(n41335) );
  NAND U50550 ( .A(n41337), .B(n41338), .Z(n41292) );
  NANDN U50551 ( .A(n41339), .B(n41340), .Z(n41338) );
  NANDN U50552 ( .A(n41341), .B(n41342), .Z(n41340) );
  NANDN U50553 ( .A(n41342), .B(n41341), .Z(n41337) );
  IV U50554 ( .A(n41343), .Z(n41341) );
  XOR U50555 ( .A(n41318), .B(n41344), .Z(N61711) );
  XNOR U50556 ( .A(n41321), .B(n41320), .Z(n41344) );
  XNOR U50557 ( .A(n41332), .B(n41345), .Z(n41320) );
  XNOR U50558 ( .A(n41336), .B(n41334), .Z(n41345) );
  XOR U50559 ( .A(n41342), .B(n41346), .Z(n41334) );
  XNOR U50560 ( .A(n41339), .B(n41343), .Z(n41346) );
  AND U50561 ( .A(n41347), .B(n41348), .Z(n41343) );
  NAND U50562 ( .A(n41349), .B(n41350), .Z(n41348) );
  NAND U50563 ( .A(n41351), .B(n41352), .Z(n41347) );
  AND U50564 ( .A(n41353), .B(n41354), .Z(n41339) );
  NAND U50565 ( .A(n41355), .B(n41356), .Z(n41354) );
  NAND U50566 ( .A(n41357), .B(n41358), .Z(n41353) );
  NANDN U50567 ( .A(n41359), .B(n41360), .Z(n41342) );
  ANDN U50568 ( .B(n41361), .A(n41362), .Z(n41336) );
  XNOR U50569 ( .A(n41327), .B(n41363), .Z(n41332) );
  XNOR U50570 ( .A(n41325), .B(n41329), .Z(n41363) );
  AND U50571 ( .A(n41364), .B(n41365), .Z(n41329) );
  NAND U50572 ( .A(n41366), .B(n41367), .Z(n41365) );
  NAND U50573 ( .A(n41368), .B(n41369), .Z(n41364) );
  AND U50574 ( .A(n41370), .B(n41371), .Z(n41325) );
  NAND U50575 ( .A(n41372), .B(n41373), .Z(n41371) );
  NAND U50576 ( .A(n41374), .B(n41375), .Z(n41370) );
  AND U50577 ( .A(n41376), .B(n41377), .Z(n41327) );
  NAND U50578 ( .A(n41378), .B(n41379), .Z(n41321) );
  XNOR U50579 ( .A(n41304), .B(n41380), .Z(n41318) );
  XNOR U50580 ( .A(n41308), .B(n41306), .Z(n41380) );
  XOR U50581 ( .A(n41314), .B(n41381), .Z(n41306) );
  XNOR U50582 ( .A(n41311), .B(n41315), .Z(n41381) );
  AND U50583 ( .A(n41382), .B(n41383), .Z(n41315) );
  NAND U50584 ( .A(n41384), .B(n41385), .Z(n41383) );
  NAND U50585 ( .A(n41386), .B(n41387), .Z(n41382) );
  AND U50586 ( .A(n41388), .B(n41389), .Z(n41311) );
  NAND U50587 ( .A(n41390), .B(n41391), .Z(n41389) );
  NAND U50588 ( .A(n41392), .B(n41393), .Z(n41388) );
  NANDN U50589 ( .A(n41394), .B(n41395), .Z(n41314) );
  ANDN U50590 ( .B(n41396), .A(n41397), .Z(n41308) );
  XNOR U50591 ( .A(n41299), .B(n41398), .Z(n41304) );
  XNOR U50592 ( .A(n41297), .B(n41301), .Z(n41398) );
  AND U50593 ( .A(n41399), .B(n41400), .Z(n41301) );
  NAND U50594 ( .A(n41401), .B(n41402), .Z(n41400) );
  NAND U50595 ( .A(n41403), .B(n41404), .Z(n41399) );
  AND U50596 ( .A(n41405), .B(n41406), .Z(n41297) );
  NAND U50597 ( .A(n41407), .B(n41408), .Z(n41406) );
  NAND U50598 ( .A(n41409), .B(n41410), .Z(n41405) );
  AND U50599 ( .A(n41411), .B(n41412), .Z(n41299) );
  XOR U50600 ( .A(n41379), .B(n41378), .Z(N61710) );
  XNOR U50601 ( .A(n41396), .B(n41397), .Z(n41378) );
  XNOR U50602 ( .A(n41411), .B(n41412), .Z(n41397) );
  XOR U50603 ( .A(n41408), .B(n41407), .Z(n41412) );
  XOR U50604 ( .A(y[2076]), .B(x[2076]), .Z(n41407) );
  XOR U50605 ( .A(n41410), .B(n41409), .Z(n41408) );
  XOR U50606 ( .A(y[2078]), .B(x[2078]), .Z(n41409) );
  XOR U50607 ( .A(y[2077]), .B(x[2077]), .Z(n41410) );
  XOR U50608 ( .A(n41402), .B(n41401), .Z(n41411) );
  XOR U50609 ( .A(n41404), .B(n41403), .Z(n41401) );
  XOR U50610 ( .A(y[2075]), .B(x[2075]), .Z(n41403) );
  XOR U50611 ( .A(y[2074]), .B(x[2074]), .Z(n41404) );
  XOR U50612 ( .A(y[2073]), .B(x[2073]), .Z(n41402) );
  XNOR U50613 ( .A(n41395), .B(n41394), .Z(n41396) );
  XNOR U50614 ( .A(n41391), .B(n41390), .Z(n41394) );
  XOR U50615 ( .A(n41393), .B(n41392), .Z(n41390) );
  XOR U50616 ( .A(y[2072]), .B(x[2072]), .Z(n41392) );
  XOR U50617 ( .A(y[2071]), .B(x[2071]), .Z(n41393) );
  XOR U50618 ( .A(y[2070]), .B(x[2070]), .Z(n41391) );
  XOR U50619 ( .A(n41385), .B(n41384), .Z(n41395) );
  XOR U50620 ( .A(n41387), .B(n41386), .Z(n41384) );
  XOR U50621 ( .A(y[2069]), .B(x[2069]), .Z(n41386) );
  XOR U50622 ( .A(y[2068]), .B(x[2068]), .Z(n41387) );
  XOR U50623 ( .A(y[2067]), .B(x[2067]), .Z(n41385) );
  XNOR U50624 ( .A(n41361), .B(n41362), .Z(n41379) );
  XNOR U50625 ( .A(n41376), .B(n41377), .Z(n41362) );
  XOR U50626 ( .A(n41373), .B(n41372), .Z(n41377) );
  XOR U50627 ( .A(y[2064]), .B(x[2064]), .Z(n41372) );
  XOR U50628 ( .A(n41375), .B(n41374), .Z(n41373) );
  XOR U50629 ( .A(y[2066]), .B(x[2066]), .Z(n41374) );
  XOR U50630 ( .A(y[2065]), .B(x[2065]), .Z(n41375) );
  XOR U50631 ( .A(n41367), .B(n41366), .Z(n41376) );
  XOR U50632 ( .A(n41369), .B(n41368), .Z(n41366) );
  XOR U50633 ( .A(y[2063]), .B(x[2063]), .Z(n41368) );
  XOR U50634 ( .A(y[2062]), .B(x[2062]), .Z(n41369) );
  XOR U50635 ( .A(y[2061]), .B(x[2061]), .Z(n41367) );
  XNOR U50636 ( .A(n41360), .B(n41359), .Z(n41361) );
  XNOR U50637 ( .A(n41356), .B(n41355), .Z(n41359) );
  XOR U50638 ( .A(n41358), .B(n41357), .Z(n41355) );
  XOR U50639 ( .A(y[2060]), .B(x[2060]), .Z(n41357) );
  XOR U50640 ( .A(y[2059]), .B(x[2059]), .Z(n41358) );
  XOR U50641 ( .A(y[2058]), .B(x[2058]), .Z(n41356) );
  XOR U50642 ( .A(n41350), .B(n41349), .Z(n41360) );
  XOR U50643 ( .A(n41352), .B(n41351), .Z(n41349) );
  XOR U50644 ( .A(y[2057]), .B(x[2057]), .Z(n41351) );
  XOR U50645 ( .A(y[2056]), .B(x[2056]), .Z(n41352) );
  XOR U50646 ( .A(y[2055]), .B(x[2055]), .Z(n41350) );
  NAND U50647 ( .A(n41413), .B(n41414), .Z(N61701) );
  NAND U50648 ( .A(n41415), .B(n41416), .Z(n41414) );
  NANDN U50649 ( .A(n41417), .B(n41418), .Z(n41416) );
  NANDN U50650 ( .A(n41418), .B(n41417), .Z(n41413) );
  XOR U50651 ( .A(n41417), .B(n41419), .Z(N61700) );
  XNOR U50652 ( .A(n41415), .B(n41418), .Z(n41419) );
  NAND U50653 ( .A(n41420), .B(n41421), .Z(n41418) );
  NAND U50654 ( .A(n41422), .B(n41423), .Z(n41421) );
  NANDN U50655 ( .A(n41424), .B(n41425), .Z(n41423) );
  NANDN U50656 ( .A(n41425), .B(n41424), .Z(n41420) );
  AND U50657 ( .A(n41426), .B(n41427), .Z(n41415) );
  NAND U50658 ( .A(n41428), .B(n41429), .Z(n41427) );
  NANDN U50659 ( .A(n41430), .B(n41431), .Z(n41429) );
  NANDN U50660 ( .A(n41431), .B(n41430), .Z(n41426) );
  IV U50661 ( .A(n41432), .Z(n41431) );
  AND U50662 ( .A(n41433), .B(n41434), .Z(n41417) );
  NAND U50663 ( .A(n41435), .B(n41436), .Z(n41434) );
  NANDN U50664 ( .A(n41437), .B(n41438), .Z(n41436) );
  NANDN U50665 ( .A(n41438), .B(n41437), .Z(n41433) );
  XOR U50666 ( .A(n41430), .B(n41439), .Z(N61699) );
  XNOR U50667 ( .A(n41428), .B(n41432), .Z(n41439) );
  XOR U50668 ( .A(n41425), .B(n41440), .Z(n41432) );
  XNOR U50669 ( .A(n41422), .B(n41424), .Z(n41440) );
  AND U50670 ( .A(n41441), .B(n41442), .Z(n41424) );
  NANDN U50671 ( .A(n41443), .B(n41444), .Z(n41442) );
  OR U50672 ( .A(n41445), .B(n41446), .Z(n41444) );
  IV U50673 ( .A(n41447), .Z(n41446) );
  NANDN U50674 ( .A(n41447), .B(n41445), .Z(n41441) );
  AND U50675 ( .A(n41448), .B(n41449), .Z(n41422) );
  NAND U50676 ( .A(n41450), .B(n41451), .Z(n41449) );
  NANDN U50677 ( .A(n41452), .B(n41453), .Z(n41451) );
  NANDN U50678 ( .A(n41453), .B(n41452), .Z(n41448) );
  IV U50679 ( .A(n41454), .Z(n41453) );
  NAND U50680 ( .A(n41455), .B(n41456), .Z(n41425) );
  NANDN U50681 ( .A(n41457), .B(n41458), .Z(n41456) );
  NANDN U50682 ( .A(n41459), .B(n41460), .Z(n41458) );
  NANDN U50683 ( .A(n41460), .B(n41459), .Z(n41455) );
  IV U50684 ( .A(n41461), .Z(n41459) );
  AND U50685 ( .A(n41462), .B(n41463), .Z(n41428) );
  NAND U50686 ( .A(n41464), .B(n41465), .Z(n41463) );
  NANDN U50687 ( .A(n41466), .B(n41467), .Z(n41465) );
  NANDN U50688 ( .A(n41467), .B(n41466), .Z(n41462) );
  XOR U50689 ( .A(n41438), .B(n41468), .Z(n41430) );
  XNOR U50690 ( .A(n41435), .B(n41437), .Z(n41468) );
  AND U50691 ( .A(n41469), .B(n41470), .Z(n41437) );
  NANDN U50692 ( .A(n41471), .B(n41472), .Z(n41470) );
  OR U50693 ( .A(n41473), .B(n41474), .Z(n41472) );
  IV U50694 ( .A(n41475), .Z(n41474) );
  NANDN U50695 ( .A(n41475), .B(n41473), .Z(n41469) );
  AND U50696 ( .A(n41476), .B(n41477), .Z(n41435) );
  NAND U50697 ( .A(n41478), .B(n41479), .Z(n41477) );
  NANDN U50698 ( .A(n41480), .B(n41481), .Z(n41479) );
  NANDN U50699 ( .A(n41481), .B(n41480), .Z(n41476) );
  IV U50700 ( .A(n41482), .Z(n41481) );
  NAND U50701 ( .A(n41483), .B(n41484), .Z(n41438) );
  NANDN U50702 ( .A(n41485), .B(n41486), .Z(n41484) );
  NANDN U50703 ( .A(n41487), .B(n41488), .Z(n41486) );
  NANDN U50704 ( .A(n41488), .B(n41487), .Z(n41483) );
  IV U50705 ( .A(n41489), .Z(n41487) );
  XOR U50706 ( .A(n41464), .B(n41490), .Z(N61698) );
  XNOR U50707 ( .A(n41467), .B(n41466), .Z(n41490) );
  XNOR U50708 ( .A(n41478), .B(n41491), .Z(n41466) );
  XNOR U50709 ( .A(n41482), .B(n41480), .Z(n41491) );
  XOR U50710 ( .A(n41488), .B(n41492), .Z(n41480) );
  XNOR U50711 ( .A(n41485), .B(n41489), .Z(n41492) );
  AND U50712 ( .A(n41493), .B(n41494), .Z(n41489) );
  NAND U50713 ( .A(n41495), .B(n41496), .Z(n41494) );
  NAND U50714 ( .A(n41497), .B(n41498), .Z(n41493) );
  AND U50715 ( .A(n41499), .B(n41500), .Z(n41485) );
  NAND U50716 ( .A(n41501), .B(n41502), .Z(n41500) );
  NAND U50717 ( .A(n41503), .B(n41504), .Z(n41499) );
  NANDN U50718 ( .A(n41505), .B(n41506), .Z(n41488) );
  ANDN U50719 ( .B(n41507), .A(n41508), .Z(n41482) );
  XNOR U50720 ( .A(n41473), .B(n41509), .Z(n41478) );
  XNOR U50721 ( .A(n41471), .B(n41475), .Z(n41509) );
  AND U50722 ( .A(n41510), .B(n41511), .Z(n41475) );
  NAND U50723 ( .A(n41512), .B(n41513), .Z(n41511) );
  NAND U50724 ( .A(n41514), .B(n41515), .Z(n41510) );
  AND U50725 ( .A(n41516), .B(n41517), .Z(n41471) );
  NAND U50726 ( .A(n41518), .B(n41519), .Z(n41517) );
  NAND U50727 ( .A(n41520), .B(n41521), .Z(n41516) );
  AND U50728 ( .A(n41522), .B(n41523), .Z(n41473) );
  NAND U50729 ( .A(n41524), .B(n41525), .Z(n41467) );
  XNOR U50730 ( .A(n41450), .B(n41526), .Z(n41464) );
  XNOR U50731 ( .A(n41454), .B(n41452), .Z(n41526) );
  XOR U50732 ( .A(n41460), .B(n41527), .Z(n41452) );
  XNOR U50733 ( .A(n41457), .B(n41461), .Z(n41527) );
  AND U50734 ( .A(n41528), .B(n41529), .Z(n41461) );
  NAND U50735 ( .A(n41530), .B(n41531), .Z(n41529) );
  NAND U50736 ( .A(n41532), .B(n41533), .Z(n41528) );
  AND U50737 ( .A(n41534), .B(n41535), .Z(n41457) );
  NAND U50738 ( .A(n41536), .B(n41537), .Z(n41535) );
  NAND U50739 ( .A(n41538), .B(n41539), .Z(n41534) );
  NANDN U50740 ( .A(n41540), .B(n41541), .Z(n41460) );
  ANDN U50741 ( .B(n41542), .A(n41543), .Z(n41454) );
  XNOR U50742 ( .A(n41445), .B(n41544), .Z(n41450) );
  XNOR U50743 ( .A(n41443), .B(n41447), .Z(n41544) );
  AND U50744 ( .A(n41545), .B(n41546), .Z(n41447) );
  NAND U50745 ( .A(n41547), .B(n41548), .Z(n41546) );
  NAND U50746 ( .A(n41549), .B(n41550), .Z(n41545) );
  AND U50747 ( .A(n41551), .B(n41552), .Z(n41443) );
  NAND U50748 ( .A(n41553), .B(n41554), .Z(n41552) );
  NAND U50749 ( .A(n41555), .B(n41556), .Z(n41551) );
  AND U50750 ( .A(n41557), .B(n41558), .Z(n41445) );
  XOR U50751 ( .A(n41525), .B(n41524), .Z(N61697) );
  XNOR U50752 ( .A(n41542), .B(n41543), .Z(n41524) );
  XNOR U50753 ( .A(n41557), .B(n41558), .Z(n41543) );
  XOR U50754 ( .A(n41554), .B(n41553), .Z(n41558) );
  XOR U50755 ( .A(y[2052]), .B(x[2052]), .Z(n41553) );
  XOR U50756 ( .A(n41556), .B(n41555), .Z(n41554) );
  XOR U50757 ( .A(y[2054]), .B(x[2054]), .Z(n41555) );
  XOR U50758 ( .A(y[2053]), .B(x[2053]), .Z(n41556) );
  XOR U50759 ( .A(n41548), .B(n41547), .Z(n41557) );
  XOR U50760 ( .A(n41550), .B(n41549), .Z(n41547) );
  XOR U50761 ( .A(y[2051]), .B(x[2051]), .Z(n41549) );
  XOR U50762 ( .A(y[2050]), .B(x[2050]), .Z(n41550) );
  XOR U50763 ( .A(y[2049]), .B(x[2049]), .Z(n41548) );
  XNOR U50764 ( .A(n41541), .B(n41540), .Z(n41542) );
  XNOR U50765 ( .A(n41537), .B(n41536), .Z(n41540) );
  XOR U50766 ( .A(n41539), .B(n41538), .Z(n41536) );
  XOR U50767 ( .A(y[2048]), .B(x[2048]), .Z(n41538) );
  XOR U50768 ( .A(y[2047]), .B(x[2047]), .Z(n41539) );
  XOR U50769 ( .A(y[2046]), .B(x[2046]), .Z(n41537) );
  XOR U50770 ( .A(n41531), .B(n41530), .Z(n41541) );
  XOR U50771 ( .A(n41533), .B(n41532), .Z(n41530) );
  XOR U50772 ( .A(y[2045]), .B(x[2045]), .Z(n41532) );
  XOR U50773 ( .A(y[2044]), .B(x[2044]), .Z(n41533) );
  XOR U50774 ( .A(y[2043]), .B(x[2043]), .Z(n41531) );
  XNOR U50775 ( .A(n41507), .B(n41508), .Z(n41525) );
  XNOR U50776 ( .A(n41522), .B(n41523), .Z(n41508) );
  XOR U50777 ( .A(n41519), .B(n41518), .Z(n41523) );
  XOR U50778 ( .A(y[2040]), .B(x[2040]), .Z(n41518) );
  XOR U50779 ( .A(n41521), .B(n41520), .Z(n41519) );
  XOR U50780 ( .A(y[2042]), .B(x[2042]), .Z(n41520) );
  XOR U50781 ( .A(y[2041]), .B(x[2041]), .Z(n41521) );
  XOR U50782 ( .A(n41513), .B(n41512), .Z(n41522) );
  XOR U50783 ( .A(n41515), .B(n41514), .Z(n41512) );
  XOR U50784 ( .A(y[2039]), .B(x[2039]), .Z(n41514) );
  XOR U50785 ( .A(y[2038]), .B(x[2038]), .Z(n41515) );
  XOR U50786 ( .A(y[2037]), .B(x[2037]), .Z(n41513) );
  XNOR U50787 ( .A(n41506), .B(n41505), .Z(n41507) );
  XNOR U50788 ( .A(n41502), .B(n41501), .Z(n41505) );
  XOR U50789 ( .A(n41504), .B(n41503), .Z(n41501) );
  XOR U50790 ( .A(y[2036]), .B(x[2036]), .Z(n41503) );
  XOR U50791 ( .A(y[2035]), .B(x[2035]), .Z(n41504) );
  XOR U50792 ( .A(y[2034]), .B(x[2034]), .Z(n41502) );
  XOR U50793 ( .A(n41496), .B(n41495), .Z(n41506) );
  XOR U50794 ( .A(n41498), .B(n41497), .Z(n41495) );
  XOR U50795 ( .A(y[2033]), .B(x[2033]), .Z(n41497) );
  XOR U50796 ( .A(y[2032]), .B(x[2032]), .Z(n41498) );
  XOR U50797 ( .A(y[2031]), .B(x[2031]), .Z(n41496) );
  NAND U50798 ( .A(n41559), .B(n41560), .Z(N61688) );
  NAND U50799 ( .A(n41561), .B(n41562), .Z(n41560) );
  NANDN U50800 ( .A(n41563), .B(n41564), .Z(n41562) );
  NANDN U50801 ( .A(n41564), .B(n41563), .Z(n41559) );
  XOR U50802 ( .A(n41563), .B(n41565), .Z(N61687) );
  XNOR U50803 ( .A(n41561), .B(n41564), .Z(n41565) );
  NAND U50804 ( .A(n41566), .B(n41567), .Z(n41564) );
  NAND U50805 ( .A(n41568), .B(n41569), .Z(n41567) );
  NANDN U50806 ( .A(n41570), .B(n41571), .Z(n41569) );
  NANDN U50807 ( .A(n41571), .B(n41570), .Z(n41566) );
  AND U50808 ( .A(n41572), .B(n41573), .Z(n41561) );
  NAND U50809 ( .A(n41574), .B(n41575), .Z(n41573) );
  NANDN U50810 ( .A(n41576), .B(n41577), .Z(n41575) );
  NANDN U50811 ( .A(n41577), .B(n41576), .Z(n41572) );
  IV U50812 ( .A(n41578), .Z(n41577) );
  AND U50813 ( .A(n41579), .B(n41580), .Z(n41563) );
  NAND U50814 ( .A(n41581), .B(n41582), .Z(n41580) );
  NANDN U50815 ( .A(n41583), .B(n41584), .Z(n41582) );
  NANDN U50816 ( .A(n41584), .B(n41583), .Z(n41579) );
  XOR U50817 ( .A(n41576), .B(n41585), .Z(N61686) );
  XNOR U50818 ( .A(n41574), .B(n41578), .Z(n41585) );
  XOR U50819 ( .A(n41571), .B(n41586), .Z(n41578) );
  XNOR U50820 ( .A(n41568), .B(n41570), .Z(n41586) );
  AND U50821 ( .A(n41587), .B(n41588), .Z(n41570) );
  NANDN U50822 ( .A(n41589), .B(n41590), .Z(n41588) );
  OR U50823 ( .A(n41591), .B(n41592), .Z(n41590) );
  IV U50824 ( .A(n41593), .Z(n41592) );
  NANDN U50825 ( .A(n41593), .B(n41591), .Z(n41587) );
  AND U50826 ( .A(n41594), .B(n41595), .Z(n41568) );
  NAND U50827 ( .A(n41596), .B(n41597), .Z(n41595) );
  NANDN U50828 ( .A(n41598), .B(n41599), .Z(n41597) );
  NANDN U50829 ( .A(n41599), .B(n41598), .Z(n41594) );
  IV U50830 ( .A(n41600), .Z(n41599) );
  NAND U50831 ( .A(n41601), .B(n41602), .Z(n41571) );
  NANDN U50832 ( .A(n41603), .B(n41604), .Z(n41602) );
  NANDN U50833 ( .A(n41605), .B(n41606), .Z(n41604) );
  NANDN U50834 ( .A(n41606), .B(n41605), .Z(n41601) );
  IV U50835 ( .A(n41607), .Z(n41605) );
  AND U50836 ( .A(n41608), .B(n41609), .Z(n41574) );
  NAND U50837 ( .A(n41610), .B(n41611), .Z(n41609) );
  NANDN U50838 ( .A(n41612), .B(n41613), .Z(n41611) );
  NANDN U50839 ( .A(n41613), .B(n41612), .Z(n41608) );
  XOR U50840 ( .A(n41584), .B(n41614), .Z(n41576) );
  XNOR U50841 ( .A(n41581), .B(n41583), .Z(n41614) );
  AND U50842 ( .A(n41615), .B(n41616), .Z(n41583) );
  NANDN U50843 ( .A(n41617), .B(n41618), .Z(n41616) );
  OR U50844 ( .A(n41619), .B(n41620), .Z(n41618) );
  IV U50845 ( .A(n41621), .Z(n41620) );
  NANDN U50846 ( .A(n41621), .B(n41619), .Z(n41615) );
  AND U50847 ( .A(n41622), .B(n41623), .Z(n41581) );
  NAND U50848 ( .A(n41624), .B(n41625), .Z(n41623) );
  NANDN U50849 ( .A(n41626), .B(n41627), .Z(n41625) );
  NANDN U50850 ( .A(n41627), .B(n41626), .Z(n41622) );
  IV U50851 ( .A(n41628), .Z(n41627) );
  NAND U50852 ( .A(n41629), .B(n41630), .Z(n41584) );
  NANDN U50853 ( .A(n41631), .B(n41632), .Z(n41630) );
  NANDN U50854 ( .A(n41633), .B(n41634), .Z(n41632) );
  NANDN U50855 ( .A(n41634), .B(n41633), .Z(n41629) );
  IV U50856 ( .A(n41635), .Z(n41633) );
  XOR U50857 ( .A(n41610), .B(n41636), .Z(N61685) );
  XNOR U50858 ( .A(n41613), .B(n41612), .Z(n41636) );
  XNOR U50859 ( .A(n41624), .B(n41637), .Z(n41612) );
  XNOR U50860 ( .A(n41628), .B(n41626), .Z(n41637) );
  XOR U50861 ( .A(n41634), .B(n41638), .Z(n41626) );
  XNOR U50862 ( .A(n41631), .B(n41635), .Z(n41638) );
  AND U50863 ( .A(n41639), .B(n41640), .Z(n41635) );
  NAND U50864 ( .A(n41641), .B(n41642), .Z(n41640) );
  NAND U50865 ( .A(n41643), .B(n41644), .Z(n41639) );
  AND U50866 ( .A(n41645), .B(n41646), .Z(n41631) );
  NAND U50867 ( .A(n41647), .B(n41648), .Z(n41646) );
  NAND U50868 ( .A(n41649), .B(n41650), .Z(n41645) );
  NANDN U50869 ( .A(n41651), .B(n41652), .Z(n41634) );
  ANDN U50870 ( .B(n41653), .A(n41654), .Z(n41628) );
  XNOR U50871 ( .A(n41619), .B(n41655), .Z(n41624) );
  XNOR U50872 ( .A(n41617), .B(n41621), .Z(n41655) );
  AND U50873 ( .A(n41656), .B(n41657), .Z(n41621) );
  NAND U50874 ( .A(n41658), .B(n41659), .Z(n41657) );
  NAND U50875 ( .A(n41660), .B(n41661), .Z(n41656) );
  AND U50876 ( .A(n41662), .B(n41663), .Z(n41617) );
  NAND U50877 ( .A(n41664), .B(n41665), .Z(n41663) );
  NAND U50878 ( .A(n41666), .B(n41667), .Z(n41662) );
  AND U50879 ( .A(n41668), .B(n41669), .Z(n41619) );
  NAND U50880 ( .A(n41670), .B(n41671), .Z(n41613) );
  XNOR U50881 ( .A(n41596), .B(n41672), .Z(n41610) );
  XNOR U50882 ( .A(n41600), .B(n41598), .Z(n41672) );
  XOR U50883 ( .A(n41606), .B(n41673), .Z(n41598) );
  XNOR U50884 ( .A(n41603), .B(n41607), .Z(n41673) );
  AND U50885 ( .A(n41674), .B(n41675), .Z(n41607) );
  NAND U50886 ( .A(n41676), .B(n41677), .Z(n41675) );
  NAND U50887 ( .A(n41678), .B(n41679), .Z(n41674) );
  AND U50888 ( .A(n41680), .B(n41681), .Z(n41603) );
  NAND U50889 ( .A(n41682), .B(n41683), .Z(n41681) );
  NAND U50890 ( .A(n41684), .B(n41685), .Z(n41680) );
  NANDN U50891 ( .A(n41686), .B(n41687), .Z(n41606) );
  ANDN U50892 ( .B(n41688), .A(n41689), .Z(n41600) );
  XNOR U50893 ( .A(n41591), .B(n41690), .Z(n41596) );
  XNOR U50894 ( .A(n41589), .B(n41593), .Z(n41690) );
  AND U50895 ( .A(n41691), .B(n41692), .Z(n41593) );
  NAND U50896 ( .A(n41693), .B(n41694), .Z(n41692) );
  NAND U50897 ( .A(n41695), .B(n41696), .Z(n41691) );
  AND U50898 ( .A(n41697), .B(n41698), .Z(n41589) );
  NAND U50899 ( .A(n41699), .B(n41700), .Z(n41698) );
  NAND U50900 ( .A(n41701), .B(n41702), .Z(n41697) );
  AND U50901 ( .A(n41703), .B(n41704), .Z(n41591) );
  XOR U50902 ( .A(n41671), .B(n41670), .Z(N61684) );
  XNOR U50903 ( .A(n41688), .B(n41689), .Z(n41670) );
  XNOR U50904 ( .A(n41703), .B(n41704), .Z(n41689) );
  XOR U50905 ( .A(n41700), .B(n41699), .Z(n41704) );
  XOR U50906 ( .A(y[2028]), .B(x[2028]), .Z(n41699) );
  XOR U50907 ( .A(n41702), .B(n41701), .Z(n41700) );
  XOR U50908 ( .A(y[2030]), .B(x[2030]), .Z(n41701) );
  XOR U50909 ( .A(y[2029]), .B(x[2029]), .Z(n41702) );
  XOR U50910 ( .A(n41694), .B(n41693), .Z(n41703) );
  XOR U50911 ( .A(n41696), .B(n41695), .Z(n41693) );
  XOR U50912 ( .A(y[2027]), .B(x[2027]), .Z(n41695) );
  XOR U50913 ( .A(y[2026]), .B(x[2026]), .Z(n41696) );
  XOR U50914 ( .A(y[2025]), .B(x[2025]), .Z(n41694) );
  XNOR U50915 ( .A(n41687), .B(n41686), .Z(n41688) );
  XNOR U50916 ( .A(n41683), .B(n41682), .Z(n41686) );
  XOR U50917 ( .A(n41685), .B(n41684), .Z(n41682) );
  XOR U50918 ( .A(y[2024]), .B(x[2024]), .Z(n41684) );
  XOR U50919 ( .A(y[2023]), .B(x[2023]), .Z(n41685) );
  XOR U50920 ( .A(y[2022]), .B(x[2022]), .Z(n41683) );
  XOR U50921 ( .A(n41677), .B(n41676), .Z(n41687) );
  XOR U50922 ( .A(n41679), .B(n41678), .Z(n41676) );
  XOR U50923 ( .A(y[2021]), .B(x[2021]), .Z(n41678) );
  XOR U50924 ( .A(y[2020]), .B(x[2020]), .Z(n41679) );
  XOR U50925 ( .A(y[2019]), .B(x[2019]), .Z(n41677) );
  XNOR U50926 ( .A(n41653), .B(n41654), .Z(n41671) );
  XNOR U50927 ( .A(n41668), .B(n41669), .Z(n41654) );
  XOR U50928 ( .A(n41665), .B(n41664), .Z(n41669) );
  XOR U50929 ( .A(y[2016]), .B(x[2016]), .Z(n41664) );
  XOR U50930 ( .A(n41667), .B(n41666), .Z(n41665) );
  XOR U50931 ( .A(y[2018]), .B(x[2018]), .Z(n41666) );
  XOR U50932 ( .A(y[2017]), .B(x[2017]), .Z(n41667) );
  XOR U50933 ( .A(n41659), .B(n41658), .Z(n41668) );
  XOR U50934 ( .A(n41661), .B(n41660), .Z(n41658) );
  XOR U50935 ( .A(y[2015]), .B(x[2015]), .Z(n41660) );
  XOR U50936 ( .A(y[2014]), .B(x[2014]), .Z(n41661) );
  XOR U50937 ( .A(y[2013]), .B(x[2013]), .Z(n41659) );
  XNOR U50938 ( .A(n41652), .B(n41651), .Z(n41653) );
  XNOR U50939 ( .A(n41648), .B(n41647), .Z(n41651) );
  XOR U50940 ( .A(n41650), .B(n41649), .Z(n41647) );
  XOR U50941 ( .A(y[2012]), .B(x[2012]), .Z(n41649) );
  XOR U50942 ( .A(y[2011]), .B(x[2011]), .Z(n41650) );
  XOR U50943 ( .A(y[2010]), .B(x[2010]), .Z(n41648) );
  XOR U50944 ( .A(n41642), .B(n41641), .Z(n41652) );
  XOR U50945 ( .A(n41644), .B(n41643), .Z(n41641) );
  XOR U50946 ( .A(y[2009]), .B(x[2009]), .Z(n41643) );
  XOR U50947 ( .A(y[2008]), .B(x[2008]), .Z(n41644) );
  XOR U50948 ( .A(y[2007]), .B(x[2007]), .Z(n41642) );
  NAND U50949 ( .A(n41705), .B(n41706), .Z(N61675) );
  NAND U50950 ( .A(n41707), .B(n41708), .Z(n41706) );
  NANDN U50951 ( .A(n41709), .B(n41710), .Z(n41708) );
  NANDN U50952 ( .A(n41710), .B(n41709), .Z(n41705) );
  XOR U50953 ( .A(n41709), .B(n41711), .Z(N61674) );
  XNOR U50954 ( .A(n41707), .B(n41710), .Z(n41711) );
  NAND U50955 ( .A(n41712), .B(n41713), .Z(n41710) );
  NAND U50956 ( .A(n41714), .B(n41715), .Z(n41713) );
  NANDN U50957 ( .A(n41716), .B(n41717), .Z(n41715) );
  NANDN U50958 ( .A(n41717), .B(n41716), .Z(n41712) );
  AND U50959 ( .A(n41718), .B(n41719), .Z(n41707) );
  NAND U50960 ( .A(n41720), .B(n41721), .Z(n41719) );
  NANDN U50961 ( .A(n41722), .B(n41723), .Z(n41721) );
  NANDN U50962 ( .A(n41723), .B(n41722), .Z(n41718) );
  IV U50963 ( .A(n41724), .Z(n41723) );
  AND U50964 ( .A(n41725), .B(n41726), .Z(n41709) );
  NAND U50965 ( .A(n41727), .B(n41728), .Z(n41726) );
  NANDN U50966 ( .A(n41729), .B(n41730), .Z(n41728) );
  NANDN U50967 ( .A(n41730), .B(n41729), .Z(n41725) );
  XOR U50968 ( .A(n41722), .B(n41731), .Z(N61673) );
  XNOR U50969 ( .A(n41720), .B(n41724), .Z(n41731) );
  XOR U50970 ( .A(n41717), .B(n41732), .Z(n41724) );
  XNOR U50971 ( .A(n41714), .B(n41716), .Z(n41732) );
  AND U50972 ( .A(n41733), .B(n41734), .Z(n41716) );
  NANDN U50973 ( .A(n41735), .B(n41736), .Z(n41734) );
  OR U50974 ( .A(n41737), .B(n41738), .Z(n41736) );
  IV U50975 ( .A(n41739), .Z(n41738) );
  NANDN U50976 ( .A(n41739), .B(n41737), .Z(n41733) );
  AND U50977 ( .A(n41740), .B(n41741), .Z(n41714) );
  NAND U50978 ( .A(n41742), .B(n41743), .Z(n41741) );
  NANDN U50979 ( .A(n41744), .B(n41745), .Z(n41743) );
  NANDN U50980 ( .A(n41745), .B(n41744), .Z(n41740) );
  IV U50981 ( .A(n41746), .Z(n41745) );
  NAND U50982 ( .A(n41747), .B(n41748), .Z(n41717) );
  NANDN U50983 ( .A(n41749), .B(n41750), .Z(n41748) );
  NANDN U50984 ( .A(n41751), .B(n41752), .Z(n41750) );
  NANDN U50985 ( .A(n41752), .B(n41751), .Z(n41747) );
  IV U50986 ( .A(n41753), .Z(n41751) );
  AND U50987 ( .A(n41754), .B(n41755), .Z(n41720) );
  NAND U50988 ( .A(n41756), .B(n41757), .Z(n41755) );
  NANDN U50989 ( .A(n41758), .B(n41759), .Z(n41757) );
  NANDN U50990 ( .A(n41759), .B(n41758), .Z(n41754) );
  XOR U50991 ( .A(n41730), .B(n41760), .Z(n41722) );
  XNOR U50992 ( .A(n41727), .B(n41729), .Z(n41760) );
  AND U50993 ( .A(n41761), .B(n41762), .Z(n41729) );
  NANDN U50994 ( .A(n41763), .B(n41764), .Z(n41762) );
  OR U50995 ( .A(n41765), .B(n41766), .Z(n41764) );
  IV U50996 ( .A(n41767), .Z(n41766) );
  NANDN U50997 ( .A(n41767), .B(n41765), .Z(n41761) );
  AND U50998 ( .A(n41768), .B(n41769), .Z(n41727) );
  NAND U50999 ( .A(n41770), .B(n41771), .Z(n41769) );
  NANDN U51000 ( .A(n41772), .B(n41773), .Z(n41771) );
  NANDN U51001 ( .A(n41773), .B(n41772), .Z(n41768) );
  IV U51002 ( .A(n41774), .Z(n41773) );
  NAND U51003 ( .A(n41775), .B(n41776), .Z(n41730) );
  NANDN U51004 ( .A(n41777), .B(n41778), .Z(n41776) );
  NANDN U51005 ( .A(n41779), .B(n41780), .Z(n41778) );
  NANDN U51006 ( .A(n41780), .B(n41779), .Z(n41775) );
  IV U51007 ( .A(n41781), .Z(n41779) );
  XOR U51008 ( .A(n41756), .B(n41782), .Z(N61672) );
  XNOR U51009 ( .A(n41759), .B(n41758), .Z(n41782) );
  XNOR U51010 ( .A(n41770), .B(n41783), .Z(n41758) );
  XNOR U51011 ( .A(n41774), .B(n41772), .Z(n41783) );
  XOR U51012 ( .A(n41780), .B(n41784), .Z(n41772) );
  XNOR U51013 ( .A(n41777), .B(n41781), .Z(n41784) );
  AND U51014 ( .A(n41785), .B(n41786), .Z(n41781) );
  NAND U51015 ( .A(n41787), .B(n41788), .Z(n41786) );
  NAND U51016 ( .A(n41789), .B(n41790), .Z(n41785) );
  AND U51017 ( .A(n41791), .B(n41792), .Z(n41777) );
  NAND U51018 ( .A(n41793), .B(n41794), .Z(n41792) );
  NAND U51019 ( .A(n41795), .B(n41796), .Z(n41791) );
  NANDN U51020 ( .A(n41797), .B(n41798), .Z(n41780) );
  ANDN U51021 ( .B(n41799), .A(n41800), .Z(n41774) );
  XNOR U51022 ( .A(n41765), .B(n41801), .Z(n41770) );
  XNOR U51023 ( .A(n41763), .B(n41767), .Z(n41801) );
  AND U51024 ( .A(n41802), .B(n41803), .Z(n41767) );
  NAND U51025 ( .A(n41804), .B(n41805), .Z(n41803) );
  NAND U51026 ( .A(n41806), .B(n41807), .Z(n41802) );
  AND U51027 ( .A(n41808), .B(n41809), .Z(n41763) );
  NAND U51028 ( .A(n41810), .B(n41811), .Z(n41809) );
  NAND U51029 ( .A(n41812), .B(n41813), .Z(n41808) );
  AND U51030 ( .A(n41814), .B(n41815), .Z(n41765) );
  NAND U51031 ( .A(n41816), .B(n41817), .Z(n41759) );
  XNOR U51032 ( .A(n41742), .B(n41818), .Z(n41756) );
  XNOR U51033 ( .A(n41746), .B(n41744), .Z(n41818) );
  XOR U51034 ( .A(n41752), .B(n41819), .Z(n41744) );
  XNOR U51035 ( .A(n41749), .B(n41753), .Z(n41819) );
  AND U51036 ( .A(n41820), .B(n41821), .Z(n41753) );
  NAND U51037 ( .A(n41822), .B(n41823), .Z(n41821) );
  NAND U51038 ( .A(n41824), .B(n41825), .Z(n41820) );
  AND U51039 ( .A(n41826), .B(n41827), .Z(n41749) );
  NAND U51040 ( .A(n41828), .B(n41829), .Z(n41827) );
  NAND U51041 ( .A(n41830), .B(n41831), .Z(n41826) );
  NANDN U51042 ( .A(n41832), .B(n41833), .Z(n41752) );
  ANDN U51043 ( .B(n41834), .A(n41835), .Z(n41746) );
  XNOR U51044 ( .A(n41737), .B(n41836), .Z(n41742) );
  XNOR U51045 ( .A(n41735), .B(n41739), .Z(n41836) );
  AND U51046 ( .A(n41837), .B(n41838), .Z(n41739) );
  NAND U51047 ( .A(n41839), .B(n41840), .Z(n41838) );
  NAND U51048 ( .A(n41841), .B(n41842), .Z(n41837) );
  AND U51049 ( .A(n41843), .B(n41844), .Z(n41735) );
  NAND U51050 ( .A(n41845), .B(n41846), .Z(n41844) );
  NAND U51051 ( .A(n41847), .B(n41848), .Z(n41843) );
  AND U51052 ( .A(n41849), .B(n41850), .Z(n41737) );
  XOR U51053 ( .A(n41817), .B(n41816), .Z(N61671) );
  XNOR U51054 ( .A(n41834), .B(n41835), .Z(n41816) );
  XNOR U51055 ( .A(n41849), .B(n41850), .Z(n41835) );
  XOR U51056 ( .A(n41846), .B(n41845), .Z(n41850) );
  XOR U51057 ( .A(y[2004]), .B(x[2004]), .Z(n41845) );
  XOR U51058 ( .A(n41848), .B(n41847), .Z(n41846) );
  XOR U51059 ( .A(y[2006]), .B(x[2006]), .Z(n41847) );
  XOR U51060 ( .A(y[2005]), .B(x[2005]), .Z(n41848) );
  XOR U51061 ( .A(n41840), .B(n41839), .Z(n41849) );
  XOR U51062 ( .A(n41842), .B(n41841), .Z(n41839) );
  XOR U51063 ( .A(y[2003]), .B(x[2003]), .Z(n41841) );
  XOR U51064 ( .A(y[2002]), .B(x[2002]), .Z(n41842) );
  XOR U51065 ( .A(y[2001]), .B(x[2001]), .Z(n41840) );
  XNOR U51066 ( .A(n41833), .B(n41832), .Z(n41834) );
  XNOR U51067 ( .A(n41829), .B(n41828), .Z(n41832) );
  XOR U51068 ( .A(n41831), .B(n41830), .Z(n41828) );
  XOR U51069 ( .A(y[2000]), .B(x[2000]), .Z(n41830) );
  XOR U51070 ( .A(y[1999]), .B(x[1999]), .Z(n41831) );
  XOR U51071 ( .A(y[1998]), .B(x[1998]), .Z(n41829) );
  XOR U51072 ( .A(n41823), .B(n41822), .Z(n41833) );
  XOR U51073 ( .A(n41825), .B(n41824), .Z(n41822) );
  XOR U51074 ( .A(y[1997]), .B(x[1997]), .Z(n41824) );
  XOR U51075 ( .A(y[1996]), .B(x[1996]), .Z(n41825) );
  XOR U51076 ( .A(y[1995]), .B(x[1995]), .Z(n41823) );
  XNOR U51077 ( .A(n41799), .B(n41800), .Z(n41817) );
  XNOR U51078 ( .A(n41814), .B(n41815), .Z(n41800) );
  XOR U51079 ( .A(n41811), .B(n41810), .Z(n41815) );
  XOR U51080 ( .A(y[1992]), .B(x[1992]), .Z(n41810) );
  XOR U51081 ( .A(n41813), .B(n41812), .Z(n41811) );
  XOR U51082 ( .A(y[1994]), .B(x[1994]), .Z(n41812) );
  XOR U51083 ( .A(y[1993]), .B(x[1993]), .Z(n41813) );
  XOR U51084 ( .A(n41805), .B(n41804), .Z(n41814) );
  XOR U51085 ( .A(n41807), .B(n41806), .Z(n41804) );
  XOR U51086 ( .A(y[1991]), .B(x[1991]), .Z(n41806) );
  XOR U51087 ( .A(y[1990]), .B(x[1990]), .Z(n41807) );
  XOR U51088 ( .A(y[1989]), .B(x[1989]), .Z(n41805) );
  XNOR U51089 ( .A(n41798), .B(n41797), .Z(n41799) );
  XNOR U51090 ( .A(n41794), .B(n41793), .Z(n41797) );
  XOR U51091 ( .A(n41796), .B(n41795), .Z(n41793) );
  XOR U51092 ( .A(y[1988]), .B(x[1988]), .Z(n41795) );
  XOR U51093 ( .A(y[1987]), .B(x[1987]), .Z(n41796) );
  XOR U51094 ( .A(y[1986]), .B(x[1986]), .Z(n41794) );
  XOR U51095 ( .A(n41788), .B(n41787), .Z(n41798) );
  XOR U51096 ( .A(n41790), .B(n41789), .Z(n41787) );
  XOR U51097 ( .A(y[1985]), .B(x[1985]), .Z(n41789) );
  XOR U51098 ( .A(y[1984]), .B(x[1984]), .Z(n41790) );
  XOR U51099 ( .A(y[1983]), .B(x[1983]), .Z(n41788) );
  NAND U51100 ( .A(n41851), .B(n41852), .Z(N61662) );
  NAND U51101 ( .A(n41853), .B(n41854), .Z(n41852) );
  NANDN U51102 ( .A(n41855), .B(n41856), .Z(n41854) );
  NANDN U51103 ( .A(n41856), .B(n41855), .Z(n41851) );
  XOR U51104 ( .A(n41855), .B(n41857), .Z(N61661) );
  XNOR U51105 ( .A(n41853), .B(n41856), .Z(n41857) );
  NAND U51106 ( .A(n41858), .B(n41859), .Z(n41856) );
  NAND U51107 ( .A(n41860), .B(n41861), .Z(n41859) );
  NANDN U51108 ( .A(n41862), .B(n41863), .Z(n41861) );
  NANDN U51109 ( .A(n41863), .B(n41862), .Z(n41858) );
  AND U51110 ( .A(n41864), .B(n41865), .Z(n41853) );
  NAND U51111 ( .A(n41866), .B(n41867), .Z(n41865) );
  NANDN U51112 ( .A(n41868), .B(n41869), .Z(n41867) );
  NANDN U51113 ( .A(n41869), .B(n41868), .Z(n41864) );
  IV U51114 ( .A(n41870), .Z(n41869) );
  AND U51115 ( .A(n41871), .B(n41872), .Z(n41855) );
  NAND U51116 ( .A(n41873), .B(n41874), .Z(n41872) );
  NANDN U51117 ( .A(n41875), .B(n41876), .Z(n41874) );
  NANDN U51118 ( .A(n41876), .B(n41875), .Z(n41871) );
  XOR U51119 ( .A(n41868), .B(n41877), .Z(N61660) );
  XNOR U51120 ( .A(n41866), .B(n41870), .Z(n41877) );
  XOR U51121 ( .A(n41863), .B(n41878), .Z(n41870) );
  XNOR U51122 ( .A(n41860), .B(n41862), .Z(n41878) );
  AND U51123 ( .A(n41879), .B(n41880), .Z(n41862) );
  NANDN U51124 ( .A(n41881), .B(n41882), .Z(n41880) );
  OR U51125 ( .A(n41883), .B(n41884), .Z(n41882) );
  IV U51126 ( .A(n41885), .Z(n41884) );
  NANDN U51127 ( .A(n41885), .B(n41883), .Z(n41879) );
  AND U51128 ( .A(n41886), .B(n41887), .Z(n41860) );
  NAND U51129 ( .A(n41888), .B(n41889), .Z(n41887) );
  NANDN U51130 ( .A(n41890), .B(n41891), .Z(n41889) );
  NANDN U51131 ( .A(n41891), .B(n41890), .Z(n41886) );
  IV U51132 ( .A(n41892), .Z(n41891) );
  NAND U51133 ( .A(n41893), .B(n41894), .Z(n41863) );
  NANDN U51134 ( .A(n41895), .B(n41896), .Z(n41894) );
  NANDN U51135 ( .A(n41897), .B(n41898), .Z(n41896) );
  NANDN U51136 ( .A(n41898), .B(n41897), .Z(n41893) );
  IV U51137 ( .A(n41899), .Z(n41897) );
  AND U51138 ( .A(n41900), .B(n41901), .Z(n41866) );
  NAND U51139 ( .A(n41902), .B(n41903), .Z(n41901) );
  NANDN U51140 ( .A(n41904), .B(n41905), .Z(n41903) );
  NANDN U51141 ( .A(n41905), .B(n41904), .Z(n41900) );
  XOR U51142 ( .A(n41876), .B(n41906), .Z(n41868) );
  XNOR U51143 ( .A(n41873), .B(n41875), .Z(n41906) );
  AND U51144 ( .A(n41907), .B(n41908), .Z(n41875) );
  NANDN U51145 ( .A(n41909), .B(n41910), .Z(n41908) );
  OR U51146 ( .A(n41911), .B(n41912), .Z(n41910) );
  IV U51147 ( .A(n41913), .Z(n41912) );
  NANDN U51148 ( .A(n41913), .B(n41911), .Z(n41907) );
  AND U51149 ( .A(n41914), .B(n41915), .Z(n41873) );
  NAND U51150 ( .A(n41916), .B(n41917), .Z(n41915) );
  NANDN U51151 ( .A(n41918), .B(n41919), .Z(n41917) );
  NANDN U51152 ( .A(n41919), .B(n41918), .Z(n41914) );
  IV U51153 ( .A(n41920), .Z(n41919) );
  NAND U51154 ( .A(n41921), .B(n41922), .Z(n41876) );
  NANDN U51155 ( .A(n41923), .B(n41924), .Z(n41922) );
  NANDN U51156 ( .A(n41925), .B(n41926), .Z(n41924) );
  NANDN U51157 ( .A(n41926), .B(n41925), .Z(n41921) );
  IV U51158 ( .A(n41927), .Z(n41925) );
  XOR U51159 ( .A(n41902), .B(n41928), .Z(N61659) );
  XNOR U51160 ( .A(n41905), .B(n41904), .Z(n41928) );
  XNOR U51161 ( .A(n41916), .B(n41929), .Z(n41904) );
  XNOR U51162 ( .A(n41920), .B(n41918), .Z(n41929) );
  XOR U51163 ( .A(n41926), .B(n41930), .Z(n41918) );
  XNOR U51164 ( .A(n41923), .B(n41927), .Z(n41930) );
  AND U51165 ( .A(n41931), .B(n41932), .Z(n41927) );
  NAND U51166 ( .A(n41933), .B(n41934), .Z(n41932) );
  NAND U51167 ( .A(n41935), .B(n41936), .Z(n41931) );
  AND U51168 ( .A(n41937), .B(n41938), .Z(n41923) );
  NAND U51169 ( .A(n41939), .B(n41940), .Z(n41938) );
  NAND U51170 ( .A(n41941), .B(n41942), .Z(n41937) );
  NANDN U51171 ( .A(n41943), .B(n41944), .Z(n41926) );
  ANDN U51172 ( .B(n41945), .A(n41946), .Z(n41920) );
  XNOR U51173 ( .A(n41911), .B(n41947), .Z(n41916) );
  XNOR U51174 ( .A(n41909), .B(n41913), .Z(n41947) );
  AND U51175 ( .A(n41948), .B(n41949), .Z(n41913) );
  NAND U51176 ( .A(n41950), .B(n41951), .Z(n41949) );
  NAND U51177 ( .A(n41952), .B(n41953), .Z(n41948) );
  AND U51178 ( .A(n41954), .B(n41955), .Z(n41909) );
  NAND U51179 ( .A(n41956), .B(n41957), .Z(n41955) );
  NAND U51180 ( .A(n41958), .B(n41959), .Z(n41954) );
  AND U51181 ( .A(n41960), .B(n41961), .Z(n41911) );
  NAND U51182 ( .A(n41962), .B(n41963), .Z(n41905) );
  XNOR U51183 ( .A(n41888), .B(n41964), .Z(n41902) );
  XNOR U51184 ( .A(n41892), .B(n41890), .Z(n41964) );
  XOR U51185 ( .A(n41898), .B(n41965), .Z(n41890) );
  XNOR U51186 ( .A(n41895), .B(n41899), .Z(n41965) );
  AND U51187 ( .A(n41966), .B(n41967), .Z(n41899) );
  NAND U51188 ( .A(n41968), .B(n41969), .Z(n41967) );
  NAND U51189 ( .A(n41970), .B(n41971), .Z(n41966) );
  AND U51190 ( .A(n41972), .B(n41973), .Z(n41895) );
  NAND U51191 ( .A(n41974), .B(n41975), .Z(n41973) );
  NAND U51192 ( .A(n41976), .B(n41977), .Z(n41972) );
  NANDN U51193 ( .A(n41978), .B(n41979), .Z(n41898) );
  ANDN U51194 ( .B(n41980), .A(n41981), .Z(n41892) );
  XNOR U51195 ( .A(n41883), .B(n41982), .Z(n41888) );
  XNOR U51196 ( .A(n41881), .B(n41885), .Z(n41982) );
  AND U51197 ( .A(n41983), .B(n41984), .Z(n41885) );
  NAND U51198 ( .A(n41985), .B(n41986), .Z(n41984) );
  NAND U51199 ( .A(n41987), .B(n41988), .Z(n41983) );
  AND U51200 ( .A(n41989), .B(n41990), .Z(n41881) );
  NAND U51201 ( .A(n41991), .B(n41992), .Z(n41990) );
  NAND U51202 ( .A(n41993), .B(n41994), .Z(n41989) );
  AND U51203 ( .A(n41995), .B(n41996), .Z(n41883) );
  XOR U51204 ( .A(n41963), .B(n41962), .Z(N61658) );
  XNOR U51205 ( .A(n41980), .B(n41981), .Z(n41962) );
  XNOR U51206 ( .A(n41995), .B(n41996), .Z(n41981) );
  XOR U51207 ( .A(n41992), .B(n41991), .Z(n41996) );
  XOR U51208 ( .A(y[1980]), .B(x[1980]), .Z(n41991) );
  XOR U51209 ( .A(n41994), .B(n41993), .Z(n41992) );
  XOR U51210 ( .A(y[1982]), .B(x[1982]), .Z(n41993) );
  XOR U51211 ( .A(y[1981]), .B(x[1981]), .Z(n41994) );
  XOR U51212 ( .A(n41986), .B(n41985), .Z(n41995) );
  XOR U51213 ( .A(n41988), .B(n41987), .Z(n41985) );
  XOR U51214 ( .A(y[1979]), .B(x[1979]), .Z(n41987) );
  XOR U51215 ( .A(y[1978]), .B(x[1978]), .Z(n41988) );
  XOR U51216 ( .A(y[1977]), .B(x[1977]), .Z(n41986) );
  XNOR U51217 ( .A(n41979), .B(n41978), .Z(n41980) );
  XNOR U51218 ( .A(n41975), .B(n41974), .Z(n41978) );
  XOR U51219 ( .A(n41977), .B(n41976), .Z(n41974) );
  XOR U51220 ( .A(y[1976]), .B(x[1976]), .Z(n41976) );
  XOR U51221 ( .A(y[1975]), .B(x[1975]), .Z(n41977) );
  XOR U51222 ( .A(y[1974]), .B(x[1974]), .Z(n41975) );
  XOR U51223 ( .A(n41969), .B(n41968), .Z(n41979) );
  XOR U51224 ( .A(n41971), .B(n41970), .Z(n41968) );
  XOR U51225 ( .A(y[1973]), .B(x[1973]), .Z(n41970) );
  XOR U51226 ( .A(y[1972]), .B(x[1972]), .Z(n41971) );
  XOR U51227 ( .A(y[1971]), .B(x[1971]), .Z(n41969) );
  XNOR U51228 ( .A(n41945), .B(n41946), .Z(n41963) );
  XNOR U51229 ( .A(n41960), .B(n41961), .Z(n41946) );
  XOR U51230 ( .A(n41957), .B(n41956), .Z(n41961) );
  XOR U51231 ( .A(y[1968]), .B(x[1968]), .Z(n41956) );
  XOR U51232 ( .A(n41959), .B(n41958), .Z(n41957) );
  XOR U51233 ( .A(y[1970]), .B(x[1970]), .Z(n41958) );
  XOR U51234 ( .A(y[1969]), .B(x[1969]), .Z(n41959) );
  XOR U51235 ( .A(n41951), .B(n41950), .Z(n41960) );
  XOR U51236 ( .A(n41953), .B(n41952), .Z(n41950) );
  XOR U51237 ( .A(y[1967]), .B(x[1967]), .Z(n41952) );
  XOR U51238 ( .A(y[1966]), .B(x[1966]), .Z(n41953) );
  XOR U51239 ( .A(y[1965]), .B(x[1965]), .Z(n41951) );
  XNOR U51240 ( .A(n41944), .B(n41943), .Z(n41945) );
  XNOR U51241 ( .A(n41940), .B(n41939), .Z(n41943) );
  XOR U51242 ( .A(n41942), .B(n41941), .Z(n41939) );
  XOR U51243 ( .A(y[1964]), .B(x[1964]), .Z(n41941) );
  XOR U51244 ( .A(y[1963]), .B(x[1963]), .Z(n41942) );
  XOR U51245 ( .A(y[1962]), .B(x[1962]), .Z(n41940) );
  XOR U51246 ( .A(n41934), .B(n41933), .Z(n41944) );
  XOR U51247 ( .A(n41936), .B(n41935), .Z(n41933) );
  XOR U51248 ( .A(y[1961]), .B(x[1961]), .Z(n41935) );
  XOR U51249 ( .A(y[1960]), .B(x[1960]), .Z(n41936) );
  XOR U51250 ( .A(y[1959]), .B(x[1959]), .Z(n41934) );
  NAND U51251 ( .A(n41997), .B(n41998), .Z(N61649) );
  NAND U51252 ( .A(n41999), .B(n42000), .Z(n41998) );
  NANDN U51253 ( .A(n42001), .B(n42002), .Z(n42000) );
  NANDN U51254 ( .A(n42002), .B(n42001), .Z(n41997) );
  XOR U51255 ( .A(n42001), .B(n42003), .Z(N61648) );
  XNOR U51256 ( .A(n41999), .B(n42002), .Z(n42003) );
  NAND U51257 ( .A(n42004), .B(n42005), .Z(n42002) );
  NAND U51258 ( .A(n42006), .B(n42007), .Z(n42005) );
  NANDN U51259 ( .A(n42008), .B(n42009), .Z(n42007) );
  NANDN U51260 ( .A(n42009), .B(n42008), .Z(n42004) );
  AND U51261 ( .A(n42010), .B(n42011), .Z(n41999) );
  NAND U51262 ( .A(n42012), .B(n42013), .Z(n42011) );
  NANDN U51263 ( .A(n42014), .B(n42015), .Z(n42013) );
  NANDN U51264 ( .A(n42015), .B(n42014), .Z(n42010) );
  IV U51265 ( .A(n42016), .Z(n42015) );
  AND U51266 ( .A(n42017), .B(n42018), .Z(n42001) );
  NAND U51267 ( .A(n42019), .B(n42020), .Z(n42018) );
  NANDN U51268 ( .A(n42021), .B(n42022), .Z(n42020) );
  NANDN U51269 ( .A(n42022), .B(n42021), .Z(n42017) );
  XOR U51270 ( .A(n42014), .B(n42023), .Z(N61647) );
  XNOR U51271 ( .A(n42012), .B(n42016), .Z(n42023) );
  XOR U51272 ( .A(n42009), .B(n42024), .Z(n42016) );
  XNOR U51273 ( .A(n42006), .B(n42008), .Z(n42024) );
  AND U51274 ( .A(n42025), .B(n42026), .Z(n42008) );
  NANDN U51275 ( .A(n42027), .B(n42028), .Z(n42026) );
  OR U51276 ( .A(n42029), .B(n42030), .Z(n42028) );
  IV U51277 ( .A(n42031), .Z(n42030) );
  NANDN U51278 ( .A(n42031), .B(n42029), .Z(n42025) );
  AND U51279 ( .A(n42032), .B(n42033), .Z(n42006) );
  NAND U51280 ( .A(n42034), .B(n42035), .Z(n42033) );
  NANDN U51281 ( .A(n42036), .B(n42037), .Z(n42035) );
  NANDN U51282 ( .A(n42037), .B(n42036), .Z(n42032) );
  IV U51283 ( .A(n42038), .Z(n42037) );
  NAND U51284 ( .A(n42039), .B(n42040), .Z(n42009) );
  NANDN U51285 ( .A(n42041), .B(n42042), .Z(n42040) );
  NANDN U51286 ( .A(n42043), .B(n42044), .Z(n42042) );
  NANDN U51287 ( .A(n42044), .B(n42043), .Z(n42039) );
  IV U51288 ( .A(n42045), .Z(n42043) );
  AND U51289 ( .A(n42046), .B(n42047), .Z(n42012) );
  NAND U51290 ( .A(n42048), .B(n42049), .Z(n42047) );
  NANDN U51291 ( .A(n42050), .B(n42051), .Z(n42049) );
  NANDN U51292 ( .A(n42051), .B(n42050), .Z(n42046) );
  XOR U51293 ( .A(n42022), .B(n42052), .Z(n42014) );
  XNOR U51294 ( .A(n42019), .B(n42021), .Z(n42052) );
  AND U51295 ( .A(n42053), .B(n42054), .Z(n42021) );
  NANDN U51296 ( .A(n42055), .B(n42056), .Z(n42054) );
  OR U51297 ( .A(n42057), .B(n42058), .Z(n42056) );
  IV U51298 ( .A(n42059), .Z(n42058) );
  NANDN U51299 ( .A(n42059), .B(n42057), .Z(n42053) );
  AND U51300 ( .A(n42060), .B(n42061), .Z(n42019) );
  NAND U51301 ( .A(n42062), .B(n42063), .Z(n42061) );
  NANDN U51302 ( .A(n42064), .B(n42065), .Z(n42063) );
  NANDN U51303 ( .A(n42065), .B(n42064), .Z(n42060) );
  IV U51304 ( .A(n42066), .Z(n42065) );
  NAND U51305 ( .A(n42067), .B(n42068), .Z(n42022) );
  NANDN U51306 ( .A(n42069), .B(n42070), .Z(n42068) );
  NANDN U51307 ( .A(n42071), .B(n42072), .Z(n42070) );
  NANDN U51308 ( .A(n42072), .B(n42071), .Z(n42067) );
  IV U51309 ( .A(n42073), .Z(n42071) );
  XOR U51310 ( .A(n42048), .B(n42074), .Z(N61646) );
  XNOR U51311 ( .A(n42051), .B(n42050), .Z(n42074) );
  XNOR U51312 ( .A(n42062), .B(n42075), .Z(n42050) );
  XNOR U51313 ( .A(n42066), .B(n42064), .Z(n42075) );
  XOR U51314 ( .A(n42072), .B(n42076), .Z(n42064) );
  XNOR U51315 ( .A(n42069), .B(n42073), .Z(n42076) );
  AND U51316 ( .A(n42077), .B(n42078), .Z(n42073) );
  NAND U51317 ( .A(n42079), .B(n42080), .Z(n42078) );
  NAND U51318 ( .A(n42081), .B(n42082), .Z(n42077) );
  AND U51319 ( .A(n42083), .B(n42084), .Z(n42069) );
  NAND U51320 ( .A(n42085), .B(n42086), .Z(n42084) );
  NAND U51321 ( .A(n42087), .B(n42088), .Z(n42083) );
  NANDN U51322 ( .A(n42089), .B(n42090), .Z(n42072) );
  ANDN U51323 ( .B(n42091), .A(n42092), .Z(n42066) );
  XNOR U51324 ( .A(n42057), .B(n42093), .Z(n42062) );
  XNOR U51325 ( .A(n42055), .B(n42059), .Z(n42093) );
  AND U51326 ( .A(n42094), .B(n42095), .Z(n42059) );
  NAND U51327 ( .A(n42096), .B(n42097), .Z(n42095) );
  NAND U51328 ( .A(n42098), .B(n42099), .Z(n42094) );
  AND U51329 ( .A(n42100), .B(n42101), .Z(n42055) );
  NAND U51330 ( .A(n42102), .B(n42103), .Z(n42101) );
  NAND U51331 ( .A(n42104), .B(n42105), .Z(n42100) );
  AND U51332 ( .A(n42106), .B(n42107), .Z(n42057) );
  NAND U51333 ( .A(n42108), .B(n42109), .Z(n42051) );
  XNOR U51334 ( .A(n42034), .B(n42110), .Z(n42048) );
  XNOR U51335 ( .A(n42038), .B(n42036), .Z(n42110) );
  XOR U51336 ( .A(n42044), .B(n42111), .Z(n42036) );
  XNOR U51337 ( .A(n42041), .B(n42045), .Z(n42111) );
  AND U51338 ( .A(n42112), .B(n42113), .Z(n42045) );
  NAND U51339 ( .A(n42114), .B(n42115), .Z(n42113) );
  NAND U51340 ( .A(n42116), .B(n42117), .Z(n42112) );
  AND U51341 ( .A(n42118), .B(n42119), .Z(n42041) );
  NAND U51342 ( .A(n42120), .B(n42121), .Z(n42119) );
  NAND U51343 ( .A(n42122), .B(n42123), .Z(n42118) );
  NANDN U51344 ( .A(n42124), .B(n42125), .Z(n42044) );
  ANDN U51345 ( .B(n42126), .A(n42127), .Z(n42038) );
  XNOR U51346 ( .A(n42029), .B(n42128), .Z(n42034) );
  XNOR U51347 ( .A(n42027), .B(n42031), .Z(n42128) );
  AND U51348 ( .A(n42129), .B(n42130), .Z(n42031) );
  NAND U51349 ( .A(n42131), .B(n42132), .Z(n42130) );
  NAND U51350 ( .A(n42133), .B(n42134), .Z(n42129) );
  AND U51351 ( .A(n42135), .B(n42136), .Z(n42027) );
  NAND U51352 ( .A(n42137), .B(n42138), .Z(n42136) );
  NAND U51353 ( .A(n42139), .B(n42140), .Z(n42135) );
  AND U51354 ( .A(n42141), .B(n42142), .Z(n42029) );
  XOR U51355 ( .A(n42109), .B(n42108), .Z(N61645) );
  XNOR U51356 ( .A(n42126), .B(n42127), .Z(n42108) );
  XNOR U51357 ( .A(n42141), .B(n42142), .Z(n42127) );
  XOR U51358 ( .A(n42138), .B(n42137), .Z(n42142) );
  XOR U51359 ( .A(y[1956]), .B(x[1956]), .Z(n42137) );
  XOR U51360 ( .A(n42140), .B(n42139), .Z(n42138) );
  XOR U51361 ( .A(y[1958]), .B(x[1958]), .Z(n42139) );
  XOR U51362 ( .A(y[1957]), .B(x[1957]), .Z(n42140) );
  XOR U51363 ( .A(n42132), .B(n42131), .Z(n42141) );
  XOR U51364 ( .A(n42134), .B(n42133), .Z(n42131) );
  XOR U51365 ( .A(y[1955]), .B(x[1955]), .Z(n42133) );
  XOR U51366 ( .A(y[1954]), .B(x[1954]), .Z(n42134) );
  XOR U51367 ( .A(y[1953]), .B(x[1953]), .Z(n42132) );
  XNOR U51368 ( .A(n42125), .B(n42124), .Z(n42126) );
  XNOR U51369 ( .A(n42121), .B(n42120), .Z(n42124) );
  XOR U51370 ( .A(n42123), .B(n42122), .Z(n42120) );
  XOR U51371 ( .A(y[1952]), .B(x[1952]), .Z(n42122) );
  XOR U51372 ( .A(y[1951]), .B(x[1951]), .Z(n42123) );
  XOR U51373 ( .A(y[1950]), .B(x[1950]), .Z(n42121) );
  XOR U51374 ( .A(n42115), .B(n42114), .Z(n42125) );
  XOR U51375 ( .A(n42117), .B(n42116), .Z(n42114) );
  XOR U51376 ( .A(y[1949]), .B(x[1949]), .Z(n42116) );
  XOR U51377 ( .A(y[1948]), .B(x[1948]), .Z(n42117) );
  XOR U51378 ( .A(y[1947]), .B(x[1947]), .Z(n42115) );
  XNOR U51379 ( .A(n42091), .B(n42092), .Z(n42109) );
  XNOR U51380 ( .A(n42106), .B(n42107), .Z(n42092) );
  XOR U51381 ( .A(n42103), .B(n42102), .Z(n42107) );
  XOR U51382 ( .A(y[1944]), .B(x[1944]), .Z(n42102) );
  XOR U51383 ( .A(n42105), .B(n42104), .Z(n42103) );
  XOR U51384 ( .A(y[1946]), .B(x[1946]), .Z(n42104) );
  XOR U51385 ( .A(y[1945]), .B(x[1945]), .Z(n42105) );
  XOR U51386 ( .A(n42097), .B(n42096), .Z(n42106) );
  XOR U51387 ( .A(n42099), .B(n42098), .Z(n42096) );
  XOR U51388 ( .A(y[1943]), .B(x[1943]), .Z(n42098) );
  XOR U51389 ( .A(y[1942]), .B(x[1942]), .Z(n42099) );
  XOR U51390 ( .A(y[1941]), .B(x[1941]), .Z(n42097) );
  XNOR U51391 ( .A(n42090), .B(n42089), .Z(n42091) );
  XNOR U51392 ( .A(n42086), .B(n42085), .Z(n42089) );
  XOR U51393 ( .A(n42088), .B(n42087), .Z(n42085) );
  XOR U51394 ( .A(y[1940]), .B(x[1940]), .Z(n42087) );
  XOR U51395 ( .A(y[1939]), .B(x[1939]), .Z(n42088) );
  XOR U51396 ( .A(y[1938]), .B(x[1938]), .Z(n42086) );
  XOR U51397 ( .A(n42080), .B(n42079), .Z(n42090) );
  XOR U51398 ( .A(n42082), .B(n42081), .Z(n42079) );
  XOR U51399 ( .A(y[1937]), .B(x[1937]), .Z(n42081) );
  XOR U51400 ( .A(y[1936]), .B(x[1936]), .Z(n42082) );
  XOR U51401 ( .A(y[1935]), .B(x[1935]), .Z(n42080) );
  NAND U51402 ( .A(n42143), .B(n42144), .Z(N61636) );
  NAND U51403 ( .A(n42145), .B(n42146), .Z(n42144) );
  NANDN U51404 ( .A(n42147), .B(n42148), .Z(n42146) );
  NANDN U51405 ( .A(n42148), .B(n42147), .Z(n42143) );
  XOR U51406 ( .A(n42147), .B(n42149), .Z(N61635) );
  XNOR U51407 ( .A(n42145), .B(n42148), .Z(n42149) );
  NAND U51408 ( .A(n42150), .B(n42151), .Z(n42148) );
  NAND U51409 ( .A(n42152), .B(n42153), .Z(n42151) );
  NANDN U51410 ( .A(n42154), .B(n42155), .Z(n42153) );
  NANDN U51411 ( .A(n42155), .B(n42154), .Z(n42150) );
  AND U51412 ( .A(n42156), .B(n42157), .Z(n42145) );
  NAND U51413 ( .A(n42158), .B(n42159), .Z(n42157) );
  NANDN U51414 ( .A(n42160), .B(n42161), .Z(n42159) );
  NANDN U51415 ( .A(n42161), .B(n42160), .Z(n42156) );
  IV U51416 ( .A(n42162), .Z(n42161) );
  AND U51417 ( .A(n42163), .B(n42164), .Z(n42147) );
  NAND U51418 ( .A(n42165), .B(n42166), .Z(n42164) );
  NANDN U51419 ( .A(n42167), .B(n42168), .Z(n42166) );
  NANDN U51420 ( .A(n42168), .B(n42167), .Z(n42163) );
  XOR U51421 ( .A(n42160), .B(n42169), .Z(N61634) );
  XNOR U51422 ( .A(n42158), .B(n42162), .Z(n42169) );
  XOR U51423 ( .A(n42155), .B(n42170), .Z(n42162) );
  XNOR U51424 ( .A(n42152), .B(n42154), .Z(n42170) );
  AND U51425 ( .A(n42171), .B(n42172), .Z(n42154) );
  NANDN U51426 ( .A(n42173), .B(n42174), .Z(n42172) );
  OR U51427 ( .A(n42175), .B(n42176), .Z(n42174) );
  IV U51428 ( .A(n42177), .Z(n42176) );
  NANDN U51429 ( .A(n42177), .B(n42175), .Z(n42171) );
  AND U51430 ( .A(n42178), .B(n42179), .Z(n42152) );
  NAND U51431 ( .A(n42180), .B(n42181), .Z(n42179) );
  NANDN U51432 ( .A(n42182), .B(n42183), .Z(n42181) );
  NANDN U51433 ( .A(n42183), .B(n42182), .Z(n42178) );
  IV U51434 ( .A(n42184), .Z(n42183) );
  NAND U51435 ( .A(n42185), .B(n42186), .Z(n42155) );
  NANDN U51436 ( .A(n42187), .B(n42188), .Z(n42186) );
  NANDN U51437 ( .A(n42189), .B(n42190), .Z(n42188) );
  NANDN U51438 ( .A(n42190), .B(n42189), .Z(n42185) );
  IV U51439 ( .A(n42191), .Z(n42189) );
  AND U51440 ( .A(n42192), .B(n42193), .Z(n42158) );
  NAND U51441 ( .A(n42194), .B(n42195), .Z(n42193) );
  NANDN U51442 ( .A(n42196), .B(n42197), .Z(n42195) );
  NANDN U51443 ( .A(n42197), .B(n42196), .Z(n42192) );
  XOR U51444 ( .A(n42168), .B(n42198), .Z(n42160) );
  XNOR U51445 ( .A(n42165), .B(n42167), .Z(n42198) );
  AND U51446 ( .A(n42199), .B(n42200), .Z(n42167) );
  NANDN U51447 ( .A(n42201), .B(n42202), .Z(n42200) );
  OR U51448 ( .A(n42203), .B(n42204), .Z(n42202) );
  IV U51449 ( .A(n42205), .Z(n42204) );
  NANDN U51450 ( .A(n42205), .B(n42203), .Z(n42199) );
  AND U51451 ( .A(n42206), .B(n42207), .Z(n42165) );
  NAND U51452 ( .A(n42208), .B(n42209), .Z(n42207) );
  NANDN U51453 ( .A(n42210), .B(n42211), .Z(n42209) );
  NANDN U51454 ( .A(n42211), .B(n42210), .Z(n42206) );
  IV U51455 ( .A(n42212), .Z(n42211) );
  NAND U51456 ( .A(n42213), .B(n42214), .Z(n42168) );
  NANDN U51457 ( .A(n42215), .B(n42216), .Z(n42214) );
  NANDN U51458 ( .A(n42217), .B(n42218), .Z(n42216) );
  NANDN U51459 ( .A(n42218), .B(n42217), .Z(n42213) );
  IV U51460 ( .A(n42219), .Z(n42217) );
  XOR U51461 ( .A(n42194), .B(n42220), .Z(N61633) );
  XNOR U51462 ( .A(n42197), .B(n42196), .Z(n42220) );
  XNOR U51463 ( .A(n42208), .B(n42221), .Z(n42196) );
  XNOR U51464 ( .A(n42212), .B(n42210), .Z(n42221) );
  XOR U51465 ( .A(n42218), .B(n42222), .Z(n42210) );
  XNOR U51466 ( .A(n42215), .B(n42219), .Z(n42222) );
  AND U51467 ( .A(n42223), .B(n42224), .Z(n42219) );
  NAND U51468 ( .A(n42225), .B(n42226), .Z(n42224) );
  NAND U51469 ( .A(n42227), .B(n42228), .Z(n42223) );
  AND U51470 ( .A(n42229), .B(n42230), .Z(n42215) );
  NAND U51471 ( .A(n42231), .B(n42232), .Z(n42230) );
  NAND U51472 ( .A(n42233), .B(n42234), .Z(n42229) );
  NANDN U51473 ( .A(n42235), .B(n42236), .Z(n42218) );
  ANDN U51474 ( .B(n42237), .A(n42238), .Z(n42212) );
  XNOR U51475 ( .A(n42203), .B(n42239), .Z(n42208) );
  XNOR U51476 ( .A(n42201), .B(n42205), .Z(n42239) );
  AND U51477 ( .A(n42240), .B(n42241), .Z(n42205) );
  NAND U51478 ( .A(n42242), .B(n42243), .Z(n42241) );
  NAND U51479 ( .A(n42244), .B(n42245), .Z(n42240) );
  AND U51480 ( .A(n42246), .B(n42247), .Z(n42201) );
  NAND U51481 ( .A(n42248), .B(n42249), .Z(n42247) );
  NAND U51482 ( .A(n42250), .B(n42251), .Z(n42246) );
  AND U51483 ( .A(n42252), .B(n42253), .Z(n42203) );
  NAND U51484 ( .A(n42254), .B(n42255), .Z(n42197) );
  XNOR U51485 ( .A(n42180), .B(n42256), .Z(n42194) );
  XNOR U51486 ( .A(n42184), .B(n42182), .Z(n42256) );
  XOR U51487 ( .A(n42190), .B(n42257), .Z(n42182) );
  XNOR U51488 ( .A(n42187), .B(n42191), .Z(n42257) );
  AND U51489 ( .A(n42258), .B(n42259), .Z(n42191) );
  NAND U51490 ( .A(n42260), .B(n42261), .Z(n42259) );
  NAND U51491 ( .A(n42262), .B(n42263), .Z(n42258) );
  AND U51492 ( .A(n42264), .B(n42265), .Z(n42187) );
  NAND U51493 ( .A(n42266), .B(n42267), .Z(n42265) );
  NAND U51494 ( .A(n42268), .B(n42269), .Z(n42264) );
  NANDN U51495 ( .A(n42270), .B(n42271), .Z(n42190) );
  ANDN U51496 ( .B(n42272), .A(n42273), .Z(n42184) );
  XNOR U51497 ( .A(n42175), .B(n42274), .Z(n42180) );
  XNOR U51498 ( .A(n42173), .B(n42177), .Z(n42274) );
  AND U51499 ( .A(n42275), .B(n42276), .Z(n42177) );
  NAND U51500 ( .A(n42277), .B(n42278), .Z(n42276) );
  NAND U51501 ( .A(n42279), .B(n42280), .Z(n42275) );
  AND U51502 ( .A(n42281), .B(n42282), .Z(n42173) );
  NAND U51503 ( .A(n42283), .B(n42284), .Z(n42282) );
  NAND U51504 ( .A(n42285), .B(n42286), .Z(n42281) );
  AND U51505 ( .A(n42287), .B(n42288), .Z(n42175) );
  XOR U51506 ( .A(n42255), .B(n42254), .Z(N61632) );
  XNOR U51507 ( .A(n42272), .B(n42273), .Z(n42254) );
  XNOR U51508 ( .A(n42287), .B(n42288), .Z(n42273) );
  XOR U51509 ( .A(n42284), .B(n42283), .Z(n42288) );
  XOR U51510 ( .A(y[1932]), .B(x[1932]), .Z(n42283) );
  XOR U51511 ( .A(n42286), .B(n42285), .Z(n42284) );
  XOR U51512 ( .A(y[1934]), .B(x[1934]), .Z(n42285) );
  XOR U51513 ( .A(y[1933]), .B(x[1933]), .Z(n42286) );
  XOR U51514 ( .A(n42278), .B(n42277), .Z(n42287) );
  XOR U51515 ( .A(n42280), .B(n42279), .Z(n42277) );
  XOR U51516 ( .A(y[1931]), .B(x[1931]), .Z(n42279) );
  XOR U51517 ( .A(y[1930]), .B(x[1930]), .Z(n42280) );
  XOR U51518 ( .A(y[1929]), .B(x[1929]), .Z(n42278) );
  XNOR U51519 ( .A(n42271), .B(n42270), .Z(n42272) );
  XNOR U51520 ( .A(n42267), .B(n42266), .Z(n42270) );
  XOR U51521 ( .A(n42269), .B(n42268), .Z(n42266) );
  XOR U51522 ( .A(y[1928]), .B(x[1928]), .Z(n42268) );
  XOR U51523 ( .A(y[1927]), .B(x[1927]), .Z(n42269) );
  XOR U51524 ( .A(y[1926]), .B(x[1926]), .Z(n42267) );
  XOR U51525 ( .A(n42261), .B(n42260), .Z(n42271) );
  XOR U51526 ( .A(n42263), .B(n42262), .Z(n42260) );
  XOR U51527 ( .A(y[1925]), .B(x[1925]), .Z(n42262) );
  XOR U51528 ( .A(y[1924]), .B(x[1924]), .Z(n42263) );
  XOR U51529 ( .A(y[1923]), .B(x[1923]), .Z(n42261) );
  XNOR U51530 ( .A(n42237), .B(n42238), .Z(n42255) );
  XNOR U51531 ( .A(n42252), .B(n42253), .Z(n42238) );
  XOR U51532 ( .A(n42249), .B(n42248), .Z(n42253) );
  XOR U51533 ( .A(y[1920]), .B(x[1920]), .Z(n42248) );
  XOR U51534 ( .A(n42251), .B(n42250), .Z(n42249) );
  XOR U51535 ( .A(y[1922]), .B(x[1922]), .Z(n42250) );
  XOR U51536 ( .A(y[1921]), .B(x[1921]), .Z(n42251) );
  XOR U51537 ( .A(n42243), .B(n42242), .Z(n42252) );
  XOR U51538 ( .A(n42245), .B(n42244), .Z(n42242) );
  XOR U51539 ( .A(y[1919]), .B(x[1919]), .Z(n42244) );
  XOR U51540 ( .A(y[1918]), .B(x[1918]), .Z(n42245) );
  XOR U51541 ( .A(y[1917]), .B(x[1917]), .Z(n42243) );
  XNOR U51542 ( .A(n42236), .B(n42235), .Z(n42237) );
  XNOR U51543 ( .A(n42232), .B(n42231), .Z(n42235) );
  XOR U51544 ( .A(n42234), .B(n42233), .Z(n42231) );
  XOR U51545 ( .A(y[1916]), .B(x[1916]), .Z(n42233) );
  XOR U51546 ( .A(y[1915]), .B(x[1915]), .Z(n42234) );
  XOR U51547 ( .A(y[1914]), .B(x[1914]), .Z(n42232) );
  XOR U51548 ( .A(n42226), .B(n42225), .Z(n42236) );
  XOR U51549 ( .A(n42228), .B(n42227), .Z(n42225) );
  XOR U51550 ( .A(y[1913]), .B(x[1913]), .Z(n42227) );
  XOR U51551 ( .A(y[1912]), .B(x[1912]), .Z(n42228) );
  XOR U51552 ( .A(y[1911]), .B(x[1911]), .Z(n42226) );
  NAND U51553 ( .A(n42289), .B(n42290), .Z(N61623) );
  NAND U51554 ( .A(n42291), .B(n42292), .Z(n42290) );
  NANDN U51555 ( .A(n42293), .B(n42294), .Z(n42292) );
  NANDN U51556 ( .A(n42294), .B(n42293), .Z(n42289) );
  XOR U51557 ( .A(n42293), .B(n42295), .Z(N61622) );
  XNOR U51558 ( .A(n42291), .B(n42294), .Z(n42295) );
  NAND U51559 ( .A(n42296), .B(n42297), .Z(n42294) );
  NAND U51560 ( .A(n42298), .B(n42299), .Z(n42297) );
  NANDN U51561 ( .A(n42300), .B(n42301), .Z(n42299) );
  NANDN U51562 ( .A(n42301), .B(n42300), .Z(n42296) );
  AND U51563 ( .A(n42302), .B(n42303), .Z(n42291) );
  NAND U51564 ( .A(n42304), .B(n42305), .Z(n42303) );
  NANDN U51565 ( .A(n42306), .B(n42307), .Z(n42305) );
  NANDN U51566 ( .A(n42307), .B(n42306), .Z(n42302) );
  IV U51567 ( .A(n42308), .Z(n42307) );
  AND U51568 ( .A(n42309), .B(n42310), .Z(n42293) );
  NAND U51569 ( .A(n42311), .B(n42312), .Z(n42310) );
  NANDN U51570 ( .A(n42313), .B(n42314), .Z(n42312) );
  NANDN U51571 ( .A(n42314), .B(n42313), .Z(n42309) );
  XOR U51572 ( .A(n42306), .B(n42315), .Z(N61621) );
  XNOR U51573 ( .A(n42304), .B(n42308), .Z(n42315) );
  XOR U51574 ( .A(n42301), .B(n42316), .Z(n42308) );
  XNOR U51575 ( .A(n42298), .B(n42300), .Z(n42316) );
  AND U51576 ( .A(n42317), .B(n42318), .Z(n42300) );
  NANDN U51577 ( .A(n42319), .B(n42320), .Z(n42318) );
  OR U51578 ( .A(n42321), .B(n42322), .Z(n42320) );
  IV U51579 ( .A(n42323), .Z(n42322) );
  NANDN U51580 ( .A(n42323), .B(n42321), .Z(n42317) );
  AND U51581 ( .A(n42324), .B(n42325), .Z(n42298) );
  NAND U51582 ( .A(n42326), .B(n42327), .Z(n42325) );
  NANDN U51583 ( .A(n42328), .B(n42329), .Z(n42327) );
  NANDN U51584 ( .A(n42329), .B(n42328), .Z(n42324) );
  IV U51585 ( .A(n42330), .Z(n42329) );
  NAND U51586 ( .A(n42331), .B(n42332), .Z(n42301) );
  NANDN U51587 ( .A(n42333), .B(n42334), .Z(n42332) );
  NANDN U51588 ( .A(n42335), .B(n42336), .Z(n42334) );
  NANDN U51589 ( .A(n42336), .B(n42335), .Z(n42331) );
  IV U51590 ( .A(n42337), .Z(n42335) );
  AND U51591 ( .A(n42338), .B(n42339), .Z(n42304) );
  NAND U51592 ( .A(n42340), .B(n42341), .Z(n42339) );
  NANDN U51593 ( .A(n42342), .B(n42343), .Z(n42341) );
  NANDN U51594 ( .A(n42343), .B(n42342), .Z(n42338) );
  XOR U51595 ( .A(n42314), .B(n42344), .Z(n42306) );
  XNOR U51596 ( .A(n42311), .B(n42313), .Z(n42344) );
  AND U51597 ( .A(n42345), .B(n42346), .Z(n42313) );
  NANDN U51598 ( .A(n42347), .B(n42348), .Z(n42346) );
  OR U51599 ( .A(n42349), .B(n42350), .Z(n42348) );
  IV U51600 ( .A(n42351), .Z(n42350) );
  NANDN U51601 ( .A(n42351), .B(n42349), .Z(n42345) );
  AND U51602 ( .A(n42352), .B(n42353), .Z(n42311) );
  NAND U51603 ( .A(n42354), .B(n42355), .Z(n42353) );
  NANDN U51604 ( .A(n42356), .B(n42357), .Z(n42355) );
  NANDN U51605 ( .A(n42357), .B(n42356), .Z(n42352) );
  IV U51606 ( .A(n42358), .Z(n42357) );
  NAND U51607 ( .A(n42359), .B(n42360), .Z(n42314) );
  NANDN U51608 ( .A(n42361), .B(n42362), .Z(n42360) );
  NANDN U51609 ( .A(n42363), .B(n42364), .Z(n42362) );
  NANDN U51610 ( .A(n42364), .B(n42363), .Z(n42359) );
  IV U51611 ( .A(n42365), .Z(n42363) );
  XOR U51612 ( .A(n42340), .B(n42366), .Z(N61620) );
  XNOR U51613 ( .A(n42343), .B(n42342), .Z(n42366) );
  XNOR U51614 ( .A(n42354), .B(n42367), .Z(n42342) );
  XNOR U51615 ( .A(n42358), .B(n42356), .Z(n42367) );
  XOR U51616 ( .A(n42364), .B(n42368), .Z(n42356) );
  XNOR U51617 ( .A(n42361), .B(n42365), .Z(n42368) );
  AND U51618 ( .A(n42369), .B(n42370), .Z(n42365) );
  NAND U51619 ( .A(n42371), .B(n42372), .Z(n42370) );
  NAND U51620 ( .A(n42373), .B(n42374), .Z(n42369) );
  AND U51621 ( .A(n42375), .B(n42376), .Z(n42361) );
  NAND U51622 ( .A(n42377), .B(n42378), .Z(n42376) );
  NAND U51623 ( .A(n42379), .B(n42380), .Z(n42375) );
  NANDN U51624 ( .A(n42381), .B(n42382), .Z(n42364) );
  ANDN U51625 ( .B(n42383), .A(n42384), .Z(n42358) );
  XNOR U51626 ( .A(n42349), .B(n42385), .Z(n42354) );
  XNOR U51627 ( .A(n42347), .B(n42351), .Z(n42385) );
  AND U51628 ( .A(n42386), .B(n42387), .Z(n42351) );
  NAND U51629 ( .A(n42388), .B(n42389), .Z(n42387) );
  NAND U51630 ( .A(n42390), .B(n42391), .Z(n42386) );
  AND U51631 ( .A(n42392), .B(n42393), .Z(n42347) );
  NAND U51632 ( .A(n42394), .B(n42395), .Z(n42393) );
  NAND U51633 ( .A(n42396), .B(n42397), .Z(n42392) );
  AND U51634 ( .A(n42398), .B(n42399), .Z(n42349) );
  NAND U51635 ( .A(n42400), .B(n42401), .Z(n42343) );
  XNOR U51636 ( .A(n42326), .B(n42402), .Z(n42340) );
  XNOR U51637 ( .A(n42330), .B(n42328), .Z(n42402) );
  XOR U51638 ( .A(n42336), .B(n42403), .Z(n42328) );
  XNOR U51639 ( .A(n42333), .B(n42337), .Z(n42403) );
  AND U51640 ( .A(n42404), .B(n42405), .Z(n42337) );
  NAND U51641 ( .A(n42406), .B(n42407), .Z(n42405) );
  NAND U51642 ( .A(n42408), .B(n42409), .Z(n42404) );
  AND U51643 ( .A(n42410), .B(n42411), .Z(n42333) );
  NAND U51644 ( .A(n42412), .B(n42413), .Z(n42411) );
  NAND U51645 ( .A(n42414), .B(n42415), .Z(n42410) );
  NANDN U51646 ( .A(n42416), .B(n42417), .Z(n42336) );
  ANDN U51647 ( .B(n42418), .A(n42419), .Z(n42330) );
  XNOR U51648 ( .A(n42321), .B(n42420), .Z(n42326) );
  XNOR U51649 ( .A(n42319), .B(n42323), .Z(n42420) );
  AND U51650 ( .A(n42421), .B(n42422), .Z(n42323) );
  NAND U51651 ( .A(n42423), .B(n42424), .Z(n42422) );
  NAND U51652 ( .A(n42425), .B(n42426), .Z(n42421) );
  AND U51653 ( .A(n42427), .B(n42428), .Z(n42319) );
  NAND U51654 ( .A(n42429), .B(n42430), .Z(n42428) );
  NAND U51655 ( .A(n42431), .B(n42432), .Z(n42427) );
  AND U51656 ( .A(n42433), .B(n42434), .Z(n42321) );
  XOR U51657 ( .A(n42401), .B(n42400), .Z(N61619) );
  XNOR U51658 ( .A(n42418), .B(n42419), .Z(n42400) );
  XNOR U51659 ( .A(n42433), .B(n42434), .Z(n42419) );
  XOR U51660 ( .A(n42430), .B(n42429), .Z(n42434) );
  XOR U51661 ( .A(y[1908]), .B(x[1908]), .Z(n42429) );
  XOR U51662 ( .A(n42432), .B(n42431), .Z(n42430) );
  XOR U51663 ( .A(y[1910]), .B(x[1910]), .Z(n42431) );
  XOR U51664 ( .A(y[1909]), .B(x[1909]), .Z(n42432) );
  XOR U51665 ( .A(n42424), .B(n42423), .Z(n42433) );
  XOR U51666 ( .A(n42426), .B(n42425), .Z(n42423) );
  XOR U51667 ( .A(y[1907]), .B(x[1907]), .Z(n42425) );
  XOR U51668 ( .A(y[1906]), .B(x[1906]), .Z(n42426) );
  XOR U51669 ( .A(y[1905]), .B(x[1905]), .Z(n42424) );
  XNOR U51670 ( .A(n42417), .B(n42416), .Z(n42418) );
  XNOR U51671 ( .A(n42413), .B(n42412), .Z(n42416) );
  XOR U51672 ( .A(n42415), .B(n42414), .Z(n42412) );
  XOR U51673 ( .A(y[1904]), .B(x[1904]), .Z(n42414) );
  XOR U51674 ( .A(y[1903]), .B(x[1903]), .Z(n42415) );
  XOR U51675 ( .A(y[1902]), .B(x[1902]), .Z(n42413) );
  XOR U51676 ( .A(n42407), .B(n42406), .Z(n42417) );
  XOR U51677 ( .A(n42409), .B(n42408), .Z(n42406) );
  XOR U51678 ( .A(y[1901]), .B(x[1901]), .Z(n42408) );
  XOR U51679 ( .A(y[1900]), .B(x[1900]), .Z(n42409) );
  XOR U51680 ( .A(y[1899]), .B(x[1899]), .Z(n42407) );
  XNOR U51681 ( .A(n42383), .B(n42384), .Z(n42401) );
  XNOR U51682 ( .A(n42398), .B(n42399), .Z(n42384) );
  XOR U51683 ( .A(n42395), .B(n42394), .Z(n42399) );
  XOR U51684 ( .A(y[1896]), .B(x[1896]), .Z(n42394) );
  XOR U51685 ( .A(n42397), .B(n42396), .Z(n42395) );
  XOR U51686 ( .A(y[1898]), .B(x[1898]), .Z(n42396) );
  XOR U51687 ( .A(y[1897]), .B(x[1897]), .Z(n42397) );
  XOR U51688 ( .A(n42389), .B(n42388), .Z(n42398) );
  XOR U51689 ( .A(n42391), .B(n42390), .Z(n42388) );
  XOR U51690 ( .A(y[1895]), .B(x[1895]), .Z(n42390) );
  XOR U51691 ( .A(y[1894]), .B(x[1894]), .Z(n42391) );
  XOR U51692 ( .A(y[1893]), .B(x[1893]), .Z(n42389) );
  XNOR U51693 ( .A(n42382), .B(n42381), .Z(n42383) );
  XNOR U51694 ( .A(n42378), .B(n42377), .Z(n42381) );
  XOR U51695 ( .A(n42380), .B(n42379), .Z(n42377) );
  XOR U51696 ( .A(y[1892]), .B(x[1892]), .Z(n42379) );
  XOR U51697 ( .A(y[1891]), .B(x[1891]), .Z(n42380) );
  XOR U51698 ( .A(y[1890]), .B(x[1890]), .Z(n42378) );
  XOR U51699 ( .A(n42372), .B(n42371), .Z(n42382) );
  XOR U51700 ( .A(n42374), .B(n42373), .Z(n42371) );
  XOR U51701 ( .A(y[1889]), .B(x[1889]), .Z(n42373) );
  XOR U51702 ( .A(y[1888]), .B(x[1888]), .Z(n42374) );
  XOR U51703 ( .A(y[1887]), .B(x[1887]), .Z(n42372) );
  NAND U51704 ( .A(n42435), .B(n42436), .Z(N61610) );
  NAND U51705 ( .A(n42437), .B(n42438), .Z(n42436) );
  NANDN U51706 ( .A(n42439), .B(n42440), .Z(n42438) );
  NANDN U51707 ( .A(n42440), .B(n42439), .Z(n42435) );
  XOR U51708 ( .A(n42439), .B(n42441), .Z(N61609) );
  XNOR U51709 ( .A(n42437), .B(n42440), .Z(n42441) );
  NAND U51710 ( .A(n42442), .B(n42443), .Z(n42440) );
  NAND U51711 ( .A(n42444), .B(n42445), .Z(n42443) );
  NANDN U51712 ( .A(n42446), .B(n42447), .Z(n42445) );
  NANDN U51713 ( .A(n42447), .B(n42446), .Z(n42442) );
  AND U51714 ( .A(n42448), .B(n42449), .Z(n42437) );
  NAND U51715 ( .A(n42450), .B(n42451), .Z(n42449) );
  NANDN U51716 ( .A(n42452), .B(n42453), .Z(n42451) );
  NANDN U51717 ( .A(n42453), .B(n42452), .Z(n42448) );
  IV U51718 ( .A(n42454), .Z(n42453) );
  AND U51719 ( .A(n42455), .B(n42456), .Z(n42439) );
  NAND U51720 ( .A(n42457), .B(n42458), .Z(n42456) );
  NANDN U51721 ( .A(n42459), .B(n42460), .Z(n42458) );
  NANDN U51722 ( .A(n42460), .B(n42459), .Z(n42455) );
  XOR U51723 ( .A(n42452), .B(n42461), .Z(N61608) );
  XNOR U51724 ( .A(n42450), .B(n42454), .Z(n42461) );
  XOR U51725 ( .A(n42447), .B(n42462), .Z(n42454) );
  XNOR U51726 ( .A(n42444), .B(n42446), .Z(n42462) );
  AND U51727 ( .A(n42463), .B(n42464), .Z(n42446) );
  NANDN U51728 ( .A(n42465), .B(n42466), .Z(n42464) );
  OR U51729 ( .A(n42467), .B(n42468), .Z(n42466) );
  IV U51730 ( .A(n42469), .Z(n42468) );
  NANDN U51731 ( .A(n42469), .B(n42467), .Z(n42463) );
  AND U51732 ( .A(n42470), .B(n42471), .Z(n42444) );
  NAND U51733 ( .A(n42472), .B(n42473), .Z(n42471) );
  NANDN U51734 ( .A(n42474), .B(n42475), .Z(n42473) );
  NANDN U51735 ( .A(n42475), .B(n42474), .Z(n42470) );
  IV U51736 ( .A(n42476), .Z(n42475) );
  NAND U51737 ( .A(n42477), .B(n42478), .Z(n42447) );
  NANDN U51738 ( .A(n42479), .B(n42480), .Z(n42478) );
  NANDN U51739 ( .A(n42481), .B(n42482), .Z(n42480) );
  NANDN U51740 ( .A(n42482), .B(n42481), .Z(n42477) );
  IV U51741 ( .A(n42483), .Z(n42481) );
  AND U51742 ( .A(n42484), .B(n42485), .Z(n42450) );
  NAND U51743 ( .A(n42486), .B(n42487), .Z(n42485) );
  NANDN U51744 ( .A(n42488), .B(n42489), .Z(n42487) );
  NANDN U51745 ( .A(n42489), .B(n42488), .Z(n42484) );
  XOR U51746 ( .A(n42460), .B(n42490), .Z(n42452) );
  XNOR U51747 ( .A(n42457), .B(n42459), .Z(n42490) );
  AND U51748 ( .A(n42491), .B(n42492), .Z(n42459) );
  NANDN U51749 ( .A(n42493), .B(n42494), .Z(n42492) );
  OR U51750 ( .A(n42495), .B(n42496), .Z(n42494) );
  IV U51751 ( .A(n42497), .Z(n42496) );
  NANDN U51752 ( .A(n42497), .B(n42495), .Z(n42491) );
  AND U51753 ( .A(n42498), .B(n42499), .Z(n42457) );
  NAND U51754 ( .A(n42500), .B(n42501), .Z(n42499) );
  NANDN U51755 ( .A(n42502), .B(n42503), .Z(n42501) );
  NANDN U51756 ( .A(n42503), .B(n42502), .Z(n42498) );
  IV U51757 ( .A(n42504), .Z(n42503) );
  NAND U51758 ( .A(n42505), .B(n42506), .Z(n42460) );
  NANDN U51759 ( .A(n42507), .B(n42508), .Z(n42506) );
  NANDN U51760 ( .A(n42509), .B(n42510), .Z(n42508) );
  NANDN U51761 ( .A(n42510), .B(n42509), .Z(n42505) );
  IV U51762 ( .A(n42511), .Z(n42509) );
  XOR U51763 ( .A(n42486), .B(n42512), .Z(N61607) );
  XNOR U51764 ( .A(n42489), .B(n42488), .Z(n42512) );
  XNOR U51765 ( .A(n42500), .B(n42513), .Z(n42488) );
  XNOR U51766 ( .A(n42504), .B(n42502), .Z(n42513) );
  XOR U51767 ( .A(n42510), .B(n42514), .Z(n42502) );
  XNOR U51768 ( .A(n42507), .B(n42511), .Z(n42514) );
  AND U51769 ( .A(n42515), .B(n42516), .Z(n42511) );
  NAND U51770 ( .A(n42517), .B(n42518), .Z(n42516) );
  NAND U51771 ( .A(n42519), .B(n42520), .Z(n42515) );
  AND U51772 ( .A(n42521), .B(n42522), .Z(n42507) );
  NAND U51773 ( .A(n42523), .B(n42524), .Z(n42522) );
  NAND U51774 ( .A(n42525), .B(n42526), .Z(n42521) );
  NANDN U51775 ( .A(n42527), .B(n42528), .Z(n42510) );
  ANDN U51776 ( .B(n42529), .A(n42530), .Z(n42504) );
  XNOR U51777 ( .A(n42495), .B(n42531), .Z(n42500) );
  XNOR U51778 ( .A(n42493), .B(n42497), .Z(n42531) );
  AND U51779 ( .A(n42532), .B(n42533), .Z(n42497) );
  NAND U51780 ( .A(n42534), .B(n42535), .Z(n42533) );
  NAND U51781 ( .A(n42536), .B(n42537), .Z(n42532) );
  AND U51782 ( .A(n42538), .B(n42539), .Z(n42493) );
  NAND U51783 ( .A(n42540), .B(n42541), .Z(n42539) );
  NAND U51784 ( .A(n42542), .B(n42543), .Z(n42538) );
  AND U51785 ( .A(n42544), .B(n42545), .Z(n42495) );
  NAND U51786 ( .A(n42546), .B(n42547), .Z(n42489) );
  XNOR U51787 ( .A(n42472), .B(n42548), .Z(n42486) );
  XNOR U51788 ( .A(n42476), .B(n42474), .Z(n42548) );
  XOR U51789 ( .A(n42482), .B(n42549), .Z(n42474) );
  XNOR U51790 ( .A(n42479), .B(n42483), .Z(n42549) );
  AND U51791 ( .A(n42550), .B(n42551), .Z(n42483) );
  NAND U51792 ( .A(n42552), .B(n42553), .Z(n42551) );
  NAND U51793 ( .A(n42554), .B(n42555), .Z(n42550) );
  AND U51794 ( .A(n42556), .B(n42557), .Z(n42479) );
  NAND U51795 ( .A(n42558), .B(n42559), .Z(n42557) );
  NAND U51796 ( .A(n42560), .B(n42561), .Z(n42556) );
  NANDN U51797 ( .A(n42562), .B(n42563), .Z(n42482) );
  ANDN U51798 ( .B(n42564), .A(n42565), .Z(n42476) );
  XNOR U51799 ( .A(n42467), .B(n42566), .Z(n42472) );
  XNOR U51800 ( .A(n42465), .B(n42469), .Z(n42566) );
  AND U51801 ( .A(n42567), .B(n42568), .Z(n42469) );
  NAND U51802 ( .A(n42569), .B(n42570), .Z(n42568) );
  NAND U51803 ( .A(n42571), .B(n42572), .Z(n42567) );
  AND U51804 ( .A(n42573), .B(n42574), .Z(n42465) );
  NAND U51805 ( .A(n42575), .B(n42576), .Z(n42574) );
  NAND U51806 ( .A(n42577), .B(n42578), .Z(n42573) );
  AND U51807 ( .A(n42579), .B(n42580), .Z(n42467) );
  XOR U51808 ( .A(n42547), .B(n42546), .Z(N61606) );
  XNOR U51809 ( .A(n42564), .B(n42565), .Z(n42546) );
  XNOR U51810 ( .A(n42579), .B(n42580), .Z(n42565) );
  XOR U51811 ( .A(n42576), .B(n42575), .Z(n42580) );
  XOR U51812 ( .A(y[1884]), .B(x[1884]), .Z(n42575) );
  XOR U51813 ( .A(n42578), .B(n42577), .Z(n42576) );
  XOR U51814 ( .A(y[1886]), .B(x[1886]), .Z(n42577) );
  XOR U51815 ( .A(y[1885]), .B(x[1885]), .Z(n42578) );
  XOR U51816 ( .A(n42570), .B(n42569), .Z(n42579) );
  XOR U51817 ( .A(n42572), .B(n42571), .Z(n42569) );
  XOR U51818 ( .A(y[1883]), .B(x[1883]), .Z(n42571) );
  XOR U51819 ( .A(y[1882]), .B(x[1882]), .Z(n42572) );
  XOR U51820 ( .A(y[1881]), .B(x[1881]), .Z(n42570) );
  XNOR U51821 ( .A(n42563), .B(n42562), .Z(n42564) );
  XNOR U51822 ( .A(n42559), .B(n42558), .Z(n42562) );
  XOR U51823 ( .A(n42561), .B(n42560), .Z(n42558) );
  XOR U51824 ( .A(y[1880]), .B(x[1880]), .Z(n42560) );
  XOR U51825 ( .A(y[1879]), .B(x[1879]), .Z(n42561) );
  XOR U51826 ( .A(y[1878]), .B(x[1878]), .Z(n42559) );
  XOR U51827 ( .A(n42553), .B(n42552), .Z(n42563) );
  XOR U51828 ( .A(n42555), .B(n42554), .Z(n42552) );
  XOR U51829 ( .A(y[1877]), .B(x[1877]), .Z(n42554) );
  XOR U51830 ( .A(y[1876]), .B(x[1876]), .Z(n42555) );
  XOR U51831 ( .A(y[1875]), .B(x[1875]), .Z(n42553) );
  XNOR U51832 ( .A(n42529), .B(n42530), .Z(n42547) );
  XNOR U51833 ( .A(n42544), .B(n42545), .Z(n42530) );
  XOR U51834 ( .A(n42541), .B(n42540), .Z(n42545) );
  XOR U51835 ( .A(y[1872]), .B(x[1872]), .Z(n42540) );
  XOR U51836 ( .A(n42543), .B(n42542), .Z(n42541) );
  XOR U51837 ( .A(y[1874]), .B(x[1874]), .Z(n42542) );
  XOR U51838 ( .A(y[1873]), .B(x[1873]), .Z(n42543) );
  XOR U51839 ( .A(n42535), .B(n42534), .Z(n42544) );
  XOR U51840 ( .A(n42537), .B(n42536), .Z(n42534) );
  XOR U51841 ( .A(y[1871]), .B(x[1871]), .Z(n42536) );
  XOR U51842 ( .A(y[1870]), .B(x[1870]), .Z(n42537) );
  XOR U51843 ( .A(y[1869]), .B(x[1869]), .Z(n42535) );
  XNOR U51844 ( .A(n42528), .B(n42527), .Z(n42529) );
  XNOR U51845 ( .A(n42524), .B(n42523), .Z(n42527) );
  XOR U51846 ( .A(n42526), .B(n42525), .Z(n42523) );
  XOR U51847 ( .A(y[1868]), .B(x[1868]), .Z(n42525) );
  XOR U51848 ( .A(y[1867]), .B(x[1867]), .Z(n42526) );
  XOR U51849 ( .A(y[1866]), .B(x[1866]), .Z(n42524) );
  XOR U51850 ( .A(n42518), .B(n42517), .Z(n42528) );
  XOR U51851 ( .A(n42520), .B(n42519), .Z(n42517) );
  XOR U51852 ( .A(y[1865]), .B(x[1865]), .Z(n42519) );
  XOR U51853 ( .A(y[1864]), .B(x[1864]), .Z(n42520) );
  XOR U51854 ( .A(y[1863]), .B(x[1863]), .Z(n42518) );
  NAND U51855 ( .A(n42581), .B(n42582), .Z(N61597) );
  NAND U51856 ( .A(n42583), .B(n42584), .Z(n42582) );
  NANDN U51857 ( .A(n42585), .B(n42586), .Z(n42584) );
  NANDN U51858 ( .A(n42586), .B(n42585), .Z(n42581) );
  XOR U51859 ( .A(n42585), .B(n42587), .Z(N61596) );
  XNOR U51860 ( .A(n42583), .B(n42586), .Z(n42587) );
  NAND U51861 ( .A(n42588), .B(n42589), .Z(n42586) );
  NAND U51862 ( .A(n42590), .B(n42591), .Z(n42589) );
  NANDN U51863 ( .A(n42592), .B(n42593), .Z(n42591) );
  NANDN U51864 ( .A(n42593), .B(n42592), .Z(n42588) );
  AND U51865 ( .A(n42594), .B(n42595), .Z(n42583) );
  NAND U51866 ( .A(n42596), .B(n42597), .Z(n42595) );
  NANDN U51867 ( .A(n42598), .B(n42599), .Z(n42597) );
  NANDN U51868 ( .A(n42599), .B(n42598), .Z(n42594) );
  IV U51869 ( .A(n42600), .Z(n42599) );
  AND U51870 ( .A(n42601), .B(n42602), .Z(n42585) );
  NAND U51871 ( .A(n42603), .B(n42604), .Z(n42602) );
  NANDN U51872 ( .A(n42605), .B(n42606), .Z(n42604) );
  NANDN U51873 ( .A(n42606), .B(n42605), .Z(n42601) );
  XOR U51874 ( .A(n42598), .B(n42607), .Z(N61595) );
  XNOR U51875 ( .A(n42596), .B(n42600), .Z(n42607) );
  XOR U51876 ( .A(n42593), .B(n42608), .Z(n42600) );
  XNOR U51877 ( .A(n42590), .B(n42592), .Z(n42608) );
  AND U51878 ( .A(n42609), .B(n42610), .Z(n42592) );
  NANDN U51879 ( .A(n42611), .B(n42612), .Z(n42610) );
  OR U51880 ( .A(n42613), .B(n42614), .Z(n42612) );
  IV U51881 ( .A(n42615), .Z(n42614) );
  NANDN U51882 ( .A(n42615), .B(n42613), .Z(n42609) );
  AND U51883 ( .A(n42616), .B(n42617), .Z(n42590) );
  NAND U51884 ( .A(n42618), .B(n42619), .Z(n42617) );
  NANDN U51885 ( .A(n42620), .B(n42621), .Z(n42619) );
  NANDN U51886 ( .A(n42621), .B(n42620), .Z(n42616) );
  IV U51887 ( .A(n42622), .Z(n42621) );
  NAND U51888 ( .A(n42623), .B(n42624), .Z(n42593) );
  NANDN U51889 ( .A(n42625), .B(n42626), .Z(n42624) );
  NANDN U51890 ( .A(n42627), .B(n42628), .Z(n42626) );
  NANDN U51891 ( .A(n42628), .B(n42627), .Z(n42623) );
  IV U51892 ( .A(n42629), .Z(n42627) );
  AND U51893 ( .A(n42630), .B(n42631), .Z(n42596) );
  NAND U51894 ( .A(n42632), .B(n42633), .Z(n42631) );
  NANDN U51895 ( .A(n42634), .B(n42635), .Z(n42633) );
  NANDN U51896 ( .A(n42635), .B(n42634), .Z(n42630) );
  XOR U51897 ( .A(n42606), .B(n42636), .Z(n42598) );
  XNOR U51898 ( .A(n42603), .B(n42605), .Z(n42636) );
  AND U51899 ( .A(n42637), .B(n42638), .Z(n42605) );
  NANDN U51900 ( .A(n42639), .B(n42640), .Z(n42638) );
  OR U51901 ( .A(n42641), .B(n42642), .Z(n42640) );
  IV U51902 ( .A(n42643), .Z(n42642) );
  NANDN U51903 ( .A(n42643), .B(n42641), .Z(n42637) );
  AND U51904 ( .A(n42644), .B(n42645), .Z(n42603) );
  NAND U51905 ( .A(n42646), .B(n42647), .Z(n42645) );
  NANDN U51906 ( .A(n42648), .B(n42649), .Z(n42647) );
  NANDN U51907 ( .A(n42649), .B(n42648), .Z(n42644) );
  IV U51908 ( .A(n42650), .Z(n42649) );
  NAND U51909 ( .A(n42651), .B(n42652), .Z(n42606) );
  NANDN U51910 ( .A(n42653), .B(n42654), .Z(n42652) );
  NANDN U51911 ( .A(n42655), .B(n42656), .Z(n42654) );
  NANDN U51912 ( .A(n42656), .B(n42655), .Z(n42651) );
  IV U51913 ( .A(n42657), .Z(n42655) );
  XOR U51914 ( .A(n42632), .B(n42658), .Z(N61594) );
  XNOR U51915 ( .A(n42635), .B(n42634), .Z(n42658) );
  XNOR U51916 ( .A(n42646), .B(n42659), .Z(n42634) );
  XNOR U51917 ( .A(n42650), .B(n42648), .Z(n42659) );
  XOR U51918 ( .A(n42656), .B(n42660), .Z(n42648) );
  XNOR U51919 ( .A(n42653), .B(n42657), .Z(n42660) );
  AND U51920 ( .A(n42661), .B(n42662), .Z(n42657) );
  NAND U51921 ( .A(n42663), .B(n42664), .Z(n42662) );
  NAND U51922 ( .A(n42665), .B(n42666), .Z(n42661) );
  AND U51923 ( .A(n42667), .B(n42668), .Z(n42653) );
  NAND U51924 ( .A(n42669), .B(n42670), .Z(n42668) );
  NAND U51925 ( .A(n42671), .B(n42672), .Z(n42667) );
  NANDN U51926 ( .A(n42673), .B(n42674), .Z(n42656) );
  ANDN U51927 ( .B(n42675), .A(n42676), .Z(n42650) );
  XNOR U51928 ( .A(n42641), .B(n42677), .Z(n42646) );
  XNOR U51929 ( .A(n42639), .B(n42643), .Z(n42677) );
  AND U51930 ( .A(n42678), .B(n42679), .Z(n42643) );
  NAND U51931 ( .A(n42680), .B(n42681), .Z(n42679) );
  NAND U51932 ( .A(n42682), .B(n42683), .Z(n42678) );
  AND U51933 ( .A(n42684), .B(n42685), .Z(n42639) );
  NAND U51934 ( .A(n42686), .B(n42687), .Z(n42685) );
  NAND U51935 ( .A(n42688), .B(n42689), .Z(n42684) );
  AND U51936 ( .A(n42690), .B(n42691), .Z(n42641) );
  NAND U51937 ( .A(n42692), .B(n42693), .Z(n42635) );
  XNOR U51938 ( .A(n42618), .B(n42694), .Z(n42632) );
  XNOR U51939 ( .A(n42622), .B(n42620), .Z(n42694) );
  XOR U51940 ( .A(n42628), .B(n42695), .Z(n42620) );
  XNOR U51941 ( .A(n42625), .B(n42629), .Z(n42695) );
  AND U51942 ( .A(n42696), .B(n42697), .Z(n42629) );
  NAND U51943 ( .A(n42698), .B(n42699), .Z(n42697) );
  NAND U51944 ( .A(n42700), .B(n42701), .Z(n42696) );
  AND U51945 ( .A(n42702), .B(n42703), .Z(n42625) );
  NAND U51946 ( .A(n42704), .B(n42705), .Z(n42703) );
  NAND U51947 ( .A(n42706), .B(n42707), .Z(n42702) );
  NANDN U51948 ( .A(n42708), .B(n42709), .Z(n42628) );
  ANDN U51949 ( .B(n42710), .A(n42711), .Z(n42622) );
  XNOR U51950 ( .A(n42613), .B(n42712), .Z(n42618) );
  XNOR U51951 ( .A(n42611), .B(n42615), .Z(n42712) );
  AND U51952 ( .A(n42713), .B(n42714), .Z(n42615) );
  NAND U51953 ( .A(n42715), .B(n42716), .Z(n42714) );
  NAND U51954 ( .A(n42717), .B(n42718), .Z(n42713) );
  AND U51955 ( .A(n42719), .B(n42720), .Z(n42611) );
  NAND U51956 ( .A(n42721), .B(n42722), .Z(n42720) );
  NAND U51957 ( .A(n42723), .B(n42724), .Z(n42719) );
  AND U51958 ( .A(n42725), .B(n42726), .Z(n42613) );
  XOR U51959 ( .A(n42693), .B(n42692), .Z(N61593) );
  XNOR U51960 ( .A(n42710), .B(n42711), .Z(n42692) );
  XNOR U51961 ( .A(n42725), .B(n42726), .Z(n42711) );
  XOR U51962 ( .A(n42722), .B(n42721), .Z(n42726) );
  XOR U51963 ( .A(y[1860]), .B(x[1860]), .Z(n42721) );
  XOR U51964 ( .A(n42724), .B(n42723), .Z(n42722) );
  XOR U51965 ( .A(y[1862]), .B(x[1862]), .Z(n42723) );
  XOR U51966 ( .A(y[1861]), .B(x[1861]), .Z(n42724) );
  XOR U51967 ( .A(n42716), .B(n42715), .Z(n42725) );
  XOR U51968 ( .A(n42718), .B(n42717), .Z(n42715) );
  XOR U51969 ( .A(y[1859]), .B(x[1859]), .Z(n42717) );
  XOR U51970 ( .A(y[1858]), .B(x[1858]), .Z(n42718) );
  XOR U51971 ( .A(y[1857]), .B(x[1857]), .Z(n42716) );
  XNOR U51972 ( .A(n42709), .B(n42708), .Z(n42710) );
  XNOR U51973 ( .A(n42705), .B(n42704), .Z(n42708) );
  XOR U51974 ( .A(n42707), .B(n42706), .Z(n42704) );
  XOR U51975 ( .A(y[1856]), .B(x[1856]), .Z(n42706) );
  XOR U51976 ( .A(y[1855]), .B(x[1855]), .Z(n42707) );
  XOR U51977 ( .A(y[1854]), .B(x[1854]), .Z(n42705) );
  XOR U51978 ( .A(n42699), .B(n42698), .Z(n42709) );
  XOR U51979 ( .A(n42701), .B(n42700), .Z(n42698) );
  XOR U51980 ( .A(y[1853]), .B(x[1853]), .Z(n42700) );
  XOR U51981 ( .A(y[1852]), .B(x[1852]), .Z(n42701) );
  XOR U51982 ( .A(y[1851]), .B(x[1851]), .Z(n42699) );
  XNOR U51983 ( .A(n42675), .B(n42676), .Z(n42693) );
  XNOR U51984 ( .A(n42690), .B(n42691), .Z(n42676) );
  XOR U51985 ( .A(n42687), .B(n42686), .Z(n42691) );
  XOR U51986 ( .A(y[1848]), .B(x[1848]), .Z(n42686) );
  XOR U51987 ( .A(n42689), .B(n42688), .Z(n42687) );
  XOR U51988 ( .A(y[1850]), .B(x[1850]), .Z(n42688) );
  XOR U51989 ( .A(y[1849]), .B(x[1849]), .Z(n42689) );
  XOR U51990 ( .A(n42681), .B(n42680), .Z(n42690) );
  XOR U51991 ( .A(n42683), .B(n42682), .Z(n42680) );
  XOR U51992 ( .A(y[1847]), .B(x[1847]), .Z(n42682) );
  XOR U51993 ( .A(y[1846]), .B(x[1846]), .Z(n42683) );
  XOR U51994 ( .A(y[1845]), .B(x[1845]), .Z(n42681) );
  XNOR U51995 ( .A(n42674), .B(n42673), .Z(n42675) );
  XNOR U51996 ( .A(n42670), .B(n42669), .Z(n42673) );
  XOR U51997 ( .A(n42672), .B(n42671), .Z(n42669) );
  XOR U51998 ( .A(y[1844]), .B(x[1844]), .Z(n42671) );
  XOR U51999 ( .A(y[1843]), .B(x[1843]), .Z(n42672) );
  XOR U52000 ( .A(y[1842]), .B(x[1842]), .Z(n42670) );
  XOR U52001 ( .A(n42664), .B(n42663), .Z(n42674) );
  XOR U52002 ( .A(n42666), .B(n42665), .Z(n42663) );
  XOR U52003 ( .A(y[1841]), .B(x[1841]), .Z(n42665) );
  XOR U52004 ( .A(y[1840]), .B(x[1840]), .Z(n42666) );
  XOR U52005 ( .A(y[1839]), .B(x[1839]), .Z(n42664) );
  NAND U52006 ( .A(n42727), .B(n42728), .Z(N61584) );
  NAND U52007 ( .A(n42729), .B(n42730), .Z(n42728) );
  NANDN U52008 ( .A(n42731), .B(n42732), .Z(n42730) );
  NANDN U52009 ( .A(n42732), .B(n42731), .Z(n42727) );
  XOR U52010 ( .A(n42731), .B(n42733), .Z(N61583) );
  XNOR U52011 ( .A(n42729), .B(n42732), .Z(n42733) );
  NAND U52012 ( .A(n42734), .B(n42735), .Z(n42732) );
  NAND U52013 ( .A(n42736), .B(n42737), .Z(n42735) );
  NANDN U52014 ( .A(n42738), .B(n42739), .Z(n42737) );
  NANDN U52015 ( .A(n42739), .B(n42738), .Z(n42734) );
  AND U52016 ( .A(n42740), .B(n42741), .Z(n42729) );
  NAND U52017 ( .A(n42742), .B(n42743), .Z(n42741) );
  NANDN U52018 ( .A(n42744), .B(n42745), .Z(n42743) );
  NANDN U52019 ( .A(n42745), .B(n42744), .Z(n42740) );
  IV U52020 ( .A(n42746), .Z(n42745) );
  AND U52021 ( .A(n42747), .B(n42748), .Z(n42731) );
  NAND U52022 ( .A(n42749), .B(n42750), .Z(n42748) );
  NANDN U52023 ( .A(n42751), .B(n42752), .Z(n42750) );
  NANDN U52024 ( .A(n42752), .B(n42751), .Z(n42747) );
  XOR U52025 ( .A(n42744), .B(n42753), .Z(N61582) );
  XNOR U52026 ( .A(n42742), .B(n42746), .Z(n42753) );
  XOR U52027 ( .A(n42739), .B(n42754), .Z(n42746) );
  XNOR U52028 ( .A(n42736), .B(n42738), .Z(n42754) );
  AND U52029 ( .A(n42755), .B(n42756), .Z(n42738) );
  NANDN U52030 ( .A(n42757), .B(n42758), .Z(n42756) );
  OR U52031 ( .A(n42759), .B(n42760), .Z(n42758) );
  IV U52032 ( .A(n42761), .Z(n42760) );
  NANDN U52033 ( .A(n42761), .B(n42759), .Z(n42755) );
  AND U52034 ( .A(n42762), .B(n42763), .Z(n42736) );
  NAND U52035 ( .A(n42764), .B(n42765), .Z(n42763) );
  NANDN U52036 ( .A(n42766), .B(n42767), .Z(n42765) );
  NANDN U52037 ( .A(n42767), .B(n42766), .Z(n42762) );
  IV U52038 ( .A(n42768), .Z(n42767) );
  NAND U52039 ( .A(n42769), .B(n42770), .Z(n42739) );
  NANDN U52040 ( .A(n42771), .B(n42772), .Z(n42770) );
  NANDN U52041 ( .A(n42773), .B(n42774), .Z(n42772) );
  NANDN U52042 ( .A(n42774), .B(n42773), .Z(n42769) );
  IV U52043 ( .A(n42775), .Z(n42773) );
  AND U52044 ( .A(n42776), .B(n42777), .Z(n42742) );
  NAND U52045 ( .A(n42778), .B(n42779), .Z(n42777) );
  NANDN U52046 ( .A(n42780), .B(n42781), .Z(n42779) );
  NANDN U52047 ( .A(n42781), .B(n42780), .Z(n42776) );
  XOR U52048 ( .A(n42752), .B(n42782), .Z(n42744) );
  XNOR U52049 ( .A(n42749), .B(n42751), .Z(n42782) );
  AND U52050 ( .A(n42783), .B(n42784), .Z(n42751) );
  NANDN U52051 ( .A(n42785), .B(n42786), .Z(n42784) );
  OR U52052 ( .A(n42787), .B(n42788), .Z(n42786) );
  IV U52053 ( .A(n42789), .Z(n42788) );
  NANDN U52054 ( .A(n42789), .B(n42787), .Z(n42783) );
  AND U52055 ( .A(n42790), .B(n42791), .Z(n42749) );
  NAND U52056 ( .A(n42792), .B(n42793), .Z(n42791) );
  NANDN U52057 ( .A(n42794), .B(n42795), .Z(n42793) );
  NANDN U52058 ( .A(n42795), .B(n42794), .Z(n42790) );
  IV U52059 ( .A(n42796), .Z(n42795) );
  NAND U52060 ( .A(n42797), .B(n42798), .Z(n42752) );
  NANDN U52061 ( .A(n42799), .B(n42800), .Z(n42798) );
  NANDN U52062 ( .A(n42801), .B(n42802), .Z(n42800) );
  NANDN U52063 ( .A(n42802), .B(n42801), .Z(n42797) );
  IV U52064 ( .A(n42803), .Z(n42801) );
  XOR U52065 ( .A(n42778), .B(n42804), .Z(N61581) );
  XNOR U52066 ( .A(n42781), .B(n42780), .Z(n42804) );
  XNOR U52067 ( .A(n42792), .B(n42805), .Z(n42780) );
  XNOR U52068 ( .A(n42796), .B(n42794), .Z(n42805) );
  XOR U52069 ( .A(n42802), .B(n42806), .Z(n42794) );
  XNOR U52070 ( .A(n42799), .B(n42803), .Z(n42806) );
  AND U52071 ( .A(n42807), .B(n42808), .Z(n42803) );
  NAND U52072 ( .A(n42809), .B(n42810), .Z(n42808) );
  NAND U52073 ( .A(n42811), .B(n42812), .Z(n42807) );
  AND U52074 ( .A(n42813), .B(n42814), .Z(n42799) );
  NAND U52075 ( .A(n42815), .B(n42816), .Z(n42814) );
  NAND U52076 ( .A(n42817), .B(n42818), .Z(n42813) );
  NANDN U52077 ( .A(n42819), .B(n42820), .Z(n42802) );
  ANDN U52078 ( .B(n42821), .A(n42822), .Z(n42796) );
  XNOR U52079 ( .A(n42787), .B(n42823), .Z(n42792) );
  XNOR U52080 ( .A(n42785), .B(n42789), .Z(n42823) );
  AND U52081 ( .A(n42824), .B(n42825), .Z(n42789) );
  NAND U52082 ( .A(n42826), .B(n42827), .Z(n42825) );
  NAND U52083 ( .A(n42828), .B(n42829), .Z(n42824) );
  AND U52084 ( .A(n42830), .B(n42831), .Z(n42785) );
  NAND U52085 ( .A(n42832), .B(n42833), .Z(n42831) );
  NAND U52086 ( .A(n42834), .B(n42835), .Z(n42830) );
  AND U52087 ( .A(n42836), .B(n42837), .Z(n42787) );
  NAND U52088 ( .A(n42838), .B(n42839), .Z(n42781) );
  XNOR U52089 ( .A(n42764), .B(n42840), .Z(n42778) );
  XNOR U52090 ( .A(n42768), .B(n42766), .Z(n42840) );
  XOR U52091 ( .A(n42774), .B(n42841), .Z(n42766) );
  XNOR U52092 ( .A(n42771), .B(n42775), .Z(n42841) );
  AND U52093 ( .A(n42842), .B(n42843), .Z(n42775) );
  NAND U52094 ( .A(n42844), .B(n42845), .Z(n42843) );
  NAND U52095 ( .A(n42846), .B(n42847), .Z(n42842) );
  AND U52096 ( .A(n42848), .B(n42849), .Z(n42771) );
  NAND U52097 ( .A(n42850), .B(n42851), .Z(n42849) );
  NAND U52098 ( .A(n42852), .B(n42853), .Z(n42848) );
  NANDN U52099 ( .A(n42854), .B(n42855), .Z(n42774) );
  ANDN U52100 ( .B(n42856), .A(n42857), .Z(n42768) );
  XNOR U52101 ( .A(n42759), .B(n42858), .Z(n42764) );
  XNOR U52102 ( .A(n42757), .B(n42761), .Z(n42858) );
  AND U52103 ( .A(n42859), .B(n42860), .Z(n42761) );
  NAND U52104 ( .A(n42861), .B(n42862), .Z(n42860) );
  NAND U52105 ( .A(n42863), .B(n42864), .Z(n42859) );
  AND U52106 ( .A(n42865), .B(n42866), .Z(n42757) );
  NAND U52107 ( .A(n42867), .B(n42868), .Z(n42866) );
  NAND U52108 ( .A(n42869), .B(n42870), .Z(n42865) );
  AND U52109 ( .A(n42871), .B(n42872), .Z(n42759) );
  XOR U52110 ( .A(n42839), .B(n42838), .Z(N61580) );
  XNOR U52111 ( .A(n42856), .B(n42857), .Z(n42838) );
  XNOR U52112 ( .A(n42871), .B(n42872), .Z(n42857) );
  XOR U52113 ( .A(n42868), .B(n42867), .Z(n42872) );
  XOR U52114 ( .A(y[1836]), .B(x[1836]), .Z(n42867) );
  XOR U52115 ( .A(n42870), .B(n42869), .Z(n42868) );
  XOR U52116 ( .A(y[1838]), .B(x[1838]), .Z(n42869) );
  XOR U52117 ( .A(y[1837]), .B(x[1837]), .Z(n42870) );
  XOR U52118 ( .A(n42862), .B(n42861), .Z(n42871) );
  XOR U52119 ( .A(n42864), .B(n42863), .Z(n42861) );
  XOR U52120 ( .A(y[1835]), .B(x[1835]), .Z(n42863) );
  XOR U52121 ( .A(y[1834]), .B(x[1834]), .Z(n42864) );
  XOR U52122 ( .A(y[1833]), .B(x[1833]), .Z(n42862) );
  XNOR U52123 ( .A(n42855), .B(n42854), .Z(n42856) );
  XNOR U52124 ( .A(n42851), .B(n42850), .Z(n42854) );
  XOR U52125 ( .A(n42853), .B(n42852), .Z(n42850) );
  XOR U52126 ( .A(y[1832]), .B(x[1832]), .Z(n42852) );
  XOR U52127 ( .A(y[1831]), .B(x[1831]), .Z(n42853) );
  XOR U52128 ( .A(y[1830]), .B(x[1830]), .Z(n42851) );
  XOR U52129 ( .A(n42845), .B(n42844), .Z(n42855) );
  XOR U52130 ( .A(n42847), .B(n42846), .Z(n42844) );
  XOR U52131 ( .A(y[1829]), .B(x[1829]), .Z(n42846) );
  XOR U52132 ( .A(y[1828]), .B(x[1828]), .Z(n42847) );
  XOR U52133 ( .A(y[1827]), .B(x[1827]), .Z(n42845) );
  XNOR U52134 ( .A(n42821), .B(n42822), .Z(n42839) );
  XNOR U52135 ( .A(n42836), .B(n42837), .Z(n42822) );
  XOR U52136 ( .A(n42833), .B(n42832), .Z(n42837) );
  XOR U52137 ( .A(y[1824]), .B(x[1824]), .Z(n42832) );
  XOR U52138 ( .A(n42835), .B(n42834), .Z(n42833) );
  XOR U52139 ( .A(y[1826]), .B(x[1826]), .Z(n42834) );
  XOR U52140 ( .A(y[1825]), .B(x[1825]), .Z(n42835) );
  XOR U52141 ( .A(n42827), .B(n42826), .Z(n42836) );
  XOR U52142 ( .A(n42829), .B(n42828), .Z(n42826) );
  XOR U52143 ( .A(y[1823]), .B(x[1823]), .Z(n42828) );
  XOR U52144 ( .A(y[1822]), .B(x[1822]), .Z(n42829) );
  XOR U52145 ( .A(y[1821]), .B(x[1821]), .Z(n42827) );
  XNOR U52146 ( .A(n42820), .B(n42819), .Z(n42821) );
  XNOR U52147 ( .A(n42816), .B(n42815), .Z(n42819) );
  XOR U52148 ( .A(n42818), .B(n42817), .Z(n42815) );
  XOR U52149 ( .A(y[1820]), .B(x[1820]), .Z(n42817) );
  XOR U52150 ( .A(y[1819]), .B(x[1819]), .Z(n42818) );
  XOR U52151 ( .A(y[1818]), .B(x[1818]), .Z(n42816) );
  XOR U52152 ( .A(n42810), .B(n42809), .Z(n42820) );
  XOR U52153 ( .A(n42812), .B(n42811), .Z(n42809) );
  XOR U52154 ( .A(y[1817]), .B(x[1817]), .Z(n42811) );
  XOR U52155 ( .A(y[1816]), .B(x[1816]), .Z(n42812) );
  XOR U52156 ( .A(y[1815]), .B(x[1815]), .Z(n42810) );
  NAND U52157 ( .A(n42873), .B(n42874), .Z(N61571) );
  NAND U52158 ( .A(n42875), .B(n42876), .Z(n42874) );
  NANDN U52159 ( .A(n42877), .B(n42878), .Z(n42876) );
  NANDN U52160 ( .A(n42878), .B(n42877), .Z(n42873) );
  XOR U52161 ( .A(n42877), .B(n42879), .Z(N61570) );
  XNOR U52162 ( .A(n42875), .B(n42878), .Z(n42879) );
  NAND U52163 ( .A(n42880), .B(n42881), .Z(n42878) );
  NAND U52164 ( .A(n42882), .B(n42883), .Z(n42881) );
  NANDN U52165 ( .A(n42884), .B(n42885), .Z(n42883) );
  NANDN U52166 ( .A(n42885), .B(n42884), .Z(n42880) );
  AND U52167 ( .A(n42886), .B(n42887), .Z(n42875) );
  NAND U52168 ( .A(n42888), .B(n42889), .Z(n42887) );
  NANDN U52169 ( .A(n42890), .B(n42891), .Z(n42889) );
  NANDN U52170 ( .A(n42891), .B(n42890), .Z(n42886) );
  IV U52171 ( .A(n42892), .Z(n42891) );
  AND U52172 ( .A(n42893), .B(n42894), .Z(n42877) );
  NAND U52173 ( .A(n42895), .B(n42896), .Z(n42894) );
  NANDN U52174 ( .A(n42897), .B(n42898), .Z(n42896) );
  NANDN U52175 ( .A(n42898), .B(n42897), .Z(n42893) );
  XOR U52176 ( .A(n42890), .B(n42899), .Z(N61569) );
  XNOR U52177 ( .A(n42888), .B(n42892), .Z(n42899) );
  XOR U52178 ( .A(n42885), .B(n42900), .Z(n42892) );
  XNOR U52179 ( .A(n42882), .B(n42884), .Z(n42900) );
  AND U52180 ( .A(n42901), .B(n42902), .Z(n42884) );
  NANDN U52181 ( .A(n42903), .B(n42904), .Z(n42902) );
  OR U52182 ( .A(n42905), .B(n42906), .Z(n42904) );
  IV U52183 ( .A(n42907), .Z(n42906) );
  NANDN U52184 ( .A(n42907), .B(n42905), .Z(n42901) );
  AND U52185 ( .A(n42908), .B(n42909), .Z(n42882) );
  NAND U52186 ( .A(n42910), .B(n42911), .Z(n42909) );
  NANDN U52187 ( .A(n42912), .B(n42913), .Z(n42911) );
  NANDN U52188 ( .A(n42913), .B(n42912), .Z(n42908) );
  IV U52189 ( .A(n42914), .Z(n42913) );
  NAND U52190 ( .A(n42915), .B(n42916), .Z(n42885) );
  NANDN U52191 ( .A(n42917), .B(n42918), .Z(n42916) );
  NANDN U52192 ( .A(n42919), .B(n42920), .Z(n42918) );
  NANDN U52193 ( .A(n42920), .B(n42919), .Z(n42915) );
  IV U52194 ( .A(n42921), .Z(n42919) );
  AND U52195 ( .A(n42922), .B(n42923), .Z(n42888) );
  NAND U52196 ( .A(n42924), .B(n42925), .Z(n42923) );
  NANDN U52197 ( .A(n42926), .B(n42927), .Z(n42925) );
  NANDN U52198 ( .A(n42927), .B(n42926), .Z(n42922) );
  XOR U52199 ( .A(n42898), .B(n42928), .Z(n42890) );
  XNOR U52200 ( .A(n42895), .B(n42897), .Z(n42928) );
  AND U52201 ( .A(n42929), .B(n42930), .Z(n42897) );
  NANDN U52202 ( .A(n42931), .B(n42932), .Z(n42930) );
  OR U52203 ( .A(n42933), .B(n42934), .Z(n42932) );
  IV U52204 ( .A(n42935), .Z(n42934) );
  NANDN U52205 ( .A(n42935), .B(n42933), .Z(n42929) );
  AND U52206 ( .A(n42936), .B(n42937), .Z(n42895) );
  NAND U52207 ( .A(n42938), .B(n42939), .Z(n42937) );
  NANDN U52208 ( .A(n42940), .B(n42941), .Z(n42939) );
  NANDN U52209 ( .A(n42941), .B(n42940), .Z(n42936) );
  IV U52210 ( .A(n42942), .Z(n42941) );
  NAND U52211 ( .A(n42943), .B(n42944), .Z(n42898) );
  NANDN U52212 ( .A(n42945), .B(n42946), .Z(n42944) );
  NANDN U52213 ( .A(n42947), .B(n42948), .Z(n42946) );
  NANDN U52214 ( .A(n42948), .B(n42947), .Z(n42943) );
  IV U52215 ( .A(n42949), .Z(n42947) );
  XOR U52216 ( .A(n42924), .B(n42950), .Z(N61568) );
  XNOR U52217 ( .A(n42927), .B(n42926), .Z(n42950) );
  XNOR U52218 ( .A(n42938), .B(n42951), .Z(n42926) );
  XNOR U52219 ( .A(n42942), .B(n42940), .Z(n42951) );
  XOR U52220 ( .A(n42948), .B(n42952), .Z(n42940) );
  XNOR U52221 ( .A(n42945), .B(n42949), .Z(n42952) );
  AND U52222 ( .A(n42953), .B(n42954), .Z(n42949) );
  NAND U52223 ( .A(n42955), .B(n42956), .Z(n42954) );
  NAND U52224 ( .A(n42957), .B(n42958), .Z(n42953) );
  AND U52225 ( .A(n42959), .B(n42960), .Z(n42945) );
  NAND U52226 ( .A(n42961), .B(n42962), .Z(n42960) );
  NAND U52227 ( .A(n42963), .B(n42964), .Z(n42959) );
  NANDN U52228 ( .A(n42965), .B(n42966), .Z(n42948) );
  ANDN U52229 ( .B(n42967), .A(n42968), .Z(n42942) );
  XNOR U52230 ( .A(n42933), .B(n42969), .Z(n42938) );
  XNOR U52231 ( .A(n42931), .B(n42935), .Z(n42969) );
  AND U52232 ( .A(n42970), .B(n42971), .Z(n42935) );
  NAND U52233 ( .A(n42972), .B(n42973), .Z(n42971) );
  NAND U52234 ( .A(n42974), .B(n42975), .Z(n42970) );
  AND U52235 ( .A(n42976), .B(n42977), .Z(n42931) );
  NAND U52236 ( .A(n42978), .B(n42979), .Z(n42977) );
  NAND U52237 ( .A(n42980), .B(n42981), .Z(n42976) );
  AND U52238 ( .A(n42982), .B(n42983), .Z(n42933) );
  NAND U52239 ( .A(n42984), .B(n42985), .Z(n42927) );
  XNOR U52240 ( .A(n42910), .B(n42986), .Z(n42924) );
  XNOR U52241 ( .A(n42914), .B(n42912), .Z(n42986) );
  XOR U52242 ( .A(n42920), .B(n42987), .Z(n42912) );
  XNOR U52243 ( .A(n42917), .B(n42921), .Z(n42987) );
  AND U52244 ( .A(n42988), .B(n42989), .Z(n42921) );
  NAND U52245 ( .A(n42990), .B(n42991), .Z(n42989) );
  NAND U52246 ( .A(n42992), .B(n42993), .Z(n42988) );
  AND U52247 ( .A(n42994), .B(n42995), .Z(n42917) );
  NAND U52248 ( .A(n42996), .B(n42997), .Z(n42995) );
  NAND U52249 ( .A(n42998), .B(n42999), .Z(n42994) );
  NANDN U52250 ( .A(n43000), .B(n43001), .Z(n42920) );
  ANDN U52251 ( .B(n43002), .A(n43003), .Z(n42914) );
  XNOR U52252 ( .A(n42905), .B(n43004), .Z(n42910) );
  XNOR U52253 ( .A(n42903), .B(n42907), .Z(n43004) );
  AND U52254 ( .A(n43005), .B(n43006), .Z(n42907) );
  NAND U52255 ( .A(n43007), .B(n43008), .Z(n43006) );
  NAND U52256 ( .A(n43009), .B(n43010), .Z(n43005) );
  AND U52257 ( .A(n43011), .B(n43012), .Z(n42903) );
  NAND U52258 ( .A(n43013), .B(n43014), .Z(n43012) );
  NAND U52259 ( .A(n43015), .B(n43016), .Z(n43011) );
  AND U52260 ( .A(n43017), .B(n43018), .Z(n42905) );
  XOR U52261 ( .A(n42985), .B(n42984), .Z(N61567) );
  XNOR U52262 ( .A(n43002), .B(n43003), .Z(n42984) );
  XNOR U52263 ( .A(n43017), .B(n43018), .Z(n43003) );
  XOR U52264 ( .A(n43014), .B(n43013), .Z(n43018) );
  XOR U52265 ( .A(y[1812]), .B(x[1812]), .Z(n43013) );
  XOR U52266 ( .A(n43016), .B(n43015), .Z(n43014) );
  XOR U52267 ( .A(y[1814]), .B(x[1814]), .Z(n43015) );
  XOR U52268 ( .A(y[1813]), .B(x[1813]), .Z(n43016) );
  XOR U52269 ( .A(n43008), .B(n43007), .Z(n43017) );
  XOR U52270 ( .A(n43010), .B(n43009), .Z(n43007) );
  XOR U52271 ( .A(y[1811]), .B(x[1811]), .Z(n43009) );
  XOR U52272 ( .A(y[1810]), .B(x[1810]), .Z(n43010) );
  XOR U52273 ( .A(y[1809]), .B(x[1809]), .Z(n43008) );
  XNOR U52274 ( .A(n43001), .B(n43000), .Z(n43002) );
  XNOR U52275 ( .A(n42997), .B(n42996), .Z(n43000) );
  XOR U52276 ( .A(n42999), .B(n42998), .Z(n42996) );
  XOR U52277 ( .A(y[1808]), .B(x[1808]), .Z(n42998) );
  XOR U52278 ( .A(y[1807]), .B(x[1807]), .Z(n42999) );
  XOR U52279 ( .A(y[1806]), .B(x[1806]), .Z(n42997) );
  XOR U52280 ( .A(n42991), .B(n42990), .Z(n43001) );
  XOR U52281 ( .A(n42993), .B(n42992), .Z(n42990) );
  XOR U52282 ( .A(y[1805]), .B(x[1805]), .Z(n42992) );
  XOR U52283 ( .A(y[1804]), .B(x[1804]), .Z(n42993) );
  XOR U52284 ( .A(y[1803]), .B(x[1803]), .Z(n42991) );
  XNOR U52285 ( .A(n42967), .B(n42968), .Z(n42985) );
  XNOR U52286 ( .A(n42982), .B(n42983), .Z(n42968) );
  XOR U52287 ( .A(n42979), .B(n42978), .Z(n42983) );
  XOR U52288 ( .A(y[1800]), .B(x[1800]), .Z(n42978) );
  XOR U52289 ( .A(n42981), .B(n42980), .Z(n42979) );
  XOR U52290 ( .A(y[1802]), .B(x[1802]), .Z(n42980) );
  XOR U52291 ( .A(y[1801]), .B(x[1801]), .Z(n42981) );
  XOR U52292 ( .A(n42973), .B(n42972), .Z(n42982) );
  XOR U52293 ( .A(n42975), .B(n42974), .Z(n42972) );
  XOR U52294 ( .A(y[1799]), .B(x[1799]), .Z(n42974) );
  XOR U52295 ( .A(y[1798]), .B(x[1798]), .Z(n42975) );
  XOR U52296 ( .A(y[1797]), .B(x[1797]), .Z(n42973) );
  XNOR U52297 ( .A(n42966), .B(n42965), .Z(n42967) );
  XNOR U52298 ( .A(n42962), .B(n42961), .Z(n42965) );
  XOR U52299 ( .A(n42964), .B(n42963), .Z(n42961) );
  XOR U52300 ( .A(y[1796]), .B(x[1796]), .Z(n42963) );
  XOR U52301 ( .A(y[1795]), .B(x[1795]), .Z(n42964) );
  XOR U52302 ( .A(y[1794]), .B(x[1794]), .Z(n42962) );
  XOR U52303 ( .A(n42956), .B(n42955), .Z(n42966) );
  XOR U52304 ( .A(n42958), .B(n42957), .Z(n42955) );
  XOR U52305 ( .A(y[1793]), .B(x[1793]), .Z(n42957) );
  XOR U52306 ( .A(y[1792]), .B(x[1792]), .Z(n42958) );
  XOR U52307 ( .A(y[1791]), .B(x[1791]), .Z(n42956) );
  NAND U52308 ( .A(n43019), .B(n43020), .Z(N61558) );
  NAND U52309 ( .A(n43021), .B(n43022), .Z(n43020) );
  NANDN U52310 ( .A(n43023), .B(n43024), .Z(n43022) );
  NANDN U52311 ( .A(n43024), .B(n43023), .Z(n43019) );
  XOR U52312 ( .A(n43023), .B(n43025), .Z(N61557) );
  XNOR U52313 ( .A(n43021), .B(n43024), .Z(n43025) );
  NAND U52314 ( .A(n43026), .B(n43027), .Z(n43024) );
  NAND U52315 ( .A(n43028), .B(n43029), .Z(n43027) );
  NANDN U52316 ( .A(n43030), .B(n43031), .Z(n43029) );
  NANDN U52317 ( .A(n43031), .B(n43030), .Z(n43026) );
  AND U52318 ( .A(n43032), .B(n43033), .Z(n43021) );
  NAND U52319 ( .A(n43034), .B(n43035), .Z(n43033) );
  NANDN U52320 ( .A(n43036), .B(n43037), .Z(n43035) );
  NANDN U52321 ( .A(n43037), .B(n43036), .Z(n43032) );
  IV U52322 ( .A(n43038), .Z(n43037) );
  AND U52323 ( .A(n43039), .B(n43040), .Z(n43023) );
  NAND U52324 ( .A(n43041), .B(n43042), .Z(n43040) );
  NANDN U52325 ( .A(n43043), .B(n43044), .Z(n43042) );
  NANDN U52326 ( .A(n43044), .B(n43043), .Z(n43039) );
  XOR U52327 ( .A(n43036), .B(n43045), .Z(N61556) );
  XNOR U52328 ( .A(n43034), .B(n43038), .Z(n43045) );
  XOR U52329 ( .A(n43031), .B(n43046), .Z(n43038) );
  XNOR U52330 ( .A(n43028), .B(n43030), .Z(n43046) );
  AND U52331 ( .A(n43047), .B(n43048), .Z(n43030) );
  NANDN U52332 ( .A(n43049), .B(n43050), .Z(n43048) );
  OR U52333 ( .A(n43051), .B(n43052), .Z(n43050) );
  IV U52334 ( .A(n43053), .Z(n43052) );
  NANDN U52335 ( .A(n43053), .B(n43051), .Z(n43047) );
  AND U52336 ( .A(n43054), .B(n43055), .Z(n43028) );
  NAND U52337 ( .A(n43056), .B(n43057), .Z(n43055) );
  NANDN U52338 ( .A(n43058), .B(n43059), .Z(n43057) );
  NANDN U52339 ( .A(n43059), .B(n43058), .Z(n43054) );
  IV U52340 ( .A(n43060), .Z(n43059) );
  NAND U52341 ( .A(n43061), .B(n43062), .Z(n43031) );
  NANDN U52342 ( .A(n43063), .B(n43064), .Z(n43062) );
  NANDN U52343 ( .A(n43065), .B(n43066), .Z(n43064) );
  NANDN U52344 ( .A(n43066), .B(n43065), .Z(n43061) );
  IV U52345 ( .A(n43067), .Z(n43065) );
  AND U52346 ( .A(n43068), .B(n43069), .Z(n43034) );
  NAND U52347 ( .A(n43070), .B(n43071), .Z(n43069) );
  NANDN U52348 ( .A(n43072), .B(n43073), .Z(n43071) );
  NANDN U52349 ( .A(n43073), .B(n43072), .Z(n43068) );
  XOR U52350 ( .A(n43044), .B(n43074), .Z(n43036) );
  XNOR U52351 ( .A(n43041), .B(n43043), .Z(n43074) );
  AND U52352 ( .A(n43075), .B(n43076), .Z(n43043) );
  NANDN U52353 ( .A(n43077), .B(n43078), .Z(n43076) );
  OR U52354 ( .A(n43079), .B(n43080), .Z(n43078) );
  IV U52355 ( .A(n43081), .Z(n43080) );
  NANDN U52356 ( .A(n43081), .B(n43079), .Z(n43075) );
  AND U52357 ( .A(n43082), .B(n43083), .Z(n43041) );
  NAND U52358 ( .A(n43084), .B(n43085), .Z(n43083) );
  NANDN U52359 ( .A(n43086), .B(n43087), .Z(n43085) );
  NANDN U52360 ( .A(n43087), .B(n43086), .Z(n43082) );
  IV U52361 ( .A(n43088), .Z(n43087) );
  NAND U52362 ( .A(n43089), .B(n43090), .Z(n43044) );
  NANDN U52363 ( .A(n43091), .B(n43092), .Z(n43090) );
  NANDN U52364 ( .A(n43093), .B(n43094), .Z(n43092) );
  NANDN U52365 ( .A(n43094), .B(n43093), .Z(n43089) );
  IV U52366 ( .A(n43095), .Z(n43093) );
  XOR U52367 ( .A(n43070), .B(n43096), .Z(N61555) );
  XNOR U52368 ( .A(n43073), .B(n43072), .Z(n43096) );
  XNOR U52369 ( .A(n43084), .B(n43097), .Z(n43072) );
  XNOR U52370 ( .A(n43088), .B(n43086), .Z(n43097) );
  XOR U52371 ( .A(n43094), .B(n43098), .Z(n43086) );
  XNOR U52372 ( .A(n43091), .B(n43095), .Z(n43098) );
  AND U52373 ( .A(n43099), .B(n43100), .Z(n43095) );
  NAND U52374 ( .A(n43101), .B(n43102), .Z(n43100) );
  NAND U52375 ( .A(n43103), .B(n43104), .Z(n43099) );
  AND U52376 ( .A(n43105), .B(n43106), .Z(n43091) );
  NAND U52377 ( .A(n43107), .B(n43108), .Z(n43106) );
  NAND U52378 ( .A(n43109), .B(n43110), .Z(n43105) );
  NANDN U52379 ( .A(n43111), .B(n43112), .Z(n43094) );
  ANDN U52380 ( .B(n43113), .A(n43114), .Z(n43088) );
  XNOR U52381 ( .A(n43079), .B(n43115), .Z(n43084) );
  XNOR U52382 ( .A(n43077), .B(n43081), .Z(n43115) );
  AND U52383 ( .A(n43116), .B(n43117), .Z(n43081) );
  NAND U52384 ( .A(n43118), .B(n43119), .Z(n43117) );
  NAND U52385 ( .A(n43120), .B(n43121), .Z(n43116) );
  AND U52386 ( .A(n43122), .B(n43123), .Z(n43077) );
  NAND U52387 ( .A(n43124), .B(n43125), .Z(n43123) );
  NAND U52388 ( .A(n43126), .B(n43127), .Z(n43122) );
  AND U52389 ( .A(n43128), .B(n43129), .Z(n43079) );
  NAND U52390 ( .A(n43130), .B(n43131), .Z(n43073) );
  XNOR U52391 ( .A(n43056), .B(n43132), .Z(n43070) );
  XNOR U52392 ( .A(n43060), .B(n43058), .Z(n43132) );
  XOR U52393 ( .A(n43066), .B(n43133), .Z(n43058) );
  XNOR U52394 ( .A(n43063), .B(n43067), .Z(n43133) );
  AND U52395 ( .A(n43134), .B(n43135), .Z(n43067) );
  NAND U52396 ( .A(n43136), .B(n43137), .Z(n43135) );
  NAND U52397 ( .A(n43138), .B(n43139), .Z(n43134) );
  AND U52398 ( .A(n43140), .B(n43141), .Z(n43063) );
  NAND U52399 ( .A(n43142), .B(n43143), .Z(n43141) );
  NAND U52400 ( .A(n43144), .B(n43145), .Z(n43140) );
  NANDN U52401 ( .A(n43146), .B(n43147), .Z(n43066) );
  ANDN U52402 ( .B(n43148), .A(n43149), .Z(n43060) );
  XNOR U52403 ( .A(n43051), .B(n43150), .Z(n43056) );
  XNOR U52404 ( .A(n43049), .B(n43053), .Z(n43150) );
  AND U52405 ( .A(n43151), .B(n43152), .Z(n43053) );
  NAND U52406 ( .A(n43153), .B(n43154), .Z(n43152) );
  NAND U52407 ( .A(n43155), .B(n43156), .Z(n43151) );
  AND U52408 ( .A(n43157), .B(n43158), .Z(n43049) );
  NAND U52409 ( .A(n43159), .B(n43160), .Z(n43158) );
  NAND U52410 ( .A(n43161), .B(n43162), .Z(n43157) );
  AND U52411 ( .A(n43163), .B(n43164), .Z(n43051) );
  XOR U52412 ( .A(n43131), .B(n43130), .Z(N61554) );
  XNOR U52413 ( .A(n43148), .B(n43149), .Z(n43130) );
  XNOR U52414 ( .A(n43163), .B(n43164), .Z(n43149) );
  XOR U52415 ( .A(n43160), .B(n43159), .Z(n43164) );
  XOR U52416 ( .A(y[1788]), .B(x[1788]), .Z(n43159) );
  XOR U52417 ( .A(n43162), .B(n43161), .Z(n43160) );
  XOR U52418 ( .A(y[1790]), .B(x[1790]), .Z(n43161) );
  XOR U52419 ( .A(y[1789]), .B(x[1789]), .Z(n43162) );
  XOR U52420 ( .A(n43154), .B(n43153), .Z(n43163) );
  XOR U52421 ( .A(n43156), .B(n43155), .Z(n43153) );
  XOR U52422 ( .A(y[1787]), .B(x[1787]), .Z(n43155) );
  XOR U52423 ( .A(y[1786]), .B(x[1786]), .Z(n43156) );
  XOR U52424 ( .A(y[1785]), .B(x[1785]), .Z(n43154) );
  XNOR U52425 ( .A(n43147), .B(n43146), .Z(n43148) );
  XNOR U52426 ( .A(n43143), .B(n43142), .Z(n43146) );
  XOR U52427 ( .A(n43145), .B(n43144), .Z(n43142) );
  XOR U52428 ( .A(y[1784]), .B(x[1784]), .Z(n43144) );
  XOR U52429 ( .A(y[1783]), .B(x[1783]), .Z(n43145) );
  XOR U52430 ( .A(y[1782]), .B(x[1782]), .Z(n43143) );
  XOR U52431 ( .A(n43137), .B(n43136), .Z(n43147) );
  XOR U52432 ( .A(n43139), .B(n43138), .Z(n43136) );
  XOR U52433 ( .A(y[1781]), .B(x[1781]), .Z(n43138) );
  XOR U52434 ( .A(y[1780]), .B(x[1780]), .Z(n43139) );
  XOR U52435 ( .A(y[1779]), .B(x[1779]), .Z(n43137) );
  XNOR U52436 ( .A(n43113), .B(n43114), .Z(n43131) );
  XNOR U52437 ( .A(n43128), .B(n43129), .Z(n43114) );
  XOR U52438 ( .A(n43125), .B(n43124), .Z(n43129) );
  XOR U52439 ( .A(y[1776]), .B(x[1776]), .Z(n43124) );
  XOR U52440 ( .A(n43127), .B(n43126), .Z(n43125) );
  XOR U52441 ( .A(y[1778]), .B(x[1778]), .Z(n43126) );
  XOR U52442 ( .A(y[1777]), .B(x[1777]), .Z(n43127) );
  XOR U52443 ( .A(n43119), .B(n43118), .Z(n43128) );
  XOR U52444 ( .A(n43121), .B(n43120), .Z(n43118) );
  XOR U52445 ( .A(y[1775]), .B(x[1775]), .Z(n43120) );
  XOR U52446 ( .A(y[1774]), .B(x[1774]), .Z(n43121) );
  XOR U52447 ( .A(y[1773]), .B(x[1773]), .Z(n43119) );
  XNOR U52448 ( .A(n43112), .B(n43111), .Z(n43113) );
  XNOR U52449 ( .A(n43108), .B(n43107), .Z(n43111) );
  XOR U52450 ( .A(n43110), .B(n43109), .Z(n43107) );
  XOR U52451 ( .A(y[1772]), .B(x[1772]), .Z(n43109) );
  XOR U52452 ( .A(y[1771]), .B(x[1771]), .Z(n43110) );
  XOR U52453 ( .A(y[1770]), .B(x[1770]), .Z(n43108) );
  XOR U52454 ( .A(n43102), .B(n43101), .Z(n43112) );
  XOR U52455 ( .A(n43104), .B(n43103), .Z(n43101) );
  XOR U52456 ( .A(y[1769]), .B(x[1769]), .Z(n43103) );
  XOR U52457 ( .A(y[1768]), .B(x[1768]), .Z(n43104) );
  XOR U52458 ( .A(y[1767]), .B(x[1767]), .Z(n43102) );
  NAND U52459 ( .A(n43165), .B(n43166), .Z(N61545) );
  NAND U52460 ( .A(n43167), .B(n43168), .Z(n43166) );
  NANDN U52461 ( .A(n43169), .B(n43170), .Z(n43168) );
  NANDN U52462 ( .A(n43170), .B(n43169), .Z(n43165) );
  XOR U52463 ( .A(n43169), .B(n43171), .Z(N61544) );
  XNOR U52464 ( .A(n43167), .B(n43170), .Z(n43171) );
  NAND U52465 ( .A(n43172), .B(n43173), .Z(n43170) );
  NAND U52466 ( .A(n43174), .B(n43175), .Z(n43173) );
  NANDN U52467 ( .A(n43176), .B(n43177), .Z(n43175) );
  NANDN U52468 ( .A(n43177), .B(n43176), .Z(n43172) );
  AND U52469 ( .A(n43178), .B(n43179), .Z(n43167) );
  NAND U52470 ( .A(n43180), .B(n43181), .Z(n43179) );
  NANDN U52471 ( .A(n43182), .B(n43183), .Z(n43181) );
  NANDN U52472 ( .A(n43183), .B(n43182), .Z(n43178) );
  IV U52473 ( .A(n43184), .Z(n43183) );
  AND U52474 ( .A(n43185), .B(n43186), .Z(n43169) );
  NAND U52475 ( .A(n43187), .B(n43188), .Z(n43186) );
  NANDN U52476 ( .A(n43189), .B(n43190), .Z(n43188) );
  NANDN U52477 ( .A(n43190), .B(n43189), .Z(n43185) );
  XOR U52478 ( .A(n43182), .B(n43191), .Z(N61543) );
  XNOR U52479 ( .A(n43180), .B(n43184), .Z(n43191) );
  XOR U52480 ( .A(n43177), .B(n43192), .Z(n43184) );
  XNOR U52481 ( .A(n43174), .B(n43176), .Z(n43192) );
  AND U52482 ( .A(n43193), .B(n43194), .Z(n43176) );
  NANDN U52483 ( .A(n43195), .B(n43196), .Z(n43194) );
  OR U52484 ( .A(n43197), .B(n43198), .Z(n43196) );
  IV U52485 ( .A(n43199), .Z(n43198) );
  NANDN U52486 ( .A(n43199), .B(n43197), .Z(n43193) );
  AND U52487 ( .A(n43200), .B(n43201), .Z(n43174) );
  NAND U52488 ( .A(n43202), .B(n43203), .Z(n43201) );
  NANDN U52489 ( .A(n43204), .B(n43205), .Z(n43203) );
  NANDN U52490 ( .A(n43205), .B(n43204), .Z(n43200) );
  IV U52491 ( .A(n43206), .Z(n43205) );
  NAND U52492 ( .A(n43207), .B(n43208), .Z(n43177) );
  NANDN U52493 ( .A(n43209), .B(n43210), .Z(n43208) );
  NANDN U52494 ( .A(n43211), .B(n43212), .Z(n43210) );
  NANDN U52495 ( .A(n43212), .B(n43211), .Z(n43207) );
  IV U52496 ( .A(n43213), .Z(n43211) );
  AND U52497 ( .A(n43214), .B(n43215), .Z(n43180) );
  NAND U52498 ( .A(n43216), .B(n43217), .Z(n43215) );
  NANDN U52499 ( .A(n43218), .B(n43219), .Z(n43217) );
  NANDN U52500 ( .A(n43219), .B(n43218), .Z(n43214) );
  XOR U52501 ( .A(n43190), .B(n43220), .Z(n43182) );
  XNOR U52502 ( .A(n43187), .B(n43189), .Z(n43220) );
  AND U52503 ( .A(n43221), .B(n43222), .Z(n43189) );
  NANDN U52504 ( .A(n43223), .B(n43224), .Z(n43222) );
  OR U52505 ( .A(n43225), .B(n43226), .Z(n43224) );
  IV U52506 ( .A(n43227), .Z(n43226) );
  NANDN U52507 ( .A(n43227), .B(n43225), .Z(n43221) );
  AND U52508 ( .A(n43228), .B(n43229), .Z(n43187) );
  NAND U52509 ( .A(n43230), .B(n43231), .Z(n43229) );
  NANDN U52510 ( .A(n43232), .B(n43233), .Z(n43231) );
  NANDN U52511 ( .A(n43233), .B(n43232), .Z(n43228) );
  IV U52512 ( .A(n43234), .Z(n43233) );
  NAND U52513 ( .A(n43235), .B(n43236), .Z(n43190) );
  NANDN U52514 ( .A(n43237), .B(n43238), .Z(n43236) );
  NANDN U52515 ( .A(n43239), .B(n43240), .Z(n43238) );
  NANDN U52516 ( .A(n43240), .B(n43239), .Z(n43235) );
  IV U52517 ( .A(n43241), .Z(n43239) );
  XOR U52518 ( .A(n43216), .B(n43242), .Z(N61542) );
  XNOR U52519 ( .A(n43219), .B(n43218), .Z(n43242) );
  XNOR U52520 ( .A(n43230), .B(n43243), .Z(n43218) );
  XNOR U52521 ( .A(n43234), .B(n43232), .Z(n43243) );
  XOR U52522 ( .A(n43240), .B(n43244), .Z(n43232) );
  XNOR U52523 ( .A(n43237), .B(n43241), .Z(n43244) );
  AND U52524 ( .A(n43245), .B(n43246), .Z(n43241) );
  NAND U52525 ( .A(n43247), .B(n43248), .Z(n43246) );
  NAND U52526 ( .A(n43249), .B(n43250), .Z(n43245) );
  AND U52527 ( .A(n43251), .B(n43252), .Z(n43237) );
  NAND U52528 ( .A(n43253), .B(n43254), .Z(n43252) );
  NAND U52529 ( .A(n43255), .B(n43256), .Z(n43251) );
  NANDN U52530 ( .A(n43257), .B(n43258), .Z(n43240) );
  ANDN U52531 ( .B(n43259), .A(n43260), .Z(n43234) );
  XNOR U52532 ( .A(n43225), .B(n43261), .Z(n43230) );
  XNOR U52533 ( .A(n43223), .B(n43227), .Z(n43261) );
  AND U52534 ( .A(n43262), .B(n43263), .Z(n43227) );
  NAND U52535 ( .A(n43264), .B(n43265), .Z(n43263) );
  NAND U52536 ( .A(n43266), .B(n43267), .Z(n43262) );
  AND U52537 ( .A(n43268), .B(n43269), .Z(n43223) );
  NAND U52538 ( .A(n43270), .B(n43271), .Z(n43269) );
  NAND U52539 ( .A(n43272), .B(n43273), .Z(n43268) );
  AND U52540 ( .A(n43274), .B(n43275), .Z(n43225) );
  NAND U52541 ( .A(n43276), .B(n43277), .Z(n43219) );
  XNOR U52542 ( .A(n43202), .B(n43278), .Z(n43216) );
  XNOR U52543 ( .A(n43206), .B(n43204), .Z(n43278) );
  XOR U52544 ( .A(n43212), .B(n43279), .Z(n43204) );
  XNOR U52545 ( .A(n43209), .B(n43213), .Z(n43279) );
  AND U52546 ( .A(n43280), .B(n43281), .Z(n43213) );
  NAND U52547 ( .A(n43282), .B(n43283), .Z(n43281) );
  NAND U52548 ( .A(n43284), .B(n43285), .Z(n43280) );
  AND U52549 ( .A(n43286), .B(n43287), .Z(n43209) );
  NAND U52550 ( .A(n43288), .B(n43289), .Z(n43287) );
  NAND U52551 ( .A(n43290), .B(n43291), .Z(n43286) );
  NANDN U52552 ( .A(n43292), .B(n43293), .Z(n43212) );
  ANDN U52553 ( .B(n43294), .A(n43295), .Z(n43206) );
  XNOR U52554 ( .A(n43197), .B(n43296), .Z(n43202) );
  XNOR U52555 ( .A(n43195), .B(n43199), .Z(n43296) );
  AND U52556 ( .A(n43297), .B(n43298), .Z(n43199) );
  NAND U52557 ( .A(n43299), .B(n43300), .Z(n43298) );
  NAND U52558 ( .A(n43301), .B(n43302), .Z(n43297) );
  AND U52559 ( .A(n43303), .B(n43304), .Z(n43195) );
  NAND U52560 ( .A(n43305), .B(n43306), .Z(n43304) );
  NAND U52561 ( .A(n43307), .B(n43308), .Z(n43303) );
  AND U52562 ( .A(n43309), .B(n43310), .Z(n43197) );
  XOR U52563 ( .A(n43277), .B(n43276), .Z(N61541) );
  XNOR U52564 ( .A(n43294), .B(n43295), .Z(n43276) );
  XNOR U52565 ( .A(n43309), .B(n43310), .Z(n43295) );
  XOR U52566 ( .A(n43306), .B(n43305), .Z(n43310) );
  XOR U52567 ( .A(y[1764]), .B(x[1764]), .Z(n43305) );
  XOR U52568 ( .A(n43308), .B(n43307), .Z(n43306) );
  XOR U52569 ( .A(y[1766]), .B(x[1766]), .Z(n43307) );
  XOR U52570 ( .A(y[1765]), .B(x[1765]), .Z(n43308) );
  XOR U52571 ( .A(n43300), .B(n43299), .Z(n43309) );
  XOR U52572 ( .A(n43302), .B(n43301), .Z(n43299) );
  XOR U52573 ( .A(y[1763]), .B(x[1763]), .Z(n43301) );
  XOR U52574 ( .A(y[1762]), .B(x[1762]), .Z(n43302) );
  XOR U52575 ( .A(y[1761]), .B(x[1761]), .Z(n43300) );
  XNOR U52576 ( .A(n43293), .B(n43292), .Z(n43294) );
  XNOR U52577 ( .A(n43289), .B(n43288), .Z(n43292) );
  XOR U52578 ( .A(n43291), .B(n43290), .Z(n43288) );
  XOR U52579 ( .A(y[1760]), .B(x[1760]), .Z(n43290) );
  XOR U52580 ( .A(y[1759]), .B(x[1759]), .Z(n43291) );
  XOR U52581 ( .A(y[1758]), .B(x[1758]), .Z(n43289) );
  XOR U52582 ( .A(n43283), .B(n43282), .Z(n43293) );
  XOR U52583 ( .A(n43285), .B(n43284), .Z(n43282) );
  XOR U52584 ( .A(y[1757]), .B(x[1757]), .Z(n43284) );
  XOR U52585 ( .A(y[1756]), .B(x[1756]), .Z(n43285) );
  XOR U52586 ( .A(y[1755]), .B(x[1755]), .Z(n43283) );
  XNOR U52587 ( .A(n43259), .B(n43260), .Z(n43277) );
  XNOR U52588 ( .A(n43274), .B(n43275), .Z(n43260) );
  XOR U52589 ( .A(n43271), .B(n43270), .Z(n43275) );
  XOR U52590 ( .A(y[1752]), .B(x[1752]), .Z(n43270) );
  XOR U52591 ( .A(n43273), .B(n43272), .Z(n43271) );
  XOR U52592 ( .A(y[1754]), .B(x[1754]), .Z(n43272) );
  XOR U52593 ( .A(y[1753]), .B(x[1753]), .Z(n43273) );
  XOR U52594 ( .A(n43265), .B(n43264), .Z(n43274) );
  XOR U52595 ( .A(n43267), .B(n43266), .Z(n43264) );
  XOR U52596 ( .A(y[1751]), .B(x[1751]), .Z(n43266) );
  XOR U52597 ( .A(y[1750]), .B(x[1750]), .Z(n43267) );
  XOR U52598 ( .A(y[1749]), .B(x[1749]), .Z(n43265) );
  XNOR U52599 ( .A(n43258), .B(n43257), .Z(n43259) );
  XNOR U52600 ( .A(n43254), .B(n43253), .Z(n43257) );
  XOR U52601 ( .A(n43256), .B(n43255), .Z(n43253) );
  XOR U52602 ( .A(y[1748]), .B(x[1748]), .Z(n43255) );
  XOR U52603 ( .A(y[1747]), .B(x[1747]), .Z(n43256) );
  XOR U52604 ( .A(y[1746]), .B(x[1746]), .Z(n43254) );
  XOR U52605 ( .A(n43248), .B(n43247), .Z(n43258) );
  XOR U52606 ( .A(n43250), .B(n43249), .Z(n43247) );
  XOR U52607 ( .A(y[1745]), .B(x[1745]), .Z(n43249) );
  XOR U52608 ( .A(y[1744]), .B(x[1744]), .Z(n43250) );
  XOR U52609 ( .A(y[1743]), .B(x[1743]), .Z(n43248) );
  NAND U52610 ( .A(n43311), .B(n43312), .Z(N61532) );
  NAND U52611 ( .A(n43313), .B(n43314), .Z(n43312) );
  NANDN U52612 ( .A(n43315), .B(n43316), .Z(n43314) );
  NANDN U52613 ( .A(n43316), .B(n43315), .Z(n43311) );
  XOR U52614 ( .A(n43315), .B(n43317), .Z(N61531) );
  XNOR U52615 ( .A(n43313), .B(n43316), .Z(n43317) );
  NAND U52616 ( .A(n43318), .B(n43319), .Z(n43316) );
  NAND U52617 ( .A(n43320), .B(n43321), .Z(n43319) );
  NANDN U52618 ( .A(n43322), .B(n43323), .Z(n43321) );
  NANDN U52619 ( .A(n43323), .B(n43322), .Z(n43318) );
  AND U52620 ( .A(n43324), .B(n43325), .Z(n43313) );
  NAND U52621 ( .A(n43326), .B(n43327), .Z(n43325) );
  NANDN U52622 ( .A(n43328), .B(n43329), .Z(n43327) );
  NANDN U52623 ( .A(n43329), .B(n43328), .Z(n43324) );
  IV U52624 ( .A(n43330), .Z(n43329) );
  AND U52625 ( .A(n43331), .B(n43332), .Z(n43315) );
  NAND U52626 ( .A(n43333), .B(n43334), .Z(n43332) );
  NANDN U52627 ( .A(n43335), .B(n43336), .Z(n43334) );
  NANDN U52628 ( .A(n43336), .B(n43335), .Z(n43331) );
  XOR U52629 ( .A(n43328), .B(n43337), .Z(N61530) );
  XNOR U52630 ( .A(n43326), .B(n43330), .Z(n43337) );
  XOR U52631 ( .A(n43323), .B(n43338), .Z(n43330) );
  XNOR U52632 ( .A(n43320), .B(n43322), .Z(n43338) );
  AND U52633 ( .A(n43339), .B(n43340), .Z(n43322) );
  NANDN U52634 ( .A(n43341), .B(n43342), .Z(n43340) );
  OR U52635 ( .A(n43343), .B(n43344), .Z(n43342) );
  IV U52636 ( .A(n43345), .Z(n43344) );
  NANDN U52637 ( .A(n43345), .B(n43343), .Z(n43339) );
  AND U52638 ( .A(n43346), .B(n43347), .Z(n43320) );
  NAND U52639 ( .A(n43348), .B(n43349), .Z(n43347) );
  NANDN U52640 ( .A(n43350), .B(n43351), .Z(n43349) );
  NANDN U52641 ( .A(n43351), .B(n43350), .Z(n43346) );
  IV U52642 ( .A(n43352), .Z(n43351) );
  NAND U52643 ( .A(n43353), .B(n43354), .Z(n43323) );
  NANDN U52644 ( .A(n43355), .B(n43356), .Z(n43354) );
  NANDN U52645 ( .A(n43357), .B(n43358), .Z(n43356) );
  NANDN U52646 ( .A(n43358), .B(n43357), .Z(n43353) );
  IV U52647 ( .A(n43359), .Z(n43357) );
  AND U52648 ( .A(n43360), .B(n43361), .Z(n43326) );
  NAND U52649 ( .A(n43362), .B(n43363), .Z(n43361) );
  NANDN U52650 ( .A(n43364), .B(n43365), .Z(n43363) );
  NANDN U52651 ( .A(n43365), .B(n43364), .Z(n43360) );
  XOR U52652 ( .A(n43336), .B(n43366), .Z(n43328) );
  XNOR U52653 ( .A(n43333), .B(n43335), .Z(n43366) );
  AND U52654 ( .A(n43367), .B(n43368), .Z(n43335) );
  NANDN U52655 ( .A(n43369), .B(n43370), .Z(n43368) );
  OR U52656 ( .A(n43371), .B(n43372), .Z(n43370) );
  IV U52657 ( .A(n43373), .Z(n43372) );
  NANDN U52658 ( .A(n43373), .B(n43371), .Z(n43367) );
  AND U52659 ( .A(n43374), .B(n43375), .Z(n43333) );
  NAND U52660 ( .A(n43376), .B(n43377), .Z(n43375) );
  NANDN U52661 ( .A(n43378), .B(n43379), .Z(n43377) );
  NANDN U52662 ( .A(n43379), .B(n43378), .Z(n43374) );
  IV U52663 ( .A(n43380), .Z(n43379) );
  NAND U52664 ( .A(n43381), .B(n43382), .Z(n43336) );
  NANDN U52665 ( .A(n43383), .B(n43384), .Z(n43382) );
  NANDN U52666 ( .A(n43385), .B(n43386), .Z(n43384) );
  NANDN U52667 ( .A(n43386), .B(n43385), .Z(n43381) );
  IV U52668 ( .A(n43387), .Z(n43385) );
  XOR U52669 ( .A(n43362), .B(n43388), .Z(N61529) );
  XNOR U52670 ( .A(n43365), .B(n43364), .Z(n43388) );
  XNOR U52671 ( .A(n43376), .B(n43389), .Z(n43364) );
  XNOR U52672 ( .A(n43380), .B(n43378), .Z(n43389) );
  XOR U52673 ( .A(n43386), .B(n43390), .Z(n43378) );
  XNOR U52674 ( .A(n43383), .B(n43387), .Z(n43390) );
  AND U52675 ( .A(n43391), .B(n43392), .Z(n43387) );
  NAND U52676 ( .A(n43393), .B(n43394), .Z(n43392) );
  NAND U52677 ( .A(n43395), .B(n43396), .Z(n43391) );
  AND U52678 ( .A(n43397), .B(n43398), .Z(n43383) );
  NAND U52679 ( .A(n43399), .B(n43400), .Z(n43398) );
  NAND U52680 ( .A(n43401), .B(n43402), .Z(n43397) );
  NANDN U52681 ( .A(n43403), .B(n43404), .Z(n43386) );
  ANDN U52682 ( .B(n43405), .A(n43406), .Z(n43380) );
  XNOR U52683 ( .A(n43371), .B(n43407), .Z(n43376) );
  XNOR U52684 ( .A(n43369), .B(n43373), .Z(n43407) );
  AND U52685 ( .A(n43408), .B(n43409), .Z(n43373) );
  NAND U52686 ( .A(n43410), .B(n43411), .Z(n43409) );
  NAND U52687 ( .A(n43412), .B(n43413), .Z(n43408) );
  AND U52688 ( .A(n43414), .B(n43415), .Z(n43369) );
  NAND U52689 ( .A(n43416), .B(n43417), .Z(n43415) );
  NAND U52690 ( .A(n43418), .B(n43419), .Z(n43414) );
  AND U52691 ( .A(n43420), .B(n43421), .Z(n43371) );
  NAND U52692 ( .A(n43422), .B(n43423), .Z(n43365) );
  XNOR U52693 ( .A(n43348), .B(n43424), .Z(n43362) );
  XNOR U52694 ( .A(n43352), .B(n43350), .Z(n43424) );
  XOR U52695 ( .A(n43358), .B(n43425), .Z(n43350) );
  XNOR U52696 ( .A(n43355), .B(n43359), .Z(n43425) );
  AND U52697 ( .A(n43426), .B(n43427), .Z(n43359) );
  NAND U52698 ( .A(n43428), .B(n43429), .Z(n43427) );
  NAND U52699 ( .A(n43430), .B(n43431), .Z(n43426) );
  AND U52700 ( .A(n43432), .B(n43433), .Z(n43355) );
  NAND U52701 ( .A(n43434), .B(n43435), .Z(n43433) );
  NAND U52702 ( .A(n43436), .B(n43437), .Z(n43432) );
  NANDN U52703 ( .A(n43438), .B(n43439), .Z(n43358) );
  ANDN U52704 ( .B(n43440), .A(n43441), .Z(n43352) );
  XNOR U52705 ( .A(n43343), .B(n43442), .Z(n43348) );
  XNOR U52706 ( .A(n43341), .B(n43345), .Z(n43442) );
  AND U52707 ( .A(n43443), .B(n43444), .Z(n43345) );
  NAND U52708 ( .A(n43445), .B(n43446), .Z(n43444) );
  NAND U52709 ( .A(n43447), .B(n43448), .Z(n43443) );
  AND U52710 ( .A(n43449), .B(n43450), .Z(n43341) );
  NAND U52711 ( .A(n43451), .B(n43452), .Z(n43450) );
  NAND U52712 ( .A(n43453), .B(n43454), .Z(n43449) );
  AND U52713 ( .A(n43455), .B(n43456), .Z(n43343) );
  XOR U52714 ( .A(n43423), .B(n43422), .Z(N61528) );
  XNOR U52715 ( .A(n43440), .B(n43441), .Z(n43422) );
  XNOR U52716 ( .A(n43455), .B(n43456), .Z(n43441) );
  XOR U52717 ( .A(n43452), .B(n43451), .Z(n43456) );
  XOR U52718 ( .A(y[1740]), .B(x[1740]), .Z(n43451) );
  XOR U52719 ( .A(n43454), .B(n43453), .Z(n43452) );
  XOR U52720 ( .A(y[1742]), .B(x[1742]), .Z(n43453) );
  XOR U52721 ( .A(y[1741]), .B(x[1741]), .Z(n43454) );
  XOR U52722 ( .A(n43446), .B(n43445), .Z(n43455) );
  XOR U52723 ( .A(n43448), .B(n43447), .Z(n43445) );
  XOR U52724 ( .A(y[1739]), .B(x[1739]), .Z(n43447) );
  XOR U52725 ( .A(y[1738]), .B(x[1738]), .Z(n43448) );
  XOR U52726 ( .A(y[1737]), .B(x[1737]), .Z(n43446) );
  XNOR U52727 ( .A(n43439), .B(n43438), .Z(n43440) );
  XNOR U52728 ( .A(n43435), .B(n43434), .Z(n43438) );
  XOR U52729 ( .A(n43437), .B(n43436), .Z(n43434) );
  XOR U52730 ( .A(y[1736]), .B(x[1736]), .Z(n43436) );
  XOR U52731 ( .A(y[1735]), .B(x[1735]), .Z(n43437) );
  XOR U52732 ( .A(y[1734]), .B(x[1734]), .Z(n43435) );
  XOR U52733 ( .A(n43429), .B(n43428), .Z(n43439) );
  XOR U52734 ( .A(n43431), .B(n43430), .Z(n43428) );
  XOR U52735 ( .A(y[1733]), .B(x[1733]), .Z(n43430) );
  XOR U52736 ( .A(y[1732]), .B(x[1732]), .Z(n43431) );
  XOR U52737 ( .A(y[1731]), .B(x[1731]), .Z(n43429) );
  XNOR U52738 ( .A(n43405), .B(n43406), .Z(n43423) );
  XNOR U52739 ( .A(n43420), .B(n43421), .Z(n43406) );
  XOR U52740 ( .A(n43417), .B(n43416), .Z(n43421) );
  XOR U52741 ( .A(y[1728]), .B(x[1728]), .Z(n43416) );
  XOR U52742 ( .A(n43419), .B(n43418), .Z(n43417) );
  XOR U52743 ( .A(y[1730]), .B(x[1730]), .Z(n43418) );
  XOR U52744 ( .A(y[1729]), .B(x[1729]), .Z(n43419) );
  XOR U52745 ( .A(n43411), .B(n43410), .Z(n43420) );
  XOR U52746 ( .A(n43413), .B(n43412), .Z(n43410) );
  XOR U52747 ( .A(y[1727]), .B(x[1727]), .Z(n43412) );
  XOR U52748 ( .A(y[1726]), .B(x[1726]), .Z(n43413) );
  XOR U52749 ( .A(y[1725]), .B(x[1725]), .Z(n43411) );
  XNOR U52750 ( .A(n43404), .B(n43403), .Z(n43405) );
  XNOR U52751 ( .A(n43400), .B(n43399), .Z(n43403) );
  XOR U52752 ( .A(n43402), .B(n43401), .Z(n43399) );
  XOR U52753 ( .A(y[1724]), .B(x[1724]), .Z(n43401) );
  XOR U52754 ( .A(y[1723]), .B(x[1723]), .Z(n43402) );
  XOR U52755 ( .A(y[1722]), .B(x[1722]), .Z(n43400) );
  XOR U52756 ( .A(n43394), .B(n43393), .Z(n43404) );
  XOR U52757 ( .A(n43396), .B(n43395), .Z(n43393) );
  XOR U52758 ( .A(y[1721]), .B(x[1721]), .Z(n43395) );
  XOR U52759 ( .A(y[1720]), .B(x[1720]), .Z(n43396) );
  XOR U52760 ( .A(y[1719]), .B(x[1719]), .Z(n43394) );
  NAND U52761 ( .A(n43457), .B(n43458), .Z(N61519) );
  NAND U52762 ( .A(n43459), .B(n43460), .Z(n43458) );
  NANDN U52763 ( .A(n43461), .B(n43462), .Z(n43460) );
  NANDN U52764 ( .A(n43462), .B(n43461), .Z(n43457) );
  XOR U52765 ( .A(n43461), .B(n43463), .Z(N61518) );
  XNOR U52766 ( .A(n43459), .B(n43462), .Z(n43463) );
  NAND U52767 ( .A(n43464), .B(n43465), .Z(n43462) );
  NAND U52768 ( .A(n43466), .B(n43467), .Z(n43465) );
  NANDN U52769 ( .A(n43468), .B(n43469), .Z(n43467) );
  NANDN U52770 ( .A(n43469), .B(n43468), .Z(n43464) );
  AND U52771 ( .A(n43470), .B(n43471), .Z(n43459) );
  NAND U52772 ( .A(n43472), .B(n43473), .Z(n43471) );
  NANDN U52773 ( .A(n43474), .B(n43475), .Z(n43473) );
  NANDN U52774 ( .A(n43475), .B(n43474), .Z(n43470) );
  IV U52775 ( .A(n43476), .Z(n43475) );
  AND U52776 ( .A(n43477), .B(n43478), .Z(n43461) );
  NAND U52777 ( .A(n43479), .B(n43480), .Z(n43478) );
  NANDN U52778 ( .A(n43481), .B(n43482), .Z(n43480) );
  NANDN U52779 ( .A(n43482), .B(n43481), .Z(n43477) );
  XOR U52780 ( .A(n43474), .B(n43483), .Z(N61517) );
  XNOR U52781 ( .A(n43472), .B(n43476), .Z(n43483) );
  XOR U52782 ( .A(n43469), .B(n43484), .Z(n43476) );
  XNOR U52783 ( .A(n43466), .B(n43468), .Z(n43484) );
  AND U52784 ( .A(n43485), .B(n43486), .Z(n43468) );
  NANDN U52785 ( .A(n43487), .B(n43488), .Z(n43486) );
  OR U52786 ( .A(n43489), .B(n43490), .Z(n43488) );
  IV U52787 ( .A(n43491), .Z(n43490) );
  NANDN U52788 ( .A(n43491), .B(n43489), .Z(n43485) );
  AND U52789 ( .A(n43492), .B(n43493), .Z(n43466) );
  NAND U52790 ( .A(n43494), .B(n43495), .Z(n43493) );
  NANDN U52791 ( .A(n43496), .B(n43497), .Z(n43495) );
  NANDN U52792 ( .A(n43497), .B(n43496), .Z(n43492) );
  IV U52793 ( .A(n43498), .Z(n43497) );
  NAND U52794 ( .A(n43499), .B(n43500), .Z(n43469) );
  NANDN U52795 ( .A(n43501), .B(n43502), .Z(n43500) );
  NANDN U52796 ( .A(n43503), .B(n43504), .Z(n43502) );
  NANDN U52797 ( .A(n43504), .B(n43503), .Z(n43499) );
  IV U52798 ( .A(n43505), .Z(n43503) );
  AND U52799 ( .A(n43506), .B(n43507), .Z(n43472) );
  NAND U52800 ( .A(n43508), .B(n43509), .Z(n43507) );
  NANDN U52801 ( .A(n43510), .B(n43511), .Z(n43509) );
  NANDN U52802 ( .A(n43511), .B(n43510), .Z(n43506) );
  XOR U52803 ( .A(n43482), .B(n43512), .Z(n43474) );
  XNOR U52804 ( .A(n43479), .B(n43481), .Z(n43512) );
  AND U52805 ( .A(n43513), .B(n43514), .Z(n43481) );
  NANDN U52806 ( .A(n43515), .B(n43516), .Z(n43514) );
  OR U52807 ( .A(n43517), .B(n43518), .Z(n43516) );
  IV U52808 ( .A(n43519), .Z(n43518) );
  NANDN U52809 ( .A(n43519), .B(n43517), .Z(n43513) );
  AND U52810 ( .A(n43520), .B(n43521), .Z(n43479) );
  NAND U52811 ( .A(n43522), .B(n43523), .Z(n43521) );
  NANDN U52812 ( .A(n43524), .B(n43525), .Z(n43523) );
  NANDN U52813 ( .A(n43525), .B(n43524), .Z(n43520) );
  IV U52814 ( .A(n43526), .Z(n43525) );
  NAND U52815 ( .A(n43527), .B(n43528), .Z(n43482) );
  NANDN U52816 ( .A(n43529), .B(n43530), .Z(n43528) );
  NANDN U52817 ( .A(n43531), .B(n43532), .Z(n43530) );
  NANDN U52818 ( .A(n43532), .B(n43531), .Z(n43527) );
  IV U52819 ( .A(n43533), .Z(n43531) );
  XOR U52820 ( .A(n43508), .B(n43534), .Z(N61516) );
  XNOR U52821 ( .A(n43511), .B(n43510), .Z(n43534) );
  XNOR U52822 ( .A(n43522), .B(n43535), .Z(n43510) );
  XNOR U52823 ( .A(n43526), .B(n43524), .Z(n43535) );
  XOR U52824 ( .A(n43532), .B(n43536), .Z(n43524) );
  XNOR U52825 ( .A(n43529), .B(n43533), .Z(n43536) );
  AND U52826 ( .A(n43537), .B(n43538), .Z(n43533) );
  NAND U52827 ( .A(n43539), .B(n43540), .Z(n43538) );
  NAND U52828 ( .A(n43541), .B(n43542), .Z(n43537) );
  AND U52829 ( .A(n43543), .B(n43544), .Z(n43529) );
  NAND U52830 ( .A(n43545), .B(n43546), .Z(n43544) );
  NAND U52831 ( .A(n43547), .B(n43548), .Z(n43543) );
  NANDN U52832 ( .A(n43549), .B(n43550), .Z(n43532) );
  ANDN U52833 ( .B(n43551), .A(n43552), .Z(n43526) );
  XNOR U52834 ( .A(n43517), .B(n43553), .Z(n43522) );
  XNOR U52835 ( .A(n43515), .B(n43519), .Z(n43553) );
  AND U52836 ( .A(n43554), .B(n43555), .Z(n43519) );
  NAND U52837 ( .A(n43556), .B(n43557), .Z(n43555) );
  NAND U52838 ( .A(n43558), .B(n43559), .Z(n43554) );
  AND U52839 ( .A(n43560), .B(n43561), .Z(n43515) );
  NAND U52840 ( .A(n43562), .B(n43563), .Z(n43561) );
  NAND U52841 ( .A(n43564), .B(n43565), .Z(n43560) );
  AND U52842 ( .A(n43566), .B(n43567), .Z(n43517) );
  NAND U52843 ( .A(n43568), .B(n43569), .Z(n43511) );
  XNOR U52844 ( .A(n43494), .B(n43570), .Z(n43508) );
  XNOR U52845 ( .A(n43498), .B(n43496), .Z(n43570) );
  XOR U52846 ( .A(n43504), .B(n43571), .Z(n43496) );
  XNOR U52847 ( .A(n43501), .B(n43505), .Z(n43571) );
  AND U52848 ( .A(n43572), .B(n43573), .Z(n43505) );
  NAND U52849 ( .A(n43574), .B(n43575), .Z(n43573) );
  NAND U52850 ( .A(n43576), .B(n43577), .Z(n43572) );
  AND U52851 ( .A(n43578), .B(n43579), .Z(n43501) );
  NAND U52852 ( .A(n43580), .B(n43581), .Z(n43579) );
  NAND U52853 ( .A(n43582), .B(n43583), .Z(n43578) );
  NANDN U52854 ( .A(n43584), .B(n43585), .Z(n43504) );
  ANDN U52855 ( .B(n43586), .A(n43587), .Z(n43498) );
  XNOR U52856 ( .A(n43489), .B(n43588), .Z(n43494) );
  XNOR U52857 ( .A(n43487), .B(n43491), .Z(n43588) );
  AND U52858 ( .A(n43589), .B(n43590), .Z(n43491) );
  NAND U52859 ( .A(n43591), .B(n43592), .Z(n43590) );
  NAND U52860 ( .A(n43593), .B(n43594), .Z(n43589) );
  AND U52861 ( .A(n43595), .B(n43596), .Z(n43487) );
  NAND U52862 ( .A(n43597), .B(n43598), .Z(n43596) );
  NAND U52863 ( .A(n43599), .B(n43600), .Z(n43595) );
  AND U52864 ( .A(n43601), .B(n43602), .Z(n43489) );
  XOR U52865 ( .A(n43569), .B(n43568), .Z(N61515) );
  XNOR U52866 ( .A(n43586), .B(n43587), .Z(n43568) );
  XNOR U52867 ( .A(n43601), .B(n43602), .Z(n43587) );
  XOR U52868 ( .A(n43598), .B(n43597), .Z(n43602) );
  XOR U52869 ( .A(y[1716]), .B(x[1716]), .Z(n43597) );
  XOR U52870 ( .A(n43600), .B(n43599), .Z(n43598) );
  XOR U52871 ( .A(y[1718]), .B(x[1718]), .Z(n43599) );
  XOR U52872 ( .A(y[1717]), .B(x[1717]), .Z(n43600) );
  XOR U52873 ( .A(n43592), .B(n43591), .Z(n43601) );
  XOR U52874 ( .A(n43594), .B(n43593), .Z(n43591) );
  XOR U52875 ( .A(y[1715]), .B(x[1715]), .Z(n43593) );
  XOR U52876 ( .A(y[1714]), .B(x[1714]), .Z(n43594) );
  XOR U52877 ( .A(y[1713]), .B(x[1713]), .Z(n43592) );
  XNOR U52878 ( .A(n43585), .B(n43584), .Z(n43586) );
  XNOR U52879 ( .A(n43581), .B(n43580), .Z(n43584) );
  XOR U52880 ( .A(n43583), .B(n43582), .Z(n43580) );
  XOR U52881 ( .A(y[1712]), .B(x[1712]), .Z(n43582) );
  XOR U52882 ( .A(y[1711]), .B(x[1711]), .Z(n43583) );
  XOR U52883 ( .A(y[1710]), .B(x[1710]), .Z(n43581) );
  XOR U52884 ( .A(n43575), .B(n43574), .Z(n43585) );
  XOR U52885 ( .A(n43577), .B(n43576), .Z(n43574) );
  XOR U52886 ( .A(y[1709]), .B(x[1709]), .Z(n43576) );
  XOR U52887 ( .A(y[1708]), .B(x[1708]), .Z(n43577) );
  XOR U52888 ( .A(y[1707]), .B(x[1707]), .Z(n43575) );
  XNOR U52889 ( .A(n43551), .B(n43552), .Z(n43569) );
  XNOR U52890 ( .A(n43566), .B(n43567), .Z(n43552) );
  XOR U52891 ( .A(n43563), .B(n43562), .Z(n43567) );
  XOR U52892 ( .A(y[1704]), .B(x[1704]), .Z(n43562) );
  XOR U52893 ( .A(n43565), .B(n43564), .Z(n43563) );
  XOR U52894 ( .A(y[1706]), .B(x[1706]), .Z(n43564) );
  XOR U52895 ( .A(y[1705]), .B(x[1705]), .Z(n43565) );
  XOR U52896 ( .A(n43557), .B(n43556), .Z(n43566) );
  XOR U52897 ( .A(n43559), .B(n43558), .Z(n43556) );
  XOR U52898 ( .A(y[1703]), .B(x[1703]), .Z(n43558) );
  XOR U52899 ( .A(y[1702]), .B(x[1702]), .Z(n43559) );
  XOR U52900 ( .A(y[1701]), .B(x[1701]), .Z(n43557) );
  XNOR U52901 ( .A(n43550), .B(n43549), .Z(n43551) );
  XNOR U52902 ( .A(n43546), .B(n43545), .Z(n43549) );
  XOR U52903 ( .A(n43548), .B(n43547), .Z(n43545) );
  XOR U52904 ( .A(y[1700]), .B(x[1700]), .Z(n43547) );
  XOR U52905 ( .A(y[1699]), .B(x[1699]), .Z(n43548) );
  XOR U52906 ( .A(y[1698]), .B(x[1698]), .Z(n43546) );
  XOR U52907 ( .A(n43540), .B(n43539), .Z(n43550) );
  XOR U52908 ( .A(n43542), .B(n43541), .Z(n43539) );
  XOR U52909 ( .A(y[1697]), .B(x[1697]), .Z(n43541) );
  XOR U52910 ( .A(y[1696]), .B(x[1696]), .Z(n43542) );
  XOR U52911 ( .A(y[1695]), .B(x[1695]), .Z(n43540) );
  NAND U52912 ( .A(n43603), .B(n43604), .Z(N61506) );
  NAND U52913 ( .A(n43605), .B(n43606), .Z(n43604) );
  NANDN U52914 ( .A(n43607), .B(n43608), .Z(n43606) );
  NANDN U52915 ( .A(n43608), .B(n43607), .Z(n43603) );
  XOR U52916 ( .A(n43607), .B(n43609), .Z(N61505) );
  XNOR U52917 ( .A(n43605), .B(n43608), .Z(n43609) );
  NAND U52918 ( .A(n43610), .B(n43611), .Z(n43608) );
  NAND U52919 ( .A(n43612), .B(n43613), .Z(n43611) );
  NANDN U52920 ( .A(n43614), .B(n43615), .Z(n43613) );
  NANDN U52921 ( .A(n43615), .B(n43614), .Z(n43610) );
  AND U52922 ( .A(n43616), .B(n43617), .Z(n43605) );
  NAND U52923 ( .A(n43618), .B(n43619), .Z(n43617) );
  NANDN U52924 ( .A(n43620), .B(n43621), .Z(n43619) );
  NANDN U52925 ( .A(n43621), .B(n43620), .Z(n43616) );
  IV U52926 ( .A(n43622), .Z(n43621) );
  AND U52927 ( .A(n43623), .B(n43624), .Z(n43607) );
  NAND U52928 ( .A(n43625), .B(n43626), .Z(n43624) );
  NANDN U52929 ( .A(n43627), .B(n43628), .Z(n43626) );
  NANDN U52930 ( .A(n43628), .B(n43627), .Z(n43623) );
  XOR U52931 ( .A(n43620), .B(n43629), .Z(N61504) );
  XNOR U52932 ( .A(n43618), .B(n43622), .Z(n43629) );
  XOR U52933 ( .A(n43615), .B(n43630), .Z(n43622) );
  XNOR U52934 ( .A(n43612), .B(n43614), .Z(n43630) );
  AND U52935 ( .A(n43631), .B(n43632), .Z(n43614) );
  NANDN U52936 ( .A(n43633), .B(n43634), .Z(n43632) );
  OR U52937 ( .A(n43635), .B(n43636), .Z(n43634) );
  IV U52938 ( .A(n43637), .Z(n43636) );
  NANDN U52939 ( .A(n43637), .B(n43635), .Z(n43631) );
  AND U52940 ( .A(n43638), .B(n43639), .Z(n43612) );
  NAND U52941 ( .A(n43640), .B(n43641), .Z(n43639) );
  NANDN U52942 ( .A(n43642), .B(n43643), .Z(n43641) );
  NANDN U52943 ( .A(n43643), .B(n43642), .Z(n43638) );
  IV U52944 ( .A(n43644), .Z(n43643) );
  NAND U52945 ( .A(n43645), .B(n43646), .Z(n43615) );
  NANDN U52946 ( .A(n43647), .B(n43648), .Z(n43646) );
  NANDN U52947 ( .A(n43649), .B(n43650), .Z(n43648) );
  NANDN U52948 ( .A(n43650), .B(n43649), .Z(n43645) );
  IV U52949 ( .A(n43651), .Z(n43649) );
  AND U52950 ( .A(n43652), .B(n43653), .Z(n43618) );
  NAND U52951 ( .A(n43654), .B(n43655), .Z(n43653) );
  NANDN U52952 ( .A(n43656), .B(n43657), .Z(n43655) );
  NANDN U52953 ( .A(n43657), .B(n43656), .Z(n43652) );
  XOR U52954 ( .A(n43628), .B(n43658), .Z(n43620) );
  XNOR U52955 ( .A(n43625), .B(n43627), .Z(n43658) );
  AND U52956 ( .A(n43659), .B(n43660), .Z(n43627) );
  NANDN U52957 ( .A(n43661), .B(n43662), .Z(n43660) );
  OR U52958 ( .A(n43663), .B(n43664), .Z(n43662) );
  IV U52959 ( .A(n43665), .Z(n43664) );
  NANDN U52960 ( .A(n43665), .B(n43663), .Z(n43659) );
  AND U52961 ( .A(n43666), .B(n43667), .Z(n43625) );
  NAND U52962 ( .A(n43668), .B(n43669), .Z(n43667) );
  NANDN U52963 ( .A(n43670), .B(n43671), .Z(n43669) );
  NANDN U52964 ( .A(n43671), .B(n43670), .Z(n43666) );
  IV U52965 ( .A(n43672), .Z(n43671) );
  NAND U52966 ( .A(n43673), .B(n43674), .Z(n43628) );
  NANDN U52967 ( .A(n43675), .B(n43676), .Z(n43674) );
  NANDN U52968 ( .A(n43677), .B(n43678), .Z(n43676) );
  NANDN U52969 ( .A(n43678), .B(n43677), .Z(n43673) );
  IV U52970 ( .A(n43679), .Z(n43677) );
  XOR U52971 ( .A(n43654), .B(n43680), .Z(N61503) );
  XNOR U52972 ( .A(n43657), .B(n43656), .Z(n43680) );
  XNOR U52973 ( .A(n43668), .B(n43681), .Z(n43656) );
  XNOR U52974 ( .A(n43672), .B(n43670), .Z(n43681) );
  XOR U52975 ( .A(n43678), .B(n43682), .Z(n43670) );
  XNOR U52976 ( .A(n43675), .B(n43679), .Z(n43682) );
  AND U52977 ( .A(n43683), .B(n43684), .Z(n43679) );
  NAND U52978 ( .A(n43685), .B(n43686), .Z(n43684) );
  NAND U52979 ( .A(n43687), .B(n43688), .Z(n43683) );
  AND U52980 ( .A(n43689), .B(n43690), .Z(n43675) );
  NAND U52981 ( .A(n43691), .B(n43692), .Z(n43690) );
  NAND U52982 ( .A(n43693), .B(n43694), .Z(n43689) );
  NANDN U52983 ( .A(n43695), .B(n43696), .Z(n43678) );
  ANDN U52984 ( .B(n43697), .A(n43698), .Z(n43672) );
  XNOR U52985 ( .A(n43663), .B(n43699), .Z(n43668) );
  XNOR U52986 ( .A(n43661), .B(n43665), .Z(n43699) );
  AND U52987 ( .A(n43700), .B(n43701), .Z(n43665) );
  NAND U52988 ( .A(n43702), .B(n43703), .Z(n43701) );
  NAND U52989 ( .A(n43704), .B(n43705), .Z(n43700) );
  AND U52990 ( .A(n43706), .B(n43707), .Z(n43661) );
  NAND U52991 ( .A(n43708), .B(n43709), .Z(n43707) );
  NAND U52992 ( .A(n43710), .B(n43711), .Z(n43706) );
  AND U52993 ( .A(n43712), .B(n43713), .Z(n43663) );
  NAND U52994 ( .A(n43714), .B(n43715), .Z(n43657) );
  XNOR U52995 ( .A(n43640), .B(n43716), .Z(n43654) );
  XNOR U52996 ( .A(n43644), .B(n43642), .Z(n43716) );
  XOR U52997 ( .A(n43650), .B(n43717), .Z(n43642) );
  XNOR U52998 ( .A(n43647), .B(n43651), .Z(n43717) );
  AND U52999 ( .A(n43718), .B(n43719), .Z(n43651) );
  NAND U53000 ( .A(n43720), .B(n43721), .Z(n43719) );
  NAND U53001 ( .A(n43722), .B(n43723), .Z(n43718) );
  AND U53002 ( .A(n43724), .B(n43725), .Z(n43647) );
  NAND U53003 ( .A(n43726), .B(n43727), .Z(n43725) );
  NAND U53004 ( .A(n43728), .B(n43729), .Z(n43724) );
  NANDN U53005 ( .A(n43730), .B(n43731), .Z(n43650) );
  ANDN U53006 ( .B(n43732), .A(n43733), .Z(n43644) );
  XNOR U53007 ( .A(n43635), .B(n43734), .Z(n43640) );
  XNOR U53008 ( .A(n43633), .B(n43637), .Z(n43734) );
  AND U53009 ( .A(n43735), .B(n43736), .Z(n43637) );
  NAND U53010 ( .A(n43737), .B(n43738), .Z(n43736) );
  NAND U53011 ( .A(n43739), .B(n43740), .Z(n43735) );
  AND U53012 ( .A(n43741), .B(n43742), .Z(n43633) );
  NAND U53013 ( .A(n43743), .B(n43744), .Z(n43742) );
  NAND U53014 ( .A(n43745), .B(n43746), .Z(n43741) );
  AND U53015 ( .A(n43747), .B(n43748), .Z(n43635) );
  XOR U53016 ( .A(n43715), .B(n43714), .Z(N61502) );
  XNOR U53017 ( .A(n43732), .B(n43733), .Z(n43714) );
  XNOR U53018 ( .A(n43747), .B(n43748), .Z(n43733) );
  XOR U53019 ( .A(n43744), .B(n43743), .Z(n43748) );
  XOR U53020 ( .A(y[1692]), .B(x[1692]), .Z(n43743) );
  XOR U53021 ( .A(n43746), .B(n43745), .Z(n43744) );
  XOR U53022 ( .A(y[1694]), .B(x[1694]), .Z(n43745) );
  XOR U53023 ( .A(y[1693]), .B(x[1693]), .Z(n43746) );
  XOR U53024 ( .A(n43738), .B(n43737), .Z(n43747) );
  XOR U53025 ( .A(n43740), .B(n43739), .Z(n43737) );
  XOR U53026 ( .A(y[1691]), .B(x[1691]), .Z(n43739) );
  XOR U53027 ( .A(y[1690]), .B(x[1690]), .Z(n43740) );
  XOR U53028 ( .A(y[1689]), .B(x[1689]), .Z(n43738) );
  XNOR U53029 ( .A(n43731), .B(n43730), .Z(n43732) );
  XNOR U53030 ( .A(n43727), .B(n43726), .Z(n43730) );
  XOR U53031 ( .A(n43729), .B(n43728), .Z(n43726) );
  XOR U53032 ( .A(y[1688]), .B(x[1688]), .Z(n43728) );
  XOR U53033 ( .A(y[1687]), .B(x[1687]), .Z(n43729) );
  XOR U53034 ( .A(y[1686]), .B(x[1686]), .Z(n43727) );
  XOR U53035 ( .A(n43721), .B(n43720), .Z(n43731) );
  XOR U53036 ( .A(n43723), .B(n43722), .Z(n43720) );
  XOR U53037 ( .A(y[1685]), .B(x[1685]), .Z(n43722) );
  XOR U53038 ( .A(y[1684]), .B(x[1684]), .Z(n43723) );
  XOR U53039 ( .A(y[1683]), .B(x[1683]), .Z(n43721) );
  XNOR U53040 ( .A(n43697), .B(n43698), .Z(n43715) );
  XNOR U53041 ( .A(n43712), .B(n43713), .Z(n43698) );
  XOR U53042 ( .A(n43709), .B(n43708), .Z(n43713) );
  XOR U53043 ( .A(y[1680]), .B(x[1680]), .Z(n43708) );
  XOR U53044 ( .A(n43711), .B(n43710), .Z(n43709) );
  XOR U53045 ( .A(y[1682]), .B(x[1682]), .Z(n43710) );
  XOR U53046 ( .A(y[1681]), .B(x[1681]), .Z(n43711) );
  XOR U53047 ( .A(n43703), .B(n43702), .Z(n43712) );
  XOR U53048 ( .A(n43705), .B(n43704), .Z(n43702) );
  XOR U53049 ( .A(y[1679]), .B(x[1679]), .Z(n43704) );
  XOR U53050 ( .A(y[1678]), .B(x[1678]), .Z(n43705) );
  XOR U53051 ( .A(y[1677]), .B(x[1677]), .Z(n43703) );
  XNOR U53052 ( .A(n43696), .B(n43695), .Z(n43697) );
  XNOR U53053 ( .A(n43692), .B(n43691), .Z(n43695) );
  XOR U53054 ( .A(n43694), .B(n43693), .Z(n43691) );
  XOR U53055 ( .A(y[1676]), .B(x[1676]), .Z(n43693) );
  XOR U53056 ( .A(y[1675]), .B(x[1675]), .Z(n43694) );
  XOR U53057 ( .A(y[1674]), .B(x[1674]), .Z(n43692) );
  XOR U53058 ( .A(n43686), .B(n43685), .Z(n43696) );
  XOR U53059 ( .A(n43688), .B(n43687), .Z(n43685) );
  XOR U53060 ( .A(y[1673]), .B(x[1673]), .Z(n43687) );
  XOR U53061 ( .A(y[1672]), .B(x[1672]), .Z(n43688) );
  XOR U53062 ( .A(y[1671]), .B(x[1671]), .Z(n43686) );
  NAND U53063 ( .A(n43749), .B(n43750), .Z(N61493) );
  NAND U53064 ( .A(n43751), .B(n43752), .Z(n43750) );
  NANDN U53065 ( .A(n43753), .B(n43754), .Z(n43752) );
  NANDN U53066 ( .A(n43754), .B(n43753), .Z(n43749) );
  XOR U53067 ( .A(n43753), .B(n43755), .Z(N61492) );
  XNOR U53068 ( .A(n43751), .B(n43754), .Z(n43755) );
  NAND U53069 ( .A(n43756), .B(n43757), .Z(n43754) );
  NAND U53070 ( .A(n43758), .B(n43759), .Z(n43757) );
  NANDN U53071 ( .A(n43760), .B(n43761), .Z(n43759) );
  NANDN U53072 ( .A(n43761), .B(n43760), .Z(n43756) );
  AND U53073 ( .A(n43762), .B(n43763), .Z(n43751) );
  NAND U53074 ( .A(n43764), .B(n43765), .Z(n43763) );
  NANDN U53075 ( .A(n43766), .B(n43767), .Z(n43765) );
  NANDN U53076 ( .A(n43767), .B(n43766), .Z(n43762) );
  IV U53077 ( .A(n43768), .Z(n43767) );
  AND U53078 ( .A(n43769), .B(n43770), .Z(n43753) );
  NAND U53079 ( .A(n43771), .B(n43772), .Z(n43770) );
  NANDN U53080 ( .A(n43773), .B(n43774), .Z(n43772) );
  NANDN U53081 ( .A(n43774), .B(n43773), .Z(n43769) );
  XOR U53082 ( .A(n43766), .B(n43775), .Z(N61491) );
  XNOR U53083 ( .A(n43764), .B(n43768), .Z(n43775) );
  XOR U53084 ( .A(n43761), .B(n43776), .Z(n43768) );
  XNOR U53085 ( .A(n43758), .B(n43760), .Z(n43776) );
  AND U53086 ( .A(n43777), .B(n43778), .Z(n43760) );
  NANDN U53087 ( .A(n43779), .B(n43780), .Z(n43778) );
  OR U53088 ( .A(n43781), .B(n43782), .Z(n43780) );
  IV U53089 ( .A(n43783), .Z(n43782) );
  NANDN U53090 ( .A(n43783), .B(n43781), .Z(n43777) );
  AND U53091 ( .A(n43784), .B(n43785), .Z(n43758) );
  NAND U53092 ( .A(n43786), .B(n43787), .Z(n43785) );
  NANDN U53093 ( .A(n43788), .B(n43789), .Z(n43787) );
  NANDN U53094 ( .A(n43789), .B(n43788), .Z(n43784) );
  IV U53095 ( .A(n43790), .Z(n43789) );
  NAND U53096 ( .A(n43791), .B(n43792), .Z(n43761) );
  NANDN U53097 ( .A(n43793), .B(n43794), .Z(n43792) );
  NANDN U53098 ( .A(n43795), .B(n43796), .Z(n43794) );
  NANDN U53099 ( .A(n43796), .B(n43795), .Z(n43791) );
  IV U53100 ( .A(n43797), .Z(n43795) );
  AND U53101 ( .A(n43798), .B(n43799), .Z(n43764) );
  NAND U53102 ( .A(n43800), .B(n43801), .Z(n43799) );
  NANDN U53103 ( .A(n43802), .B(n43803), .Z(n43801) );
  NANDN U53104 ( .A(n43803), .B(n43802), .Z(n43798) );
  XOR U53105 ( .A(n43774), .B(n43804), .Z(n43766) );
  XNOR U53106 ( .A(n43771), .B(n43773), .Z(n43804) );
  AND U53107 ( .A(n43805), .B(n43806), .Z(n43773) );
  NANDN U53108 ( .A(n43807), .B(n43808), .Z(n43806) );
  OR U53109 ( .A(n43809), .B(n43810), .Z(n43808) );
  IV U53110 ( .A(n43811), .Z(n43810) );
  NANDN U53111 ( .A(n43811), .B(n43809), .Z(n43805) );
  AND U53112 ( .A(n43812), .B(n43813), .Z(n43771) );
  NAND U53113 ( .A(n43814), .B(n43815), .Z(n43813) );
  NANDN U53114 ( .A(n43816), .B(n43817), .Z(n43815) );
  NANDN U53115 ( .A(n43817), .B(n43816), .Z(n43812) );
  IV U53116 ( .A(n43818), .Z(n43817) );
  NAND U53117 ( .A(n43819), .B(n43820), .Z(n43774) );
  NANDN U53118 ( .A(n43821), .B(n43822), .Z(n43820) );
  NANDN U53119 ( .A(n43823), .B(n43824), .Z(n43822) );
  NANDN U53120 ( .A(n43824), .B(n43823), .Z(n43819) );
  IV U53121 ( .A(n43825), .Z(n43823) );
  XOR U53122 ( .A(n43800), .B(n43826), .Z(N61490) );
  XNOR U53123 ( .A(n43803), .B(n43802), .Z(n43826) );
  XNOR U53124 ( .A(n43814), .B(n43827), .Z(n43802) );
  XNOR U53125 ( .A(n43818), .B(n43816), .Z(n43827) );
  XOR U53126 ( .A(n43824), .B(n43828), .Z(n43816) );
  XNOR U53127 ( .A(n43821), .B(n43825), .Z(n43828) );
  AND U53128 ( .A(n43829), .B(n43830), .Z(n43825) );
  NAND U53129 ( .A(n43831), .B(n43832), .Z(n43830) );
  NAND U53130 ( .A(n43833), .B(n43834), .Z(n43829) );
  AND U53131 ( .A(n43835), .B(n43836), .Z(n43821) );
  NAND U53132 ( .A(n43837), .B(n43838), .Z(n43836) );
  NAND U53133 ( .A(n43839), .B(n43840), .Z(n43835) );
  NANDN U53134 ( .A(n43841), .B(n43842), .Z(n43824) );
  ANDN U53135 ( .B(n43843), .A(n43844), .Z(n43818) );
  XNOR U53136 ( .A(n43809), .B(n43845), .Z(n43814) );
  XNOR U53137 ( .A(n43807), .B(n43811), .Z(n43845) );
  AND U53138 ( .A(n43846), .B(n43847), .Z(n43811) );
  NAND U53139 ( .A(n43848), .B(n43849), .Z(n43847) );
  NAND U53140 ( .A(n43850), .B(n43851), .Z(n43846) );
  AND U53141 ( .A(n43852), .B(n43853), .Z(n43807) );
  NAND U53142 ( .A(n43854), .B(n43855), .Z(n43853) );
  NAND U53143 ( .A(n43856), .B(n43857), .Z(n43852) );
  AND U53144 ( .A(n43858), .B(n43859), .Z(n43809) );
  NAND U53145 ( .A(n43860), .B(n43861), .Z(n43803) );
  XNOR U53146 ( .A(n43786), .B(n43862), .Z(n43800) );
  XNOR U53147 ( .A(n43790), .B(n43788), .Z(n43862) );
  XOR U53148 ( .A(n43796), .B(n43863), .Z(n43788) );
  XNOR U53149 ( .A(n43793), .B(n43797), .Z(n43863) );
  AND U53150 ( .A(n43864), .B(n43865), .Z(n43797) );
  NAND U53151 ( .A(n43866), .B(n43867), .Z(n43865) );
  NAND U53152 ( .A(n43868), .B(n43869), .Z(n43864) );
  AND U53153 ( .A(n43870), .B(n43871), .Z(n43793) );
  NAND U53154 ( .A(n43872), .B(n43873), .Z(n43871) );
  NAND U53155 ( .A(n43874), .B(n43875), .Z(n43870) );
  NANDN U53156 ( .A(n43876), .B(n43877), .Z(n43796) );
  ANDN U53157 ( .B(n43878), .A(n43879), .Z(n43790) );
  XNOR U53158 ( .A(n43781), .B(n43880), .Z(n43786) );
  XNOR U53159 ( .A(n43779), .B(n43783), .Z(n43880) );
  AND U53160 ( .A(n43881), .B(n43882), .Z(n43783) );
  NAND U53161 ( .A(n43883), .B(n43884), .Z(n43882) );
  NAND U53162 ( .A(n43885), .B(n43886), .Z(n43881) );
  AND U53163 ( .A(n43887), .B(n43888), .Z(n43779) );
  NAND U53164 ( .A(n43889), .B(n43890), .Z(n43888) );
  NAND U53165 ( .A(n43891), .B(n43892), .Z(n43887) );
  AND U53166 ( .A(n43893), .B(n43894), .Z(n43781) );
  XOR U53167 ( .A(n43861), .B(n43860), .Z(N61489) );
  XNOR U53168 ( .A(n43878), .B(n43879), .Z(n43860) );
  XNOR U53169 ( .A(n43893), .B(n43894), .Z(n43879) );
  XOR U53170 ( .A(n43890), .B(n43889), .Z(n43894) );
  XOR U53171 ( .A(y[1668]), .B(x[1668]), .Z(n43889) );
  XOR U53172 ( .A(n43892), .B(n43891), .Z(n43890) );
  XOR U53173 ( .A(y[1670]), .B(x[1670]), .Z(n43891) );
  XOR U53174 ( .A(y[1669]), .B(x[1669]), .Z(n43892) );
  XOR U53175 ( .A(n43884), .B(n43883), .Z(n43893) );
  XOR U53176 ( .A(n43886), .B(n43885), .Z(n43883) );
  XOR U53177 ( .A(y[1667]), .B(x[1667]), .Z(n43885) );
  XOR U53178 ( .A(y[1666]), .B(x[1666]), .Z(n43886) );
  XOR U53179 ( .A(y[1665]), .B(x[1665]), .Z(n43884) );
  XNOR U53180 ( .A(n43877), .B(n43876), .Z(n43878) );
  XNOR U53181 ( .A(n43873), .B(n43872), .Z(n43876) );
  XOR U53182 ( .A(n43875), .B(n43874), .Z(n43872) );
  XOR U53183 ( .A(y[1664]), .B(x[1664]), .Z(n43874) );
  XOR U53184 ( .A(y[1663]), .B(x[1663]), .Z(n43875) );
  XOR U53185 ( .A(y[1662]), .B(x[1662]), .Z(n43873) );
  XOR U53186 ( .A(n43867), .B(n43866), .Z(n43877) );
  XOR U53187 ( .A(n43869), .B(n43868), .Z(n43866) );
  XOR U53188 ( .A(y[1661]), .B(x[1661]), .Z(n43868) );
  XOR U53189 ( .A(y[1660]), .B(x[1660]), .Z(n43869) );
  XOR U53190 ( .A(y[1659]), .B(x[1659]), .Z(n43867) );
  XNOR U53191 ( .A(n43843), .B(n43844), .Z(n43861) );
  XNOR U53192 ( .A(n43858), .B(n43859), .Z(n43844) );
  XOR U53193 ( .A(n43855), .B(n43854), .Z(n43859) );
  XOR U53194 ( .A(y[1656]), .B(x[1656]), .Z(n43854) );
  XOR U53195 ( .A(n43857), .B(n43856), .Z(n43855) );
  XOR U53196 ( .A(y[1658]), .B(x[1658]), .Z(n43856) );
  XOR U53197 ( .A(y[1657]), .B(x[1657]), .Z(n43857) );
  XOR U53198 ( .A(n43849), .B(n43848), .Z(n43858) );
  XOR U53199 ( .A(n43851), .B(n43850), .Z(n43848) );
  XOR U53200 ( .A(y[1655]), .B(x[1655]), .Z(n43850) );
  XOR U53201 ( .A(y[1654]), .B(x[1654]), .Z(n43851) );
  XOR U53202 ( .A(y[1653]), .B(x[1653]), .Z(n43849) );
  XNOR U53203 ( .A(n43842), .B(n43841), .Z(n43843) );
  XNOR U53204 ( .A(n43838), .B(n43837), .Z(n43841) );
  XOR U53205 ( .A(n43840), .B(n43839), .Z(n43837) );
  XOR U53206 ( .A(y[1652]), .B(x[1652]), .Z(n43839) );
  XOR U53207 ( .A(y[1651]), .B(x[1651]), .Z(n43840) );
  XOR U53208 ( .A(y[1650]), .B(x[1650]), .Z(n43838) );
  XOR U53209 ( .A(n43832), .B(n43831), .Z(n43842) );
  XOR U53210 ( .A(n43834), .B(n43833), .Z(n43831) );
  XOR U53211 ( .A(y[1649]), .B(x[1649]), .Z(n43833) );
  XOR U53212 ( .A(y[1648]), .B(x[1648]), .Z(n43834) );
  XOR U53213 ( .A(y[1647]), .B(x[1647]), .Z(n43832) );
  NAND U53214 ( .A(n43895), .B(n43896), .Z(N61480) );
  NAND U53215 ( .A(n43897), .B(n43898), .Z(n43896) );
  NANDN U53216 ( .A(n43899), .B(n43900), .Z(n43898) );
  NANDN U53217 ( .A(n43900), .B(n43899), .Z(n43895) );
  XOR U53218 ( .A(n43899), .B(n43901), .Z(N61479) );
  XNOR U53219 ( .A(n43897), .B(n43900), .Z(n43901) );
  NAND U53220 ( .A(n43902), .B(n43903), .Z(n43900) );
  NAND U53221 ( .A(n43904), .B(n43905), .Z(n43903) );
  NANDN U53222 ( .A(n43906), .B(n43907), .Z(n43905) );
  NANDN U53223 ( .A(n43907), .B(n43906), .Z(n43902) );
  AND U53224 ( .A(n43908), .B(n43909), .Z(n43897) );
  NAND U53225 ( .A(n43910), .B(n43911), .Z(n43909) );
  NANDN U53226 ( .A(n43912), .B(n43913), .Z(n43911) );
  NANDN U53227 ( .A(n43913), .B(n43912), .Z(n43908) );
  IV U53228 ( .A(n43914), .Z(n43913) );
  AND U53229 ( .A(n43915), .B(n43916), .Z(n43899) );
  NAND U53230 ( .A(n43917), .B(n43918), .Z(n43916) );
  NANDN U53231 ( .A(n43919), .B(n43920), .Z(n43918) );
  NANDN U53232 ( .A(n43920), .B(n43919), .Z(n43915) );
  XOR U53233 ( .A(n43912), .B(n43921), .Z(N61478) );
  XNOR U53234 ( .A(n43910), .B(n43914), .Z(n43921) );
  XOR U53235 ( .A(n43907), .B(n43922), .Z(n43914) );
  XNOR U53236 ( .A(n43904), .B(n43906), .Z(n43922) );
  AND U53237 ( .A(n43923), .B(n43924), .Z(n43906) );
  NANDN U53238 ( .A(n43925), .B(n43926), .Z(n43924) );
  OR U53239 ( .A(n43927), .B(n43928), .Z(n43926) );
  IV U53240 ( .A(n43929), .Z(n43928) );
  NANDN U53241 ( .A(n43929), .B(n43927), .Z(n43923) );
  AND U53242 ( .A(n43930), .B(n43931), .Z(n43904) );
  NAND U53243 ( .A(n43932), .B(n43933), .Z(n43931) );
  NANDN U53244 ( .A(n43934), .B(n43935), .Z(n43933) );
  NANDN U53245 ( .A(n43935), .B(n43934), .Z(n43930) );
  IV U53246 ( .A(n43936), .Z(n43935) );
  NAND U53247 ( .A(n43937), .B(n43938), .Z(n43907) );
  NANDN U53248 ( .A(n43939), .B(n43940), .Z(n43938) );
  NANDN U53249 ( .A(n43941), .B(n43942), .Z(n43940) );
  NANDN U53250 ( .A(n43942), .B(n43941), .Z(n43937) );
  IV U53251 ( .A(n43943), .Z(n43941) );
  AND U53252 ( .A(n43944), .B(n43945), .Z(n43910) );
  NAND U53253 ( .A(n43946), .B(n43947), .Z(n43945) );
  NANDN U53254 ( .A(n43948), .B(n43949), .Z(n43947) );
  NANDN U53255 ( .A(n43949), .B(n43948), .Z(n43944) );
  XOR U53256 ( .A(n43920), .B(n43950), .Z(n43912) );
  XNOR U53257 ( .A(n43917), .B(n43919), .Z(n43950) );
  AND U53258 ( .A(n43951), .B(n43952), .Z(n43919) );
  NANDN U53259 ( .A(n43953), .B(n43954), .Z(n43952) );
  OR U53260 ( .A(n43955), .B(n43956), .Z(n43954) );
  IV U53261 ( .A(n43957), .Z(n43956) );
  NANDN U53262 ( .A(n43957), .B(n43955), .Z(n43951) );
  AND U53263 ( .A(n43958), .B(n43959), .Z(n43917) );
  NAND U53264 ( .A(n43960), .B(n43961), .Z(n43959) );
  NANDN U53265 ( .A(n43962), .B(n43963), .Z(n43961) );
  NANDN U53266 ( .A(n43963), .B(n43962), .Z(n43958) );
  IV U53267 ( .A(n43964), .Z(n43963) );
  NAND U53268 ( .A(n43965), .B(n43966), .Z(n43920) );
  NANDN U53269 ( .A(n43967), .B(n43968), .Z(n43966) );
  NANDN U53270 ( .A(n43969), .B(n43970), .Z(n43968) );
  NANDN U53271 ( .A(n43970), .B(n43969), .Z(n43965) );
  IV U53272 ( .A(n43971), .Z(n43969) );
  XOR U53273 ( .A(n43946), .B(n43972), .Z(N61477) );
  XNOR U53274 ( .A(n43949), .B(n43948), .Z(n43972) );
  XNOR U53275 ( .A(n43960), .B(n43973), .Z(n43948) );
  XNOR U53276 ( .A(n43964), .B(n43962), .Z(n43973) );
  XOR U53277 ( .A(n43970), .B(n43974), .Z(n43962) );
  XNOR U53278 ( .A(n43967), .B(n43971), .Z(n43974) );
  AND U53279 ( .A(n43975), .B(n43976), .Z(n43971) );
  NAND U53280 ( .A(n43977), .B(n43978), .Z(n43976) );
  NAND U53281 ( .A(n43979), .B(n43980), .Z(n43975) );
  AND U53282 ( .A(n43981), .B(n43982), .Z(n43967) );
  NAND U53283 ( .A(n43983), .B(n43984), .Z(n43982) );
  NAND U53284 ( .A(n43985), .B(n43986), .Z(n43981) );
  NANDN U53285 ( .A(n43987), .B(n43988), .Z(n43970) );
  ANDN U53286 ( .B(n43989), .A(n43990), .Z(n43964) );
  XNOR U53287 ( .A(n43955), .B(n43991), .Z(n43960) );
  XNOR U53288 ( .A(n43953), .B(n43957), .Z(n43991) );
  AND U53289 ( .A(n43992), .B(n43993), .Z(n43957) );
  NAND U53290 ( .A(n43994), .B(n43995), .Z(n43993) );
  NAND U53291 ( .A(n43996), .B(n43997), .Z(n43992) );
  AND U53292 ( .A(n43998), .B(n43999), .Z(n43953) );
  NAND U53293 ( .A(n44000), .B(n44001), .Z(n43999) );
  NAND U53294 ( .A(n44002), .B(n44003), .Z(n43998) );
  AND U53295 ( .A(n44004), .B(n44005), .Z(n43955) );
  NAND U53296 ( .A(n44006), .B(n44007), .Z(n43949) );
  XNOR U53297 ( .A(n43932), .B(n44008), .Z(n43946) );
  XNOR U53298 ( .A(n43936), .B(n43934), .Z(n44008) );
  XOR U53299 ( .A(n43942), .B(n44009), .Z(n43934) );
  XNOR U53300 ( .A(n43939), .B(n43943), .Z(n44009) );
  AND U53301 ( .A(n44010), .B(n44011), .Z(n43943) );
  NAND U53302 ( .A(n44012), .B(n44013), .Z(n44011) );
  NAND U53303 ( .A(n44014), .B(n44015), .Z(n44010) );
  AND U53304 ( .A(n44016), .B(n44017), .Z(n43939) );
  NAND U53305 ( .A(n44018), .B(n44019), .Z(n44017) );
  NAND U53306 ( .A(n44020), .B(n44021), .Z(n44016) );
  NANDN U53307 ( .A(n44022), .B(n44023), .Z(n43942) );
  ANDN U53308 ( .B(n44024), .A(n44025), .Z(n43936) );
  XNOR U53309 ( .A(n43927), .B(n44026), .Z(n43932) );
  XNOR U53310 ( .A(n43925), .B(n43929), .Z(n44026) );
  AND U53311 ( .A(n44027), .B(n44028), .Z(n43929) );
  NAND U53312 ( .A(n44029), .B(n44030), .Z(n44028) );
  NAND U53313 ( .A(n44031), .B(n44032), .Z(n44027) );
  AND U53314 ( .A(n44033), .B(n44034), .Z(n43925) );
  NAND U53315 ( .A(n44035), .B(n44036), .Z(n44034) );
  NAND U53316 ( .A(n44037), .B(n44038), .Z(n44033) );
  AND U53317 ( .A(n44039), .B(n44040), .Z(n43927) );
  XOR U53318 ( .A(n44007), .B(n44006), .Z(N61476) );
  XNOR U53319 ( .A(n44024), .B(n44025), .Z(n44006) );
  XNOR U53320 ( .A(n44039), .B(n44040), .Z(n44025) );
  XOR U53321 ( .A(n44036), .B(n44035), .Z(n44040) );
  XOR U53322 ( .A(y[1644]), .B(x[1644]), .Z(n44035) );
  XOR U53323 ( .A(n44038), .B(n44037), .Z(n44036) );
  XOR U53324 ( .A(y[1646]), .B(x[1646]), .Z(n44037) );
  XOR U53325 ( .A(y[1645]), .B(x[1645]), .Z(n44038) );
  XOR U53326 ( .A(n44030), .B(n44029), .Z(n44039) );
  XOR U53327 ( .A(n44032), .B(n44031), .Z(n44029) );
  XOR U53328 ( .A(y[1643]), .B(x[1643]), .Z(n44031) );
  XOR U53329 ( .A(y[1642]), .B(x[1642]), .Z(n44032) );
  XOR U53330 ( .A(y[1641]), .B(x[1641]), .Z(n44030) );
  XNOR U53331 ( .A(n44023), .B(n44022), .Z(n44024) );
  XNOR U53332 ( .A(n44019), .B(n44018), .Z(n44022) );
  XOR U53333 ( .A(n44021), .B(n44020), .Z(n44018) );
  XOR U53334 ( .A(y[1640]), .B(x[1640]), .Z(n44020) );
  XOR U53335 ( .A(y[1639]), .B(x[1639]), .Z(n44021) );
  XOR U53336 ( .A(y[1638]), .B(x[1638]), .Z(n44019) );
  XOR U53337 ( .A(n44013), .B(n44012), .Z(n44023) );
  XOR U53338 ( .A(n44015), .B(n44014), .Z(n44012) );
  XOR U53339 ( .A(y[1637]), .B(x[1637]), .Z(n44014) );
  XOR U53340 ( .A(y[1636]), .B(x[1636]), .Z(n44015) );
  XOR U53341 ( .A(y[1635]), .B(x[1635]), .Z(n44013) );
  XNOR U53342 ( .A(n43989), .B(n43990), .Z(n44007) );
  XNOR U53343 ( .A(n44004), .B(n44005), .Z(n43990) );
  XOR U53344 ( .A(n44001), .B(n44000), .Z(n44005) );
  XOR U53345 ( .A(y[1632]), .B(x[1632]), .Z(n44000) );
  XOR U53346 ( .A(n44003), .B(n44002), .Z(n44001) );
  XOR U53347 ( .A(y[1634]), .B(x[1634]), .Z(n44002) );
  XOR U53348 ( .A(y[1633]), .B(x[1633]), .Z(n44003) );
  XOR U53349 ( .A(n43995), .B(n43994), .Z(n44004) );
  XOR U53350 ( .A(n43997), .B(n43996), .Z(n43994) );
  XOR U53351 ( .A(y[1631]), .B(x[1631]), .Z(n43996) );
  XOR U53352 ( .A(y[1630]), .B(x[1630]), .Z(n43997) );
  XOR U53353 ( .A(y[1629]), .B(x[1629]), .Z(n43995) );
  XNOR U53354 ( .A(n43988), .B(n43987), .Z(n43989) );
  XNOR U53355 ( .A(n43984), .B(n43983), .Z(n43987) );
  XOR U53356 ( .A(n43986), .B(n43985), .Z(n43983) );
  XOR U53357 ( .A(y[1628]), .B(x[1628]), .Z(n43985) );
  XOR U53358 ( .A(y[1627]), .B(x[1627]), .Z(n43986) );
  XOR U53359 ( .A(y[1626]), .B(x[1626]), .Z(n43984) );
  XOR U53360 ( .A(n43978), .B(n43977), .Z(n43988) );
  XOR U53361 ( .A(n43980), .B(n43979), .Z(n43977) );
  XOR U53362 ( .A(y[1625]), .B(x[1625]), .Z(n43979) );
  XOR U53363 ( .A(y[1624]), .B(x[1624]), .Z(n43980) );
  XOR U53364 ( .A(y[1623]), .B(x[1623]), .Z(n43978) );
  NAND U53365 ( .A(n44041), .B(n44042), .Z(N61467) );
  NAND U53366 ( .A(n44043), .B(n44044), .Z(n44042) );
  NANDN U53367 ( .A(n44045), .B(n44046), .Z(n44044) );
  NANDN U53368 ( .A(n44046), .B(n44045), .Z(n44041) );
  XOR U53369 ( .A(n44045), .B(n44047), .Z(N61466) );
  XNOR U53370 ( .A(n44043), .B(n44046), .Z(n44047) );
  NAND U53371 ( .A(n44048), .B(n44049), .Z(n44046) );
  NAND U53372 ( .A(n44050), .B(n44051), .Z(n44049) );
  NANDN U53373 ( .A(n44052), .B(n44053), .Z(n44051) );
  NANDN U53374 ( .A(n44053), .B(n44052), .Z(n44048) );
  AND U53375 ( .A(n44054), .B(n44055), .Z(n44043) );
  NAND U53376 ( .A(n44056), .B(n44057), .Z(n44055) );
  NANDN U53377 ( .A(n44058), .B(n44059), .Z(n44057) );
  NANDN U53378 ( .A(n44059), .B(n44058), .Z(n44054) );
  IV U53379 ( .A(n44060), .Z(n44059) );
  AND U53380 ( .A(n44061), .B(n44062), .Z(n44045) );
  NAND U53381 ( .A(n44063), .B(n44064), .Z(n44062) );
  NANDN U53382 ( .A(n44065), .B(n44066), .Z(n44064) );
  NANDN U53383 ( .A(n44066), .B(n44065), .Z(n44061) );
  XOR U53384 ( .A(n44058), .B(n44067), .Z(N61465) );
  XNOR U53385 ( .A(n44056), .B(n44060), .Z(n44067) );
  XOR U53386 ( .A(n44053), .B(n44068), .Z(n44060) );
  XNOR U53387 ( .A(n44050), .B(n44052), .Z(n44068) );
  AND U53388 ( .A(n44069), .B(n44070), .Z(n44052) );
  NANDN U53389 ( .A(n44071), .B(n44072), .Z(n44070) );
  OR U53390 ( .A(n44073), .B(n44074), .Z(n44072) );
  IV U53391 ( .A(n44075), .Z(n44074) );
  NANDN U53392 ( .A(n44075), .B(n44073), .Z(n44069) );
  AND U53393 ( .A(n44076), .B(n44077), .Z(n44050) );
  NAND U53394 ( .A(n44078), .B(n44079), .Z(n44077) );
  NANDN U53395 ( .A(n44080), .B(n44081), .Z(n44079) );
  NANDN U53396 ( .A(n44081), .B(n44080), .Z(n44076) );
  IV U53397 ( .A(n44082), .Z(n44081) );
  NAND U53398 ( .A(n44083), .B(n44084), .Z(n44053) );
  NANDN U53399 ( .A(n44085), .B(n44086), .Z(n44084) );
  NANDN U53400 ( .A(n44087), .B(n44088), .Z(n44086) );
  NANDN U53401 ( .A(n44088), .B(n44087), .Z(n44083) );
  IV U53402 ( .A(n44089), .Z(n44087) );
  AND U53403 ( .A(n44090), .B(n44091), .Z(n44056) );
  NAND U53404 ( .A(n44092), .B(n44093), .Z(n44091) );
  NANDN U53405 ( .A(n44094), .B(n44095), .Z(n44093) );
  NANDN U53406 ( .A(n44095), .B(n44094), .Z(n44090) );
  XOR U53407 ( .A(n44066), .B(n44096), .Z(n44058) );
  XNOR U53408 ( .A(n44063), .B(n44065), .Z(n44096) );
  AND U53409 ( .A(n44097), .B(n44098), .Z(n44065) );
  NANDN U53410 ( .A(n44099), .B(n44100), .Z(n44098) );
  OR U53411 ( .A(n44101), .B(n44102), .Z(n44100) );
  IV U53412 ( .A(n44103), .Z(n44102) );
  NANDN U53413 ( .A(n44103), .B(n44101), .Z(n44097) );
  AND U53414 ( .A(n44104), .B(n44105), .Z(n44063) );
  NAND U53415 ( .A(n44106), .B(n44107), .Z(n44105) );
  NANDN U53416 ( .A(n44108), .B(n44109), .Z(n44107) );
  NANDN U53417 ( .A(n44109), .B(n44108), .Z(n44104) );
  IV U53418 ( .A(n44110), .Z(n44109) );
  NAND U53419 ( .A(n44111), .B(n44112), .Z(n44066) );
  NANDN U53420 ( .A(n44113), .B(n44114), .Z(n44112) );
  NANDN U53421 ( .A(n44115), .B(n44116), .Z(n44114) );
  NANDN U53422 ( .A(n44116), .B(n44115), .Z(n44111) );
  IV U53423 ( .A(n44117), .Z(n44115) );
  XOR U53424 ( .A(n44092), .B(n44118), .Z(N61464) );
  XNOR U53425 ( .A(n44095), .B(n44094), .Z(n44118) );
  XNOR U53426 ( .A(n44106), .B(n44119), .Z(n44094) );
  XNOR U53427 ( .A(n44110), .B(n44108), .Z(n44119) );
  XOR U53428 ( .A(n44116), .B(n44120), .Z(n44108) );
  XNOR U53429 ( .A(n44113), .B(n44117), .Z(n44120) );
  AND U53430 ( .A(n44121), .B(n44122), .Z(n44117) );
  NAND U53431 ( .A(n44123), .B(n44124), .Z(n44122) );
  NAND U53432 ( .A(n44125), .B(n44126), .Z(n44121) );
  AND U53433 ( .A(n44127), .B(n44128), .Z(n44113) );
  NAND U53434 ( .A(n44129), .B(n44130), .Z(n44128) );
  NAND U53435 ( .A(n44131), .B(n44132), .Z(n44127) );
  NANDN U53436 ( .A(n44133), .B(n44134), .Z(n44116) );
  ANDN U53437 ( .B(n44135), .A(n44136), .Z(n44110) );
  XNOR U53438 ( .A(n44101), .B(n44137), .Z(n44106) );
  XNOR U53439 ( .A(n44099), .B(n44103), .Z(n44137) );
  AND U53440 ( .A(n44138), .B(n44139), .Z(n44103) );
  NAND U53441 ( .A(n44140), .B(n44141), .Z(n44139) );
  NAND U53442 ( .A(n44142), .B(n44143), .Z(n44138) );
  AND U53443 ( .A(n44144), .B(n44145), .Z(n44099) );
  NAND U53444 ( .A(n44146), .B(n44147), .Z(n44145) );
  NAND U53445 ( .A(n44148), .B(n44149), .Z(n44144) );
  AND U53446 ( .A(n44150), .B(n44151), .Z(n44101) );
  NAND U53447 ( .A(n44152), .B(n44153), .Z(n44095) );
  XNOR U53448 ( .A(n44078), .B(n44154), .Z(n44092) );
  XNOR U53449 ( .A(n44082), .B(n44080), .Z(n44154) );
  XOR U53450 ( .A(n44088), .B(n44155), .Z(n44080) );
  XNOR U53451 ( .A(n44085), .B(n44089), .Z(n44155) );
  AND U53452 ( .A(n44156), .B(n44157), .Z(n44089) );
  NAND U53453 ( .A(n44158), .B(n44159), .Z(n44157) );
  NAND U53454 ( .A(n44160), .B(n44161), .Z(n44156) );
  AND U53455 ( .A(n44162), .B(n44163), .Z(n44085) );
  NAND U53456 ( .A(n44164), .B(n44165), .Z(n44163) );
  NAND U53457 ( .A(n44166), .B(n44167), .Z(n44162) );
  NANDN U53458 ( .A(n44168), .B(n44169), .Z(n44088) );
  ANDN U53459 ( .B(n44170), .A(n44171), .Z(n44082) );
  XNOR U53460 ( .A(n44073), .B(n44172), .Z(n44078) );
  XNOR U53461 ( .A(n44071), .B(n44075), .Z(n44172) );
  AND U53462 ( .A(n44173), .B(n44174), .Z(n44075) );
  NAND U53463 ( .A(n44175), .B(n44176), .Z(n44174) );
  NAND U53464 ( .A(n44177), .B(n44178), .Z(n44173) );
  AND U53465 ( .A(n44179), .B(n44180), .Z(n44071) );
  NAND U53466 ( .A(n44181), .B(n44182), .Z(n44180) );
  NAND U53467 ( .A(n44183), .B(n44184), .Z(n44179) );
  AND U53468 ( .A(n44185), .B(n44186), .Z(n44073) );
  XOR U53469 ( .A(n44153), .B(n44152), .Z(N61463) );
  XNOR U53470 ( .A(n44170), .B(n44171), .Z(n44152) );
  XNOR U53471 ( .A(n44185), .B(n44186), .Z(n44171) );
  XOR U53472 ( .A(n44182), .B(n44181), .Z(n44186) );
  XOR U53473 ( .A(y[1620]), .B(x[1620]), .Z(n44181) );
  XOR U53474 ( .A(n44184), .B(n44183), .Z(n44182) );
  XOR U53475 ( .A(y[1622]), .B(x[1622]), .Z(n44183) );
  XOR U53476 ( .A(y[1621]), .B(x[1621]), .Z(n44184) );
  XOR U53477 ( .A(n44176), .B(n44175), .Z(n44185) );
  XOR U53478 ( .A(n44178), .B(n44177), .Z(n44175) );
  XOR U53479 ( .A(y[1619]), .B(x[1619]), .Z(n44177) );
  XOR U53480 ( .A(y[1618]), .B(x[1618]), .Z(n44178) );
  XOR U53481 ( .A(y[1617]), .B(x[1617]), .Z(n44176) );
  XNOR U53482 ( .A(n44169), .B(n44168), .Z(n44170) );
  XNOR U53483 ( .A(n44165), .B(n44164), .Z(n44168) );
  XOR U53484 ( .A(n44167), .B(n44166), .Z(n44164) );
  XOR U53485 ( .A(y[1616]), .B(x[1616]), .Z(n44166) );
  XOR U53486 ( .A(y[1615]), .B(x[1615]), .Z(n44167) );
  XOR U53487 ( .A(y[1614]), .B(x[1614]), .Z(n44165) );
  XOR U53488 ( .A(n44159), .B(n44158), .Z(n44169) );
  XOR U53489 ( .A(n44161), .B(n44160), .Z(n44158) );
  XOR U53490 ( .A(y[1613]), .B(x[1613]), .Z(n44160) );
  XOR U53491 ( .A(y[1612]), .B(x[1612]), .Z(n44161) );
  XOR U53492 ( .A(y[1611]), .B(x[1611]), .Z(n44159) );
  XNOR U53493 ( .A(n44135), .B(n44136), .Z(n44153) );
  XNOR U53494 ( .A(n44150), .B(n44151), .Z(n44136) );
  XOR U53495 ( .A(n44147), .B(n44146), .Z(n44151) );
  XOR U53496 ( .A(y[1608]), .B(x[1608]), .Z(n44146) );
  XOR U53497 ( .A(n44149), .B(n44148), .Z(n44147) );
  XOR U53498 ( .A(y[1610]), .B(x[1610]), .Z(n44148) );
  XOR U53499 ( .A(y[1609]), .B(x[1609]), .Z(n44149) );
  XOR U53500 ( .A(n44141), .B(n44140), .Z(n44150) );
  XOR U53501 ( .A(n44143), .B(n44142), .Z(n44140) );
  XOR U53502 ( .A(y[1607]), .B(x[1607]), .Z(n44142) );
  XOR U53503 ( .A(y[1606]), .B(x[1606]), .Z(n44143) );
  XOR U53504 ( .A(y[1605]), .B(x[1605]), .Z(n44141) );
  XNOR U53505 ( .A(n44134), .B(n44133), .Z(n44135) );
  XNOR U53506 ( .A(n44130), .B(n44129), .Z(n44133) );
  XOR U53507 ( .A(n44132), .B(n44131), .Z(n44129) );
  XOR U53508 ( .A(y[1604]), .B(x[1604]), .Z(n44131) );
  XOR U53509 ( .A(y[1603]), .B(x[1603]), .Z(n44132) );
  XOR U53510 ( .A(y[1602]), .B(x[1602]), .Z(n44130) );
  XOR U53511 ( .A(n44124), .B(n44123), .Z(n44134) );
  XOR U53512 ( .A(n44126), .B(n44125), .Z(n44123) );
  XOR U53513 ( .A(y[1601]), .B(x[1601]), .Z(n44125) );
  XOR U53514 ( .A(y[1600]), .B(x[1600]), .Z(n44126) );
  XOR U53515 ( .A(y[1599]), .B(x[1599]), .Z(n44124) );
  NAND U53516 ( .A(n44187), .B(n44188), .Z(N61454) );
  NAND U53517 ( .A(n44189), .B(n44190), .Z(n44188) );
  NANDN U53518 ( .A(n44191), .B(n44192), .Z(n44190) );
  NANDN U53519 ( .A(n44192), .B(n44191), .Z(n44187) );
  XOR U53520 ( .A(n44191), .B(n44193), .Z(N61453) );
  XNOR U53521 ( .A(n44189), .B(n44192), .Z(n44193) );
  NAND U53522 ( .A(n44194), .B(n44195), .Z(n44192) );
  NAND U53523 ( .A(n44196), .B(n44197), .Z(n44195) );
  NANDN U53524 ( .A(n44198), .B(n44199), .Z(n44197) );
  NANDN U53525 ( .A(n44199), .B(n44198), .Z(n44194) );
  AND U53526 ( .A(n44200), .B(n44201), .Z(n44189) );
  NAND U53527 ( .A(n44202), .B(n44203), .Z(n44201) );
  NANDN U53528 ( .A(n44204), .B(n44205), .Z(n44203) );
  NANDN U53529 ( .A(n44205), .B(n44204), .Z(n44200) );
  IV U53530 ( .A(n44206), .Z(n44205) );
  AND U53531 ( .A(n44207), .B(n44208), .Z(n44191) );
  NAND U53532 ( .A(n44209), .B(n44210), .Z(n44208) );
  NANDN U53533 ( .A(n44211), .B(n44212), .Z(n44210) );
  NANDN U53534 ( .A(n44212), .B(n44211), .Z(n44207) );
  XOR U53535 ( .A(n44204), .B(n44213), .Z(N61452) );
  XNOR U53536 ( .A(n44202), .B(n44206), .Z(n44213) );
  XOR U53537 ( .A(n44199), .B(n44214), .Z(n44206) );
  XNOR U53538 ( .A(n44196), .B(n44198), .Z(n44214) );
  AND U53539 ( .A(n44215), .B(n44216), .Z(n44198) );
  NANDN U53540 ( .A(n44217), .B(n44218), .Z(n44216) );
  OR U53541 ( .A(n44219), .B(n44220), .Z(n44218) );
  IV U53542 ( .A(n44221), .Z(n44220) );
  NANDN U53543 ( .A(n44221), .B(n44219), .Z(n44215) );
  AND U53544 ( .A(n44222), .B(n44223), .Z(n44196) );
  NAND U53545 ( .A(n44224), .B(n44225), .Z(n44223) );
  NANDN U53546 ( .A(n44226), .B(n44227), .Z(n44225) );
  NANDN U53547 ( .A(n44227), .B(n44226), .Z(n44222) );
  IV U53548 ( .A(n44228), .Z(n44227) );
  NAND U53549 ( .A(n44229), .B(n44230), .Z(n44199) );
  NANDN U53550 ( .A(n44231), .B(n44232), .Z(n44230) );
  NANDN U53551 ( .A(n44233), .B(n44234), .Z(n44232) );
  NANDN U53552 ( .A(n44234), .B(n44233), .Z(n44229) );
  IV U53553 ( .A(n44235), .Z(n44233) );
  AND U53554 ( .A(n44236), .B(n44237), .Z(n44202) );
  NAND U53555 ( .A(n44238), .B(n44239), .Z(n44237) );
  NANDN U53556 ( .A(n44240), .B(n44241), .Z(n44239) );
  NANDN U53557 ( .A(n44241), .B(n44240), .Z(n44236) );
  XOR U53558 ( .A(n44212), .B(n44242), .Z(n44204) );
  XNOR U53559 ( .A(n44209), .B(n44211), .Z(n44242) );
  AND U53560 ( .A(n44243), .B(n44244), .Z(n44211) );
  NANDN U53561 ( .A(n44245), .B(n44246), .Z(n44244) );
  OR U53562 ( .A(n44247), .B(n44248), .Z(n44246) );
  IV U53563 ( .A(n44249), .Z(n44248) );
  NANDN U53564 ( .A(n44249), .B(n44247), .Z(n44243) );
  AND U53565 ( .A(n44250), .B(n44251), .Z(n44209) );
  NAND U53566 ( .A(n44252), .B(n44253), .Z(n44251) );
  NANDN U53567 ( .A(n44254), .B(n44255), .Z(n44253) );
  NANDN U53568 ( .A(n44255), .B(n44254), .Z(n44250) );
  IV U53569 ( .A(n44256), .Z(n44255) );
  NAND U53570 ( .A(n44257), .B(n44258), .Z(n44212) );
  NANDN U53571 ( .A(n44259), .B(n44260), .Z(n44258) );
  NANDN U53572 ( .A(n44261), .B(n44262), .Z(n44260) );
  NANDN U53573 ( .A(n44262), .B(n44261), .Z(n44257) );
  IV U53574 ( .A(n44263), .Z(n44261) );
  XOR U53575 ( .A(n44238), .B(n44264), .Z(N61451) );
  XNOR U53576 ( .A(n44241), .B(n44240), .Z(n44264) );
  XNOR U53577 ( .A(n44252), .B(n44265), .Z(n44240) );
  XNOR U53578 ( .A(n44256), .B(n44254), .Z(n44265) );
  XOR U53579 ( .A(n44262), .B(n44266), .Z(n44254) );
  XNOR U53580 ( .A(n44259), .B(n44263), .Z(n44266) );
  AND U53581 ( .A(n44267), .B(n44268), .Z(n44263) );
  NAND U53582 ( .A(n44269), .B(n44270), .Z(n44268) );
  NAND U53583 ( .A(n44271), .B(n44272), .Z(n44267) );
  AND U53584 ( .A(n44273), .B(n44274), .Z(n44259) );
  NAND U53585 ( .A(n44275), .B(n44276), .Z(n44274) );
  NAND U53586 ( .A(n44277), .B(n44278), .Z(n44273) );
  NANDN U53587 ( .A(n44279), .B(n44280), .Z(n44262) );
  ANDN U53588 ( .B(n44281), .A(n44282), .Z(n44256) );
  XNOR U53589 ( .A(n44247), .B(n44283), .Z(n44252) );
  XNOR U53590 ( .A(n44245), .B(n44249), .Z(n44283) );
  AND U53591 ( .A(n44284), .B(n44285), .Z(n44249) );
  NAND U53592 ( .A(n44286), .B(n44287), .Z(n44285) );
  NAND U53593 ( .A(n44288), .B(n44289), .Z(n44284) );
  AND U53594 ( .A(n44290), .B(n44291), .Z(n44245) );
  NAND U53595 ( .A(n44292), .B(n44293), .Z(n44291) );
  NAND U53596 ( .A(n44294), .B(n44295), .Z(n44290) );
  AND U53597 ( .A(n44296), .B(n44297), .Z(n44247) );
  NAND U53598 ( .A(n44298), .B(n44299), .Z(n44241) );
  XNOR U53599 ( .A(n44224), .B(n44300), .Z(n44238) );
  XNOR U53600 ( .A(n44228), .B(n44226), .Z(n44300) );
  XOR U53601 ( .A(n44234), .B(n44301), .Z(n44226) );
  XNOR U53602 ( .A(n44231), .B(n44235), .Z(n44301) );
  AND U53603 ( .A(n44302), .B(n44303), .Z(n44235) );
  NAND U53604 ( .A(n44304), .B(n44305), .Z(n44303) );
  NAND U53605 ( .A(n44306), .B(n44307), .Z(n44302) );
  AND U53606 ( .A(n44308), .B(n44309), .Z(n44231) );
  NAND U53607 ( .A(n44310), .B(n44311), .Z(n44309) );
  NAND U53608 ( .A(n44312), .B(n44313), .Z(n44308) );
  NANDN U53609 ( .A(n44314), .B(n44315), .Z(n44234) );
  ANDN U53610 ( .B(n44316), .A(n44317), .Z(n44228) );
  XNOR U53611 ( .A(n44219), .B(n44318), .Z(n44224) );
  XNOR U53612 ( .A(n44217), .B(n44221), .Z(n44318) );
  AND U53613 ( .A(n44319), .B(n44320), .Z(n44221) );
  NAND U53614 ( .A(n44321), .B(n44322), .Z(n44320) );
  NAND U53615 ( .A(n44323), .B(n44324), .Z(n44319) );
  AND U53616 ( .A(n44325), .B(n44326), .Z(n44217) );
  NAND U53617 ( .A(n44327), .B(n44328), .Z(n44326) );
  NAND U53618 ( .A(n44329), .B(n44330), .Z(n44325) );
  AND U53619 ( .A(n44331), .B(n44332), .Z(n44219) );
  XOR U53620 ( .A(n44299), .B(n44298), .Z(N61450) );
  XNOR U53621 ( .A(n44316), .B(n44317), .Z(n44298) );
  XNOR U53622 ( .A(n44331), .B(n44332), .Z(n44317) );
  XOR U53623 ( .A(n44328), .B(n44327), .Z(n44332) );
  XOR U53624 ( .A(y[1596]), .B(x[1596]), .Z(n44327) );
  XOR U53625 ( .A(n44330), .B(n44329), .Z(n44328) );
  XOR U53626 ( .A(y[1598]), .B(x[1598]), .Z(n44329) );
  XOR U53627 ( .A(y[1597]), .B(x[1597]), .Z(n44330) );
  XOR U53628 ( .A(n44322), .B(n44321), .Z(n44331) );
  XOR U53629 ( .A(n44324), .B(n44323), .Z(n44321) );
  XOR U53630 ( .A(y[1595]), .B(x[1595]), .Z(n44323) );
  XOR U53631 ( .A(y[1594]), .B(x[1594]), .Z(n44324) );
  XOR U53632 ( .A(y[1593]), .B(x[1593]), .Z(n44322) );
  XNOR U53633 ( .A(n44315), .B(n44314), .Z(n44316) );
  XNOR U53634 ( .A(n44311), .B(n44310), .Z(n44314) );
  XOR U53635 ( .A(n44313), .B(n44312), .Z(n44310) );
  XOR U53636 ( .A(y[1592]), .B(x[1592]), .Z(n44312) );
  XOR U53637 ( .A(y[1591]), .B(x[1591]), .Z(n44313) );
  XOR U53638 ( .A(y[1590]), .B(x[1590]), .Z(n44311) );
  XOR U53639 ( .A(n44305), .B(n44304), .Z(n44315) );
  XOR U53640 ( .A(n44307), .B(n44306), .Z(n44304) );
  XOR U53641 ( .A(y[1589]), .B(x[1589]), .Z(n44306) );
  XOR U53642 ( .A(y[1588]), .B(x[1588]), .Z(n44307) );
  XOR U53643 ( .A(y[1587]), .B(x[1587]), .Z(n44305) );
  XNOR U53644 ( .A(n44281), .B(n44282), .Z(n44299) );
  XNOR U53645 ( .A(n44296), .B(n44297), .Z(n44282) );
  XOR U53646 ( .A(n44293), .B(n44292), .Z(n44297) );
  XOR U53647 ( .A(y[1584]), .B(x[1584]), .Z(n44292) );
  XOR U53648 ( .A(n44295), .B(n44294), .Z(n44293) );
  XOR U53649 ( .A(y[1586]), .B(x[1586]), .Z(n44294) );
  XOR U53650 ( .A(y[1585]), .B(x[1585]), .Z(n44295) );
  XOR U53651 ( .A(n44287), .B(n44286), .Z(n44296) );
  XOR U53652 ( .A(n44289), .B(n44288), .Z(n44286) );
  XOR U53653 ( .A(y[1583]), .B(x[1583]), .Z(n44288) );
  XOR U53654 ( .A(y[1582]), .B(x[1582]), .Z(n44289) );
  XOR U53655 ( .A(y[1581]), .B(x[1581]), .Z(n44287) );
  XNOR U53656 ( .A(n44280), .B(n44279), .Z(n44281) );
  XNOR U53657 ( .A(n44276), .B(n44275), .Z(n44279) );
  XOR U53658 ( .A(n44278), .B(n44277), .Z(n44275) );
  XOR U53659 ( .A(y[1580]), .B(x[1580]), .Z(n44277) );
  XOR U53660 ( .A(y[1579]), .B(x[1579]), .Z(n44278) );
  XOR U53661 ( .A(y[1578]), .B(x[1578]), .Z(n44276) );
  XOR U53662 ( .A(n44270), .B(n44269), .Z(n44280) );
  XOR U53663 ( .A(n44272), .B(n44271), .Z(n44269) );
  XOR U53664 ( .A(y[1577]), .B(x[1577]), .Z(n44271) );
  XOR U53665 ( .A(y[1576]), .B(x[1576]), .Z(n44272) );
  XOR U53666 ( .A(y[1575]), .B(x[1575]), .Z(n44270) );
  NAND U53667 ( .A(n44333), .B(n44334), .Z(N61441) );
  NAND U53668 ( .A(n44335), .B(n44336), .Z(n44334) );
  NANDN U53669 ( .A(n44337), .B(n44338), .Z(n44336) );
  NANDN U53670 ( .A(n44338), .B(n44337), .Z(n44333) );
  XOR U53671 ( .A(n44337), .B(n44339), .Z(N61440) );
  XNOR U53672 ( .A(n44335), .B(n44338), .Z(n44339) );
  NAND U53673 ( .A(n44340), .B(n44341), .Z(n44338) );
  NAND U53674 ( .A(n44342), .B(n44343), .Z(n44341) );
  NANDN U53675 ( .A(n44344), .B(n44345), .Z(n44343) );
  NANDN U53676 ( .A(n44345), .B(n44344), .Z(n44340) );
  AND U53677 ( .A(n44346), .B(n44347), .Z(n44335) );
  NAND U53678 ( .A(n44348), .B(n44349), .Z(n44347) );
  NANDN U53679 ( .A(n44350), .B(n44351), .Z(n44349) );
  NANDN U53680 ( .A(n44351), .B(n44350), .Z(n44346) );
  IV U53681 ( .A(n44352), .Z(n44351) );
  AND U53682 ( .A(n44353), .B(n44354), .Z(n44337) );
  NAND U53683 ( .A(n44355), .B(n44356), .Z(n44354) );
  NANDN U53684 ( .A(n44357), .B(n44358), .Z(n44356) );
  NANDN U53685 ( .A(n44358), .B(n44357), .Z(n44353) );
  XOR U53686 ( .A(n44350), .B(n44359), .Z(N61439) );
  XNOR U53687 ( .A(n44348), .B(n44352), .Z(n44359) );
  XOR U53688 ( .A(n44345), .B(n44360), .Z(n44352) );
  XNOR U53689 ( .A(n44342), .B(n44344), .Z(n44360) );
  AND U53690 ( .A(n44361), .B(n44362), .Z(n44344) );
  NANDN U53691 ( .A(n44363), .B(n44364), .Z(n44362) );
  OR U53692 ( .A(n44365), .B(n44366), .Z(n44364) );
  IV U53693 ( .A(n44367), .Z(n44366) );
  NANDN U53694 ( .A(n44367), .B(n44365), .Z(n44361) );
  AND U53695 ( .A(n44368), .B(n44369), .Z(n44342) );
  NAND U53696 ( .A(n44370), .B(n44371), .Z(n44369) );
  NANDN U53697 ( .A(n44372), .B(n44373), .Z(n44371) );
  NANDN U53698 ( .A(n44373), .B(n44372), .Z(n44368) );
  IV U53699 ( .A(n44374), .Z(n44373) );
  NAND U53700 ( .A(n44375), .B(n44376), .Z(n44345) );
  NANDN U53701 ( .A(n44377), .B(n44378), .Z(n44376) );
  NANDN U53702 ( .A(n44379), .B(n44380), .Z(n44378) );
  NANDN U53703 ( .A(n44380), .B(n44379), .Z(n44375) );
  IV U53704 ( .A(n44381), .Z(n44379) );
  AND U53705 ( .A(n44382), .B(n44383), .Z(n44348) );
  NAND U53706 ( .A(n44384), .B(n44385), .Z(n44383) );
  NANDN U53707 ( .A(n44386), .B(n44387), .Z(n44385) );
  NANDN U53708 ( .A(n44387), .B(n44386), .Z(n44382) );
  XOR U53709 ( .A(n44358), .B(n44388), .Z(n44350) );
  XNOR U53710 ( .A(n44355), .B(n44357), .Z(n44388) );
  AND U53711 ( .A(n44389), .B(n44390), .Z(n44357) );
  NANDN U53712 ( .A(n44391), .B(n44392), .Z(n44390) );
  OR U53713 ( .A(n44393), .B(n44394), .Z(n44392) );
  IV U53714 ( .A(n44395), .Z(n44394) );
  NANDN U53715 ( .A(n44395), .B(n44393), .Z(n44389) );
  AND U53716 ( .A(n44396), .B(n44397), .Z(n44355) );
  NAND U53717 ( .A(n44398), .B(n44399), .Z(n44397) );
  NANDN U53718 ( .A(n44400), .B(n44401), .Z(n44399) );
  NANDN U53719 ( .A(n44401), .B(n44400), .Z(n44396) );
  IV U53720 ( .A(n44402), .Z(n44401) );
  NAND U53721 ( .A(n44403), .B(n44404), .Z(n44358) );
  NANDN U53722 ( .A(n44405), .B(n44406), .Z(n44404) );
  NANDN U53723 ( .A(n44407), .B(n44408), .Z(n44406) );
  NANDN U53724 ( .A(n44408), .B(n44407), .Z(n44403) );
  IV U53725 ( .A(n44409), .Z(n44407) );
  XOR U53726 ( .A(n44384), .B(n44410), .Z(N61438) );
  XNOR U53727 ( .A(n44387), .B(n44386), .Z(n44410) );
  XNOR U53728 ( .A(n44398), .B(n44411), .Z(n44386) );
  XNOR U53729 ( .A(n44402), .B(n44400), .Z(n44411) );
  XOR U53730 ( .A(n44408), .B(n44412), .Z(n44400) );
  XNOR U53731 ( .A(n44405), .B(n44409), .Z(n44412) );
  AND U53732 ( .A(n44413), .B(n44414), .Z(n44409) );
  NAND U53733 ( .A(n44415), .B(n44416), .Z(n44414) );
  NAND U53734 ( .A(n44417), .B(n44418), .Z(n44413) );
  AND U53735 ( .A(n44419), .B(n44420), .Z(n44405) );
  NAND U53736 ( .A(n44421), .B(n44422), .Z(n44420) );
  NAND U53737 ( .A(n44423), .B(n44424), .Z(n44419) );
  NANDN U53738 ( .A(n44425), .B(n44426), .Z(n44408) );
  ANDN U53739 ( .B(n44427), .A(n44428), .Z(n44402) );
  XNOR U53740 ( .A(n44393), .B(n44429), .Z(n44398) );
  XNOR U53741 ( .A(n44391), .B(n44395), .Z(n44429) );
  AND U53742 ( .A(n44430), .B(n44431), .Z(n44395) );
  NAND U53743 ( .A(n44432), .B(n44433), .Z(n44431) );
  NAND U53744 ( .A(n44434), .B(n44435), .Z(n44430) );
  AND U53745 ( .A(n44436), .B(n44437), .Z(n44391) );
  NAND U53746 ( .A(n44438), .B(n44439), .Z(n44437) );
  NAND U53747 ( .A(n44440), .B(n44441), .Z(n44436) );
  AND U53748 ( .A(n44442), .B(n44443), .Z(n44393) );
  NAND U53749 ( .A(n44444), .B(n44445), .Z(n44387) );
  XNOR U53750 ( .A(n44370), .B(n44446), .Z(n44384) );
  XNOR U53751 ( .A(n44374), .B(n44372), .Z(n44446) );
  XOR U53752 ( .A(n44380), .B(n44447), .Z(n44372) );
  XNOR U53753 ( .A(n44377), .B(n44381), .Z(n44447) );
  AND U53754 ( .A(n44448), .B(n44449), .Z(n44381) );
  NAND U53755 ( .A(n44450), .B(n44451), .Z(n44449) );
  NAND U53756 ( .A(n44452), .B(n44453), .Z(n44448) );
  AND U53757 ( .A(n44454), .B(n44455), .Z(n44377) );
  NAND U53758 ( .A(n44456), .B(n44457), .Z(n44455) );
  NAND U53759 ( .A(n44458), .B(n44459), .Z(n44454) );
  NANDN U53760 ( .A(n44460), .B(n44461), .Z(n44380) );
  ANDN U53761 ( .B(n44462), .A(n44463), .Z(n44374) );
  XNOR U53762 ( .A(n44365), .B(n44464), .Z(n44370) );
  XNOR U53763 ( .A(n44363), .B(n44367), .Z(n44464) );
  AND U53764 ( .A(n44465), .B(n44466), .Z(n44367) );
  NAND U53765 ( .A(n44467), .B(n44468), .Z(n44466) );
  NAND U53766 ( .A(n44469), .B(n44470), .Z(n44465) );
  AND U53767 ( .A(n44471), .B(n44472), .Z(n44363) );
  NAND U53768 ( .A(n44473), .B(n44474), .Z(n44472) );
  NAND U53769 ( .A(n44475), .B(n44476), .Z(n44471) );
  AND U53770 ( .A(n44477), .B(n44478), .Z(n44365) );
  XOR U53771 ( .A(n44445), .B(n44444), .Z(N61437) );
  XNOR U53772 ( .A(n44462), .B(n44463), .Z(n44444) );
  XNOR U53773 ( .A(n44477), .B(n44478), .Z(n44463) );
  XOR U53774 ( .A(n44474), .B(n44473), .Z(n44478) );
  XOR U53775 ( .A(y[1572]), .B(x[1572]), .Z(n44473) );
  XOR U53776 ( .A(n44476), .B(n44475), .Z(n44474) );
  XOR U53777 ( .A(y[1574]), .B(x[1574]), .Z(n44475) );
  XOR U53778 ( .A(y[1573]), .B(x[1573]), .Z(n44476) );
  XOR U53779 ( .A(n44468), .B(n44467), .Z(n44477) );
  XOR U53780 ( .A(n44470), .B(n44469), .Z(n44467) );
  XOR U53781 ( .A(y[1571]), .B(x[1571]), .Z(n44469) );
  XOR U53782 ( .A(y[1570]), .B(x[1570]), .Z(n44470) );
  XOR U53783 ( .A(y[1569]), .B(x[1569]), .Z(n44468) );
  XNOR U53784 ( .A(n44461), .B(n44460), .Z(n44462) );
  XNOR U53785 ( .A(n44457), .B(n44456), .Z(n44460) );
  XOR U53786 ( .A(n44459), .B(n44458), .Z(n44456) );
  XOR U53787 ( .A(y[1568]), .B(x[1568]), .Z(n44458) );
  XOR U53788 ( .A(y[1567]), .B(x[1567]), .Z(n44459) );
  XOR U53789 ( .A(y[1566]), .B(x[1566]), .Z(n44457) );
  XOR U53790 ( .A(n44451), .B(n44450), .Z(n44461) );
  XOR U53791 ( .A(n44453), .B(n44452), .Z(n44450) );
  XOR U53792 ( .A(y[1565]), .B(x[1565]), .Z(n44452) );
  XOR U53793 ( .A(y[1564]), .B(x[1564]), .Z(n44453) );
  XOR U53794 ( .A(y[1563]), .B(x[1563]), .Z(n44451) );
  XNOR U53795 ( .A(n44427), .B(n44428), .Z(n44445) );
  XNOR U53796 ( .A(n44442), .B(n44443), .Z(n44428) );
  XOR U53797 ( .A(n44439), .B(n44438), .Z(n44443) );
  XOR U53798 ( .A(y[1560]), .B(x[1560]), .Z(n44438) );
  XOR U53799 ( .A(n44441), .B(n44440), .Z(n44439) );
  XOR U53800 ( .A(y[1562]), .B(x[1562]), .Z(n44440) );
  XOR U53801 ( .A(y[1561]), .B(x[1561]), .Z(n44441) );
  XOR U53802 ( .A(n44433), .B(n44432), .Z(n44442) );
  XOR U53803 ( .A(n44435), .B(n44434), .Z(n44432) );
  XOR U53804 ( .A(y[1559]), .B(x[1559]), .Z(n44434) );
  XOR U53805 ( .A(y[1558]), .B(x[1558]), .Z(n44435) );
  XOR U53806 ( .A(y[1557]), .B(x[1557]), .Z(n44433) );
  XNOR U53807 ( .A(n44426), .B(n44425), .Z(n44427) );
  XNOR U53808 ( .A(n44422), .B(n44421), .Z(n44425) );
  XOR U53809 ( .A(n44424), .B(n44423), .Z(n44421) );
  XOR U53810 ( .A(y[1556]), .B(x[1556]), .Z(n44423) );
  XOR U53811 ( .A(y[1555]), .B(x[1555]), .Z(n44424) );
  XOR U53812 ( .A(y[1554]), .B(x[1554]), .Z(n44422) );
  XOR U53813 ( .A(n44416), .B(n44415), .Z(n44426) );
  XOR U53814 ( .A(n44418), .B(n44417), .Z(n44415) );
  XOR U53815 ( .A(y[1553]), .B(x[1553]), .Z(n44417) );
  XOR U53816 ( .A(y[1552]), .B(x[1552]), .Z(n44418) );
  XOR U53817 ( .A(y[1551]), .B(x[1551]), .Z(n44416) );
  NAND U53818 ( .A(n44479), .B(n44480), .Z(N61428) );
  NAND U53819 ( .A(n44481), .B(n44482), .Z(n44480) );
  NANDN U53820 ( .A(n44483), .B(n44484), .Z(n44482) );
  NANDN U53821 ( .A(n44484), .B(n44483), .Z(n44479) );
  XOR U53822 ( .A(n44483), .B(n44485), .Z(N61427) );
  XNOR U53823 ( .A(n44481), .B(n44484), .Z(n44485) );
  NAND U53824 ( .A(n44486), .B(n44487), .Z(n44484) );
  NAND U53825 ( .A(n44488), .B(n44489), .Z(n44487) );
  NANDN U53826 ( .A(n44490), .B(n44491), .Z(n44489) );
  NANDN U53827 ( .A(n44491), .B(n44490), .Z(n44486) );
  AND U53828 ( .A(n44492), .B(n44493), .Z(n44481) );
  NAND U53829 ( .A(n44494), .B(n44495), .Z(n44493) );
  NANDN U53830 ( .A(n44496), .B(n44497), .Z(n44495) );
  NANDN U53831 ( .A(n44497), .B(n44496), .Z(n44492) );
  IV U53832 ( .A(n44498), .Z(n44497) );
  AND U53833 ( .A(n44499), .B(n44500), .Z(n44483) );
  NAND U53834 ( .A(n44501), .B(n44502), .Z(n44500) );
  NANDN U53835 ( .A(n44503), .B(n44504), .Z(n44502) );
  NANDN U53836 ( .A(n44504), .B(n44503), .Z(n44499) );
  XOR U53837 ( .A(n44496), .B(n44505), .Z(N61426) );
  XNOR U53838 ( .A(n44494), .B(n44498), .Z(n44505) );
  XOR U53839 ( .A(n44491), .B(n44506), .Z(n44498) );
  XNOR U53840 ( .A(n44488), .B(n44490), .Z(n44506) );
  AND U53841 ( .A(n44507), .B(n44508), .Z(n44490) );
  NANDN U53842 ( .A(n44509), .B(n44510), .Z(n44508) );
  OR U53843 ( .A(n44511), .B(n44512), .Z(n44510) );
  IV U53844 ( .A(n44513), .Z(n44512) );
  NANDN U53845 ( .A(n44513), .B(n44511), .Z(n44507) );
  AND U53846 ( .A(n44514), .B(n44515), .Z(n44488) );
  NAND U53847 ( .A(n44516), .B(n44517), .Z(n44515) );
  NANDN U53848 ( .A(n44518), .B(n44519), .Z(n44517) );
  NANDN U53849 ( .A(n44519), .B(n44518), .Z(n44514) );
  IV U53850 ( .A(n44520), .Z(n44519) );
  NAND U53851 ( .A(n44521), .B(n44522), .Z(n44491) );
  NANDN U53852 ( .A(n44523), .B(n44524), .Z(n44522) );
  NANDN U53853 ( .A(n44525), .B(n44526), .Z(n44524) );
  NANDN U53854 ( .A(n44526), .B(n44525), .Z(n44521) );
  IV U53855 ( .A(n44527), .Z(n44525) );
  AND U53856 ( .A(n44528), .B(n44529), .Z(n44494) );
  NAND U53857 ( .A(n44530), .B(n44531), .Z(n44529) );
  NANDN U53858 ( .A(n44532), .B(n44533), .Z(n44531) );
  NANDN U53859 ( .A(n44533), .B(n44532), .Z(n44528) );
  XOR U53860 ( .A(n44504), .B(n44534), .Z(n44496) );
  XNOR U53861 ( .A(n44501), .B(n44503), .Z(n44534) );
  AND U53862 ( .A(n44535), .B(n44536), .Z(n44503) );
  NANDN U53863 ( .A(n44537), .B(n44538), .Z(n44536) );
  OR U53864 ( .A(n44539), .B(n44540), .Z(n44538) );
  IV U53865 ( .A(n44541), .Z(n44540) );
  NANDN U53866 ( .A(n44541), .B(n44539), .Z(n44535) );
  AND U53867 ( .A(n44542), .B(n44543), .Z(n44501) );
  NAND U53868 ( .A(n44544), .B(n44545), .Z(n44543) );
  NANDN U53869 ( .A(n44546), .B(n44547), .Z(n44545) );
  NANDN U53870 ( .A(n44547), .B(n44546), .Z(n44542) );
  IV U53871 ( .A(n44548), .Z(n44547) );
  NAND U53872 ( .A(n44549), .B(n44550), .Z(n44504) );
  NANDN U53873 ( .A(n44551), .B(n44552), .Z(n44550) );
  NANDN U53874 ( .A(n44553), .B(n44554), .Z(n44552) );
  NANDN U53875 ( .A(n44554), .B(n44553), .Z(n44549) );
  IV U53876 ( .A(n44555), .Z(n44553) );
  XOR U53877 ( .A(n44530), .B(n44556), .Z(N61425) );
  XNOR U53878 ( .A(n44533), .B(n44532), .Z(n44556) );
  XNOR U53879 ( .A(n44544), .B(n44557), .Z(n44532) );
  XNOR U53880 ( .A(n44548), .B(n44546), .Z(n44557) );
  XOR U53881 ( .A(n44554), .B(n44558), .Z(n44546) );
  XNOR U53882 ( .A(n44551), .B(n44555), .Z(n44558) );
  AND U53883 ( .A(n44559), .B(n44560), .Z(n44555) );
  NAND U53884 ( .A(n44561), .B(n44562), .Z(n44560) );
  NAND U53885 ( .A(n44563), .B(n44564), .Z(n44559) );
  AND U53886 ( .A(n44565), .B(n44566), .Z(n44551) );
  NAND U53887 ( .A(n44567), .B(n44568), .Z(n44566) );
  NAND U53888 ( .A(n44569), .B(n44570), .Z(n44565) );
  NANDN U53889 ( .A(n44571), .B(n44572), .Z(n44554) );
  ANDN U53890 ( .B(n44573), .A(n44574), .Z(n44548) );
  XNOR U53891 ( .A(n44539), .B(n44575), .Z(n44544) );
  XNOR U53892 ( .A(n44537), .B(n44541), .Z(n44575) );
  AND U53893 ( .A(n44576), .B(n44577), .Z(n44541) );
  NAND U53894 ( .A(n44578), .B(n44579), .Z(n44577) );
  NAND U53895 ( .A(n44580), .B(n44581), .Z(n44576) );
  AND U53896 ( .A(n44582), .B(n44583), .Z(n44537) );
  NAND U53897 ( .A(n44584), .B(n44585), .Z(n44583) );
  NAND U53898 ( .A(n44586), .B(n44587), .Z(n44582) );
  AND U53899 ( .A(n44588), .B(n44589), .Z(n44539) );
  NAND U53900 ( .A(n44590), .B(n44591), .Z(n44533) );
  XNOR U53901 ( .A(n44516), .B(n44592), .Z(n44530) );
  XNOR U53902 ( .A(n44520), .B(n44518), .Z(n44592) );
  XOR U53903 ( .A(n44526), .B(n44593), .Z(n44518) );
  XNOR U53904 ( .A(n44523), .B(n44527), .Z(n44593) );
  AND U53905 ( .A(n44594), .B(n44595), .Z(n44527) );
  NAND U53906 ( .A(n44596), .B(n44597), .Z(n44595) );
  NAND U53907 ( .A(n44598), .B(n44599), .Z(n44594) );
  AND U53908 ( .A(n44600), .B(n44601), .Z(n44523) );
  NAND U53909 ( .A(n44602), .B(n44603), .Z(n44601) );
  NAND U53910 ( .A(n44604), .B(n44605), .Z(n44600) );
  NANDN U53911 ( .A(n44606), .B(n44607), .Z(n44526) );
  ANDN U53912 ( .B(n44608), .A(n44609), .Z(n44520) );
  XNOR U53913 ( .A(n44511), .B(n44610), .Z(n44516) );
  XNOR U53914 ( .A(n44509), .B(n44513), .Z(n44610) );
  AND U53915 ( .A(n44611), .B(n44612), .Z(n44513) );
  NAND U53916 ( .A(n44613), .B(n44614), .Z(n44612) );
  NAND U53917 ( .A(n44615), .B(n44616), .Z(n44611) );
  AND U53918 ( .A(n44617), .B(n44618), .Z(n44509) );
  NAND U53919 ( .A(n44619), .B(n44620), .Z(n44618) );
  NAND U53920 ( .A(n44621), .B(n44622), .Z(n44617) );
  AND U53921 ( .A(n44623), .B(n44624), .Z(n44511) );
  XOR U53922 ( .A(n44591), .B(n44590), .Z(N61424) );
  XNOR U53923 ( .A(n44608), .B(n44609), .Z(n44590) );
  XNOR U53924 ( .A(n44623), .B(n44624), .Z(n44609) );
  XOR U53925 ( .A(n44620), .B(n44619), .Z(n44624) );
  XOR U53926 ( .A(y[1548]), .B(x[1548]), .Z(n44619) );
  XOR U53927 ( .A(n44622), .B(n44621), .Z(n44620) );
  XOR U53928 ( .A(y[1550]), .B(x[1550]), .Z(n44621) );
  XOR U53929 ( .A(y[1549]), .B(x[1549]), .Z(n44622) );
  XOR U53930 ( .A(n44614), .B(n44613), .Z(n44623) );
  XOR U53931 ( .A(n44616), .B(n44615), .Z(n44613) );
  XOR U53932 ( .A(y[1547]), .B(x[1547]), .Z(n44615) );
  XOR U53933 ( .A(y[1546]), .B(x[1546]), .Z(n44616) );
  XOR U53934 ( .A(y[1545]), .B(x[1545]), .Z(n44614) );
  XNOR U53935 ( .A(n44607), .B(n44606), .Z(n44608) );
  XNOR U53936 ( .A(n44603), .B(n44602), .Z(n44606) );
  XOR U53937 ( .A(n44605), .B(n44604), .Z(n44602) );
  XOR U53938 ( .A(y[1544]), .B(x[1544]), .Z(n44604) );
  XOR U53939 ( .A(y[1543]), .B(x[1543]), .Z(n44605) );
  XOR U53940 ( .A(y[1542]), .B(x[1542]), .Z(n44603) );
  XOR U53941 ( .A(n44597), .B(n44596), .Z(n44607) );
  XOR U53942 ( .A(n44599), .B(n44598), .Z(n44596) );
  XOR U53943 ( .A(y[1541]), .B(x[1541]), .Z(n44598) );
  XOR U53944 ( .A(y[1540]), .B(x[1540]), .Z(n44599) );
  XOR U53945 ( .A(y[1539]), .B(x[1539]), .Z(n44597) );
  XNOR U53946 ( .A(n44573), .B(n44574), .Z(n44591) );
  XNOR U53947 ( .A(n44588), .B(n44589), .Z(n44574) );
  XOR U53948 ( .A(n44585), .B(n44584), .Z(n44589) );
  XOR U53949 ( .A(y[1536]), .B(x[1536]), .Z(n44584) );
  XOR U53950 ( .A(n44587), .B(n44586), .Z(n44585) );
  XOR U53951 ( .A(y[1538]), .B(x[1538]), .Z(n44586) );
  XOR U53952 ( .A(y[1537]), .B(x[1537]), .Z(n44587) );
  XOR U53953 ( .A(n44579), .B(n44578), .Z(n44588) );
  XOR U53954 ( .A(n44581), .B(n44580), .Z(n44578) );
  XOR U53955 ( .A(y[1535]), .B(x[1535]), .Z(n44580) );
  XOR U53956 ( .A(y[1534]), .B(x[1534]), .Z(n44581) );
  XOR U53957 ( .A(y[1533]), .B(x[1533]), .Z(n44579) );
  XNOR U53958 ( .A(n44572), .B(n44571), .Z(n44573) );
  XNOR U53959 ( .A(n44568), .B(n44567), .Z(n44571) );
  XOR U53960 ( .A(n44570), .B(n44569), .Z(n44567) );
  XOR U53961 ( .A(y[1532]), .B(x[1532]), .Z(n44569) );
  XOR U53962 ( .A(y[1531]), .B(x[1531]), .Z(n44570) );
  XOR U53963 ( .A(y[1530]), .B(x[1530]), .Z(n44568) );
  XOR U53964 ( .A(n44562), .B(n44561), .Z(n44572) );
  XOR U53965 ( .A(n44564), .B(n44563), .Z(n44561) );
  XOR U53966 ( .A(y[1529]), .B(x[1529]), .Z(n44563) );
  XOR U53967 ( .A(y[1528]), .B(x[1528]), .Z(n44564) );
  XOR U53968 ( .A(y[1527]), .B(x[1527]), .Z(n44562) );
  NAND U53969 ( .A(n44625), .B(n44626), .Z(N61415) );
  NAND U53970 ( .A(n44627), .B(n44628), .Z(n44626) );
  NANDN U53971 ( .A(n44629), .B(n44630), .Z(n44628) );
  NANDN U53972 ( .A(n44630), .B(n44629), .Z(n44625) );
  XOR U53973 ( .A(n44629), .B(n44631), .Z(N61414) );
  XNOR U53974 ( .A(n44627), .B(n44630), .Z(n44631) );
  NAND U53975 ( .A(n44632), .B(n44633), .Z(n44630) );
  NAND U53976 ( .A(n44634), .B(n44635), .Z(n44633) );
  NANDN U53977 ( .A(n44636), .B(n44637), .Z(n44635) );
  NANDN U53978 ( .A(n44637), .B(n44636), .Z(n44632) );
  AND U53979 ( .A(n44638), .B(n44639), .Z(n44627) );
  NAND U53980 ( .A(n44640), .B(n44641), .Z(n44639) );
  NANDN U53981 ( .A(n44642), .B(n44643), .Z(n44641) );
  NANDN U53982 ( .A(n44643), .B(n44642), .Z(n44638) );
  IV U53983 ( .A(n44644), .Z(n44643) );
  AND U53984 ( .A(n44645), .B(n44646), .Z(n44629) );
  NAND U53985 ( .A(n44647), .B(n44648), .Z(n44646) );
  NANDN U53986 ( .A(n44649), .B(n44650), .Z(n44648) );
  NANDN U53987 ( .A(n44650), .B(n44649), .Z(n44645) );
  XOR U53988 ( .A(n44642), .B(n44651), .Z(N61413) );
  XNOR U53989 ( .A(n44640), .B(n44644), .Z(n44651) );
  XOR U53990 ( .A(n44637), .B(n44652), .Z(n44644) );
  XNOR U53991 ( .A(n44634), .B(n44636), .Z(n44652) );
  AND U53992 ( .A(n44653), .B(n44654), .Z(n44636) );
  NANDN U53993 ( .A(n44655), .B(n44656), .Z(n44654) );
  OR U53994 ( .A(n44657), .B(n44658), .Z(n44656) );
  IV U53995 ( .A(n44659), .Z(n44658) );
  NANDN U53996 ( .A(n44659), .B(n44657), .Z(n44653) );
  AND U53997 ( .A(n44660), .B(n44661), .Z(n44634) );
  NAND U53998 ( .A(n44662), .B(n44663), .Z(n44661) );
  NANDN U53999 ( .A(n44664), .B(n44665), .Z(n44663) );
  NANDN U54000 ( .A(n44665), .B(n44664), .Z(n44660) );
  IV U54001 ( .A(n44666), .Z(n44665) );
  NAND U54002 ( .A(n44667), .B(n44668), .Z(n44637) );
  NANDN U54003 ( .A(n44669), .B(n44670), .Z(n44668) );
  NANDN U54004 ( .A(n44671), .B(n44672), .Z(n44670) );
  NANDN U54005 ( .A(n44672), .B(n44671), .Z(n44667) );
  IV U54006 ( .A(n44673), .Z(n44671) );
  AND U54007 ( .A(n44674), .B(n44675), .Z(n44640) );
  NAND U54008 ( .A(n44676), .B(n44677), .Z(n44675) );
  NANDN U54009 ( .A(n44678), .B(n44679), .Z(n44677) );
  NANDN U54010 ( .A(n44679), .B(n44678), .Z(n44674) );
  XOR U54011 ( .A(n44650), .B(n44680), .Z(n44642) );
  XNOR U54012 ( .A(n44647), .B(n44649), .Z(n44680) );
  AND U54013 ( .A(n44681), .B(n44682), .Z(n44649) );
  NANDN U54014 ( .A(n44683), .B(n44684), .Z(n44682) );
  OR U54015 ( .A(n44685), .B(n44686), .Z(n44684) );
  IV U54016 ( .A(n44687), .Z(n44686) );
  NANDN U54017 ( .A(n44687), .B(n44685), .Z(n44681) );
  AND U54018 ( .A(n44688), .B(n44689), .Z(n44647) );
  NAND U54019 ( .A(n44690), .B(n44691), .Z(n44689) );
  NANDN U54020 ( .A(n44692), .B(n44693), .Z(n44691) );
  NANDN U54021 ( .A(n44693), .B(n44692), .Z(n44688) );
  IV U54022 ( .A(n44694), .Z(n44693) );
  NAND U54023 ( .A(n44695), .B(n44696), .Z(n44650) );
  NANDN U54024 ( .A(n44697), .B(n44698), .Z(n44696) );
  NANDN U54025 ( .A(n44699), .B(n44700), .Z(n44698) );
  NANDN U54026 ( .A(n44700), .B(n44699), .Z(n44695) );
  IV U54027 ( .A(n44701), .Z(n44699) );
  XOR U54028 ( .A(n44676), .B(n44702), .Z(N61412) );
  XNOR U54029 ( .A(n44679), .B(n44678), .Z(n44702) );
  XNOR U54030 ( .A(n44690), .B(n44703), .Z(n44678) );
  XNOR U54031 ( .A(n44694), .B(n44692), .Z(n44703) );
  XOR U54032 ( .A(n44700), .B(n44704), .Z(n44692) );
  XNOR U54033 ( .A(n44697), .B(n44701), .Z(n44704) );
  AND U54034 ( .A(n44705), .B(n44706), .Z(n44701) );
  NAND U54035 ( .A(n44707), .B(n44708), .Z(n44706) );
  NAND U54036 ( .A(n44709), .B(n44710), .Z(n44705) );
  AND U54037 ( .A(n44711), .B(n44712), .Z(n44697) );
  NAND U54038 ( .A(n44713), .B(n44714), .Z(n44712) );
  NAND U54039 ( .A(n44715), .B(n44716), .Z(n44711) );
  NANDN U54040 ( .A(n44717), .B(n44718), .Z(n44700) );
  ANDN U54041 ( .B(n44719), .A(n44720), .Z(n44694) );
  XNOR U54042 ( .A(n44685), .B(n44721), .Z(n44690) );
  XNOR U54043 ( .A(n44683), .B(n44687), .Z(n44721) );
  AND U54044 ( .A(n44722), .B(n44723), .Z(n44687) );
  NAND U54045 ( .A(n44724), .B(n44725), .Z(n44723) );
  NAND U54046 ( .A(n44726), .B(n44727), .Z(n44722) );
  AND U54047 ( .A(n44728), .B(n44729), .Z(n44683) );
  NAND U54048 ( .A(n44730), .B(n44731), .Z(n44729) );
  NAND U54049 ( .A(n44732), .B(n44733), .Z(n44728) );
  AND U54050 ( .A(n44734), .B(n44735), .Z(n44685) );
  NAND U54051 ( .A(n44736), .B(n44737), .Z(n44679) );
  XNOR U54052 ( .A(n44662), .B(n44738), .Z(n44676) );
  XNOR U54053 ( .A(n44666), .B(n44664), .Z(n44738) );
  XOR U54054 ( .A(n44672), .B(n44739), .Z(n44664) );
  XNOR U54055 ( .A(n44669), .B(n44673), .Z(n44739) );
  AND U54056 ( .A(n44740), .B(n44741), .Z(n44673) );
  NAND U54057 ( .A(n44742), .B(n44743), .Z(n44741) );
  NAND U54058 ( .A(n44744), .B(n44745), .Z(n44740) );
  AND U54059 ( .A(n44746), .B(n44747), .Z(n44669) );
  NAND U54060 ( .A(n44748), .B(n44749), .Z(n44747) );
  NAND U54061 ( .A(n44750), .B(n44751), .Z(n44746) );
  NANDN U54062 ( .A(n44752), .B(n44753), .Z(n44672) );
  ANDN U54063 ( .B(n44754), .A(n44755), .Z(n44666) );
  XNOR U54064 ( .A(n44657), .B(n44756), .Z(n44662) );
  XNOR U54065 ( .A(n44655), .B(n44659), .Z(n44756) );
  AND U54066 ( .A(n44757), .B(n44758), .Z(n44659) );
  NAND U54067 ( .A(n44759), .B(n44760), .Z(n44758) );
  NAND U54068 ( .A(n44761), .B(n44762), .Z(n44757) );
  AND U54069 ( .A(n44763), .B(n44764), .Z(n44655) );
  NAND U54070 ( .A(n44765), .B(n44766), .Z(n44764) );
  NAND U54071 ( .A(n44767), .B(n44768), .Z(n44763) );
  AND U54072 ( .A(n44769), .B(n44770), .Z(n44657) );
  XOR U54073 ( .A(n44737), .B(n44736), .Z(N61411) );
  XNOR U54074 ( .A(n44754), .B(n44755), .Z(n44736) );
  XNOR U54075 ( .A(n44769), .B(n44770), .Z(n44755) );
  XOR U54076 ( .A(n44766), .B(n44765), .Z(n44770) );
  XOR U54077 ( .A(y[1524]), .B(x[1524]), .Z(n44765) );
  XOR U54078 ( .A(n44768), .B(n44767), .Z(n44766) );
  XOR U54079 ( .A(y[1526]), .B(x[1526]), .Z(n44767) );
  XOR U54080 ( .A(y[1525]), .B(x[1525]), .Z(n44768) );
  XOR U54081 ( .A(n44760), .B(n44759), .Z(n44769) );
  XOR U54082 ( .A(n44762), .B(n44761), .Z(n44759) );
  XOR U54083 ( .A(y[1523]), .B(x[1523]), .Z(n44761) );
  XOR U54084 ( .A(y[1522]), .B(x[1522]), .Z(n44762) );
  XOR U54085 ( .A(y[1521]), .B(x[1521]), .Z(n44760) );
  XNOR U54086 ( .A(n44753), .B(n44752), .Z(n44754) );
  XNOR U54087 ( .A(n44749), .B(n44748), .Z(n44752) );
  XOR U54088 ( .A(n44751), .B(n44750), .Z(n44748) );
  XOR U54089 ( .A(y[1520]), .B(x[1520]), .Z(n44750) );
  XOR U54090 ( .A(y[1519]), .B(x[1519]), .Z(n44751) );
  XOR U54091 ( .A(y[1518]), .B(x[1518]), .Z(n44749) );
  XOR U54092 ( .A(n44743), .B(n44742), .Z(n44753) );
  XOR U54093 ( .A(n44745), .B(n44744), .Z(n44742) );
  XOR U54094 ( .A(y[1517]), .B(x[1517]), .Z(n44744) );
  XOR U54095 ( .A(y[1516]), .B(x[1516]), .Z(n44745) );
  XOR U54096 ( .A(y[1515]), .B(x[1515]), .Z(n44743) );
  XNOR U54097 ( .A(n44719), .B(n44720), .Z(n44737) );
  XNOR U54098 ( .A(n44734), .B(n44735), .Z(n44720) );
  XOR U54099 ( .A(n44731), .B(n44730), .Z(n44735) );
  XOR U54100 ( .A(y[1512]), .B(x[1512]), .Z(n44730) );
  XOR U54101 ( .A(n44733), .B(n44732), .Z(n44731) );
  XOR U54102 ( .A(y[1514]), .B(x[1514]), .Z(n44732) );
  XOR U54103 ( .A(y[1513]), .B(x[1513]), .Z(n44733) );
  XOR U54104 ( .A(n44725), .B(n44724), .Z(n44734) );
  XOR U54105 ( .A(n44727), .B(n44726), .Z(n44724) );
  XOR U54106 ( .A(y[1511]), .B(x[1511]), .Z(n44726) );
  XOR U54107 ( .A(y[1510]), .B(x[1510]), .Z(n44727) );
  XOR U54108 ( .A(y[1509]), .B(x[1509]), .Z(n44725) );
  XNOR U54109 ( .A(n44718), .B(n44717), .Z(n44719) );
  XNOR U54110 ( .A(n44714), .B(n44713), .Z(n44717) );
  XOR U54111 ( .A(n44716), .B(n44715), .Z(n44713) );
  XOR U54112 ( .A(y[1508]), .B(x[1508]), .Z(n44715) );
  XOR U54113 ( .A(y[1507]), .B(x[1507]), .Z(n44716) );
  XOR U54114 ( .A(y[1506]), .B(x[1506]), .Z(n44714) );
  XOR U54115 ( .A(n44708), .B(n44707), .Z(n44718) );
  XOR U54116 ( .A(n44710), .B(n44709), .Z(n44707) );
  XOR U54117 ( .A(y[1505]), .B(x[1505]), .Z(n44709) );
  XOR U54118 ( .A(y[1504]), .B(x[1504]), .Z(n44710) );
  XOR U54119 ( .A(y[1503]), .B(x[1503]), .Z(n44708) );
  NAND U54120 ( .A(n44771), .B(n44772), .Z(N61402) );
  NAND U54121 ( .A(n44773), .B(n44774), .Z(n44772) );
  NANDN U54122 ( .A(n44775), .B(n44776), .Z(n44774) );
  NANDN U54123 ( .A(n44776), .B(n44775), .Z(n44771) );
  XOR U54124 ( .A(n44775), .B(n44777), .Z(N61401) );
  XNOR U54125 ( .A(n44773), .B(n44776), .Z(n44777) );
  NAND U54126 ( .A(n44778), .B(n44779), .Z(n44776) );
  NAND U54127 ( .A(n44780), .B(n44781), .Z(n44779) );
  NANDN U54128 ( .A(n44782), .B(n44783), .Z(n44781) );
  NANDN U54129 ( .A(n44783), .B(n44782), .Z(n44778) );
  AND U54130 ( .A(n44784), .B(n44785), .Z(n44773) );
  NAND U54131 ( .A(n44786), .B(n44787), .Z(n44785) );
  NANDN U54132 ( .A(n44788), .B(n44789), .Z(n44787) );
  NANDN U54133 ( .A(n44789), .B(n44788), .Z(n44784) );
  IV U54134 ( .A(n44790), .Z(n44789) );
  AND U54135 ( .A(n44791), .B(n44792), .Z(n44775) );
  NAND U54136 ( .A(n44793), .B(n44794), .Z(n44792) );
  NANDN U54137 ( .A(n44795), .B(n44796), .Z(n44794) );
  NANDN U54138 ( .A(n44796), .B(n44795), .Z(n44791) );
  XOR U54139 ( .A(n44788), .B(n44797), .Z(N61400) );
  XNOR U54140 ( .A(n44786), .B(n44790), .Z(n44797) );
  XOR U54141 ( .A(n44783), .B(n44798), .Z(n44790) );
  XNOR U54142 ( .A(n44780), .B(n44782), .Z(n44798) );
  AND U54143 ( .A(n44799), .B(n44800), .Z(n44782) );
  NANDN U54144 ( .A(n44801), .B(n44802), .Z(n44800) );
  OR U54145 ( .A(n44803), .B(n44804), .Z(n44802) );
  IV U54146 ( .A(n44805), .Z(n44804) );
  NANDN U54147 ( .A(n44805), .B(n44803), .Z(n44799) );
  AND U54148 ( .A(n44806), .B(n44807), .Z(n44780) );
  NAND U54149 ( .A(n44808), .B(n44809), .Z(n44807) );
  NANDN U54150 ( .A(n44810), .B(n44811), .Z(n44809) );
  NANDN U54151 ( .A(n44811), .B(n44810), .Z(n44806) );
  IV U54152 ( .A(n44812), .Z(n44811) );
  NAND U54153 ( .A(n44813), .B(n44814), .Z(n44783) );
  NANDN U54154 ( .A(n44815), .B(n44816), .Z(n44814) );
  NANDN U54155 ( .A(n44817), .B(n44818), .Z(n44816) );
  NANDN U54156 ( .A(n44818), .B(n44817), .Z(n44813) );
  IV U54157 ( .A(n44819), .Z(n44817) );
  AND U54158 ( .A(n44820), .B(n44821), .Z(n44786) );
  NAND U54159 ( .A(n44822), .B(n44823), .Z(n44821) );
  NANDN U54160 ( .A(n44824), .B(n44825), .Z(n44823) );
  NANDN U54161 ( .A(n44825), .B(n44824), .Z(n44820) );
  XOR U54162 ( .A(n44796), .B(n44826), .Z(n44788) );
  XNOR U54163 ( .A(n44793), .B(n44795), .Z(n44826) );
  AND U54164 ( .A(n44827), .B(n44828), .Z(n44795) );
  NANDN U54165 ( .A(n44829), .B(n44830), .Z(n44828) );
  OR U54166 ( .A(n44831), .B(n44832), .Z(n44830) );
  IV U54167 ( .A(n44833), .Z(n44832) );
  NANDN U54168 ( .A(n44833), .B(n44831), .Z(n44827) );
  AND U54169 ( .A(n44834), .B(n44835), .Z(n44793) );
  NAND U54170 ( .A(n44836), .B(n44837), .Z(n44835) );
  NANDN U54171 ( .A(n44838), .B(n44839), .Z(n44837) );
  NANDN U54172 ( .A(n44839), .B(n44838), .Z(n44834) );
  IV U54173 ( .A(n44840), .Z(n44839) );
  NAND U54174 ( .A(n44841), .B(n44842), .Z(n44796) );
  NANDN U54175 ( .A(n44843), .B(n44844), .Z(n44842) );
  NANDN U54176 ( .A(n44845), .B(n44846), .Z(n44844) );
  NANDN U54177 ( .A(n44846), .B(n44845), .Z(n44841) );
  IV U54178 ( .A(n44847), .Z(n44845) );
  XOR U54179 ( .A(n44822), .B(n44848), .Z(N61399) );
  XNOR U54180 ( .A(n44825), .B(n44824), .Z(n44848) );
  XNOR U54181 ( .A(n44836), .B(n44849), .Z(n44824) );
  XNOR U54182 ( .A(n44840), .B(n44838), .Z(n44849) );
  XOR U54183 ( .A(n44846), .B(n44850), .Z(n44838) );
  XNOR U54184 ( .A(n44843), .B(n44847), .Z(n44850) );
  AND U54185 ( .A(n44851), .B(n44852), .Z(n44847) );
  NAND U54186 ( .A(n44853), .B(n44854), .Z(n44852) );
  NAND U54187 ( .A(n44855), .B(n44856), .Z(n44851) );
  AND U54188 ( .A(n44857), .B(n44858), .Z(n44843) );
  NAND U54189 ( .A(n44859), .B(n44860), .Z(n44858) );
  NAND U54190 ( .A(n44861), .B(n44862), .Z(n44857) );
  NANDN U54191 ( .A(n44863), .B(n44864), .Z(n44846) );
  ANDN U54192 ( .B(n44865), .A(n44866), .Z(n44840) );
  XNOR U54193 ( .A(n44831), .B(n44867), .Z(n44836) );
  XNOR U54194 ( .A(n44829), .B(n44833), .Z(n44867) );
  AND U54195 ( .A(n44868), .B(n44869), .Z(n44833) );
  NAND U54196 ( .A(n44870), .B(n44871), .Z(n44869) );
  NAND U54197 ( .A(n44872), .B(n44873), .Z(n44868) );
  AND U54198 ( .A(n44874), .B(n44875), .Z(n44829) );
  NAND U54199 ( .A(n44876), .B(n44877), .Z(n44875) );
  NAND U54200 ( .A(n44878), .B(n44879), .Z(n44874) );
  AND U54201 ( .A(n44880), .B(n44881), .Z(n44831) );
  NAND U54202 ( .A(n44882), .B(n44883), .Z(n44825) );
  XNOR U54203 ( .A(n44808), .B(n44884), .Z(n44822) );
  XNOR U54204 ( .A(n44812), .B(n44810), .Z(n44884) );
  XOR U54205 ( .A(n44818), .B(n44885), .Z(n44810) );
  XNOR U54206 ( .A(n44815), .B(n44819), .Z(n44885) );
  AND U54207 ( .A(n44886), .B(n44887), .Z(n44819) );
  NAND U54208 ( .A(n44888), .B(n44889), .Z(n44887) );
  NAND U54209 ( .A(n44890), .B(n44891), .Z(n44886) );
  AND U54210 ( .A(n44892), .B(n44893), .Z(n44815) );
  NAND U54211 ( .A(n44894), .B(n44895), .Z(n44893) );
  NAND U54212 ( .A(n44896), .B(n44897), .Z(n44892) );
  NANDN U54213 ( .A(n44898), .B(n44899), .Z(n44818) );
  ANDN U54214 ( .B(n44900), .A(n44901), .Z(n44812) );
  XNOR U54215 ( .A(n44803), .B(n44902), .Z(n44808) );
  XNOR U54216 ( .A(n44801), .B(n44805), .Z(n44902) );
  AND U54217 ( .A(n44903), .B(n44904), .Z(n44805) );
  NAND U54218 ( .A(n44905), .B(n44906), .Z(n44904) );
  NAND U54219 ( .A(n44907), .B(n44908), .Z(n44903) );
  AND U54220 ( .A(n44909), .B(n44910), .Z(n44801) );
  NAND U54221 ( .A(n44911), .B(n44912), .Z(n44910) );
  NAND U54222 ( .A(n44913), .B(n44914), .Z(n44909) );
  AND U54223 ( .A(n44915), .B(n44916), .Z(n44803) );
  XOR U54224 ( .A(n44883), .B(n44882), .Z(N61398) );
  XNOR U54225 ( .A(n44900), .B(n44901), .Z(n44882) );
  XNOR U54226 ( .A(n44915), .B(n44916), .Z(n44901) );
  XOR U54227 ( .A(n44912), .B(n44911), .Z(n44916) );
  XOR U54228 ( .A(y[1500]), .B(x[1500]), .Z(n44911) );
  XOR U54229 ( .A(n44914), .B(n44913), .Z(n44912) );
  XOR U54230 ( .A(y[1502]), .B(x[1502]), .Z(n44913) );
  XOR U54231 ( .A(y[1501]), .B(x[1501]), .Z(n44914) );
  XOR U54232 ( .A(n44906), .B(n44905), .Z(n44915) );
  XOR U54233 ( .A(n44908), .B(n44907), .Z(n44905) );
  XOR U54234 ( .A(y[1499]), .B(x[1499]), .Z(n44907) );
  XOR U54235 ( .A(y[1498]), .B(x[1498]), .Z(n44908) );
  XOR U54236 ( .A(y[1497]), .B(x[1497]), .Z(n44906) );
  XNOR U54237 ( .A(n44899), .B(n44898), .Z(n44900) );
  XNOR U54238 ( .A(n44895), .B(n44894), .Z(n44898) );
  XOR U54239 ( .A(n44897), .B(n44896), .Z(n44894) );
  XOR U54240 ( .A(y[1496]), .B(x[1496]), .Z(n44896) );
  XOR U54241 ( .A(y[1495]), .B(x[1495]), .Z(n44897) );
  XOR U54242 ( .A(y[1494]), .B(x[1494]), .Z(n44895) );
  XOR U54243 ( .A(n44889), .B(n44888), .Z(n44899) );
  XOR U54244 ( .A(n44891), .B(n44890), .Z(n44888) );
  XOR U54245 ( .A(y[1493]), .B(x[1493]), .Z(n44890) );
  XOR U54246 ( .A(y[1492]), .B(x[1492]), .Z(n44891) );
  XOR U54247 ( .A(y[1491]), .B(x[1491]), .Z(n44889) );
  XNOR U54248 ( .A(n44865), .B(n44866), .Z(n44883) );
  XNOR U54249 ( .A(n44880), .B(n44881), .Z(n44866) );
  XOR U54250 ( .A(n44877), .B(n44876), .Z(n44881) );
  XOR U54251 ( .A(y[1488]), .B(x[1488]), .Z(n44876) );
  XOR U54252 ( .A(n44879), .B(n44878), .Z(n44877) );
  XOR U54253 ( .A(y[1490]), .B(x[1490]), .Z(n44878) );
  XOR U54254 ( .A(y[1489]), .B(x[1489]), .Z(n44879) );
  XOR U54255 ( .A(n44871), .B(n44870), .Z(n44880) );
  XOR U54256 ( .A(n44873), .B(n44872), .Z(n44870) );
  XOR U54257 ( .A(y[1487]), .B(x[1487]), .Z(n44872) );
  XOR U54258 ( .A(y[1486]), .B(x[1486]), .Z(n44873) );
  XOR U54259 ( .A(y[1485]), .B(x[1485]), .Z(n44871) );
  XNOR U54260 ( .A(n44864), .B(n44863), .Z(n44865) );
  XNOR U54261 ( .A(n44860), .B(n44859), .Z(n44863) );
  XOR U54262 ( .A(n44862), .B(n44861), .Z(n44859) );
  XOR U54263 ( .A(y[1484]), .B(x[1484]), .Z(n44861) );
  XOR U54264 ( .A(y[1483]), .B(x[1483]), .Z(n44862) );
  XOR U54265 ( .A(y[1482]), .B(x[1482]), .Z(n44860) );
  XOR U54266 ( .A(n44854), .B(n44853), .Z(n44864) );
  XOR U54267 ( .A(n44856), .B(n44855), .Z(n44853) );
  XOR U54268 ( .A(y[1481]), .B(x[1481]), .Z(n44855) );
  XOR U54269 ( .A(y[1480]), .B(x[1480]), .Z(n44856) );
  XOR U54270 ( .A(y[1479]), .B(x[1479]), .Z(n44854) );
  NAND U54271 ( .A(n44917), .B(n44918), .Z(N61389) );
  NAND U54272 ( .A(n44919), .B(n44920), .Z(n44918) );
  NANDN U54273 ( .A(n44921), .B(n44922), .Z(n44920) );
  NANDN U54274 ( .A(n44922), .B(n44921), .Z(n44917) );
  XOR U54275 ( .A(n44921), .B(n44923), .Z(N61388) );
  XNOR U54276 ( .A(n44919), .B(n44922), .Z(n44923) );
  NAND U54277 ( .A(n44924), .B(n44925), .Z(n44922) );
  NAND U54278 ( .A(n44926), .B(n44927), .Z(n44925) );
  NANDN U54279 ( .A(n44928), .B(n44929), .Z(n44927) );
  NANDN U54280 ( .A(n44929), .B(n44928), .Z(n44924) );
  AND U54281 ( .A(n44930), .B(n44931), .Z(n44919) );
  NAND U54282 ( .A(n44932), .B(n44933), .Z(n44931) );
  NANDN U54283 ( .A(n44934), .B(n44935), .Z(n44933) );
  NANDN U54284 ( .A(n44935), .B(n44934), .Z(n44930) );
  IV U54285 ( .A(n44936), .Z(n44935) );
  AND U54286 ( .A(n44937), .B(n44938), .Z(n44921) );
  NAND U54287 ( .A(n44939), .B(n44940), .Z(n44938) );
  NANDN U54288 ( .A(n44941), .B(n44942), .Z(n44940) );
  NANDN U54289 ( .A(n44942), .B(n44941), .Z(n44937) );
  XOR U54290 ( .A(n44934), .B(n44943), .Z(N61387) );
  XNOR U54291 ( .A(n44932), .B(n44936), .Z(n44943) );
  XOR U54292 ( .A(n44929), .B(n44944), .Z(n44936) );
  XNOR U54293 ( .A(n44926), .B(n44928), .Z(n44944) );
  AND U54294 ( .A(n44945), .B(n44946), .Z(n44928) );
  NANDN U54295 ( .A(n44947), .B(n44948), .Z(n44946) );
  OR U54296 ( .A(n44949), .B(n44950), .Z(n44948) );
  IV U54297 ( .A(n44951), .Z(n44950) );
  NANDN U54298 ( .A(n44951), .B(n44949), .Z(n44945) );
  AND U54299 ( .A(n44952), .B(n44953), .Z(n44926) );
  NAND U54300 ( .A(n44954), .B(n44955), .Z(n44953) );
  NANDN U54301 ( .A(n44956), .B(n44957), .Z(n44955) );
  NANDN U54302 ( .A(n44957), .B(n44956), .Z(n44952) );
  IV U54303 ( .A(n44958), .Z(n44957) );
  NAND U54304 ( .A(n44959), .B(n44960), .Z(n44929) );
  NANDN U54305 ( .A(n44961), .B(n44962), .Z(n44960) );
  NANDN U54306 ( .A(n44963), .B(n44964), .Z(n44962) );
  NANDN U54307 ( .A(n44964), .B(n44963), .Z(n44959) );
  IV U54308 ( .A(n44965), .Z(n44963) );
  AND U54309 ( .A(n44966), .B(n44967), .Z(n44932) );
  NAND U54310 ( .A(n44968), .B(n44969), .Z(n44967) );
  NANDN U54311 ( .A(n44970), .B(n44971), .Z(n44969) );
  NANDN U54312 ( .A(n44971), .B(n44970), .Z(n44966) );
  XOR U54313 ( .A(n44942), .B(n44972), .Z(n44934) );
  XNOR U54314 ( .A(n44939), .B(n44941), .Z(n44972) );
  AND U54315 ( .A(n44973), .B(n44974), .Z(n44941) );
  NANDN U54316 ( .A(n44975), .B(n44976), .Z(n44974) );
  OR U54317 ( .A(n44977), .B(n44978), .Z(n44976) );
  IV U54318 ( .A(n44979), .Z(n44978) );
  NANDN U54319 ( .A(n44979), .B(n44977), .Z(n44973) );
  AND U54320 ( .A(n44980), .B(n44981), .Z(n44939) );
  NAND U54321 ( .A(n44982), .B(n44983), .Z(n44981) );
  NANDN U54322 ( .A(n44984), .B(n44985), .Z(n44983) );
  NANDN U54323 ( .A(n44985), .B(n44984), .Z(n44980) );
  IV U54324 ( .A(n44986), .Z(n44985) );
  NAND U54325 ( .A(n44987), .B(n44988), .Z(n44942) );
  NANDN U54326 ( .A(n44989), .B(n44990), .Z(n44988) );
  NANDN U54327 ( .A(n44991), .B(n44992), .Z(n44990) );
  NANDN U54328 ( .A(n44992), .B(n44991), .Z(n44987) );
  IV U54329 ( .A(n44993), .Z(n44991) );
  XOR U54330 ( .A(n44968), .B(n44994), .Z(N61386) );
  XNOR U54331 ( .A(n44971), .B(n44970), .Z(n44994) );
  XNOR U54332 ( .A(n44982), .B(n44995), .Z(n44970) );
  XNOR U54333 ( .A(n44986), .B(n44984), .Z(n44995) );
  XOR U54334 ( .A(n44992), .B(n44996), .Z(n44984) );
  XNOR U54335 ( .A(n44989), .B(n44993), .Z(n44996) );
  AND U54336 ( .A(n44997), .B(n44998), .Z(n44993) );
  NAND U54337 ( .A(n44999), .B(n45000), .Z(n44998) );
  NAND U54338 ( .A(n45001), .B(n45002), .Z(n44997) );
  AND U54339 ( .A(n45003), .B(n45004), .Z(n44989) );
  NAND U54340 ( .A(n45005), .B(n45006), .Z(n45004) );
  NAND U54341 ( .A(n45007), .B(n45008), .Z(n45003) );
  NANDN U54342 ( .A(n45009), .B(n45010), .Z(n44992) );
  ANDN U54343 ( .B(n45011), .A(n45012), .Z(n44986) );
  XNOR U54344 ( .A(n44977), .B(n45013), .Z(n44982) );
  XNOR U54345 ( .A(n44975), .B(n44979), .Z(n45013) );
  AND U54346 ( .A(n45014), .B(n45015), .Z(n44979) );
  NAND U54347 ( .A(n45016), .B(n45017), .Z(n45015) );
  NAND U54348 ( .A(n45018), .B(n45019), .Z(n45014) );
  AND U54349 ( .A(n45020), .B(n45021), .Z(n44975) );
  NAND U54350 ( .A(n45022), .B(n45023), .Z(n45021) );
  NAND U54351 ( .A(n45024), .B(n45025), .Z(n45020) );
  AND U54352 ( .A(n45026), .B(n45027), .Z(n44977) );
  NAND U54353 ( .A(n45028), .B(n45029), .Z(n44971) );
  XNOR U54354 ( .A(n44954), .B(n45030), .Z(n44968) );
  XNOR U54355 ( .A(n44958), .B(n44956), .Z(n45030) );
  XOR U54356 ( .A(n44964), .B(n45031), .Z(n44956) );
  XNOR U54357 ( .A(n44961), .B(n44965), .Z(n45031) );
  AND U54358 ( .A(n45032), .B(n45033), .Z(n44965) );
  NAND U54359 ( .A(n45034), .B(n45035), .Z(n45033) );
  NAND U54360 ( .A(n45036), .B(n45037), .Z(n45032) );
  AND U54361 ( .A(n45038), .B(n45039), .Z(n44961) );
  NAND U54362 ( .A(n45040), .B(n45041), .Z(n45039) );
  NAND U54363 ( .A(n45042), .B(n45043), .Z(n45038) );
  NANDN U54364 ( .A(n45044), .B(n45045), .Z(n44964) );
  ANDN U54365 ( .B(n45046), .A(n45047), .Z(n44958) );
  XNOR U54366 ( .A(n44949), .B(n45048), .Z(n44954) );
  XNOR U54367 ( .A(n44947), .B(n44951), .Z(n45048) );
  AND U54368 ( .A(n45049), .B(n45050), .Z(n44951) );
  NAND U54369 ( .A(n45051), .B(n45052), .Z(n45050) );
  NAND U54370 ( .A(n45053), .B(n45054), .Z(n45049) );
  AND U54371 ( .A(n45055), .B(n45056), .Z(n44947) );
  NAND U54372 ( .A(n45057), .B(n45058), .Z(n45056) );
  NAND U54373 ( .A(n45059), .B(n45060), .Z(n45055) );
  AND U54374 ( .A(n45061), .B(n45062), .Z(n44949) );
  XOR U54375 ( .A(n45029), .B(n45028), .Z(N61385) );
  XNOR U54376 ( .A(n45046), .B(n45047), .Z(n45028) );
  XNOR U54377 ( .A(n45061), .B(n45062), .Z(n45047) );
  XOR U54378 ( .A(n45058), .B(n45057), .Z(n45062) );
  XOR U54379 ( .A(y[1476]), .B(x[1476]), .Z(n45057) );
  XOR U54380 ( .A(n45060), .B(n45059), .Z(n45058) );
  XOR U54381 ( .A(y[1478]), .B(x[1478]), .Z(n45059) );
  XOR U54382 ( .A(y[1477]), .B(x[1477]), .Z(n45060) );
  XOR U54383 ( .A(n45052), .B(n45051), .Z(n45061) );
  XOR U54384 ( .A(n45054), .B(n45053), .Z(n45051) );
  XOR U54385 ( .A(y[1475]), .B(x[1475]), .Z(n45053) );
  XOR U54386 ( .A(y[1474]), .B(x[1474]), .Z(n45054) );
  XOR U54387 ( .A(y[1473]), .B(x[1473]), .Z(n45052) );
  XNOR U54388 ( .A(n45045), .B(n45044), .Z(n45046) );
  XNOR U54389 ( .A(n45041), .B(n45040), .Z(n45044) );
  XOR U54390 ( .A(n45043), .B(n45042), .Z(n45040) );
  XOR U54391 ( .A(y[1472]), .B(x[1472]), .Z(n45042) );
  XOR U54392 ( .A(y[1471]), .B(x[1471]), .Z(n45043) );
  XOR U54393 ( .A(y[1470]), .B(x[1470]), .Z(n45041) );
  XOR U54394 ( .A(n45035), .B(n45034), .Z(n45045) );
  XOR U54395 ( .A(n45037), .B(n45036), .Z(n45034) );
  XOR U54396 ( .A(y[1469]), .B(x[1469]), .Z(n45036) );
  XOR U54397 ( .A(y[1468]), .B(x[1468]), .Z(n45037) );
  XOR U54398 ( .A(y[1467]), .B(x[1467]), .Z(n45035) );
  XNOR U54399 ( .A(n45011), .B(n45012), .Z(n45029) );
  XNOR U54400 ( .A(n45026), .B(n45027), .Z(n45012) );
  XOR U54401 ( .A(n45023), .B(n45022), .Z(n45027) );
  XOR U54402 ( .A(y[1464]), .B(x[1464]), .Z(n45022) );
  XOR U54403 ( .A(n45025), .B(n45024), .Z(n45023) );
  XOR U54404 ( .A(y[1466]), .B(x[1466]), .Z(n45024) );
  XOR U54405 ( .A(y[1465]), .B(x[1465]), .Z(n45025) );
  XOR U54406 ( .A(n45017), .B(n45016), .Z(n45026) );
  XOR U54407 ( .A(n45019), .B(n45018), .Z(n45016) );
  XOR U54408 ( .A(y[1463]), .B(x[1463]), .Z(n45018) );
  XOR U54409 ( .A(y[1462]), .B(x[1462]), .Z(n45019) );
  XOR U54410 ( .A(y[1461]), .B(x[1461]), .Z(n45017) );
  XNOR U54411 ( .A(n45010), .B(n45009), .Z(n45011) );
  XNOR U54412 ( .A(n45006), .B(n45005), .Z(n45009) );
  XOR U54413 ( .A(n45008), .B(n45007), .Z(n45005) );
  XOR U54414 ( .A(y[1460]), .B(x[1460]), .Z(n45007) );
  XOR U54415 ( .A(y[1459]), .B(x[1459]), .Z(n45008) );
  XOR U54416 ( .A(y[1458]), .B(x[1458]), .Z(n45006) );
  XOR U54417 ( .A(n45000), .B(n44999), .Z(n45010) );
  XOR U54418 ( .A(n45002), .B(n45001), .Z(n44999) );
  XOR U54419 ( .A(y[1457]), .B(x[1457]), .Z(n45001) );
  XOR U54420 ( .A(y[1456]), .B(x[1456]), .Z(n45002) );
  XOR U54421 ( .A(y[1455]), .B(x[1455]), .Z(n45000) );
  NAND U54422 ( .A(n45063), .B(n45064), .Z(N61376) );
  NAND U54423 ( .A(n45065), .B(n45066), .Z(n45064) );
  NANDN U54424 ( .A(n45067), .B(n45068), .Z(n45066) );
  NANDN U54425 ( .A(n45068), .B(n45067), .Z(n45063) );
  XOR U54426 ( .A(n45067), .B(n45069), .Z(N61375) );
  XNOR U54427 ( .A(n45065), .B(n45068), .Z(n45069) );
  NAND U54428 ( .A(n45070), .B(n45071), .Z(n45068) );
  NAND U54429 ( .A(n45072), .B(n45073), .Z(n45071) );
  NANDN U54430 ( .A(n45074), .B(n45075), .Z(n45073) );
  NANDN U54431 ( .A(n45075), .B(n45074), .Z(n45070) );
  AND U54432 ( .A(n45076), .B(n45077), .Z(n45065) );
  NAND U54433 ( .A(n45078), .B(n45079), .Z(n45077) );
  NANDN U54434 ( .A(n45080), .B(n45081), .Z(n45079) );
  NANDN U54435 ( .A(n45081), .B(n45080), .Z(n45076) );
  IV U54436 ( .A(n45082), .Z(n45081) );
  AND U54437 ( .A(n45083), .B(n45084), .Z(n45067) );
  NAND U54438 ( .A(n45085), .B(n45086), .Z(n45084) );
  NANDN U54439 ( .A(n45087), .B(n45088), .Z(n45086) );
  NANDN U54440 ( .A(n45088), .B(n45087), .Z(n45083) );
  XOR U54441 ( .A(n45080), .B(n45089), .Z(N61374) );
  XNOR U54442 ( .A(n45078), .B(n45082), .Z(n45089) );
  XOR U54443 ( .A(n45075), .B(n45090), .Z(n45082) );
  XNOR U54444 ( .A(n45072), .B(n45074), .Z(n45090) );
  AND U54445 ( .A(n45091), .B(n45092), .Z(n45074) );
  NANDN U54446 ( .A(n45093), .B(n45094), .Z(n45092) );
  OR U54447 ( .A(n45095), .B(n45096), .Z(n45094) );
  IV U54448 ( .A(n45097), .Z(n45096) );
  NANDN U54449 ( .A(n45097), .B(n45095), .Z(n45091) );
  AND U54450 ( .A(n45098), .B(n45099), .Z(n45072) );
  NAND U54451 ( .A(n45100), .B(n45101), .Z(n45099) );
  NANDN U54452 ( .A(n45102), .B(n45103), .Z(n45101) );
  NANDN U54453 ( .A(n45103), .B(n45102), .Z(n45098) );
  IV U54454 ( .A(n45104), .Z(n45103) );
  NAND U54455 ( .A(n45105), .B(n45106), .Z(n45075) );
  NANDN U54456 ( .A(n45107), .B(n45108), .Z(n45106) );
  NANDN U54457 ( .A(n45109), .B(n45110), .Z(n45108) );
  NANDN U54458 ( .A(n45110), .B(n45109), .Z(n45105) );
  IV U54459 ( .A(n45111), .Z(n45109) );
  AND U54460 ( .A(n45112), .B(n45113), .Z(n45078) );
  NAND U54461 ( .A(n45114), .B(n45115), .Z(n45113) );
  NANDN U54462 ( .A(n45116), .B(n45117), .Z(n45115) );
  NANDN U54463 ( .A(n45117), .B(n45116), .Z(n45112) );
  XOR U54464 ( .A(n45088), .B(n45118), .Z(n45080) );
  XNOR U54465 ( .A(n45085), .B(n45087), .Z(n45118) );
  AND U54466 ( .A(n45119), .B(n45120), .Z(n45087) );
  NANDN U54467 ( .A(n45121), .B(n45122), .Z(n45120) );
  OR U54468 ( .A(n45123), .B(n45124), .Z(n45122) );
  IV U54469 ( .A(n45125), .Z(n45124) );
  NANDN U54470 ( .A(n45125), .B(n45123), .Z(n45119) );
  AND U54471 ( .A(n45126), .B(n45127), .Z(n45085) );
  NAND U54472 ( .A(n45128), .B(n45129), .Z(n45127) );
  NANDN U54473 ( .A(n45130), .B(n45131), .Z(n45129) );
  NANDN U54474 ( .A(n45131), .B(n45130), .Z(n45126) );
  IV U54475 ( .A(n45132), .Z(n45131) );
  NAND U54476 ( .A(n45133), .B(n45134), .Z(n45088) );
  NANDN U54477 ( .A(n45135), .B(n45136), .Z(n45134) );
  NANDN U54478 ( .A(n45137), .B(n45138), .Z(n45136) );
  NANDN U54479 ( .A(n45138), .B(n45137), .Z(n45133) );
  IV U54480 ( .A(n45139), .Z(n45137) );
  XOR U54481 ( .A(n45114), .B(n45140), .Z(N61373) );
  XNOR U54482 ( .A(n45117), .B(n45116), .Z(n45140) );
  XNOR U54483 ( .A(n45128), .B(n45141), .Z(n45116) );
  XNOR U54484 ( .A(n45132), .B(n45130), .Z(n45141) );
  XOR U54485 ( .A(n45138), .B(n45142), .Z(n45130) );
  XNOR U54486 ( .A(n45135), .B(n45139), .Z(n45142) );
  AND U54487 ( .A(n45143), .B(n45144), .Z(n45139) );
  NAND U54488 ( .A(n45145), .B(n45146), .Z(n45144) );
  NAND U54489 ( .A(n45147), .B(n45148), .Z(n45143) );
  AND U54490 ( .A(n45149), .B(n45150), .Z(n45135) );
  NAND U54491 ( .A(n45151), .B(n45152), .Z(n45150) );
  NAND U54492 ( .A(n45153), .B(n45154), .Z(n45149) );
  NANDN U54493 ( .A(n45155), .B(n45156), .Z(n45138) );
  ANDN U54494 ( .B(n45157), .A(n45158), .Z(n45132) );
  XNOR U54495 ( .A(n45123), .B(n45159), .Z(n45128) );
  XNOR U54496 ( .A(n45121), .B(n45125), .Z(n45159) );
  AND U54497 ( .A(n45160), .B(n45161), .Z(n45125) );
  NAND U54498 ( .A(n45162), .B(n45163), .Z(n45161) );
  NAND U54499 ( .A(n45164), .B(n45165), .Z(n45160) );
  AND U54500 ( .A(n45166), .B(n45167), .Z(n45121) );
  NAND U54501 ( .A(n45168), .B(n45169), .Z(n45167) );
  NAND U54502 ( .A(n45170), .B(n45171), .Z(n45166) );
  AND U54503 ( .A(n45172), .B(n45173), .Z(n45123) );
  NAND U54504 ( .A(n45174), .B(n45175), .Z(n45117) );
  XNOR U54505 ( .A(n45100), .B(n45176), .Z(n45114) );
  XNOR U54506 ( .A(n45104), .B(n45102), .Z(n45176) );
  XOR U54507 ( .A(n45110), .B(n45177), .Z(n45102) );
  XNOR U54508 ( .A(n45107), .B(n45111), .Z(n45177) );
  AND U54509 ( .A(n45178), .B(n45179), .Z(n45111) );
  NAND U54510 ( .A(n45180), .B(n45181), .Z(n45179) );
  NAND U54511 ( .A(n45182), .B(n45183), .Z(n45178) );
  AND U54512 ( .A(n45184), .B(n45185), .Z(n45107) );
  NAND U54513 ( .A(n45186), .B(n45187), .Z(n45185) );
  NAND U54514 ( .A(n45188), .B(n45189), .Z(n45184) );
  NANDN U54515 ( .A(n45190), .B(n45191), .Z(n45110) );
  ANDN U54516 ( .B(n45192), .A(n45193), .Z(n45104) );
  XNOR U54517 ( .A(n45095), .B(n45194), .Z(n45100) );
  XNOR U54518 ( .A(n45093), .B(n45097), .Z(n45194) );
  AND U54519 ( .A(n45195), .B(n45196), .Z(n45097) );
  NAND U54520 ( .A(n45197), .B(n45198), .Z(n45196) );
  NAND U54521 ( .A(n45199), .B(n45200), .Z(n45195) );
  AND U54522 ( .A(n45201), .B(n45202), .Z(n45093) );
  NAND U54523 ( .A(n45203), .B(n45204), .Z(n45202) );
  NAND U54524 ( .A(n45205), .B(n45206), .Z(n45201) );
  AND U54525 ( .A(n45207), .B(n45208), .Z(n45095) );
  XOR U54526 ( .A(n45175), .B(n45174), .Z(N61372) );
  XNOR U54527 ( .A(n45192), .B(n45193), .Z(n45174) );
  XNOR U54528 ( .A(n45207), .B(n45208), .Z(n45193) );
  XOR U54529 ( .A(n45204), .B(n45203), .Z(n45208) );
  XOR U54530 ( .A(y[1452]), .B(x[1452]), .Z(n45203) );
  XOR U54531 ( .A(n45206), .B(n45205), .Z(n45204) );
  XOR U54532 ( .A(y[1454]), .B(x[1454]), .Z(n45205) );
  XOR U54533 ( .A(y[1453]), .B(x[1453]), .Z(n45206) );
  XOR U54534 ( .A(n45198), .B(n45197), .Z(n45207) );
  XOR U54535 ( .A(n45200), .B(n45199), .Z(n45197) );
  XOR U54536 ( .A(y[1451]), .B(x[1451]), .Z(n45199) );
  XOR U54537 ( .A(y[1450]), .B(x[1450]), .Z(n45200) );
  XOR U54538 ( .A(y[1449]), .B(x[1449]), .Z(n45198) );
  XNOR U54539 ( .A(n45191), .B(n45190), .Z(n45192) );
  XNOR U54540 ( .A(n45187), .B(n45186), .Z(n45190) );
  XOR U54541 ( .A(n45189), .B(n45188), .Z(n45186) );
  XOR U54542 ( .A(y[1448]), .B(x[1448]), .Z(n45188) );
  XOR U54543 ( .A(y[1447]), .B(x[1447]), .Z(n45189) );
  XOR U54544 ( .A(y[1446]), .B(x[1446]), .Z(n45187) );
  XOR U54545 ( .A(n45181), .B(n45180), .Z(n45191) );
  XOR U54546 ( .A(n45183), .B(n45182), .Z(n45180) );
  XOR U54547 ( .A(y[1445]), .B(x[1445]), .Z(n45182) );
  XOR U54548 ( .A(y[1444]), .B(x[1444]), .Z(n45183) );
  XOR U54549 ( .A(y[1443]), .B(x[1443]), .Z(n45181) );
  XNOR U54550 ( .A(n45157), .B(n45158), .Z(n45175) );
  XNOR U54551 ( .A(n45172), .B(n45173), .Z(n45158) );
  XOR U54552 ( .A(n45169), .B(n45168), .Z(n45173) );
  XOR U54553 ( .A(y[1440]), .B(x[1440]), .Z(n45168) );
  XOR U54554 ( .A(n45171), .B(n45170), .Z(n45169) );
  XOR U54555 ( .A(y[1442]), .B(x[1442]), .Z(n45170) );
  XOR U54556 ( .A(y[1441]), .B(x[1441]), .Z(n45171) );
  XOR U54557 ( .A(n45163), .B(n45162), .Z(n45172) );
  XOR U54558 ( .A(n45165), .B(n45164), .Z(n45162) );
  XOR U54559 ( .A(y[1439]), .B(x[1439]), .Z(n45164) );
  XOR U54560 ( .A(y[1438]), .B(x[1438]), .Z(n45165) );
  XOR U54561 ( .A(y[1437]), .B(x[1437]), .Z(n45163) );
  XNOR U54562 ( .A(n45156), .B(n45155), .Z(n45157) );
  XNOR U54563 ( .A(n45152), .B(n45151), .Z(n45155) );
  XOR U54564 ( .A(n45154), .B(n45153), .Z(n45151) );
  XOR U54565 ( .A(y[1436]), .B(x[1436]), .Z(n45153) );
  XOR U54566 ( .A(y[1435]), .B(x[1435]), .Z(n45154) );
  XOR U54567 ( .A(y[1434]), .B(x[1434]), .Z(n45152) );
  XOR U54568 ( .A(n45146), .B(n45145), .Z(n45156) );
  XOR U54569 ( .A(n45148), .B(n45147), .Z(n45145) );
  XOR U54570 ( .A(y[1433]), .B(x[1433]), .Z(n45147) );
  XOR U54571 ( .A(y[1432]), .B(x[1432]), .Z(n45148) );
  XOR U54572 ( .A(y[1431]), .B(x[1431]), .Z(n45146) );
  NAND U54573 ( .A(n45209), .B(n45210), .Z(N61363) );
  NAND U54574 ( .A(n45211), .B(n45212), .Z(n45210) );
  NANDN U54575 ( .A(n45213), .B(n45214), .Z(n45212) );
  NANDN U54576 ( .A(n45214), .B(n45213), .Z(n45209) );
  XOR U54577 ( .A(n45213), .B(n45215), .Z(N61362) );
  XNOR U54578 ( .A(n45211), .B(n45214), .Z(n45215) );
  NAND U54579 ( .A(n45216), .B(n45217), .Z(n45214) );
  NAND U54580 ( .A(n45218), .B(n45219), .Z(n45217) );
  NANDN U54581 ( .A(n45220), .B(n45221), .Z(n45219) );
  NANDN U54582 ( .A(n45221), .B(n45220), .Z(n45216) );
  AND U54583 ( .A(n45222), .B(n45223), .Z(n45211) );
  NAND U54584 ( .A(n45224), .B(n45225), .Z(n45223) );
  NANDN U54585 ( .A(n45226), .B(n45227), .Z(n45225) );
  NANDN U54586 ( .A(n45227), .B(n45226), .Z(n45222) );
  IV U54587 ( .A(n45228), .Z(n45227) );
  AND U54588 ( .A(n45229), .B(n45230), .Z(n45213) );
  NAND U54589 ( .A(n45231), .B(n45232), .Z(n45230) );
  NANDN U54590 ( .A(n45233), .B(n45234), .Z(n45232) );
  NANDN U54591 ( .A(n45234), .B(n45233), .Z(n45229) );
  XOR U54592 ( .A(n45226), .B(n45235), .Z(N61361) );
  XNOR U54593 ( .A(n45224), .B(n45228), .Z(n45235) );
  XOR U54594 ( .A(n45221), .B(n45236), .Z(n45228) );
  XNOR U54595 ( .A(n45218), .B(n45220), .Z(n45236) );
  AND U54596 ( .A(n45237), .B(n45238), .Z(n45220) );
  NANDN U54597 ( .A(n45239), .B(n45240), .Z(n45238) );
  OR U54598 ( .A(n45241), .B(n45242), .Z(n45240) );
  IV U54599 ( .A(n45243), .Z(n45242) );
  NANDN U54600 ( .A(n45243), .B(n45241), .Z(n45237) );
  AND U54601 ( .A(n45244), .B(n45245), .Z(n45218) );
  NAND U54602 ( .A(n45246), .B(n45247), .Z(n45245) );
  NANDN U54603 ( .A(n45248), .B(n45249), .Z(n45247) );
  NANDN U54604 ( .A(n45249), .B(n45248), .Z(n45244) );
  IV U54605 ( .A(n45250), .Z(n45249) );
  NAND U54606 ( .A(n45251), .B(n45252), .Z(n45221) );
  NANDN U54607 ( .A(n45253), .B(n45254), .Z(n45252) );
  NANDN U54608 ( .A(n45255), .B(n45256), .Z(n45254) );
  NANDN U54609 ( .A(n45256), .B(n45255), .Z(n45251) );
  IV U54610 ( .A(n45257), .Z(n45255) );
  AND U54611 ( .A(n45258), .B(n45259), .Z(n45224) );
  NAND U54612 ( .A(n45260), .B(n45261), .Z(n45259) );
  NANDN U54613 ( .A(n45262), .B(n45263), .Z(n45261) );
  NANDN U54614 ( .A(n45263), .B(n45262), .Z(n45258) );
  XOR U54615 ( .A(n45234), .B(n45264), .Z(n45226) );
  XNOR U54616 ( .A(n45231), .B(n45233), .Z(n45264) );
  AND U54617 ( .A(n45265), .B(n45266), .Z(n45233) );
  NANDN U54618 ( .A(n45267), .B(n45268), .Z(n45266) );
  OR U54619 ( .A(n45269), .B(n45270), .Z(n45268) );
  IV U54620 ( .A(n45271), .Z(n45270) );
  NANDN U54621 ( .A(n45271), .B(n45269), .Z(n45265) );
  AND U54622 ( .A(n45272), .B(n45273), .Z(n45231) );
  NAND U54623 ( .A(n45274), .B(n45275), .Z(n45273) );
  NANDN U54624 ( .A(n45276), .B(n45277), .Z(n45275) );
  NANDN U54625 ( .A(n45277), .B(n45276), .Z(n45272) );
  IV U54626 ( .A(n45278), .Z(n45277) );
  NAND U54627 ( .A(n45279), .B(n45280), .Z(n45234) );
  NANDN U54628 ( .A(n45281), .B(n45282), .Z(n45280) );
  NANDN U54629 ( .A(n45283), .B(n45284), .Z(n45282) );
  NANDN U54630 ( .A(n45284), .B(n45283), .Z(n45279) );
  IV U54631 ( .A(n45285), .Z(n45283) );
  XOR U54632 ( .A(n45260), .B(n45286), .Z(N61360) );
  XNOR U54633 ( .A(n45263), .B(n45262), .Z(n45286) );
  XNOR U54634 ( .A(n45274), .B(n45287), .Z(n45262) );
  XNOR U54635 ( .A(n45278), .B(n45276), .Z(n45287) );
  XOR U54636 ( .A(n45284), .B(n45288), .Z(n45276) );
  XNOR U54637 ( .A(n45281), .B(n45285), .Z(n45288) );
  AND U54638 ( .A(n45289), .B(n45290), .Z(n45285) );
  NAND U54639 ( .A(n45291), .B(n45292), .Z(n45290) );
  NAND U54640 ( .A(n45293), .B(n45294), .Z(n45289) );
  AND U54641 ( .A(n45295), .B(n45296), .Z(n45281) );
  NAND U54642 ( .A(n45297), .B(n45298), .Z(n45296) );
  NAND U54643 ( .A(n45299), .B(n45300), .Z(n45295) );
  NANDN U54644 ( .A(n45301), .B(n45302), .Z(n45284) );
  ANDN U54645 ( .B(n45303), .A(n45304), .Z(n45278) );
  XNOR U54646 ( .A(n45269), .B(n45305), .Z(n45274) );
  XNOR U54647 ( .A(n45267), .B(n45271), .Z(n45305) );
  AND U54648 ( .A(n45306), .B(n45307), .Z(n45271) );
  NAND U54649 ( .A(n45308), .B(n45309), .Z(n45307) );
  NAND U54650 ( .A(n45310), .B(n45311), .Z(n45306) );
  AND U54651 ( .A(n45312), .B(n45313), .Z(n45267) );
  NAND U54652 ( .A(n45314), .B(n45315), .Z(n45313) );
  NAND U54653 ( .A(n45316), .B(n45317), .Z(n45312) );
  AND U54654 ( .A(n45318), .B(n45319), .Z(n45269) );
  NAND U54655 ( .A(n45320), .B(n45321), .Z(n45263) );
  XNOR U54656 ( .A(n45246), .B(n45322), .Z(n45260) );
  XNOR U54657 ( .A(n45250), .B(n45248), .Z(n45322) );
  XOR U54658 ( .A(n45256), .B(n45323), .Z(n45248) );
  XNOR U54659 ( .A(n45253), .B(n45257), .Z(n45323) );
  AND U54660 ( .A(n45324), .B(n45325), .Z(n45257) );
  NAND U54661 ( .A(n45326), .B(n45327), .Z(n45325) );
  NAND U54662 ( .A(n45328), .B(n45329), .Z(n45324) );
  AND U54663 ( .A(n45330), .B(n45331), .Z(n45253) );
  NAND U54664 ( .A(n45332), .B(n45333), .Z(n45331) );
  NAND U54665 ( .A(n45334), .B(n45335), .Z(n45330) );
  NANDN U54666 ( .A(n45336), .B(n45337), .Z(n45256) );
  ANDN U54667 ( .B(n45338), .A(n45339), .Z(n45250) );
  XNOR U54668 ( .A(n45241), .B(n45340), .Z(n45246) );
  XNOR U54669 ( .A(n45239), .B(n45243), .Z(n45340) );
  AND U54670 ( .A(n45341), .B(n45342), .Z(n45243) );
  NAND U54671 ( .A(n45343), .B(n45344), .Z(n45342) );
  NAND U54672 ( .A(n45345), .B(n45346), .Z(n45341) );
  AND U54673 ( .A(n45347), .B(n45348), .Z(n45239) );
  NAND U54674 ( .A(n45349), .B(n45350), .Z(n45348) );
  NAND U54675 ( .A(n45351), .B(n45352), .Z(n45347) );
  AND U54676 ( .A(n45353), .B(n45354), .Z(n45241) );
  XOR U54677 ( .A(n45321), .B(n45320), .Z(N61359) );
  XNOR U54678 ( .A(n45338), .B(n45339), .Z(n45320) );
  XNOR U54679 ( .A(n45353), .B(n45354), .Z(n45339) );
  XOR U54680 ( .A(n45350), .B(n45349), .Z(n45354) );
  XOR U54681 ( .A(y[1428]), .B(x[1428]), .Z(n45349) );
  XOR U54682 ( .A(n45352), .B(n45351), .Z(n45350) );
  XOR U54683 ( .A(y[1430]), .B(x[1430]), .Z(n45351) );
  XOR U54684 ( .A(y[1429]), .B(x[1429]), .Z(n45352) );
  XOR U54685 ( .A(n45344), .B(n45343), .Z(n45353) );
  XOR U54686 ( .A(n45346), .B(n45345), .Z(n45343) );
  XOR U54687 ( .A(y[1427]), .B(x[1427]), .Z(n45345) );
  XOR U54688 ( .A(y[1426]), .B(x[1426]), .Z(n45346) );
  XOR U54689 ( .A(y[1425]), .B(x[1425]), .Z(n45344) );
  XNOR U54690 ( .A(n45337), .B(n45336), .Z(n45338) );
  XNOR U54691 ( .A(n45333), .B(n45332), .Z(n45336) );
  XOR U54692 ( .A(n45335), .B(n45334), .Z(n45332) );
  XOR U54693 ( .A(y[1424]), .B(x[1424]), .Z(n45334) );
  XOR U54694 ( .A(y[1423]), .B(x[1423]), .Z(n45335) );
  XOR U54695 ( .A(y[1422]), .B(x[1422]), .Z(n45333) );
  XOR U54696 ( .A(n45327), .B(n45326), .Z(n45337) );
  XOR U54697 ( .A(n45329), .B(n45328), .Z(n45326) );
  XOR U54698 ( .A(y[1421]), .B(x[1421]), .Z(n45328) );
  XOR U54699 ( .A(y[1420]), .B(x[1420]), .Z(n45329) );
  XOR U54700 ( .A(y[1419]), .B(x[1419]), .Z(n45327) );
  XNOR U54701 ( .A(n45303), .B(n45304), .Z(n45321) );
  XNOR U54702 ( .A(n45318), .B(n45319), .Z(n45304) );
  XOR U54703 ( .A(n45315), .B(n45314), .Z(n45319) );
  XOR U54704 ( .A(y[1416]), .B(x[1416]), .Z(n45314) );
  XOR U54705 ( .A(n45317), .B(n45316), .Z(n45315) );
  XOR U54706 ( .A(y[1418]), .B(x[1418]), .Z(n45316) );
  XOR U54707 ( .A(y[1417]), .B(x[1417]), .Z(n45317) );
  XOR U54708 ( .A(n45309), .B(n45308), .Z(n45318) );
  XOR U54709 ( .A(n45311), .B(n45310), .Z(n45308) );
  XOR U54710 ( .A(y[1415]), .B(x[1415]), .Z(n45310) );
  XOR U54711 ( .A(y[1414]), .B(x[1414]), .Z(n45311) );
  XOR U54712 ( .A(y[1413]), .B(x[1413]), .Z(n45309) );
  XNOR U54713 ( .A(n45302), .B(n45301), .Z(n45303) );
  XNOR U54714 ( .A(n45298), .B(n45297), .Z(n45301) );
  XOR U54715 ( .A(n45300), .B(n45299), .Z(n45297) );
  XOR U54716 ( .A(y[1412]), .B(x[1412]), .Z(n45299) );
  XOR U54717 ( .A(y[1411]), .B(x[1411]), .Z(n45300) );
  XOR U54718 ( .A(y[1410]), .B(x[1410]), .Z(n45298) );
  XOR U54719 ( .A(n45292), .B(n45291), .Z(n45302) );
  XOR U54720 ( .A(n45294), .B(n45293), .Z(n45291) );
  XOR U54721 ( .A(y[1409]), .B(x[1409]), .Z(n45293) );
  XOR U54722 ( .A(y[1408]), .B(x[1408]), .Z(n45294) );
  XOR U54723 ( .A(y[1407]), .B(x[1407]), .Z(n45292) );
  NAND U54724 ( .A(n45355), .B(n45356), .Z(N61350) );
  NAND U54725 ( .A(n45357), .B(n45358), .Z(n45356) );
  NANDN U54726 ( .A(n45359), .B(n45360), .Z(n45358) );
  NANDN U54727 ( .A(n45360), .B(n45359), .Z(n45355) );
  XOR U54728 ( .A(n45359), .B(n45361), .Z(N61349) );
  XNOR U54729 ( .A(n45357), .B(n45360), .Z(n45361) );
  NAND U54730 ( .A(n45362), .B(n45363), .Z(n45360) );
  NAND U54731 ( .A(n45364), .B(n45365), .Z(n45363) );
  NANDN U54732 ( .A(n45366), .B(n45367), .Z(n45365) );
  NANDN U54733 ( .A(n45367), .B(n45366), .Z(n45362) );
  AND U54734 ( .A(n45368), .B(n45369), .Z(n45357) );
  NAND U54735 ( .A(n45370), .B(n45371), .Z(n45369) );
  NANDN U54736 ( .A(n45372), .B(n45373), .Z(n45371) );
  NANDN U54737 ( .A(n45373), .B(n45372), .Z(n45368) );
  IV U54738 ( .A(n45374), .Z(n45373) );
  AND U54739 ( .A(n45375), .B(n45376), .Z(n45359) );
  NAND U54740 ( .A(n45377), .B(n45378), .Z(n45376) );
  NANDN U54741 ( .A(n45379), .B(n45380), .Z(n45378) );
  NANDN U54742 ( .A(n45380), .B(n45379), .Z(n45375) );
  XOR U54743 ( .A(n45372), .B(n45381), .Z(N61348) );
  XNOR U54744 ( .A(n45370), .B(n45374), .Z(n45381) );
  XOR U54745 ( .A(n45367), .B(n45382), .Z(n45374) );
  XNOR U54746 ( .A(n45364), .B(n45366), .Z(n45382) );
  AND U54747 ( .A(n45383), .B(n45384), .Z(n45366) );
  NANDN U54748 ( .A(n45385), .B(n45386), .Z(n45384) );
  OR U54749 ( .A(n45387), .B(n45388), .Z(n45386) );
  IV U54750 ( .A(n45389), .Z(n45388) );
  NANDN U54751 ( .A(n45389), .B(n45387), .Z(n45383) );
  AND U54752 ( .A(n45390), .B(n45391), .Z(n45364) );
  NAND U54753 ( .A(n45392), .B(n45393), .Z(n45391) );
  NANDN U54754 ( .A(n45394), .B(n45395), .Z(n45393) );
  NANDN U54755 ( .A(n45395), .B(n45394), .Z(n45390) );
  IV U54756 ( .A(n45396), .Z(n45395) );
  NAND U54757 ( .A(n45397), .B(n45398), .Z(n45367) );
  NANDN U54758 ( .A(n45399), .B(n45400), .Z(n45398) );
  NANDN U54759 ( .A(n45401), .B(n45402), .Z(n45400) );
  NANDN U54760 ( .A(n45402), .B(n45401), .Z(n45397) );
  IV U54761 ( .A(n45403), .Z(n45401) );
  AND U54762 ( .A(n45404), .B(n45405), .Z(n45370) );
  NAND U54763 ( .A(n45406), .B(n45407), .Z(n45405) );
  NANDN U54764 ( .A(n45408), .B(n45409), .Z(n45407) );
  NANDN U54765 ( .A(n45409), .B(n45408), .Z(n45404) );
  XOR U54766 ( .A(n45380), .B(n45410), .Z(n45372) );
  XNOR U54767 ( .A(n45377), .B(n45379), .Z(n45410) );
  AND U54768 ( .A(n45411), .B(n45412), .Z(n45379) );
  NANDN U54769 ( .A(n45413), .B(n45414), .Z(n45412) );
  OR U54770 ( .A(n45415), .B(n45416), .Z(n45414) );
  IV U54771 ( .A(n45417), .Z(n45416) );
  NANDN U54772 ( .A(n45417), .B(n45415), .Z(n45411) );
  AND U54773 ( .A(n45418), .B(n45419), .Z(n45377) );
  NAND U54774 ( .A(n45420), .B(n45421), .Z(n45419) );
  NANDN U54775 ( .A(n45422), .B(n45423), .Z(n45421) );
  NANDN U54776 ( .A(n45423), .B(n45422), .Z(n45418) );
  IV U54777 ( .A(n45424), .Z(n45423) );
  NAND U54778 ( .A(n45425), .B(n45426), .Z(n45380) );
  NANDN U54779 ( .A(n45427), .B(n45428), .Z(n45426) );
  NANDN U54780 ( .A(n45429), .B(n45430), .Z(n45428) );
  NANDN U54781 ( .A(n45430), .B(n45429), .Z(n45425) );
  IV U54782 ( .A(n45431), .Z(n45429) );
  XOR U54783 ( .A(n45406), .B(n45432), .Z(N61347) );
  XNOR U54784 ( .A(n45409), .B(n45408), .Z(n45432) );
  XNOR U54785 ( .A(n45420), .B(n45433), .Z(n45408) );
  XNOR U54786 ( .A(n45424), .B(n45422), .Z(n45433) );
  XOR U54787 ( .A(n45430), .B(n45434), .Z(n45422) );
  XNOR U54788 ( .A(n45427), .B(n45431), .Z(n45434) );
  AND U54789 ( .A(n45435), .B(n45436), .Z(n45431) );
  NAND U54790 ( .A(n45437), .B(n45438), .Z(n45436) );
  NAND U54791 ( .A(n45439), .B(n45440), .Z(n45435) );
  AND U54792 ( .A(n45441), .B(n45442), .Z(n45427) );
  NAND U54793 ( .A(n45443), .B(n45444), .Z(n45442) );
  NAND U54794 ( .A(n45445), .B(n45446), .Z(n45441) );
  NANDN U54795 ( .A(n45447), .B(n45448), .Z(n45430) );
  ANDN U54796 ( .B(n45449), .A(n45450), .Z(n45424) );
  XNOR U54797 ( .A(n45415), .B(n45451), .Z(n45420) );
  XNOR U54798 ( .A(n45413), .B(n45417), .Z(n45451) );
  AND U54799 ( .A(n45452), .B(n45453), .Z(n45417) );
  NAND U54800 ( .A(n45454), .B(n45455), .Z(n45453) );
  NAND U54801 ( .A(n45456), .B(n45457), .Z(n45452) );
  AND U54802 ( .A(n45458), .B(n45459), .Z(n45413) );
  NAND U54803 ( .A(n45460), .B(n45461), .Z(n45459) );
  NAND U54804 ( .A(n45462), .B(n45463), .Z(n45458) );
  AND U54805 ( .A(n45464), .B(n45465), .Z(n45415) );
  NAND U54806 ( .A(n45466), .B(n45467), .Z(n45409) );
  XNOR U54807 ( .A(n45392), .B(n45468), .Z(n45406) );
  XNOR U54808 ( .A(n45396), .B(n45394), .Z(n45468) );
  XOR U54809 ( .A(n45402), .B(n45469), .Z(n45394) );
  XNOR U54810 ( .A(n45399), .B(n45403), .Z(n45469) );
  AND U54811 ( .A(n45470), .B(n45471), .Z(n45403) );
  NAND U54812 ( .A(n45472), .B(n45473), .Z(n45471) );
  NAND U54813 ( .A(n45474), .B(n45475), .Z(n45470) );
  AND U54814 ( .A(n45476), .B(n45477), .Z(n45399) );
  NAND U54815 ( .A(n45478), .B(n45479), .Z(n45477) );
  NAND U54816 ( .A(n45480), .B(n45481), .Z(n45476) );
  NANDN U54817 ( .A(n45482), .B(n45483), .Z(n45402) );
  ANDN U54818 ( .B(n45484), .A(n45485), .Z(n45396) );
  XNOR U54819 ( .A(n45387), .B(n45486), .Z(n45392) );
  XNOR U54820 ( .A(n45385), .B(n45389), .Z(n45486) );
  AND U54821 ( .A(n45487), .B(n45488), .Z(n45389) );
  NAND U54822 ( .A(n45489), .B(n45490), .Z(n45488) );
  NAND U54823 ( .A(n45491), .B(n45492), .Z(n45487) );
  AND U54824 ( .A(n45493), .B(n45494), .Z(n45385) );
  NAND U54825 ( .A(n45495), .B(n45496), .Z(n45494) );
  NAND U54826 ( .A(n45497), .B(n45498), .Z(n45493) );
  AND U54827 ( .A(n45499), .B(n45500), .Z(n45387) );
  XOR U54828 ( .A(n45467), .B(n45466), .Z(N61346) );
  XNOR U54829 ( .A(n45484), .B(n45485), .Z(n45466) );
  XNOR U54830 ( .A(n45499), .B(n45500), .Z(n45485) );
  XOR U54831 ( .A(n45496), .B(n45495), .Z(n45500) );
  XOR U54832 ( .A(y[1404]), .B(x[1404]), .Z(n45495) );
  XOR U54833 ( .A(n45498), .B(n45497), .Z(n45496) );
  XOR U54834 ( .A(y[1406]), .B(x[1406]), .Z(n45497) );
  XOR U54835 ( .A(y[1405]), .B(x[1405]), .Z(n45498) );
  XOR U54836 ( .A(n45490), .B(n45489), .Z(n45499) );
  XOR U54837 ( .A(n45492), .B(n45491), .Z(n45489) );
  XOR U54838 ( .A(y[1403]), .B(x[1403]), .Z(n45491) );
  XOR U54839 ( .A(y[1402]), .B(x[1402]), .Z(n45492) );
  XOR U54840 ( .A(y[1401]), .B(x[1401]), .Z(n45490) );
  XNOR U54841 ( .A(n45483), .B(n45482), .Z(n45484) );
  XNOR U54842 ( .A(n45479), .B(n45478), .Z(n45482) );
  XOR U54843 ( .A(n45481), .B(n45480), .Z(n45478) );
  XOR U54844 ( .A(y[1400]), .B(x[1400]), .Z(n45480) );
  XOR U54845 ( .A(y[1399]), .B(x[1399]), .Z(n45481) );
  XOR U54846 ( .A(y[1398]), .B(x[1398]), .Z(n45479) );
  XOR U54847 ( .A(n45473), .B(n45472), .Z(n45483) );
  XOR U54848 ( .A(n45475), .B(n45474), .Z(n45472) );
  XOR U54849 ( .A(y[1397]), .B(x[1397]), .Z(n45474) );
  XOR U54850 ( .A(y[1396]), .B(x[1396]), .Z(n45475) );
  XOR U54851 ( .A(y[1395]), .B(x[1395]), .Z(n45473) );
  XNOR U54852 ( .A(n45449), .B(n45450), .Z(n45467) );
  XNOR U54853 ( .A(n45464), .B(n45465), .Z(n45450) );
  XOR U54854 ( .A(n45461), .B(n45460), .Z(n45465) );
  XOR U54855 ( .A(y[1392]), .B(x[1392]), .Z(n45460) );
  XOR U54856 ( .A(n45463), .B(n45462), .Z(n45461) );
  XOR U54857 ( .A(y[1394]), .B(x[1394]), .Z(n45462) );
  XOR U54858 ( .A(y[1393]), .B(x[1393]), .Z(n45463) );
  XOR U54859 ( .A(n45455), .B(n45454), .Z(n45464) );
  XOR U54860 ( .A(n45457), .B(n45456), .Z(n45454) );
  XOR U54861 ( .A(y[1391]), .B(x[1391]), .Z(n45456) );
  XOR U54862 ( .A(y[1390]), .B(x[1390]), .Z(n45457) );
  XOR U54863 ( .A(y[1389]), .B(x[1389]), .Z(n45455) );
  XNOR U54864 ( .A(n45448), .B(n45447), .Z(n45449) );
  XNOR U54865 ( .A(n45444), .B(n45443), .Z(n45447) );
  XOR U54866 ( .A(n45446), .B(n45445), .Z(n45443) );
  XOR U54867 ( .A(y[1388]), .B(x[1388]), .Z(n45445) );
  XOR U54868 ( .A(y[1387]), .B(x[1387]), .Z(n45446) );
  XOR U54869 ( .A(y[1386]), .B(x[1386]), .Z(n45444) );
  XOR U54870 ( .A(n45438), .B(n45437), .Z(n45448) );
  XOR U54871 ( .A(n45440), .B(n45439), .Z(n45437) );
  XOR U54872 ( .A(y[1385]), .B(x[1385]), .Z(n45439) );
  XOR U54873 ( .A(y[1384]), .B(x[1384]), .Z(n45440) );
  XOR U54874 ( .A(y[1383]), .B(x[1383]), .Z(n45438) );
  NAND U54875 ( .A(n45501), .B(n45502), .Z(N61337) );
  NAND U54876 ( .A(n45503), .B(n45504), .Z(n45502) );
  NANDN U54877 ( .A(n45505), .B(n45506), .Z(n45504) );
  NANDN U54878 ( .A(n45506), .B(n45505), .Z(n45501) );
  XOR U54879 ( .A(n45505), .B(n45507), .Z(N61336) );
  XNOR U54880 ( .A(n45503), .B(n45506), .Z(n45507) );
  NAND U54881 ( .A(n45508), .B(n45509), .Z(n45506) );
  NAND U54882 ( .A(n45510), .B(n45511), .Z(n45509) );
  NANDN U54883 ( .A(n45512), .B(n45513), .Z(n45511) );
  NANDN U54884 ( .A(n45513), .B(n45512), .Z(n45508) );
  AND U54885 ( .A(n45514), .B(n45515), .Z(n45503) );
  NAND U54886 ( .A(n45516), .B(n45517), .Z(n45515) );
  NANDN U54887 ( .A(n45518), .B(n45519), .Z(n45517) );
  NANDN U54888 ( .A(n45519), .B(n45518), .Z(n45514) );
  IV U54889 ( .A(n45520), .Z(n45519) );
  AND U54890 ( .A(n45521), .B(n45522), .Z(n45505) );
  NAND U54891 ( .A(n45523), .B(n45524), .Z(n45522) );
  NANDN U54892 ( .A(n45525), .B(n45526), .Z(n45524) );
  NANDN U54893 ( .A(n45526), .B(n45525), .Z(n45521) );
  XOR U54894 ( .A(n45518), .B(n45527), .Z(N61335) );
  XNOR U54895 ( .A(n45516), .B(n45520), .Z(n45527) );
  XOR U54896 ( .A(n45513), .B(n45528), .Z(n45520) );
  XNOR U54897 ( .A(n45510), .B(n45512), .Z(n45528) );
  AND U54898 ( .A(n45529), .B(n45530), .Z(n45512) );
  NANDN U54899 ( .A(n45531), .B(n45532), .Z(n45530) );
  OR U54900 ( .A(n45533), .B(n45534), .Z(n45532) );
  IV U54901 ( .A(n45535), .Z(n45534) );
  NANDN U54902 ( .A(n45535), .B(n45533), .Z(n45529) );
  AND U54903 ( .A(n45536), .B(n45537), .Z(n45510) );
  NAND U54904 ( .A(n45538), .B(n45539), .Z(n45537) );
  NANDN U54905 ( .A(n45540), .B(n45541), .Z(n45539) );
  NANDN U54906 ( .A(n45541), .B(n45540), .Z(n45536) );
  IV U54907 ( .A(n45542), .Z(n45541) );
  NAND U54908 ( .A(n45543), .B(n45544), .Z(n45513) );
  NANDN U54909 ( .A(n45545), .B(n45546), .Z(n45544) );
  NANDN U54910 ( .A(n45547), .B(n45548), .Z(n45546) );
  NANDN U54911 ( .A(n45548), .B(n45547), .Z(n45543) );
  IV U54912 ( .A(n45549), .Z(n45547) );
  AND U54913 ( .A(n45550), .B(n45551), .Z(n45516) );
  NAND U54914 ( .A(n45552), .B(n45553), .Z(n45551) );
  NANDN U54915 ( .A(n45554), .B(n45555), .Z(n45553) );
  NANDN U54916 ( .A(n45555), .B(n45554), .Z(n45550) );
  XOR U54917 ( .A(n45526), .B(n45556), .Z(n45518) );
  XNOR U54918 ( .A(n45523), .B(n45525), .Z(n45556) );
  AND U54919 ( .A(n45557), .B(n45558), .Z(n45525) );
  NANDN U54920 ( .A(n45559), .B(n45560), .Z(n45558) );
  OR U54921 ( .A(n45561), .B(n45562), .Z(n45560) );
  IV U54922 ( .A(n45563), .Z(n45562) );
  NANDN U54923 ( .A(n45563), .B(n45561), .Z(n45557) );
  AND U54924 ( .A(n45564), .B(n45565), .Z(n45523) );
  NAND U54925 ( .A(n45566), .B(n45567), .Z(n45565) );
  NANDN U54926 ( .A(n45568), .B(n45569), .Z(n45567) );
  NANDN U54927 ( .A(n45569), .B(n45568), .Z(n45564) );
  IV U54928 ( .A(n45570), .Z(n45569) );
  NAND U54929 ( .A(n45571), .B(n45572), .Z(n45526) );
  NANDN U54930 ( .A(n45573), .B(n45574), .Z(n45572) );
  NANDN U54931 ( .A(n45575), .B(n45576), .Z(n45574) );
  NANDN U54932 ( .A(n45576), .B(n45575), .Z(n45571) );
  IV U54933 ( .A(n45577), .Z(n45575) );
  XOR U54934 ( .A(n45552), .B(n45578), .Z(N61334) );
  XNOR U54935 ( .A(n45555), .B(n45554), .Z(n45578) );
  XNOR U54936 ( .A(n45566), .B(n45579), .Z(n45554) );
  XNOR U54937 ( .A(n45570), .B(n45568), .Z(n45579) );
  XOR U54938 ( .A(n45576), .B(n45580), .Z(n45568) );
  XNOR U54939 ( .A(n45573), .B(n45577), .Z(n45580) );
  AND U54940 ( .A(n45581), .B(n45582), .Z(n45577) );
  NAND U54941 ( .A(n45583), .B(n45584), .Z(n45582) );
  NAND U54942 ( .A(n45585), .B(n45586), .Z(n45581) );
  AND U54943 ( .A(n45587), .B(n45588), .Z(n45573) );
  NAND U54944 ( .A(n45589), .B(n45590), .Z(n45588) );
  NAND U54945 ( .A(n45591), .B(n45592), .Z(n45587) );
  NANDN U54946 ( .A(n45593), .B(n45594), .Z(n45576) );
  ANDN U54947 ( .B(n45595), .A(n45596), .Z(n45570) );
  XNOR U54948 ( .A(n45561), .B(n45597), .Z(n45566) );
  XNOR U54949 ( .A(n45559), .B(n45563), .Z(n45597) );
  AND U54950 ( .A(n45598), .B(n45599), .Z(n45563) );
  NAND U54951 ( .A(n45600), .B(n45601), .Z(n45599) );
  NAND U54952 ( .A(n45602), .B(n45603), .Z(n45598) );
  AND U54953 ( .A(n45604), .B(n45605), .Z(n45559) );
  NAND U54954 ( .A(n45606), .B(n45607), .Z(n45605) );
  NAND U54955 ( .A(n45608), .B(n45609), .Z(n45604) );
  AND U54956 ( .A(n45610), .B(n45611), .Z(n45561) );
  NAND U54957 ( .A(n45612), .B(n45613), .Z(n45555) );
  XNOR U54958 ( .A(n45538), .B(n45614), .Z(n45552) );
  XNOR U54959 ( .A(n45542), .B(n45540), .Z(n45614) );
  XOR U54960 ( .A(n45548), .B(n45615), .Z(n45540) );
  XNOR U54961 ( .A(n45545), .B(n45549), .Z(n45615) );
  AND U54962 ( .A(n45616), .B(n45617), .Z(n45549) );
  NAND U54963 ( .A(n45618), .B(n45619), .Z(n45617) );
  NAND U54964 ( .A(n45620), .B(n45621), .Z(n45616) );
  AND U54965 ( .A(n45622), .B(n45623), .Z(n45545) );
  NAND U54966 ( .A(n45624), .B(n45625), .Z(n45623) );
  NAND U54967 ( .A(n45626), .B(n45627), .Z(n45622) );
  NANDN U54968 ( .A(n45628), .B(n45629), .Z(n45548) );
  ANDN U54969 ( .B(n45630), .A(n45631), .Z(n45542) );
  XNOR U54970 ( .A(n45533), .B(n45632), .Z(n45538) );
  XNOR U54971 ( .A(n45531), .B(n45535), .Z(n45632) );
  AND U54972 ( .A(n45633), .B(n45634), .Z(n45535) );
  NAND U54973 ( .A(n45635), .B(n45636), .Z(n45634) );
  NAND U54974 ( .A(n45637), .B(n45638), .Z(n45633) );
  AND U54975 ( .A(n45639), .B(n45640), .Z(n45531) );
  NAND U54976 ( .A(n45641), .B(n45642), .Z(n45640) );
  NAND U54977 ( .A(n45643), .B(n45644), .Z(n45639) );
  AND U54978 ( .A(n45645), .B(n45646), .Z(n45533) );
  XOR U54979 ( .A(n45613), .B(n45612), .Z(N61333) );
  XNOR U54980 ( .A(n45630), .B(n45631), .Z(n45612) );
  XNOR U54981 ( .A(n45645), .B(n45646), .Z(n45631) );
  XOR U54982 ( .A(n45642), .B(n45641), .Z(n45646) );
  XOR U54983 ( .A(y[1380]), .B(x[1380]), .Z(n45641) );
  XOR U54984 ( .A(n45644), .B(n45643), .Z(n45642) );
  XOR U54985 ( .A(y[1382]), .B(x[1382]), .Z(n45643) );
  XOR U54986 ( .A(y[1381]), .B(x[1381]), .Z(n45644) );
  XOR U54987 ( .A(n45636), .B(n45635), .Z(n45645) );
  XOR U54988 ( .A(n45638), .B(n45637), .Z(n45635) );
  XOR U54989 ( .A(y[1379]), .B(x[1379]), .Z(n45637) );
  XOR U54990 ( .A(y[1378]), .B(x[1378]), .Z(n45638) );
  XOR U54991 ( .A(y[1377]), .B(x[1377]), .Z(n45636) );
  XNOR U54992 ( .A(n45629), .B(n45628), .Z(n45630) );
  XNOR U54993 ( .A(n45625), .B(n45624), .Z(n45628) );
  XOR U54994 ( .A(n45627), .B(n45626), .Z(n45624) );
  XOR U54995 ( .A(y[1376]), .B(x[1376]), .Z(n45626) );
  XOR U54996 ( .A(y[1375]), .B(x[1375]), .Z(n45627) );
  XOR U54997 ( .A(y[1374]), .B(x[1374]), .Z(n45625) );
  XOR U54998 ( .A(n45619), .B(n45618), .Z(n45629) );
  XOR U54999 ( .A(n45621), .B(n45620), .Z(n45618) );
  XOR U55000 ( .A(y[1373]), .B(x[1373]), .Z(n45620) );
  XOR U55001 ( .A(y[1372]), .B(x[1372]), .Z(n45621) );
  XOR U55002 ( .A(y[1371]), .B(x[1371]), .Z(n45619) );
  XNOR U55003 ( .A(n45595), .B(n45596), .Z(n45613) );
  XNOR U55004 ( .A(n45610), .B(n45611), .Z(n45596) );
  XOR U55005 ( .A(n45607), .B(n45606), .Z(n45611) );
  XOR U55006 ( .A(y[1368]), .B(x[1368]), .Z(n45606) );
  XOR U55007 ( .A(n45609), .B(n45608), .Z(n45607) );
  XOR U55008 ( .A(y[1370]), .B(x[1370]), .Z(n45608) );
  XOR U55009 ( .A(y[1369]), .B(x[1369]), .Z(n45609) );
  XOR U55010 ( .A(n45601), .B(n45600), .Z(n45610) );
  XOR U55011 ( .A(n45603), .B(n45602), .Z(n45600) );
  XOR U55012 ( .A(y[1367]), .B(x[1367]), .Z(n45602) );
  XOR U55013 ( .A(y[1366]), .B(x[1366]), .Z(n45603) );
  XOR U55014 ( .A(y[1365]), .B(x[1365]), .Z(n45601) );
  XNOR U55015 ( .A(n45594), .B(n45593), .Z(n45595) );
  XNOR U55016 ( .A(n45590), .B(n45589), .Z(n45593) );
  XOR U55017 ( .A(n45592), .B(n45591), .Z(n45589) );
  XOR U55018 ( .A(y[1364]), .B(x[1364]), .Z(n45591) );
  XOR U55019 ( .A(y[1363]), .B(x[1363]), .Z(n45592) );
  XOR U55020 ( .A(y[1362]), .B(x[1362]), .Z(n45590) );
  XOR U55021 ( .A(n45584), .B(n45583), .Z(n45594) );
  XOR U55022 ( .A(n45586), .B(n45585), .Z(n45583) );
  XOR U55023 ( .A(y[1361]), .B(x[1361]), .Z(n45585) );
  XOR U55024 ( .A(y[1360]), .B(x[1360]), .Z(n45586) );
  XOR U55025 ( .A(y[1359]), .B(x[1359]), .Z(n45584) );
  NAND U55026 ( .A(n45647), .B(n45648), .Z(N61324) );
  NAND U55027 ( .A(n45649), .B(n45650), .Z(n45648) );
  NANDN U55028 ( .A(n45651), .B(n45652), .Z(n45650) );
  NANDN U55029 ( .A(n45652), .B(n45651), .Z(n45647) );
  XOR U55030 ( .A(n45651), .B(n45653), .Z(N61323) );
  XNOR U55031 ( .A(n45649), .B(n45652), .Z(n45653) );
  NAND U55032 ( .A(n45654), .B(n45655), .Z(n45652) );
  NAND U55033 ( .A(n45656), .B(n45657), .Z(n45655) );
  NANDN U55034 ( .A(n45658), .B(n45659), .Z(n45657) );
  NANDN U55035 ( .A(n45659), .B(n45658), .Z(n45654) );
  AND U55036 ( .A(n45660), .B(n45661), .Z(n45649) );
  NAND U55037 ( .A(n45662), .B(n45663), .Z(n45661) );
  NANDN U55038 ( .A(n45664), .B(n45665), .Z(n45663) );
  NANDN U55039 ( .A(n45665), .B(n45664), .Z(n45660) );
  IV U55040 ( .A(n45666), .Z(n45665) );
  AND U55041 ( .A(n45667), .B(n45668), .Z(n45651) );
  NAND U55042 ( .A(n45669), .B(n45670), .Z(n45668) );
  NANDN U55043 ( .A(n45671), .B(n45672), .Z(n45670) );
  NANDN U55044 ( .A(n45672), .B(n45671), .Z(n45667) );
  XOR U55045 ( .A(n45664), .B(n45673), .Z(N61322) );
  XNOR U55046 ( .A(n45662), .B(n45666), .Z(n45673) );
  XOR U55047 ( .A(n45659), .B(n45674), .Z(n45666) );
  XNOR U55048 ( .A(n45656), .B(n45658), .Z(n45674) );
  AND U55049 ( .A(n45675), .B(n45676), .Z(n45658) );
  NANDN U55050 ( .A(n45677), .B(n45678), .Z(n45676) );
  OR U55051 ( .A(n45679), .B(n45680), .Z(n45678) );
  IV U55052 ( .A(n45681), .Z(n45680) );
  NANDN U55053 ( .A(n45681), .B(n45679), .Z(n45675) );
  AND U55054 ( .A(n45682), .B(n45683), .Z(n45656) );
  NAND U55055 ( .A(n45684), .B(n45685), .Z(n45683) );
  NANDN U55056 ( .A(n45686), .B(n45687), .Z(n45685) );
  NANDN U55057 ( .A(n45687), .B(n45686), .Z(n45682) );
  IV U55058 ( .A(n45688), .Z(n45687) );
  NAND U55059 ( .A(n45689), .B(n45690), .Z(n45659) );
  NANDN U55060 ( .A(n45691), .B(n45692), .Z(n45690) );
  NANDN U55061 ( .A(n45693), .B(n45694), .Z(n45692) );
  NANDN U55062 ( .A(n45694), .B(n45693), .Z(n45689) );
  IV U55063 ( .A(n45695), .Z(n45693) );
  AND U55064 ( .A(n45696), .B(n45697), .Z(n45662) );
  NAND U55065 ( .A(n45698), .B(n45699), .Z(n45697) );
  NANDN U55066 ( .A(n45700), .B(n45701), .Z(n45699) );
  NANDN U55067 ( .A(n45701), .B(n45700), .Z(n45696) );
  XOR U55068 ( .A(n45672), .B(n45702), .Z(n45664) );
  XNOR U55069 ( .A(n45669), .B(n45671), .Z(n45702) );
  AND U55070 ( .A(n45703), .B(n45704), .Z(n45671) );
  NANDN U55071 ( .A(n45705), .B(n45706), .Z(n45704) );
  OR U55072 ( .A(n45707), .B(n45708), .Z(n45706) );
  IV U55073 ( .A(n45709), .Z(n45708) );
  NANDN U55074 ( .A(n45709), .B(n45707), .Z(n45703) );
  AND U55075 ( .A(n45710), .B(n45711), .Z(n45669) );
  NAND U55076 ( .A(n45712), .B(n45713), .Z(n45711) );
  NANDN U55077 ( .A(n45714), .B(n45715), .Z(n45713) );
  NANDN U55078 ( .A(n45715), .B(n45714), .Z(n45710) );
  IV U55079 ( .A(n45716), .Z(n45715) );
  NAND U55080 ( .A(n45717), .B(n45718), .Z(n45672) );
  NANDN U55081 ( .A(n45719), .B(n45720), .Z(n45718) );
  NANDN U55082 ( .A(n45721), .B(n45722), .Z(n45720) );
  NANDN U55083 ( .A(n45722), .B(n45721), .Z(n45717) );
  IV U55084 ( .A(n45723), .Z(n45721) );
  XOR U55085 ( .A(n45698), .B(n45724), .Z(N61321) );
  XNOR U55086 ( .A(n45701), .B(n45700), .Z(n45724) );
  XNOR U55087 ( .A(n45712), .B(n45725), .Z(n45700) );
  XNOR U55088 ( .A(n45716), .B(n45714), .Z(n45725) );
  XOR U55089 ( .A(n45722), .B(n45726), .Z(n45714) );
  XNOR U55090 ( .A(n45719), .B(n45723), .Z(n45726) );
  AND U55091 ( .A(n45727), .B(n45728), .Z(n45723) );
  NAND U55092 ( .A(n45729), .B(n45730), .Z(n45728) );
  NAND U55093 ( .A(n45731), .B(n45732), .Z(n45727) );
  AND U55094 ( .A(n45733), .B(n45734), .Z(n45719) );
  NAND U55095 ( .A(n45735), .B(n45736), .Z(n45734) );
  NAND U55096 ( .A(n45737), .B(n45738), .Z(n45733) );
  NANDN U55097 ( .A(n45739), .B(n45740), .Z(n45722) );
  ANDN U55098 ( .B(n45741), .A(n45742), .Z(n45716) );
  XNOR U55099 ( .A(n45707), .B(n45743), .Z(n45712) );
  XNOR U55100 ( .A(n45705), .B(n45709), .Z(n45743) );
  AND U55101 ( .A(n45744), .B(n45745), .Z(n45709) );
  NAND U55102 ( .A(n45746), .B(n45747), .Z(n45745) );
  NAND U55103 ( .A(n45748), .B(n45749), .Z(n45744) );
  AND U55104 ( .A(n45750), .B(n45751), .Z(n45705) );
  NAND U55105 ( .A(n45752), .B(n45753), .Z(n45751) );
  NAND U55106 ( .A(n45754), .B(n45755), .Z(n45750) );
  AND U55107 ( .A(n45756), .B(n45757), .Z(n45707) );
  NAND U55108 ( .A(n45758), .B(n45759), .Z(n45701) );
  XNOR U55109 ( .A(n45684), .B(n45760), .Z(n45698) );
  XNOR U55110 ( .A(n45688), .B(n45686), .Z(n45760) );
  XOR U55111 ( .A(n45694), .B(n45761), .Z(n45686) );
  XNOR U55112 ( .A(n45691), .B(n45695), .Z(n45761) );
  AND U55113 ( .A(n45762), .B(n45763), .Z(n45695) );
  NAND U55114 ( .A(n45764), .B(n45765), .Z(n45763) );
  NAND U55115 ( .A(n45766), .B(n45767), .Z(n45762) );
  AND U55116 ( .A(n45768), .B(n45769), .Z(n45691) );
  NAND U55117 ( .A(n45770), .B(n45771), .Z(n45769) );
  NAND U55118 ( .A(n45772), .B(n45773), .Z(n45768) );
  NANDN U55119 ( .A(n45774), .B(n45775), .Z(n45694) );
  ANDN U55120 ( .B(n45776), .A(n45777), .Z(n45688) );
  XNOR U55121 ( .A(n45679), .B(n45778), .Z(n45684) );
  XNOR U55122 ( .A(n45677), .B(n45681), .Z(n45778) );
  AND U55123 ( .A(n45779), .B(n45780), .Z(n45681) );
  NAND U55124 ( .A(n45781), .B(n45782), .Z(n45780) );
  NAND U55125 ( .A(n45783), .B(n45784), .Z(n45779) );
  AND U55126 ( .A(n45785), .B(n45786), .Z(n45677) );
  NAND U55127 ( .A(n45787), .B(n45788), .Z(n45786) );
  NAND U55128 ( .A(n45789), .B(n45790), .Z(n45785) );
  AND U55129 ( .A(n45791), .B(n45792), .Z(n45679) );
  XOR U55130 ( .A(n45759), .B(n45758), .Z(N61320) );
  XNOR U55131 ( .A(n45776), .B(n45777), .Z(n45758) );
  XNOR U55132 ( .A(n45791), .B(n45792), .Z(n45777) );
  XOR U55133 ( .A(n45788), .B(n45787), .Z(n45792) );
  XOR U55134 ( .A(y[1356]), .B(x[1356]), .Z(n45787) );
  XOR U55135 ( .A(n45790), .B(n45789), .Z(n45788) );
  XOR U55136 ( .A(y[1358]), .B(x[1358]), .Z(n45789) );
  XOR U55137 ( .A(y[1357]), .B(x[1357]), .Z(n45790) );
  XOR U55138 ( .A(n45782), .B(n45781), .Z(n45791) );
  XOR U55139 ( .A(n45784), .B(n45783), .Z(n45781) );
  XOR U55140 ( .A(y[1355]), .B(x[1355]), .Z(n45783) );
  XOR U55141 ( .A(y[1354]), .B(x[1354]), .Z(n45784) );
  XOR U55142 ( .A(y[1353]), .B(x[1353]), .Z(n45782) );
  XNOR U55143 ( .A(n45775), .B(n45774), .Z(n45776) );
  XNOR U55144 ( .A(n45771), .B(n45770), .Z(n45774) );
  XOR U55145 ( .A(n45773), .B(n45772), .Z(n45770) );
  XOR U55146 ( .A(y[1352]), .B(x[1352]), .Z(n45772) );
  XOR U55147 ( .A(y[1351]), .B(x[1351]), .Z(n45773) );
  XOR U55148 ( .A(y[1350]), .B(x[1350]), .Z(n45771) );
  XOR U55149 ( .A(n45765), .B(n45764), .Z(n45775) );
  XOR U55150 ( .A(n45767), .B(n45766), .Z(n45764) );
  XOR U55151 ( .A(y[1349]), .B(x[1349]), .Z(n45766) );
  XOR U55152 ( .A(y[1348]), .B(x[1348]), .Z(n45767) );
  XOR U55153 ( .A(y[1347]), .B(x[1347]), .Z(n45765) );
  XNOR U55154 ( .A(n45741), .B(n45742), .Z(n45759) );
  XNOR U55155 ( .A(n45756), .B(n45757), .Z(n45742) );
  XOR U55156 ( .A(n45753), .B(n45752), .Z(n45757) );
  XOR U55157 ( .A(y[1344]), .B(x[1344]), .Z(n45752) );
  XOR U55158 ( .A(n45755), .B(n45754), .Z(n45753) );
  XOR U55159 ( .A(y[1346]), .B(x[1346]), .Z(n45754) );
  XOR U55160 ( .A(y[1345]), .B(x[1345]), .Z(n45755) );
  XOR U55161 ( .A(n45747), .B(n45746), .Z(n45756) );
  XOR U55162 ( .A(n45749), .B(n45748), .Z(n45746) );
  XOR U55163 ( .A(y[1343]), .B(x[1343]), .Z(n45748) );
  XOR U55164 ( .A(y[1342]), .B(x[1342]), .Z(n45749) );
  XOR U55165 ( .A(y[1341]), .B(x[1341]), .Z(n45747) );
  XNOR U55166 ( .A(n45740), .B(n45739), .Z(n45741) );
  XNOR U55167 ( .A(n45736), .B(n45735), .Z(n45739) );
  XOR U55168 ( .A(n45738), .B(n45737), .Z(n45735) );
  XOR U55169 ( .A(y[1340]), .B(x[1340]), .Z(n45737) );
  XOR U55170 ( .A(y[1339]), .B(x[1339]), .Z(n45738) );
  XOR U55171 ( .A(y[1338]), .B(x[1338]), .Z(n45736) );
  XOR U55172 ( .A(n45730), .B(n45729), .Z(n45740) );
  XOR U55173 ( .A(n45732), .B(n45731), .Z(n45729) );
  XOR U55174 ( .A(y[1337]), .B(x[1337]), .Z(n45731) );
  XOR U55175 ( .A(y[1336]), .B(x[1336]), .Z(n45732) );
  XOR U55176 ( .A(y[1335]), .B(x[1335]), .Z(n45730) );
  NAND U55177 ( .A(n45793), .B(n45794), .Z(N61311) );
  NAND U55178 ( .A(n45795), .B(n45796), .Z(n45794) );
  NANDN U55179 ( .A(n45797), .B(n45798), .Z(n45796) );
  NANDN U55180 ( .A(n45798), .B(n45797), .Z(n45793) );
  XOR U55181 ( .A(n45797), .B(n45799), .Z(N61310) );
  XNOR U55182 ( .A(n45795), .B(n45798), .Z(n45799) );
  NAND U55183 ( .A(n45800), .B(n45801), .Z(n45798) );
  NAND U55184 ( .A(n45802), .B(n45803), .Z(n45801) );
  NANDN U55185 ( .A(n45804), .B(n45805), .Z(n45803) );
  NANDN U55186 ( .A(n45805), .B(n45804), .Z(n45800) );
  AND U55187 ( .A(n45806), .B(n45807), .Z(n45795) );
  NAND U55188 ( .A(n45808), .B(n45809), .Z(n45807) );
  NANDN U55189 ( .A(n45810), .B(n45811), .Z(n45809) );
  NANDN U55190 ( .A(n45811), .B(n45810), .Z(n45806) );
  IV U55191 ( .A(n45812), .Z(n45811) );
  AND U55192 ( .A(n45813), .B(n45814), .Z(n45797) );
  NAND U55193 ( .A(n45815), .B(n45816), .Z(n45814) );
  NANDN U55194 ( .A(n45817), .B(n45818), .Z(n45816) );
  NANDN U55195 ( .A(n45818), .B(n45817), .Z(n45813) );
  XOR U55196 ( .A(n45810), .B(n45819), .Z(N61309) );
  XNOR U55197 ( .A(n45808), .B(n45812), .Z(n45819) );
  XOR U55198 ( .A(n45805), .B(n45820), .Z(n45812) );
  XNOR U55199 ( .A(n45802), .B(n45804), .Z(n45820) );
  AND U55200 ( .A(n45821), .B(n45822), .Z(n45804) );
  NANDN U55201 ( .A(n45823), .B(n45824), .Z(n45822) );
  OR U55202 ( .A(n45825), .B(n45826), .Z(n45824) );
  IV U55203 ( .A(n45827), .Z(n45826) );
  NANDN U55204 ( .A(n45827), .B(n45825), .Z(n45821) );
  AND U55205 ( .A(n45828), .B(n45829), .Z(n45802) );
  NAND U55206 ( .A(n45830), .B(n45831), .Z(n45829) );
  NANDN U55207 ( .A(n45832), .B(n45833), .Z(n45831) );
  NANDN U55208 ( .A(n45833), .B(n45832), .Z(n45828) );
  IV U55209 ( .A(n45834), .Z(n45833) );
  NAND U55210 ( .A(n45835), .B(n45836), .Z(n45805) );
  NANDN U55211 ( .A(n45837), .B(n45838), .Z(n45836) );
  NANDN U55212 ( .A(n45839), .B(n45840), .Z(n45838) );
  NANDN U55213 ( .A(n45840), .B(n45839), .Z(n45835) );
  IV U55214 ( .A(n45841), .Z(n45839) );
  AND U55215 ( .A(n45842), .B(n45843), .Z(n45808) );
  NAND U55216 ( .A(n45844), .B(n45845), .Z(n45843) );
  NANDN U55217 ( .A(n45846), .B(n45847), .Z(n45845) );
  NANDN U55218 ( .A(n45847), .B(n45846), .Z(n45842) );
  XOR U55219 ( .A(n45818), .B(n45848), .Z(n45810) );
  XNOR U55220 ( .A(n45815), .B(n45817), .Z(n45848) );
  AND U55221 ( .A(n45849), .B(n45850), .Z(n45817) );
  NANDN U55222 ( .A(n45851), .B(n45852), .Z(n45850) );
  OR U55223 ( .A(n45853), .B(n45854), .Z(n45852) );
  IV U55224 ( .A(n45855), .Z(n45854) );
  NANDN U55225 ( .A(n45855), .B(n45853), .Z(n45849) );
  AND U55226 ( .A(n45856), .B(n45857), .Z(n45815) );
  NAND U55227 ( .A(n45858), .B(n45859), .Z(n45857) );
  NANDN U55228 ( .A(n45860), .B(n45861), .Z(n45859) );
  NANDN U55229 ( .A(n45861), .B(n45860), .Z(n45856) );
  IV U55230 ( .A(n45862), .Z(n45861) );
  NAND U55231 ( .A(n45863), .B(n45864), .Z(n45818) );
  NANDN U55232 ( .A(n45865), .B(n45866), .Z(n45864) );
  NANDN U55233 ( .A(n45867), .B(n45868), .Z(n45866) );
  NANDN U55234 ( .A(n45868), .B(n45867), .Z(n45863) );
  IV U55235 ( .A(n45869), .Z(n45867) );
  XOR U55236 ( .A(n45844), .B(n45870), .Z(N61308) );
  XNOR U55237 ( .A(n45847), .B(n45846), .Z(n45870) );
  XNOR U55238 ( .A(n45858), .B(n45871), .Z(n45846) );
  XNOR U55239 ( .A(n45862), .B(n45860), .Z(n45871) );
  XOR U55240 ( .A(n45868), .B(n45872), .Z(n45860) );
  XNOR U55241 ( .A(n45865), .B(n45869), .Z(n45872) );
  AND U55242 ( .A(n45873), .B(n45874), .Z(n45869) );
  NAND U55243 ( .A(n45875), .B(n45876), .Z(n45874) );
  NAND U55244 ( .A(n45877), .B(n45878), .Z(n45873) );
  AND U55245 ( .A(n45879), .B(n45880), .Z(n45865) );
  NAND U55246 ( .A(n45881), .B(n45882), .Z(n45880) );
  NAND U55247 ( .A(n45883), .B(n45884), .Z(n45879) );
  NANDN U55248 ( .A(n45885), .B(n45886), .Z(n45868) );
  ANDN U55249 ( .B(n45887), .A(n45888), .Z(n45862) );
  XNOR U55250 ( .A(n45853), .B(n45889), .Z(n45858) );
  XNOR U55251 ( .A(n45851), .B(n45855), .Z(n45889) );
  AND U55252 ( .A(n45890), .B(n45891), .Z(n45855) );
  NAND U55253 ( .A(n45892), .B(n45893), .Z(n45891) );
  NAND U55254 ( .A(n45894), .B(n45895), .Z(n45890) );
  AND U55255 ( .A(n45896), .B(n45897), .Z(n45851) );
  NAND U55256 ( .A(n45898), .B(n45899), .Z(n45897) );
  NAND U55257 ( .A(n45900), .B(n45901), .Z(n45896) );
  AND U55258 ( .A(n45902), .B(n45903), .Z(n45853) );
  NAND U55259 ( .A(n45904), .B(n45905), .Z(n45847) );
  XNOR U55260 ( .A(n45830), .B(n45906), .Z(n45844) );
  XNOR U55261 ( .A(n45834), .B(n45832), .Z(n45906) );
  XOR U55262 ( .A(n45840), .B(n45907), .Z(n45832) );
  XNOR U55263 ( .A(n45837), .B(n45841), .Z(n45907) );
  AND U55264 ( .A(n45908), .B(n45909), .Z(n45841) );
  NAND U55265 ( .A(n45910), .B(n45911), .Z(n45909) );
  NAND U55266 ( .A(n45912), .B(n45913), .Z(n45908) );
  AND U55267 ( .A(n45914), .B(n45915), .Z(n45837) );
  NAND U55268 ( .A(n45916), .B(n45917), .Z(n45915) );
  NAND U55269 ( .A(n45918), .B(n45919), .Z(n45914) );
  NANDN U55270 ( .A(n45920), .B(n45921), .Z(n45840) );
  ANDN U55271 ( .B(n45922), .A(n45923), .Z(n45834) );
  XNOR U55272 ( .A(n45825), .B(n45924), .Z(n45830) );
  XNOR U55273 ( .A(n45823), .B(n45827), .Z(n45924) );
  AND U55274 ( .A(n45925), .B(n45926), .Z(n45827) );
  NAND U55275 ( .A(n45927), .B(n45928), .Z(n45926) );
  NAND U55276 ( .A(n45929), .B(n45930), .Z(n45925) );
  AND U55277 ( .A(n45931), .B(n45932), .Z(n45823) );
  NAND U55278 ( .A(n45933), .B(n45934), .Z(n45932) );
  NAND U55279 ( .A(n45935), .B(n45936), .Z(n45931) );
  AND U55280 ( .A(n45937), .B(n45938), .Z(n45825) );
  XOR U55281 ( .A(n45905), .B(n45904), .Z(N61307) );
  XNOR U55282 ( .A(n45922), .B(n45923), .Z(n45904) );
  XNOR U55283 ( .A(n45937), .B(n45938), .Z(n45923) );
  XOR U55284 ( .A(n45934), .B(n45933), .Z(n45938) );
  XOR U55285 ( .A(y[1332]), .B(x[1332]), .Z(n45933) );
  XOR U55286 ( .A(n45936), .B(n45935), .Z(n45934) );
  XOR U55287 ( .A(y[1334]), .B(x[1334]), .Z(n45935) );
  XOR U55288 ( .A(y[1333]), .B(x[1333]), .Z(n45936) );
  XOR U55289 ( .A(n45928), .B(n45927), .Z(n45937) );
  XOR U55290 ( .A(n45930), .B(n45929), .Z(n45927) );
  XOR U55291 ( .A(y[1331]), .B(x[1331]), .Z(n45929) );
  XOR U55292 ( .A(y[1330]), .B(x[1330]), .Z(n45930) );
  XOR U55293 ( .A(y[1329]), .B(x[1329]), .Z(n45928) );
  XNOR U55294 ( .A(n45921), .B(n45920), .Z(n45922) );
  XNOR U55295 ( .A(n45917), .B(n45916), .Z(n45920) );
  XOR U55296 ( .A(n45919), .B(n45918), .Z(n45916) );
  XOR U55297 ( .A(y[1328]), .B(x[1328]), .Z(n45918) );
  XOR U55298 ( .A(y[1327]), .B(x[1327]), .Z(n45919) );
  XOR U55299 ( .A(y[1326]), .B(x[1326]), .Z(n45917) );
  XOR U55300 ( .A(n45911), .B(n45910), .Z(n45921) );
  XOR U55301 ( .A(n45913), .B(n45912), .Z(n45910) );
  XOR U55302 ( .A(y[1325]), .B(x[1325]), .Z(n45912) );
  XOR U55303 ( .A(y[1324]), .B(x[1324]), .Z(n45913) );
  XOR U55304 ( .A(y[1323]), .B(x[1323]), .Z(n45911) );
  XNOR U55305 ( .A(n45887), .B(n45888), .Z(n45905) );
  XNOR U55306 ( .A(n45902), .B(n45903), .Z(n45888) );
  XOR U55307 ( .A(n45899), .B(n45898), .Z(n45903) );
  XOR U55308 ( .A(y[1320]), .B(x[1320]), .Z(n45898) );
  XOR U55309 ( .A(n45901), .B(n45900), .Z(n45899) );
  XOR U55310 ( .A(y[1322]), .B(x[1322]), .Z(n45900) );
  XOR U55311 ( .A(y[1321]), .B(x[1321]), .Z(n45901) );
  XOR U55312 ( .A(n45893), .B(n45892), .Z(n45902) );
  XOR U55313 ( .A(n45895), .B(n45894), .Z(n45892) );
  XOR U55314 ( .A(y[1319]), .B(x[1319]), .Z(n45894) );
  XOR U55315 ( .A(y[1318]), .B(x[1318]), .Z(n45895) );
  XOR U55316 ( .A(y[1317]), .B(x[1317]), .Z(n45893) );
  XNOR U55317 ( .A(n45886), .B(n45885), .Z(n45887) );
  XNOR U55318 ( .A(n45882), .B(n45881), .Z(n45885) );
  XOR U55319 ( .A(n45884), .B(n45883), .Z(n45881) );
  XOR U55320 ( .A(y[1316]), .B(x[1316]), .Z(n45883) );
  XOR U55321 ( .A(y[1315]), .B(x[1315]), .Z(n45884) );
  XOR U55322 ( .A(y[1314]), .B(x[1314]), .Z(n45882) );
  XOR U55323 ( .A(n45876), .B(n45875), .Z(n45886) );
  XOR U55324 ( .A(n45878), .B(n45877), .Z(n45875) );
  XOR U55325 ( .A(y[1313]), .B(x[1313]), .Z(n45877) );
  XOR U55326 ( .A(y[1312]), .B(x[1312]), .Z(n45878) );
  XOR U55327 ( .A(y[1311]), .B(x[1311]), .Z(n45876) );
  NAND U55328 ( .A(n45939), .B(n45940), .Z(N61298) );
  NAND U55329 ( .A(n45941), .B(n45942), .Z(n45940) );
  NANDN U55330 ( .A(n45943), .B(n45944), .Z(n45942) );
  NANDN U55331 ( .A(n45944), .B(n45943), .Z(n45939) );
  XOR U55332 ( .A(n45943), .B(n45945), .Z(N61297) );
  XNOR U55333 ( .A(n45941), .B(n45944), .Z(n45945) );
  NAND U55334 ( .A(n45946), .B(n45947), .Z(n45944) );
  NAND U55335 ( .A(n45948), .B(n45949), .Z(n45947) );
  NANDN U55336 ( .A(n45950), .B(n45951), .Z(n45949) );
  NANDN U55337 ( .A(n45951), .B(n45950), .Z(n45946) );
  AND U55338 ( .A(n45952), .B(n45953), .Z(n45941) );
  NAND U55339 ( .A(n45954), .B(n45955), .Z(n45953) );
  NANDN U55340 ( .A(n45956), .B(n45957), .Z(n45955) );
  NANDN U55341 ( .A(n45957), .B(n45956), .Z(n45952) );
  IV U55342 ( .A(n45958), .Z(n45957) );
  AND U55343 ( .A(n45959), .B(n45960), .Z(n45943) );
  NAND U55344 ( .A(n45961), .B(n45962), .Z(n45960) );
  NANDN U55345 ( .A(n45963), .B(n45964), .Z(n45962) );
  NANDN U55346 ( .A(n45964), .B(n45963), .Z(n45959) );
  XOR U55347 ( .A(n45956), .B(n45965), .Z(N61296) );
  XNOR U55348 ( .A(n45954), .B(n45958), .Z(n45965) );
  XOR U55349 ( .A(n45951), .B(n45966), .Z(n45958) );
  XNOR U55350 ( .A(n45948), .B(n45950), .Z(n45966) );
  AND U55351 ( .A(n45967), .B(n45968), .Z(n45950) );
  NANDN U55352 ( .A(n45969), .B(n45970), .Z(n45968) );
  OR U55353 ( .A(n45971), .B(n45972), .Z(n45970) );
  IV U55354 ( .A(n45973), .Z(n45972) );
  NANDN U55355 ( .A(n45973), .B(n45971), .Z(n45967) );
  AND U55356 ( .A(n45974), .B(n45975), .Z(n45948) );
  NAND U55357 ( .A(n45976), .B(n45977), .Z(n45975) );
  NANDN U55358 ( .A(n45978), .B(n45979), .Z(n45977) );
  NANDN U55359 ( .A(n45979), .B(n45978), .Z(n45974) );
  IV U55360 ( .A(n45980), .Z(n45979) );
  NAND U55361 ( .A(n45981), .B(n45982), .Z(n45951) );
  NANDN U55362 ( .A(n45983), .B(n45984), .Z(n45982) );
  NANDN U55363 ( .A(n45985), .B(n45986), .Z(n45984) );
  NANDN U55364 ( .A(n45986), .B(n45985), .Z(n45981) );
  IV U55365 ( .A(n45987), .Z(n45985) );
  AND U55366 ( .A(n45988), .B(n45989), .Z(n45954) );
  NAND U55367 ( .A(n45990), .B(n45991), .Z(n45989) );
  NANDN U55368 ( .A(n45992), .B(n45993), .Z(n45991) );
  NANDN U55369 ( .A(n45993), .B(n45992), .Z(n45988) );
  XOR U55370 ( .A(n45964), .B(n45994), .Z(n45956) );
  XNOR U55371 ( .A(n45961), .B(n45963), .Z(n45994) );
  AND U55372 ( .A(n45995), .B(n45996), .Z(n45963) );
  NANDN U55373 ( .A(n45997), .B(n45998), .Z(n45996) );
  OR U55374 ( .A(n45999), .B(n46000), .Z(n45998) );
  IV U55375 ( .A(n46001), .Z(n46000) );
  NANDN U55376 ( .A(n46001), .B(n45999), .Z(n45995) );
  AND U55377 ( .A(n46002), .B(n46003), .Z(n45961) );
  NAND U55378 ( .A(n46004), .B(n46005), .Z(n46003) );
  NANDN U55379 ( .A(n46006), .B(n46007), .Z(n46005) );
  NANDN U55380 ( .A(n46007), .B(n46006), .Z(n46002) );
  IV U55381 ( .A(n46008), .Z(n46007) );
  NAND U55382 ( .A(n46009), .B(n46010), .Z(n45964) );
  NANDN U55383 ( .A(n46011), .B(n46012), .Z(n46010) );
  NANDN U55384 ( .A(n46013), .B(n46014), .Z(n46012) );
  NANDN U55385 ( .A(n46014), .B(n46013), .Z(n46009) );
  IV U55386 ( .A(n46015), .Z(n46013) );
  XOR U55387 ( .A(n45990), .B(n46016), .Z(N61295) );
  XNOR U55388 ( .A(n45993), .B(n45992), .Z(n46016) );
  XNOR U55389 ( .A(n46004), .B(n46017), .Z(n45992) );
  XNOR U55390 ( .A(n46008), .B(n46006), .Z(n46017) );
  XOR U55391 ( .A(n46014), .B(n46018), .Z(n46006) );
  XNOR U55392 ( .A(n46011), .B(n46015), .Z(n46018) );
  AND U55393 ( .A(n46019), .B(n46020), .Z(n46015) );
  NAND U55394 ( .A(n46021), .B(n46022), .Z(n46020) );
  NAND U55395 ( .A(n46023), .B(n46024), .Z(n46019) );
  AND U55396 ( .A(n46025), .B(n46026), .Z(n46011) );
  NAND U55397 ( .A(n46027), .B(n46028), .Z(n46026) );
  NAND U55398 ( .A(n46029), .B(n46030), .Z(n46025) );
  NANDN U55399 ( .A(n46031), .B(n46032), .Z(n46014) );
  ANDN U55400 ( .B(n46033), .A(n46034), .Z(n46008) );
  XNOR U55401 ( .A(n45999), .B(n46035), .Z(n46004) );
  XNOR U55402 ( .A(n45997), .B(n46001), .Z(n46035) );
  AND U55403 ( .A(n46036), .B(n46037), .Z(n46001) );
  NAND U55404 ( .A(n46038), .B(n46039), .Z(n46037) );
  NAND U55405 ( .A(n46040), .B(n46041), .Z(n46036) );
  AND U55406 ( .A(n46042), .B(n46043), .Z(n45997) );
  NAND U55407 ( .A(n46044), .B(n46045), .Z(n46043) );
  NAND U55408 ( .A(n46046), .B(n46047), .Z(n46042) );
  AND U55409 ( .A(n46048), .B(n46049), .Z(n45999) );
  NAND U55410 ( .A(n46050), .B(n46051), .Z(n45993) );
  XNOR U55411 ( .A(n45976), .B(n46052), .Z(n45990) );
  XNOR U55412 ( .A(n45980), .B(n45978), .Z(n46052) );
  XOR U55413 ( .A(n45986), .B(n46053), .Z(n45978) );
  XNOR U55414 ( .A(n45983), .B(n45987), .Z(n46053) );
  AND U55415 ( .A(n46054), .B(n46055), .Z(n45987) );
  NAND U55416 ( .A(n46056), .B(n46057), .Z(n46055) );
  NAND U55417 ( .A(n46058), .B(n46059), .Z(n46054) );
  AND U55418 ( .A(n46060), .B(n46061), .Z(n45983) );
  NAND U55419 ( .A(n46062), .B(n46063), .Z(n46061) );
  NAND U55420 ( .A(n46064), .B(n46065), .Z(n46060) );
  NANDN U55421 ( .A(n46066), .B(n46067), .Z(n45986) );
  ANDN U55422 ( .B(n46068), .A(n46069), .Z(n45980) );
  XNOR U55423 ( .A(n45971), .B(n46070), .Z(n45976) );
  XNOR U55424 ( .A(n45969), .B(n45973), .Z(n46070) );
  AND U55425 ( .A(n46071), .B(n46072), .Z(n45973) );
  NAND U55426 ( .A(n46073), .B(n46074), .Z(n46072) );
  NAND U55427 ( .A(n46075), .B(n46076), .Z(n46071) );
  AND U55428 ( .A(n46077), .B(n46078), .Z(n45969) );
  NAND U55429 ( .A(n46079), .B(n46080), .Z(n46078) );
  NAND U55430 ( .A(n46081), .B(n46082), .Z(n46077) );
  AND U55431 ( .A(n46083), .B(n46084), .Z(n45971) );
  XOR U55432 ( .A(n46051), .B(n46050), .Z(N61294) );
  XNOR U55433 ( .A(n46068), .B(n46069), .Z(n46050) );
  XNOR U55434 ( .A(n46083), .B(n46084), .Z(n46069) );
  XOR U55435 ( .A(n46080), .B(n46079), .Z(n46084) );
  XOR U55436 ( .A(y[1308]), .B(x[1308]), .Z(n46079) );
  XOR U55437 ( .A(n46082), .B(n46081), .Z(n46080) );
  XOR U55438 ( .A(y[1310]), .B(x[1310]), .Z(n46081) );
  XOR U55439 ( .A(y[1309]), .B(x[1309]), .Z(n46082) );
  XOR U55440 ( .A(n46074), .B(n46073), .Z(n46083) );
  XOR U55441 ( .A(n46076), .B(n46075), .Z(n46073) );
  XOR U55442 ( .A(y[1307]), .B(x[1307]), .Z(n46075) );
  XOR U55443 ( .A(y[1306]), .B(x[1306]), .Z(n46076) );
  XOR U55444 ( .A(y[1305]), .B(x[1305]), .Z(n46074) );
  XNOR U55445 ( .A(n46067), .B(n46066), .Z(n46068) );
  XNOR U55446 ( .A(n46063), .B(n46062), .Z(n46066) );
  XOR U55447 ( .A(n46065), .B(n46064), .Z(n46062) );
  XOR U55448 ( .A(y[1304]), .B(x[1304]), .Z(n46064) );
  XOR U55449 ( .A(y[1303]), .B(x[1303]), .Z(n46065) );
  XOR U55450 ( .A(y[1302]), .B(x[1302]), .Z(n46063) );
  XOR U55451 ( .A(n46057), .B(n46056), .Z(n46067) );
  XOR U55452 ( .A(n46059), .B(n46058), .Z(n46056) );
  XOR U55453 ( .A(y[1301]), .B(x[1301]), .Z(n46058) );
  XOR U55454 ( .A(y[1300]), .B(x[1300]), .Z(n46059) );
  XOR U55455 ( .A(y[1299]), .B(x[1299]), .Z(n46057) );
  XNOR U55456 ( .A(n46033), .B(n46034), .Z(n46051) );
  XNOR U55457 ( .A(n46048), .B(n46049), .Z(n46034) );
  XOR U55458 ( .A(n46045), .B(n46044), .Z(n46049) );
  XOR U55459 ( .A(y[1296]), .B(x[1296]), .Z(n46044) );
  XOR U55460 ( .A(n46047), .B(n46046), .Z(n46045) );
  XOR U55461 ( .A(y[1298]), .B(x[1298]), .Z(n46046) );
  XOR U55462 ( .A(y[1297]), .B(x[1297]), .Z(n46047) );
  XOR U55463 ( .A(n46039), .B(n46038), .Z(n46048) );
  XOR U55464 ( .A(n46041), .B(n46040), .Z(n46038) );
  XOR U55465 ( .A(y[1295]), .B(x[1295]), .Z(n46040) );
  XOR U55466 ( .A(y[1294]), .B(x[1294]), .Z(n46041) );
  XOR U55467 ( .A(y[1293]), .B(x[1293]), .Z(n46039) );
  XNOR U55468 ( .A(n46032), .B(n46031), .Z(n46033) );
  XNOR U55469 ( .A(n46028), .B(n46027), .Z(n46031) );
  XOR U55470 ( .A(n46030), .B(n46029), .Z(n46027) );
  XOR U55471 ( .A(y[1292]), .B(x[1292]), .Z(n46029) );
  XOR U55472 ( .A(y[1291]), .B(x[1291]), .Z(n46030) );
  XOR U55473 ( .A(y[1290]), .B(x[1290]), .Z(n46028) );
  XOR U55474 ( .A(n46022), .B(n46021), .Z(n46032) );
  XOR U55475 ( .A(n46024), .B(n46023), .Z(n46021) );
  XOR U55476 ( .A(y[1289]), .B(x[1289]), .Z(n46023) );
  XOR U55477 ( .A(y[1288]), .B(x[1288]), .Z(n46024) );
  XOR U55478 ( .A(y[1287]), .B(x[1287]), .Z(n46022) );
  NAND U55479 ( .A(n46085), .B(n46086), .Z(N61285) );
  NAND U55480 ( .A(n46087), .B(n46088), .Z(n46086) );
  NANDN U55481 ( .A(n46089), .B(n46090), .Z(n46088) );
  NANDN U55482 ( .A(n46090), .B(n46089), .Z(n46085) );
  XOR U55483 ( .A(n46089), .B(n46091), .Z(N61284) );
  XNOR U55484 ( .A(n46087), .B(n46090), .Z(n46091) );
  NAND U55485 ( .A(n46092), .B(n46093), .Z(n46090) );
  NAND U55486 ( .A(n46094), .B(n46095), .Z(n46093) );
  NANDN U55487 ( .A(n46096), .B(n46097), .Z(n46095) );
  NANDN U55488 ( .A(n46097), .B(n46096), .Z(n46092) );
  AND U55489 ( .A(n46098), .B(n46099), .Z(n46087) );
  NAND U55490 ( .A(n46100), .B(n46101), .Z(n46099) );
  NANDN U55491 ( .A(n46102), .B(n46103), .Z(n46101) );
  NANDN U55492 ( .A(n46103), .B(n46102), .Z(n46098) );
  IV U55493 ( .A(n46104), .Z(n46103) );
  AND U55494 ( .A(n46105), .B(n46106), .Z(n46089) );
  NAND U55495 ( .A(n46107), .B(n46108), .Z(n46106) );
  NANDN U55496 ( .A(n46109), .B(n46110), .Z(n46108) );
  NANDN U55497 ( .A(n46110), .B(n46109), .Z(n46105) );
  XOR U55498 ( .A(n46102), .B(n46111), .Z(N61283) );
  XNOR U55499 ( .A(n46100), .B(n46104), .Z(n46111) );
  XOR U55500 ( .A(n46097), .B(n46112), .Z(n46104) );
  XNOR U55501 ( .A(n46094), .B(n46096), .Z(n46112) );
  AND U55502 ( .A(n46113), .B(n46114), .Z(n46096) );
  NANDN U55503 ( .A(n46115), .B(n46116), .Z(n46114) );
  OR U55504 ( .A(n46117), .B(n46118), .Z(n46116) );
  IV U55505 ( .A(n46119), .Z(n46118) );
  NANDN U55506 ( .A(n46119), .B(n46117), .Z(n46113) );
  AND U55507 ( .A(n46120), .B(n46121), .Z(n46094) );
  NAND U55508 ( .A(n46122), .B(n46123), .Z(n46121) );
  NANDN U55509 ( .A(n46124), .B(n46125), .Z(n46123) );
  NANDN U55510 ( .A(n46125), .B(n46124), .Z(n46120) );
  IV U55511 ( .A(n46126), .Z(n46125) );
  NAND U55512 ( .A(n46127), .B(n46128), .Z(n46097) );
  NANDN U55513 ( .A(n46129), .B(n46130), .Z(n46128) );
  NANDN U55514 ( .A(n46131), .B(n46132), .Z(n46130) );
  NANDN U55515 ( .A(n46132), .B(n46131), .Z(n46127) );
  IV U55516 ( .A(n46133), .Z(n46131) );
  AND U55517 ( .A(n46134), .B(n46135), .Z(n46100) );
  NAND U55518 ( .A(n46136), .B(n46137), .Z(n46135) );
  NANDN U55519 ( .A(n46138), .B(n46139), .Z(n46137) );
  NANDN U55520 ( .A(n46139), .B(n46138), .Z(n46134) );
  XOR U55521 ( .A(n46110), .B(n46140), .Z(n46102) );
  XNOR U55522 ( .A(n46107), .B(n46109), .Z(n46140) );
  AND U55523 ( .A(n46141), .B(n46142), .Z(n46109) );
  NANDN U55524 ( .A(n46143), .B(n46144), .Z(n46142) );
  OR U55525 ( .A(n46145), .B(n46146), .Z(n46144) );
  IV U55526 ( .A(n46147), .Z(n46146) );
  NANDN U55527 ( .A(n46147), .B(n46145), .Z(n46141) );
  AND U55528 ( .A(n46148), .B(n46149), .Z(n46107) );
  NAND U55529 ( .A(n46150), .B(n46151), .Z(n46149) );
  NANDN U55530 ( .A(n46152), .B(n46153), .Z(n46151) );
  NANDN U55531 ( .A(n46153), .B(n46152), .Z(n46148) );
  IV U55532 ( .A(n46154), .Z(n46153) );
  NAND U55533 ( .A(n46155), .B(n46156), .Z(n46110) );
  NANDN U55534 ( .A(n46157), .B(n46158), .Z(n46156) );
  NANDN U55535 ( .A(n46159), .B(n46160), .Z(n46158) );
  NANDN U55536 ( .A(n46160), .B(n46159), .Z(n46155) );
  IV U55537 ( .A(n46161), .Z(n46159) );
  XOR U55538 ( .A(n46136), .B(n46162), .Z(N61282) );
  XNOR U55539 ( .A(n46139), .B(n46138), .Z(n46162) );
  XNOR U55540 ( .A(n46150), .B(n46163), .Z(n46138) );
  XNOR U55541 ( .A(n46154), .B(n46152), .Z(n46163) );
  XOR U55542 ( .A(n46160), .B(n46164), .Z(n46152) );
  XNOR U55543 ( .A(n46157), .B(n46161), .Z(n46164) );
  AND U55544 ( .A(n46165), .B(n46166), .Z(n46161) );
  NAND U55545 ( .A(n46167), .B(n46168), .Z(n46166) );
  NAND U55546 ( .A(n46169), .B(n46170), .Z(n46165) );
  AND U55547 ( .A(n46171), .B(n46172), .Z(n46157) );
  NAND U55548 ( .A(n46173), .B(n46174), .Z(n46172) );
  NAND U55549 ( .A(n46175), .B(n46176), .Z(n46171) );
  NANDN U55550 ( .A(n46177), .B(n46178), .Z(n46160) );
  ANDN U55551 ( .B(n46179), .A(n46180), .Z(n46154) );
  XNOR U55552 ( .A(n46145), .B(n46181), .Z(n46150) );
  XNOR U55553 ( .A(n46143), .B(n46147), .Z(n46181) );
  AND U55554 ( .A(n46182), .B(n46183), .Z(n46147) );
  NAND U55555 ( .A(n46184), .B(n46185), .Z(n46183) );
  NAND U55556 ( .A(n46186), .B(n46187), .Z(n46182) );
  AND U55557 ( .A(n46188), .B(n46189), .Z(n46143) );
  NAND U55558 ( .A(n46190), .B(n46191), .Z(n46189) );
  NAND U55559 ( .A(n46192), .B(n46193), .Z(n46188) );
  AND U55560 ( .A(n46194), .B(n46195), .Z(n46145) );
  NAND U55561 ( .A(n46196), .B(n46197), .Z(n46139) );
  XNOR U55562 ( .A(n46122), .B(n46198), .Z(n46136) );
  XNOR U55563 ( .A(n46126), .B(n46124), .Z(n46198) );
  XOR U55564 ( .A(n46132), .B(n46199), .Z(n46124) );
  XNOR U55565 ( .A(n46129), .B(n46133), .Z(n46199) );
  AND U55566 ( .A(n46200), .B(n46201), .Z(n46133) );
  NAND U55567 ( .A(n46202), .B(n46203), .Z(n46201) );
  NAND U55568 ( .A(n46204), .B(n46205), .Z(n46200) );
  AND U55569 ( .A(n46206), .B(n46207), .Z(n46129) );
  NAND U55570 ( .A(n46208), .B(n46209), .Z(n46207) );
  NAND U55571 ( .A(n46210), .B(n46211), .Z(n46206) );
  NANDN U55572 ( .A(n46212), .B(n46213), .Z(n46132) );
  ANDN U55573 ( .B(n46214), .A(n46215), .Z(n46126) );
  XNOR U55574 ( .A(n46117), .B(n46216), .Z(n46122) );
  XNOR U55575 ( .A(n46115), .B(n46119), .Z(n46216) );
  AND U55576 ( .A(n46217), .B(n46218), .Z(n46119) );
  NAND U55577 ( .A(n46219), .B(n46220), .Z(n46218) );
  NAND U55578 ( .A(n46221), .B(n46222), .Z(n46217) );
  AND U55579 ( .A(n46223), .B(n46224), .Z(n46115) );
  NAND U55580 ( .A(n46225), .B(n46226), .Z(n46224) );
  NAND U55581 ( .A(n46227), .B(n46228), .Z(n46223) );
  AND U55582 ( .A(n46229), .B(n46230), .Z(n46117) );
  XOR U55583 ( .A(n46197), .B(n46196), .Z(N61281) );
  XNOR U55584 ( .A(n46214), .B(n46215), .Z(n46196) );
  XNOR U55585 ( .A(n46229), .B(n46230), .Z(n46215) );
  XOR U55586 ( .A(n46226), .B(n46225), .Z(n46230) );
  XOR U55587 ( .A(y[1284]), .B(x[1284]), .Z(n46225) );
  XOR U55588 ( .A(n46228), .B(n46227), .Z(n46226) );
  XOR U55589 ( .A(y[1286]), .B(x[1286]), .Z(n46227) );
  XOR U55590 ( .A(y[1285]), .B(x[1285]), .Z(n46228) );
  XOR U55591 ( .A(n46220), .B(n46219), .Z(n46229) );
  XOR U55592 ( .A(n46222), .B(n46221), .Z(n46219) );
  XOR U55593 ( .A(y[1283]), .B(x[1283]), .Z(n46221) );
  XOR U55594 ( .A(y[1282]), .B(x[1282]), .Z(n46222) );
  XOR U55595 ( .A(y[1281]), .B(x[1281]), .Z(n46220) );
  XNOR U55596 ( .A(n46213), .B(n46212), .Z(n46214) );
  XNOR U55597 ( .A(n46209), .B(n46208), .Z(n46212) );
  XOR U55598 ( .A(n46211), .B(n46210), .Z(n46208) );
  XOR U55599 ( .A(y[1280]), .B(x[1280]), .Z(n46210) );
  XOR U55600 ( .A(y[1279]), .B(x[1279]), .Z(n46211) );
  XOR U55601 ( .A(y[1278]), .B(x[1278]), .Z(n46209) );
  XOR U55602 ( .A(n46203), .B(n46202), .Z(n46213) );
  XOR U55603 ( .A(n46205), .B(n46204), .Z(n46202) );
  XOR U55604 ( .A(y[1277]), .B(x[1277]), .Z(n46204) );
  XOR U55605 ( .A(y[1276]), .B(x[1276]), .Z(n46205) );
  XOR U55606 ( .A(y[1275]), .B(x[1275]), .Z(n46203) );
  XNOR U55607 ( .A(n46179), .B(n46180), .Z(n46197) );
  XNOR U55608 ( .A(n46194), .B(n46195), .Z(n46180) );
  XOR U55609 ( .A(n46191), .B(n46190), .Z(n46195) );
  XOR U55610 ( .A(y[1272]), .B(x[1272]), .Z(n46190) );
  XOR U55611 ( .A(n46193), .B(n46192), .Z(n46191) );
  XOR U55612 ( .A(y[1274]), .B(x[1274]), .Z(n46192) );
  XOR U55613 ( .A(y[1273]), .B(x[1273]), .Z(n46193) );
  XOR U55614 ( .A(n46185), .B(n46184), .Z(n46194) );
  XOR U55615 ( .A(n46187), .B(n46186), .Z(n46184) );
  XOR U55616 ( .A(y[1271]), .B(x[1271]), .Z(n46186) );
  XOR U55617 ( .A(y[1270]), .B(x[1270]), .Z(n46187) );
  XOR U55618 ( .A(y[1269]), .B(x[1269]), .Z(n46185) );
  XNOR U55619 ( .A(n46178), .B(n46177), .Z(n46179) );
  XNOR U55620 ( .A(n46174), .B(n46173), .Z(n46177) );
  XOR U55621 ( .A(n46176), .B(n46175), .Z(n46173) );
  XOR U55622 ( .A(y[1268]), .B(x[1268]), .Z(n46175) );
  XOR U55623 ( .A(y[1267]), .B(x[1267]), .Z(n46176) );
  XOR U55624 ( .A(y[1266]), .B(x[1266]), .Z(n46174) );
  XOR U55625 ( .A(n46168), .B(n46167), .Z(n46178) );
  XOR U55626 ( .A(n46170), .B(n46169), .Z(n46167) );
  XOR U55627 ( .A(y[1265]), .B(x[1265]), .Z(n46169) );
  XOR U55628 ( .A(y[1264]), .B(x[1264]), .Z(n46170) );
  XOR U55629 ( .A(y[1263]), .B(x[1263]), .Z(n46168) );
  NAND U55630 ( .A(n46231), .B(n46232), .Z(N61272) );
  NAND U55631 ( .A(n46233), .B(n46234), .Z(n46232) );
  NANDN U55632 ( .A(n46235), .B(n46236), .Z(n46234) );
  NANDN U55633 ( .A(n46236), .B(n46235), .Z(n46231) );
  XOR U55634 ( .A(n46235), .B(n46237), .Z(N61271) );
  XNOR U55635 ( .A(n46233), .B(n46236), .Z(n46237) );
  NAND U55636 ( .A(n46238), .B(n46239), .Z(n46236) );
  NAND U55637 ( .A(n46240), .B(n46241), .Z(n46239) );
  NANDN U55638 ( .A(n46242), .B(n46243), .Z(n46241) );
  NANDN U55639 ( .A(n46243), .B(n46242), .Z(n46238) );
  AND U55640 ( .A(n46244), .B(n46245), .Z(n46233) );
  NAND U55641 ( .A(n46246), .B(n46247), .Z(n46245) );
  NANDN U55642 ( .A(n46248), .B(n46249), .Z(n46247) );
  NANDN U55643 ( .A(n46249), .B(n46248), .Z(n46244) );
  IV U55644 ( .A(n46250), .Z(n46249) );
  AND U55645 ( .A(n46251), .B(n46252), .Z(n46235) );
  NAND U55646 ( .A(n46253), .B(n46254), .Z(n46252) );
  NANDN U55647 ( .A(n46255), .B(n46256), .Z(n46254) );
  NANDN U55648 ( .A(n46256), .B(n46255), .Z(n46251) );
  XOR U55649 ( .A(n46248), .B(n46257), .Z(N61270) );
  XNOR U55650 ( .A(n46246), .B(n46250), .Z(n46257) );
  XOR U55651 ( .A(n46243), .B(n46258), .Z(n46250) );
  XNOR U55652 ( .A(n46240), .B(n46242), .Z(n46258) );
  AND U55653 ( .A(n46259), .B(n46260), .Z(n46242) );
  NANDN U55654 ( .A(n46261), .B(n46262), .Z(n46260) );
  OR U55655 ( .A(n46263), .B(n46264), .Z(n46262) );
  IV U55656 ( .A(n46265), .Z(n46264) );
  NANDN U55657 ( .A(n46265), .B(n46263), .Z(n46259) );
  AND U55658 ( .A(n46266), .B(n46267), .Z(n46240) );
  NAND U55659 ( .A(n46268), .B(n46269), .Z(n46267) );
  NANDN U55660 ( .A(n46270), .B(n46271), .Z(n46269) );
  NANDN U55661 ( .A(n46271), .B(n46270), .Z(n46266) );
  IV U55662 ( .A(n46272), .Z(n46271) );
  NAND U55663 ( .A(n46273), .B(n46274), .Z(n46243) );
  NANDN U55664 ( .A(n46275), .B(n46276), .Z(n46274) );
  NANDN U55665 ( .A(n46277), .B(n46278), .Z(n46276) );
  NANDN U55666 ( .A(n46278), .B(n46277), .Z(n46273) );
  IV U55667 ( .A(n46279), .Z(n46277) );
  AND U55668 ( .A(n46280), .B(n46281), .Z(n46246) );
  NAND U55669 ( .A(n46282), .B(n46283), .Z(n46281) );
  NANDN U55670 ( .A(n46284), .B(n46285), .Z(n46283) );
  NANDN U55671 ( .A(n46285), .B(n46284), .Z(n46280) );
  XOR U55672 ( .A(n46256), .B(n46286), .Z(n46248) );
  XNOR U55673 ( .A(n46253), .B(n46255), .Z(n46286) );
  AND U55674 ( .A(n46287), .B(n46288), .Z(n46255) );
  NANDN U55675 ( .A(n46289), .B(n46290), .Z(n46288) );
  OR U55676 ( .A(n46291), .B(n46292), .Z(n46290) );
  IV U55677 ( .A(n46293), .Z(n46292) );
  NANDN U55678 ( .A(n46293), .B(n46291), .Z(n46287) );
  AND U55679 ( .A(n46294), .B(n46295), .Z(n46253) );
  NAND U55680 ( .A(n46296), .B(n46297), .Z(n46295) );
  NANDN U55681 ( .A(n46298), .B(n46299), .Z(n46297) );
  NANDN U55682 ( .A(n46299), .B(n46298), .Z(n46294) );
  IV U55683 ( .A(n46300), .Z(n46299) );
  NAND U55684 ( .A(n46301), .B(n46302), .Z(n46256) );
  NANDN U55685 ( .A(n46303), .B(n46304), .Z(n46302) );
  NANDN U55686 ( .A(n46305), .B(n46306), .Z(n46304) );
  NANDN U55687 ( .A(n46306), .B(n46305), .Z(n46301) );
  IV U55688 ( .A(n46307), .Z(n46305) );
  XOR U55689 ( .A(n46282), .B(n46308), .Z(N61269) );
  XNOR U55690 ( .A(n46285), .B(n46284), .Z(n46308) );
  XNOR U55691 ( .A(n46296), .B(n46309), .Z(n46284) );
  XNOR U55692 ( .A(n46300), .B(n46298), .Z(n46309) );
  XOR U55693 ( .A(n46306), .B(n46310), .Z(n46298) );
  XNOR U55694 ( .A(n46303), .B(n46307), .Z(n46310) );
  AND U55695 ( .A(n46311), .B(n46312), .Z(n46307) );
  NAND U55696 ( .A(n46313), .B(n46314), .Z(n46312) );
  NAND U55697 ( .A(n46315), .B(n46316), .Z(n46311) );
  AND U55698 ( .A(n46317), .B(n46318), .Z(n46303) );
  NAND U55699 ( .A(n46319), .B(n46320), .Z(n46318) );
  NAND U55700 ( .A(n46321), .B(n46322), .Z(n46317) );
  NANDN U55701 ( .A(n46323), .B(n46324), .Z(n46306) );
  ANDN U55702 ( .B(n46325), .A(n46326), .Z(n46300) );
  XNOR U55703 ( .A(n46291), .B(n46327), .Z(n46296) );
  XNOR U55704 ( .A(n46289), .B(n46293), .Z(n46327) );
  AND U55705 ( .A(n46328), .B(n46329), .Z(n46293) );
  NAND U55706 ( .A(n46330), .B(n46331), .Z(n46329) );
  NAND U55707 ( .A(n46332), .B(n46333), .Z(n46328) );
  AND U55708 ( .A(n46334), .B(n46335), .Z(n46289) );
  NAND U55709 ( .A(n46336), .B(n46337), .Z(n46335) );
  NAND U55710 ( .A(n46338), .B(n46339), .Z(n46334) );
  AND U55711 ( .A(n46340), .B(n46341), .Z(n46291) );
  NAND U55712 ( .A(n46342), .B(n46343), .Z(n46285) );
  XNOR U55713 ( .A(n46268), .B(n46344), .Z(n46282) );
  XNOR U55714 ( .A(n46272), .B(n46270), .Z(n46344) );
  XOR U55715 ( .A(n46278), .B(n46345), .Z(n46270) );
  XNOR U55716 ( .A(n46275), .B(n46279), .Z(n46345) );
  AND U55717 ( .A(n46346), .B(n46347), .Z(n46279) );
  NAND U55718 ( .A(n46348), .B(n46349), .Z(n46347) );
  NAND U55719 ( .A(n46350), .B(n46351), .Z(n46346) );
  AND U55720 ( .A(n46352), .B(n46353), .Z(n46275) );
  NAND U55721 ( .A(n46354), .B(n46355), .Z(n46353) );
  NAND U55722 ( .A(n46356), .B(n46357), .Z(n46352) );
  NANDN U55723 ( .A(n46358), .B(n46359), .Z(n46278) );
  ANDN U55724 ( .B(n46360), .A(n46361), .Z(n46272) );
  XNOR U55725 ( .A(n46263), .B(n46362), .Z(n46268) );
  XNOR U55726 ( .A(n46261), .B(n46265), .Z(n46362) );
  AND U55727 ( .A(n46363), .B(n46364), .Z(n46265) );
  NAND U55728 ( .A(n46365), .B(n46366), .Z(n46364) );
  NAND U55729 ( .A(n46367), .B(n46368), .Z(n46363) );
  AND U55730 ( .A(n46369), .B(n46370), .Z(n46261) );
  NAND U55731 ( .A(n46371), .B(n46372), .Z(n46370) );
  NAND U55732 ( .A(n46373), .B(n46374), .Z(n46369) );
  AND U55733 ( .A(n46375), .B(n46376), .Z(n46263) );
  XOR U55734 ( .A(n46343), .B(n46342), .Z(N61268) );
  XNOR U55735 ( .A(n46360), .B(n46361), .Z(n46342) );
  XNOR U55736 ( .A(n46375), .B(n46376), .Z(n46361) );
  XOR U55737 ( .A(n46372), .B(n46371), .Z(n46376) );
  XOR U55738 ( .A(y[1260]), .B(x[1260]), .Z(n46371) );
  XOR U55739 ( .A(n46374), .B(n46373), .Z(n46372) );
  XOR U55740 ( .A(y[1262]), .B(x[1262]), .Z(n46373) );
  XOR U55741 ( .A(y[1261]), .B(x[1261]), .Z(n46374) );
  XOR U55742 ( .A(n46366), .B(n46365), .Z(n46375) );
  XOR U55743 ( .A(n46368), .B(n46367), .Z(n46365) );
  XOR U55744 ( .A(y[1259]), .B(x[1259]), .Z(n46367) );
  XOR U55745 ( .A(y[1258]), .B(x[1258]), .Z(n46368) );
  XOR U55746 ( .A(y[1257]), .B(x[1257]), .Z(n46366) );
  XNOR U55747 ( .A(n46359), .B(n46358), .Z(n46360) );
  XNOR U55748 ( .A(n46355), .B(n46354), .Z(n46358) );
  XOR U55749 ( .A(n46357), .B(n46356), .Z(n46354) );
  XOR U55750 ( .A(y[1256]), .B(x[1256]), .Z(n46356) );
  XOR U55751 ( .A(y[1255]), .B(x[1255]), .Z(n46357) );
  XOR U55752 ( .A(y[1254]), .B(x[1254]), .Z(n46355) );
  XOR U55753 ( .A(n46349), .B(n46348), .Z(n46359) );
  XOR U55754 ( .A(n46351), .B(n46350), .Z(n46348) );
  XOR U55755 ( .A(y[1253]), .B(x[1253]), .Z(n46350) );
  XOR U55756 ( .A(y[1252]), .B(x[1252]), .Z(n46351) );
  XOR U55757 ( .A(y[1251]), .B(x[1251]), .Z(n46349) );
  XNOR U55758 ( .A(n46325), .B(n46326), .Z(n46343) );
  XNOR U55759 ( .A(n46340), .B(n46341), .Z(n46326) );
  XOR U55760 ( .A(n46337), .B(n46336), .Z(n46341) );
  XOR U55761 ( .A(y[1248]), .B(x[1248]), .Z(n46336) );
  XOR U55762 ( .A(n46339), .B(n46338), .Z(n46337) );
  XOR U55763 ( .A(y[1250]), .B(x[1250]), .Z(n46338) );
  XOR U55764 ( .A(y[1249]), .B(x[1249]), .Z(n46339) );
  XOR U55765 ( .A(n46331), .B(n46330), .Z(n46340) );
  XOR U55766 ( .A(n46333), .B(n46332), .Z(n46330) );
  XOR U55767 ( .A(y[1247]), .B(x[1247]), .Z(n46332) );
  XOR U55768 ( .A(y[1246]), .B(x[1246]), .Z(n46333) );
  XOR U55769 ( .A(y[1245]), .B(x[1245]), .Z(n46331) );
  XNOR U55770 ( .A(n46324), .B(n46323), .Z(n46325) );
  XNOR U55771 ( .A(n46320), .B(n46319), .Z(n46323) );
  XOR U55772 ( .A(n46322), .B(n46321), .Z(n46319) );
  XOR U55773 ( .A(y[1244]), .B(x[1244]), .Z(n46321) );
  XOR U55774 ( .A(y[1243]), .B(x[1243]), .Z(n46322) );
  XOR U55775 ( .A(y[1242]), .B(x[1242]), .Z(n46320) );
  XOR U55776 ( .A(n46314), .B(n46313), .Z(n46324) );
  XOR U55777 ( .A(n46316), .B(n46315), .Z(n46313) );
  XOR U55778 ( .A(y[1241]), .B(x[1241]), .Z(n46315) );
  XOR U55779 ( .A(y[1240]), .B(x[1240]), .Z(n46316) );
  XOR U55780 ( .A(y[1239]), .B(x[1239]), .Z(n46314) );
  NAND U55781 ( .A(n46377), .B(n46378), .Z(N61259) );
  NAND U55782 ( .A(n46379), .B(n46380), .Z(n46378) );
  NANDN U55783 ( .A(n46381), .B(n46382), .Z(n46380) );
  NANDN U55784 ( .A(n46382), .B(n46381), .Z(n46377) );
  XOR U55785 ( .A(n46381), .B(n46383), .Z(N61258) );
  XNOR U55786 ( .A(n46379), .B(n46382), .Z(n46383) );
  NAND U55787 ( .A(n46384), .B(n46385), .Z(n46382) );
  NAND U55788 ( .A(n46386), .B(n46387), .Z(n46385) );
  NANDN U55789 ( .A(n46388), .B(n46389), .Z(n46387) );
  NANDN U55790 ( .A(n46389), .B(n46388), .Z(n46384) );
  AND U55791 ( .A(n46390), .B(n46391), .Z(n46379) );
  NAND U55792 ( .A(n46392), .B(n46393), .Z(n46391) );
  NANDN U55793 ( .A(n46394), .B(n46395), .Z(n46393) );
  NANDN U55794 ( .A(n46395), .B(n46394), .Z(n46390) );
  IV U55795 ( .A(n46396), .Z(n46395) );
  AND U55796 ( .A(n46397), .B(n46398), .Z(n46381) );
  NAND U55797 ( .A(n46399), .B(n46400), .Z(n46398) );
  NANDN U55798 ( .A(n46401), .B(n46402), .Z(n46400) );
  NANDN U55799 ( .A(n46402), .B(n46401), .Z(n46397) );
  XOR U55800 ( .A(n46394), .B(n46403), .Z(N61257) );
  XNOR U55801 ( .A(n46392), .B(n46396), .Z(n46403) );
  XOR U55802 ( .A(n46389), .B(n46404), .Z(n46396) );
  XNOR U55803 ( .A(n46386), .B(n46388), .Z(n46404) );
  AND U55804 ( .A(n46405), .B(n46406), .Z(n46388) );
  NANDN U55805 ( .A(n46407), .B(n46408), .Z(n46406) );
  OR U55806 ( .A(n46409), .B(n46410), .Z(n46408) );
  IV U55807 ( .A(n46411), .Z(n46410) );
  NANDN U55808 ( .A(n46411), .B(n46409), .Z(n46405) );
  AND U55809 ( .A(n46412), .B(n46413), .Z(n46386) );
  NAND U55810 ( .A(n46414), .B(n46415), .Z(n46413) );
  NANDN U55811 ( .A(n46416), .B(n46417), .Z(n46415) );
  NANDN U55812 ( .A(n46417), .B(n46416), .Z(n46412) );
  IV U55813 ( .A(n46418), .Z(n46417) );
  NAND U55814 ( .A(n46419), .B(n46420), .Z(n46389) );
  NANDN U55815 ( .A(n46421), .B(n46422), .Z(n46420) );
  NANDN U55816 ( .A(n46423), .B(n46424), .Z(n46422) );
  NANDN U55817 ( .A(n46424), .B(n46423), .Z(n46419) );
  IV U55818 ( .A(n46425), .Z(n46423) );
  AND U55819 ( .A(n46426), .B(n46427), .Z(n46392) );
  NAND U55820 ( .A(n46428), .B(n46429), .Z(n46427) );
  NANDN U55821 ( .A(n46430), .B(n46431), .Z(n46429) );
  NANDN U55822 ( .A(n46431), .B(n46430), .Z(n46426) );
  XOR U55823 ( .A(n46402), .B(n46432), .Z(n46394) );
  XNOR U55824 ( .A(n46399), .B(n46401), .Z(n46432) );
  AND U55825 ( .A(n46433), .B(n46434), .Z(n46401) );
  NANDN U55826 ( .A(n46435), .B(n46436), .Z(n46434) );
  OR U55827 ( .A(n46437), .B(n46438), .Z(n46436) );
  IV U55828 ( .A(n46439), .Z(n46438) );
  NANDN U55829 ( .A(n46439), .B(n46437), .Z(n46433) );
  AND U55830 ( .A(n46440), .B(n46441), .Z(n46399) );
  NAND U55831 ( .A(n46442), .B(n46443), .Z(n46441) );
  NANDN U55832 ( .A(n46444), .B(n46445), .Z(n46443) );
  NANDN U55833 ( .A(n46445), .B(n46444), .Z(n46440) );
  IV U55834 ( .A(n46446), .Z(n46445) );
  NAND U55835 ( .A(n46447), .B(n46448), .Z(n46402) );
  NANDN U55836 ( .A(n46449), .B(n46450), .Z(n46448) );
  NANDN U55837 ( .A(n46451), .B(n46452), .Z(n46450) );
  NANDN U55838 ( .A(n46452), .B(n46451), .Z(n46447) );
  IV U55839 ( .A(n46453), .Z(n46451) );
  XOR U55840 ( .A(n46428), .B(n46454), .Z(N61256) );
  XNOR U55841 ( .A(n46431), .B(n46430), .Z(n46454) );
  XNOR U55842 ( .A(n46442), .B(n46455), .Z(n46430) );
  XNOR U55843 ( .A(n46446), .B(n46444), .Z(n46455) );
  XOR U55844 ( .A(n46452), .B(n46456), .Z(n46444) );
  XNOR U55845 ( .A(n46449), .B(n46453), .Z(n46456) );
  AND U55846 ( .A(n46457), .B(n46458), .Z(n46453) );
  NAND U55847 ( .A(n46459), .B(n46460), .Z(n46458) );
  NAND U55848 ( .A(n46461), .B(n46462), .Z(n46457) );
  AND U55849 ( .A(n46463), .B(n46464), .Z(n46449) );
  NAND U55850 ( .A(n46465), .B(n46466), .Z(n46464) );
  NAND U55851 ( .A(n46467), .B(n46468), .Z(n46463) );
  NANDN U55852 ( .A(n46469), .B(n46470), .Z(n46452) );
  ANDN U55853 ( .B(n46471), .A(n46472), .Z(n46446) );
  XNOR U55854 ( .A(n46437), .B(n46473), .Z(n46442) );
  XNOR U55855 ( .A(n46435), .B(n46439), .Z(n46473) );
  AND U55856 ( .A(n46474), .B(n46475), .Z(n46439) );
  NAND U55857 ( .A(n46476), .B(n46477), .Z(n46475) );
  NAND U55858 ( .A(n46478), .B(n46479), .Z(n46474) );
  AND U55859 ( .A(n46480), .B(n46481), .Z(n46435) );
  NAND U55860 ( .A(n46482), .B(n46483), .Z(n46481) );
  NAND U55861 ( .A(n46484), .B(n46485), .Z(n46480) );
  AND U55862 ( .A(n46486), .B(n46487), .Z(n46437) );
  NAND U55863 ( .A(n46488), .B(n46489), .Z(n46431) );
  XNOR U55864 ( .A(n46414), .B(n46490), .Z(n46428) );
  XNOR U55865 ( .A(n46418), .B(n46416), .Z(n46490) );
  XOR U55866 ( .A(n46424), .B(n46491), .Z(n46416) );
  XNOR U55867 ( .A(n46421), .B(n46425), .Z(n46491) );
  AND U55868 ( .A(n46492), .B(n46493), .Z(n46425) );
  NAND U55869 ( .A(n46494), .B(n46495), .Z(n46493) );
  NAND U55870 ( .A(n46496), .B(n46497), .Z(n46492) );
  AND U55871 ( .A(n46498), .B(n46499), .Z(n46421) );
  NAND U55872 ( .A(n46500), .B(n46501), .Z(n46499) );
  NAND U55873 ( .A(n46502), .B(n46503), .Z(n46498) );
  NANDN U55874 ( .A(n46504), .B(n46505), .Z(n46424) );
  ANDN U55875 ( .B(n46506), .A(n46507), .Z(n46418) );
  XNOR U55876 ( .A(n46409), .B(n46508), .Z(n46414) );
  XNOR U55877 ( .A(n46407), .B(n46411), .Z(n46508) );
  AND U55878 ( .A(n46509), .B(n46510), .Z(n46411) );
  NAND U55879 ( .A(n46511), .B(n46512), .Z(n46510) );
  NAND U55880 ( .A(n46513), .B(n46514), .Z(n46509) );
  AND U55881 ( .A(n46515), .B(n46516), .Z(n46407) );
  NAND U55882 ( .A(n46517), .B(n46518), .Z(n46516) );
  NAND U55883 ( .A(n46519), .B(n46520), .Z(n46515) );
  AND U55884 ( .A(n46521), .B(n46522), .Z(n46409) );
  XOR U55885 ( .A(n46489), .B(n46488), .Z(N61255) );
  XNOR U55886 ( .A(n46506), .B(n46507), .Z(n46488) );
  XNOR U55887 ( .A(n46521), .B(n46522), .Z(n46507) );
  XOR U55888 ( .A(n46518), .B(n46517), .Z(n46522) );
  XOR U55889 ( .A(y[1236]), .B(x[1236]), .Z(n46517) );
  XOR U55890 ( .A(n46520), .B(n46519), .Z(n46518) );
  XOR U55891 ( .A(y[1238]), .B(x[1238]), .Z(n46519) );
  XOR U55892 ( .A(y[1237]), .B(x[1237]), .Z(n46520) );
  XOR U55893 ( .A(n46512), .B(n46511), .Z(n46521) );
  XOR U55894 ( .A(n46514), .B(n46513), .Z(n46511) );
  XOR U55895 ( .A(y[1235]), .B(x[1235]), .Z(n46513) );
  XOR U55896 ( .A(y[1234]), .B(x[1234]), .Z(n46514) );
  XOR U55897 ( .A(y[1233]), .B(x[1233]), .Z(n46512) );
  XNOR U55898 ( .A(n46505), .B(n46504), .Z(n46506) );
  XNOR U55899 ( .A(n46501), .B(n46500), .Z(n46504) );
  XOR U55900 ( .A(n46503), .B(n46502), .Z(n46500) );
  XOR U55901 ( .A(y[1232]), .B(x[1232]), .Z(n46502) );
  XOR U55902 ( .A(y[1231]), .B(x[1231]), .Z(n46503) );
  XOR U55903 ( .A(y[1230]), .B(x[1230]), .Z(n46501) );
  XOR U55904 ( .A(n46495), .B(n46494), .Z(n46505) );
  XOR U55905 ( .A(n46497), .B(n46496), .Z(n46494) );
  XOR U55906 ( .A(y[1229]), .B(x[1229]), .Z(n46496) );
  XOR U55907 ( .A(y[1228]), .B(x[1228]), .Z(n46497) );
  XOR U55908 ( .A(y[1227]), .B(x[1227]), .Z(n46495) );
  XNOR U55909 ( .A(n46471), .B(n46472), .Z(n46489) );
  XNOR U55910 ( .A(n46486), .B(n46487), .Z(n46472) );
  XOR U55911 ( .A(n46483), .B(n46482), .Z(n46487) );
  XOR U55912 ( .A(y[1224]), .B(x[1224]), .Z(n46482) );
  XOR U55913 ( .A(n46485), .B(n46484), .Z(n46483) );
  XOR U55914 ( .A(y[1226]), .B(x[1226]), .Z(n46484) );
  XOR U55915 ( .A(y[1225]), .B(x[1225]), .Z(n46485) );
  XOR U55916 ( .A(n46477), .B(n46476), .Z(n46486) );
  XOR U55917 ( .A(n46479), .B(n46478), .Z(n46476) );
  XOR U55918 ( .A(y[1223]), .B(x[1223]), .Z(n46478) );
  XOR U55919 ( .A(y[1222]), .B(x[1222]), .Z(n46479) );
  XOR U55920 ( .A(y[1221]), .B(x[1221]), .Z(n46477) );
  XNOR U55921 ( .A(n46470), .B(n46469), .Z(n46471) );
  XNOR U55922 ( .A(n46466), .B(n46465), .Z(n46469) );
  XOR U55923 ( .A(n46468), .B(n46467), .Z(n46465) );
  XOR U55924 ( .A(y[1220]), .B(x[1220]), .Z(n46467) );
  XOR U55925 ( .A(y[1219]), .B(x[1219]), .Z(n46468) );
  XOR U55926 ( .A(y[1218]), .B(x[1218]), .Z(n46466) );
  XOR U55927 ( .A(n46460), .B(n46459), .Z(n46470) );
  XOR U55928 ( .A(n46462), .B(n46461), .Z(n46459) );
  XOR U55929 ( .A(y[1217]), .B(x[1217]), .Z(n46461) );
  XOR U55930 ( .A(y[1216]), .B(x[1216]), .Z(n46462) );
  XOR U55931 ( .A(y[1215]), .B(x[1215]), .Z(n46460) );
  NAND U55932 ( .A(n46523), .B(n46524), .Z(N61246) );
  NAND U55933 ( .A(n46525), .B(n46526), .Z(n46524) );
  NANDN U55934 ( .A(n46527), .B(n46528), .Z(n46526) );
  NANDN U55935 ( .A(n46528), .B(n46527), .Z(n46523) );
  XOR U55936 ( .A(n46527), .B(n46529), .Z(N61245) );
  XNOR U55937 ( .A(n46525), .B(n46528), .Z(n46529) );
  NAND U55938 ( .A(n46530), .B(n46531), .Z(n46528) );
  NAND U55939 ( .A(n46532), .B(n46533), .Z(n46531) );
  NANDN U55940 ( .A(n46534), .B(n46535), .Z(n46533) );
  NANDN U55941 ( .A(n46535), .B(n46534), .Z(n46530) );
  AND U55942 ( .A(n46536), .B(n46537), .Z(n46525) );
  NAND U55943 ( .A(n46538), .B(n46539), .Z(n46537) );
  NANDN U55944 ( .A(n46540), .B(n46541), .Z(n46539) );
  NANDN U55945 ( .A(n46541), .B(n46540), .Z(n46536) );
  IV U55946 ( .A(n46542), .Z(n46541) );
  AND U55947 ( .A(n46543), .B(n46544), .Z(n46527) );
  NAND U55948 ( .A(n46545), .B(n46546), .Z(n46544) );
  NANDN U55949 ( .A(n46547), .B(n46548), .Z(n46546) );
  NANDN U55950 ( .A(n46548), .B(n46547), .Z(n46543) );
  XOR U55951 ( .A(n46540), .B(n46549), .Z(N61244) );
  XNOR U55952 ( .A(n46538), .B(n46542), .Z(n46549) );
  XOR U55953 ( .A(n46535), .B(n46550), .Z(n46542) );
  XNOR U55954 ( .A(n46532), .B(n46534), .Z(n46550) );
  AND U55955 ( .A(n46551), .B(n46552), .Z(n46534) );
  NANDN U55956 ( .A(n46553), .B(n46554), .Z(n46552) );
  OR U55957 ( .A(n46555), .B(n46556), .Z(n46554) );
  IV U55958 ( .A(n46557), .Z(n46556) );
  NANDN U55959 ( .A(n46557), .B(n46555), .Z(n46551) );
  AND U55960 ( .A(n46558), .B(n46559), .Z(n46532) );
  NAND U55961 ( .A(n46560), .B(n46561), .Z(n46559) );
  NANDN U55962 ( .A(n46562), .B(n46563), .Z(n46561) );
  NANDN U55963 ( .A(n46563), .B(n46562), .Z(n46558) );
  IV U55964 ( .A(n46564), .Z(n46563) );
  NAND U55965 ( .A(n46565), .B(n46566), .Z(n46535) );
  NANDN U55966 ( .A(n46567), .B(n46568), .Z(n46566) );
  NANDN U55967 ( .A(n46569), .B(n46570), .Z(n46568) );
  NANDN U55968 ( .A(n46570), .B(n46569), .Z(n46565) );
  IV U55969 ( .A(n46571), .Z(n46569) );
  AND U55970 ( .A(n46572), .B(n46573), .Z(n46538) );
  NAND U55971 ( .A(n46574), .B(n46575), .Z(n46573) );
  NANDN U55972 ( .A(n46576), .B(n46577), .Z(n46575) );
  NANDN U55973 ( .A(n46577), .B(n46576), .Z(n46572) );
  XOR U55974 ( .A(n46548), .B(n46578), .Z(n46540) );
  XNOR U55975 ( .A(n46545), .B(n46547), .Z(n46578) );
  AND U55976 ( .A(n46579), .B(n46580), .Z(n46547) );
  NANDN U55977 ( .A(n46581), .B(n46582), .Z(n46580) );
  OR U55978 ( .A(n46583), .B(n46584), .Z(n46582) );
  IV U55979 ( .A(n46585), .Z(n46584) );
  NANDN U55980 ( .A(n46585), .B(n46583), .Z(n46579) );
  AND U55981 ( .A(n46586), .B(n46587), .Z(n46545) );
  NAND U55982 ( .A(n46588), .B(n46589), .Z(n46587) );
  NANDN U55983 ( .A(n46590), .B(n46591), .Z(n46589) );
  NANDN U55984 ( .A(n46591), .B(n46590), .Z(n46586) );
  IV U55985 ( .A(n46592), .Z(n46591) );
  NAND U55986 ( .A(n46593), .B(n46594), .Z(n46548) );
  NANDN U55987 ( .A(n46595), .B(n46596), .Z(n46594) );
  NANDN U55988 ( .A(n46597), .B(n46598), .Z(n46596) );
  NANDN U55989 ( .A(n46598), .B(n46597), .Z(n46593) );
  IV U55990 ( .A(n46599), .Z(n46597) );
  XOR U55991 ( .A(n46574), .B(n46600), .Z(N61243) );
  XNOR U55992 ( .A(n46577), .B(n46576), .Z(n46600) );
  XNOR U55993 ( .A(n46588), .B(n46601), .Z(n46576) );
  XNOR U55994 ( .A(n46592), .B(n46590), .Z(n46601) );
  XOR U55995 ( .A(n46598), .B(n46602), .Z(n46590) );
  XNOR U55996 ( .A(n46595), .B(n46599), .Z(n46602) );
  AND U55997 ( .A(n46603), .B(n46604), .Z(n46599) );
  NAND U55998 ( .A(n46605), .B(n46606), .Z(n46604) );
  NAND U55999 ( .A(n46607), .B(n46608), .Z(n46603) );
  AND U56000 ( .A(n46609), .B(n46610), .Z(n46595) );
  NAND U56001 ( .A(n46611), .B(n46612), .Z(n46610) );
  NAND U56002 ( .A(n46613), .B(n46614), .Z(n46609) );
  NANDN U56003 ( .A(n46615), .B(n46616), .Z(n46598) );
  ANDN U56004 ( .B(n46617), .A(n46618), .Z(n46592) );
  XNOR U56005 ( .A(n46583), .B(n46619), .Z(n46588) );
  XNOR U56006 ( .A(n46581), .B(n46585), .Z(n46619) );
  AND U56007 ( .A(n46620), .B(n46621), .Z(n46585) );
  NAND U56008 ( .A(n46622), .B(n46623), .Z(n46621) );
  NAND U56009 ( .A(n46624), .B(n46625), .Z(n46620) );
  AND U56010 ( .A(n46626), .B(n46627), .Z(n46581) );
  NAND U56011 ( .A(n46628), .B(n46629), .Z(n46627) );
  NAND U56012 ( .A(n46630), .B(n46631), .Z(n46626) );
  AND U56013 ( .A(n46632), .B(n46633), .Z(n46583) );
  NAND U56014 ( .A(n46634), .B(n46635), .Z(n46577) );
  XNOR U56015 ( .A(n46560), .B(n46636), .Z(n46574) );
  XNOR U56016 ( .A(n46564), .B(n46562), .Z(n46636) );
  XOR U56017 ( .A(n46570), .B(n46637), .Z(n46562) );
  XNOR U56018 ( .A(n46567), .B(n46571), .Z(n46637) );
  AND U56019 ( .A(n46638), .B(n46639), .Z(n46571) );
  NAND U56020 ( .A(n46640), .B(n46641), .Z(n46639) );
  NAND U56021 ( .A(n46642), .B(n46643), .Z(n46638) );
  AND U56022 ( .A(n46644), .B(n46645), .Z(n46567) );
  NAND U56023 ( .A(n46646), .B(n46647), .Z(n46645) );
  NAND U56024 ( .A(n46648), .B(n46649), .Z(n46644) );
  NANDN U56025 ( .A(n46650), .B(n46651), .Z(n46570) );
  ANDN U56026 ( .B(n46652), .A(n46653), .Z(n46564) );
  XNOR U56027 ( .A(n46555), .B(n46654), .Z(n46560) );
  XNOR U56028 ( .A(n46553), .B(n46557), .Z(n46654) );
  AND U56029 ( .A(n46655), .B(n46656), .Z(n46557) );
  NAND U56030 ( .A(n46657), .B(n46658), .Z(n46656) );
  NAND U56031 ( .A(n46659), .B(n46660), .Z(n46655) );
  AND U56032 ( .A(n46661), .B(n46662), .Z(n46553) );
  NAND U56033 ( .A(n46663), .B(n46664), .Z(n46662) );
  NAND U56034 ( .A(n46665), .B(n46666), .Z(n46661) );
  AND U56035 ( .A(n46667), .B(n46668), .Z(n46555) );
  XOR U56036 ( .A(n46635), .B(n46634), .Z(N61242) );
  XNOR U56037 ( .A(n46652), .B(n46653), .Z(n46634) );
  XNOR U56038 ( .A(n46667), .B(n46668), .Z(n46653) );
  XOR U56039 ( .A(n46664), .B(n46663), .Z(n46668) );
  XOR U56040 ( .A(y[1212]), .B(x[1212]), .Z(n46663) );
  XOR U56041 ( .A(n46666), .B(n46665), .Z(n46664) );
  XOR U56042 ( .A(y[1214]), .B(x[1214]), .Z(n46665) );
  XOR U56043 ( .A(y[1213]), .B(x[1213]), .Z(n46666) );
  XOR U56044 ( .A(n46658), .B(n46657), .Z(n46667) );
  XOR U56045 ( .A(n46660), .B(n46659), .Z(n46657) );
  XOR U56046 ( .A(y[1211]), .B(x[1211]), .Z(n46659) );
  XOR U56047 ( .A(y[1210]), .B(x[1210]), .Z(n46660) );
  XOR U56048 ( .A(y[1209]), .B(x[1209]), .Z(n46658) );
  XNOR U56049 ( .A(n46651), .B(n46650), .Z(n46652) );
  XNOR U56050 ( .A(n46647), .B(n46646), .Z(n46650) );
  XOR U56051 ( .A(n46649), .B(n46648), .Z(n46646) );
  XOR U56052 ( .A(y[1208]), .B(x[1208]), .Z(n46648) );
  XOR U56053 ( .A(y[1207]), .B(x[1207]), .Z(n46649) );
  XOR U56054 ( .A(y[1206]), .B(x[1206]), .Z(n46647) );
  XOR U56055 ( .A(n46641), .B(n46640), .Z(n46651) );
  XOR U56056 ( .A(n46643), .B(n46642), .Z(n46640) );
  XOR U56057 ( .A(y[1205]), .B(x[1205]), .Z(n46642) );
  XOR U56058 ( .A(y[1204]), .B(x[1204]), .Z(n46643) );
  XOR U56059 ( .A(y[1203]), .B(x[1203]), .Z(n46641) );
  XNOR U56060 ( .A(n46617), .B(n46618), .Z(n46635) );
  XNOR U56061 ( .A(n46632), .B(n46633), .Z(n46618) );
  XOR U56062 ( .A(n46629), .B(n46628), .Z(n46633) );
  XOR U56063 ( .A(y[1200]), .B(x[1200]), .Z(n46628) );
  XOR U56064 ( .A(n46631), .B(n46630), .Z(n46629) );
  XOR U56065 ( .A(y[1202]), .B(x[1202]), .Z(n46630) );
  XOR U56066 ( .A(y[1201]), .B(x[1201]), .Z(n46631) );
  XOR U56067 ( .A(n46623), .B(n46622), .Z(n46632) );
  XOR U56068 ( .A(n46625), .B(n46624), .Z(n46622) );
  XOR U56069 ( .A(y[1199]), .B(x[1199]), .Z(n46624) );
  XOR U56070 ( .A(y[1198]), .B(x[1198]), .Z(n46625) );
  XOR U56071 ( .A(y[1197]), .B(x[1197]), .Z(n46623) );
  XNOR U56072 ( .A(n46616), .B(n46615), .Z(n46617) );
  XNOR U56073 ( .A(n46612), .B(n46611), .Z(n46615) );
  XOR U56074 ( .A(n46614), .B(n46613), .Z(n46611) );
  XOR U56075 ( .A(y[1196]), .B(x[1196]), .Z(n46613) );
  XOR U56076 ( .A(y[1195]), .B(x[1195]), .Z(n46614) );
  XOR U56077 ( .A(y[1194]), .B(x[1194]), .Z(n46612) );
  XOR U56078 ( .A(n46606), .B(n46605), .Z(n46616) );
  XOR U56079 ( .A(n46608), .B(n46607), .Z(n46605) );
  XOR U56080 ( .A(y[1193]), .B(x[1193]), .Z(n46607) );
  XOR U56081 ( .A(y[1192]), .B(x[1192]), .Z(n46608) );
  XOR U56082 ( .A(y[1191]), .B(x[1191]), .Z(n46606) );
  NAND U56083 ( .A(n46669), .B(n46670), .Z(N61233) );
  NAND U56084 ( .A(n46671), .B(n46672), .Z(n46670) );
  NANDN U56085 ( .A(n46673), .B(n46674), .Z(n46672) );
  NANDN U56086 ( .A(n46674), .B(n46673), .Z(n46669) );
  XOR U56087 ( .A(n46673), .B(n46675), .Z(N61232) );
  XNOR U56088 ( .A(n46671), .B(n46674), .Z(n46675) );
  NAND U56089 ( .A(n46676), .B(n46677), .Z(n46674) );
  NAND U56090 ( .A(n46678), .B(n46679), .Z(n46677) );
  NANDN U56091 ( .A(n46680), .B(n46681), .Z(n46679) );
  NANDN U56092 ( .A(n46681), .B(n46680), .Z(n46676) );
  AND U56093 ( .A(n46682), .B(n46683), .Z(n46671) );
  NAND U56094 ( .A(n46684), .B(n46685), .Z(n46683) );
  NANDN U56095 ( .A(n46686), .B(n46687), .Z(n46685) );
  NANDN U56096 ( .A(n46687), .B(n46686), .Z(n46682) );
  IV U56097 ( .A(n46688), .Z(n46687) );
  AND U56098 ( .A(n46689), .B(n46690), .Z(n46673) );
  NAND U56099 ( .A(n46691), .B(n46692), .Z(n46690) );
  NANDN U56100 ( .A(n46693), .B(n46694), .Z(n46692) );
  NANDN U56101 ( .A(n46694), .B(n46693), .Z(n46689) );
  XOR U56102 ( .A(n46686), .B(n46695), .Z(N61231) );
  XNOR U56103 ( .A(n46684), .B(n46688), .Z(n46695) );
  XOR U56104 ( .A(n46681), .B(n46696), .Z(n46688) );
  XNOR U56105 ( .A(n46678), .B(n46680), .Z(n46696) );
  AND U56106 ( .A(n46697), .B(n46698), .Z(n46680) );
  NANDN U56107 ( .A(n46699), .B(n46700), .Z(n46698) );
  OR U56108 ( .A(n46701), .B(n46702), .Z(n46700) );
  IV U56109 ( .A(n46703), .Z(n46702) );
  NANDN U56110 ( .A(n46703), .B(n46701), .Z(n46697) );
  AND U56111 ( .A(n46704), .B(n46705), .Z(n46678) );
  NAND U56112 ( .A(n46706), .B(n46707), .Z(n46705) );
  NANDN U56113 ( .A(n46708), .B(n46709), .Z(n46707) );
  NANDN U56114 ( .A(n46709), .B(n46708), .Z(n46704) );
  IV U56115 ( .A(n46710), .Z(n46709) );
  NAND U56116 ( .A(n46711), .B(n46712), .Z(n46681) );
  NANDN U56117 ( .A(n46713), .B(n46714), .Z(n46712) );
  NANDN U56118 ( .A(n46715), .B(n46716), .Z(n46714) );
  NANDN U56119 ( .A(n46716), .B(n46715), .Z(n46711) );
  IV U56120 ( .A(n46717), .Z(n46715) );
  AND U56121 ( .A(n46718), .B(n46719), .Z(n46684) );
  NAND U56122 ( .A(n46720), .B(n46721), .Z(n46719) );
  NANDN U56123 ( .A(n46722), .B(n46723), .Z(n46721) );
  NANDN U56124 ( .A(n46723), .B(n46722), .Z(n46718) );
  XOR U56125 ( .A(n46694), .B(n46724), .Z(n46686) );
  XNOR U56126 ( .A(n46691), .B(n46693), .Z(n46724) );
  AND U56127 ( .A(n46725), .B(n46726), .Z(n46693) );
  NANDN U56128 ( .A(n46727), .B(n46728), .Z(n46726) );
  OR U56129 ( .A(n46729), .B(n46730), .Z(n46728) );
  IV U56130 ( .A(n46731), .Z(n46730) );
  NANDN U56131 ( .A(n46731), .B(n46729), .Z(n46725) );
  AND U56132 ( .A(n46732), .B(n46733), .Z(n46691) );
  NAND U56133 ( .A(n46734), .B(n46735), .Z(n46733) );
  NANDN U56134 ( .A(n46736), .B(n46737), .Z(n46735) );
  NANDN U56135 ( .A(n46737), .B(n46736), .Z(n46732) );
  IV U56136 ( .A(n46738), .Z(n46737) );
  NAND U56137 ( .A(n46739), .B(n46740), .Z(n46694) );
  NANDN U56138 ( .A(n46741), .B(n46742), .Z(n46740) );
  NANDN U56139 ( .A(n46743), .B(n46744), .Z(n46742) );
  NANDN U56140 ( .A(n46744), .B(n46743), .Z(n46739) );
  IV U56141 ( .A(n46745), .Z(n46743) );
  XOR U56142 ( .A(n46720), .B(n46746), .Z(N61230) );
  XNOR U56143 ( .A(n46723), .B(n46722), .Z(n46746) );
  XNOR U56144 ( .A(n46734), .B(n46747), .Z(n46722) );
  XNOR U56145 ( .A(n46738), .B(n46736), .Z(n46747) );
  XOR U56146 ( .A(n46744), .B(n46748), .Z(n46736) );
  XNOR U56147 ( .A(n46741), .B(n46745), .Z(n46748) );
  AND U56148 ( .A(n46749), .B(n46750), .Z(n46745) );
  NAND U56149 ( .A(n46751), .B(n46752), .Z(n46750) );
  NAND U56150 ( .A(n46753), .B(n46754), .Z(n46749) );
  AND U56151 ( .A(n46755), .B(n46756), .Z(n46741) );
  NAND U56152 ( .A(n46757), .B(n46758), .Z(n46756) );
  NAND U56153 ( .A(n46759), .B(n46760), .Z(n46755) );
  NANDN U56154 ( .A(n46761), .B(n46762), .Z(n46744) );
  ANDN U56155 ( .B(n46763), .A(n46764), .Z(n46738) );
  XNOR U56156 ( .A(n46729), .B(n46765), .Z(n46734) );
  XNOR U56157 ( .A(n46727), .B(n46731), .Z(n46765) );
  AND U56158 ( .A(n46766), .B(n46767), .Z(n46731) );
  NAND U56159 ( .A(n46768), .B(n46769), .Z(n46767) );
  NAND U56160 ( .A(n46770), .B(n46771), .Z(n46766) );
  AND U56161 ( .A(n46772), .B(n46773), .Z(n46727) );
  NAND U56162 ( .A(n46774), .B(n46775), .Z(n46773) );
  NAND U56163 ( .A(n46776), .B(n46777), .Z(n46772) );
  AND U56164 ( .A(n46778), .B(n46779), .Z(n46729) );
  NAND U56165 ( .A(n46780), .B(n46781), .Z(n46723) );
  XNOR U56166 ( .A(n46706), .B(n46782), .Z(n46720) );
  XNOR U56167 ( .A(n46710), .B(n46708), .Z(n46782) );
  XOR U56168 ( .A(n46716), .B(n46783), .Z(n46708) );
  XNOR U56169 ( .A(n46713), .B(n46717), .Z(n46783) );
  AND U56170 ( .A(n46784), .B(n46785), .Z(n46717) );
  NAND U56171 ( .A(n46786), .B(n46787), .Z(n46785) );
  NAND U56172 ( .A(n46788), .B(n46789), .Z(n46784) );
  AND U56173 ( .A(n46790), .B(n46791), .Z(n46713) );
  NAND U56174 ( .A(n46792), .B(n46793), .Z(n46791) );
  NAND U56175 ( .A(n46794), .B(n46795), .Z(n46790) );
  NANDN U56176 ( .A(n46796), .B(n46797), .Z(n46716) );
  ANDN U56177 ( .B(n46798), .A(n46799), .Z(n46710) );
  XNOR U56178 ( .A(n46701), .B(n46800), .Z(n46706) );
  XNOR U56179 ( .A(n46699), .B(n46703), .Z(n46800) );
  AND U56180 ( .A(n46801), .B(n46802), .Z(n46703) );
  NAND U56181 ( .A(n46803), .B(n46804), .Z(n46802) );
  NAND U56182 ( .A(n46805), .B(n46806), .Z(n46801) );
  AND U56183 ( .A(n46807), .B(n46808), .Z(n46699) );
  NAND U56184 ( .A(n46809), .B(n46810), .Z(n46808) );
  NAND U56185 ( .A(n46811), .B(n46812), .Z(n46807) );
  AND U56186 ( .A(n46813), .B(n46814), .Z(n46701) );
  XOR U56187 ( .A(n46781), .B(n46780), .Z(N61229) );
  XNOR U56188 ( .A(n46798), .B(n46799), .Z(n46780) );
  XNOR U56189 ( .A(n46813), .B(n46814), .Z(n46799) );
  XOR U56190 ( .A(n46810), .B(n46809), .Z(n46814) );
  XOR U56191 ( .A(y[1188]), .B(x[1188]), .Z(n46809) );
  XOR U56192 ( .A(n46812), .B(n46811), .Z(n46810) );
  XOR U56193 ( .A(y[1190]), .B(x[1190]), .Z(n46811) );
  XOR U56194 ( .A(y[1189]), .B(x[1189]), .Z(n46812) );
  XOR U56195 ( .A(n46804), .B(n46803), .Z(n46813) );
  XOR U56196 ( .A(n46806), .B(n46805), .Z(n46803) );
  XOR U56197 ( .A(y[1187]), .B(x[1187]), .Z(n46805) );
  XOR U56198 ( .A(y[1186]), .B(x[1186]), .Z(n46806) );
  XOR U56199 ( .A(y[1185]), .B(x[1185]), .Z(n46804) );
  XNOR U56200 ( .A(n46797), .B(n46796), .Z(n46798) );
  XNOR U56201 ( .A(n46793), .B(n46792), .Z(n46796) );
  XOR U56202 ( .A(n46795), .B(n46794), .Z(n46792) );
  XOR U56203 ( .A(y[1184]), .B(x[1184]), .Z(n46794) );
  XOR U56204 ( .A(y[1183]), .B(x[1183]), .Z(n46795) );
  XOR U56205 ( .A(y[1182]), .B(x[1182]), .Z(n46793) );
  XOR U56206 ( .A(n46787), .B(n46786), .Z(n46797) );
  XOR U56207 ( .A(n46789), .B(n46788), .Z(n46786) );
  XOR U56208 ( .A(y[1181]), .B(x[1181]), .Z(n46788) );
  XOR U56209 ( .A(y[1180]), .B(x[1180]), .Z(n46789) );
  XOR U56210 ( .A(y[1179]), .B(x[1179]), .Z(n46787) );
  XNOR U56211 ( .A(n46763), .B(n46764), .Z(n46781) );
  XNOR U56212 ( .A(n46778), .B(n46779), .Z(n46764) );
  XOR U56213 ( .A(n46775), .B(n46774), .Z(n46779) );
  XOR U56214 ( .A(y[1176]), .B(x[1176]), .Z(n46774) );
  XOR U56215 ( .A(n46777), .B(n46776), .Z(n46775) );
  XOR U56216 ( .A(y[1178]), .B(x[1178]), .Z(n46776) );
  XOR U56217 ( .A(y[1177]), .B(x[1177]), .Z(n46777) );
  XOR U56218 ( .A(n46769), .B(n46768), .Z(n46778) );
  XOR U56219 ( .A(n46771), .B(n46770), .Z(n46768) );
  XOR U56220 ( .A(y[1175]), .B(x[1175]), .Z(n46770) );
  XOR U56221 ( .A(y[1174]), .B(x[1174]), .Z(n46771) );
  XOR U56222 ( .A(y[1173]), .B(x[1173]), .Z(n46769) );
  XNOR U56223 ( .A(n46762), .B(n46761), .Z(n46763) );
  XNOR U56224 ( .A(n46758), .B(n46757), .Z(n46761) );
  XOR U56225 ( .A(n46760), .B(n46759), .Z(n46757) );
  XOR U56226 ( .A(y[1172]), .B(x[1172]), .Z(n46759) );
  XOR U56227 ( .A(y[1171]), .B(x[1171]), .Z(n46760) );
  XOR U56228 ( .A(y[1170]), .B(x[1170]), .Z(n46758) );
  XOR U56229 ( .A(n46752), .B(n46751), .Z(n46762) );
  XOR U56230 ( .A(n46754), .B(n46753), .Z(n46751) );
  XOR U56231 ( .A(y[1169]), .B(x[1169]), .Z(n46753) );
  XOR U56232 ( .A(y[1168]), .B(x[1168]), .Z(n46754) );
  XOR U56233 ( .A(y[1167]), .B(x[1167]), .Z(n46752) );
  NAND U56234 ( .A(n46815), .B(n46816), .Z(N61220) );
  NAND U56235 ( .A(n46817), .B(n46818), .Z(n46816) );
  NANDN U56236 ( .A(n46819), .B(n46820), .Z(n46818) );
  NANDN U56237 ( .A(n46820), .B(n46819), .Z(n46815) );
  XOR U56238 ( .A(n46819), .B(n46821), .Z(N61219) );
  XNOR U56239 ( .A(n46817), .B(n46820), .Z(n46821) );
  NAND U56240 ( .A(n46822), .B(n46823), .Z(n46820) );
  NAND U56241 ( .A(n46824), .B(n46825), .Z(n46823) );
  NANDN U56242 ( .A(n46826), .B(n46827), .Z(n46825) );
  NANDN U56243 ( .A(n46827), .B(n46826), .Z(n46822) );
  AND U56244 ( .A(n46828), .B(n46829), .Z(n46817) );
  NAND U56245 ( .A(n46830), .B(n46831), .Z(n46829) );
  NANDN U56246 ( .A(n46832), .B(n46833), .Z(n46831) );
  NANDN U56247 ( .A(n46833), .B(n46832), .Z(n46828) );
  IV U56248 ( .A(n46834), .Z(n46833) );
  AND U56249 ( .A(n46835), .B(n46836), .Z(n46819) );
  NAND U56250 ( .A(n46837), .B(n46838), .Z(n46836) );
  NANDN U56251 ( .A(n46839), .B(n46840), .Z(n46838) );
  NANDN U56252 ( .A(n46840), .B(n46839), .Z(n46835) );
  XOR U56253 ( .A(n46832), .B(n46841), .Z(N61218) );
  XNOR U56254 ( .A(n46830), .B(n46834), .Z(n46841) );
  XOR U56255 ( .A(n46827), .B(n46842), .Z(n46834) );
  XNOR U56256 ( .A(n46824), .B(n46826), .Z(n46842) );
  AND U56257 ( .A(n46843), .B(n46844), .Z(n46826) );
  NANDN U56258 ( .A(n46845), .B(n46846), .Z(n46844) );
  OR U56259 ( .A(n46847), .B(n46848), .Z(n46846) );
  IV U56260 ( .A(n46849), .Z(n46848) );
  NANDN U56261 ( .A(n46849), .B(n46847), .Z(n46843) );
  AND U56262 ( .A(n46850), .B(n46851), .Z(n46824) );
  NAND U56263 ( .A(n46852), .B(n46853), .Z(n46851) );
  NANDN U56264 ( .A(n46854), .B(n46855), .Z(n46853) );
  NANDN U56265 ( .A(n46855), .B(n46854), .Z(n46850) );
  IV U56266 ( .A(n46856), .Z(n46855) );
  NAND U56267 ( .A(n46857), .B(n46858), .Z(n46827) );
  NANDN U56268 ( .A(n46859), .B(n46860), .Z(n46858) );
  NANDN U56269 ( .A(n46861), .B(n46862), .Z(n46860) );
  NANDN U56270 ( .A(n46862), .B(n46861), .Z(n46857) );
  IV U56271 ( .A(n46863), .Z(n46861) );
  AND U56272 ( .A(n46864), .B(n46865), .Z(n46830) );
  NAND U56273 ( .A(n46866), .B(n46867), .Z(n46865) );
  NANDN U56274 ( .A(n46868), .B(n46869), .Z(n46867) );
  NANDN U56275 ( .A(n46869), .B(n46868), .Z(n46864) );
  XOR U56276 ( .A(n46840), .B(n46870), .Z(n46832) );
  XNOR U56277 ( .A(n46837), .B(n46839), .Z(n46870) );
  AND U56278 ( .A(n46871), .B(n46872), .Z(n46839) );
  NANDN U56279 ( .A(n46873), .B(n46874), .Z(n46872) );
  OR U56280 ( .A(n46875), .B(n46876), .Z(n46874) );
  IV U56281 ( .A(n46877), .Z(n46876) );
  NANDN U56282 ( .A(n46877), .B(n46875), .Z(n46871) );
  AND U56283 ( .A(n46878), .B(n46879), .Z(n46837) );
  NAND U56284 ( .A(n46880), .B(n46881), .Z(n46879) );
  NANDN U56285 ( .A(n46882), .B(n46883), .Z(n46881) );
  NANDN U56286 ( .A(n46883), .B(n46882), .Z(n46878) );
  IV U56287 ( .A(n46884), .Z(n46883) );
  NAND U56288 ( .A(n46885), .B(n46886), .Z(n46840) );
  NANDN U56289 ( .A(n46887), .B(n46888), .Z(n46886) );
  NANDN U56290 ( .A(n46889), .B(n46890), .Z(n46888) );
  NANDN U56291 ( .A(n46890), .B(n46889), .Z(n46885) );
  IV U56292 ( .A(n46891), .Z(n46889) );
  XOR U56293 ( .A(n46866), .B(n46892), .Z(N61217) );
  XNOR U56294 ( .A(n46869), .B(n46868), .Z(n46892) );
  XNOR U56295 ( .A(n46880), .B(n46893), .Z(n46868) );
  XNOR U56296 ( .A(n46884), .B(n46882), .Z(n46893) );
  XOR U56297 ( .A(n46890), .B(n46894), .Z(n46882) );
  XNOR U56298 ( .A(n46887), .B(n46891), .Z(n46894) );
  AND U56299 ( .A(n46895), .B(n46896), .Z(n46891) );
  NAND U56300 ( .A(n46897), .B(n46898), .Z(n46896) );
  NAND U56301 ( .A(n46899), .B(n46900), .Z(n46895) );
  AND U56302 ( .A(n46901), .B(n46902), .Z(n46887) );
  NAND U56303 ( .A(n46903), .B(n46904), .Z(n46902) );
  NAND U56304 ( .A(n46905), .B(n46906), .Z(n46901) );
  NANDN U56305 ( .A(n46907), .B(n46908), .Z(n46890) );
  ANDN U56306 ( .B(n46909), .A(n46910), .Z(n46884) );
  XNOR U56307 ( .A(n46875), .B(n46911), .Z(n46880) );
  XNOR U56308 ( .A(n46873), .B(n46877), .Z(n46911) );
  AND U56309 ( .A(n46912), .B(n46913), .Z(n46877) );
  NAND U56310 ( .A(n46914), .B(n46915), .Z(n46913) );
  NAND U56311 ( .A(n46916), .B(n46917), .Z(n46912) );
  AND U56312 ( .A(n46918), .B(n46919), .Z(n46873) );
  NAND U56313 ( .A(n46920), .B(n46921), .Z(n46919) );
  NAND U56314 ( .A(n46922), .B(n46923), .Z(n46918) );
  AND U56315 ( .A(n46924), .B(n46925), .Z(n46875) );
  NAND U56316 ( .A(n46926), .B(n46927), .Z(n46869) );
  XNOR U56317 ( .A(n46852), .B(n46928), .Z(n46866) );
  XNOR U56318 ( .A(n46856), .B(n46854), .Z(n46928) );
  XOR U56319 ( .A(n46862), .B(n46929), .Z(n46854) );
  XNOR U56320 ( .A(n46859), .B(n46863), .Z(n46929) );
  AND U56321 ( .A(n46930), .B(n46931), .Z(n46863) );
  NAND U56322 ( .A(n46932), .B(n46933), .Z(n46931) );
  NAND U56323 ( .A(n46934), .B(n46935), .Z(n46930) );
  AND U56324 ( .A(n46936), .B(n46937), .Z(n46859) );
  NAND U56325 ( .A(n46938), .B(n46939), .Z(n46937) );
  NAND U56326 ( .A(n46940), .B(n46941), .Z(n46936) );
  NANDN U56327 ( .A(n46942), .B(n46943), .Z(n46862) );
  ANDN U56328 ( .B(n46944), .A(n46945), .Z(n46856) );
  XNOR U56329 ( .A(n46847), .B(n46946), .Z(n46852) );
  XNOR U56330 ( .A(n46845), .B(n46849), .Z(n46946) );
  AND U56331 ( .A(n46947), .B(n46948), .Z(n46849) );
  NAND U56332 ( .A(n46949), .B(n46950), .Z(n46948) );
  NAND U56333 ( .A(n46951), .B(n46952), .Z(n46947) );
  AND U56334 ( .A(n46953), .B(n46954), .Z(n46845) );
  NAND U56335 ( .A(n46955), .B(n46956), .Z(n46954) );
  NAND U56336 ( .A(n46957), .B(n46958), .Z(n46953) );
  AND U56337 ( .A(n46959), .B(n46960), .Z(n46847) );
  XOR U56338 ( .A(n46927), .B(n46926), .Z(N61216) );
  XNOR U56339 ( .A(n46944), .B(n46945), .Z(n46926) );
  XNOR U56340 ( .A(n46959), .B(n46960), .Z(n46945) );
  XOR U56341 ( .A(n46956), .B(n46955), .Z(n46960) );
  XOR U56342 ( .A(y[1164]), .B(x[1164]), .Z(n46955) );
  XOR U56343 ( .A(n46958), .B(n46957), .Z(n46956) );
  XOR U56344 ( .A(y[1166]), .B(x[1166]), .Z(n46957) );
  XOR U56345 ( .A(y[1165]), .B(x[1165]), .Z(n46958) );
  XOR U56346 ( .A(n46950), .B(n46949), .Z(n46959) );
  XOR U56347 ( .A(n46952), .B(n46951), .Z(n46949) );
  XOR U56348 ( .A(y[1163]), .B(x[1163]), .Z(n46951) );
  XOR U56349 ( .A(y[1162]), .B(x[1162]), .Z(n46952) );
  XOR U56350 ( .A(y[1161]), .B(x[1161]), .Z(n46950) );
  XNOR U56351 ( .A(n46943), .B(n46942), .Z(n46944) );
  XNOR U56352 ( .A(n46939), .B(n46938), .Z(n46942) );
  XOR U56353 ( .A(n46941), .B(n46940), .Z(n46938) );
  XOR U56354 ( .A(y[1160]), .B(x[1160]), .Z(n46940) );
  XOR U56355 ( .A(y[1159]), .B(x[1159]), .Z(n46941) );
  XOR U56356 ( .A(y[1158]), .B(x[1158]), .Z(n46939) );
  XOR U56357 ( .A(n46933), .B(n46932), .Z(n46943) );
  XOR U56358 ( .A(n46935), .B(n46934), .Z(n46932) );
  XOR U56359 ( .A(y[1157]), .B(x[1157]), .Z(n46934) );
  XOR U56360 ( .A(y[1156]), .B(x[1156]), .Z(n46935) );
  XOR U56361 ( .A(y[1155]), .B(x[1155]), .Z(n46933) );
  XNOR U56362 ( .A(n46909), .B(n46910), .Z(n46927) );
  XNOR U56363 ( .A(n46924), .B(n46925), .Z(n46910) );
  XOR U56364 ( .A(n46921), .B(n46920), .Z(n46925) );
  XOR U56365 ( .A(y[1152]), .B(x[1152]), .Z(n46920) );
  XOR U56366 ( .A(n46923), .B(n46922), .Z(n46921) );
  XOR U56367 ( .A(y[1154]), .B(x[1154]), .Z(n46922) );
  XOR U56368 ( .A(y[1153]), .B(x[1153]), .Z(n46923) );
  XOR U56369 ( .A(n46915), .B(n46914), .Z(n46924) );
  XOR U56370 ( .A(n46917), .B(n46916), .Z(n46914) );
  XOR U56371 ( .A(y[1151]), .B(x[1151]), .Z(n46916) );
  XOR U56372 ( .A(y[1150]), .B(x[1150]), .Z(n46917) );
  XOR U56373 ( .A(y[1149]), .B(x[1149]), .Z(n46915) );
  XNOR U56374 ( .A(n46908), .B(n46907), .Z(n46909) );
  XNOR U56375 ( .A(n46904), .B(n46903), .Z(n46907) );
  XOR U56376 ( .A(n46906), .B(n46905), .Z(n46903) );
  XOR U56377 ( .A(y[1148]), .B(x[1148]), .Z(n46905) );
  XOR U56378 ( .A(y[1147]), .B(x[1147]), .Z(n46906) );
  XOR U56379 ( .A(y[1146]), .B(x[1146]), .Z(n46904) );
  XOR U56380 ( .A(n46898), .B(n46897), .Z(n46908) );
  XOR U56381 ( .A(n46900), .B(n46899), .Z(n46897) );
  XOR U56382 ( .A(y[1145]), .B(x[1145]), .Z(n46899) );
  XOR U56383 ( .A(y[1144]), .B(x[1144]), .Z(n46900) );
  XOR U56384 ( .A(y[1143]), .B(x[1143]), .Z(n46898) );
  NAND U56385 ( .A(n46961), .B(n46962), .Z(N61207) );
  NAND U56386 ( .A(n46963), .B(n46964), .Z(n46962) );
  NANDN U56387 ( .A(n46965), .B(n46966), .Z(n46964) );
  NANDN U56388 ( .A(n46966), .B(n46965), .Z(n46961) );
  XOR U56389 ( .A(n46965), .B(n46967), .Z(N61206) );
  XNOR U56390 ( .A(n46963), .B(n46966), .Z(n46967) );
  NAND U56391 ( .A(n46968), .B(n46969), .Z(n46966) );
  NAND U56392 ( .A(n46970), .B(n46971), .Z(n46969) );
  NANDN U56393 ( .A(n46972), .B(n46973), .Z(n46971) );
  NANDN U56394 ( .A(n46973), .B(n46972), .Z(n46968) );
  AND U56395 ( .A(n46974), .B(n46975), .Z(n46963) );
  NAND U56396 ( .A(n46976), .B(n46977), .Z(n46975) );
  NANDN U56397 ( .A(n46978), .B(n46979), .Z(n46977) );
  NANDN U56398 ( .A(n46979), .B(n46978), .Z(n46974) );
  IV U56399 ( .A(n46980), .Z(n46979) );
  AND U56400 ( .A(n46981), .B(n46982), .Z(n46965) );
  NAND U56401 ( .A(n46983), .B(n46984), .Z(n46982) );
  NANDN U56402 ( .A(n46985), .B(n46986), .Z(n46984) );
  NANDN U56403 ( .A(n46986), .B(n46985), .Z(n46981) );
  XOR U56404 ( .A(n46978), .B(n46987), .Z(N61205) );
  XNOR U56405 ( .A(n46976), .B(n46980), .Z(n46987) );
  XOR U56406 ( .A(n46973), .B(n46988), .Z(n46980) );
  XNOR U56407 ( .A(n46970), .B(n46972), .Z(n46988) );
  AND U56408 ( .A(n46989), .B(n46990), .Z(n46972) );
  NANDN U56409 ( .A(n46991), .B(n46992), .Z(n46990) );
  OR U56410 ( .A(n46993), .B(n46994), .Z(n46992) );
  IV U56411 ( .A(n46995), .Z(n46994) );
  NANDN U56412 ( .A(n46995), .B(n46993), .Z(n46989) );
  AND U56413 ( .A(n46996), .B(n46997), .Z(n46970) );
  NAND U56414 ( .A(n46998), .B(n46999), .Z(n46997) );
  NANDN U56415 ( .A(n47000), .B(n47001), .Z(n46999) );
  NANDN U56416 ( .A(n47001), .B(n47000), .Z(n46996) );
  IV U56417 ( .A(n47002), .Z(n47001) );
  NAND U56418 ( .A(n47003), .B(n47004), .Z(n46973) );
  NANDN U56419 ( .A(n47005), .B(n47006), .Z(n47004) );
  NANDN U56420 ( .A(n47007), .B(n47008), .Z(n47006) );
  NANDN U56421 ( .A(n47008), .B(n47007), .Z(n47003) );
  IV U56422 ( .A(n47009), .Z(n47007) );
  AND U56423 ( .A(n47010), .B(n47011), .Z(n46976) );
  NAND U56424 ( .A(n47012), .B(n47013), .Z(n47011) );
  NANDN U56425 ( .A(n47014), .B(n47015), .Z(n47013) );
  NANDN U56426 ( .A(n47015), .B(n47014), .Z(n47010) );
  XOR U56427 ( .A(n46986), .B(n47016), .Z(n46978) );
  XNOR U56428 ( .A(n46983), .B(n46985), .Z(n47016) );
  AND U56429 ( .A(n47017), .B(n47018), .Z(n46985) );
  NANDN U56430 ( .A(n47019), .B(n47020), .Z(n47018) );
  OR U56431 ( .A(n47021), .B(n47022), .Z(n47020) );
  IV U56432 ( .A(n47023), .Z(n47022) );
  NANDN U56433 ( .A(n47023), .B(n47021), .Z(n47017) );
  AND U56434 ( .A(n47024), .B(n47025), .Z(n46983) );
  NAND U56435 ( .A(n47026), .B(n47027), .Z(n47025) );
  NANDN U56436 ( .A(n47028), .B(n47029), .Z(n47027) );
  NANDN U56437 ( .A(n47029), .B(n47028), .Z(n47024) );
  IV U56438 ( .A(n47030), .Z(n47029) );
  NAND U56439 ( .A(n47031), .B(n47032), .Z(n46986) );
  NANDN U56440 ( .A(n47033), .B(n47034), .Z(n47032) );
  NANDN U56441 ( .A(n47035), .B(n47036), .Z(n47034) );
  NANDN U56442 ( .A(n47036), .B(n47035), .Z(n47031) );
  IV U56443 ( .A(n47037), .Z(n47035) );
  XOR U56444 ( .A(n47012), .B(n47038), .Z(N61204) );
  XNOR U56445 ( .A(n47015), .B(n47014), .Z(n47038) );
  XNOR U56446 ( .A(n47026), .B(n47039), .Z(n47014) );
  XNOR U56447 ( .A(n47030), .B(n47028), .Z(n47039) );
  XOR U56448 ( .A(n47036), .B(n47040), .Z(n47028) );
  XNOR U56449 ( .A(n47033), .B(n47037), .Z(n47040) );
  AND U56450 ( .A(n47041), .B(n47042), .Z(n47037) );
  NAND U56451 ( .A(n47043), .B(n47044), .Z(n47042) );
  NAND U56452 ( .A(n47045), .B(n47046), .Z(n47041) );
  AND U56453 ( .A(n47047), .B(n47048), .Z(n47033) );
  NAND U56454 ( .A(n47049), .B(n47050), .Z(n47048) );
  NAND U56455 ( .A(n47051), .B(n47052), .Z(n47047) );
  NANDN U56456 ( .A(n47053), .B(n47054), .Z(n47036) );
  ANDN U56457 ( .B(n47055), .A(n47056), .Z(n47030) );
  XNOR U56458 ( .A(n47021), .B(n47057), .Z(n47026) );
  XNOR U56459 ( .A(n47019), .B(n47023), .Z(n47057) );
  AND U56460 ( .A(n47058), .B(n47059), .Z(n47023) );
  NAND U56461 ( .A(n47060), .B(n47061), .Z(n47059) );
  NAND U56462 ( .A(n47062), .B(n47063), .Z(n47058) );
  AND U56463 ( .A(n47064), .B(n47065), .Z(n47019) );
  NAND U56464 ( .A(n47066), .B(n47067), .Z(n47065) );
  NAND U56465 ( .A(n47068), .B(n47069), .Z(n47064) );
  AND U56466 ( .A(n47070), .B(n47071), .Z(n47021) );
  NAND U56467 ( .A(n47072), .B(n47073), .Z(n47015) );
  XNOR U56468 ( .A(n46998), .B(n47074), .Z(n47012) );
  XNOR U56469 ( .A(n47002), .B(n47000), .Z(n47074) );
  XOR U56470 ( .A(n47008), .B(n47075), .Z(n47000) );
  XNOR U56471 ( .A(n47005), .B(n47009), .Z(n47075) );
  AND U56472 ( .A(n47076), .B(n47077), .Z(n47009) );
  NAND U56473 ( .A(n47078), .B(n47079), .Z(n47077) );
  NAND U56474 ( .A(n47080), .B(n47081), .Z(n47076) );
  AND U56475 ( .A(n47082), .B(n47083), .Z(n47005) );
  NAND U56476 ( .A(n47084), .B(n47085), .Z(n47083) );
  NAND U56477 ( .A(n47086), .B(n47087), .Z(n47082) );
  NANDN U56478 ( .A(n47088), .B(n47089), .Z(n47008) );
  ANDN U56479 ( .B(n47090), .A(n47091), .Z(n47002) );
  XNOR U56480 ( .A(n46993), .B(n47092), .Z(n46998) );
  XNOR U56481 ( .A(n46991), .B(n46995), .Z(n47092) );
  AND U56482 ( .A(n47093), .B(n47094), .Z(n46995) );
  NAND U56483 ( .A(n47095), .B(n47096), .Z(n47094) );
  NAND U56484 ( .A(n47097), .B(n47098), .Z(n47093) );
  AND U56485 ( .A(n47099), .B(n47100), .Z(n46991) );
  NAND U56486 ( .A(n47101), .B(n47102), .Z(n47100) );
  NAND U56487 ( .A(n47103), .B(n47104), .Z(n47099) );
  AND U56488 ( .A(n47105), .B(n47106), .Z(n46993) );
  XOR U56489 ( .A(n47073), .B(n47072), .Z(N61203) );
  XNOR U56490 ( .A(n47090), .B(n47091), .Z(n47072) );
  XNOR U56491 ( .A(n47105), .B(n47106), .Z(n47091) );
  XOR U56492 ( .A(n47102), .B(n47101), .Z(n47106) );
  XOR U56493 ( .A(y[1140]), .B(x[1140]), .Z(n47101) );
  XOR U56494 ( .A(n47104), .B(n47103), .Z(n47102) );
  XOR U56495 ( .A(y[1142]), .B(x[1142]), .Z(n47103) );
  XOR U56496 ( .A(y[1141]), .B(x[1141]), .Z(n47104) );
  XOR U56497 ( .A(n47096), .B(n47095), .Z(n47105) );
  XOR U56498 ( .A(n47098), .B(n47097), .Z(n47095) );
  XOR U56499 ( .A(y[1139]), .B(x[1139]), .Z(n47097) );
  XOR U56500 ( .A(y[1138]), .B(x[1138]), .Z(n47098) );
  XOR U56501 ( .A(y[1137]), .B(x[1137]), .Z(n47096) );
  XNOR U56502 ( .A(n47089), .B(n47088), .Z(n47090) );
  XNOR U56503 ( .A(n47085), .B(n47084), .Z(n47088) );
  XOR U56504 ( .A(n47087), .B(n47086), .Z(n47084) );
  XOR U56505 ( .A(y[1136]), .B(x[1136]), .Z(n47086) );
  XOR U56506 ( .A(y[1135]), .B(x[1135]), .Z(n47087) );
  XOR U56507 ( .A(y[1134]), .B(x[1134]), .Z(n47085) );
  XOR U56508 ( .A(n47079), .B(n47078), .Z(n47089) );
  XOR U56509 ( .A(n47081), .B(n47080), .Z(n47078) );
  XOR U56510 ( .A(y[1133]), .B(x[1133]), .Z(n47080) );
  XOR U56511 ( .A(y[1132]), .B(x[1132]), .Z(n47081) );
  XOR U56512 ( .A(y[1131]), .B(x[1131]), .Z(n47079) );
  XNOR U56513 ( .A(n47055), .B(n47056), .Z(n47073) );
  XNOR U56514 ( .A(n47070), .B(n47071), .Z(n47056) );
  XOR U56515 ( .A(n47067), .B(n47066), .Z(n47071) );
  XOR U56516 ( .A(y[1128]), .B(x[1128]), .Z(n47066) );
  XOR U56517 ( .A(n47069), .B(n47068), .Z(n47067) );
  XOR U56518 ( .A(y[1130]), .B(x[1130]), .Z(n47068) );
  XOR U56519 ( .A(y[1129]), .B(x[1129]), .Z(n47069) );
  XOR U56520 ( .A(n47061), .B(n47060), .Z(n47070) );
  XOR U56521 ( .A(n47063), .B(n47062), .Z(n47060) );
  XOR U56522 ( .A(y[1127]), .B(x[1127]), .Z(n47062) );
  XOR U56523 ( .A(y[1126]), .B(x[1126]), .Z(n47063) );
  XOR U56524 ( .A(y[1125]), .B(x[1125]), .Z(n47061) );
  XNOR U56525 ( .A(n47054), .B(n47053), .Z(n47055) );
  XNOR U56526 ( .A(n47050), .B(n47049), .Z(n47053) );
  XOR U56527 ( .A(n47052), .B(n47051), .Z(n47049) );
  XOR U56528 ( .A(y[1124]), .B(x[1124]), .Z(n47051) );
  XOR U56529 ( .A(y[1123]), .B(x[1123]), .Z(n47052) );
  XOR U56530 ( .A(y[1122]), .B(x[1122]), .Z(n47050) );
  XOR U56531 ( .A(n47044), .B(n47043), .Z(n47054) );
  XOR U56532 ( .A(n47046), .B(n47045), .Z(n47043) );
  XOR U56533 ( .A(y[1121]), .B(x[1121]), .Z(n47045) );
  XOR U56534 ( .A(y[1120]), .B(x[1120]), .Z(n47046) );
  XOR U56535 ( .A(y[1119]), .B(x[1119]), .Z(n47044) );
  NAND U56536 ( .A(n47107), .B(n47108), .Z(N61194) );
  NAND U56537 ( .A(n47109), .B(n47110), .Z(n47108) );
  NANDN U56538 ( .A(n47111), .B(n47112), .Z(n47110) );
  NANDN U56539 ( .A(n47112), .B(n47111), .Z(n47107) );
  XOR U56540 ( .A(n47111), .B(n47113), .Z(N61193) );
  XNOR U56541 ( .A(n47109), .B(n47112), .Z(n47113) );
  NAND U56542 ( .A(n47114), .B(n47115), .Z(n47112) );
  NAND U56543 ( .A(n47116), .B(n47117), .Z(n47115) );
  NANDN U56544 ( .A(n47118), .B(n47119), .Z(n47117) );
  NANDN U56545 ( .A(n47119), .B(n47118), .Z(n47114) );
  AND U56546 ( .A(n47120), .B(n47121), .Z(n47109) );
  NAND U56547 ( .A(n47122), .B(n47123), .Z(n47121) );
  NANDN U56548 ( .A(n47124), .B(n47125), .Z(n47123) );
  NANDN U56549 ( .A(n47125), .B(n47124), .Z(n47120) );
  IV U56550 ( .A(n47126), .Z(n47125) );
  AND U56551 ( .A(n47127), .B(n47128), .Z(n47111) );
  NAND U56552 ( .A(n47129), .B(n47130), .Z(n47128) );
  NANDN U56553 ( .A(n47131), .B(n47132), .Z(n47130) );
  NANDN U56554 ( .A(n47132), .B(n47131), .Z(n47127) );
  XOR U56555 ( .A(n47124), .B(n47133), .Z(N61192) );
  XNOR U56556 ( .A(n47122), .B(n47126), .Z(n47133) );
  XOR U56557 ( .A(n47119), .B(n47134), .Z(n47126) );
  XNOR U56558 ( .A(n47116), .B(n47118), .Z(n47134) );
  AND U56559 ( .A(n47135), .B(n47136), .Z(n47118) );
  NANDN U56560 ( .A(n47137), .B(n47138), .Z(n47136) );
  OR U56561 ( .A(n47139), .B(n47140), .Z(n47138) );
  IV U56562 ( .A(n47141), .Z(n47140) );
  NANDN U56563 ( .A(n47141), .B(n47139), .Z(n47135) );
  AND U56564 ( .A(n47142), .B(n47143), .Z(n47116) );
  NAND U56565 ( .A(n47144), .B(n47145), .Z(n47143) );
  NANDN U56566 ( .A(n47146), .B(n47147), .Z(n47145) );
  NANDN U56567 ( .A(n47147), .B(n47146), .Z(n47142) );
  IV U56568 ( .A(n47148), .Z(n47147) );
  NAND U56569 ( .A(n47149), .B(n47150), .Z(n47119) );
  NANDN U56570 ( .A(n47151), .B(n47152), .Z(n47150) );
  NANDN U56571 ( .A(n47153), .B(n47154), .Z(n47152) );
  NANDN U56572 ( .A(n47154), .B(n47153), .Z(n47149) );
  IV U56573 ( .A(n47155), .Z(n47153) );
  AND U56574 ( .A(n47156), .B(n47157), .Z(n47122) );
  NAND U56575 ( .A(n47158), .B(n47159), .Z(n47157) );
  NANDN U56576 ( .A(n47160), .B(n47161), .Z(n47159) );
  NANDN U56577 ( .A(n47161), .B(n47160), .Z(n47156) );
  XOR U56578 ( .A(n47132), .B(n47162), .Z(n47124) );
  XNOR U56579 ( .A(n47129), .B(n47131), .Z(n47162) );
  AND U56580 ( .A(n47163), .B(n47164), .Z(n47131) );
  NANDN U56581 ( .A(n47165), .B(n47166), .Z(n47164) );
  OR U56582 ( .A(n47167), .B(n47168), .Z(n47166) );
  IV U56583 ( .A(n47169), .Z(n47168) );
  NANDN U56584 ( .A(n47169), .B(n47167), .Z(n47163) );
  AND U56585 ( .A(n47170), .B(n47171), .Z(n47129) );
  NAND U56586 ( .A(n47172), .B(n47173), .Z(n47171) );
  NANDN U56587 ( .A(n47174), .B(n47175), .Z(n47173) );
  NANDN U56588 ( .A(n47175), .B(n47174), .Z(n47170) );
  IV U56589 ( .A(n47176), .Z(n47175) );
  NAND U56590 ( .A(n47177), .B(n47178), .Z(n47132) );
  NANDN U56591 ( .A(n47179), .B(n47180), .Z(n47178) );
  NANDN U56592 ( .A(n47181), .B(n47182), .Z(n47180) );
  NANDN U56593 ( .A(n47182), .B(n47181), .Z(n47177) );
  IV U56594 ( .A(n47183), .Z(n47181) );
  XOR U56595 ( .A(n47158), .B(n47184), .Z(N61191) );
  XNOR U56596 ( .A(n47161), .B(n47160), .Z(n47184) );
  XNOR U56597 ( .A(n47172), .B(n47185), .Z(n47160) );
  XNOR U56598 ( .A(n47176), .B(n47174), .Z(n47185) );
  XOR U56599 ( .A(n47182), .B(n47186), .Z(n47174) );
  XNOR U56600 ( .A(n47179), .B(n47183), .Z(n47186) );
  AND U56601 ( .A(n47187), .B(n47188), .Z(n47183) );
  NAND U56602 ( .A(n47189), .B(n47190), .Z(n47188) );
  NAND U56603 ( .A(n47191), .B(n47192), .Z(n47187) );
  AND U56604 ( .A(n47193), .B(n47194), .Z(n47179) );
  NAND U56605 ( .A(n47195), .B(n47196), .Z(n47194) );
  NAND U56606 ( .A(n47197), .B(n47198), .Z(n47193) );
  NANDN U56607 ( .A(n47199), .B(n47200), .Z(n47182) );
  ANDN U56608 ( .B(n47201), .A(n47202), .Z(n47176) );
  XNOR U56609 ( .A(n47167), .B(n47203), .Z(n47172) );
  XNOR U56610 ( .A(n47165), .B(n47169), .Z(n47203) );
  AND U56611 ( .A(n47204), .B(n47205), .Z(n47169) );
  NAND U56612 ( .A(n47206), .B(n47207), .Z(n47205) );
  NAND U56613 ( .A(n47208), .B(n47209), .Z(n47204) );
  AND U56614 ( .A(n47210), .B(n47211), .Z(n47165) );
  NAND U56615 ( .A(n47212), .B(n47213), .Z(n47211) );
  NAND U56616 ( .A(n47214), .B(n47215), .Z(n47210) );
  AND U56617 ( .A(n47216), .B(n47217), .Z(n47167) );
  NAND U56618 ( .A(n47218), .B(n47219), .Z(n47161) );
  XNOR U56619 ( .A(n47144), .B(n47220), .Z(n47158) );
  XNOR U56620 ( .A(n47148), .B(n47146), .Z(n47220) );
  XOR U56621 ( .A(n47154), .B(n47221), .Z(n47146) );
  XNOR U56622 ( .A(n47151), .B(n47155), .Z(n47221) );
  AND U56623 ( .A(n47222), .B(n47223), .Z(n47155) );
  NAND U56624 ( .A(n47224), .B(n47225), .Z(n47223) );
  NAND U56625 ( .A(n47226), .B(n47227), .Z(n47222) );
  AND U56626 ( .A(n47228), .B(n47229), .Z(n47151) );
  NAND U56627 ( .A(n47230), .B(n47231), .Z(n47229) );
  NAND U56628 ( .A(n47232), .B(n47233), .Z(n47228) );
  NANDN U56629 ( .A(n47234), .B(n47235), .Z(n47154) );
  ANDN U56630 ( .B(n47236), .A(n47237), .Z(n47148) );
  XNOR U56631 ( .A(n47139), .B(n47238), .Z(n47144) );
  XNOR U56632 ( .A(n47137), .B(n47141), .Z(n47238) );
  AND U56633 ( .A(n47239), .B(n47240), .Z(n47141) );
  NAND U56634 ( .A(n47241), .B(n47242), .Z(n47240) );
  NAND U56635 ( .A(n47243), .B(n47244), .Z(n47239) );
  AND U56636 ( .A(n47245), .B(n47246), .Z(n47137) );
  NAND U56637 ( .A(n47247), .B(n47248), .Z(n47246) );
  NAND U56638 ( .A(n47249), .B(n47250), .Z(n47245) );
  AND U56639 ( .A(n47251), .B(n47252), .Z(n47139) );
  XOR U56640 ( .A(n47219), .B(n47218), .Z(N61190) );
  XNOR U56641 ( .A(n47236), .B(n47237), .Z(n47218) );
  XNOR U56642 ( .A(n47251), .B(n47252), .Z(n47237) );
  XOR U56643 ( .A(n47248), .B(n47247), .Z(n47252) );
  XOR U56644 ( .A(y[1116]), .B(x[1116]), .Z(n47247) );
  XOR U56645 ( .A(n47250), .B(n47249), .Z(n47248) );
  XOR U56646 ( .A(y[1118]), .B(x[1118]), .Z(n47249) );
  XOR U56647 ( .A(y[1117]), .B(x[1117]), .Z(n47250) );
  XOR U56648 ( .A(n47242), .B(n47241), .Z(n47251) );
  XOR U56649 ( .A(n47244), .B(n47243), .Z(n47241) );
  XOR U56650 ( .A(y[1115]), .B(x[1115]), .Z(n47243) );
  XOR U56651 ( .A(y[1114]), .B(x[1114]), .Z(n47244) );
  XOR U56652 ( .A(y[1113]), .B(x[1113]), .Z(n47242) );
  XNOR U56653 ( .A(n47235), .B(n47234), .Z(n47236) );
  XNOR U56654 ( .A(n47231), .B(n47230), .Z(n47234) );
  XOR U56655 ( .A(n47233), .B(n47232), .Z(n47230) );
  XOR U56656 ( .A(y[1112]), .B(x[1112]), .Z(n47232) );
  XOR U56657 ( .A(y[1111]), .B(x[1111]), .Z(n47233) );
  XOR U56658 ( .A(y[1110]), .B(x[1110]), .Z(n47231) );
  XOR U56659 ( .A(n47225), .B(n47224), .Z(n47235) );
  XOR U56660 ( .A(n47227), .B(n47226), .Z(n47224) );
  XOR U56661 ( .A(y[1109]), .B(x[1109]), .Z(n47226) );
  XOR U56662 ( .A(y[1108]), .B(x[1108]), .Z(n47227) );
  XOR U56663 ( .A(y[1107]), .B(x[1107]), .Z(n47225) );
  XNOR U56664 ( .A(n47201), .B(n47202), .Z(n47219) );
  XNOR U56665 ( .A(n47216), .B(n47217), .Z(n47202) );
  XOR U56666 ( .A(n47213), .B(n47212), .Z(n47217) );
  XOR U56667 ( .A(y[1104]), .B(x[1104]), .Z(n47212) );
  XOR U56668 ( .A(n47215), .B(n47214), .Z(n47213) );
  XOR U56669 ( .A(y[1106]), .B(x[1106]), .Z(n47214) );
  XOR U56670 ( .A(y[1105]), .B(x[1105]), .Z(n47215) );
  XOR U56671 ( .A(n47207), .B(n47206), .Z(n47216) );
  XOR U56672 ( .A(n47209), .B(n47208), .Z(n47206) );
  XOR U56673 ( .A(y[1103]), .B(x[1103]), .Z(n47208) );
  XOR U56674 ( .A(y[1102]), .B(x[1102]), .Z(n47209) );
  XOR U56675 ( .A(y[1101]), .B(x[1101]), .Z(n47207) );
  XNOR U56676 ( .A(n47200), .B(n47199), .Z(n47201) );
  XNOR U56677 ( .A(n47196), .B(n47195), .Z(n47199) );
  XOR U56678 ( .A(n47198), .B(n47197), .Z(n47195) );
  XOR U56679 ( .A(y[1100]), .B(x[1100]), .Z(n47197) );
  XOR U56680 ( .A(y[1099]), .B(x[1099]), .Z(n47198) );
  XOR U56681 ( .A(y[1098]), .B(x[1098]), .Z(n47196) );
  XOR U56682 ( .A(n47190), .B(n47189), .Z(n47200) );
  XOR U56683 ( .A(n47192), .B(n47191), .Z(n47189) );
  XOR U56684 ( .A(y[1097]), .B(x[1097]), .Z(n47191) );
  XOR U56685 ( .A(y[1096]), .B(x[1096]), .Z(n47192) );
  XOR U56686 ( .A(y[1095]), .B(x[1095]), .Z(n47190) );
  NAND U56687 ( .A(n47253), .B(n47254), .Z(N61181) );
  NAND U56688 ( .A(n47255), .B(n47256), .Z(n47254) );
  NANDN U56689 ( .A(n47257), .B(n47258), .Z(n47256) );
  NANDN U56690 ( .A(n47258), .B(n47257), .Z(n47253) );
  XOR U56691 ( .A(n47257), .B(n47259), .Z(N61180) );
  XNOR U56692 ( .A(n47255), .B(n47258), .Z(n47259) );
  NAND U56693 ( .A(n47260), .B(n47261), .Z(n47258) );
  NAND U56694 ( .A(n47262), .B(n47263), .Z(n47261) );
  NANDN U56695 ( .A(n47264), .B(n47265), .Z(n47263) );
  NANDN U56696 ( .A(n47265), .B(n47264), .Z(n47260) );
  AND U56697 ( .A(n47266), .B(n47267), .Z(n47255) );
  NAND U56698 ( .A(n47268), .B(n47269), .Z(n47267) );
  NANDN U56699 ( .A(n47270), .B(n47271), .Z(n47269) );
  NANDN U56700 ( .A(n47271), .B(n47270), .Z(n47266) );
  IV U56701 ( .A(n47272), .Z(n47271) );
  AND U56702 ( .A(n47273), .B(n47274), .Z(n47257) );
  NAND U56703 ( .A(n47275), .B(n47276), .Z(n47274) );
  NANDN U56704 ( .A(n47277), .B(n47278), .Z(n47276) );
  NANDN U56705 ( .A(n47278), .B(n47277), .Z(n47273) );
  XOR U56706 ( .A(n47270), .B(n47279), .Z(N61179) );
  XNOR U56707 ( .A(n47268), .B(n47272), .Z(n47279) );
  XOR U56708 ( .A(n47265), .B(n47280), .Z(n47272) );
  XNOR U56709 ( .A(n47262), .B(n47264), .Z(n47280) );
  AND U56710 ( .A(n47281), .B(n47282), .Z(n47264) );
  NANDN U56711 ( .A(n47283), .B(n47284), .Z(n47282) );
  OR U56712 ( .A(n47285), .B(n47286), .Z(n47284) );
  IV U56713 ( .A(n47287), .Z(n47286) );
  NANDN U56714 ( .A(n47287), .B(n47285), .Z(n47281) );
  AND U56715 ( .A(n47288), .B(n47289), .Z(n47262) );
  NAND U56716 ( .A(n47290), .B(n47291), .Z(n47289) );
  NANDN U56717 ( .A(n47292), .B(n47293), .Z(n47291) );
  NANDN U56718 ( .A(n47293), .B(n47292), .Z(n47288) );
  IV U56719 ( .A(n47294), .Z(n47293) );
  NAND U56720 ( .A(n47295), .B(n47296), .Z(n47265) );
  NANDN U56721 ( .A(n47297), .B(n47298), .Z(n47296) );
  NANDN U56722 ( .A(n47299), .B(n47300), .Z(n47298) );
  NANDN U56723 ( .A(n47300), .B(n47299), .Z(n47295) );
  IV U56724 ( .A(n47301), .Z(n47299) );
  AND U56725 ( .A(n47302), .B(n47303), .Z(n47268) );
  NAND U56726 ( .A(n47304), .B(n47305), .Z(n47303) );
  NANDN U56727 ( .A(n47306), .B(n47307), .Z(n47305) );
  NANDN U56728 ( .A(n47307), .B(n47306), .Z(n47302) );
  XOR U56729 ( .A(n47278), .B(n47308), .Z(n47270) );
  XNOR U56730 ( .A(n47275), .B(n47277), .Z(n47308) );
  AND U56731 ( .A(n47309), .B(n47310), .Z(n47277) );
  NANDN U56732 ( .A(n47311), .B(n47312), .Z(n47310) );
  OR U56733 ( .A(n47313), .B(n47314), .Z(n47312) );
  IV U56734 ( .A(n47315), .Z(n47314) );
  NANDN U56735 ( .A(n47315), .B(n47313), .Z(n47309) );
  AND U56736 ( .A(n47316), .B(n47317), .Z(n47275) );
  NAND U56737 ( .A(n47318), .B(n47319), .Z(n47317) );
  NANDN U56738 ( .A(n47320), .B(n47321), .Z(n47319) );
  NANDN U56739 ( .A(n47321), .B(n47320), .Z(n47316) );
  IV U56740 ( .A(n47322), .Z(n47321) );
  NAND U56741 ( .A(n47323), .B(n47324), .Z(n47278) );
  NANDN U56742 ( .A(n47325), .B(n47326), .Z(n47324) );
  NANDN U56743 ( .A(n47327), .B(n47328), .Z(n47326) );
  NANDN U56744 ( .A(n47328), .B(n47327), .Z(n47323) );
  IV U56745 ( .A(n47329), .Z(n47327) );
  XOR U56746 ( .A(n47304), .B(n47330), .Z(N61178) );
  XNOR U56747 ( .A(n47307), .B(n47306), .Z(n47330) );
  XNOR U56748 ( .A(n47318), .B(n47331), .Z(n47306) );
  XNOR U56749 ( .A(n47322), .B(n47320), .Z(n47331) );
  XOR U56750 ( .A(n47328), .B(n47332), .Z(n47320) );
  XNOR U56751 ( .A(n47325), .B(n47329), .Z(n47332) );
  AND U56752 ( .A(n47333), .B(n47334), .Z(n47329) );
  NAND U56753 ( .A(n47335), .B(n47336), .Z(n47334) );
  NAND U56754 ( .A(n47337), .B(n47338), .Z(n47333) );
  AND U56755 ( .A(n47339), .B(n47340), .Z(n47325) );
  NAND U56756 ( .A(n47341), .B(n47342), .Z(n47340) );
  NAND U56757 ( .A(n47343), .B(n47344), .Z(n47339) );
  NANDN U56758 ( .A(n47345), .B(n47346), .Z(n47328) );
  ANDN U56759 ( .B(n47347), .A(n47348), .Z(n47322) );
  XNOR U56760 ( .A(n47313), .B(n47349), .Z(n47318) );
  XNOR U56761 ( .A(n47311), .B(n47315), .Z(n47349) );
  AND U56762 ( .A(n47350), .B(n47351), .Z(n47315) );
  NAND U56763 ( .A(n47352), .B(n47353), .Z(n47351) );
  NAND U56764 ( .A(n47354), .B(n47355), .Z(n47350) );
  AND U56765 ( .A(n47356), .B(n47357), .Z(n47311) );
  NAND U56766 ( .A(n47358), .B(n47359), .Z(n47357) );
  NAND U56767 ( .A(n47360), .B(n47361), .Z(n47356) );
  AND U56768 ( .A(n47362), .B(n47363), .Z(n47313) );
  NAND U56769 ( .A(n47364), .B(n47365), .Z(n47307) );
  XNOR U56770 ( .A(n47290), .B(n47366), .Z(n47304) );
  XNOR U56771 ( .A(n47294), .B(n47292), .Z(n47366) );
  XOR U56772 ( .A(n47300), .B(n47367), .Z(n47292) );
  XNOR U56773 ( .A(n47297), .B(n47301), .Z(n47367) );
  AND U56774 ( .A(n47368), .B(n47369), .Z(n47301) );
  NAND U56775 ( .A(n47370), .B(n47371), .Z(n47369) );
  NAND U56776 ( .A(n47372), .B(n47373), .Z(n47368) );
  AND U56777 ( .A(n47374), .B(n47375), .Z(n47297) );
  NAND U56778 ( .A(n47376), .B(n47377), .Z(n47375) );
  NAND U56779 ( .A(n47378), .B(n47379), .Z(n47374) );
  NANDN U56780 ( .A(n47380), .B(n47381), .Z(n47300) );
  ANDN U56781 ( .B(n47382), .A(n47383), .Z(n47294) );
  XNOR U56782 ( .A(n47285), .B(n47384), .Z(n47290) );
  XNOR U56783 ( .A(n47283), .B(n47287), .Z(n47384) );
  AND U56784 ( .A(n47385), .B(n47386), .Z(n47287) );
  NAND U56785 ( .A(n47387), .B(n47388), .Z(n47386) );
  NAND U56786 ( .A(n47389), .B(n47390), .Z(n47385) );
  AND U56787 ( .A(n47391), .B(n47392), .Z(n47283) );
  NAND U56788 ( .A(n47393), .B(n47394), .Z(n47392) );
  NAND U56789 ( .A(n47395), .B(n47396), .Z(n47391) );
  AND U56790 ( .A(n47397), .B(n47398), .Z(n47285) );
  XOR U56791 ( .A(n47365), .B(n47364), .Z(N61177) );
  XNOR U56792 ( .A(n47382), .B(n47383), .Z(n47364) );
  XNOR U56793 ( .A(n47397), .B(n47398), .Z(n47383) );
  XOR U56794 ( .A(n47394), .B(n47393), .Z(n47398) );
  XOR U56795 ( .A(y[1092]), .B(x[1092]), .Z(n47393) );
  XOR U56796 ( .A(n47396), .B(n47395), .Z(n47394) );
  XOR U56797 ( .A(y[1094]), .B(x[1094]), .Z(n47395) );
  XOR U56798 ( .A(y[1093]), .B(x[1093]), .Z(n47396) );
  XOR U56799 ( .A(n47388), .B(n47387), .Z(n47397) );
  XOR U56800 ( .A(n47390), .B(n47389), .Z(n47387) );
  XOR U56801 ( .A(y[1091]), .B(x[1091]), .Z(n47389) );
  XOR U56802 ( .A(y[1090]), .B(x[1090]), .Z(n47390) );
  XOR U56803 ( .A(y[1089]), .B(x[1089]), .Z(n47388) );
  XNOR U56804 ( .A(n47381), .B(n47380), .Z(n47382) );
  XNOR U56805 ( .A(n47377), .B(n47376), .Z(n47380) );
  XOR U56806 ( .A(n47379), .B(n47378), .Z(n47376) );
  XOR U56807 ( .A(y[1088]), .B(x[1088]), .Z(n47378) );
  XOR U56808 ( .A(y[1087]), .B(x[1087]), .Z(n47379) );
  XOR U56809 ( .A(y[1086]), .B(x[1086]), .Z(n47377) );
  XOR U56810 ( .A(n47371), .B(n47370), .Z(n47381) );
  XOR U56811 ( .A(n47373), .B(n47372), .Z(n47370) );
  XOR U56812 ( .A(y[1085]), .B(x[1085]), .Z(n47372) );
  XOR U56813 ( .A(y[1084]), .B(x[1084]), .Z(n47373) );
  XOR U56814 ( .A(y[1083]), .B(x[1083]), .Z(n47371) );
  XNOR U56815 ( .A(n47347), .B(n47348), .Z(n47365) );
  XNOR U56816 ( .A(n47362), .B(n47363), .Z(n47348) );
  XOR U56817 ( .A(n47359), .B(n47358), .Z(n47363) );
  XOR U56818 ( .A(y[1080]), .B(x[1080]), .Z(n47358) );
  XOR U56819 ( .A(n47361), .B(n47360), .Z(n47359) );
  XOR U56820 ( .A(y[1082]), .B(x[1082]), .Z(n47360) );
  XOR U56821 ( .A(y[1081]), .B(x[1081]), .Z(n47361) );
  XOR U56822 ( .A(n47353), .B(n47352), .Z(n47362) );
  XOR U56823 ( .A(n47355), .B(n47354), .Z(n47352) );
  XOR U56824 ( .A(y[1079]), .B(x[1079]), .Z(n47354) );
  XOR U56825 ( .A(y[1078]), .B(x[1078]), .Z(n47355) );
  XOR U56826 ( .A(y[1077]), .B(x[1077]), .Z(n47353) );
  XNOR U56827 ( .A(n47346), .B(n47345), .Z(n47347) );
  XNOR U56828 ( .A(n47342), .B(n47341), .Z(n47345) );
  XOR U56829 ( .A(n47344), .B(n47343), .Z(n47341) );
  XOR U56830 ( .A(y[1076]), .B(x[1076]), .Z(n47343) );
  XOR U56831 ( .A(y[1075]), .B(x[1075]), .Z(n47344) );
  XOR U56832 ( .A(y[1074]), .B(x[1074]), .Z(n47342) );
  XOR U56833 ( .A(n47336), .B(n47335), .Z(n47346) );
  XOR U56834 ( .A(n47338), .B(n47337), .Z(n47335) );
  XOR U56835 ( .A(y[1073]), .B(x[1073]), .Z(n47337) );
  XOR U56836 ( .A(y[1072]), .B(x[1072]), .Z(n47338) );
  XOR U56837 ( .A(y[1071]), .B(x[1071]), .Z(n47336) );
  NAND U56838 ( .A(n47399), .B(n47400), .Z(N61168) );
  NAND U56839 ( .A(n47401), .B(n47402), .Z(n47400) );
  NANDN U56840 ( .A(n47403), .B(n47404), .Z(n47402) );
  NANDN U56841 ( .A(n47404), .B(n47403), .Z(n47399) );
  XOR U56842 ( .A(n47403), .B(n47405), .Z(N61167) );
  XNOR U56843 ( .A(n47401), .B(n47404), .Z(n47405) );
  NAND U56844 ( .A(n47406), .B(n47407), .Z(n47404) );
  NAND U56845 ( .A(n47408), .B(n47409), .Z(n47407) );
  NANDN U56846 ( .A(n47410), .B(n47411), .Z(n47409) );
  NANDN U56847 ( .A(n47411), .B(n47410), .Z(n47406) );
  AND U56848 ( .A(n47412), .B(n47413), .Z(n47401) );
  NAND U56849 ( .A(n47414), .B(n47415), .Z(n47413) );
  NANDN U56850 ( .A(n47416), .B(n47417), .Z(n47415) );
  NANDN U56851 ( .A(n47417), .B(n47416), .Z(n47412) );
  IV U56852 ( .A(n47418), .Z(n47417) );
  AND U56853 ( .A(n47419), .B(n47420), .Z(n47403) );
  NAND U56854 ( .A(n47421), .B(n47422), .Z(n47420) );
  NANDN U56855 ( .A(n47423), .B(n47424), .Z(n47422) );
  NANDN U56856 ( .A(n47424), .B(n47423), .Z(n47419) );
  XOR U56857 ( .A(n47416), .B(n47425), .Z(N61166) );
  XNOR U56858 ( .A(n47414), .B(n47418), .Z(n47425) );
  XOR U56859 ( .A(n47411), .B(n47426), .Z(n47418) );
  XNOR U56860 ( .A(n47408), .B(n47410), .Z(n47426) );
  AND U56861 ( .A(n47427), .B(n47428), .Z(n47410) );
  NANDN U56862 ( .A(n47429), .B(n47430), .Z(n47428) );
  OR U56863 ( .A(n47431), .B(n47432), .Z(n47430) );
  IV U56864 ( .A(n47433), .Z(n47432) );
  NANDN U56865 ( .A(n47433), .B(n47431), .Z(n47427) );
  AND U56866 ( .A(n47434), .B(n47435), .Z(n47408) );
  NAND U56867 ( .A(n47436), .B(n47437), .Z(n47435) );
  NANDN U56868 ( .A(n47438), .B(n47439), .Z(n47437) );
  NANDN U56869 ( .A(n47439), .B(n47438), .Z(n47434) );
  IV U56870 ( .A(n47440), .Z(n47439) );
  NAND U56871 ( .A(n47441), .B(n47442), .Z(n47411) );
  NANDN U56872 ( .A(n47443), .B(n47444), .Z(n47442) );
  NANDN U56873 ( .A(n47445), .B(n47446), .Z(n47444) );
  NANDN U56874 ( .A(n47446), .B(n47445), .Z(n47441) );
  IV U56875 ( .A(n47447), .Z(n47445) );
  AND U56876 ( .A(n47448), .B(n47449), .Z(n47414) );
  NAND U56877 ( .A(n47450), .B(n47451), .Z(n47449) );
  NANDN U56878 ( .A(n47452), .B(n47453), .Z(n47451) );
  NANDN U56879 ( .A(n47453), .B(n47452), .Z(n47448) );
  XOR U56880 ( .A(n47424), .B(n47454), .Z(n47416) );
  XNOR U56881 ( .A(n47421), .B(n47423), .Z(n47454) );
  AND U56882 ( .A(n47455), .B(n47456), .Z(n47423) );
  NANDN U56883 ( .A(n47457), .B(n47458), .Z(n47456) );
  OR U56884 ( .A(n47459), .B(n47460), .Z(n47458) );
  IV U56885 ( .A(n47461), .Z(n47460) );
  NANDN U56886 ( .A(n47461), .B(n47459), .Z(n47455) );
  AND U56887 ( .A(n47462), .B(n47463), .Z(n47421) );
  NAND U56888 ( .A(n47464), .B(n47465), .Z(n47463) );
  NANDN U56889 ( .A(n47466), .B(n47467), .Z(n47465) );
  NANDN U56890 ( .A(n47467), .B(n47466), .Z(n47462) );
  IV U56891 ( .A(n47468), .Z(n47467) );
  NAND U56892 ( .A(n47469), .B(n47470), .Z(n47424) );
  NANDN U56893 ( .A(n47471), .B(n47472), .Z(n47470) );
  NANDN U56894 ( .A(n47473), .B(n47474), .Z(n47472) );
  NANDN U56895 ( .A(n47474), .B(n47473), .Z(n47469) );
  IV U56896 ( .A(n47475), .Z(n47473) );
  XOR U56897 ( .A(n47450), .B(n47476), .Z(N61165) );
  XNOR U56898 ( .A(n47453), .B(n47452), .Z(n47476) );
  XNOR U56899 ( .A(n47464), .B(n47477), .Z(n47452) );
  XNOR U56900 ( .A(n47468), .B(n47466), .Z(n47477) );
  XOR U56901 ( .A(n47474), .B(n47478), .Z(n47466) );
  XNOR U56902 ( .A(n47471), .B(n47475), .Z(n47478) );
  AND U56903 ( .A(n47479), .B(n47480), .Z(n47475) );
  NAND U56904 ( .A(n47481), .B(n47482), .Z(n47480) );
  NAND U56905 ( .A(n47483), .B(n47484), .Z(n47479) );
  AND U56906 ( .A(n47485), .B(n47486), .Z(n47471) );
  NAND U56907 ( .A(n47487), .B(n47488), .Z(n47486) );
  NAND U56908 ( .A(n47489), .B(n47490), .Z(n47485) );
  NANDN U56909 ( .A(n47491), .B(n47492), .Z(n47474) );
  ANDN U56910 ( .B(n47493), .A(n47494), .Z(n47468) );
  XNOR U56911 ( .A(n47459), .B(n47495), .Z(n47464) );
  XNOR U56912 ( .A(n47457), .B(n47461), .Z(n47495) );
  AND U56913 ( .A(n47496), .B(n47497), .Z(n47461) );
  NAND U56914 ( .A(n47498), .B(n47499), .Z(n47497) );
  NAND U56915 ( .A(n47500), .B(n47501), .Z(n47496) );
  AND U56916 ( .A(n47502), .B(n47503), .Z(n47457) );
  NAND U56917 ( .A(n47504), .B(n47505), .Z(n47503) );
  NAND U56918 ( .A(n47506), .B(n47507), .Z(n47502) );
  AND U56919 ( .A(n47508), .B(n47509), .Z(n47459) );
  NAND U56920 ( .A(n47510), .B(n47511), .Z(n47453) );
  XNOR U56921 ( .A(n47436), .B(n47512), .Z(n47450) );
  XNOR U56922 ( .A(n47440), .B(n47438), .Z(n47512) );
  XOR U56923 ( .A(n47446), .B(n47513), .Z(n47438) );
  XNOR U56924 ( .A(n47443), .B(n47447), .Z(n47513) );
  AND U56925 ( .A(n47514), .B(n47515), .Z(n47447) );
  NAND U56926 ( .A(n47516), .B(n47517), .Z(n47515) );
  NAND U56927 ( .A(n47518), .B(n47519), .Z(n47514) );
  AND U56928 ( .A(n47520), .B(n47521), .Z(n47443) );
  NAND U56929 ( .A(n47522), .B(n47523), .Z(n47521) );
  NAND U56930 ( .A(n47524), .B(n47525), .Z(n47520) );
  NANDN U56931 ( .A(n47526), .B(n47527), .Z(n47446) );
  ANDN U56932 ( .B(n47528), .A(n47529), .Z(n47440) );
  XNOR U56933 ( .A(n47431), .B(n47530), .Z(n47436) );
  XNOR U56934 ( .A(n47429), .B(n47433), .Z(n47530) );
  AND U56935 ( .A(n47531), .B(n47532), .Z(n47433) );
  NAND U56936 ( .A(n47533), .B(n47534), .Z(n47532) );
  NAND U56937 ( .A(n47535), .B(n47536), .Z(n47531) );
  AND U56938 ( .A(n47537), .B(n47538), .Z(n47429) );
  NAND U56939 ( .A(n47539), .B(n47540), .Z(n47538) );
  NAND U56940 ( .A(n47541), .B(n47542), .Z(n47537) );
  AND U56941 ( .A(n47543), .B(n47544), .Z(n47431) );
  XOR U56942 ( .A(n47511), .B(n47510), .Z(N61164) );
  XNOR U56943 ( .A(n47528), .B(n47529), .Z(n47510) );
  XNOR U56944 ( .A(n47543), .B(n47544), .Z(n47529) );
  XOR U56945 ( .A(n47540), .B(n47539), .Z(n47544) );
  XOR U56946 ( .A(y[1068]), .B(x[1068]), .Z(n47539) );
  XOR U56947 ( .A(n47542), .B(n47541), .Z(n47540) );
  XOR U56948 ( .A(y[1070]), .B(x[1070]), .Z(n47541) );
  XOR U56949 ( .A(y[1069]), .B(x[1069]), .Z(n47542) );
  XOR U56950 ( .A(n47534), .B(n47533), .Z(n47543) );
  XOR U56951 ( .A(n47536), .B(n47535), .Z(n47533) );
  XOR U56952 ( .A(y[1067]), .B(x[1067]), .Z(n47535) );
  XOR U56953 ( .A(y[1066]), .B(x[1066]), .Z(n47536) );
  XOR U56954 ( .A(y[1065]), .B(x[1065]), .Z(n47534) );
  XNOR U56955 ( .A(n47527), .B(n47526), .Z(n47528) );
  XNOR U56956 ( .A(n47523), .B(n47522), .Z(n47526) );
  XOR U56957 ( .A(n47525), .B(n47524), .Z(n47522) );
  XOR U56958 ( .A(y[1064]), .B(x[1064]), .Z(n47524) );
  XOR U56959 ( .A(y[1063]), .B(x[1063]), .Z(n47525) );
  XOR U56960 ( .A(y[1062]), .B(x[1062]), .Z(n47523) );
  XOR U56961 ( .A(n47517), .B(n47516), .Z(n47527) );
  XOR U56962 ( .A(n47519), .B(n47518), .Z(n47516) );
  XOR U56963 ( .A(y[1061]), .B(x[1061]), .Z(n47518) );
  XOR U56964 ( .A(y[1060]), .B(x[1060]), .Z(n47519) );
  XOR U56965 ( .A(y[1059]), .B(x[1059]), .Z(n47517) );
  XNOR U56966 ( .A(n47493), .B(n47494), .Z(n47511) );
  XNOR U56967 ( .A(n47508), .B(n47509), .Z(n47494) );
  XOR U56968 ( .A(n47505), .B(n47504), .Z(n47509) );
  XOR U56969 ( .A(y[1056]), .B(x[1056]), .Z(n47504) );
  XOR U56970 ( .A(n47507), .B(n47506), .Z(n47505) );
  XOR U56971 ( .A(y[1058]), .B(x[1058]), .Z(n47506) );
  XOR U56972 ( .A(y[1057]), .B(x[1057]), .Z(n47507) );
  XOR U56973 ( .A(n47499), .B(n47498), .Z(n47508) );
  XOR U56974 ( .A(n47501), .B(n47500), .Z(n47498) );
  XOR U56975 ( .A(y[1055]), .B(x[1055]), .Z(n47500) );
  XOR U56976 ( .A(y[1054]), .B(x[1054]), .Z(n47501) );
  XOR U56977 ( .A(y[1053]), .B(x[1053]), .Z(n47499) );
  XNOR U56978 ( .A(n47492), .B(n47491), .Z(n47493) );
  XNOR U56979 ( .A(n47488), .B(n47487), .Z(n47491) );
  XOR U56980 ( .A(n47490), .B(n47489), .Z(n47487) );
  XOR U56981 ( .A(y[1052]), .B(x[1052]), .Z(n47489) );
  XOR U56982 ( .A(y[1051]), .B(x[1051]), .Z(n47490) );
  XOR U56983 ( .A(y[1050]), .B(x[1050]), .Z(n47488) );
  XOR U56984 ( .A(n47482), .B(n47481), .Z(n47492) );
  XOR U56985 ( .A(n47484), .B(n47483), .Z(n47481) );
  XOR U56986 ( .A(y[1049]), .B(x[1049]), .Z(n47483) );
  XOR U56987 ( .A(y[1048]), .B(x[1048]), .Z(n47484) );
  XOR U56988 ( .A(y[1047]), .B(x[1047]), .Z(n47482) );
  NAND U56989 ( .A(n47545), .B(n47546), .Z(N61155) );
  NAND U56990 ( .A(n47547), .B(n47548), .Z(n47546) );
  NANDN U56991 ( .A(n47549), .B(n47550), .Z(n47548) );
  NANDN U56992 ( .A(n47550), .B(n47549), .Z(n47545) );
  XOR U56993 ( .A(n47549), .B(n47551), .Z(N61154) );
  XNOR U56994 ( .A(n47547), .B(n47550), .Z(n47551) );
  NAND U56995 ( .A(n47552), .B(n47553), .Z(n47550) );
  NAND U56996 ( .A(n47554), .B(n47555), .Z(n47553) );
  NANDN U56997 ( .A(n47556), .B(n47557), .Z(n47555) );
  NANDN U56998 ( .A(n47557), .B(n47556), .Z(n47552) );
  AND U56999 ( .A(n47558), .B(n47559), .Z(n47547) );
  NAND U57000 ( .A(n47560), .B(n47561), .Z(n47559) );
  NANDN U57001 ( .A(n47562), .B(n47563), .Z(n47561) );
  NANDN U57002 ( .A(n47563), .B(n47562), .Z(n47558) );
  IV U57003 ( .A(n47564), .Z(n47563) );
  AND U57004 ( .A(n47565), .B(n47566), .Z(n47549) );
  NAND U57005 ( .A(n47567), .B(n47568), .Z(n47566) );
  NANDN U57006 ( .A(n47569), .B(n47570), .Z(n47568) );
  NANDN U57007 ( .A(n47570), .B(n47569), .Z(n47565) );
  XOR U57008 ( .A(n47562), .B(n47571), .Z(N61153) );
  XNOR U57009 ( .A(n47560), .B(n47564), .Z(n47571) );
  XOR U57010 ( .A(n47557), .B(n47572), .Z(n47564) );
  XNOR U57011 ( .A(n47554), .B(n47556), .Z(n47572) );
  AND U57012 ( .A(n47573), .B(n47574), .Z(n47556) );
  NANDN U57013 ( .A(n47575), .B(n47576), .Z(n47574) );
  OR U57014 ( .A(n47577), .B(n47578), .Z(n47576) );
  IV U57015 ( .A(n47579), .Z(n47578) );
  NANDN U57016 ( .A(n47579), .B(n47577), .Z(n47573) );
  AND U57017 ( .A(n47580), .B(n47581), .Z(n47554) );
  NAND U57018 ( .A(n47582), .B(n47583), .Z(n47581) );
  NANDN U57019 ( .A(n47584), .B(n47585), .Z(n47583) );
  NANDN U57020 ( .A(n47585), .B(n47584), .Z(n47580) );
  IV U57021 ( .A(n47586), .Z(n47585) );
  NAND U57022 ( .A(n47587), .B(n47588), .Z(n47557) );
  NANDN U57023 ( .A(n47589), .B(n47590), .Z(n47588) );
  NANDN U57024 ( .A(n47591), .B(n47592), .Z(n47590) );
  NANDN U57025 ( .A(n47592), .B(n47591), .Z(n47587) );
  IV U57026 ( .A(n47593), .Z(n47591) );
  AND U57027 ( .A(n47594), .B(n47595), .Z(n47560) );
  NAND U57028 ( .A(n47596), .B(n47597), .Z(n47595) );
  NANDN U57029 ( .A(n47598), .B(n47599), .Z(n47597) );
  NANDN U57030 ( .A(n47599), .B(n47598), .Z(n47594) );
  XOR U57031 ( .A(n47570), .B(n47600), .Z(n47562) );
  XNOR U57032 ( .A(n47567), .B(n47569), .Z(n47600) );
  AND U57033 ( .A(n47601), .B(n47602), .Z(n47569) );
  NANDN U57034 ( .A(n47603), .B(n47604), .Z(n47602) );
  OR U57035 ( .A(n47605), .B(n47606), .Z(n47604) );
  IV U57036 ( .A(n47607), .Z(n47606) );
  NANDN U57037 ( .A(n47607), .B(n47605), .Z(n47601) );
  AND U57038 ( .A(n47608), .B(n47609), .Z(n47567) );
  NAND U57039 ( .A(n47610), .B(n47611), .Z(n47609) );
  NANDN U57040 ( .A(n47612), .B(n47613), .Z(n47611) );
  NANDN U57041 ( .A(n47613), .B(n47612), .Z(n47608) );
  IV U57042 ( .A(n47614), .Z(n47613) );
  NAND U57043 ( .A(n47615), .B(n47616), .Z(n47570) );
  NANDN U57044 ( .A(n47617), .B(n47618), .Z(n47616) );
  NANDN U57045 ( .A(n47619), .B(n47620), .Z(n47618) );
  NANDN U57046 ( .A(n47620), .B(n47619), .Z(n47615) );
  IV U57047 ( .A(n47621), .Z(n47619) );
  XOR U57048 ( .A(n47596), .B(n47622), .Z(N61152) );
  XNOR U57049 ( .A(n47599), .B(n47598), .Z(n47622) );
  XNOR U57050 ( .A(n47610), .B(n47623), .Z(n47598) );
  XNOR U57051 ( .A(n47614), .B(n47612), .Z(n47623) );
  XOR U57052 ( .A(n47620), .B(n47624), .Z(n47612) );
  XNOR U57053 ( .A(n47617), .B(n47621), .Z(n47624) );
  AND U57054 ( .A(n47625), .B(n47626), .Z(n47621) );
  NAND U57055 ( .A(n47627), .B(n47628), .Z(n47626) );
  NAND U57056 ( .A(n47629), .B(n47630), .Z(n47625) );
  AND U57057 ( .A(n47631), .B(n47632), .Z(n47617) );
  NAND U57058 ( .A(n47633), .B(n47634), .Z(n47632) );
  NAND U57059 ( .A(n47635), .B(n47636), .Z(n47631) );
  NANDN U57060 ( .A(n47637), .B(n47638), .Z(n47620) );
  ANDN U57061 ( .B(n47639), .A(n47640), .Z(n47614) );
  XNOR U57062 ( .A(n47605), .B(n47641), .Z(n47610) );
  XNOR U57063 ( .A(n47603), .B(n47607), .Z(n47641) );
  AND U57064 ( .A(n47642), .B(n47643), .Z(n47607) );
  NAND U57065 ( .A(n47644), .B(n47645), .Z(n47643) );
  NAND U57066 ( .A(n47646), .B(n47647), .Z(n47642) );
  AND U57067 ( .A(n47648), .B(n47649), .Z(n47603) );
  NAND U57068 ( .A(n47650), .B(n47651), .Z(n47649) );
  NAND U57069 ( .A(n47652), .B(n47653), .Z(n47648) );
  AND U57070 ( .A(n47654), .B(n47655), .Z(n47605) );
  NAND U57071 ( .A(n47656), .B(n47657), .Z(n47599) );
  XNOR U57072 ( .A(n47582), .B(n47658), .Z(n47596) );
  XNOR U57073 ( .A(n47586), .B(n47584), .Z(n47658) );
  XOR U57074 ( .A(n47592), .B(n47659), .Z(n47584) );
  XNOR U57075 ( .A(n47589), .B(n47593), .Z(n47659) );
  AND U57076 ( .A(n47660), .B(n47661), .Z(n47593) );
  NAND U57077 ( .A(n47662), .B(n47663), .Z(n47661) );
  NAND U57078 ( .A(n47664), .B(n47665), .Z(n47660) );
  AND U57079 ( .A(n47666), .B(n47667), .Z(n47589) );
  NAND U57080 ( .A(n47668), .B(n47669), .Z(n47667) );
  NAND U57081 ( .A(n47670), .B(n47671), .Z(n47666) );
  NANDN U57082 ( .A(n47672), .B(n47673), .Z(n47592) );
  ANDN U57083 ( .B(n47674), .A(n47675), .Z(n47586) );
  XNOR U57084 ( .A(n47577), .B(n47676), .Z(n47582) );
  XNOR U57085 ( .A(n47575), .B(n47579), .Z(n47676) );
  AND U57086 ( .A(n47677), .B(n47678), .Z(n47579) );
  NAND U57087 ( .A(n47679), .B(n47680), .Z(n47678) );
  NAND U57088 ( .A(n47681), .B(n47682), .Z(n47677) );
  AND U57089 ( .A(n47683), .B(n47684), .Z(n47575) );
  NAND U57090 ( .A(n47685), .B(n47686), .Z(n47684) );
  NAND U57091 ( .A(n47687), .B(n47688), .Z(n47683) );
  AND U57092 ( .A(n47689), .B(n47690), .Z(n47577) );
  XOR U57093 ( .A(n47657), .B(n47656), .Z(N61151) );
  XNOR U57094 ( .A(n47674), .B(n47675), .Z(n47656) );
  XNOR U57095 ( .A(n47689), .B(n47690), .Z(n47675) );
  XOR U57096 ( .A(n47686), .B(n47685), .Z(n47690) );
  XOR U57097 ( .A(y[1044]), .B(x[1044]), .Z(n47685) );
  XOR U57098 ( .A(n47688), .B(n47687), .Z(n47686) );
  XOR U57099 ( .A(y[1046]), .B(x[1046]), .Z(n47687) );
  XOR U57100 ( .A(y[1045]), .B(x[1045]), .Z(n47688) );
  XOR U57101 ( .A(n47680), .B(n47679), .Z(n47689) );
  XOR U57102 ( .A(n47682), .B(n47681), .Z(n47679) );
  XOR U57103 ( .A(y[1043]), .B(x[1043]), .Z(n47681) );
  XOR U57104 ( .A(y[1042]), .B(x[1042]), .Z(n47682) );
  XOR U57105 ( .A(y[1041]), .B(x[1041]), .Z(n47680) );
  XNOR U57106 ( .A(n47673), .B(n47672), .Z(n47674) );
  XNOR U57107 ( .A(n47669), .B(n47668), .Z(n47672) );
  XOR U57108 ( .A(n47671), .B(n47670), .Z(n47668) );
  XOR U57109 ( .A(y[1040]), .B(x[1040]), .Z(n47670) );
  XOR U57110 ( .A(y[1039]), .B(x[1039]), .Z(n47671) );
  XOR U57111 ( .A(y[1038]), .B(x[1038]), .Z(n47669) );
  XOR U57112 ( .A(n47663), .B(n47662), .Z(n47673) );
  XOR U57113 ( .A(n47665), .B(n47664), .Z(n47662) );
  XOR U57114 ( .A(y[1037]), .B(x[1037]), .Z(n47664) );
  XOR U57115 ( .A(y[1036]), .B(x[1036]), .Z(n47665) );
  XOR U57116 ( .A(y[1035]), .B(x[1035]), .Z(n47663) );
  XNOR U57117 ( .A(n47639), .B(n47640), .Z(n47657) );
  XNOR U57118 ( .A(n47654), .B(n47655), .Z(n47640) );
  XOR U57119 ( .A(n47651), .B(n47650), .Z(n47655) );
  XOR U57120 ( .A(y[1032]), .B(x[1032]), .Z(n47650) );
  XOR U57121 ( .A(n47653), .B(n47652), .Z(n47651) );
  XOR U57122 ( .A(y[1034]), .B(x[1034]), .Z(n47652) );
  XOR U57123 ( .A(y[1033]), .B(x[1033]), .Z(n47653) );
  XOR U57124 ( .A(n47645), .B(n47644), .Z(n47654) );
  XOR U57125 ( .A(n47647), .B(n47646), .Z(n47644) );
  XOR U57126 ( .A(y[1031]), .B(x[1031]), .Z(n47646) );
  XOR U57127 ( .A(y[1030]), .B(x[1030]), .Z(n47647) );
  XOR U57128 ( .A(y[1029]), .B(x[1029]), .Z(n47645) );
  XNOR U57129 ( .A(n47638), .B(n47637), .Z(n47639) );
  XNOR U57130 ( .A(n47634), .B(n47633), .Z(n47637) );
  XOR U57131 ( .A(n47636), .B(n47635), .Z(n47633) );
  XOR U57132 ( .A(y[1028]), .B(x[1028]), .Z(n47635) );
  XOR U57133 ( .A(y[1027]), .B(x[1027]), .Z(n47636) );
  XOR U57134 ( .A(y[1026]), .B(x[1026]), .Z(n47634) );
  XOR U57135 ( .A(n47628), .B(n47627), .Z(n47638) );
  XOR U57136 ( .A(n47630), .B(n47629), .Z(n47627) );
  XOR U57137 ( .A(y[1025]), .B(x[1025]), .Z(n47629) );
  XOR U57138 ( .A(y[1024]), .B(x[1024]), .Z(n47630) );
  XOR U57139 ( .A(y[1023]), .B(x[1023]), .Z(n47628) );
  NAND U57140 ( .A(n47691), .B(n47692), .Z(N61142) );
  NAND U57141 ( .A(n47693), .B(n47694), .Z(n47692) );
  NANDN U57142 ( .A(n47695), .B(n47696), .Z(n47694) );
  NANDN U57143 ( .A(n47696), .B(n47695), .Z(n47691) );
  XOR U57144 ( .A(n47695), .B(n47697), .Z(N61141) );
  XNOR U57145 ( .A(n47693), .B(n47696), .Z(n47697) );
  NAND U57146 ( .A(n47698), .B(n47699), .Z(n47696) );
  NAND U57147 ( .A(n47700), .B(n47701), .Z(n47699) );
  NANDN U57148 ( .A(n47702), .B(n47703), .Z(n47701) );
  NANDN U57149 ( .A(n47703), .B(n47702), .Z(n47698) );
  AND U57150 ( .A(n47704), .B(n47705), .Z(n47693) );
  NAND U57151 ( .A(n47706), .B(n47707), .Z(n47705) );
  NANDN U57152 ( .A(n47708), .B(n47709), .Z(n47707) );
  NANDN U57153 ( .A(n47709), .B(n47708), .Z(n47704) );
  IV U57154 ( .A(n47710), .Z(n47709) );
  AND U57155 ( .A(n47711), .B(n47712), .Z(n47695) );
  NAND U57156 ( .A(n47713), .B(n47714), .Z(n47712) );
  NANDN U57157 ( .A(n47715), .B(n47716), .Z(n47714) );
  NANDN U57158 ( .A(n47716), .B(n47715), .Z(n47711) );
  XOR U57159 ( .A(n47708), .B(n47717), .Z(N61140) );
  XNOR U57160 ( .A(n47706), .B(n47710), .Z(n47717) );
  XOR U57161 ( .A(n47703), .B(n47718), .Z(n47710) );
  XNOR U57162 ( .A(n47700), .B(n47702), .Z(n47718) );
  AND U57163 ( .A(n47719), .B(n47720), .Z(n47702) );
  NANDN U57164 ( .A(n47721), .B(n47722), .Z(n47720) );
  OR U57165 ( .A(n47723), .B(n47724), .Z(n47722) );
  IV U57166 ( .A(n47725), .Z(n47724) );
  NANDN U57167 ( .A(n47725), .B(n47723), .Z(n47719) );
  AND U57168 ( .A(n47726), .B(n47727), .Z(n47700) );
  NAND U57169 ( .A(n47728), .B(n47729), .Z(n47727) );
  NANDN U57170 ( .A(n47730), .B(n47731), .Z(n47729) );
  NANDN U57171 ( .A(n47731), .B(n47730), .Z(n47726) );
  IV U57172 ( .A(n47732), .Z(n47731) );
  NAND U57173 ( .A(n47733), .B(n47734), .Z(n47703) );
  NANDN U57174 ( .A(n47735), .B(n47736), .Z(n47734) );
  NANDN U57175 ( .A(n47737), .B(n47738), .Z(n47736) );
  NANDN U57176 ( .A(n47738), .B(n47737), .Z(n47733) );
  IV U57177 ( .A(n47739), .Z(n47737) );
  AND U57178 ( .A(n47740), .B(n47741), .Z(n47706) );
  NAND U57179 ( .A(n47742), .B(n47743), .Z(n47741) );
  NANDN U57180 ( .A(n47744), .B(n47745), .Z(n47743) );
  NANDN U57181 ( .A(n47745), .B(n47744), .Z(n47740) );
  XOR U57182 ( .A(n47716), .B(n47746), .Z(n47708) );
  XNOR U57183 ( .A(n47713), .B(n47715), .Z(n47746) );
  AND U57184 ( .A(n47747), .B(n47748), .Z(n47715) );
  NANDN U57185 ( .A(n47749), .B(n47750), .Z(n47748) );
  OR U57186 ( .A(n47751), .B(n47752), .Z(n47750) );
  IV U57187 ( .A(n47753), .Z(n47752) );
  NANDN U57188 ( .A(n47753), .B(n47751), .Z(n47747) );
  AND U57189 ( .A(n47754), .B(n47755), .Z(n47713) );
  NAND U57190 ( .A(n47756), .B(n47757), .Z(n47755) );
  NANDN U57191 ( .A(n47758), .B(n47759), .Z(n47757) );
  NANDN U57192 ( .A(n47759), .B(n47758), .Z(n47754) );
  IV U57193 ( .A(n47760), .Z(n47759) );
  NAND U57194 ( .A(n47761), .B(n47762), .Z(n47716) );
  NANDN U57195 ( .A(n47763), .B(n47764), .Z(n47762) );
  NANDN U57196 ( .A(n47765), .B(n47766), .Z(n47764) );
  NANDN U57197 ( .A(n47766), .B(n47765), .Z(n47761) );
  IV U57198 ( .A(n47767), .Z(n47765) );
  XOR U57199 ( .A(n47742), .B(n47768), .Z(N61139) );
  XNOR U57200 ( .A(n47745), .B(n47744), .Z(n47768) );
  XNOR U57201 ( .A(n47756), .B(n47769), .Z(n47744) );
  XNOR U57202 ( .A(n47760), .B(n47758), .Z(n47769) );
  XOR U57203 ( .A(n47766), .B(n47770), .Z(n47758) );
  XNOR U57204 ( .A(n47763), .B(n47767), .Z(n47770) );
  AND U57205 ( .A(n47771), .B(n47772), .Z(n47767) );
  NAND U57206 ( .A(n47773), .B(n47774), .Z(n47772) );
  NAND U57207 ( .A(n47775), .B(n47776), .Z(n47771) );
  AND U57208 ( .A(n47777), .B(n47778), .Z(n47763) );
  NAND U57209 ( .A(n47779), .B(n47780), .Z(n47778) );
  NAND U57210 ( .A(n47781), .B(n47782), .Z(n47777) );
  NANDN U57211 ( .A(n47783), .B(n47784), .Z(n47766) );
  ANDN U57212 ( .B(n47785), .A(n47786), .Z(n47760) );
  XNOR U57213 ( .A(n47751), .B(n47787), .Z(n47756) );
  XNOR U57214 ( .A(n47749), .B(n47753), .Z(n47787) );
  AND U57215 ( .A(n47788), .B(n47789), .Z(n47753) );
  NAND U57216 ( .A(n47790), .B(n47791), .Z(n47789) );
  NAND U57217 ( .A(n47792), .B(n47793), .Z(n47788) );
  AND U57218 ( .A(n47794), .B(n47795), .Z(n47749) );
  NAND U57219 ( .A(n47796), .B(n47797), .Z(n47795) );
  NAND U57220 ( .A(n47798), .B(n47799), .Z(n47794) );
  AND U57221 ( .A(n47800), .B(n47801), .Z(n47751) );
  NAND U57222 ( .A(n47802), .B(n47803), .Z(n47745) );
  XNOR U57223 ( .A(n47728), .B(n47804), .Z(n47742) );
  XNOR U57224 ( .A(n47732), .B(n47730), .Z(n47804) );
  XOR U57225 ( .A(n47738), .B(n47805), .Z(n47730) );
  XNOR U57226 ( .A(n47735), .B(n47739), .Z(n47805) );
  AND U57227 ( .A(n47806), .B(n47807), .Z(n47739) );
  NAND U57228 ( .A(n47808), .B(n47809), .Z(n47807) );
  NAND U57229 ( .A(n47810), .B(n47811), .Z(n47806) );
  AND U57230 ( .A(n47812), .B(n47813), .Z(n47735) );
  NAND U57231 ( .A(n47814), .B(n47815), .Z(n47813) );
  NAND U57232 ( .A(n47816), .B(n47817), .Z(n47812) );
  NANDN U57233 ( .A(n47818), .B(n47819), .Z(n47738) );
  ANDN U57234 ( .B(n47820), .A(n47821), .Z(n47732) );
  XNOR U57235 ( .A(n47723), .B(n47822), .Z(n47728) );
  XNOR U57236 ( .A(n47721), .B(n47725), .Z(n47822) );
  AND U57237 ( .A(n47823), .B(n47824), .Z(n47725) );
  NAND U57238 ( .A(n47825), .B(n47826), .Z(n47824) );
  NAND U57239 ( .A(n47827), .B(n47828), .Z(n47823) );
  AND U57240 ( .A(n47829), .B(n47830), .Z(n47721) );
  NAND U57241 ( .A(n47831), .B(n47832), .Z(n47830) );
  NAND U57242 ( .A(n47833), .B(n47834), .Z(n47829) );
  AND U57243 ( .A(n47835), .B(n47836), .Z(n47723) );
  XOR U57244 ( .A(n47803), .B(n47802), .Z(N61138) );
  XNOR U57245 ( .A(n47820), .B(n47821), .Z(n47802) );
  XNOR U57246 ( .A(n47835), .B(n47836), .Z(n47821) );
  XOR U57247 ( .A(n47832), .B(n47831), .Z(n47836) );
  XOR U57248 ( .A(y[1020]), .B(x[1020]), .Z(n47831) );
  XOR U57249 ( .A(n47834), .B(n47833), .Z(n47832) );
  XOR U57250 ( .A(y[1022]), .B(x[1022]), .Z(n47833) );
  XOR U57251 ( .A(y[1021]), .B(x[1021]), .Z(n47834) );
  XOR U57252 ( .A(n47826), .B(n47825), .Z(n47835) );
  XOR U57253 ( .A(n47828), .B(n47827), .Z(n47825) );
  XOR U57254 ( .A(y[1019]), .B(x[1019]), .Z(n47827) );
  XOR U57255 ( .A(y[1018]), .B(x[1018]), .Z(n47828) );
  XOR U57256 ( .A(y[1017]), .B(x[1017]), .Z(n47826) );
  XNOR U57257 ( .A(n47819), .B(n47818), .Z(n47820) );
  XNOR U57258 ( .A(n47815), .B(n47814), .Z(n47818) );
  XOR U57259 ( .A(n47817), .B(n47816), .Z(n47814) );
  XOR U57260 ( .A(y[1016]), .B(x[1016]), .Z(n47816) );
  XOR U57261 ( .A(y[1015]), .B(x[1015]), .Z(n47817) );
  XOR U57262 ( .A(y[1014]), .B(x[1014]), .Z(n47815) );
  XOR U57263 ( .A(n47809), .B(n47808), .Z(n47819) );
  XOR U57264 ( .A(n47811), .B(n47810), .Z(n47808) );
  XOR U57265 ( .A(y[1013]), .B(x[1013]), .Z(n47810) );
  XOR U57266 ( .A(y[1012]), .B(x[1012]), .Z(n47811) );
  XOR U57267 ( .A(y[1011]), .B(x[1011]), .Z(n47809) );
  XNOR U57268 ( .A(n47785), .B(n47786), .Z(n47803) );
  XNOR U57269 ( .A(n47800), .B(n47801), .Z(n47786) );
  XOR U57270 ( .A(n47797), .B(n47796), .Z(n47801) );
  XOR U57271 ( .A(y[1008]), .B(x[1008]), .Z(n47796) );
  XOR U57272 ( .A(n47799), .B(n47798), .Z(n47797) );
  XOR U57273 ( .A(y[1010]), .B(x[1010]), .Z(n47798) );
  XOR U57274 ( .A(y[1009]), .B(x[1009]), .Z(n47799) );
  XOR U57275 ( .A(n47791), .B(n47790), .Z(n47800) );
  XOR U57276 ( .A(n47793), .B(n47792), .Z(n47790) );
  XOR U57277 ( .A(y[1007]), .B(x[1007]), .Z(n47792) );
  XOR U57278 ( .A(y[1006]), .B(x[1006]), .Z(n47793) );
  XOR U57279 ( .A(y[1005]), .B(x[1005]), .Z(n47791) );
  XNOR U57280 ( .A(n47784), .B(n47783), .Z(n47785) );
  XNOR U57281 ( .A(n47780), .B(n47779), .Z(n47783) );
  XOR U57282 ( .A(n47782), .B(n47781), .Z(n47779) );
  XOR U57283 ( .A(y[1004]), .B(x[1004]), .Z(n47781) );
  XOR U57284 ( .A(y[1003]), .B(x[1003]), .Z(n47782) );
  XOR U57285 ( .A(y[1002]), .B(x[1002]), .Z(n47780) );
  XOR U57286 ( .A(n47774), .B(n47773), .Z(n47784) );
  XOR U57287 ( .A(n47776), .B(n47775), .Z(n47773) );
  XOR U57288 ( .A(y[1001]), .B(x[1001]), .Z(n47775) );
  XOR U57289 ( .A(y[1000]), .B(x[1000]), .Z(n47776) );
  XOR U57290 ( .A(y[999]), .B(x[999]), .Z(n47774) );
  NAND U57291 ( .A(n47837), .B(n47838), .Z(N61129) );
  NAND U57292 ( .A(n47839), .B(n47840), .Z(n47838) );
  NANDN U57293 ( .A(n47841), .B(n47842), .Z(n47840) );
  NANDN U57294 ( .A(n47842), .B(n47841), .Z(n47837) );
  XOR U57295 ( .A(n47841), .B(n47843), .Z(N61128) );
  XNOR U57296 ( .A(n47839), .B(n47842), .Z(n47843) );
  NAND U57297 ( .A(n47844), .B(n47845), .Z(n47842) );
  NAND U57298 ( .A(n47846), .B(n47847), .Z(n47845) );
  NANDN U57299 ( .A(n47848), .B(n47849), .Z(n47847) );
  NANDN U57300 ( .A(n47849), .B(n47848), .Z(n47844) );
  AND U57301 ( .A(n47850), .B(n47851), .Z(n47839) );
  NAND U57302 ( .A(n47852), .B(n47853), .Z(n47851) );
  NANDN U57303 ( .A(n47854), .B(n47855), .Z(n47853) );
  NANDN U57304 ( .A(n47855), .B(n47854), .Z(n47850) );
  IV U57305 ( .A(n47856), .Z(n47855) );
  AND U57306 ( .A(n47857), .B(n47858), .Z(n47841) );
  NAND U57307 ( .A(n47859), .B(n47860), .Z(n47858) );
  NANDN U57308 ( .A(n47861), .B(n47862), .Z(n47860) );
  NANDN U57309 ( .A(n47862), .B(n47861), .Z(n47857) );
  XOR U57310 ( .A(n47854), .B(n47863), .Z(N61127) );
  XNOR U57311 ( .A(n47852), .B(n47856), .Z(n47863) );
  XOR U57312 ( .A(n47849), .B(n47864), .Z(n47856) );
  XNOR U57313 ( .A(n47846), .B(n47848), .Z(n47864) );
  AND U57314 ( .A(n47865), .B(n47866), .Z(n47848) );
  NANDN U57315 ( .A(n47867), .B(n47868), .Z(n47866) );
  OR U57316 ( .A(n47869), .B(n47870), .Z(n47868) );
  IV U57317 ( .A(n47871), .Z(n47870) );
  NANDN U57318 ( .A(n47871), .B(n47869), .Z(n47865) );
  AND U57319 ( .A(n47872), .B(n47873), .Z(n47846) );
  NAND U57320 ( .A(n47874), .B(n47875), .Z(n47873) );
  NANDN U57321 ( .A(n47876), .B(n47877), .Z(n47875) );
  NANDN U57322 ( .A(n47877), .B(n47876), .Z(n47872) );
  IV U57323 ( .A(n47878), .Z(n47877) );
  NAND U57324 ( .A(n47879), .B(n47880), .Z(n47849) );
  NANDN U57325 ( .A(n47881), .B(n47882), .Z(n47880) );
  NANDN U57326 ( .A(n47883), .B(n47884), .Z(n47882) );
  NANDN U57327 ( .A(n47884), .B(n47883), .Z(n47879) );
  IV U57328 ( .A(n47885), .Z(n47883) );
  AND U57329 ( .A(n47886), .B(n47887), .Z(n47852) );
  NAND U57330 ( .A(n47888), .B(n47889), .Z(n47887) );
  NANDN U57331 ( .A(n47890), .B(n47891), .Z(n47889) );
  NANDN U57332 ( .A(n47891), .B(n47890), .Z(n47886) );
  XOR U57333 ( .A(n47862), .B(n47892), .Z(n47854) );
  XNOR U57334 ( .A(n47859), .B(n47861), .Z(n47892) );
  AND U57335 ( .A(n47893), .B(n47894), .Z(n47861) );
  NANDN U57336 ( .A(n47895), .B(n47896), .Z(n47894) );
  OR U57337 ( .A(n47897), .B(n47898), .Z(n47896) );
  IV U57338 ( .A(n47899), .Z(n47898) );
  NANDN U57339 ( .A(n47899), .B(n47897), .Z(n47893) );
  AND U57340 ( .A(n47900), .B(n47901), .Z(n47859) );
  NAND U57341 ( .A(n47902), .B(n47903), .Z(n47901) );
  NANDN U57342 ( .A(n47904), .B(n47905), .Z(n47903) );
  NANDN U57343 ( .A(n47905), .B(n47904), .Z(n47900) );
  IV U57344 ( .A(n47906), .Z(n47905) );
  NAND U57345 ( .A(n47907), .B(n47908), .Z(n47862) );
  NANDN U57346 ( .A(n47909), .B(n47910), .Z(n47908) );
  NANDN U57347 ( .A(n47911), .B(n47912), .Z(n47910) );
  NANDN U57348 ( .A(n47912), .B(n47911), .Z(n47907) );
  IV U57349 ( .A(n47913), .Z(n47911) );
  XOR U57350 ( .A(n47888), .B(n47914), .Z(N61126) );
  XNOR U57351 ( .A(n47891), .B(n47890), .Z(n47914) );
  XNOR U57352 ( .A(n47902), .B(n47915), .Z(n47890) );
  XNOR U57353 ( .A(n47906), .B(n47904), .Z(n47915) );
  XOR U57354 ( .A(n47912), .B(n47916), .Z(n47904) );
  XNOR U57355 ( .A(n47909), .B(n47913), .Z(n47916) );
  AND U57356 ( .A(n47917), .B(n47918), .Z(n47913) );
  NAND U57357 ( .A(n47919), .B(n47920), .Z(n47918) );
  NAND U57358 ( .A(n47921), .B(n47922), .Z(n47917) );
  AND U57359 ( .A(n47923), .B(n47924), .Z(n47909) );
  NAND U57360 ( .A(n47925), .B(n47926), .Z(n47924) );
  NAND U57361 ( .A(n47927), .B(n47928), .Z(n47923) );
  NANDN U57362 ( .A(n47929), .B(n47930), .Z(n47912) );
  ANDN U57363 ( .B(n47931), .A(n47932), .Z(n47906) );
  XNOR U57364 ( .A(n47897), .B(n47933), .Z(n47902) );
  XNOR U57365 ( .A(n47895), .B(n47899), .Z(n47933) );
  AND U57366 ( .A(n47934), .B(n47935), .Z(n47899) );
  NAND U57367 ( .A(n47936), .B(n47937), .Z(n47935) );
  NAND U57368 ( .A(n47938), .B(n47939), .Z(n47934) );
  AND U57369 ( .A(n47940), .B(n47941), .Z(n47895) );
  NAND U57370 ( .A(n47942), .B(n47943), .Z(n47941) );
  NAND U57371 ( .A(n47944), .B(n47945), .Z(n47940) );
  AND U57372 ( .A(n47946), .B(n47947), .Z(n47897) );
  NAND U57373 ( .A(n47948), .B(n47949), .Z(n47891) );
  XNOR U57374 ( .A(n47874), .B(n47950), .Z(n47888) );
  XNOR U57375 ( .A(n47878), .B(n47876), .Z(n47950) );
  XOR U57376 ( .A(n47884), .B(n47951), .Z(n47876) );
  XNOR U57377 ( .A(n47881), .B(n47885), .Z(n47951) );
  AND U57378 ( .A(n47952), .B(n47953), .Z(n47885) );
  NAND U57379 ( .A(n47954), .B(n47955), .Z(n47953) );
  NAND U57380 ( .A(n47956), .B(n47957), .Z(n47952) );
  AND U57381 ( .A(n47958), .B(n47959), .Z(n47881) );
  NAND U57382 ( .A(n47960), .B(n47961), .Z(n47959) );
  NAND U57383 ( .A(n47962), .B(n47963), .Z(n47958) );
  NANDN U57384 ( .A(n47964), .B(n47965), .Z(n47884) );
  ANDN U57385 ( .B(n47966), .A(n47967), .Z(n47878) );
  XNOR U57386 ( .A(n47869), .B(n47968), .Z(n47874) );
  XNOR U57387 ( .A(n47867), .B(n47871), .Z(n47968) );
  AND U57388 ( .A(n47969), .B(n47970), .Z(n47871) );
  NAND U57389 ( .A(n47971), .B(n47972), .Z(n47970) );
  NAND U57390 ( .A(n47973), .B(n47974), .Z(n47969) );
  AND U57391 ( .A(n47975), .B(n47976), .Z(n47867) );
  NAND U57392 ( .A(n47977), .B(n47978), .Z(n47976) );
  NAND U57393 ( .A(n47979), .B(n47980), .Z(n47975) );
  AND U57394 ( .A(n47981), .B(n47982), .Z(n47869) );
  XOR U57395 ( .A(n47949), .B(n47948), .Z(N61125) );
  XNOR U57396 ( .A(n47966), .B(n47967), .Z(n47948) );
  XNOR U57397 ( .A(n47981), .B(n47982), .Z(n47967) );
  XOR U57398 ( .A(n47978), .B(n47977), .Z(n47982) );
  XOR U57399 ( .A(y[996]), .B(x[996]), .Z(n47977) );
  XOR U57400 ( .A(n47980), .B(n47979), .Z(n47978) );
  XOR U57401 ( .A(y[998]), .B(x[998]), .Z(n47979) );
  XOR U57402 ( .A(y[997]), .B(x[997]), .Z(n47980) );
  XOR U57403 ( .A(n47972), .B(n47971), .Z(n47981) );
  XOR U57404 ( .A(n47974), .B(n47973), .Z(n47971) );
  XOR U57405 ( .A(y[995]), .B(x[995]), .Z(n47973) );
  XOR U57406 ( .A(y[994]), .B(x[994]), .Z(n47974) );
  XOR U57407 ( .A(y[993]), .B(x[993]), .Z(n47972) );
  XNOR U57408 ( .A(n47965), .B(n47964), .Z(n47966) );
  XNOR U57409 ( .A(n47961), .B(n47960), .Z(n47964) );
  XOR U57410 ( .A(n47963), .B(n47962), .Z(n47960) );
  XOR U57411 ( .A(y[992]), .B(x[992]), .Z(n47962) );
  XOR U57412 ( .A(y[991]), .B(x[991]), .Z(n47963) );
  XOR U57413 ( .A(y[990]), .B(x[990]), .Z(n47961) );
  XOR U57414 ( .A(n47955), .B(n47954), .Z(n47965) );
  XOR U57415 ( .A(n47957), .B(n47956), .Z(n47954) );
  XOR U57416 ( .A(y[989]), .B(x[989]), .Z(n47956) );
  XOR U57417 ( .A(y[988]), .B(x[988]), .Z(n47957) );
  XOR U57418 ( .A(y[987]), .B(x[987]), .Z(n47955) );
  XNOR U57419 ( .A(n47931), .B(n47932), .Z(n47949) );
  XNOR U57420 ( .A(n47946), .B(n47947), .Z(n47932) );
  XOR U57421 ( .A(n47943), .B(n47942), .Z(n47947) );
  XOR U57422 ( .A(y[984]), .B(x[984]), .Z(n47942) );
  XOR U57423 ( .A(n47945), .B(n47944), .Z(n47943) );
  XOR U57424 ( .A(y[986]), .B(x[986]), .Z(n47944) );
  XOR U57425 ( .A(y[985]), .B(x[985]), .Z(n47945) );
  XOR U57426 ( .A(n47937), .B(n47936), .Z(n47946) );
  XOR U57427 ( .A(n47939), .B(n47938), .Z(n47936) );
  XOR U57428 ( .A(y[983]), .B(x[983]), .Z(n47938) );
  XOR U57429 ( .A(y[982]), .B(x[982]), .Z(n47939) );
  XOR U57430 ( .A(y[981]), .B(x[981]), .Z(n47937) );
  XNOR U57431 ( .A(n47930), .B(n47929), .Z(n47931) );
  XNOR U57432 ( .A(n47926), .B(n47925), .Z(n47929) );
  XOR U57433 ( .A(n47928), .B(n47927), .Z(n47925) );
  XOR U57434 ( .A(y[980]), .B(x[980]), .Z(n47927) );
  XOR U57435 ( .A(y[979]), .B(x[979]), .Z(n47928) );
  XOR U57436 ( .A(y[978]), .B(x[978]), .Z(n47926) );
  XOR U57437 ( .A(n47920), .B(n47919), .Z(n47930) );
  XOR U57438 ( .A(n47922), .B(n47921), .Z(n47919) );
  XOR U57439 ( .A(y[977]), .B(x[977]), .Z(n47921) );
  XOR U57440 ( .A(y[976]), .B(x[976]), .Z(n47922) );
  XOR U57441 ( .A(y[975]), .B(x[975]), .Z(n47920) );
  NAND U57442 ( .A(n47983), .B(n47984), .Z(N61116) );
  NAND U57443 ( .A(n47985), .B(n47986), .Z(n47984) );
  NANDN U57444 ( .A(n47987), .B(n47988), .Z(n47986) );
  NANDN U57445 ( .A(n47988), .B(n47987), .Z(n47983) );
  XOR U57446 ( .A(n47987), .B(n47989), .Z(N61115) );
  XNOR U57447 ( .A(n47985), .B(n47988), .Z(n47989) );
  NAND U57448 ( .A(n47990), .B(n47991), .Z(n47988) );
  NAND U57449 ( .A(n47992), .B(n47993), .Z(n47991) );
  NANDN U57450 ( .A(n47994), .B(n47995), .Z(n47993) );
  NANDN U57451 ( .A(n47995), .B(n47994), .Z(n47990) );
  AND U57452 ( .A(n47996), .B(n47997), .Z(n47985) );
  NAND U57453 ( .A(n47998), .B(n47999), .Z(n47997) );
  NANDN U57454 ( .A(n48000), .B(n48001), .Z(n47999) );
  NANDN U57455 ( .A(n48001), .B(n48000), .Z(n47996) );
  IV U57456 ( .A(n48002), .Z(n48001) );
  AND U57457 ( .A(n48003), .B(n48004), .Z(n47987) );
  NAND U57458 ( .A(n48005), .B(n48006), .Z(n48004) );
  NANDN U57459 ( .A(n48007), .B(n48008), .Z(n48006) );
  NANDN U57460 ( .A(n48008), .B(n48007), .Z(n48003) );
  XOR U57461 ( .A(n48000), .B(n48009), .Z(N61114) );
  XNOR U57462 ( .A(n47998), .B(n48002), .Z(n48009) );
  XOR U57463 ( .A(n47995), .B(n48010), .Z(n48002) );
  XNOR U57464 ( .A(n47992), .B(n47994), .Z(n48010) );
  AND U57465 ( .A(n48011), .B(n48012), .Z(n47994) );
  NANDN U57466 ( .A(n48013), .B(n48014), .Z(n48012) );
  OR U57467 ( .A(n48015), .B(n48016), .Z(n48014) );
  IV U57468 ( .A(n48017), .Z(n48016) );
  NANDN U57469 ( .A(n48017), .B(n48015), .Z(n48011) );
  AND U57470 ( .A(n48018), .B(n48019), .Z(n47992) );
  NAND U57471 ( .A(n48020), .B(n48021), .Z(n48019) );
  NANDN U57472 ( .A(n48022), .B(n48023), .Z(n48021) );
  NANDN U57473 ( .A(n48023), .B(n48022), .Z(n48018) );
  IV U57474 ( .A(n48024), .Z(n48023) );
  NAND U57475 ( .A(n48025), .B(n48026), .Z(n47995) );
  NANDN U57476 ( .A(n48027), .B(n48028), .Z(n48026) );
  NANDN U57477 ( .A(n48029), .B(n48030), .Z(n48028) );
  NANDN U57478 ( .A(n48030), .B(n48029), .Z(n48025) );
  IV U57479 ( .A(n48031), .Z(n48029) );
  AND U57480 ( .A(n48032), .B(n48033), .Z(n47998) );
  NAND U57481 ( .A(n48034), .B(n48035), .Z(n48033) );
  NANDN U57482 ( .A(n48036), .B(n48037), .Z(n48035) );
  NANDN U57483 ( .A(n48037), .B(n48036), .Z(n48032) );
  XOR U57484 ( .A(n48008), .B(n48038), .Z(n48000) );
  XNOR U57485 ( .A(n48005), .B(n48007), .Z(n48038) );
  AND U57486 ( .A(n48039), .B(n48040), .Z(n48007) );
  NANDN U57487 ( .A(n48041), .B(n48042), .Z(n48040) );
  OR U57488 ( .A(n48043), .B(n48044), .Z(n48042) );
  IV U57489 ( .A(n48045), .Z(n48044) );
  NANDN U57490 ( .A(n48045), .B(n48043), .Z(n48039) );
  AND U57491 ( .A(n48046), .B(n48047), .Z(n48005) );
  NAND U57492 ( .A(n48048), .B(n48049), .Z(n48047) );
  NANDN U57493 ( .A(n48050), .B(n48051), .Z(n48049) );
  NANDN U57494 ( .A(n48051), .B(n48050), .Z(n48046) );
  IV U57495 ( .A(n48052), .Z(n48051) );
  NAND U57496 ( .A(n48053), .B(n48054), .Z(n48008) );
  NANDN U57497 ( .A(n48055), .B(n48056), .Z(n48054) );
  NANDN U57498 ( .A(n48057), .B(n48058), .Z(n48056) );
  NANDN U57499 ( .A(n48058), .B(n48057), .Z(n48053) );
  IV U57500 ( .A(n48059), .Z(n48057) );
  XOR U57501 ( .A(n48034), .B(n48060), .Z(N61113) );
  XNOR U57502 ( .A(n48037), .B(n48036), .Z(n48060) );
  XNOR U57503 ( .A(n48048), .B(n48061), .Z(n48036) );
  XNOR U57504 ( .A(n48052), .B(n48050), .Z(n48061) );
  XOR U57505 ( .A(n48058), .B(n48062), .Z(n48050) );
  XNOR U57506 ( .A(n48055), .B(n48059), .Z(n48062) );
  AND U57507 ( .A(n48063), .B(n48064), .Z(n48059) );
  NAND U57508 ( .A(n48065), .B(n48066), .Z(n48064) );
  NAND U57509 ( .A(n48067), .B(n48068), .Z(n48063) );
  AND U57510 ( .A(n48069), .B(n48070), .Z(n48055) );
  NAND U57511 ( .A(n48071), .B(n48072), .Z(n48070) );
  NAND U57512 ( .A(n48073), .B(n48074), .Z(n48069) );
  NANDN U57513 ( .A(n48075), .B(n48076), .Z(n48058) );
  ANDN U57514 ( .B(n48077), .A(n48078), .Z(n48052) );
  XNOR U57515 ( .A(n48043), .B(n48079), .Z(n48048) );
  XNOR U57516 ( .A(n48041), .B(n48045), .Z(n48079) );
  AND U57517 ( .A(n48080), .B(n48081), .Z(n48045) );
  NAND U57518 ( .A(n48082), .B(n48083), .Z(n48081) );
  NAND U57519 ( .A(n48084), .B(n48085), .Z(n48080) );
  AND U57520 ( .A(n48086), .B(n48087), .Z(n48041) );
  NAND U57521 ( .A(n48088), .B(n48089), .Z(n48087) );
  NAND U57522 ( .A(n48090), .B(n48091), .Z(n48086) );
  AND U57523 ( .A(n48092), .B(n48093), .Z(n48043) );
  NAND U57524 ( .A(n48094), .B(n48095), .Z(n48037) );
  XNOR U57525 ( .A(n48020), .B(n48096), .Z(n48034) );
  XNOR U57526 ( .A(n48024), .B(n48022), .Z(n48096) );
  XOR U57527 ( .A(n48030), .B(n48097), .Z(n48022) );
  XNOR U57528 ( .A(n48027), .B(n48031), .Z(n48097) );
  AND U57529 ( .A(n48098), .B(n48099), .Z(n48031) );
  NAND U57530 ( .A(n48100), .B(n48101), .Z(n48099) );
  NAND U57531 ( .A(n48102), .B(n48103), .Z(n48098) );
  AND U57532 ( .A(n48104), .B(n48105), .Z(n48027) );
  NAND U57533 ( .A(n48106), .B(n48107), .Z(n48105) );
  NAND U57534 ( .A(n48108), .B(n48109), .Z(n48104) );
  NANDN U57535 ( .A(n48110), .B(n48111), .Z(n48030) );
  ANDN U57536 ( .B(n48112), .A(n48113), .Z(n48024) );
  XNOR U57537 ( .A(n48015), .B(n48114), .Z(n48020) );
  XNOR U57538 ( .A(n48013), .B(n48017), .Z(n48114) );
  AND U57539 ( .A(n48115), .B(n48116), .Z(n48017) );
  NAND U57540 ( .A(n48117), .B(n48118), .Z(n48116) );
  NAND U57541 ( .A(n48119), .B(n48120), .Z(n48115) );
  AND U57542 ( .A(n48121), .B(n48122), .Z(n48013) );
  NAND U57543 ( .A(n48123), .B(n48124), .Z(n48122) );
  NAND U57544 ( .A(n48125), .B(n48126), .Z(n48121) );
  AND U57545 ( .A(n48127), .B(n48128), .Z(n48015) );
  XOR U57546 ( .A(n48095), .B(n48094), .Z(N61112) );
  XNOR U57547 ( .A(n48112), .B(n48113), .Z(n48094) );
  XNOR U57548 ( .A(n48127), .B(n48128), .Z(n48113) );
  XOR U57549 ( .A(n48124), .B(n48123), .Z(n48128) );
  XOR U57550 ( .A(y[972]), .B(x[972]), .Z(n48123) );
  XOR U57551 ( .A(n48126), .B(n48125), .Z(n48124) );
  XOR U57552 ( .A(y[974]), .B(x[974]), .Z(n48125) );
  XOR U57553 ( .A(y[973]), .B(x[973]), .Z(n48126) );
  XOR U57554 ( .A(n48118), .B(n48117), .Z(n48127) );
  XOR U57555 ( .A(n48120), .B(n48119), .Z(n48117) );
  XOR U57556 ( .A(y[971]), .B(x[971]), .Z(n48119) );
  XOR U57557 ( .A(y[970]), .B(x[970]), .Z(n48120) );
  XOR U57558 ( .A(y[969]), .B(x[969]), .Z(n48118) );
  XNOR U57559 ( .A(n48111), .B(n48110), .Z(n48112) );
  XNOR U57560 ( .A(n48107), .B(n48106), .Z(n48110) );
  XOR U57561 ( .A(n48109), .B(n48108), .Z(n48106) );
  XOR U57562 ( .A(y[968]), .B(x[968]), .Z(n48108) );
  XOR U57563 ( .A(y[967]), .B(x[967]), .Z(n48109) );
  XOR U57564 ( .A(y[966]), .B(x[966]), .Z(n48107) );
  XOR U57565 ( .A(n48101), .B(n48100), .Z(n48111) );
  XOR U57566 ( .A(n48103), .B(n48102), .Z(n48100) );
  XOR U57567 ( .A(y[965]), .B(x[965]), .Z(n48102) );
  XOR U57568 ( .A(y[964]), .B(x[964]), .Z(n48103) );
  XOR U57569 ( .A(y[963]), .B(x[963]), .Z(n48101) );
  XNOR U57570 ( .A(n48077), .B(n48078), .Z(n48095) );
  XNOR U57571 ( .A(n48092), .B(n48093), .Z(n48078) );
  XOR U57572 ( .A(n48089), .B(n48088), .Z(n48093) );
  XOR U57573 ( .A(y[960]), .B(x[960]), .Z(n48088) );
  XOR U57574 ( .A(n48091), .B(n48090), .Z(n48089) );
  XOR U57575 ( .A(y[962]), .B(x[962]), .Z(n48090) );
  XOR U57576 ( .A(y[961]), .B(x[961]), .Z(n48091) );
  XOR U57577 ( .A(n48083), .B(n48082), .Z(n48092) );
  XOR U57578 ( .A(n48085), .B(n48084), .Z(n48082) );
  XOR U57579 ( .A(y[959]), .B(x[959]), .Z(n48084) );
  XOR U57580 ( .A(y[958]), .B(x[958]), .Z(n48085) );
  XOR U57581 ( .A(y[957]), .B(x[957]), .Z(n48083) );
  XNOR U57582 ( .A(n48076), .B(n48075), .Z(n48077) );
  XNOR U57583 ( .A(n48072), .B(n48071), .Z(n48075) );
  XOR U57584 ( .A(n48074), .B(n48073), .Z(n48071) );
  XOR U57585 ( .A(y[956]), .B(x[956]), .Z(n48073) );
  XOR U57586 ( .A(y[955]), .B(x[955]), .Z(n48074) );
  XOR U57587 ( .A(y[954]), .B(x[954]), .Z(n48072) );
  XOR U57588 ( .A(n48066), .B(n48065), .Z(n48076) );
  XOR U57589 ( .A(n48068), .B(n48067), .Z(n48065) );
  XOR U57590 ( .A(y[953]), .B(x[953]), .Z(n48067) );
  XOR U57591 ( .A(y[952]), .B(x[952]), .Z(n48068) );
  XOR U57592 ( .A(y[951]), .B(x[951]), .Z(n48066) );
  NAND U57593 ( .A(n48129), .B(n48130), .Z(N61103) );
  NAND U57594 ( .A(n48131), .B(n48132), .Z(n48130) );
  NANDN U57595 ( .A(n48133), .B(n48134), .Z(n48132) );
  NANDN U57596 ( .A(n48134), .B(n48133), .Z(n48129) );
  XOR U57597 ( .A(n48133), .B(n48135), .Z(N61102) );
  XNOR U57598 ( .A(n48131), .B(n48134), .Z(n48135) );
  NAND U57599 ( .A(n48136), .B(n48137), .Z(n48134) );
  NAND U57600 ( .A(n48138), .B(n48139), .Z(n48137) );
  NANDN U57601 ( .A(n48140), .B(n48141), .Z(n48139) );
  NANDN U57602 ( .A(n48141), .B(n48140), .Z(n48136) );
  AND U57603 ( .A(n48142), .B(n48143), .Z(n48131) );
  NAND U57604 ( .A(n48144), .B(n48145), .Z(n48143) );
  NANDN U57605 ( .A(n48146), .B(n48147), .Z(n48145) );
  NANDN U57606 ( .A(n48147), .B(n48146), .Z(n48142) );
  IV U57607 ( .A(n48148), .Z(n48147) );
  AND U57608 ( .A(n48149), .B(n48150), .Z(n48133) );
  NAND U57609 ( .A(n48151), .B(n48152), .Z(n48150) );
  NANDN U57610 ( .A(n48153), .B(n48154), .Z(n48152) );
  NANDN U57611 ( .A(n48154), .B(n48153), .Z(n48149) );
  XOR U57612 ( .A(n48146), .B(n48155), .Z(N61101) );
  XNOR U57613 ( .A(n48144), .B(n48148), .Z(n48155) );
  XOR U57614 ( .A(n48141), .B(n48156), .Z(n48148) );
  XNOR U57615 ( .A(n48138), .B(n48140), .Z(n48156) );
  AND U57616 ( .A(n48157), .B(n48158), .Z(n48140) );
  NANDN U57617 ( .A(n48159), .B(n48160), .Z(n48158) );
  OR U57618 ( .A(n48161), .B(n48162), .Z(n48160) );
  IV U57619 ( .A(n48163), .Z(n48162) );
  NANDN U57620 ( .A(n48163), .B(n48161), .Z(n48157) );
  AND U57621 ( .A(n48164), .B(n48165), .Z(n48138) );
  NAND U57622 ( .A(n48166), .B(n48167), .Z(n48165) );
  NANDN U57623 ( .A(n48168), .B(n48169), .Z(n48167) );
  NANDN U57624 ( .A(n48169), .B(n48168), .Z(n48164) );
  IV U57625 ( .A(n48170), .Z(n48169) );
  NAND U57626 ( .A(n48171), .B(n48172), .Z(n48141) );
  NANDN U57627 ( .A(n48173), .B(n48174), .Z(n48172) );
  NANDN U57628 ( .A(n48175), .B(n48176), .Z(n48174) );
  NANDN U57629 ( .A(n48176), .B(n48175), .Z(n48171) );
  IV U57630 ( .A(n48177), .Z(n48175) );
  AND U57631 ( .A(n48178), .B(n48179), .Z(n48144) );
  NAND U57632 ( .A(n48180), .B(n48181), .Z(n48179) );
  NANDN U57633 ( .A(n48182), .B(n48183), .Z(n48181) );
  NANDN U57634 ( .A(n48183), .B(n48182), .Z(n48178) );
  XOR U57635 ( .A(n48154), .B(n48184), .Z(n48146) );
  XNOR U57636 ( .A(n48151), .B(n48153), .Z(n48184) );
  AND U57637 ( .A(n48185), .B(n48186), .Z(n48153) );
  NANDN U57638 ( .A(n48187), .B(n48188), .Z(n48186) );
  OR U57639 ( .A(n48189), .B(n48190), .Z(n48188) );
  IV U57640 ( .A(n48191), .Z(n48190) );
  NANDN U57641 ( .A(n48191), .B(n48189), .Z(n48185) );
  AND U57642 ( .A(n48192), .B(n48193), .Z(n48151) );
  NAND U57643 ( .A(n48194), .B(n48195), .Z(n48193) );
  NANDN U57644 ( .A(n48196), .B(n48197), .Z(n48195) );
  NANDN U57645 ( .A(n48197), .B(n48196), .Z(n48192) );
  IV U57646 ( .A(n48198), .Z(n48197) );
  NAND U57647 ( .A(n48199), .B(n48200), .Z(n48154) );
  NANDN U57648 ( .A(n48201), .B(n48202), .Z(n48200) );
  NANDN U57649 ( .A(n48203), .B(n48204), .Z(n48202) );
  NANDN U57650 ( .A(n48204), .B(n48203), .Z(n48199) );
  IV U57651 ( .A(n48205), .Z(n48203) );
  XOR U57652 ( .A(n48180), .B(n48206), .Z(N61100) );
  XNOR U57653 ( .A(n48183), .B(n48182), .Z(n48206) );
  XNOR U57654 ( .A(n48194), .B(n48207), .Z(n48182) );
  XNOR U57655 ( .A(n48198), .B(n48196), .Z(n48207) );
  XOR U57656 ( .A(n48204), .B(n48208), .Z(n48196) );
  XNOR U57657 ( .A(n48201), .B(n48205), .Z(n48208) );
  AND U57658 ( .A(n48209), .B(n48210), .Z(n48205) );
  NAND U57659 ( .A(n48211), .B(n48212), .Z(n48210) );
  NAND U57660 ( .A(n48213), .B(n48214), .Z(n48209) );
  AND U57661 ( .A(n48215), .B(n48216), .Z(n48201) );
  NAND U57662 ( .A(n48217), .B(n48218), .Z(n48216) );
  NAND U57663 ( .A(n48219), .B(n48220), .Z(n48215) );
  NANDN U57664 ( .A(n48221), .B(n48222), .Z(n48204) );
  ANDN U57665 ( .B(n48223), .A(n48224), .Z(n48198) );
  XNOR U57666 ( .A(n48189), .B(n48225), .Z(n48194) );
  XNOR U57667 ( .A(n48187), .B(n48191), .Z(n48225) );
  AND U57668 ( .A(n48226), .B(n48227), .Z(n48191) );
  NAND U57669 ( .A(n48228), .B(n48229), .Z(n48227) );
  NAND U57670 ( .A(n48230), .B(n48231), .Z(n48226) );
  AND U57671 ( .A(n48232), .B(n48233), .Z(n48187) );
  NAND U57672 ( .A(n48234), .B(n48235), .Z(n48233) );
  NAND U57673 ( .A(n48236), .B(n48237), .Z(n48232) );
  AND U57674 ( .A(n48238), .B(n48239), .Z(n48189) );
  NAND U57675 ( .A(n48240), .B(n48241), .Z(n48183) );
  XNOR U57676 ( .A(n48166), .B(n48242), .Z(n48180) );
  XNOR U57677 ( .A(n48170), .B(n48168), .Z(n48242) );
  XOR U57678 ( .A(n48176), .B(n48243), .Z(n48168) );
  XNOR U57679 ( .A(n48173), .B(n48177), .Z(n48243) );
  AND U57680 ( .A(n48244), .B(n48245), .Z(n48177) );
  NAND U57681 ( .A(n48246), .B(n48247), .Z(n48245) );
  NAND U57682 ( .A(n48248), .B(n48249), .Z(n48244) );
  AND U57683 ( .A(n48250), .B(n48251), .Z(n48173) );
  NAND U57684 ( .A(n48252), .B(n48253), .Z(n48251) );
  NAND U57685 ( .A(n48254), .B(n48255), .Z(n48250) );
  NANDN U57686 ( .A(n48256), .B(n48257), .Z(n48176) );
  ANDN U57687 ( .B(n48258), .A(n48259), .Z(n48170) );
  XNOR U57688 ( .A(n48161), .B(n48260), .Z(n48166) );
  XNOR U57689 ( .A(n48159), .B(n48163), .Z(n48260) );
  AND U57690 ( .A(n48261), .B(n48262), .Z(n48163) );
  NAND U57691 ( .A(n48263), .B(n48264), .Z(n48262) );
  NAND U57692 ( .A(n48265), .B(n48266), .Z(n48261) );
  AND U57693 ( .A(n48267), .B(n48268), .Z(n48159) );
  NAND U57694 ( .A(n48269), .B(n48270), .Z(n48268) );
  NAND U57695 ( .A(n48271), .B(n48272), .Z(n48267) );
  AND U57696 ( .A(n48273), .B(n48274), .Z(n48161) );
  XOR U57697 ( .A(n48241), .B(n48240), .Z(N61099) );
  XNOR U57698 ( .A(n48258), .B(n48259), .Z(n48240) );
  XNOR U57699 ( .A(n48273), .B(n48274), .Z(n48259) );
  XOR U57700 ( .A(n48270), .B(n48269), .Z(n48274) );
  XOR U57701 ( .A(y[948]), .B(x[948]), .Z(n48269) );
  XOR U57702 ( .A(n48272), .B(n48271), .Z(n48270) );
  XOR U57703 ( .A(y[950]), .B(x[950]), .Z(n48271) );
  XOR U57704 ( .A(y[949]), .B(x[949]), .Z(n48272) );
  XOR U57705 ( .A(n48264), .B(n48263), .Z(n48273) );
  XOR U57706 ( .A(n48266), .B(n48265), .Z(n48263) );
  XOR U57707 ( .A(y[947]), .B(x[947]), .Z(n48265) );
  XOR U57708 ( .A(y[946]), .B(x[946]), .Z(n48266) );
  XOR U57709 ( .A(y[945]), .B(x[945]), .Z(n48264) );
  XNOR U57710 ( .A(n48257), .B(n48256), .Z(n48258) );
  XNOR U57711 ( .A(n48253), .B(n48252), .Z(n48256) );
  XOR U57712 ( .A(n48255), .B(n48254), .Z(n48252) );
  XOR U57713 ( .A(y[944]), .B(x[944]), .Z(n48254) );
  XOR U57714 ( .A(y[943]), .B(x[943]), .Z(n48255) );
  XOR U57715 ( .A(y[942]), .B(x[942]), .Z(n48253) );
  XOR U57716 ( .A(n48247), .B(n48246), .Z(n48257) );
  XOR U57717 ( .A(n48249), .B(n48248), .Z(n48246) );
  XOR U57718 ( .A(y[941]), .B(x[941]), .Z(n48248) );
  XOR U57719 ( .A(y[940]), .B(x[940]), .Z(n48249) );
  XOR U57720 ( .A(y[939]), .B(x[939]), .Z(n48247) );
  XNOR U57721 ( .A(n48223), .B(n48224), .Z(n48241) );
  XNOR U57722 ( .A(n48238), .B(n48239), .Z(n48224) );
  XOR U57723 ( .A(n48235), .B(n48234), .Z(n48239) );
  XOR U57724 ( .A(y[936]), .B(x[936]), .Z(n48234) );
  XOR U57725 ( .A(n48237), .B(n48236), .Z(n48235) );
  XOR U57726 ( .A(y[938]), .B(x[938]), .Z(n48236) );
  XOR U57727 ( .A(y[937]), .B(x[937]), .Z(n48237) );
  XOR U57728 ( .A(n48229), .B(n48228), .Z(n48238) );
  XOR U57729 ( .A(n48231), .B(n48230), .Z(n48228) );
  XOR U57730 ( .A(y[935]), .B(x[935]), .Z(n48230) );
  XOR U57731 ( .A(y[934]), .B(x[934]), .Z(n48231) );
  XOR U57732 ( .A(y[933]), .B(x[933]), .Z(n48229) );
  XNOR U57733 ( .A(n48222), .B(n48221), .Z(n48223) );
  XNOR U57734 ( .A(n48218), .B(n48217), .Z(n48221) );
  XOR U57735 ( .A(n48220), .B(n48219), .Z(n48217) );
  XOR U57736 ( .A(y[932]), .B(x[932]), .Z(n48219) );
  XOR U57737 ( .A(y[931]), .B(x[931]), .Z(n48220) );
  XOR U57738 ( .A(y[930]), .B(x[930]), .Z(n48218) );
  XOR U57739 ( .A(n48212), .B(n48211), .Z(n48222) );
  XOR U57740 ( .A(n48214), .B(n48213), .Z(n48211) );
  XOR U57741 ( .A(y[929]), .B(x[929]), .Z(n48213) );
  XOR U57742 ( .A(y[928]), .B(x[928]), .Z(n48214) );
  XOR U57743 ( .A(y[927]), .B(x[927]), .Z(n48212) );
  NAND U57744 ( .A(n48275), .B(n48276), .Z(N61090) );
  NAND U57745 ( .A(n48277), .B(n48278), .Z(n48276) );
  NANDN U57746 ( .A(n48279), .B(n48280), .Z(n48278) );
  NANDN U57747 ( .A(n48280), .B(n48279), .Z(n48275) );
  XOR U57748 ( .A(n48279), .B(n48281), .Z(N61089) );
  XNOR U57749 ( .A(n48277), .B(n48280), .Z(n48281) );
  NAND U57750 ( .A(n48282), .B(n48283), .Z(n48280) );
  NAND U57751 ( .A(n48284), .B(n48285), .Z(n48283) );
  NANDN U57752 ( .A(n48286), .B(n48287), .Z(n48285) );
  NANDN U57753 ( .A(n48287), .B(n48286), .Z(n48282) );
  AND U57754 ( .A(n48288), .B(n48289), .Z(n48277) );
  NAND U57755 ( .A(n48290), .B(n48291), .Z(n48289) );
  NANDN U57756 ( .A(n48292), .B(n48293), .Z(n48291) );
  NANDN U57757 ( .A(n48293), .B(n48292), .Z(n48288) );
  IV U57758 ( .A(n48294), .Z(n48293) );
  AND U57759 ( .A(n48295), .B(n48296), .Z(n48279) );
  NAND U57760 ( .A(n48297), .B(n48298), .Z(n48296) );
  NANDN U57761 ( .A(n48299), .B(n48300), .Z(n48298) );
  NANDN U57762 ( .A(n48300), .B(n48299), .Z(n48295) );
  XOR U57763 ( .A(n48292), .B(n48301), .Z(N61088) );
  XNOR U57764 ( .A(n48290), .B(n48294), .Z(n48301) );
  XOR U57765 ( .A(n48287), .B(n48302), .Z(n48294) );
  XNOR U57766 ( .A(n48284), .B(n48286), .Z(n48302) );
  AND U57767 ( .A(n48303), .B(n48304), .Z(n48286) );
  NANDN U57768 ( .A(n48305), .B(n48306), .Z(n48304) );
  OR U57769 ( .A(n48307), .B(n48308), .Z(n48306) );
  IV U57770 ( .A(n48309), .Z(n48308) );
  NANDN U57771 ( .A(n48309), .B(n48307), .Z(n48303) );
  AND U57772 ( .A(n48310), .B(n48311), .Z(n48284) );
  NAND U57773 ( .A(n48312), .B(n48313), .Z(n48311) );
  NANDN U57774 ( .A(n48314), .B(n48315), .Z(n48313) );
  NANDN U57775 ( .A(n48315), .B(n48314), .Z(n48310) );
  IV U57776 ( .A(n48316), .Z(n48315) );
  NAND U57777 ( .A(n48317), .B(n48318), .Z(n48287) );
  NANDN U57778 ( .A(n48319), .B(n48320), .Z(n48318) );
  NANDN U57779 ( .A(n48321), .B(n48322), .Z(n48320) );
  NANDN U57780 ( .A(n48322), .B(n48321), .Z(n48317) );
  IV U57781 ( .A(n48323), .Z(n48321) );
  AND U57782 ( .A(n48324), .B(n48325), .Z(n48290) );
  NAND U57783 ( .A(n48326), .B(n48327), .Z(n48325) );
  NANDN U57784 ( .A(n48328), .B(n48329), .Z(n48327) );
  NANDN U57785 ( .A(n48329), .B(n48328), .Z(n48324) );
  XOR U57786 ( .A(n48300), .B(n48330), .Z(n48292) );
  XNOR U57787 ( .A(n48297), .B(n48299), .Z(n48330) );
  AND U57788 ( .A(n48331), .B(n48332), .Z(n48299) );
  NANDN U57789 ( .A(n48333), .B(n48334), .Z(n48332) );
  OR U57790 ( .A(n48335), .B(n48336), .Z(n48334) );
  IV U57791 ( .A(n48337), .Z(n48336) );
  NANDN U57792 ( .A(n48337), .B(n48335), .Z(n48331) );
  AND U57793 ( .A(n48338), .B(n48339), .Z(n48297) );
  NAND U57794 ( .A(n48340), .B(n48341), .Z(n48339) );
  NANDN U57795 ( .A(n48342), .B(n48343), .Z(n48341) );
  NANDN U57796 ( .A(n48343), .B(n48342), .Z(n48338) );
  IV U57797 ( .A(n48344), .Z(n48343) );
  NAND U57798 ( .A(n48345), .B(n48346), .Z(n48300) );
  NANDN U57799 ( .A(n48347), .B(n48348), .Z(n48346) );
  NANDN U57800 ( .A(n48349), .B(n48350), .Z(n48348) );
  NANDN U57801 ( .A(n48350), .B(n48349), .Z(n48345) );
  IV U57802 ( .A(n48351), .Z(n48349) );
  XOR U57803 ( .A(n48326), .B(n48352), .Z(N61087) );
  XNOR U57804 ( .A(n48329), .B(n48328), .Z(n48352) );
  XNOR U57805 ( .A(n48340), .B(n48353), .Z(n48328) );
  XNOR U57806 ( .A(n48344), .B(n48342), .Z(n48353) );
  XOR U57807 ( .A(n48350), .B(n48354), .Z(n48342) );
  XNOR U57808 ( .A(n48347), .B(n48351), .Z(n48354) );
  AND U57809 ( .A(n48355), .B(n48356), .Z(n48351) );
  NAND U57810 ( .A(n48357), .B(n48358), .Z(n48356) );
  NAND U57811 ( .A(n48359), .B(n48360), .Z(n48355) );
  AND U57812 ( .A(n48361), .B(n48362), .Z(n48347) );
  NAND U57813 ( .A(n48363), .B(n48364), .Z(n48362) );
  NAND U57814 ( .A(n48365), .B(n48366), .Z(n48361) );
  NANDN U57815 ( .A(n48367), .B(n48368), .Z(n48350) );
  ANDN U57816 ( .B(n48369), .A(n48370), .Z(n48344) );
  XNOR U57817 ( .A(n48335), .B(n48371), .Z(n48340) );
  XNOR U57818 ( .A(n48333), .B(n48337), .Z(n48371) );
  AND U57819 ( .A(n48372), .B(n48373), .Z(n48337) );
  NAND U57820 ( .A(n48374), .B(n48375), .Z(n48373) );
  NAND U57821 ( .A(n48376), .B(n48377), .Z(n48372) );
  AND U57822 ( .A(n48378), .B(n48379), .Z(n48333) );
  NAND U57823 ( .A(n48380), .B(n48381), .Z(n48379) );
  NAND U57824 ( .A(n48382), .B(n48383), .Z(n48378) );
  AND U57825 ( .A(n48384), .B(n48385), .Z(n48335) );
  NAND U57826 ( .A(n48386), .B(n48387), .Z(n48329) );
  XNOR U57827 ( .A(n48312), .B(n48388), .Z(n48326) );
  XNOR U57828 ( .A(n48316), .B(n48314), .Z(n48388) );
  XOR U57829 ( .A(n48322), .B(n48389), .Z(n48314) );
  XNOR U57830 ( .A(n48319), .B(n48323), .Z(n48389) );
  AND U57831 ( .A(n48390), .B(n48391), .Z(n48323) );
  NAND U57832 ( .A(n48392), .B(n48393), .Z(n48391) );
  NAND U57833 ( .A(n48394), .B(n48395), .Z(n48390) );
  AND U57834 ( .A(n48396), .B(n48397), .Z(n48319) );
  NAND U57835 ( .A(n48398), .B(n48399), .Z(n48397) );
  NAND U57836 ( .A(n48400), .B(n48401), .Z(n48396) );
  NANDN U57837 ( .A(n48402), .B(n48403), .Z(n48322) );
  ANDN U57838 ( .B(n48404), .A(n48405), .Z(n48316) );
  XNOR U57839 ( .A(n48307), .B(n48406), .Z(n48312) );
  XNOR U57840 ( .A(n48305), .B(n48309), .Z(n48406) );
  AND U57841 ( .A(n48407), .B(n48408), .Z(n48309) );
  NAND U57842 ( .A(n48409), .B(n48410), .Z(n48408) );
  NAND U57843 ( .A(n48411), .B(n48412), .Z(n48407) );
  AND U57844 ( .A(n48413), .B(n48414), .Z(n48305) );
  NAND U57845 ( .A(n48415), .B(n48416), .Z(n48414) );
  NAND U57846 ( .A(n48417), .B(n48418), .Z(n48413) );
  AND U57847 ( .A(n48419), .B(n48420), .Z(n48307) );
  XOR U57848 ( .A(n48387), .B(n48386), .Z(N61086) );
  XNOR U57849 ( .A(n48404), .B(n48405), .Z(n48386) );
  XNOR U57850 ( .A(n48419), .B(n48420), .Z(n48405) );
  XOR U57851 ( .A(n48416), .B(n48415), .Z(n48420) );
  XOR U57852 ( .A(y[924]), .B(x[924]), .Z(n48415) );
  XOR U57853 ( .A(n48418), .B(n48417), .Z(n48416) );
  XOR U57854 ( .A(y[926]), .B(x[926]), .Z(n48417) );
  XOR U57855 ( .A(y[925]), .B(x[925]), .Z(n48418) );
  XOR U57856 ( .A(n48410), .B(n48409), .Z(n48419) );
  XOR U57857 ( .A(n48412), .B(n48411), .Z(n48409) );
  XOR U57858 ( .A(y[923]), .B(x[923]), .Z(n48411) );
  XOR U57859 ( .A(y[922]), .B(x[922]), .Z(n48412) );
  XOR U57860 ( .A(y[921]), .B(x[921]), .Z(n48410) );
  XNOR U57861 ( .A(n48403), .B(n48402), .Z(n48404) );
  XNOR U57862 ( .A(n48399), .B(n48398), .Z(n48402) );
  XOR U57863 ( .A(n48401), .B(n48400), .Z(n48398) );
  XOR U57864 ( .A(y[920]), .B(x[920]), .Z(n48400) );
  XOR U57865 ( .A(y[919]), .B(x[919]), .Z(n48401) );
  XOR U57866 ( .A(y[918]), .B(x[918]), .Z(n48399) );
  XOR U57867 ( .A(n48393), .B(n48392), .Z(n48403) );
  XOR U57868 ( .A(n48395), .B(n48394), .Z(n48392) );
  XOR U57869 ( .A(y[917]), .B(x[917]), .Z(n48394) );
  XOR U57870 ( .A(y[916]), .B(x[916]), .Z(n48395) );
  XOR U57871 ( .A(y[915]), .B(x[915]), .Z(n48393) );
  XNOR U57872 ( .A(n48369), .B(n48370), .Z(n48387) );
  XNOR U57873 ( .A(n48384), .B(n48385), .Z(n48370) );
  XOR U57874 ( .A(n48381), .B(n48380), .Z(n48385) );
  XOR U57875 ( .A(y[912]), .B(x[912]), .Z(n48380) );
  XOR U57876 ( .A(n48383), .B(n48382), .Z(n48381) );
  XOR U57877 ( .A(y[914]), .B(x[914]), .Z(n48382) );
  XOR U57878 ( .A(y[913]), .B(x[913]), .Z(n48383) );
  XOR U57879 ( .A(n48375), .B(n48374), .Z(n48384) );
  XOR U57880 ( .A(n48377), .B(n48376), .Z(n48374) );
  XOR U57881 ( .A(y[911]), .B(x[911]), .Z(n48376) );
  XOR U57882 ( .A(y[910]), .B(x[910]), .Z(n48377) );
  XOR U57883 ( .A(y[909]), .B(x[909]), .Z(n48375) );
  XNOR U57884 ( .A(n48368), .B(n48367), .Z(n48369) );
  XNOR U57885 ( .A(n48364), .B(n48363), .Z(n48367) );
  XOR U57886 ( .A(n48366), .B(n48365), .Z(n48363) );
  XOR U57887 ( .A(y[908]), .B(x[908]), .Z(n48365) );
  XOR U57888 ( .A(y[907]), .B(x[907]), .Z(n48366) );
  XOR U57889 ( .A(y[906]), .B(x[906]), .Z(n48364) );
  XOR U57890 ( .A(n48358), .B(n48357), .Z(n48368) );
  XOR U57891 ( .A(n48360), .B(n48359), .Z(n48357) );
  XOR U57892 ( .A(y[905]), .B(x[905]), .Z(n48359) );
  XOR U57893 ( .A(y[904]), .B(x[904]), .Z(n48360) );
  XOR U57894 ( .A(y[903]), .B(x[903]), .Z(n48358) );
  NAND U57895 ( .A(n48421), .B(n48422), .Z(N61077) );
  NAND U57896 ( .A(n48423), .B(n48424), .Z(n48422) );
  NANDN U57897 ( .A(n48425), .B(n48426), .Z(n48424) );
  NANDN U57898 ( .A(n48426), .B(n48425), .Z(n48421) );
  XOR U57899 ( .A(n48425), .B(n48427), .Z(N61076) );
  XNOR U57900 ( .A(n48423), .B(n48426), .Z(n48427) );
  NAND U57901 ( .A(n48428), .B(n48429), .Z(n48426) );
  NAND U57902 ( .A(n48430), .B(n48431), .Z(n48429) );
  NANDN U57903 ( .A(n48432), .B(n48433), .Z(n48431) );
  NANDN U57904 ( .A(n48433), .B(n48432), .Z(n48428) );
  AND U57905 ( .A(n48434), .B(n48435), .Z(n48423) );
  NAND U57906 ( .A(n48436), .B(n48437), .Z(n48435) );
  NANDN U57907 ( .A(n48438), .B(n48439), .Z(n48437) );
  NANDN U57908 ( .A(n48439), .B(n48438), .Z(n48434) );
  IV U57909 ( .A(n48440), .Z(n48439) );
  AND U57910 ( .A(n48441), .B(n48442), .Z(n48425) );
  NAND U57911 ( .A(n48443), .B(n48444), .Z(n48442) );
  NANDN U57912 ( .A(n48445), .B(n48446), .Z(n48444) );
  NANDN U57913 ( .A(n48446), .B(n48445), .Z(n48441) );
  XOR U57914 ( .A(n48438), .B(n48447), .Z(N61075) );
  XNOR U57915 ( .A(n48436), .B(n48440), .Z(n48447) );
  XOR U57916 ( .A(n48433), .B(n48448), .Z(n48440) );
  XNOR U57917 ( .A(n48430), .B(n48432), .Z(n48448) );
  AND U57918 ( .A(n48449), .B(n48450), .Z(n48432) );
  NANDN U57919 ( .A(n48451), .B(n48452), .Z(n48450) );
  OR U57920 ( .A(n48453), .B(n48454), .Z(n48452) );
  IV U57921 ( .A(n48455), .Z(n48454) );
  NANDN U57922 ( .A(n48455), .B(n48453), .Z(n48449) );
  AND U57923 ( .A(n48456), .B(n48457), .Z(n48430) );
  NAND U57924 ( .A(n48458), .B(n48459), .Z(n48457) );
  NANDN U57925 ( .A(n48460), .B(n48461), .Z(n48459) );
  NANDN U57926 ( .A(n48461), .B(n48460), .Z(n48456) );
  IV U57927 ( .A(n48462), .Z(n48461) );
  NAND U57928 ( .A(n48463), .B(n48464), .Z(n48433) );
  NANDN U57929 ( .A(n48465), .B(n48466), .Z(n48464) );
  NANDN U57930 ( .A(n48467), .B(n48468), .Z(n48466) );
  NANDN U57931 ( .A(n48468), .B(n48467), .Z(n48463) );
  IV U57932 ( .A(n48469), .Z(n48467) );
  AND U57933 ( .A(n48470), .B(n48471), .Z(n48436) );
  NAND U57934 ( .A(n48472), .B(n48473), .Z(n48471) );
  NANDN U57935 ( .A(n48474), .B(n48475), .Z(n48473) );
  NANDN U57936 ( .A(n48475), .B(n48474), .Z(n48470) );
  XOR U57937 ( .A(n48446), .B(n48476), .Z(n48438) );
  XNOR U57938 ( .A(n48443), .B(n48445), .Z(n48476) );
  AND U57939 ( .A(n48477), .B(n48478), .Z(n48445) );
  NANDN U57940 ( .A(n48479), .B(n48480), .Z(n48478) );
  OR U57941 ( .A(n48481), .B(n48482), .Z(n48480) );
  IV U57942 ( .A(n48483), .Z(n48482) );
  NANDN U57943 ( .A(n48483), .B(n48481), .Z(n48477) );
  AND U57944 ( .A(n48484), .B(n48485), .Z(n48443) );
  NAND U57945 ( .A(n48486), .B(n48487), .Z(n48485) );
  NANDN U57946 ( .A(n48488), .B(n48489), .Z(n48487) );
  NANDN U57947 ( .A(n48489), .B(n48488), .Z(n48484) );
  IV U57948 ( .A(n48490), .Z(n48489) );
  NAND U57949 ( .A(n48491), .B(n48492), .Z(n48446) );
  NANDN U57950 ( .A(n48493), .B(n48494), .Z(n48492) );
  NANDN U57951 ( .A(n48495), .B(n48496), .Z(n48494) );
  NANDN U57952 ( .A(n48496), .B(n48495), .Z(n48491) );
  IV U57953 ( .A(n48497), .Z(n48495) );
  XOR U57954 ( .A(n48472), .B(n48498), .Z(N61074) );
  XNOR U57955 ( .A(n48475), .B(n48474), .Z(n48498) );
  XNOR U57956 ( .A(n48486), .B(n48499), .Z(n48474) );
  XNOR U57957 ( .A(n48490), .B(n48488), .Z(n48499) );
  XOR U57958 ( .A(n48496), .B(n48500), .Z(n48488) );
  XNOR U57959 ( .A(n48493), .B(n48497), .Z(n48500) );
  AND U57960 ( .A(n48501), .B(n48502), .Z(n48497) );
  NAND U57961 ( .A(n48503), .B(n48504), .Z(n48502) );
  NAND U57962 ( .A(n48505), .B(n48506), .Z(n48501) );
  AND U57963 ( .A(n48507), .B(n48508), .Z(n48493) );
  NAND U57964 ( .A(n48509), .B(n48510), .Z(n48508) );
  NAND U57965 ( .A(n48511), .B(n48512), .Z(n48507) );
  NANDN U57966 ( .A(n48513), .B(n48514), .Z(n48496) );
  ANDN U57967 ( .B(n48515), .A(n48516), .Z(n48490) );
  XNOR U57968 ( .A(n48481), .B(n48517), .Z(n48486) );
  XNOR U57969 ( .A(n48479), .B(n48483), .Z(n48517) );
  AND U57970 ( .A(n48518), .B(n48519), .Z(n48483) );
  NAND U57971 ( .A(n48520), .B(n48521), .Z(n48519) );
  NAND U57972 ( .A(n48522), .B(n48523), .Z(n48518) );
  AND U57973 ( .A(n48524), .B(n48525), .Z(n48479) );
  NAND U57974 ( .A(n48526), .B(n48527), .Z(n48525) );
  NAND U57975 ( .A(n48528), .B(n48529), .Z(n48524) );
  AND U57976 ( .A(n48530), .B(n48531), .Z(n48481) );
  NAND U57977 ( .A(n48532), .B(n48533), .Z(n48475) );
  XNOR U57978 ( .A(n48458), .B(n48534), .Z(n48472) );
  XNOR U57979 ( .A(n48462), .B(n48460), .Z(n48534) );
  XOR U57980 ( .A(n48468), .B(n48535), .Z(n48460) );
  XNOR U57981 ( .A(n48465), .B(n48469), .Z(n48535) );
  AND U57982 ( .A(n48536), .B(n48537), .Z(n48469) );
  NAND U57983 ( .A(n48538), .B(n48539), .Z(n48537) );
  NAND U57984 ( .A(n48540), .B(n48541), .Z(n48536) );
  AND U57985 ( .A(n48542), .B(n48543), .Z(n48465) );
  NAND U57986 ( .A(n48544), .B(n48545), .Z(n48543) );
  NAND U57987 ( .A(n48546), .B(n48547), .Z(n48542) );
  NANDN U57988 ( .A(n48548), .B(n48549), .Z(n48468) );
  ANDN U57989 ( .B(n48550), .A(n48551), .Z(n48462) );
  XNOR U57990 ( .A(n48453), .B(n48552), .Z(n48458) );
  XNOR U57991 ( .A(n48451), .B(n48455), .Z(n48552) );
  AND U57992 ( .A(n48553), .B(n48554), .Z(n48455) );
  NAND U57993 ( .A(n48555), .B(n48556), .Z(n48554) );
  NAND U57994 ( .A(n48557), .B(n48558), .Z(n48553) );
  AND U57995 ( .A(n48559), .B(n48560), .Z(n48451) );
  NAND U57996 ( .A(n48561), .B(n48562), .Z(n48560) );
  NAND U57997 ( .A(n48563), .B(n48564), .Z(n48559) );
  AND U57998 ( .A(n48565), .B(n48566), .Z(n48453) );
  XOR U57999 ( .A(n48533), .B(n48532), .Z(N61073) );
  XNOR U58000 ( .A(n48550), .B(n48551), .Z(n48532) );
  XNOR U58001 ( .A(n48565), .B(n48566), .Z(n48551) );
  XOR U58002 ( .A(n48562), .B(n48561), .Z(n48566) );
  XOR U58003 ( .A(y[900]), .B(x[900]), .Z(n48561) );
  XOR U58004 ( .A(n48564), .B(n48563), .Z(n48562) );
  XOR U58005 ( .A(y[902]), .B(x[902]), .Z(n48563) );
  XOR U58006 ( .A(y[901]), .B(x[901]), .Z(n48564) );
  XOR U58007 ( .A(n48556), .B(n48555), .Z(n48565) );
  XOR U58008 ( .A(n48558), .B(n48557), .Z(n48555) );
  XOR U58009 ( .A(y[899]), .B(x[899]), .Z(n48557) );
  XOR U58010 ( .A(y[898]), .B(x[898]), .Z(n48558) );
  XOR U58011 ( .A(y[897]), .B(x[897]), .Z(n48556) );
  XNOR U58012 ( .A(n48549), .B(n48548), .Z(n48550) );
  XNOR U58013 ( .A(n48545), .B(n48544), .Z(n48548) );
  XOR U58014 ( .A(n48547), .B(n48546), .Z(n48544) );
  XOR U58015 ( .A(y[896]), .B(x[896]), .Z(n48546) );
  XOR U58016 ( .A(y[895]), .B(x[895]), .Z(n48547) );
  XOR U58017 ( .A(y[894]), .B(x[894]), .Z(n48545) );
  XOR U58018 ( .A(n48539), .B(n48538), .Z(n48549) );
  XOR U58019 ( .A(n48541), .B(n48540), .Z(n48538) );
  XOR U58020 ( .A(y[893]), .B(x[893]), .Z(n48540) );
  XOR U58021 ( .A(y[892]), .B(x[892]), .Z(n48541) );
  XOR U58022 ( .A(y[891]), .B(x[891]), .Z(n48539) );
  XNOR U58023 ( .A(n48515), .B(n48516), .Z(n48533) );
  XNOR U58024 ( .A(n48530), .B(n48531), .Z(n48516) );
  XOR U58025 ( .A(n48527), .B(n48526), .Z(n48531) );
  XOR U58026 ( .A(y[888]), .B(x[888]), .Z(n48526) );
  XOR U58027 ( .A(n48529), .B(n48528), .Z(n48527) );
  XOR U58028 ( .A(y[890]), .B(x[890]), .Z(n48528) );
  XOR U58029 ( .A(y[889]), .B(x[889]), .Z(n48529) );
  XOR U58030 ( .A(n48521), .B(n48520), .Z(n48530) );
  XOR U58031 ( .A(n48523), .B(n48522), .Z(n48520) );
  XOR U58032 ( .A(y[887]), .B(x[887]), .Z(n48522) );
  XOR U58033 ( .A(y[886]), .B(x[886]), .Z(n48523) );
  XOR U58034 ( .A(y[885]), .B(x[885]), .Z(n48521) );
  XNOR U58035 ( .A(n48514), .B(n48513), .Z(n48515) );
  XNOR U58036 ( .A(n48510), .B(n48509), .Z(n48513) );
  XOR U58037 ( .A(n48512), .B(n48511), .Z(n48509) );
  XOR U58038 ( .A(y[884]), .B(x[884]), .Z(n48511) );
  XOR U58039 ( .A(y[883]), .B(x[883]), .Z(n48512) );
  XOR U58040 ( .A(y[882]), .B(x[882]), .Z(n48510) );
  XOR U58041 ( .A(n48504), .B(n48503), .Z(n48514) );
  XOR U58042 ( .A(n48506), .B(n48505), .Z(n48503) );
  XOR U58043 ( .A(y[881]), .B(x[881]), .Z(n48505) );
  XOR U58044 ( .A(y[880]), .B(x[880]), .Z(n48506) );
  XOR U58045 ( .A(y[879]), .B(x[879]), .Z(n48504) );
  NAND U58046 ( .A(n48567), .B(n48568), .Z(N61064) );
  NAND U58047 ( .A(n48569), .B(n48570), .Z(n48568) );
  NANDN U58048 ( .A(n48571), .B(n48572), .Z(n48570) );
  NANDN U58049 ( .A(n48572), .B(n48571), .Z(n48567) );
  XOR U58050 ( .A(n48571), .B(n48573), .Z(N61063) );
  XNOR U58051 ( .A(n48569), .B(n48572), .Z(n48573) );
  NAND U58052 ( .A(n48574), .B(n48575), .Z(n48572) );
  NAND U58053 ( .A(n48576), .B(n48577), .Z(n48575) );
  NANDN U58054 ( .A(n48578), .B(n48579), .Z(n48577) );
  NANDN U58055 ( .A(n48579), .B(n48578), .Z(n48574) );
  AND U58056 ( .A(n48580), .B(n48581), .Z(n48569) );
  NAND U58057 ( .A(n48582), .B(n48583), .Z(n48581) );
  NANDN U58058 ( .A(n48584), .B(n48585), .Z(n48583) );
  NANDN U58059 ( .A(n48585), .B(n48584), .Z(n48580) );
  IV U58060 ( .A(n48586), .Z(n48585) );
  AND U58061 ( .A(n48587), .B(n48588), .Z(n48571) );
  NAND U58062 ( .A(n48589), .B(n48590), .Z(n48588) );
  NANDN U58063 ( .A(n48591), .B(n48592), .Z(n48590) );
  NANDN U58064 ( .A(n48592), .B(n48591), .Z(n48587) );
  XOR U58065 ( .A(n48584), .B(n48593), .Z(N61062) );
  XNOR U58066 ( .A(n48582), .B(n48586), .Z(n48593) );
  XOR U58067 ( .A(n48579), .B(n48594), .Z(n48586) );
  XNOR U58068 ( .A(n48576), .B(n48578), .Z(n48594) );
  AND U58069 ( .A(n48595), .B(n48596), .Z(n48578) );
  NANDN U58070 ( .A(n48597), .B(n48598), .Z(n48596) );
  OR U58071 ( .A(n48599), .B(n48600), .Z(n48598) );
  IV U58072 ( .A(n48601), .Z(n48600) );
  NANDN U58073 ( .A(n48601), .B(n48599), .Z(n48595) );
  AND U58074 ( .A(n48602), .B(n48603), .Z(n48576) );
  NAND U58075 ( .A(n48604), .B(n48605), .Z(n48603) );
  NANDN U58076 ( .A(n48606), .B(n48607), .Z(n48605) );
  NANDN U58077 ( .A(n48607), .B(n48606), .Z(n48602) );
  IV U58078 ( .A(n48608), .Z(n48607) );
  NAND U58079 ( .A(n48609), .B(n48610), .Z(n48579) );
  NANDN U58080 ( .A(n48611), .B(n48612), .Z(n48610) );
  NANDN U58081 ( .A(n48613), .B(n48614), .Z(n48612) );
  NANDN U58082 ( .A(n48614), .B(n48613), .Z(n48609) );
  IV U58083 ( .A(n48615), .Z(n48613) );
  AND U58084 ( .A(n48616), .B(n48617), .Z(n48582) );
  NAND U58085 ( .A(n48618), .B(n48619), .Z(n48617) );
  NANDN U58086 ( .A(n48620), .B(n48621), .Z(n48619) );
  NANDN U58087 ( .A(n48621), .B(n48620), .Z(n48616) );
  XOR U58088 ( .A(n48592), .B(n48622), .Z(n48584) );
  XNOR U58089 ( .A(n48589), .B(n48591), .Z(n48622) );
  AND U58090 ( .A(n48623), .B(n48624), .Z(n48591) );
  NANDN U58091 ( .A(n48625), .B(n48626), .Z(n48624) );
  OR U58092 ( .A(n48627), .B(n48628), .Z(n48626) );
  IV U58093 ( .A(n48629), .Z(n48628) );
  NANDN U58094 ( .A(n48629), .B(n48627), .Z(n48623) );
  AND U58095 ( .A(n48630), .B(n48631), .Z(n48589) );
  NAND U58096 ( .A(n48632), .B(n48633), .Z(n48631) );
  NANDN U58097 ( .A(n48634), .B(n48635), .Z(n48633) );
  NANDN U58098 ( .A(n48635), .B(n48634), .Z(n48630) );
  IV U58099 ( .A(n48636), .Z(n48635) );
  NAND U58100 ( .A(n48637), .B(n48638), .Z(n48592) );
  NANDN U58101 ( .A(n48639), .B(n48640), .Z(n48638) );
  NANDN U58102 ( .A(n48641), .B(n48642), .Z(n48640) );
  NANDN U58103 ( .A(n48642), .B(n48641), .Z(n48637) );
  IV U58104 ( .A(n48643), .Z(n48641) );
  XOR U58105 ( .A(n48618), .B(n48644), .Z(N61061) );
  XNOR U58106 ( .A(n48621), .B(n48620), .Z(n48644) );
  XNOR U58107 ( .A(n48632), .B(n48645), .Z(n48620) );
  XNOR U58108 ( .A(n48636), .B(n48634), .Z(n48645) );
  XOR U58109 ( .A(n48642), .B(n48646), .Z(n48634) );
  XNOR U58110 ( .A(n48639), .B(n48643), .Z(n48646) );
  AND U58111 ( .A(n48647), .B(n48648), .Z(n48643) );
  NAND U58112 ( .A(n48649), .B(n48650), .Z(n48648) );
  NAND U58113 ( .A(n48651), .B(n48652), .Z(n48647) );
  AND U58114 ( .A(n48653), .B(n48654), .Z(n48639) );
  NAND U58115 ( .A(n48655), .B(n48656), .Z(n48654) );
  NAND U58116 ( .A(n48657), .B(n48658), .Z(n48653) );
  NANDN U58117 ( .A(n48659), .B(n48660), .Z(n48642) );
  ANDN U58118 ( .B(n48661), .A(n48662), .Z(n48636) );
  XNOR U58119 ( .A(n48627), .B(n48663), .Z(n48632) );
  XNOR U58120 ( .A(n48625), .B(n48629), .Z(n48663) );
  AND U58121 ( .A(n48664), .B(n48665), .Z(n48629) );
  NAND U58122 ( .A(n48666), .B(n48667), .Z(n48665) );
  NAND U58123 ( .A(n48668), .B(n48669), .Z(n48664) );
  AND U58124 ( .A(n48670), .B(n48671), .Z(n48625) );
  NAND U58125 ( .A(n48672), .B(n48673), .Z(n48671) );
  NAND U58126 ( .A(n48674), .B(n48675), .Z(n48670) );
  AND U58127 ( .A(n48676), .B(n48677), .Z(n48627) );
  NAND U58128 ( .A(n48678), .B(n48679), .Z(n48621) );
  XNOR U58129 ( .A(n48604), .B(n48680), .Z(n48618) );
  XNOR U58130 ( .A(n48608), .B(n48606), .Z(n48680) );
  XOR U58131 ( .A(n48614), .B(n48681), .Z(n48606) );
  XNOR U58132 ( .A(n48611), .B(n48615), .Z(n48681) );
  AND U58133 ( .A(n48682), .B(n48683), .Z(n48615) );
  NAND U58134 ( .A(n48684), .B(n48685), .Z(n48683) );
  NAND U58135 ( .A(n48686), .B(n48687), .Z(n48682) );
  AND U58136 ( .A(n48688), .B(n48689), .Z(n48611) );
  NAND U58137 ( .A(n48690), .B(n48691), .Z(n48689) );
  NAND U58138 ( .A(n48692), .B(n48693), .Z(n48688) );
  NANDN U58139 ( .A(n48694), .B(n48695), .Z(n48614) );
  ANDN U58140 ( .B(n48696), .A(n48697), .Z(n48608) );
  XNOR U58141 ( .A(n48599), .B(n48698), .Z(n48604) );
  XNOR U58142 ( .A(n48597), .B(n48601), .Z(n48698) );
  AND U58143 ( .A(n48699), .B(n48700), .Z(n48601) );
  NAND U58144 ( .A(n48701), .B(n48702), .Z(n48700) );
  NAND U58145 ( .A(n48703), .B(n48704), .Z(n48699) );
  AND U58146 ( .A(n48705), .B(n48706), .Z(n48597) );
  NAND U58147 ( .A(n48707), .B(n48708), .Z(n48706) );
  NAND U58148 ( .A(n48709), .B(n48710), .Z(n48705) );
  AND U58149 ( .A(n48711), .B(n48712), .Z(n48599) );
  XOR U58150 ( .A(n48679), .B(n48678), .Z(N61060) );
  XNOR U58151 ( .A(n48696), .B(n48697), .Z(n48678) );
  XNOR U58152 ( .A(n48711), .B(n48712), .Z(n48697) );
  XOR U58153 ( .A(n48708), .B(n48707), .Z(n48712) );
  XOR U58154 ( .A(y[876]), .B(x[876]), .Z(n48707) );
  XOR U58155 ( .A(n48710), .B(n48709), .Z(n48708) );
  XOR U58156 ( .A(y[878]), .B(x[878]), .Z(n48709) );
  XOR U58157 ( .A(y[877]), .B(x[877]), .Z(n48710) );
  XOR U58158 ( .A(n48702), .B(n48701), .Z(n48711) );
  XOR U58159 ( .A(n48704), .B(n48703), .Z(n48701) );
  XOR U58160 ( .A(y[875]), .B(x[875]), .Z(n48703) );
  XOR U58161 ( .A(y[874]), .B(x[874]), .Z(n48704) );
  XOR U58162 ( .A(y[873]), .B(x[873]), .Z(n48702) );
  XNOR U58163 ( .A(n48695), .B(n48694), .Z(n48696) );
  XNOR U58164 ( .A(n48691), .B(n48690), .Z(n48694) );
  XOR U58165 ( .A(n48693), .B(n48692), .Z(n48690) );
  XOR U58166 ( .A(y[872]), .B(x[872]), .Z(n48692) );
  XOR U58167 ( .A(y[871]), .B(x[871]), .Z(n48693) );
  XOR U58168 ( .A(y[870]), .B(x[870]), .Z(n48691) );
  XOR U58169 ( .A(n48685), .B(n48684), .Z(n48695) );
  XOR U58170 ( .A(n48687), .B(n48686), .Z(n48684) );
  XOR U58171 ( .A(y[869]), .B(x[869]), .Z(n48686) );
  XOR U58172 ( .A(y[868]), .B(x[868]), .Z(n48687) );
  XOR U58173 ( .A(y[867]), .B(x[867]), .Z(n48685) );
  XNOR U58174 ( .A(n48661), .B(n48662), .Z(n48679) );
  XNOR U58175 ( .A(n48676), .B(n48677), .Z(n48662) );
  XOR U58176 ( .A(n48673), .B(n48672), .Z(n48677) );
  XOR U58177 ( .A(y[864]), .B(x[864]), .Z(n48672) );
  XOR U58178 ( .A(n48675), .B(n48674), .Z(n48673) );
  XOR U58179 ( .A(y[866]), .B(x[866]), .Z(n48674) );
  XOR U58180 ( .A(y[865]), .B(x[865]), .Z(n48675) );
  XOR U58181 ( .A(n48667), .B(n48666), .Z(n48676) );
  XOR U58182 ( .A(n48669), .B(n48668), .Z(n48666) );
  XOR U58183 ( .A(y[863]), .B(x[863]), .Z(n48668) );
  XOR U58184 ( .A(y[862]), .B(x[862]), .Z(n48669) );
  XOR U58185 ( .A(y[861]), .B(x[861]), .Z(n48667) );
  XNOR U58186 ( .A(n48660), .B(n48659), .Z(n48661) );
  XNOR U58187 ( .A(n48656), .B(n48655), .Z(n48659) );
  XOR U58188 ( .A(n48658), .B(n48657), .Z(n48655) );
  XOR U58189 ( .A(y[860]), .B(x[860]), .Z(n48657) );
  XOR U58190 ( .A(y[859]), .B(x[859]), .Z(n48658) );
  XOR U58191 ( .A(y[858]), .B(x[858]), .Z(n48656) );
  XOR U58192 ( .A(n48650), .B(n48649), .Z(n48660) );
  XOR U58193 ( .A(n48652), .B(n48651), .Z(n48649) );
  XOR U58194 ( .A(y[857]), .B(x[857]), .Z(n48651) );
  XOR U58195 ( .A(y[856]), .B(x[856]), .Z(n48652) );
  XOR U58196 ( .A(y[855]), .B(x[855]), .Z(n48650) );
  NAND U58197 ( .A(n48713), .B(n48714), .Z(N61051) );
  NAND U58198 ( .A(n48715), .B(n48716), .Z(n48714) );
  NANDN U58199 ( .A(n48717), .B(n48718), .Z(n48716) );
  NANDN U58200 ( .A(n48718), .B(n48717), .Z(n48713) );
  XOR U58201 ( .A(n48717), .B(n48719), .Z(N61050) );
  XNOR U58202 ( .A(n48715), .B(n48718), .Z(n48719) );
  NAND U58203 ( .A(n48720), .B(n48721), .Z(n48718) );
  NAND U58204 ( .A(n48722), .B(n48723), .Z(n48721) );
  NANDN U58205 ( .A(n48724), .B(n48725), .Z(n48723) );
  NANDN U58206 ( .A(n48725), .B(n48724), .Z(n48720) );
  AND U58207 ( .A(n48726), .B(n48727), .Z(n48715) );
  NAND U58208 ( .A(n48728), .B(n48729), .Z(n48727) );
  NANDN U58209 ( .A(n48730), .B(n48731), .Z(n48729) );
  NANDN U58210 ( .A(n48731), .B(n48730), .Z(n48726) );
  IV U58211 ( .A(n48732), .Z(n48731) );
  AND U58212 ( .A(n48733), .B(n48734), .Z(n48717) );
  NAND U58213 ( .A(n48735), .B(n48736), .Z(n48734) );
  NANDN U58214 ( .A(n48737), .B(n48738), .Z(n48736) );
  NANDN U58215 ( .A(n48738), .B(n48737), .Z(n48733) );
  XOR U58216 ( .A(n48730), .B(n48739), .Z(N61049) );
  XNOR U58217 ( .A(n48728), .B(n48732), .Z(n48739) );
  XOR U58218 ( .A(n48725), .B(n48740), .Z(n48732) );
  XNOR U58219 ( .A(n48722), .B(n48724), .Z(n48740) );
  AND U58220 ( .A(n48741), .B(n48742), .Z(n48724) );
  NANDN U58221 ( .A(n48743), .B(n48744), .Z(n48742) );
  OR U58222 ( .A(n48745), .B(n48746), .Z(n48744) );
  IV U58223 ( .A(n48747), .Z(n48746) );
  NANDN U58224 ( .A(n48747), .B(n48745), .Z(n48741) );
  AND U58225 ( .A(n48748), .B(n48749), .Z(n48722) );
  NAND U58226 ( .A(n48750), .B(n48751), .Z(n48749) );
  NANDN U58227 ( .A(n48752), .B(n48753), .Z(n48751) );
  NANDN U58228 ( .A(n48753), .B(n48752), .Z(n48748) );
  IV U58229 ( .A(n48754), .Z(n48753) );
  NAND U58230 ( .A(n48755), .B(n48756), .Z(n48725) );
  NANDN U58231 ( .A(n48757), .B(n48758), .Z(n48756) );
  NANDN U58232 ( .A(n48759), .B(n48760), .Z(n48758) );
  NANDN U58233 ( .A(n48760), .B(n48759), .Z(n48755) );
  IV U58234 ( .A(n48761), .Z(n48759) );
  AND U58235 ( .A(n48762), .B(n48763), .Z(n48728) );
  NAND U58236 ( .A(n48764), .B(n48765), .Z(n48763) );
  NANDN U58237 ( .A(n48766), .B(n48767), .Z(n48765) );
  NANDN U58238 ( .A(n48767), .B(n48766), .Z(n48762) );
  XOR U58239 ( .A(n48738), .B(n48768), .Z(n48730) );
  XNOR U58240 ( .A(n48735), .B(n48737), .Z(n48768) );
  AND U58241 ( .A(n48769), .B(n48770), .Z(n48737) );
  NANDN U58242 ( .A(n48771), .B(n48772), .Z(n48770) );
  OR U58243 ( .A(n48773), .B(n48774), .Z(n48772) );
  IV U58244 ( .A(n48775), .Z(n48774) );
  NANDN U58245 ( .A(n48775), .B(n48773), .Z(n48769) );
  AND U58246 ( .A(n48776), .B(n48777), .Z(n48735) );
  NAND U58247 ( .A(n48778), .B(n48779), .Z(n48777) );
  NANDN U58248 ( .A(n48780), .B(n48781), .Z(n48779) );
  NANDN U58249 ( .A(n48781), .B(n48780), .Z(n48776) );
  IV U58250 ( .A(n48782), .Z(n48781) );
  NAND U58251 ( .A(n48783), .B(n48784), .Z(n48738) );
  NANDN U58252 ( .A(n48785), .B(n48786), .Z(n48784) );
  NANDN U58253 ( .A(n48787), .B(n48788), .Z(n48786) );
  NANDN U58254 ( .A(n48788), .B(n48787), .Z(n48783) );
  IV U58255 ( .A(n48789), .Z(n48787) );
  XOR U58256 ( .A(n48764), .B(n48790), .Z(N61048) );
  XNOR U58257 ( .A(n48767), .B(n48766), .Z(n48790) );
  XNOR U58258 ( .A(n48778), .B(n48791), .Z(n48766) );
  XNOR U58259 ( .A(n48782), .B(n48780), .Z(n48791) );
  XOR U58260 ( .A(n48788), .B(n48792), .Z(n48780) );
  XNOR U58261 ( .A(n48785), .B(n48789), .Z(n48792) );
  AND U58262 ( .A(n48793), .B(n48794), .Z(n48789) );
  NAND U58263 ( .A(n48795), .B(n48796), .Z(n48794) );
  NAND U58264 ( .A(n48797), .B(n48798), .Z(n48793) );
  AND U58265 ( .A(n48799), .B(n48800), .Z(n48785) );
  NAND U58266 ( .A(n48801), .B(n48802), .Z(n48800) );
  NAND U58267 ( .A(n48803), .B(n48804), .Z(n48799) );
  NANDN U58268 ( .A(n48805), .B(n48806), .Z(n48788) );
  ANDN U58269 ( .B(n48807), .A(n48808), .Z(n48782) );
  XNOR U58270 ( .A(n48773), .B(n48809), .Z(n48778) );
  XNOR U58271 ( .A(n48771), .B(n48775), .Z(n48809) );
  AND U58272 ( .A(n48810), .B(n48811), .Z(n48775) );
  NAND U58273 ( .A(n48812), .B(n48813), .Z(n48811) );
  NAND U58274 ( .A(n48814), .B(n48815), .Z(n48810) );
  AND U58275 ( .A(n48816), .B(n48817), .Z(n48771) );
  NAND U58276 ( .A(n48818), .B(n48819), .Z(n48817) );
  NAND U58277 ( .A(n48820), .B(n48821), .Z(n48816) );
  AND U58278 ( .A(n48822), .B(n48823), .Z(n48773) );
  NAND U58279 ( .A(n48824), .B(n48825), .Z(n48767) );
  XNOR U58280 ( .A(n48750), .B(n48826), .Z(n48764) );
  XNOR U58281 ( .A(n48754), .B(n48752), .Z(n48826) );
  XOR U58282 ( .A(n48760), .B(n48827), .Z(n48752) );
  XNOR U58283 ( .A(n48757), .B(n48761), .Z(n48827) );
  AND U58284 ( .A(n48828), .B(n48829), .Z(n48761) );
  NAND U58285 ( .A(n48830), .B(n48831), .Z(n48829) );
  NAND U58286 ( .A(n48832), .B(n48833), .Z(n48828) );
  AND U58287 ( .A(n48834), .B(n48835), .Z(n48757) );
  NAND U58288 ( .A(n48836), .B(n48837), .Z(n48835) );
  NAND U58289 ( .A(n48838), .B(n48839), .Z(n48834) );
  NANDN U58290 ( .A(n48840), .B(n48841), .Z(n48760) );
  ANDN U58291 ( .B(n48842), .A(n48843), .Z(n48754) );
  XNOR U58292 ( .A(n48745), .B(n48844), .Z(n48750) );
  XNOR U58293 ( .A(n48743), .B(n48747), .Z(n48844) );
  AND U58294 ( .A(n48845), .B(n48846), .Z(n48747) );
  NAND U58295 ( .A(n48847), .B(n48848), .Z(n48846) );
  NAND U58296 ( .A(n48849), .B(n48850), .Z(n48845) );
  AND U58297 ( .A(n48851), .B(n48852), .Z(n48743) );
  NAND U58298 ( .A(n48853), .B(n48854), .Z(n48852) );
  NAND U58299 ( .A(n48855), .B(n48856), .Z(n48851) );
  AND U58300 ( .A(n48857), .B(n48858), .Z(n48745) );
  XOR U58301 ( .A(n48825), .B(n48824), .Z(N61047) );
  XNOR U58302 ( .A(n48842), .B(n48843), .Z(n48824) );
  XNOR U58303 ( .A(n48857), .B(n48858), .Z(n48843) );
  XOR U58304 ( .A(n48854), .B(n48853), .Z(n48858) );
  XOR U58305 ( .A(y[852]), .B(x[852]), .Z(n48853) );
  XOR U58306 ( .A(n48856), .B(n48855), .Z(n48854) );
  XOR U58307 ( .A(y[854]), .B(x[854]), .Z(n48855) );
  XOR U58308 ( .A(y[853]), .B(x[853]), .Z(n48856) );
  XOR U58309 ( .A(n48848), .B(n48847), .Z(n48857) );
  XOR U58310 ( .A(n48850), .B(n48849), .Z(n48847) );
  XOR U58311 ( .A(y[851]), .B(x[851]), .Z(n48849) );
  XOR U58312 ( .A(y[850]), .B(x[850]), .Z(n48850) );
  XOR U58313 ( .A(y[849]), .B(x[849]), .Z(n48848) );
  XNOR U58314 ( .A(n48841), .B(n48840), .Z(n48842) );
  XNOR U58315 ( .A(n48837), .B(n48836), .Z(n48840) );
  XOR U58316 ( .A(n48839), .B(n48838), .Z(n48836) );
  XOR U58317 ( .A(y[848]), .B(x[848]), .Z(n48838) );
  XOR U58318 ( .A(y[847]), .B(x[847]), .Z(n48839) );
  XOR U58319 ( .A(y[846]), .B(x[846]), .Z(n48837) );
  XOR U58320 ( .A(n48831), .B(n48830), .Z(n48841) );
  XOR U58321 ( .A(n48833), .B(n48832), .Z(n48830) );
  XOR U58322 ( .A(y[845]), .B(x[845]), .Z(n48832) );
  XOR U58323 ( .A(y[844]), .B(x[844]), .Z(n48833) );
  XOR U58324 ( .A(y[843]), .B(x[843]), .Z(n48831) );
  XNOR U58325 ( .A(n48807), .B(n48808), .Z(n48825) );
  XNOR U58326 ( .A(n48822), .B(n48823), .Z(n48808) );
  XOR U58327 ( .A(n48819), .B(n48818), .Z(n48823) );
  XOR U58328 ( .A(y[840]), .B(x[840]), .Z(n48818) );
  XOR U58329 ( .A(n48821), .B(n48820), .Z(n48819) );
  XOR U58330 ( .A(y[842]), .B(x[842]), .Z(n48820) );
  XOR U58331 ( .A(y[841]), .B(x[841]), .Z(n48821) );
  XOR U58332 ( .A(n48813), .B(n48812), .Z(n48822) );
  XOR U58333 ( .A(n48815), .B(n48814), .Z(n48812) );
  XOR U58334 ( .A(y[839]), .B(x[839]), .Z(n48814) );
  XOR U58335 ( .A(y[838]), .B(x[838]), .Z(n48815) );
  XOR U58336 ( .A(y[837]), .B(x[837]), .Z(n48813) );
  XNOR U58337 ( .A(n48806), .B(n48805), .Z(n48807) );
  XNOR U58338 ( .A(n48802), .B(n48801), .Z(n48805) );
  XOR U58339 ( .A(n48804), .B(n48803), .Z(n48801) );
  XOR U58340 ( .A(y[836]), .B(x[836]), .Z(n48803) );
  XOR U58341 ( .A(y[835]), .B(x[835]), .Z(n48804) );
  XOR U58342 ( .A(y[834]), .B(x[834]), .Z(n48802) );
  XOR U58343 ( .A(n48796), .B(n48795), .Z(n48806) );
  XOR U58344 ( .A(n48798), .B(n48797), .Z(n48795) );
  XOR U58345 ( .A(y[833]), .B(x[833]), .Z(n48797) );
  XOR U58346 ( .A(y[832]), .B(x[832]), .Z(n48798) );
  XOR U58347 ( .A(y[831]), .B(x[831]), .Z(n48796) );
  NAND U58348 ( .A(n48859), .B(n48860), .Z(N61038) );
  NAND U58349 ( .A(n48861), .B(n48862), .Z(n48860) );
  NANDN U58350 ( .A(n48863), .B(n48864), .Z(n48862) );
  NANDN U58351 ( .A(n48864), .B(n48863), .Z(n48859) );
  XOR U58352 ( .A(n48863), .B(n48865), .Z(N61037) );
  XNOR U58353 ( .A(n48861), .B(n48864), .Z(n48865) );
  NAND U58354 ( .A(n48866), .B(n48867), .Z(n48864) );
  NAND U58355 ( .A(n48868), .B(n48869), .Z(n48867) );
  NANDN U58356 ( .A(n48870), .B(n48871), .Z(n48869) );
  NANDN U58357 ( .A(n48871), .B(n48870), .Z(n48866) );
  AND U58358 ( .A(n48872), .B(n48873), .Z(n48861) );
  NAND U58359 ( .A(n48874), .B(n48875), .Z(n48873) );
  NANDN U58360 ( .A(n48876), .B(n48877), .Z(n48875) );
  NANDN U58361 ( .A(n48877), .B(n48876), .Z(n48872) );
  IV U58362 ( .A(n48878), .Z(n48877) );
  AND U58363 ( .A(n48879), .B(n48880), .Z(n48863) );
  NAND U58364 ( .A(n48881), .B(n48882), .Z(n48880) );
  NANDN U58365 ( .A(n48883), .B(n48884), .Z(n48882) );
  NANDN U58366 ( .A(n48884), .B(n48883), .Z(n48879) );
  XOR U58367 ( .A(n48876), .B(n48885), .Z(N61036) );
  XNOR U58368 ( .A(n48874), .B(n48878), .Z(n48885) );
  XOR U58369 ( .A(n48871), .B(n48886), .Z(n48878) );
  XNOR U58370 ( .A(n48868), .B(n48870), .Z(n48886) );
  AND U58371 ( .A(n48887), .B(n48888), .Z(n48870) );
  NANDN U58372 ( .A(n48889), .B(n48890), .Z(n48888) );
  OR U58373 ( .A(n48891), .B(n48892), .Z(n48890) );
  IV U58374 ( .A(n48893), .Z(n48892) );
  NANDN U58375 ( .A(n48893), .B(n48891), .Z(n48887) );
  AND U58376 ( .A(n48894), .B(n48895), .Z(n48868) );
  NAND U58377 ( .A(n48896), .B(n48897), .Z(n48895) );
  NANDN U58378 ( .A(n48898), .B(n48899), .Z(n48897) );
  NANDN U58379 ( .A(n48899), .B(n48898), .Z(n48894) );
  IV U58380 ( .A(n48900), .Z(n48899) );
  NAND U58381 ( .A(n48901), .B(n48902), .Z(n48871) );
  NANDN U58382 ( .A(n48903), .B(n48904), .Z(n48902) );
  NANDN U58383 ( .A(n48905), .B(n48906), .Z(n48904) );
  NANDN U58384 ( .A(n48906), .B(n48905), .Z(n48901) );
  IV U58385 ( .A(n48907), .Z(n48905) );
  AND U58386 ( .A(n48908), .B(n48909), .Z(n48874) );
  NAND U58387 ( .A(n48910), .B(n48911), .Z(n48909) );
  NANDN U58388 ( .A(n48912), .B(n48913), .Z(n48911) );
  NANDN U58389 ( .A(n48913), .B(n48912), .Z(n48908) );
  XOR U58390 ( .A(n48884), .B(n48914), .Z(n48876) );
  XNOR U58391 ( .A(n48881), .B(n48883), .Z(n48914) );
  AND U58392 ( .A(n48915), .B(n48916), .Z(n48883) );
  NANDN U58393 ( .A(n48917), .B(n48918), .Z(n48916) );
  OR U58394 ( .A(n48919), .B(n48920), .Z(n48918) );
  IV U58395 ( .A(n48921), .Z(n48920) );
  NANDN U58396 ( .A(n48921), .B(n48919), .Z(n48915) );
  AND U58397 ( .A(n48922), .B(n48923), .Z(n48881) );
  NAND U58398 ( .A(n48924), .B(n48925), .Z(n48923) );
  NANDN U58399 ( .A(n48926), .B(n48927), .Z(n48925) );
  NANDN U58400 ( .A(n48927), .B(n48926), .Z(n48922) );
  IV U58401 ( .A(n48928), .Z(n48927) );
  NAND U58402 ( .A(n48929), .B(n48930), .Z(n48884) );
  NANDN U58403 ( .A(n48931), .B(n48932), .Z(n48930) );
  NANDN U58404 ( .A(n48933), .B(n48934), .Z(n48932) );
  NANDN U58405 ( .A(n48934), .B(n48933), .Z(n48929) );
  IV U58406 ( .A(n48935), .Z(n48933) );
  XOR U58407 ( .A(n48910), .B(n48936), .Z(N61035) );
  XNOR U58408 ( .A(n48913), .B(n48912), .Z(n48936) );
  XNOR U58409 ( .A(n48924), .B(n48937), .Z(n48912) );
  XNOR U58410 ( .A(n48928), .B(n48926), .Z(n48937) );
  XOR U58411 ( .A(n48934), .B(n48938), .Z(n48926) );
  XNOR U58412 ( .A(n48931), .B(n48935), .Z(n48938) );
  AND U58413 ( .A(n48939), .B(n48940), .Z(n48935) );
  NAND U58414 ( .A(n48941), .B(n48942), .Z(n48940) );
  NAND U58415 ( .A(n48943), .B(n48944), .Z(n48939) );
  AND U58416 ( .A(n48945), .B(n48946), .Z(n48931) );
  NAND U58417 ( .A(n48947), .B(n48948), .Z(n48946) );
  NAND U58418 ( .A(n48949), .B(n48950), .Z(n48945) );
  NANDN U58419 ( .A(n48951), .B(n48952), .Z(n48934) );
  ANDN U58420 ( .B(n48953), .A(n48954), .Z(n48928) );
  XNOR U58421 ( .A(n48919), .B(n48955), .Z(n48924) );
  XNOR U58422 ( .A(n48917), .B(n48921), .Z(n48955) );
  AND U58423 ( .A(n48956), .B(n48957), .Z(n48921) );
  NAND U58424 ( .A(n48958), .B(n48959), .Z(n48957) );
  NAND U58425 ( .A(n48960), .B(n48961), .Z(n48956) );
  AND U58426 ( .A(n48962), .B(n48963), .Z(n48917) );
  NAND U58427 ( .A(n48964), .B(n48965), .Z(n48963) );
  NAND U58428 ( .A(n48966), .B(n48967), .Z(n48962) );
  AND U58429 ( .A(n48968), .B(n48969), .Z(n48919) );
  NAND U58430 ( .A(n48970), .B(n48971), .Z(n48913) );
  XNOR U58431 ( .A(n48896), .B(n48972), .Z(n48910) );
  XNOR U58432 ( .A(n48900), .B(n48898), .Z(n48972) );
  XOR U58433 ( .A(n48906), .B(n48973), .Z(n48898) );
  XNOR U58434 ( .A(n48903), .B(n48907), .Z(n48973) );
  AND U58435 ( .A(n48974), .B(n48975), .Z(n48907) );
  NAND U58436 ( .A(n48976), .B(n48977), .Z(n48975) );
  NAND U58437 ( .A(n48978), .B(n48979), .Z(n48974) );
  AND U58438 ( .A(n48980), .B(n48981), .Z(n48903) );
  NAND U58439 ( .A(n48982), .B(n48983), .Z(n48981) );
  NAND U58440 ( .A(n48984), .B(n48985), .Z(n48980) );
  NANDN U58441 ( .A(n48986), .B(n48987), .Z(n48906) );
  ANDN U58442 ( .B(n48988), .A(n48989), .Z(n48900) );
  XNOR U58443 ( .A(n48891), .B(n48990), .Z(n48896) );
  XNOR U58444 ( .A(n48889), .B(n48893), .Z(n48990) );
  AND U58445 ( .A(n48991), .B(n48992), .Z(n48893) );
  NAND U58446 ( .A(n48993), .B(n48994), .Z(n48992) );
  NAND U58447 ( .A(n48995), .B(n48996), .Z(n48991) );
  AND U58448 ( .A(n48997), .B(n48998), .Z(n48889) );
  NAND U58449 ( .A(n48999), .B(n49000), .Z(n48998) );
  NAND U58450 ( .A(n49001), .B(n49002), .Z(n48997) );
  AND U58451 ( .A(n49003), .B(n49004), .Z(n48891) );
  XOR U58452 ( .A(n48971), .B(n48970), .Z(N61034) );
  XNOR U58453 ( .A(n48988), .B(n48989), .Z(n48970) );
  XNOR U58454 ( .A(n49003), .B(n49004), .Z(n48989) );
  XOR U58455 ( .A(n49000), .B(n48999), .Z(n49004) );
  XOR U58456 ( .A(y[828]), .B(x[828]), .Z(n48999) );
  XOR U58457 ( .A(n49002), .B(n49001), .Z(n49000) );
  XOR U58458 ( .A(y[830]), .B(x[830]), .Z(n49001) );
  XOR U58459 ( .A(y[829]), .B(x[829]), .Z(n49002) );
  XOR U58460 ( .A(n48994), .B(n48993), .Z(n49003) );
  XOR U58461 ( .A(n48996), .B(n48995), .Z(n48993) );
  XOR U58462 ( .A(y[827]), .B(x[827]), .Z(n48995) );
  XOR U58463 ( .A(y[826]), .B(x[826]), .Z(n48996) );
  XOR U58464 ( .A(y[825]), .B(x[825]), .Z(n48994) );
  XNOR U58465 ( .A(n48987), .B(n48986), .Z(n48988) );
  XNOR U58466 ( .A(n48983), .B(n48982), .Z(n48986) );
  XOR U58467 ( .A(n48985), .B(n48984), .Z(n48982) );
  XOR U58468 ( .A(y[824]), .B(x[824]), .Z(n48984) );
  XOR U58469 ( .A(y[823]), .B(x[823]), .Z(n48985) );
  XOR U58470 ( .A(y[822]), .B(x[822]), .Z(n48983) );
  XOR U58471 ( .A(n48977), .B(n48976), .Z(n48987) );
  XOR U58472 ( .A(n48979), .B(n48978), .Z(n48976) );
  XOR U58473 ( .A(y[821]), .B(x[821]), .Z(n48978) );
  XOR U58474 ( .A(y[820]), .B(x[820]), .Z(n48979) );
  XOR U58475 ( .A(y[819]), .B(x[819]), .Z(n48977) );
  XNOR U58476 ( .A(n48953), .B(n48954), .Z(n48971) );
  XNOR U58477 ( .A(n48968), .B(n48969), .Z(n48954) );
  XOR U58478 ( .A(n48965), .B(n48964), .Z(n48969) );
  XOR U58479 ( .A(y[816]), .B(x[816]), .Z(n48964) );
  XOR U58480 ( .A(n48967), .B(n48966), .Z(n48965) );
  XOR U58481 ( .A(y[818]), .B(x[818]), .Z(n48966) );
  XOR U58482 ( .A(y[817]), .B(x[817]), .Z(n48967) );
  XOR U58483 ( .A(n48959), .B(n48958), .Z(n48968) );
  XOR U58484 ( .A(n48961), .B(n48960), .Z(n48958) );
  XOR U58485 ( .A(y[815]), .B(x[815]), .Z(n48960) );
  XOR U58486 ( .A(y[814]), .B(x[814]), .Z(n48961) );
  XOR U58487 ( .A(y[813]), .B(x[813]), .Z(n48959) );
  XNOR U58488 ( .A(n48952), .B(n48951), .Z(n48953) );
  XNOR U58489 ( .A(n48948), .B(n48947), .Z(n48951) );
  XOR U58490 ( .A(n48950), .B(n48949), .Z(n48947) );
  XOR U58491 ( .A(y[812]), .B(x[812]), .Z(n48949) );
  XOR U58492 ( .A(y[811]), .B(x[811]), .Z(n48950) );
  XOR U58493 ( .A(y[810]), .B(x[810]), .Z(n48948) );
  XOR U58494 ( .A(n48942), .B(n48941), .Z(n48952) );
  XOR U58495 ( .A(n48944), .B(n48943), .Z(n48941) );
  XOR U58496 ( .A(y[809]), .B(x[809]), .Z(n48943) );
  XOR U58497 ( .A(y[808]), .B(x[808]), .Z(n48944) );
  XOR U58498 ( .A(y[807]), .B(x[807]), .Z(n48942) );
  NAND U58499 ( .A(n49005), .B(n49006), .Z(N61025) );
  NAND U58500 ( .A(n49007), .B(n49008), .Z(n49006) );
  NANDN U58501 ( .A(n49009), .B(n49010), .Z(n49008) );
  NANDN U58502 ( .A(n49010), .B(n49009), .Z(n49005) );
  XOR U58503 ( .A(n49009), .B(n49011), .Z(N61024) );
  XNOR U58504 ( .A(n49007), .B(n49010), .Z(n49011) );
  NAND U58505 ( .A(n49012), .B(n49013), .Z(n49010) );
  NAND U58506 ( .A(n49014), .B(n49015), .Z(n49013) );
  NANDN U58507 ( .A(n49016), .B(n49017), .Z(n49015) );
  NANDN U58508 ( .A(n49017), .B(n49016), .Z(n49012) );
  AND U58509 ( .A(n49018), .B(n49019), .Z(n49007) );
  NAND U58510 ( .A(n49020), .B(n49021), .Z(n49019) );
  NANDN U58511 ( .A(n49022), .B(n49023), .Z(n49021) );
  NANDN U58512 ( .A(n49023), .B(n49022), .Z(n49018) );
  IV U58513 ( .A(n49024), .Z(n49023) );
  AND U58514 ( .A(n49025), .B(n49026), .Z(n49009) );
  NAND U58515 ( .A(n49027), .B(n49028), .Z(n49026) );
  NANDN U58516 ( .A(n49029), .B(n49030), .Z(n49028) );
  NANDN U58517 ( .A(n49030), .B(n49029), .Z(n49025) );
  XOR U58518 ( .A(n49022), .B(n49031), .Z(N61023) );
  XNOR U58519 ( .A(n49020), .B(n49024), .Z(n49031) );
  XOR U58520 ( .A(n49017), .B(n49032), .Z(n49024) );
  XNOR U58521 ( .A(n49014), .B(n49016), .Z(n49032) );
  AND U58522 ( .A(n49033), .B(n49034), .Z(n49016) );
  NANDN U58523 ( .A(n49035), .B(n49036), .Z(n49034) );
  OR U58524 ( .A(n49037), .B(n49038), .Z(n49036) );
  IV U58525 ( .A(n49039), .Z(n49038) );
  NANDN U58526 ( .A(n49039), .B(n49037), .Z(n49033) );
  AND U58527 ( .A(n49040), .B(n49041), .Z(n49014) );
  NAND U58528 ( .A(n49042), .B(n49043), .Z(n49041) );
  NANDN U58529 ( .A(n49044), .B(n49045), .Z(n49043) );
  NANDN U58530 ( .A(n49045), .B(n49044), .Z(n49040) );
  IV U58531 ( .A(n49046), .Z(n49045) );
  NAND U58532 ( .A(n49047), .B(n49048), .Z(n49017) );
  NANDN U58533 ( .A(n49049), .B(n49050), .Z(n49048) );
  NANDN U58534 ( .A(n49051), .B(n49052), .Z(n49050) );
  NANDN U58535 ( .A(n49052), .B(n49051), .Z(n49047) );
  IV U58536 ( .A(n49053), .Z(n49051) );
  AND U58537 ( .A(n49054), .B(n49055), .Z(n49020) );
  NAND U58538 ( .A(n49056), .B(n49057), .Z(n49055) );
  NANDN U58539 ( .A(n49058), .B(n49059), .Z(n49057) );
  NANDN U58540 ( .A(n49059), .B(n49058), .Z(n49054) );
  XOR U58541 ( .A(n49030), .B(n49060), .Z(n49022) );
  XNOR U58542 ( .A(n49027), .B(n49029), .Z(n49060) );
  AND U58543 ( .A(n49061), .B(n49062), .Z(n49029) );
  NANDN U58544 ( .A(n49063), .B(n49064), .Z(n49062) );
  OR U58545 ( .A(n49065), .B(n49066), .Z(n49064) );
  IV U58546 ( .A(n49067), .Z(n49066) );
  NANDN U58547 ( .A(n49067), .B(n49065), .Z(n49061) );
  AND U58548 ( .A(n49068), .B(n49069), .Z(n49027) );
  NAND U58549 ( .A(n49070), .B(n49071), .Z(n49069) );
  NANDN U58550 ( .A(n49072), .B(n49073), .Z(n49071) );
  NANDN U58551 ( .A(n49073), .B(n49072), .Z(n49068) );
  IV U58552 ( .A(n49074), .Z(n49073) );
  NAND U58553 ( .A(n49075), .B(n49076), .Z(n49030) );
  NANDN U58554 ( .A(n49077), .B(n49078), .Z(n49076) );
  NANDN U58555 ( .A(n49079), .B(n49080), .Z(n49078) );
  NANDN U58556 ( .A(n49080), .B(n49079), .Z(n49075) );
  IV U58557 ( .A(n49081), .Z(n49079) );
  XOR U58558 ( .A(n49056), .B(n49082), .Z(N61022) );
  XNOR U58559 ( .A(n49059), .B(n49058), .Z(n49082) );
  XNOR U58560 ( .A(n49070), .B(n49083), .Z(n49058) );
  XNOR U58561 ( .A(n49074), .B(n49072), .Z(n49083) );
  XOR U58562 ( .A(n49080), .B(n49084), .Z(n49072) );
  XNOR U58563 ( .A(n49077), .B(n49081), .Z(n49084) );
  AND U58564 ( .A(n49085), .B(n49086), .Z(n49081) );
  NAND U58565 ( .A(n49087), .B(n49088), .Z(n49086) );
  NAND U58566 ( .A(n49089), .B(n49090), .Z(n49085) );
  AND U58567 ( .A(n49091), .B(n49092), .Z(n49077) );
  NAND U58568 ( .A(n49093), .B(n49094), .Z(n49092) );
  NAND U58569 ( .A(n49095), .B(n49096), .Z(n49091) );
  NANDN U58570 ( .A(n49097), .B(n49098), .Z(n49080) );
  ANDN U58571 ( .B(n49099), .A(n49100), .Z(n49074) );
  XNOR U58572 ( .A(n49065), .B(n49101), .Z(n49070) );
  XNOR U58573 ( .A(n49063), .B(n49067), .Z(n49101) );
  AND U58574 ( .A(n49102), .B(n49103), .Z(n49067) );
  NAND U58575 ( .A(n49104), .B(n49105), .Z(n49103) );
  NAND U58576 ( .A(n49106), .B(n49107), .Z(n49102) );
  AND U58577 ( .A(n49108), .B(n49109), .Z(n49063) );
  NAND U58578 ( .A(n49110), .B(n49111), .Z(n49109) );
  NAND U58579 ( .A(n49112), .B(n49113), .Z(n49108) );
  AND U58580 ( .A(n49114), .B(n49115), .Z(n49065) );
  NAND U58581 ( .A(n49116), .B(n49117), .Z(n49059) );
  XNOR U58582 ( .A(n49042), .B(n49118), .Z(n49056) );
  XNOR U58583 ( .A(n49046), .B(n49044), .Z(n49118) );
  XOR U58584 ( .A(n49052), .B(n49119), .Z(n49044) );
  XNOR U58585 ( .A(n49049), .B(n49053), .Z(n49119) );
  AND U58586 ( .A(n49120), .B(n49121), .Z(n49053) );
  NAND U58587 ( .A(n49122), .B(n49123), .Z(n49121) );
  NAND U58588 ( .A(n49124), .B(n49125), .Z(n49120) );
  AND U58589 ( .A(n49126), .B(n49127), .Z(n49049) );
  NAND U58590 ( .A(n49128), .B(n49129), .Z(n49127) );
  NAND U58591 ( .A(n49130), .B(n49131), .Z(n49126) );
  NANDN U58592 ( .A(n49132), .B(n49133), .Z(n49052) );
  ANDN U58593 ( .B(n49134), .A(n49135), .Z(n49046) );
  XNOR U58594 ( .A(n49037), .B(n49136), .Z(n49042) );
  XNOR U58595 ( .A(n49035), .B(n49039), .Z(n49136) );
  AND U58596 ( .A(n49137), .B(n49138), .Z(n49039) );
  NAND U58597 ( .A(n49139), .B(n49140), .Z(n49138) );
  NAND U58598 ( .A(n49141), .B(n49142), .Z(n49137) );
  AND U58599 ( .A(n49143), .B(n49144), .Z(n49035) );
  NAND U58600 ( .A(n49145), .B(n49146), .Z(n49144) );
  NAND U58601 ( .A(n49147), .B(n49148), .Z(n49143) );
  AND U58602 ( .A(n49149), .B(n49150), .Z(n49037) );
  XOR U58603 ( .A(n49117), .B(n49116), .Z(N61021) );
  XNOR U58604 ( .A(n49134), .B(n49135), .Z(n49116) );
  XNOR U58605 ( .A(n49149), .B(n49150), .Z(n49135) );
  XOR U58606 ( .A(n49146), .B(n49145), .Z(n49150) );
  XOR U58607 ( .A(y[804]), .B(x[804]), .Z(n49145) );
  XOR U58608 ( .A(n49148), .B(n49147), .Z(n49146) );
  XOR U58609 ( .A(y[806]), .B(x[806]), .Z(n49147) );
  XOR U58610 ( .A(y[805]), .B(x[805]), .Z(n49148) );
  XOR U58611 ( .A(n49140), .B(n49139), .Z(n49149) );
  XOR U58612 ( .A(n49142), .B(n49141), .Z(n49139) );
  XOR U58613 ( .A(y[803]), .B(x[803]), .Z(n49141) );
  XOR U58614 ( .A(y[802]), .B(x[802]), .Z(n49142) );
  XOR U58615 ( .A(y[801]), .B(x[801]), .Z(n49140) );
  XNOR U58616 ( .A(n49133), .B(n49132), .Z(n49134) );
  XNOR U58617 ( .A(n49129), .B(n49128), .Z(n49132) );
  XOR U58618 ( .A(n49131), .B(n49130), .Z(n49128) );
  XOR U58619 ( .A(y[800]), .B(x[800]), .Z(n49130) );
  XOR U58620 ( .A(y[799]), .B(x[799]), .Z(n49131) );
  XOR U58621 ( .A(y[798]), .B(x[798]), .Z(n49129) );
  XOR U58622 ( .A(n49123), .B(n49122), .Z(n49133) );
  XOR U58623 ( .A(n49125), .B(n49124), .Z(n49122) );
  XOR U58624 ( .A(y[797]), .B(x[797]), .Z(n49124) );
  XOR U58625 ( .A(y[796]), .B(x[796]), .Z(n49125) );
  XOR U58626 ( .A(y[795]), .B(x[795]), .Z(n49123) );
  XNOR U58627 ( .A(n49099), .B(n49100), .Z(n49117) );
  XNOR U58628 ( .A(n49114), .B(n49115), .Z(n49100) );
  XOR U58629 ( .A(n49111), .B(n49110), .Z(n49115) );
  XOR U58630 ( .A(y[792]), .B(x[792]), .Z(n49110) );
  XOR U58631 ( .A(n49113), .B(n49112), .Z(n49111) );
  XOR U58632 ( .A(y[794]), .B(x[794]), .Z(n49112) );
  XOR U58633 ( .A(y[793]), .B(x[793]), .Z(n49113) );
  XOR U58634 ( .A(n49105), .B(n49104), .Z(n49114) );
  XOR U58635 ( .A(n49107), .B(n49106), .Z(n49104) );
  XOR U58636 ( .A(y[791]), .B(x[791]), .Z(n49106) );
  XOR U58637 ( .A(y[790]), .B(x[790]), .Z(n49107) );
  XOR U58638 ( .A(y[789]), .B(x[789]), .Z(n49105) );
  XNOR U58639 ( .A(n49098), .B(n49097), .Z(n49099) );
  XNOR U58640 ( .A(n49094), .B(n49093), .Z(n49097) );
  XOR U58641 ( .A(n49096), .B(n49095), .Z(n49093) );
  XOR U58642 ( .A(y[788]), .B(x[788]), .Z(n49095) );
  XOR U58643 ( .A(y[787]), .B(x[787]), .Z(n49096) );
  XOR U58644 ( .A(y[786]), .B(x[786]), .Z(n49094) );
  XOR U58645 ( .A(n49088), .B(n49087), .Z(n49098) );
  XOR U58646 ( .A(n49090), .B(n49089), .Z(n49087) );
  XOR U58647 ( .A(y[785]), .B(x[785]), .Z(n49089) );
  XOR U58648 ( .A(y[784]), .B(x[784]), .Z(n49090) );
  XOR U58649 ( .A(y[783]), .B(x[783]), .Z(n49088) );
  NAND U58650 ( .A(n49151), .B(n49152), .Z(N61012) );
  NAND U58651 ( .A(n49153), .B(n49154), .Z(n49152) );
  NANDN U58652 ( .A(n49155), .B(n49156), .Z(n49154) );
  NANDN U58653 ( .A(n49156), .B(n49155), .Z(n49151) );
  XOR U58654 ( .A(n49155), .B(n49157), .Z(N61011) );
  XNOR U58655 ( .A(n49153), .B(n49156), .Z(n49157) );
  NAND U58656 ( .A(n49158), .B(n49159), .Z(n49156) );
  NAND U58657 ( .A(n49160), .B(n49161), .Z(n49159) );
  NANDN U58658 ( .A(n49162), .B(n49163), .Z(n49161) );
  NANDN U58659 ( .A(n49163), .B(n49162), .Z(n49158) );
  AND U58660 ( .A(n49164), .B(n49165), .Z(n49153) );
  NAND U58661 ( .A(n49166), .B(n49167), .Z(n49165) );
  NANDN U58662 ( .A(n49168), .B(n49169), .Z(n49167) );
  NANDN U58663 ( .A(n49169), .B(n49168), .Z(n49164) );
  IV U58664 ( .A(n49170), .Z(n49169) );
  AND U58665 ( .A(n49171), .B(n49172), .Z(n49155) );
  NAND U58666 ( .A(n49173), .B(n49174), .Z(n49172) );
  NANDN U58667 ( .A(n49175), .B(n49176), .Z(n49174) );
  NANDN U58668 ( .A(n49176), .B(n49175), .Z(n49171) );
  XOR U58669 ( .A(n49168), .B(n49177), .Z(N61010) );
  XNOR U58670 ( .A(n49166), .B(n49170), .Z(n49177) );
  XOR U58671 ( .A(n49163), .B(n49178), .Z(n49170) );
  XNOR U58672 ( .A(n49160), .B(n49162), .Z(n49178) );
  AND U58673 ( .A(n49179), .B(n49180), .Z(n49162) );
  NANDN U58674 ( .A(n49181), .B(n49182), .Z(n49180) );
  OR U58675 ( .A(n49183), .B(n49184), .Z(n49182) );
  IV U58676 ( .A(n49185), .Z(n49184) );
  NANDN U58677 ( .A(n49185), .B(n49183), .Z(n49179) );
  AND U58678 ( .A(n49186), .B(n49187), .Z(n49160) );
  NAND U58679 ( .A(n49188), .B(n49189), .Z(n49187) );
  NANDN U58680 ( .A(n49190), .B(n49191), .Z(n49189) );
  NANDN U58681 ( .A(n49191), .B(n49190), .Z(n49186) );
  IV U58682 ( .A(n49192), .Z(n49191) );
  NAND U58683 ( .A(n49193), .B(n49194), .Z(n49163) );
  NANDN U58684 ( .A(n49195), .B(n49196), .Z(n49194) );
  NANDN U58685 ( .A(n49197), .B(n49198), .Z(n49196) );
  NANDN U58686 ( .A(n49198), .B(n49197), .Z(n49193) );
  IV U58687 ( .A(n49199), .Z(n49197) );
  AND U58688 ( .A(n49200), .B(n49201), .Z(n49166) );
  NAND U58689 ( .A(n49202), .B(n49203), .Z(n49201) );
  NANDN U58690 ( .A(n49204), .B(n49205), .Z(n49203) );
  NANDN U58691 ( .A(n49205), .B(n49204), .Z(n49200) );
  XOR U58692 ( .A(n49176), .B(n49206), .Z(n49168) );
  XNOR U58693 ( .A(n49173), .B(n49175), .Z(n49206) );
  AND U58694 ( .A(n49207), .B(n49208), .Z(n49175) );
  NANDN U58695 ( .A(n49209), .B(n49210), .Z(n49208) );
  OR U58696 ( .A(n49211), .B(n49212), .Z(n49210) );
  IV U58697 ( .A(n49213), .Z(n49212) );
  NANDN U58698 ( .A(n49213), .B(n49211), .Z(n49207) );
  AND U58699 ( .A(n49214), .B(n49215), .Z(n49173) );
  NAND U58700 ( .A(n49216), .B(n49217), .Z(n49215) );
  NANDN U58701 ( .A(n49218), .B(n49219), .Z(n49217) );
  NANDN U58702 ( .A(n49219), .B(n49218), .Z(n49214) );
  IV U58703 ( .A(n49220), .Z(n49219) );
  NAND U58704 ( .A(n49221), .B(n49222), .Z(n49176) );
  NANDN U58705 ( .A(n49223), .B(n49224), .Z(n49222) );
  NANDN U58706 ( .A(n49225), .B(n49226), .Z(n49224) );
  NANDN U58707 ( .A(n49226), .B(n49225), .Z(n49221) );
  IV U58708 ( .A(n49227), .Z(n49225) );
  XOR U58709 ( .A(n49202), .B(n49228), .Z(N61009) );
  XNOR U58710 ( .A(n49205), .B(n49204), .Z(n49228) );
  XNOR U58711 ( .A(n49216), .B(n49229), .Z(n49204) );
  XNOR U58712 ( .A(n49220), .B(n49218), .Z(n49229) );
  XOR U58713 ( .A(n49226), .B(n49230), .Z(n49218) );
  XNOR U58714 ( .A(n49223), .B(n49227), .Z(n49230) );
  AND U58715 ( .A(n49231), .B(n49232), .Z(n49227) );
  NAND U58716 ( .A(n49233), .B(n49234), .Z(n49232) );
  NAND U58717 ( .A(n49235), .B(n49236), .Z(n49231) );
  AND U58718 ( .A(n49237), .B(n49238), .Z(n49223) );
  NAND U58719 ( .A(n49239), .B(n49240), .Z(n49238) );
  NAND U58720 ( .A(n49241), .B(n49242), .Z(n49237) );
  NANDN U58721 ( .A(n49243), .B(n49244), .Z(n49226) );
  ANDN U58722 ( .B(n49245), .A(n49246), .Z(n49220) );
  XNOR U58723 ( .A(n49211), .B(n49247), .Z(n49216) );
  XNOR U58724 ( .A(n49209), .B(n49213), .Z(n49247) );
  AND U58725 ( .A(n49248), .B(n49249), .Z(n49213) );
  NAND U58726 ( .A(n49250), .B(n49251), .Z(n49249) );
  NAND U58727 ( .A(n49252), .B(n49253), .Z(n49248) );
  AND U58728 ( .A(n49254), .B(n49255), .Z(n49209) );
  NAND U58729 ( .A(n49256), .B(n49257), .Z(n49255) );
  NAND U58730 ( .A(n49258), .B(n49259), .Z(n49254) );
  AND U58731 ( .A(n49260), .B(n49261), .Z(n49211) );
  NAND U58732 ( .A(n49262), .B(n49263), .Z(n49205) );
  XNOR U58733 ( .A(n49188), .B(n49264), .Z(n49202) );
  XNOR U58734 ( .A(n49192), .B(n49190), .Z(n49264) );
  XOR U58735 ( .A(n49198), .B(n49265), .Z(n49190) );
  XNOR U58736 ( .A(n49195), .B(n49199), .Z(n49265) );
  AND U58737 ( .A(n49266), .B(n49267), .Z(n49199) );
  NAND U58738 ( .A(n49268), .B(n49269), .Z(n49267) );
  NAND U58739 ( .A(n49270), .B(n49271), .Z(n49266) );
  AND U58740 ( .A(n49272), .B(n49273), .Z(n49195) );
  NAND U58741 ( .A(n49274), .B(n49275), .Z(n49273) );
  NAND U58742 ( .A(n49276), .B(n49277), .Z(n49272) );
  NANDN U58743 ( .A(n49278), .B(n49279), .Z(n49198) );
  ANDN U58744 ( .B(n49280), .A(n49281), .Z(n49192) );
  XNOR U58745 ( .A(n49183), .B(n49282), .Z(n49188) );
  XNOR U58746 ( .A(n49181), .B(n49185), .Z(n49282) );
  AND U58747 ( .A(n49283), .B(n49284), .Z(n49185) );
  NAND U58748 ( .A(n49285), .B(n49286), .Z(n49284) );
  NAND U58749 ( .A(n49287), .B(n49288), .Z(n49283) );
  AND U58750 ( .A(n49289), .B(n49290), .Z(n49181) );
  NAND U58751 ( .A(n49291), .B(n49292), .Z(n49290) );
  NAND U58752 ( .A(n49293), .B(n49294), .Z(n49289) );
  AND U58753 ( .A(n49295), .B(n49296), .Z(n49183) );
  XOR U58754 ( .A(n49263), .B(n49262), .Z(N61008) );
  XNOR U58755 ( .A(n49280), .B(n49281), .Z(n49262) );
  XNOR U58756 ( .A(n49295), .B(n49296), .Z(n49281) );
  XOR U58757 ( .A(n49292), .B(n49291), .Z(n49296) );
  XOR U58758 ( .A(y[780]), .B(x[780]), .Z(n49291) );
  XOR U58759 ( .A(n49294), .B(n49293), .Z(n49292) );
  XOR U58760 ( .A(y[782]), .B(x[782]), .Z(n49293) );
  XOR U58761 ( .A(y[781]), .B(x[781]), .Z(n49294) );
  XOR U58762 ( .A(n49286), .B(n49285), .Z(n49295) );
  XOR U58763 ( .A(n49288), .B(n49287), .Z(n49285) );
  XOR U58764 ( .A(y[779]), .B(x[779]), .Z(n49287) );
  XOR U58765 ( .A(y[778]), .B(x[778]), .Z(n49288) );
  XOR U58766 ( .A(y[777]), .B(x[777]), .Z(n49286) );
  XNOR U58767 ( .A(n49279), .B(n49278), .Z(n49280) );
  XNOR U58768 ( .A(n49275), .B(n49274), .Z(n49278) );
  XOR U58769 ( .A(n49277), .B(n49276), .Z(n49274) );
  XOR U58770 ( .A(y[776]), .B(x[776]), .Z(n49276) );
  XOR U58771 ( .A(y[775]), .B(x[775]), .Z(n49277) );
  XOR U58772 ( .A(y[774]), .B(x[774]), .Z(n49275) );
  XOR U58773 ( .A(n49269), .B(n49268), .Z(n49279) );
  XOR U58774 ( .A(n49271), .B(n49270), .Z(n49268) );
  XOR U58775 ( .A(y[773]), .B(x[773]), .Z(n49270) );
  XOR U58776 ( .A(y[772]), .B(x[772]), .Z(n49271) );
  XOR U58777 ( .A(y[771]), .B(x[771]), .Z(n49269) );
  XNOR U58778 ( .A(n49245), .B(n49246), .Z(n49263) );
  XNOR U58779 ( .A(n49260), .B(n49261), .Z(n49246) );
  XOR U58780 ( .A(n49257), .B(n49256), .Z(n49261) );
  XOR U58781 ( .A(y[768]), .B(x[768]), .Z(n49256) );
  XOR U58782 ( .A(n49259), .B(n49258), .Z(n49257) );
  XOR U58783 ( .A(y[770]), .B(x[770]), .Z(n49258) );
  XOR U58784 ( .A(y[769]), .B(x[769]), .Z(n49259) );
  XOR U58785 ( .A(n49251), .B(n49250), .Z(n49260) );
  XOR U58786 ( .A(n49253), .B(n49252), .Z(n49250) );
  XOR U58787 ( .A(y[767]), .B(x[767]), .Z(n49252) );
  XOR U58788 ( .A(y[766]), .B(x[766]), .Z(n49253) );
  XOR U58789 ( .A(y[765]), .B(x[765]), .Z(n49251) );
  XNOR U58790 ( .A(n49244), .B(n49243), .Z(n49245) );
  XNOR U58791 ( .A(n49240), .B(n49239), .Z(n49243) );
  XOR U58792 ( .A(n49242), .B(n49241), .Z(n49239) );
  XOR U58793 ( .A(y[764]), .B(x[764]), .Z(n49241) );
  XOR U58794 ( .A(y[763]), .B(x[763]), .Z(n49242) );
  XOR U58795 ( .A(y[762]), .B(x[762]), .Z(n49240) );
  XOR U58796 ( .A(n49234), .B(n49233), .Z(n49244) );
  XOR U58797 ( .A(n49236), .B(n49235), .Z(n49233) );
  XOR U58798 ( .A(y[761]), .B(x[761]), .Z(n49235) );
  XOR U58799 ( .A(y[760]), .B(x[760]), .Z(n49236) );
  XOR U58800 ( .A(y[759]), .B(x[759]), .Z(n49234) );
  NAND U58801 ( .A(n49297), .B(n49298), .Z(N60999) );
  NAND U58802 ( .A(n49299), .B(n49300), .Z(n49298) );
  NANDN U58803 ( .A(n49301), .B(n49302), .Z(n49300) );
  NANDN U58804 ( .A(n49302), .B(n49301), .Z(n49297) );
  XOR U58805 ( .A(n49301), .B(n49303), .Z(N60998) );
  XNOR U58806 ( .A(n49299), .B(n49302), .Z(n49303) );
  NAND U58807 ( .A(n49304), .B(n49305), .Z(n49302) );
  NAND U58808 ( .A(n49306), .B(n49307), .Z(n49305) );
  NANDN U58809 ( .A(n49308), .B(n49309), .Z(n49307) );
  NANDN U58810 ( .A(n49309), .B(n49308), .Z(n49304) );
  AND U58811 ( .A(n49310), .B(n49311), .Z(n49299) );
  NAND U58812 ( .A(n49312), .B(n49313), .Z(n49311) );
  NANDN U58813 ( .A(n49314), .B(n49315), .Z(n49313) );
  NANDN U58814 ( .A(n49315), .B(n49314), .Z(n49310) );
  IV U58815 ( .A(n49316), .Z(n49315) );
  AND U58816 ( .A(n49317), .B(n49318), .Z(n49301) );
  NAND U58817 ( .A(n49319), .B(n49320), .Z(n49318) );
  NANDN U58818 ( .A(n49321), .B(n49322), .Z(n49320) );
  NANDN U58819 ( .A(n49322), .B(n49321), .Z(n49317) );
  XOR U58820 ( .A(n49314), .B(n49323), .Z(N60997) );
  XNOR U58821 ( .A(n49312), .B(n49316), .Z(n49323) );
  XOR U58822 ( .A(n49309), .B(n49324), .Z(n49316) );
  XNOR U58823 ( .A(n49306), .B(n49308), .Z(n49324) );
  AND U58824 ( .A(n49325), .B(n49326), .Z(n49308) );
  NANDN U58825 ( .A(n49327), .B(n49328), .Z(n49326) );
  OR U58826 ( .A(n49329), .B(n49330), .Z(n49328) );
  IV U58827 ( .A(n49331), .Z(n49330) );
  NANDN U58828 ( .A(n49331), .B(n49329), .Z(n49325) );
  AND U58829 ( .A(n49332), .B(n49333), .Z(n49306) );
  NAND U58830 ( .A(n49334), .B(n49335), .Z(n49333) );
  NANDN U58831 ( .A(n49336), .B(n49337), .Z(n49335) );
  NANDN U58832 ( .A(n49337), .B(n49336), .Z(n49332) );
  IV U58833 ( .A(n49338), .Z(n49337) );
  NAND U58834 ( .A(n49339), .B(n49340), .Z(n49309) );
  NANDN U58835 ( .A(n49341), .B(n49342), .Z(n49340) );
  NANDN U58836 ( .A(n49343), .B(n49344), .Z(n49342) );
  NANDN U58837 ( .A(n49344), .B(n49343), .Z(n49339) );
  IV U58838 ( .A(n49345), .Z(n49343) );
  AND U58839 ( .A(n49346), .B(n49347), .Z(n49312) );
  NAND U58840 ( .A(n49348), .B(n49349), .Z(n49347) );
  NANDN U58841 ( .A(n49350), .B(n49351), .Z(n49349) );
  NANDN U58842 ( .A(n49351), .B(n49350), .Z(n49346) );
  XOR U58843 ( .A(n49322), .B(n49352), .Z(n49314) );
  XNOR U58844 ( .A(n49319), .B(n49321), .Z(n49352) );
  AND U58845 ( .A(n49353), .B(n49354), .Z(n49321) );
  NANDN U58846 ( .A(n49355), .B(n49356), .Z(n49354) );
  OR U58847 ( .A(n49357), .B(n49358), .Z(n49356) );
  IV U58848 ( .A(n49359), .Z(n49358) );
  NANDN U58849 ( .A(n49359), .B(n49357), .Z(n49353) );
  AND U58850 ( .A(n49360), .B(n49361), .Z(n49319) );
  NAND U58851 ( .A(n49362), .B(n49363), .Z(n49361) );
  NANDN U58852 ( .A(n49364), .B(n49365), .Z(n49363) );
  NANDN U58853 ( .A(n49365), .B(n49364), .Z(n49360) );
  IV U58854 ( .A(n49366), .Z(n49365) );
  NAND U58855 ( .A(n49367), .B(n49368), .Z(n49322) );
  NANDN U58856 ( .A(n49369), .B(n49370), .Z(n49368) );
  NANDN U58857 ( .A(n49371), .B(n49372), .Z(n49370) );
  NANDN U58858 ( .A(n49372), .B(n49371), .Z(n49367) );
  IV U58859 ( .A(n49373), .Z(n49371) );
  XOR U58860 ( .A(n49348), .B(n49374), .Z(N60996) );
  XNOR U58861 ( .A(n49351), .B(n49350), .Z(n49374) );
  XNOR U58862 ( .A(n49362), .B(n49375), .Z(n49350) );
  XNOR U58863 ( .A(n49366), .B(n49364), .Z(n49375) );
  XOR U58864 ( .A(n49372), .B(n49376), .Z(n49364) );
  XNOR U58865 ( .A(n49369), .B(n49373), .Z(n49376) );
  AND U58866 ( .A(n49377), .B(n49378), .Z(n49373) );
  NAND U58867 ( .A(n49379), .B(n49380), .Z(n49378) );
  NAND U58868 ( .A(n49381), .B(n49382), .Z(n49377) );
  AND U58869 ( .A(n49383), .B(n49384), .Z(n49369) );
  NAND U58870 ( .A(n49385), .B(n49386), .Z(n49384) );
  NAND U58871 ( .A(n49387), .B(n49388), .Z(n49383) );
  NANDN U58872 ( .A(n49389), .B(n49390), .Z(n49372) );
  ANDN U58873 ( .B(n49391), .A(n49392), .Z(n49366) );
  XNOR U58874 ( .A(n49357), .B(n49393), .Z(n49362) );
  XNOR U58875 ( .A(n49355), .B(n49359), .Z(n49393) );
  AND U58876 ( .A(n49394), .B(n49395), .Z(n49359) );
  NAND U58877 ( .A(n49396), .B(n49397), .Z(n49395) );
  NAND U58878 ( .A(n49398), .B(n49399), .Z(n49394) );
  AND U58879 ( .A(n49400), .B(n49401), .Z(n49355) );
  NAND U58880 ( .A(n49402), .B(n49403), .Z(n49401) );
  NAND U58881 ( .A(n49404), .B(n49405), .Z(n49400) );
  AND U58882 ( .A(n49406), .B(n49407), .Z(n49357) );
  NAND U58883 ( .A(n49408), .B(n49409), .Z(n49351) );
  XNOR U58884 ( .A(n49334), .B(n49410), .Z(n49348) );
  XNOR U58885 ( .A(n49338), .B(n49336), .Z(n49410) );
  XOR U58886 ( .A(n49344), .B(n49411), .Z(n49336) );
  XNOR U58887 ( .A(n49341), .B(n49345), .Z(n49411) );
  AND U58888 ( .A(n49412), .B(n49413), .Z(n49345) );
  NAND U58889 ( .A(n49414), .B(n49415), .Z(n49413) );
  NAND U58890 ( .A(n49416), .B(n49417), .Z(n49412) );
  AND U58891 ( .A(n49418), .B(n49419), .Z(n49341) );
  NAND U58892 ( .A(n49420), .B(n49421), .Z(n49419) );
  NAND U58893 ( .A(n49422), .B(n49423), .Z(n49418) );
  NANDN U58894 ( .A(n49424), .B(n49425), .Z(n49344) );
  ANDN U58895 ( .B(n49426), .A(n49427), .Z(n49338) );
  XNOR U58896 ( .A(n49329), .B(n49428), .Z(n49334) );
  XNOR U58897 ( .A(n49327), .B(n49331), .Z(n49428) );
  AND U58898 ( .A(n49429), .B(n49430), .Z(n49331) );
  NAND U58899 ( .A(n49431), .B(n49432), .Z(n49430) );
  NAND U58900 ( .A(n49433), .B(n49434), .Z(n49429) );
  AND U58901 ( .A(n49435), .B(n49436), .Z(n49327) );
  NAND U58902 ( .A(n49437), .B(n49438), .Z(n49436) );
  NAND U58903 ( .A(n49439), .B(n49440), .Z(n49435) );
  AND U58904 ( .A(n49441), .B(n49442), .Z(n49329) );
  XOR U58905 ( .A(n49409), .B(n49408), .Z(N60995) );
  XNOR U58906 ( .A(n49426), .B(n49427), .Z(n49408) );
  XNOR U58907 ( .A(n49441), .B(n49442), .Z(n49427) );
  XOR U58908 ( .A(n49438), .B(n49437), .Z(n49442) );
  XOR U58909 ( .A(y[756]), .B(x[756]), .Z(n49437) );
  XOR U58910 ( .A(n49440), .B(n49439), .Z(n49438) );
  XOR U58911 ( .A(y[758]), .B(x[758]), .Z(n49439) );
  XOR U58912 ( .A(y[757]), .B(x[757]), .Z(n49440) );
  XOR U58913 ( .A(n49432), .B(n49431), .Z(n49441) );
  XOR U58914 ( .A(n49434), .B(n49433), .Z(n49431) );
  XOR U58915 ( .A(y[755]), .B(x[755]), .Z(n49433) );
  XOR U58916 ( .A(y[754]), .B(x[754]), .Z(n49434) );
  XOR U58917 ( .A(y[753]), .B(x[753]), .Z(n49432) );
  XNOR U58918 ( .A(n49425), .B(n49424), .Z(n49426) );
  XNOR U58919 ( .A(n49421), .B(n49420), .Z(n49424) );
  XOR U58920 ( .A(n49423), .B(n49422), .Z(n49420) );
  XOR U58921 ( .A(y[752]), .B(x[752]), .Z(n49422) );
  XOR U58922 ( .A(y[751]), .B(x[751]), .Z(n49423) );
  XOR U58923 ( .A(y[750]), .B(x[750]), .Z(n49421) );
  XOR U58924 ( .A(n49415), .B(n49414), .Z(n49425) );
  XOR U58925 ( .A(n49417), .B(n49416), .Z(n49414) );
  XOR U58926 ( .A(y[749]), .B(x[749]), .Z(n49416) );
  XOR U58927 ( .A(y[748]), .B(x[748]), .Z(n49417) );
  XOR U58928 ( .A(y[747]), .B(x[747]), .Z(n49415) );
  XNOR U58929 ( .A(n49391), .B(n49392), .Z(n49409) );
  XNOR U58930 ( .A(n49406), .B(n49407), .Z(n49392) );
  XOR U58931 ( .A(n49403), .B(n49402), .Z(n49407) );
  XOR U58932 ( .A(y[744]), .B(x[744]), .Z(n49402) );
  XOR U58933 ( .A(n49405), .B(n49404), .Z(n49403) );
  XOR U58934 ( .A(y[746]), .B(x[746]), .Z(n49404) );
  XOR U58935 ( .A(y[745]), .B(x[745]), .Z(n49405) );
  XOR U58936 ( .A(n49397), .B(n49396), .Z(n49406) );
  XOR U58937 ( .A(n49399), .B(n49398), .Z(n49396) );
  XOR U58938 ( .A(y[743]), .B(x[743]), .Z(n49398) );
  XOR U58939 ( .A(y[742]), .B(x[742]), .Z(n49399) );
  XOR U58940 ( .A(y[741]), .B(x[741]), .Z(n49397) );
  XNOR U58941 ( .A(n49390), .B(n49389), .Z(n49391) );
  XNOR U58942 ( .A(n49386), .B(n49385), .Z(n49389) );
  XOR U58943 ( .A(n49388), .B(n49387), .Z(n49385) );
  XOR U58944 ( .A(y[740]), .B(x[740]), .Z(n49387) );
  XOR U58945 ( .A(y[739]), .B(x[739]), .Z(n49388) );
  XOR U58946 ( .A(y[738]), .B(x[738]), .Z(n49386) );
  XOR U58947 ( .A(n49380), .B(n49379), .Z(n49390) );
  XOR U58948 ( .A(n49382), .B(n49381), .Z(n49379) );
  XOR U58949 ( .A(y[737]), .B(x[737]), .Z(n49381) );
  XOR U58950 ( .A(y[736]), .B(x[736]), .Z(n49382) );
  XOR U58951 ( .A(y[735]), .B(x[735]), .Z(n49380) );
  NAND U58952 ( .A(n49443), .B(n49444), .Z(N60986) );
  NAND U58953 ( .A(n49445), .B(n49446), .Z(n49444) );
  NANDN U58954 ( .A(n49447), .B(n49448), .Z(n49446) );
  NANDN U58955 ( .A(n49448), .B(n49447), .Z(n49443) );
  XOR U58956 ( .A(n49447), .B(n49449), .Z(N60985) );
  XNOR U58957 ( .A(n49445), .B(n49448), .Z(n49449) );
  NAND U58958 ( .A(n49450), .B(n49451), .Z(n49448) );
  NAND U58959 ( .A(n49452), .B(n49453), .Z(n49451) );
  NANDN U58960 ( .A(n49454), .B(n49455), .Z(n49453) );
  NANDN U58961 ( .A(n49455), .B(n49454), .Z(n49450) );
  AND U58962 ( .A(n49456), .B(n49457), .Z(n49445) );
  NAND U58963 ( .A(n49458), .B(n49459), .Z(n49457) );
  NANDN U58964 ( .A(n49460), .B(n49461), .Z(n49459) );
  NANDN U58965 ( .A(n49461), .B(n49460), .Z(n49456) );
  IV U58966 ( .A(n49462), .Z(n49461) );
  AND U58967 ( .A(n49463), .B(n49464), .Z(n49447) );
  NAND U58968 ( .A(n49465), .B(n49466), .Z(n49464) );
  NANDN U58969 ( .A(n49467), .B(n49468), .Z(n49466) );
  NANDN U58970 ( .A(n49468), .B(n49467), .Z(n49463) );
  XOR U58971 ( .A(n49460), .B(n49469), .Z(N60984) );
  XNOR U58972 ( .A(n49458), .B(n49462), .Z(n49469) );
  XOR U58973 ( .A(n49455), .B(n49470), .Z(n49462) );
  XNOR U58974 ( .A(n49452), .B(n49454), .Z(n49470) );
  AND U58975 ( .A(n49471), .B(n49472), .Z(n49454) );
  NANDN U58976 ( .A(n49473), .B(n49474), .Z(n49472) );
  OR U58977 ( .A(n49475), .B(n49476), .Z(n49474) );
  IV U58978 ( .A(n49477), .Z(n49476) );
  NANDN U58979 ( .A(n49477), .B(n49475), .Z(n49471) );
  AND U58980 ( .A(n49478), .B(n49479), .Z(n49452) );
  NAND U58981 ( .A(n49480), .B(n49481), .Z(n49479) );
  NANDN U58982 ( .A(n49482), .B(n49483), .Z(n49481) );
  NANDN U58983 ( .A(n49483), .B(n49482), .Z(n49478) );
  IV U58984 ( .A(n49484), .Z(n49483) );
  NAND U58985 ( .A(n49485), .B(n49486), .Z(n49455) );
  NANDN U58986 ( .A(n49487), .B(n49488), .Z(n49486) );
  NANDN U58987 ( .A(n49489), .B(n49490), .Z(n49488) );
  NANDN U58988 ( .A(n49490), .B(n49489), .Z(n49485) );
  IV U58989 ( .A(n49491), .Z(n49489) );
  AND U58990 ( .A(n49492), .B(n49493), .Z(n49458) );
  NAND U58991 ( .A(n49494), .B(n49495), .Z(n49493) );
  NANDN U58992 ( .A(n49496), .B(n49497), .Z(n49495) );
  NANDN U58993 ( .A(n49497), .B(n49496), .Z(n49492) );
  XOR U58994 ( .A(n49468), .B(n49498), .Z(n49460) );
  XNOR U58995 ( .A(n49465), .B(n49467), .Z(n49498) );
  AND U58996 ( .A(n49499), .B(n49500), .Z(n49467) );
  NANDN U58997 ( .A(n49501), .B(n49502), .Z(n49500) );
  OR U58998 ( .A(n49503), .B(n49504), .Z(n49502) );
  IV U58999 ( .A(n49505), .Z(n49504) );
  NANDN U59000 ( .A(n49505), .B(n49503), .Z(n49499) );
  AND U59001 ( .A(n49506), .B(n49507), .Z(n49465) );
  NAND U59002 ( .A(n49508), .B(n49509), .Z(n49507) );
  NANDN U59003 ( .A(n49510), .B(n49511), .Z(n49509) );
  NANDN U59004 ( .A(n49511), .B(n49510), .Z(n49506) );
  IV U59005 ( .A(n49512), .Z(n49511) );
  NAND U59006 ( .A(n49513), .B(n49514), .Z(n49468) );
  NANDN U59007 ( .A(n49515), .B(n49516), .Z(n49514) );
  NANDN U59008 ( .A(n49517), .B(n49518), .Z(n49516) );
  NANDN U59009 ( .A(n49518), .B(n49517), .Z(n49513) );
  IV U59010 ( .A(n49519), .Z(n49517) );
  XOR U59011 ( .A(n49494), .B(n49520), .Z(N60983) );
  XNOR U59012 ( .A(n49497), .B(n49496), .Z(n49520) );
  XNOR U59013 ( .A(n49508), .B(n49521), .Z(n49496) );
  XNOR U59014 ( .A(n49512), .B(n49510), .Z(n49521) );
  XOR U59015 ( .A(n49518), .B(n49522), .Z(n49510) );
  XNOR U59016 ( .A(n49515), .B(n49519), .Z(n49522) );
  AND U59017 ( .A(n49523), .B(n49524), .Z(n49519) );
  NAND U59018 ( .A(n49525), .B(n49526), .Z(n49524) );
  NAND U59019 ( .A(n49527), .B(n49528), .Z(n49523) );
  AND U59020 ( .A(n49529), .B(n49530), .Z(n49515) );
  NAND U59021 ( .A(n49531), .B(n49532), .Z(n49530) );
  NAND U59022 ( .A(n49533), .B(n49534), .Z(n49529) );
  NANDN U59023 ( .A(n49535), .B(n49536), .Z(n49518) );
  ANDN U59024 ( .B(n49537), .A(n49538), .Z(n49512) );
  XNOR U59025 ( .A(n49503), .B(n49539), .Z(n49508) );
  XNOR U59026 ( .A(n49501), .B(n49505), .Z(n49539) );
  AND U59027 ( .A(n49540), .B(n49541), .Z(n49505) );
  NAND U59028 ( .A(n49542), .B(n49543), .Z(n49541) );
  NAND U59029 ( .A(n49544), .B(n49545), .Z(n49540) );
  AND U59030 ( .A(n49546), .B(n49547), .Z(n49501) );
  NAND U59031 ( .A(n49548), .B(n49549), .Z(n49547) );
  NAND U59032 ( .A(n49550), .B(n49551), .Z(n49546) );
  AND U59033 ( .A(n49552), .B(n49553), .Z(n49503) );
  NAND U59034 ( .A(n49554), .B(n49555), .Z(n49497) );
  XNOR U59035 ( .A(n49480), .B(n49556), .Z(n49494) );
  XNOR U59036 ( .A(n49484), .B(n49482), .Z(n49556) );
  XOR U59037 ( .A(n49490), .B(n49557), .Z(n49482) );
  XNOR U59038 ( .A(n49487), .B(n49491), .Z(n49557) );
  AND U59039 ( .A(n49558), .B(n49559), .Z(n49491) );
  NAND U59040 ( .A(n49560), .B(n49561), .Z(n49559) );
  NAND U59041 ( .A(n49562), .B(n49563), .Z(n49558) );
  AND U59042 ( .A(n49564), .B(n49565), .Z(n49487) );
  NAND U59043 ( .A(n49566), .B(n49567), .Z(n49565) );
  NAND U59044 ( .A(n49568), .B(n49569), .Z(n49564) );
  NANDN U59045 ( .A(n49570), .B(n49571), .Z(n49490) );
  ANDN U59046 ( .B(n49572), .A(n49573), .Z(n49484) );
  XNOR U59047 ( .A(n49475), .B(n49574), .Z(n49480) );
  XNOR U59048 ( .A(n49473), .B(n49477), .Z(n49574) );
  AND U59049 ( .A(n49575), .B(n49576), .Z(n49477) );
  NAND U59050 ( .A(n49577), .B(n49578), .Z(n49576) );
  NAND U59051 ( .A(n49579), .B(n49580), .Z(n49575) );
  AND U59052 ( .A(n49581), .B(n49582), .Z(n49473) );
  NAND U59053 ( .A(n49583), .B(n49584), .Z(n49582) );
  NAND U59054 ( .A(n49585), .B(n49586), .Z(n49581) );
  AND U59055 ( .A(n49587), .B(n49588), .Z(n49475) );
  XOR U59056 ( .A(n49555), .B(n49554), .Z(N60982) );
  XNOR U59057 ( .A(n49572), .B(n49573), .Z(n49554) );
  XNOR U59058 ( .A(n49587), .B(n49588), .Z(n49573) );
  XOR U59059 ( .A(n49584), .B(n49583), .Z(n49588) );
  XOR U59060 ( .A(y[732]), .B(x[732]), .Z(n49583) );
  XOR U59061 ( .A(n49586), .B(n49585), .Z(n49584) );
  XOR U59062 ( .A(y[734]), .B(x[734]), .Z(n49585) );
  XOR U59063 ( .A(y[733]), .B(x[733]), .Z(n49586) );
  XOR U59064 ( .A(n49578), .B(n49577), .Z(n49587) );
  XOR U59065 ( .A(n49580), .B(n49579), .Z(n49577) );
  XOR U59066 ( .A(y[731]), .B(x[731]), .Z(n49579) );
  XOR U59067 ( .A(y[730]), .B(x[730]), .Z(n49580) );
  XOR U59068 ( .A(y[729]), .B(x[729]), .Z(n49578) );
  XNOR U59069 ( .A(n49571), .B(n49570), .Z(n49572) );
  XNOR U59070 ( .A(n49567), .B(n49566), .Z(n49570) );
  XOR U59071 ( .A(n49569), .B(n49568), .Z(n49566) );
  XOR U59072 ( .A(y[728]), .B(x[728]), .Z(n49568) );
  XOR U59073 ( .A(y[727]), .B(x[727]), .Z(n49569) );
  XOR U59074 ( .A(y[726]), .B(x[726]), .Z(n49567) );
  XOR U59075 ( .A(n49561), .B(n49560), .Z(n49571) );
  XOR U59076 ( .A(n49563), .B(n49562), .Z(n49560) );
  XOR U59077 ( .A(y[725]), .B(x[725]), .Z(n49562) );
  XOR U59078 ( .A(y[724]), .B(x[724]), .Z(n49563) );
  XOR U59079 ( .A(y[723]), .B(x[723]), .Z(n49561) );
  XNOR U59080 ( .A(n49537), .B(n49538), .Z(n49555) );
  XNOR U59081 ( .A(n49552), .B(n49553), .Z(n49538) );
  XOR U59082 ( .A(n49549), .B(n49548), .Z(n49553) );
  XOR U59083 ( .A(y[720]), .B(x[720]), .Z(n49548) );
  XOR U59084 ( .A(n49551), .B(n49550), .Z(n49549) );
  XOR U59085 ( .A(y[722]), .B(x[722]), .Z(n49550) );
  XOR U59086 ( .A(y[721]), .B(x[721]), .Z(n49551) );
  XOR U59087 ( .A(n49543), .B(n49542), .Z(n49552) );
  XOR U59088 ( .A(n49545), .B(n49544), .Z(n49542) );
  XOR U59089 ( .A(y[719]), .B(x[719]), .Z(n49544) );
  XOR U59090 ( .A(y[718]), .B(x[718]), .Z(n49545) );
  XOR U59091 ( .A(y[717]), .B(x[717]), .Z(n49543) );
  XNOR U59092 ( .A(n49536), .B(n49535), .Z(n49537) );
  XNOR U59093 ( .A(n49532), .B(n49531), .Z(n49535) );
  XOR U59094 ( .A(n49534), .B(n49533), .Z(n49531) );
  XOR U59095 ( .A(y[716]), .B(x[716]), .Z(n49533) );
  XOR U59096 ( .A(y[715]), .B(x[715]), .Z(n49534) );
  XOR U59097 ( .A(y[714]), .B(x[714]), .Z(n49532) );
  XOR U59098 ( .A(n49526), .B(n49525), .Z(n49536) );
  XOR U59099 ( .A(n49528), .B(n49527), .Z(n49525) );
  XOR U59100 ( .A(y[713]), .B(x[713]), .Z(n49527) );
  XOR U59101 ( .A(y[712]), .B(x[712]), .Z(n49528) );
  XOR U59102 ( .A(y[711]), .B(x[711]), .Z(n49526) );
  NAND U59103 ( .A(n49589), .B(n49590), .Z(N60973) );
  NAND U59104 ( .A(n49591), .B(n49592), .Z(n49590) );
  NANDN U59105 ( .A(n49593), .B(n49594), .Z(n49592) );
  NANDN U59106 ( .A(n49594), .B(n49593), .Z(n49589) );
  XOR U59107 ( .A(n49593), .B(n49595), .Z(N60972) );
  XNOR U59108 ( .A(n49591), .B(n49594), .Z(n49595) );
  NAND U59109 ( .A(n49596), .B(n49597), .Z(n49594) );
  NAND U59110 ( .A(n49598), .B(n49599), .Z(n49597) );
  NANDN U59111 ( .A(n49600), .B(n49601), .Z(n49599) );
  NANDN U59112 ( .A(n49601), .B(n49600), .Z(n49596) );
  AND U59113 ( .A(n49602), .B(n49603), .Z(n49591) );
  NAND U59114 ( .A(n49604), .B(n49605), .Z(n49603) );
  NANDN U59115 ( .A(n49606), .B(n49607), .Z(n49605) );
  NANDN U59116 ( .A(n49607), .B(n49606), .Z(n49602) );
  IV U59117 ( .A(n49608), .Z(n49607) );
  AND U59118 ( .A(n49609), .B(n49610), .Z(n49593) );
  NAND U59119 ( .A(n49611), .B(n49612), .Z(n49610) );
  NANDN U59120 ( .A(n49613), .B(n49614), .Z(n49612) );
  NANDN U59121 ( .A(n49614), .B(n49613), .Z(n49609) );
  XOR U59122 ( .A(n49606), .B(n49615), .Z(N60971) );
  XNOR U59123 ( .A(n49604), .B(n49608), .Z(n49615) );
  XOR U59124 ( .A(n49601), .B(n49616), .Z(n49608) );
  XNOR U59125 ( .A(n49598), .B(n49600), .Z(n49616) );
  AND U59126 ( .A(n49617), .B(n49618), .Z(n49600) );
  NANDN U59127 ( .A(n49619), .B(n49620), .Z(n49618) );
  OR U59128 ( .A(n49621), .B(n49622), .Z(n49620) );
  IV U59129 ( .A(n49623), .Z(n49622) );
  NANDN U59130 ( .A(n49623), .B(n49621), .Z(n49617) );
  AND U59131 ( .A(n49624), .B(n49625), .Z(n49598) );
  NAND U59132 ( .A(n49626), .B(n49627), .Z(n49625) );
  NANDN U59133 ( .A(n49628), .B(n49629), .Z(n49627) );
  NANDN U59134 ( .A(n49629), .B(n49628), .Z(n49624) );
  IV U59135 ( .A(n49630), .Z(n49629) );
  NAND U59136 ( .A(n49631), .B(n49632), .Z(n49601) );
  NANDN U59137 ( .A(n49633), .B(n49634), .Z(n49632) );
  NANDN U59138 ( .A(n49635), .B(n49636), .Z(n49634) );
  NANDN U59139 ( .A(n49636), .B(n49635), .Z(n49631) );
  IV U59140 ( .A(n49637), .Z(n49635) );
  AND U59141 ( .A(n49638), .B(n49639), .Z(n49604) );
  NAND U59142 ( .A(n49640), .B(n49641), .Z(n49639) );
  NANDN U59143 ( .A(n49642), .B(n49643), .Z(n49641) );
  NANDN U59144 ( .A(n49643), .B(n49642), .Z(n49638) );
  XOR U59145 ( .A(n49614), .B(n49644), .Z(n49606) );
  XNOR U59146 ( .A(n49611), .B(n49613), .Z(n49644) );
  AND U59147 ( .A(n49645), .B(n49646), .Z(n49613) );
  NANDN U59148 ( .A(n49647), .B(n49648), .Z(n49646) );
  OR U59149 ( .A(n49649), .B(n49650), .Z(n49648) );
  IV U59150 ( .A(n49651), .Z(n49650) );
  NANDN U59151 ( .A(n49651), .B(n49649), .Z(n49645) );
  AND U59152 ( .A(n49652), .B(n49653), .Z(n49611) );
  NAND U59153 ( .A(n49654), .B(n49655), .Z(n49653) );
  NANDN U59154 ( .A(n49656), .B(n49657), .Z(n49655) );
  NANDN U59155 ( .A(n49657), .B(n49656), .Z(n49652) );
  IV U59156 ( .A(n49658), .Z(n49657) );
  NAND U59157 ( .A(n49659), .B(n49660), .Z(n49614) );
  NANDN U59158 ( .A(n49661), .B(n49662), .Z(n49660) );
  NANDN U59159 ( .A(n49663), .B(n49664), .Z(n49662) );
  NANDN U59160 ( .A(n49664), .B(n49663), .Z(n49659) );
  IV U59161 ( .A(n49665), .Z(n49663) );
  XOR U59162 ( .A(n49640), .B(n49666), .Z(N60970) );
  XNOR U59163 ( .A(n49643), .B(n49642), .Z(n49666) );
  XNOR U59164 ( .A(n49654), .B(n49667), .Z(n49642) );
  XNOR U59165 ( .A(n49658), .B(n49656), .Z(n49667) );
  XOR U59166 ( .A(n49664), .B(n49668), .Z(n49656) );
  XNOR U59167 ( .A(n49661), .B(n49665), .Z(n49668) );
  AND U59168 ( .A(n49669), .B(n49670), .Z(n49665) );
  NAND U59169 ( .A(n49671), .B(n49672), .Z(n49670) );
  NAND U59170 ( .A(n49673), .B(n49674), .Z(n49669) );
  AND U59171 ( .A(n49675), .B(n49676), .Z(n49661) );
  NAND U59172 ( .A(n49677), .B(n49678), .Z(n49676) );
  NAND U59173 ( .A(n49679), .B(n49680), .Z(n49675) );
  NANDN U59174 ( .A(n49681), .B(n49682), .Z(n49664) );
  ANDN U59175 ( .B(n49683), .A(n49684), .Z(n49658) );
  XNOR U59176 ( .A(n49649), .B(n49685), .Z(n49654) );
  XNOR U59177 ( .A(n49647), .B(n49651), .Z(n49685) );
  AND U59178 ( .A(n49686), .B(n49687), .Z(n49651) );
  NAND U59179 ( .A(n49688), .B(n49689), .Z(n49687) );
  NAND U59180 ( .A(n49690), .B(n49691), .Z(n49686) );
  AND U59181 ( .A(n49692), .B(n49693), .Z(n49647) );
  NAND U59182 ( .A(n49694), .B(n49695), .Z(n49693) );
  NAND U59183 ( .A(n49696), .B(n49697), .Z(n49692) );
  AND U59184 ( .A(n49698), .B(n49699), .Z(n49649) );
  NAND U59185 ( .A(n49700), .B(n49701), .Z(n49643) );
  XNOR U59186 ( .A(n49626), .B(n49702), .Z(n49640) );
  XNOR U59187 ( .A(n49630), .B(n49628), .Z(n49702) );
  XOR U59188 ( .A(n49636), .B(n49703), .Z(n49628) );
  XNOR U59189 ( .A(n49633), .B(n49637), .Z(n49703) );
  AND U59190 ( .A(n49704), .B(n49705), .Z(n49637) );
  NAND U59191 ( .A(n49706), .B(n49707), .Z(n49705) );
  NAND U59192 ( .A(n49708), .B(n49709), .Z(n49704) );
  AND U59193 ( .A(n49710), .B(n49711), .Z(n49633) );
  NAND U59194 ( .A(n49712), .B(n49713), .Z(n49711) );
  NAND U59195 ( .A(n49714), .B(n49715), .Z(n49710) );
  NANDN U59196 ( .A(n49716), .B(n49717), .Z(n49636) );
  ANDN U59197 ( .B(n49718), .A(n49719), .Z(n49630) );
  XNOR U59198 ( .A(n49621), .B(n49720), .Z(n49626) );
  XNOR U59199 ( .A(n49619), .B(n49623), .Z(n49720) );
  AND U59200 ( .A(n49721), .B(n49722), .Z(n49623) );
  NAND U59201 ( .A(n49723), .B(n49724), .Z(n49722) );
  NAND U59202 ( .A(n49725), .B(n49726), .Z(n49721) );
  AND U59203 ( .A(n49727), .B(n49728), .Z(n49619) );
  NAND U59204 ( .A(n49729), .B(n49730), .Z(n49728) );
  NAND U59205 ( .A(n49731), .B(n49732), .Z(n49727) );
  AND U59206 ( .A(n49733), .B(n49734), .Z(n49621) );
  XOR U59207 ( .A(n49701), .B(n49700), .Z(N60969) );
  XNOR U59208 ( .A(n49718), .B(n49719), .Z(n49700) );
  XNOR U59209 ( .A(n49733), .B(n49734), .Z(n49719) );
  XOR U59210 ( .A(n49730), .B(n49729), .Z(n49734) );
  XOR U59211 ( .A(y[708]), .B(x[708]), .Z(n49729) );
  XOR U59212 ( .A(n49732), .B(n49731), .Z(n49730) );
  XOR U59213 ( .A(y[710]), .B(x[710]), .Z(n49731) );
  XOR U59214 ( .A(y[709]), .B(x[709]), .Z(n49732) );
  XOR U59215 ( .A(n49724), .B(n49723), .Z(n49733) );
  XOR U59216 ( .A(n49726), .B(n49725), .Z(n49723) );
  XOR U59217 ( .A(y[707]), .B(x[707]), .Z(n49725) );
  XOR U59218 ( .A(y[706]), .B(x[706]), .Z(n49726) );
  XOR U59219 ( .A(y[705]), .B(x[705]), .Z(n49724) );
  XNOR U59220 ( .A(n49717), .B(n49716), .Z(n49718) );
  XNOR U59221 ( .A(n49713), .B(n49712), .Z(n49716) );
  XOR U59222 ( .A(n49715), .B(n49714), .Z(n49712) );
  XOR U59223 ( .A(y[704]), .B(x[704]), .Z(n49714) );
  XOR U59224 ( .A(y[703]), .B(x[703]), .Z(n49715) );
  XOR U59225 ( .A(y[702]), .B(x[702]), .Z(n49713) );
  XOR U59226 ( .A(n49707), .B(n49706), .Z(n49717) );
  XOR U59227 ( .A(n49709), .B(n49708), .Z(n49706) );
  XOR U59228 ( .A(y[701]), .B(x[701]), .Z(n49708) );
  XOR U59229 ( .A(y[700]), .B(x[700]), .Z(n49709) );
  XOR U59230 ( .A(y[699]), .B(x[699]), .Z(n49707) );
  XNOR U59231 ( .A(n49683), .B(n49684), .Z(n49701) );
  XNOR U59232 ( .A(n49698), .B(n49699), .Z(n49684) );
  XOR U59233 ( .A(n49695), .B(n49694), .Z(n49699) );
  XOR U59234 ( .A(y[696]), .B(x[696]), .Z(n49694) );
  XOR U59235 ( .A(n49697), .B(n49696), .Z(n49695) );
  XOR U59236 ( .A(y[698]), .B(x[698]), .Z(n49696) );
  XOR U59237 ( .A(y[697]), .B(x[697]), .Z(n49697) );
  XOR U59238 ( .A(n49689), .B(n49688), .Z(n49698) );
  XOR U59239 ( .A(n49691), .B(n49690), .Z(n49688) );
  XOR U59240 ( .A(y[695]), .B(x[695]), .Z(n49690) );
  XOR U59241 ( .A(y[694]), .B(x[694]), .Z(n49691) );
  XOR U59242 ( .A(y[693]), .B(x[693]), .Z(n49689) );
  XNOR U59243 ( .A(n49682), .B(n49681), .Z(n49683) );
  XNOR U59244 ( .A(n49678), .B(n49677), .Z(n49681) );
  XOR U59245 ( .A(n49680), .B(n49679), .Z(n49677) );
  XOR U59246 ( .A(y[692]), .B(x[692]), .Z(n49679) );
  XOR U59247 ( .A(y[691]), .B(x[691]), .Z(n49680) );
  XOR U59248 ( .A(y[690]), .B(x[690]), .Z(n49678) );
  XOR U59249 ( .A(n49672), .B(n49671), .Z(n49682) );
  XOR U59250 ( .A(n49674), .B(n49673), .Z(n49671) );
  XOR U59251 ( .A(y[689]), .B(x[689]), .Z(n49673) );
  XOR U59252 ( .A(y[688]), .B(x[688]), .Z(n49674) );
  XOR U59253 ( .A(y[687]), .B(x[687]), .Z(n49672) );
  NAND U59254 ( .A(n49735), .B(n49736), .Z(N60960) );
  NAND U59255 ( .A(n49737), .B(n49738), .Z(n49736) );
  NANDN U59256 ( .A(n49739), .B(n49740), .Z(n49738) );
  NANDN U59257 ( .A(n49740), .B(n49739), .Z(n49735) );
  XOR U59258 ( .A(n49739), .B(n49741), .Z(N60959) );
  XNOR U59259 ( .A(n49737), .B(n49740), .Z(n49741) );
  NAND U59260 ( .A(n49742), .B(n49743), .Z(n49740) );
  NAND U59261 ( .A(n49744), .B(n49745), .Z(n49743) );
  NANDN U59262 ( .A(n49746), .B(n49747), .Z(n49745) );
  NANDN U59263 ( .A(n49747), .B(n49746), .Z(n49742) );
  AND U59264 ( .A(n49748), .B(n49749), .Z(n49737) );
  NAND U59265 ( .A(n49750), .B(n49751), .Z(n49749) );
  NANDN U59266 ( .A(n49752), .B(n49753), .Z(n49751) );
  NANDN U59267 ( .A(n49753), .B(n49752), .Z(n49748) );
  IV U59268 ( .A(n49754), .Z(n49753) );
  AND U59269 ( .A(n49755), .B(n49756), .Z(n49739) );
  NAND U59270 ( .A(n49757), .B(n49758), .Z(n49756) );
  NANDN U59271 ( .A(n49759), .B(n49760), .Z(n49758) );
  NANDN U59272 ( .A(n49760), .B(n49759), .Z(n49755) );
  XOR U59273 ( .A(n49752), .B(n49761), .Z(N60958) );
  XNOR U59274 ( .A(n49750), .B(n49754), .Z(n49761) );
  XOR U59275 ( .A(n49747), .B(n49762), .Z(n49754) );
  XNOR U59276 ( .A(n49744), .B(n49746), .Z(n49762) );
  AND U59277 ( .A(n49763), .B(n49764), .Z(n49746) );
  NANDN U59278 ( .A(n49765), .B(n49766), .Z(n49764) );
  OR U59279 ( .A(n49767), .B(n49768), .Z(n49766) );
  IV U59280 ( .A(n49769), .Z(n49768) );
  NANDN U59281 ( .A(n49769), .B(n49767), .Z(n49763) );
  AND U59282 ( .A(n49770), .B(n49771), .Z(n49744) );
  NAND U59283 ( .A(n49772), .B(n49773), .Z(n49771) );
  NANDN U59284 ( .A(n49774), .B(n49775), .Z(n49773) );
  NANDN U59285 ( .A(n49775), .B(n49774), .Z(n49770) );
  IV U59286 ( .A(n49776), .Z(n49775) );
  NAND U59287 ( .A(n49777), .B(n49778), .Z(n49747) );
  NANDN U59288 ( .A(n49779), .B(n49780), .Z(n49778) );
  NANDN U59289 ( .A(n49781), .B(n49782), .Z(n49780) );
  NANDN U59290 ( .A(n49782), .B(n49781), .Z(n49777) );
  IV U59291 ( .A(n49783), .Z(n49781) );
  AND U59292 ( .A(n49784), .B(n49785), .Z(n49750) );
  NAND U59293 ( .A(n49786), .B(n49787), .Z(n49785) );
  NANDN U59294 ( .A(n49788), .B(n49789), .Z(n49787) );
  NANDN U59295 ( .A(n49789), .B(n49788), .Z(n49784) );
  XOR U59296 ( .A(n49760), .B(n49790), .Z(n49752) );
  XNOR U59297 ( .A(n49757), .B(n49759), .Z(n49790) );
  AND U59298 ( .A(n49791), .B(n49792), .Z(n49759) );
  NANDN U59299 ( .A(n49793), .B(n49794), .Z(n49792) );
  OR U59300 ( .A(n49795), .B(n49796), .Z(n49794) );
  IV U59301 ( .A(n49797), .Z(n49796) );
  NANDN U59302 ( .A(n49797), .B(n49795), .Z(n49791) );
  AND U59303 ( .A(n49798), .B(n49799), .Z(n49757) );
  NAND U59304 ( .A(n49800), .B(n49801), .Z(n49799) );
  NANDN U59305 ( .A(n49802), .B(n49803), .Z(n49801) );
  NANDN U59306 ( .A(n49803), .B(n49802), .Z(n49798) );
  IV U59307 ( .A(n49804), .Z(n49803) );
  NAND U59308 ( .A(n49805), .B(n49806), .Z(n49760) );
  NANDN U59309 ( .A(n49807), .B(n49808), .Z(n49806) );
  NANDN U59310 ( .A(n49809), .B(n49810), .Z(n49808) );
  NANDN U59311 ( .A(n49810), .B(n49809), .Z(n49805) );
  IV U59312 ( .A(n49811), .Z(n49809) );
  XOR U59313 ( .A(n49786), .B(n49812), .Z(N60957) );
  XNOR U59314 ( .A(n49789), .B(n49788), .Z(n49812) );
  XNOR U59315 ( .A(n49800), .B(n49813), .Z(n49788) );
  XNOR U59316 ( .A(n49804), .B(n49802), .Z(n49813) );
  XOR U59317 ( .A(n49810), .B(n49814), .Z(n49802) );
  XNOR U59318 ( .A(n49807), .B(n49811), .Z(n49814) );
  AND U59319 ( .A(n49815), .B(n49816), .Z(n49811) );
  NAND U59320 ( .A(n49817), .B(n49818), .Z(n49816) );
  NAND U59321 ( .A(n49819), .B(n49820), .Z(n49815) );
  AND U59322 ( .A(n49821), .B(n49822), .Z(n49807) );
  NAND U59323 ( .A(n49823), .B(n49824), .Z(n49822) );
  NAND U59324 ( .A(n49825), .B(n49826), .Z(n49821) );
  NANDN U59325 ( .A(n49827), .B(n49828), .Z(n49810) );
  ANDN U59326 ( .B(n49829), .A(n49830), .Z(n49804) );
  XNOR U59327 ( .A(n49795), .B(n49831), .Z(n49800) );
  XNOR U59328 ( .A(n49793), .B(n49797), .Z(n49831) );
  AND U59329 ( .A(n49832), .B(n49833), .Z(n49797) );
  NAND U59330 ( .A(n49834), .B(n49835), .Z(n49833) );
  NAND U59331 ( .A(n49836), .B(n49837), .Z(n49832) );
  AND U59332 ( .A(n49838), .B(n49839), .Z(n49793) );
  NAND U59333 ( .A(n49840), .B(n49841), .Z(n49839) );
  NAND U59334 ( .A(n49842), .B(n49843), .Z(n49838) );
  AND U59335 ( .A(n49844), .B(n49845), .Z(n49795) );
  NAND U59336 ( .A(n49846), .B(n49847), .Z(n49789) );
  XNOR U59337 ( .A(n49772), .B(n49848), .Z(n49786) );
  XNOR U59338 ( .A(n49776), .B(n49774), .Z(n49848) );
  XOR U59339 ( .A(n49782), .B(n49849), .Z(n49774) );
  XNOR U59340 ( .A(n49779), .B(n49783), .Z(n49849) );
  AND U59341 ( .A(n49850), .B(n49851), .Z(n49783) );
  NAND U59342 ( .A(n49852), .B(n49853), .Z(n49851) );
  NAND U59343 ( .A(n49854), .B(n49855), .Z(n49850) );
  AND U59344 ( .A(n49856), .B(n49857), .Z(n49779) );
  NAND U59345 ( .A(n49858), .B(n49859), .Z(n49857) );
  NAND U59346 ( .A(n49860), .B(n49861), .Z(n49856) );
  NANDN U59347 ( .A(n49862), .B(n49863), .Z(n49782) );
  ANDN U59348 ( .B(n49864), .A(n49865), .Z(n49776) );
  XNOR U59349 ( .A(n49767), .B(n49866), .Z(n49772) );
  XNOR U59350 ( .A(n49765), .B(n49769), .Z(n49866) );
  AND U59351 ( .A(n49867), .B(n49868), .Z(n49769) );
  NAND U59352 ( .A(n49869), .B(n49870), .Z(n49868) );
  NAND U59353 ( .A(n49871), .B(n49872), .Z(n49867) );
  AND U59354 ( .A(n49873), .B(n49874), .Z(n49765) );
  NAND U59355 ( .A(n49875), .B(n49876), .Z(n49874) );
  NAND U59356 ( .A(n49877), .B(n49878), .Z(n49873) );
  AND U59357 ( .A(n49879), .B(n49880), .Z(n49767) );
  XOR U59358 ( .A(n49847), .B(n49846), .Z(N60956) );
  XNOR U59359 ( .A(n49864), .B(n49865), .Z(n49846) );
  XNOR U59360 ( .A(n49879), .B(n49880), .Z(n49865) );
  XOR U59361 ( .A(n49876), .B(n49875), .Z(n49880) );
  XOR U59362 ( .A(y[684]), .B(x[684]), .Z(n49875) );
  XOR U59363 ( .A(n49878), .B(n49877), .Z(n49876) );
  XOR U59364 ( .A(y[686]), .B(x[686]), .Z(n49877) );
  XOR U59365 ( .A(y[685]), .B(x[685]), .Z(n49878) );
  XOR U59366 ( .A(n49870), .B(n49869), .Z(n49879) );
  XOR U59367 ( .A(n49872), .B(n49871), .Z(n49869) );
  XOR U59368 ( .A(y[683]), .B(x[683]), .Z(n49871) );
  XOR U59369 ( .A(y[682]), .B(x[682]), .Z(n49872) );
  XOR U59370 ( .A(y[681]), .B(x[681]), .Z(n49870) );
  XNOR U59371 ( .A(n49863), .B(n49862), .Z(n49864) );
  XNOR U59372 ( .A(n49859), .B(n49858), .Z(n49862) );
  XOR U59373 ( .A(n49861), .B(n49860), .Z(n49858) );
  XOR U59374 ( .A(y[680]), .B(x[680]), .Z(n49860) );
  XOR U59375 ( .A(y[679]), .B(x[679]), .Z(n49861) );
  XOR U59376 ( .A(y[678]), .B(x[678]), .Z(n49859) );
  XOR U59377 ( .A(n49853), .B(n49852), .Z(n49863) );
  XOR U59378 ( .A(n49855), .B(n49854), .Z(n49852) );
  XOR U59379 ( .A(y[677]), .B(x[677]), .Z(n49854) );
  XOR U59380 ( .A(y[676]), .B(x[676]), .Z(n49855) );
  XOR U59381 ( .A(y[675]), .B(x[675]), .Z(n49853) );
  XNOR U59382 ( .A(n49829), .B(n49830), .Z(n49847) );
  XNOR U59383 ( .A(n49844), .B(n49845), .Z(n49830) );
  XOR U59384 ( .A(n49841), .B(n49840), .Z(n49845) );
  XOR U59385 ( .A(y[672]), .B(x[672]), .Z(n49840) );
  XOR U59386 ( .A(n49843), .B(n49842), .Z(n49841) );
  XOR U59387 ( .A(y[674]), .B(x[674]), .Z(n49842) );
  XOR U59388 ( .A(y[673]), .B(x[673]), .Z(n49843) );
  XOR U59389 ( .A(n49835), .B(n49834), .Z(n49844) );
  XOR U59390 ( .A(n49837), .B(n49836), .Z(n49834) );
  XOR U59391 ( .A(y[671]), .B(x[671]), .Z(n49836) );
  XOR U59392 ( .A(y[670]), .B(x[670]), .Z(n49837) );
  XOR U59393 ( .A(y[669]), .B(x[669]), .Z(n49835) );
  XNOR U59394 ( .A(n49828), .B(n49827), .Z(n49829) );
  XNOR U59395 ( .A(n49824), .B(n49823), .Z(n49827) );
  XOR U59396 ( .A(n49826), .B(n49825), .Z(n49823) );
  XOR U59397 ( .A(y[668]), .B(x[668]), .Z(n49825) );
  XOR U59398 ( .A(y[667]), .B(x[667]), .Z(n49826) );
  XOR U59399 ( .A(y[666]), .B(x[666]), .Z(n49824) );
  XOR U59400 ( .A(n49818), .B(n49817), .Z(n49828) );
  XOR U59401 ( .A(n49820), .B(n49819), .Z(n49817) );
  XOR U59402 ( .A(y[665]), .B(x[665]), .Z(n49819) );
  XOR U59403 ( .A(y[664]), .B(x[664]), .Z(n49820) );
  XOR U59404 ( .A(y[663]), .B(x[663]), .Z(n49818) );
  NAND U59405 ( .A(n49881), .B(n49882), .Z(N60947) );
  NAND U59406 ( .A(n49883), .B(n49884), .Z(n49882) );
  NANDN U59407 ( .A(n49885), .B(n49886), .Z(n49884) );
  NANDN U59408 ( .A(n49886), .B(n49885), .Z(n49881) );
  XOR U59409 ( .A(n49885), .B(n49887), .Z(N60946) );
  XNOR U59410 ( .A(n49883), .B(n49886), .Z(n49887) );
  NAND U59411 ( .A(n49888), .B(n49889), .Z(n49886) );
  NAND U59412 ( .A(n49890), .B(n49891), .Z(n49889) );
  NANDN U59413 ( .A(n49892), .B(n49893), .Z(n49891) );
  NANDN U59414 ( .A(n49893), .B(n49892), .Z(n49888) );
  AND U59415 ( .A(n49894), .B(n49895), .Z(n49883) );
  NAND U59416 ( .A(n49896), .B(n49897), .Z(n49895) );
  NANDN U59417 ( .A(n49898), .B(n49899), .Z(n49897) );
  NANDN U59418 ( .A(n49899), .B(n49898), .Z(n49894) );
  IV U59419 ( .A(n49900), .Z(n49899) );
  AND U59420 ( .A(n49901), .B(n49902), .Z(n49885) );
  NAND U59421 ( .A(n49903), .B(n49904), .Z(n49902) );
  NANDN U59422 ( .A(n49905), .B(n49906), .Z(n49904) );
  NANDN U59423 ( .A(n49906), .B(n49905), .Z(n49901) );
  XOR U59424 ( .A(n49898), .B(n49907), .Z(N60945) );
  XNOR U59425 ( .A(n49896), .B(n49900), .Z(n49907) );
  XOR U59426 ( .A(n49893), .B(n49908), .Z(n49900) );
  XNOR U59427 ( .A(n49890), .B(n49892), .Z(n49908) );
  AND U59428 ( .A(n49909), .B(n49910), .Z(n49892) );
  NANDN U59429 ( .A(n49911), .B(n49912), .Z(n49910) );
  OR U59430 ( .A(n49913), .B(n49914), .Z(n49912) );
  IV U59431 ( .A(n49915), .Z(n49914) );
  NANDN U59432 ( .A(n49915), .B(n49913), .Z(n49909) );
  AND U59433 ( .A(n49916), .B(n49917), .Z(n49890) );
  NAND U59434 ( .A(n49918), .B(n49919), .Z(n49917) );
  NANDN U59435 ( .A(n49920), .B(n49921), .Z(n49919) );
  NANDN U59436 ( .A(n49921), .B(n49920), .Z(n49916) );
  IV U59437 ( .A(n49922), .Z(n49921) );
  NAND U59438 ( .A(n49923), .B(n49924), .Z(n49893) );
  NANDN U59439 ( .A(n49925), .B(n49926), .Z(n49924) );
  NANDN U59440 ( .A(n49927), .B(n49928), .Z(n49926) );
  NANDN U59441 ( .A(n49928), .B(n49927), .Z(n49923) );
  IV U59442 ( .A(n49929), .Z(n49927) );
  AND U59443 ( .A(n49930), .B(n49931), .Z(n49896) );
  NAND U59444 ( .A(n49932), .B(n49933), .Z(n49931) );
  NANDN U59445 ( .A(n49934), .B(n49935), .Z(n49933) );
  NANDN U59446 ( .A(n49935), .B(n49934), .Z(n49930) );
  XOR U59447 ( .A(n49906), .B(n49936), .Z(n49898) );
  XNOR U59448 ( .A(n49903), .B(n49905), .Z(n49936) );
  AND U59449 ( .A(n49937), .B(n49938), .Z(n49905) );
  NANDN U59450 ( .A(n49939), .B(n49940), .Z(n49938) );
  OR U59451 ( .A(n49941), .B(n49942), .Z(n49940) );
  IV U59452 ( .A(n49943), .Z(n49942) );
  NANDN U59453 ( .A(n49943), .B(n49941), .Z(n49937) );
  AND U59454 ( .A(n49944), .B(n49945), .Z(n49903) );
  NAND U59455 ( .A(n49946), .B(n49947), .Z(n49945) );
  NANDN U59456 ( .A(n49948), .B(n49949), .Z(n49947) );
  NANDN U59457 ( .A(n49949), .B(n49948), .Z(n49944) );
  IV U59458 ( .A(n49950), .Z(n49949) );
  NAND U59459 ( .A(n49951), .B(n49952), .Z(n49906) );
  NANDN U59460 ( .A(n49953), .B(n49954), .Z(n49952) );
  NANDN U59461 ( .A(n49955), .B(n49956), .Z(n49954) );
  NANDN U59462 ( .A(n49956), .B(n49955), .Z(n49951) );
  IV U59463 ( .A(n49957), .Z(n49955) );
  XOR U59464 ( .A(n49932), .B(n49958), .Z(N60944) );
  XNOR U59465 ( .A(n49935), .B(n49934), .Z(n49958) );
  XNOR U59466 ( .A(n49946), .B(n49959), .Z(n49934) );
  XNOR U59467 ( .A(n49950), .B(n49948), .Z(n49959) );
  XOR U59468 ( .A(n49956), .B(n49960), .Z(n49948) );
  XNOR U59469 ( .A(n49953), .B(n49957), .Z(n49960) );
  AND U59470 ( .A(n49961), .B(n49962), .Z(n49957) );
  NAND U59471 ( .A(n49963), .B(n49964), .Z(n49962) );
  NAND U59472 ( .A(n49965), .B(n49966), .Z(n49961) );
  AND U59473 ( .A(n49967), .B(n49968), .Z(n49953) );
  NAND U59474 ( .A(n49969), .B(n49970), .Z(n49968) );
  NAND U59475 ( .A(n49971), .B(n49972), .Z(n49967) );
  NANDN U59476 ( .A(n49973), .B(n49974), .Z(n49956) );
  ANDN U59477 ( .B(n49975), .A(n49976), .Z(n49950) );
  XNOR U59478 ( .A(n49941), .B(n49977), .Z(n49946) );
  XNOR U59479 ( .A(n49939), .B(n49943), .Z(n49977) );
  AND U59480 ( .A(n49978), .B(n49979), .Z(n49943) );
  NAND U59481 ( .A(n49980), .B(n49981), .Z(n49979) );
  NAND U59482 ( .A(n49982), .B(n49983), .Z(n49978) );
  AND U59483 ( .A(n49984), .B(n49985), .Z(n49939) );
  NAND U59484 ( .A(n49986), .B(n49987), .Z(n49985) );
  NAND U59485 ( .A(n49988), .B(n49989), .Z(n49984) );
  AND U59486 ( .A(n49990), .B(n49991), .Z(n49941) );
  NAND U59487 ( .A(n49992), .B(n49993), .Z(n49935) );
  XNOR U59488 ( .A(n49918), .B(n49994), .Z(n49932) );
  XNOR U59489 ( .A(n49922), .B(n49920), .Z(n49994) );
  XOR U59490 ( .A(n49928), .B(n49995), .Z(n49920) );
  XNOR U59491 ( .A(n49925), .B(n49929), .Z(n49995) );
  AND U59492 ( .A(n49996), .B(n49997), .Z(n49929) );
  NAND U59493 ( .A(n49998), .B(n49999), .Z(n49997) );
  NAND U59494 ( .A(n50000), .B(n50001), .Z(n49996) );
  AND U59495 ( .A(n50002), .B(n50003), .Z(n49925) );
  NAND U59496 ( .A(n50004), .B(n50005), .Z(n50003) );
  NAND U59497 ( .A(n50006), .B(n50007), .Z(n50002) );
  NANDN U59498 ( .A(n50008), .B(n50009), .Z(n49928) );
  ANDN U59499 ( .B(n50010), .A(n50011), .Z(n49922) );
  XNOR U59500 ( .A(n49913), .B(n50012), .Z(n49918) );
  XNOR U59501 ( .A(n49911), .B(n49915), .Z(n50012) );
  AND U59502 ( .A(n50013), .B(n50014), .Z(n49915) );
  NAND U59503 ( .A(n50015), .B(n50016), .Z(n50014) );
  NAND U59504 ( .A(n50017), .B(n50018), .Z(n50013) );
  AND U59505 ( .A(n50019), .B(n50020), .Z(n49911) );
  NAND U59506 ( .A(n50021), .B(n50022), .Z(n50020) );
  NAND U59507 ( .A(n50023), .B(n50024), .Z(n50019) );
  AND U59508 ( .A(n50025), .B(n50026), .Z(n49913) );
  XOR U59509 ( .A(n49993), .B(n49992), .Z(N60943) );
  XNOR U59510 ( .A(n50010), .B(n50011), .Z(n49992) );
  XNOR U59511 ( .A(n50025), .B(n50026), .Z(n50011) );
  XOR U59512 ( .A(n50022), .B(n50021), .Z(n50026) );
  XOR U59513 ( .A(y[660]), .B(x[660]), .Z(n50021) );
  XOR U59514 ( .A(n50024), .B(n50023), .Z(n50022) );
  XOR U59515 ( .A(y[662]), .B(x[662]), .Z(n50023) );
  XOR U59516 ( .A(y[661]), .B(x[661]), .Z(n50024) );
  XOR U59517 ( .A(n50016), .B(n50015), .Z(n50025) );
  XOR U59518 ( .A(n50018), .B(n50017), .Z(n50015) );
  XOR U59519 ( .A(y[659]), .B(x[659]), .Z(n50017) );
  XOR U59520 ( .A(y[658]), .B(x[658]), .Z(n50018) );
  XOR U59521 ( .A(y[657]), .B(x[657]), .Z(n50016) );
  XNOR U59522 ( .A(n50009), .B(n50008), .Z(n50010) );
  XNOR U59523 ( .A(n50005), .B(n50004), .Z(n50008) );
  XOR U59524 ( .A(n50007), .B(n50006), .Z(n50004) );
  XOR U59525 ( .A(y[656]), .B(x[656]), .Z(n50006) );
  XOR U59526 ( .A(y[655]), .B(x[655]), .Z(n50007) );
  XOR U59527 ( .A(y[654]), .B(x[654]), .Z(n50005) );
  XOR U59528 ( .A(n49999), .B(n49998), .Z(n50009) );
  XOR U59529 ( .A(n50001), .B(n50000), .Z(n49998) );
  XOR U59530 ( .A(y[653]), .B(x[653]), .Z(n50000) );
  XOR U59531 ( .A(y[652]), .B(x[652]), .Z(n50001) );
  XOR U59532 ( .A(y[651]), .B(x[651]), .Z(n49999) );
  XNOR U59533 ( .A(n49975), .B(n49976), .Z(n49993) );
  XNOR U59534 ( .A(n49990), .B(n49991), .Z(n49976) );
  XOR U59535 ( .A(n49987), .B(n49986), .Z(n49991) );
  XOR U59536 ( .A(y[648]), .B(x[648]), .Z(n49986) );
  XOR U59537 ( .A(n49989), .B(n49988), .Z(n49987) );
  XOR U59538 ( .A(y[650]), .B(x[650]), .Z(n49988) );
  XOR U59539 ( .A(y[649]), .B(x[649]), .Z(n49989) );
  XOR U59540 ( .A(n49981), .B(n49980), .Z(n49990) );
  XOR U59541 ( .A(n49983), .B(n49982), .Z(n49980) );
  XOR U59542 ( .A(y[647]), .B(x[647]), .Z(n49982) );
  XOR U59543 ( .A(y[646]), .B(x[646]), .Z(n49983) );
  XOR U59544 ( .A(y[645]), .B(x[645]), .Z(n49981) );
  XNOR U59545 ( .A(n49974), .B(n49973), .Z(n49975) );
  XNOR U59546 ( .A(n49970), .B(n49969), .Z(n49973) );
  XOR U59547 ( .A(n49972), .B(n49971), .Z(n49969) );
  XOR U59548 ( .A(y[644]), .B(x[644]), .Z(n49971) );
  XOR U59549 ( .A(y[643]), .B(x[643]), .Z(n49972) );
  XOR U59550 ( .A(y[642]), .B(x[642]), .Z(n49970) );
  XOR U59551 ( .A(n49964), .B(n49963), .Z(n49974) );
  XOR U59552 ( .A(n49966), .B(n49965), .Z(n49963) );
  XOR U59553 ( .A(y[641]), .B(x[641]), .Z(n49965) );
  XOR U59554 ( .A(y[640]), .B(x[640]), .Z(n49966) );
  XOR U59555 ( .A(y[639]), .B(x[639]), .Z(n49964) );
  NAND U59556 ( .A(n50027), .B(n50028), .Z(N60934) );
  NAND U59557 ( .A(n50029), .B(n50030), .Z(n50028) );
  NANDN U59558 ( .A(n50031), .B(n50032), .Z(n50030) );
  NANDN U59559 ( .A(n50032), .B(n50031), .Z(n50027) );
  XOR U59560 ( .A(n50031), .B(n50033), .Z(N60933) );
  XNOR U59561 ( .A(n50029), .B(n50032), .Z(n50033) );
  NAND U59562 ( .A(n50034), .B(n50035), .Z(n50032) );
  NAND U59563 ( .A(n50036), .B(n50037), .Z(n50035) );
  NANDN U59564 ( .A(n50038), .B(n50039), .Z(n50037) );
  NANDN U59565 ( .A(n50039), .B(n50038), .Z(n50034) );
  AND U59566 ( .A(n50040), .B(n50041), .Z(n50029) );
  NAND U59567 ( .A(n50042), .B(n50043), .Z(n50041) );
  NANDN U59568 ( .A(n50044), .B(n50045), .Z(n50043) );
  NANDN U59569 ( .A(n50045), .B(n50044), .Z(n50040) );
  IV U59570 ( .A(n50046), .Z(n50045) );
  AND U59571 ( .A(n50047), .B(n50048), .Z(n50031) );
  NAND U59572 ( .A(n50049), .B(n50050), .Z(n50048) );
  NANDN U59573 ( .A(n50051), .B(n50052), .Z(n50050) );
  NANDN U59574 ( .A(n50052), .B(n50051), .Z(n50047) );
  XOR U59575 ( .A(n50044), .B(n50053), .Z(N60932) );
  XNOR U59576 ( .A(n50042), .B(n50046), .Z(n50053) );
  XOR U59577 ( .A(n50039), .B(n50054), .Z(n50046) );
  XNOR U59578 ( .A(n50036), .B(n50038), .Z(n50054) );
  AND U59579 ( .A(n50055), .B(n50056), .Z(n50038) );
  NANDN U59580 ( .A(n50057), .B(n50058), .Z(n50056) );
  OR U59581 ( .A(n50059), .B(n50060), .Z(n50058) );
  IV U59582 ( .A(n50061), .Z(n50060) );
  NANDN U59583 ( .A(n50061), .B(n50059), .Z(n50055) );
  AND U59584 ( .A(n50062), .B(n50063), .Z(n50036) );
  NAND U59585 ( .A(n50064), .B(n50065), .Z(n50063) );
  NANDN U59586 ( .A(n50066), .B(n50067), .Z(n50065) );
  NANDN U59587 ( .A(n50067), .B(n50066), .Z(n50062) );
  IV U59588 ( .A(n50068), .Z(n50067) );
  NAND U59589 ( .A(n50069), .B(n50070), .Z(n50039) );
  NANDN U59590 ( .A(n50071), .B(n50072), .Z(n50070) );
  NANDN U59591 ( .A(n50073), .B(n50074), .Z(n50072) );
  NANDN U59592 ( .A(n50074), .B(n50073), .Z(n50069) );
  IV U59593 ( .A(n50075), .Z(n50073) );
  AND U59594 ( .A(n50076), .B(n50077), .Z(n50042) );
  NAND U59595 ( .A(n50078), .B(n50079), .Z(n50077) );
  NANDN U59596 ( .A(n50080), .B(n50081), .Z(n50079) );
  NANDN U59597 ( .A(n50081), .B(n50080), .Z(n50076) );
  XOR U59598 ( .A(n50052), .B(n50082), .Z(n50044) );
  XNOR U59599 ( .A(n50049), .B(n50051), .Z(n50082) );
  AND U59600 ( .A(n50083), .B(n50084), .Z(n50051) );
  NANDN U59601 ( .A(n50085), .B(n50086), .Z(n50084) );
  OR U59602 ( .A(n50087), .B(n50088), .Z(n50086) );
  IV U59603 ( .A(n50089), .Z(n50088) );
  NANDN U59604 ( .A(n50089), .B(n50087), .Z(n50083) );
  AND U59605 ( .A(n50090), .B(n50091), .Z(n50049) );
  NAND U59606 ( .A(n50092), .B(n50093), .Z(n50091) );
  NANDN U59607 ( .A(n50094), .B(n50095), .Z(n50093) );
  NANDN U59608 ( .A(n50095), .B(n50094), .Z(n50090) );
  IV U59609 ( .A(n50096), .Z(n50095) );
  NAND U59610 ( .A(n50097), .B(n50098), .Z(n50052) );
  NANDN U59611 ( .A(n50099), .B(n50100), .Z(n50098) );
  NANDN U59612 ( .A(n50101), .B(n50102), .Z(n50100) );
  NANDN U59613 ( .A(n50102), .B(n50101), .Z(n50097) );
  IV U59614 ( .A(n50103), .Z(n50101) );
  XOR U59615 ( .A(n50078), .B(n50104), .Z(N60931) );
  XNOR U59616 ( .A(n50081), .B(n50080), .Z(n50104) );
  XNOR U59617 ( .A(n50092), .B(n50105), .Z(n50080) );
  XNOR U59618 ( .A(n50096), .B(n50094), .Z(n50105) );
  XOR U59619 ( .A(n50102), .B(n50106), .Z(n50094) );
  XNOR U59620 ( .A(n50099), .B(n50103), .Z(n50106) );
  AND U59621 ( .A(n50107), .B(n50108), .Z(n50103) );
  NAND U59622 ( .A(n50109), .B(n50110), .Z(n50108) );
  NAND U59623 ( .A(n50111), .B(n50112), .Z(n50107) );
  AND U59624 ( .A(n50113), .B(n50114), .Z(n50099) );
  NAND U59625 ( .A(n50115), .B(n50116), .Z(n50114) );
  NAND U59626 ( .A(n50117), .B(n50118), .Z(n50113) );
  NANDN U59627 ( .A(n50119), .B(n50120), .Z(n50102) );
  ANDN U59628 ( .B(n50121), .A(n50122), .Z(n50096) );
  XNOR U59629 ( .A(n50087), .B(n50123), .Z(n50092) );
  XNOR U59630 ( .A(n50085), .B(n50089), .Z(n50123) );
  AND U59631 ( .A(n50124), .B(n50125), .Z(n50089) );
  NAND U59632 ( .A(n50126), .B(n50127), .Z(n50125) );
  NAND U59633 ( .A(n50128), .B(n50129), .Z(n50124) );
  AND U59634 ( .A(n50130), .B(n50131), .Z(n50085) );
  NAND U59635 ( .A(n50132), .B(n50133), .Z(n50131) );
  NAND U59636 ( .A(n50134), .B(n50135), .Z(n50130) );
  AND U59637 ( .A(n50136), .B(n50137), .Z(n50087) );
  NAND U59638 ( .A(n50138), .B(n50139), .Z(n50081) );
  XNOR U59639 ( .A(n50064), .B(n50140), .Z(n50078) );
  XNOR U59640 ( .A(n50068), .B(n50066), .Z(n50140) );
  XOR U59641 ( .A(n50074), .B(n50141), .Z(n50066) );
  XNOR U59642 ( .A(n50071), .B(n50075), .Z(n50141) );
  AND U59643 ( .A(n50142), .B(n50143), .Z(n50075) );
  NAND U59644 ( .A(n50144), .B(n50145), .Z(n50143) );
  NAND U59645 ( .A(n50146), .B(n50147), .Z(n50142) );
  AND U59646 ( .A(n50148), .B(n50149), .Z(n50071) );
  NAND U59647 ( .A(n50150), .B(n50151), .Z(n50149) );
  NAND U59648 ( .A(n50152), .B(n50153), .Z(n50148) );
  NANDN U59649 ( .A(n50154), .B(n50155), .Z(n50074) );
  ANDN U59650 ( .B(n50156), .A(n50157), .Z(n50068) );
  XNOR U59651 ( .A(n50059), .B(n50158), .Z(n50064) );
  XNOR U59652 ( .A(n50057), .B(n50061), .Z(n50158) );
  AND U59653 ( .A(n50159), .B(n50160), .Z(n50061) );
  NAND U59654 ( .A(n50161), .B(n50162), .Z(n50160) );
  NAND U59655 ( .A(n50163), .B(n50164), .Z(n50159) );
  AND U59656 ( .A(n50165), .B(n50166), .Z(n50057) );
  NAND U59657 ( .A(n50167), .B(n50168), .Z(n50166) );
  NAND U59658 ( .A(n50169), .B(n50170), .Z(n50165) );
  AND U59659 ( .A(n50171), .B(n50172), .Z(n50059) );
  XOR U59660 ( .A(n50139), .B(n50138), .Z(N60930) );
  XNOR U59661 ( .A(n50156), .B(n50157), .Z(n50138) );
  XNOR U59662 ( .A(n50171), .B(n50172), .Z(n50157) );
  XOR U59663 ( .A(n50168), .B(n50167), .Z(n50172) );
  XOR U59664 ( .A(y[636]), .B(x[636]), .Z(n50167) );
  XOR U59665 ( .A(n50170), .B(n50169), .Z(n50168) );
  XOR U59666 ( .A(y[638]), .B(x[638]), .Z(n50169) );
  XOR U59667 ( .A(y[637]), .B(x[637]), .Z(n50170) );
  XOR U59668 ( .A(n50162), .B(n50161), .Z(n50171) );
  XOR U59669 ( .A(n50164), .B(n50163), .Z(n50161) );
  XOR U59670 ( .A(y[635]), .B(x[635]), .Z(n50163) );
  XOR U59671 ( .A(y[634]), .B(x[634]), .Z(n50164) );
  XOR U59672 ( .A(y[633]), .B(x[633]), .Z(n50162) );
  XNOR U59673 ( .A(n50155), .B(n50154), .Z(n50156) );
  XNOR U59674 ( .A(n50151), .B(n50150), .Z(n50154) );
  XOR U59675 ( .A(n50153), .B(n50152), .Z(n50150) );
  XOR U59676 ( .A(y[632]), .B(x[632]), .Z(n50152) );
  XOR U59677 ( .A(y[631]), .B(x[631]), .Z(n50153) );
  XOR U59678 ( .A(y[630]), .B(x[630]), .Z(n50151) );
  XOR U59679 ( .A(n50145), .B(n50144), .Z(n50155) );
  XOR U59680 ( .A(n50147), .B(n50146), .Z(n50144) );
  XOR U59681 ( .A(y[629]), .B(x[629]), .Z(n50146) );
  XOR U59682 ( .A(y[628]), .B(x[628]), .Z(n50147) );
  XOR U59683 ( .A(y[627]), .B(x[627]), .Z(n50145) );
  XNOR U59684 ( .A(n50121), .B(n50122), .Z(n50139) );
  XNOR U59685 ( .A(n50136), .B(n50137), .Z(n50122) );
  XOR U59686 ( .A(n50133), .B(n50132), .Z(n50137) );
  XOR U59687 ( .A(y[624]), .B(x[624]), .Z(n50132) );
  XOR U59688 ( .A(n50135), .B(n50134), .Z(n50133) );
  XOR U59689 ( .A(y[626]), .B(x[626]), .Z(n50134) );
  XOR U59690 ( .A(y[625]), .B(x[625]), .Z(n50135) );
  XOR U59691 ( .A(n50127), .B(n50126), .Z(n50136) );
  XOR U59692 ( .A(n50129), .B(n50128), .Z(n50126) );
  XOR U59693 ( .A(y[623]), .B(x[623]), .Z(n50128) );
  XOR U59694 ( .A(y[622]), .B(x[622]), .Z(n50129) );
  XOR U59695 ( .A(y[621]), .B(x[621]), .Z(n50127) );
  XNOR U59696 ( .A(n50120), .B(n50119), .Z(n50121) );
  XNOR U59697 ( .A(n50116), .B(n50115), .Z(n50119) );
  XOR U59698 ( .A(n50118), .B(n50117), .Z(n50115) );
  XOR U59699 ( .A(y[620]), .B(x[620]), .Z(n50117) );
  XOR U59700 ( .A(y[619]), .B(x[619]), .Z(n50118) );
  XOR U59701 ( .A(y[618]), .B(x[618]), .Z(n50116) );
  XOR U59702 ( .A(n50110), .B(n50109), .Z(n50120) );
  XOR U59703 ( .A(n50112), .B(n50111), .Z(n50109) );
  XOR U59704 ( .A(y[617]), .B(x[617]), .Z(n50111) );
  XOR U59705 ( .A(y[616]), .B(x[616]), .Z(n50112) );
  XOR U59706 ( .A(y[615]), .B(x[615]), .Z(n50110) );
  NAND U59707 ( .A(n50173), .B(n50174), .Z(N60921) );
  NAND U59708 ( .A(n50175), .B(n50176), .Z(n50174) );
  NANDN U59709 ( .A(n50177), .B(n50178), .Z(n50176) );
  NANDN U59710 ( .A(n50178), .B(n50177), .Z(n50173) );
  XOR U59711 ( .A(n50177), .B(n50179), .Z(N60920) );
  XNOR U59712 ( .A(n50175), .B(n50178), .Z(n50179) );
  NAND U59713 ( .A(n50180), .B(n50181), .Z(n50178) );
  NAND U59714 ( .A(n50182), .B(n50183), .Z(n50181) );
  NANDN U59715 ( .A(n50184), .B(n50185), .Z(n50183) );
  NANDN U59716 ( .A(n50185), .B(n50184), .Z(n50180) );
  AND U59717 ( .A(n50186), .B(n50187), .Z(n50175) );
  NAND U59718 ( .A(n50188), .B(n50189), .Z(n50187) );
  NANDN U59719 ( .A(n50190), .B(n50191), .Z(n50189) );
  NANDN U59720 ( .A(n50191), .B(n50190), .Z(n50186) );
  IV U59721 ( .A(n50192), .Z(n50191) );
  AND U59722 ( .A(n50193), .B(n50194), .Z(n50177) );
  NAND U59723 ( .A(n50195), .B(n50196), .Z(n50194) );
  NANDN U59724 ( .A(n50197), .B(n50198), .Z(n50196) );
  NANDN U59725 ( .A(n50198), .B(n50197), .Z(n50193) );
  XOR U59726 ( .A(n50190), .B(n50199), .Z(N60919) );
  XNOR U59727 ( .A(n50188), .B(n50192), .Z(n50199) );
  XOR U59728 ( .A(n50185), .B(n50200), .Z(n50192) );
  XNOR U59729 ( .A(n50182), .B(n50184), .Z(n50200) );
  AND U59730 ( .A(n50201), .B(n50202), .Z(n50184) );
  NANDN U59731 ( .A(n50203), .B(n50204), .Z(n50202) );
  OR U59732 ( .A(n50205), .B(n50206), .Z(n50204) );
  IV U59733 ( .A(n50207), .Z(n50206) );
  NANDN U59734 ( .A(n50207), .B(n50205), .Z(n50201) );
  AND U59735 ( .A(n50208), .B(n50209), .Z(n50182) );
  NAND U59736 ( .A(n50210), .B(n50211), .Z(n50209) );
  NANDN U59737 ( .A(n50212), .B(n50213), .Z(n50211) );
  NANDN U59738 ( .A(n50213), .B(n50212), .Z(n50208) );
  IV U59739 ( .A(n50214), .Z(n50213) );
  NAND U59740 ( .A(n50215), .B(n50216), .Z(n50185) );
  NANDN U59741 ( .A(n50217), .B(n50218), .Z(n50216) );
  NANDN U59742 ( .A(n50219), .B(n50220), .Z(n50218) );
  NANDN U59743 ( .A(n50220), .B(n50219), .Z(n50215) );
  IV U59744 ( .A(n50221), .Z(n50219) );
  AND U59745 ( .A(n50222), .B(n50223), .Z(n50188) );
  NAND U59746 ( .A(n50224), .B(n50225), .Z(n50223) );
  NANDN U59747 ( .A(n50226), .B(n50227), .Z(n50225) );
  NANDN U59748 ( .A(n50227), .B(n50226), .Z(n50222) );
  XOR U59749 ( .A(n50198), .B(n50228), .Z(n50190) );
  XNOR U59750 ( .A(n50195), .B(n50197), .Z(n50228) );
  AND U59751 ( .A(n50229), .B(n50230), .Z(n50197) );
  NANDN U59752 ( .A(n50231), .B(n50232), .Z(n50230) );
  OR U59753 ( .A(n50233), .B(n50234), .Z(n50232) );
  IV U59754 ( .A(n50235), .Z(n50234) );
  NANDN U59755 ( .A(n50235), .B(n50233), .Z(n50229) );
  AND U59756 ( .A(n50236), .B(n50237), .Z(n50195) );
  NAND U59757 ( .A(n50238), .B(n50239), .Z(n50237) );
  NANDN U59758 ( .A(n50240), .B(n50241), .Z(n50239) );
  NANDN U59759 ( .A(n50241), .B(n50240), .Z(n50236) );
  IV U59760 ( .A(n50242), .Z(n50241) );
  NAND U59761 ( .A(n50243), .B(n50244), .Z(n50198) );
  NANDN U59762 ( .A(n50245), .B(n50246), .Z(n50244) );
  NANDN U59763 ( .A(n50247), .B(n50248), .Z(n50246) );
  NANDN U59764 ( .A(n50248), .B(n50247), .Z(n50243) );
  IV U59765 ( .A(n50249), .Z(n50247) );
  XOR U59766 ( .A(n50224), .B(n50250), .Z(N60918) );
  XNOR U59767 ( .A(n50227), .B(n50226), .Z(n50250) );
  XNOR U59768 ( .A(n50238), .B(n50251), .Z(n50226) );
  XNOR U59769 ( .A(n50242), .B(n50240), .Z(n50251) );
  XOR U59770 ( .A(n50248), .B(n50252), .Z(n50240) );
  XNOR U59771 ( .A(n50245), .B(n50249), .Z(n50252) );
  AND U59772 ( .A(n50253), .B(n50254), .Z(n50249) );
  NAND U59773 ( .A(n50255), .B(n50256), .Z(n50254) );
  NAND U59774 ( .A(n50257), .B(n50258), .Z(n50253) );
  AND U59775 ( .A(n50259), .B(n50260), .Z(n50245) );
  NAND U59776 ( .A(n50261), .B(n50262), .Z(n50260) );
  NAND U59777 ( .A(n50263), .B(n50264), .Z(n50259) );
  NANDN U59778 ( .A(n50265), .B(n50266), .Z(n50248) );
  ANDN U59779 ( .B(n50267), .A(n50268), .Z(n50242) );
  XNOR U59780 ( .A(n50233), .B(n50269), .Z(n50238) );
  XNOR U59781 ( .A(n50231), .B(n50235), .Z(n50269) );
  AND U59782 ( .A(n50270), .B(n50271), .Z(n50235) );
  NAND U59783 ( .A(n50272), .B(n50273), .Z(n50271) );
  NAND U59784 ( .A(n50274), .B(n50275), .Z(n50270) );
  AND U59785 ( .A(n50276), .B(n50277), .Z(n50231) );
  NAND U59786 ( .A(n50278), .B(n50279), .Z(n50277) );
  NAND U59787 ( .A(n50280), .B(n50281), .Z(n50276) );
  AND U59788 ( .A(n50282), .B(n50283), .Z(n50233) );
  NAND U59789 ( .A(n50284), .B(n50285), .Z(n50227) );
  XNOR U59790 ( .A(n50210), .B(n50286), .Z(n50224) );
  XNOR U59791 ( .A(n50214), .B(n50212), .Z(n50286) );
  XOR U59792 ( .A(n50220), .B(n50287), .Z(n50212) );
  XNOR U59793 ( .A(n50217), .B(n50221), .Z(n50287) );
  AND U59794 ( .A(n50288), .B(n50289), .Z(n50221) );
  NAND U59795 ( .A(n50290), .B(n50291), .Z(n50289) );
  NAND U59796 ( .A(n50292), .B(n50293), .Z(n50288) );
  AND U59797 ( .A(n50294), .B(n50295), .Z(n50217) );
  NAND U59798 ( .A(n50296), .B(n50297), .Z(n50295) );
  NAND U59799 ( .A(n50298), .B(n50299), .Z(n50294) );
  NANDN U59800 ( .A(n50300), .B(n50301), .Z(n50220) );
  ANDN U59801 ( .B(n50302), .A(n50303), .Z(n50214) );
  XNOR U59802 ( .A(n50205), .B(n50304), .Z(n50210) );
  XNOR U59803 ( .A(n50203), .B(n50207), .Z(n50304) );
  AND U59804 ( .A(n50305), .B(n50306), .Z(n50207) );
  NAND U59805 ( .A(n50307), .B(n50308), .Z(n50306) );
  NAND U59806 ( .A(n50309), .B(n50310), .Z(n50305) );
  AND U59807 ( .A(n50311), .B(n50312), .Z(n50203) );
  NAND U59808 ( .A(n50313), .B(n50314), .Z(n50312) );
  NAND U59809 ( .A(n50315), .B(n50316), .Z(n50311) );
  AND U59810 ( .A(n50317), .B(n50318), .Z(n50205) );
  XOR U59811 ( .A(n50285), .B(n50284), .Z(N60917) );
  XNOR U59812 ( .A(n50302), .B(n50303), .Z(n50284) );
  XNOR U59813 ( .A(n50317), .B(n50318), .Z(n50303) );
  XOR U59814 ( .A(n50314), .B(n50313), .Z(n50318) );
  XOR U59815 ( .A(y[612]), .B(x[612]), .Z(n50313) );
  XOR U59816 ( .A(n50316), .B(n50315), .Z(n50314) );
  XOR U59817 ( .A(y[614]), .B(x[614]), .Z(n50315) );
  XOR U59818 ( .A(y[613]), .B(x[613]), .Z(n50316) );
  XOR U59819 ( .A(n50308), .B(n50307), .Z(n50317) );
  XOR U59820 ( .A(n50310), .B(n50309), .Z(n50307) );
  XOR U59821 ( .A(y[611]), .B(x[611]), .Z(n50309) );
  XOR U59822 ( .A(y[610]), .B(x[610]), .Z(n50310) );
  XOR U59823 ( .A(y[609]), .B(x[609]), .Z(n50308) );
  XNOR U59824 ( .A(n50301), .B(n50300), .Z(n50302) );
  XNOR U59825 ( .A(n50297), .B(n50296), .Z(n50300) );
  XOR U59826 ( .A(n50299), .B(n50298), .Z(n50296) );
  XOR U59827 ( .A(y[608]), .B(x[608]), .Z(n50298) );
  XOR U59828 ( .A(y[607]), .B(x[607]), .Z(n50299) );
  XOR U59829 ( .A(y[606]), .B(x[606]), .Z(n50297) );
  XOR U59830 ( .A(n50291), .B(n50290), .Z(n50301) );
  XOR U59831 ( .A(n50293), .B(n50292), .Z(n50290) );
  XOR U59832 ( .A(y[605]), .B(x[605]), .Z(n50292) );
  XOR U59833 ( .A(y[604]), .B(x[604]), .Z(n50293) );
  XOR U59834 ( .A(y[603]), .B(x[603]), .Z(n50291) );
  XNOR U59835 ( .A(n50267), .B(n50268), .Z(n50285) );
  XNOR U59836 ( .A(n50282), .B(n50283), .Z(n50268) );
  XOR U59837 ( .A(n50279), .B(n50278), .Z(n50283) );
  XOR U59838 ( .A(y[600]), .B(x[600]), .Z(n50278) );
  XOR U59839 ( .A(n50281), .B(n50280), .Z(n50279) );
  XOR U59840 ( .A(y[602]), .B(x[602]), .Z(n50280) );
  XOR U59841 ( .A(y[601]), .B(x[601]), .Z(n50281) );
  XOR U59842 ( .A(n50273), .B(n50272), .Z(n50282) );
  XOR U59843 ( .A(n50275), .B(n50274), .Z(n50272) );
  XOR U59844 ( .A(y[599]), .B(x[599]), .Z(n50274) );
  XOR U59845 ( .A(y[598]), .B(x[598]), .Z(n50275) );
  XOR U59846 ( .A(y[597]), .B(x[597]), .Z(n50273) );
  XNOR U59847 ( .A(n50266), .B(n50265), .Z(n50267) );
  XNOR U59848 ( .A(n50262), .B(n50261), .Z(n50265) );
  XOR U59849 ( .A(n50264), .B(n50263), .Z(n50261) );
  XOR U59850 ( .A(y[596]), .B(x[596]), .Z(n50263) );
  XOR U59851 ( .A(y[595]), .B(x[595]), .Z(n50264) );
  XOR U59852 ( .A(y[594]), .B(x[594]), .Z(n50262) );
  XOR U59853 ( .A(n50256), .B(n50255), .Z(n50266) );
  XOR U59854 ( .A(n50258), .B(n50257), .Z(n50255) );
  XOR U59855 ( .A(y[593]), .B(x[593]), .Z(n50257) );
  XOR U59856 ( .A(y[592]), .B(x[592]), .Z(n50258) );
  XOR U59857 ( .A(y[591]), .B(x[591]), .Z(n50256) );
  NAND U59858 ( .A(n50319), .B(n50320), .Z(N60908) );
  NAND U59859 ( .A(n50321), .B(n50322), .Z(n50320) );
  NANDN U59860 ( .A(n50323), .B(n50324), .Z(n50322) );
  NANDN U59861 ( .A(n50324), .B(n50323), .Z(n50319) );
  XOR U59862 ( .A(n50323), .B(n50325), .Z(N60907) );
  XNOR U59863 ( .A(n50321), .B(n50324), .Z(n50325) );
  NAND U59864 ( .A(n50326), .B(n50327), .Z(n50324) );
  NAND U59865 ( .A(n50328), .B(n50329), .Z(n50327) );
  NANDN U59866 ( .A(n50330), .B(n50331), .Z(n50329) );
  NANDN U59867 ( .A(n50331), .B(n50330), .Z(n50326) );
  AND U59868 ( .A(n50332), .B(n50333), .Z(n50321) );
  NAND U59869 ( .A(n50334), .B(n50335), .Z(n50333) );
  NANDN U59870 ( .A(n50336), .B(n50337), .Z(n50335) );
  NANDN U59871 ( .A(n50337), .B(n50336), .Z(n50332) );
  IV U59872 ( .A(n50338), .Z(n50337) );
  AND U59873 ( .A(n50339), .B(n50340), .Z(n50323) );
  NAND U59874 ( .A(n50341), .B(n50342), .Z(n50340) );
  NANDN U59875 ( .A(n50343), .B(n50344), .Z(n50342) );
  NANDN U59876 ( .A(n50344), .B(n50343), .Z(n50339) );
  XOR U59877 ( .A(n50336), .B(n50345), .Z(N60906) );
  XNOR U59878 ( .A(n50334), .B(n50338), .Z(n50345) );
  XOR U59879 ( .A(n50331), .B(n50346), .Z(n50338) );
  XNOR U59880 ( .A(n50328), .B(n50330), .Z(n50346) );
  AND U59881 ( .A(n50347), .B(n50348), .Z(n50330) );
  NANDN U59882 ( .A(n50349), .B(n50350), .Z(n50348) );
  OR U59883 ( .A(n50351), .B(n50352), .Z(n50350) );
  IV U59884 ( .A(n50353), .Z(n50352) );
  NANDN U59885 ( .A(n50353), .B(n50351), .Z(n50347) );
  AND U59886 ( .A(n50354), .B(n50355), .Z(n50328) );
  NAND U59887 ( .A(n50356), .B(n50357), .Z(n50355) );
  NANDN U59888 ( .A(n50358), .B(n50359), .Z(n50357) );
  NANDN U59889 ( .A(n50359), .B(n50358), .Z(n50354) );
  IV U59890 ( .A(n50360), .Z(n50359) );
  NAND U59891 ( .A(n50361), .B(n50362), .Z(n50331) );
  NANDN U59892 ( .A(n50363), .B(n50364), .Z(n50362) );
  NANDN U59893 ( .A(n50365), .B(n50366), .Z(n50364) );
  NANDN U59894 ( .A(n50366), .B(n50365), .Z(n50361) );
  IV U59895 ( .A(n50367), .Z(n50365) );
  AND U59896 ( .A(n50368), .B(n50369), .Z(n50334) );
  NAND U59897 ( .A(n50370), .B(n50371), .Z(n50369) );
  NANDN U59898 ( .A(n50372), .B(n50373), .Z(n50371) );
  NANDN U59899 ( .A(n50373), .B(n50372), .Z(n50368) );
  XOR U59900 ( .A(n50344), .B(n50374), .Z(n50336) );
  XNOR U59901 ( .A(n50341), .B(n50343), .Z(n50374) );
  AND U59902 ( .A(n50375), .B(n50376), .Z(n50343) );
  NANDN U59903 ( .A(n50377), .B(n50378), .Z(n50376) );
  OR U59904 ( .A(n50379), .B(n50380), .Z(n50378) );
  IV U59905 ( .A(n50381), .Z(n50380) );
  NANDN U59906 ( .A(n50381), .B(n50379), .Z(n50375) );
  AND U59907 ( .A(n50382), .B(n50383), .Z(n50341) );
  NAND U59908 ( .A(n50384), .B(n50385), .Z(n50383) );
  NANDN U59909 ( .A(n50386), .B(n50387), .Z(n50385) );
  NANDN U59910 ( .A(n50387), .B(n50386), .Z(n50382) );
  IV U59911 ( .A(n50388), .Z(n50387) );
  NAND U59912 ( .A(n50389), .B(n50390), .Z(n50344) );
  NANDN U59913 ( .A(n50391), .B(n50392), .Z(n50390) );
  NANDN U59914 ( .A(n50393), .B(n50394), .Z(n50392) );
  NANDN U59915 ( .A(n50394), .B(n50393), .Z(n50389) );
  IV U59916 ( .A(n50395), .Z(n50393) );
  XOR U59917 ( .A(n50370), .B(n50396), .Z(N60905) );
  XNOR U59918 ( .A(n50373), .B(n50372), .Z(n50396) );
  XNOR U59919 ( .A(n50384), .B(n50397), .Z(n50372) );
  XNOR U59920 ( .A(n50388), .B(n50386), .Z(n50397) );
  XOR U59921 ( .A(n50394), .B(n50398), .Z(n50386) );
  XNOR U59922 ( .A(n50391), .B(n50395), .Z(n50398) );
  AND U59923 ( .A(n50399), .B(n50400), .Z(n50395) );
  NAND U59924 ( .A(n50401), .B(n50402), .Z(n50400) );
  NAND U59925 ( .A(n50403), .B(n50404), .Z(n50399) );
  AND U59926 ( .A(n50405), .B(n50406), .Z(n50391) );
  NAND U59927 ( .A(n50407), .B(n50408), .Z(n50406) );
  NAND U59928 ( .A(n50409), .B(n50410), .Z(n50405) );
  NANDN U59929 ( .A(n50411), .B(n50412), .Z(n50394) );
  ANDN U59930 ( .B(n50413), .A(n50414), .Z(n50388) );
  XNOR U59931 ( .A(n50379), .B(n50415), .Z(n50384) );
  XNOR U59932 ( .A(n50377), .B(n50381), .Z(n50415) );
  AND U59933 ( .A(n50416), .B(n50417), .Z(n50381) );
  NAND U59934 ( .A(n50418), .B(n50419), .Z(n50417) );
  NAND U59935 ( .A(n50420), .B(n50421), .Z(n50416) );
  AND U59936 ( .A(n50422), .B(n50423), .Z(n50377) );
  NAND U59937 ( .A(n50424), .B(n50425), .Z(n50423) );
  NAND U59938 ( .A(n50426), .B(n50427), .Z(n50422) );
  AND U59939 ( .A(n50428), .B(n50429), .Z(n50379) );
  NAND U59940 ( .A(n50430), .B(n50431), .Z(n50373) );
  XNOR U59941 ( .A(n50356), .B(n50432), .Z(n50370) );
  XNOR U59942 ( .A(n50360), .B(n50358), .Z(n50432) );
  XOR U59943 ( .A(n50366), .B(n50433), .Z(n50358) );
  XNOR U59944 ( .A(n50363), .B(n50367), .Z(n50433) );
  AND U59945 ( .A(n50434), .B(n50435), .Z(n50367) );
  NAND U59946 ( .A(n50436), .B(n50437), .Z(n50435) );
  NAND U59947 ( .A(n50438), .B(n50439), .Z(n50434) );
  AND U59948 ( .A(n50440), .B(n50441), .Z(n50363) );
  NAND U59949 ( .A(n50442), .B(n50443), .Z(n50441) );
  NAND U59950 ( .A(n50444), .B(n50445), .Z(n50440) );
  NANDN U59951 ( .A(n50446), .B(n50447), .Z(n50366) );
  ANDN U59952 ( .B(n50448), .A(n50449), .Z(n50360) );
  XNOR U59953 ( .A(n50351), .B(n50450), .Z(n50356) );
  XNOR U59954 ( .A(n50349), .B(n50353), .Z(n50450) );
  AND U59955 ( .A(n50451), .B(n50452), .Z(n50353) );
  NAND U59956 ( .A(n50453), .B(n50454), .Z(n50452) );
  NAND U59957 ( .A(n50455), .B(n50456), .Z(n50451) );
  AND U59958 ( .A(n50457), .B(n50458), .Z(n50349) );
  NAND U59959 ( .A(n50459), .B(n50460), .Z(n50458) );
  NAND U59960 ( .A(n50461), .B(n50462), .Z(n50457) );
  AND U59961 ( .A(n50463), .B(n50464), .Z(n50351) );
  XOR U59962 ( .A(n50431), .B(n50430), .Z(N60904) );
  XNOR U59963 ( .A(n50448), .B(n50449), .Z(n50430) );
  XNOR U59964 ( .A(n50463), .B(n50464), .Z(n50449) );
  XOR U59965 ( .A(n50460), .B(n50459), .Z(n50464) );
  XOR U59966 ( .A(y[588]), .B(x[588]), .Z(n50459) );
  XOR U59967 ( .A(n50462), .B(n50461), .Z(n50460) );
  XOR U59968 ( .A(y[590]), .B(x[590]), .Z(n50461) );
  XOR U59969 ( .A(y[589]), .B(x[589]), .Z(n50462) );
  XOR U59970 ( .A(n50454), .B(n50453), .Z(n50463) );
  XOR U59971 ( .A(n50456), .B(n50455), .Z(n50453) );
  XOR U59972 ( .A(y[587]), .B(x[587]), .Z(n50455) );
  XOR U59973 ( .A(y[586]), .B(x[586]), .Z(n50456) );
  XOR U59974 ( .A(y[585]), .B(x[585]), .Z(n50454) );
  XNOR U59975 ( .A(n50447), .B(n50446), .Z(n50448) );
  XNOR U59976 ( .A(n50443), .B(n50442), .Z(n50446) );
  XOR U59977 ( .A(n50445), .B(n50444), .Z(n50442) );
  XOR U59978 ( .A(y[584]), .B(x[584]), .Z(n50444) );
  XOR U59979 ( .A(y[583]), .B(x[583]), .Z(n50445) );
  XOR U59980 ( .A(y[582]), .B(x[582]), .Z(n50443) );
  XOR U59981 ( .A(n50437), .B(n50436), .Z(n50447) );
  XOR U59982 ( .A(n50439), .B(n50438), .Z(n50436) );
  XOR U59983 ( .A(y[581]), .B(x[581]), .Z(n50438) );
  XOR U59984 ( .A(y[580]), .B(x[580]), .Z(n50439) );
  XOR U59985 ( .A(y[579]), .B(x[579]), .Z(n50437) );
  XNOR U59986 ( .A(n50413), .B(n50414), .Z(n50431) );
  XNOR U59987 ( .A(n50428), .B(n50429), .Z(n50414) );
  XOR U59988 ( .A(n50425), .B(n50424), .Z(n50429) );
  XOR U59989 ( .A(y[576]), .B(x[576]), .Z(n50424) );
  XOR U59990 ( .A(n50427), .B(n50426), .Z(n50425) );
  XOR U59991 ( .A(y[578]), .B(x[578]), .Z(n50426) );
  XOR U59992 ( .A(y[577]), .B(x[577]), .Z(n50427) );
  XOR U59993 ( .A(n50419), .B(n50418), .Z(n50428) );
  XOR U59994 ( .A(n50421), .B(n50420), .Z(n50418) );
  XOR U59995 ( .A(y[575]), .B(x[575]), .Z(n50420) );
  XOR U59996 ( .A(y[574]), .B(x[574]), .Z(n50421) );
  XOR U59997 ( .A(y[573]), .B(x[573]), .Z(n50419) );
  XNOR U59998 ( .A(n50412), .B(n50411), .Z(n50413) );
  XNOR U59999 ( .A(n50408), .B(n50407), .Z(n50411) );
  XOR U60000 ( .A(n50410), .B(n50409), .Z(n50407) );
  XOR U60001 ( .A(y[572]), .B(x[572]), .Z(n50409) );
  XOR U60002 ( .A(y[571]), .B(x[571]), .Z(n50410) );
  XOR U60003 ( .A(y[570]), .B(x[570]), .Z(n50408) );
  XOR U60004 ( .A(n50402), .B(n50401), .Z(n50412) );
  XOR U60005 ( .A(n50404), .B(n50403), .Z(n50401) );
  XOR U60006 ( .A(y[569]), .B(x[569]), .Z(n50403) );
  XOR U60007 ( .A(y[568]), .B(x[568]), .Z(n50404) );
  XOR U60008 ( .A(y[567]), .B(x[567]), .Z(n50402) );
  NAND U60009 ( .A(n50465), .B(n50466), .Z(N60895) );
  NAND U60010 ( .A(n50467), .B(n50468), .Z(n50466) );
  NANDN U60011 ( .A(n50469), .B(n50470), .Z(n50468) );
  NANDN U60012 ( .A(n50470), .B(n50469), .Z(n50465) );
  XOR U60013 ( .A(n50469), .B(n50471), .Z(N60894) );
  XNOR U60014 ( .A(n50467), .B(n50470), .Z(n50471) );
  NAND U60015 ( .A(n50472), .B(n50473), .Z(n50470) );
  NAND U60016 ( .A(n50474), .B(n50475), .Z(n50473) );
  NANDN U60017 ( .A(n50476), .B(n50477), .Z(n50475) );
  NANDN U60018 ( .A(n50477), .B(n50476), .Z(n50472) );
  AND U60019 ( .A(n50478), .B(n50479), .Z(n50467) );
  NAND U60020 ( .A(n50480), .B(n50481), .Z(n50479) );
  NANDN U60021 ( .A(n50482), .B(n50483), .Z(n50481) );
  NANDN U60022 ( .A(n50483), .B(n50482), .Z(n50478) );
  IV U60023 ( .A(n50484), .Z(n50483) );
  AND U60024 ( .A(n50485), .B(n50486), .Z(n50469) );
  NAND U60025 ( .A(n50487), .B(n50488), .Z(n50486) );
  NANDN U60026 ( .A(n50489), .B(n50490), .Z(n50488) );
  NANDN U60027 ( .A(n50490), .B(n50489), .Z(n50485) );
  XOR U60028 ( .A(n50482), .B(n50491), .Z(N60893) );
  XNOR U60029 ( .A(n50480), .B(n50484), .Z(n50491) );
  XOR U60030 ( .A(n50477), .B(n50492), .Z(n50484) );
  XNOR U60031 ( .A(n50474), .B(n50476), .Z(n50492) );
  AND U60032 ( .A(n50493), .B(n50494), .Z(n50476) );
  NANDN U60033 ( .A(n50495), .B(n50496), .Z(n50494) );
  OR U60034 ( .A(n50497), .B(n50498), .Z(n50496) );
  IV U60035 ( .A(n50499), .Z(n50498) );
  NANDN U60036 ( .A(n50499), .B(n50497), .Z(n50493) );
  AND U60037 ( .A(n50500), .B(n50501), .Z(n50474) );
  NAND U60038 ( .A(n50502), .B(n50503), .Z(n50501) );
  NANDN U60039 ( .A(n50504), .B(n50505), .Z(n50503) );
  NANDN U60040 ( .A(n50505), .B(n50504), .Z(n50500) );
  IV U60041 ( .A(n50506), .Z(n50505) );
  NAND U60042 ( .A(n50507), .B(n50508), .Z(n50477) );
  NANDN U60043 ( .A(n50509), .B(n50510), .Z(n50508) );
  NANDN U60044 ( .A(n50511), .B(n50512), .Z(n50510) );
  NANDN U60045 ( .A(n50512), .B(n50511), .Z(n50507) );
  IV U60046 ( .A(n50513), .Z(n50511) );
  AND U60047 ( .A(n50514), .B(n50515), .Z(n50480) );
  NAND U60048 ( .A(n50516), .B(n50517), .Z(n50515) );
  NANDN U60049 ( .A(n50518), .B(n50519), .Z(n50517) );
  NANDN U60050 ( .A(n50519), .B(n50518), .Z(n50514) );
  XOR U60051 ( .A(n50490), .B(n50520), .Z(n50482) );
  XNOR U60052 ( .A(n50487), .B(n50489), .Z(n50520) );
  AND U60053 ( .A(n50521), .B(n50522), .Z(n50489) );
  NANDN U60054 ( .A(n50523), .B(n50524), .Z(n50522) );
  OR U60055 ( .A(n50525), .B(n50526), .Z(n50524) );
  IV U60056 ( .A(n50527), .Z(n50526) );
  NANDN U60057 ( .A(n50527), .B(n50525), .Z(n50521) );
  AND U60058 ( .A(n50528), .B(n50529), .Z(n50487) );
  NAND U60059 ( .A(n50530), .B(n50531), .Z(n50529) );
  NANDN U60060 ( .A(n50532), .B(n50533), .Z(n50531) );
  NANDN U60061 ( .A(n50533), .B(n50532), .Z(n50528) );
  IV U60062 ( .A(n50534), .Z(n50533) );
  NAND U60063 ( .A(n50535), .B(n50536), .Z(n50490) );
  NANDN U60064 ( .A(n50537), .B(n50538), .Z(n50536) );
  NANDN U60065 ( .A(n50539), .B(n50540), .Z(n50538) );
  NANDN U60066 ( .A(n50540), .B(n50539), .Z(n50535) );
  IV U60067 ( .A(n50541), .Z(n50539) );
  XOR U60068 ( .A(n50516), .B(n50542), .Z(N60892) );
  XNOR U60069 ( .A(n50519), .B(n50518), .Z(n50542) );
  XNOR U60070 ( .A(n50530), .B(n50543), .Z(n50518) );
  XNOR U60071 ( .A(n50534), .B(n50532), .Z(n50543) );
  XOR U60072 ( .A(n50540), .B(n50544), .Z(n50532) );
  XNOR U60073 ( .A(n50537), .B(n50541), .Z(n50544) );
  AND U60074 ( .A(n50545), .B(n50546), .Z(n50541) );
  NAND U60075 ( .A(n50547), .B(n50548), .Z(n50546) );
  NAND U60076 ( .A(n50549), .B(n50550), .Z(n50545) );
  AND U60077 ( .A(n50551), .B(n50552), .Z(n50537) );
  NAND U60078 ( .A(n50553), .B(n50554), .Z(n50552) );
  NAND U60079 ( .A(n50555), .B(n50556), .Z(n50551) );
  NANDN U60080 ( .A(n50557), .B(n50558), .Z(n50540) );
  ANDN U60081 ( .B(n50559), .A(n50560), .Z(n50534) );
  XNOR U60082 ( .A(n50525), .B(n50561), .Z(n50530) );
  XNOR U60083 ( .A(n50523), .B(n50527), .Z(n50561) );
  AND U60084 ( .A(n50562), .B(n50563), .Z(n50527) );
  NAND U60085 ( .A(n50564), .B(n50565), .Z(n50563) );
  NAND U60086 ( .A(n50566), .B(n50567), .Z(n50562) );
  AND U60087 ( .A(n50568), .B(n50569), .Z(n50523) );
  NAND U60088 ( .A(n50570), .B(n50571), .Z(n50569) );
  NAND U60089 ( .A(n50572), .B(n50573), .Z(n50568) );
  AND U60090 ( .A(n50574), .B(n50575), .Z(n50525) );
  NAND U60091 ( .A(n50576), .B(n50577), .Z(n50519) );
  XNOR U60092 ( .A(n50502), .B(n50578), .Z(n50516) );
  XNOR U60093 ( .A(n50506), .B(n50504), .Z(n50578) );
  XOR U60094 ( .A(n50512), .B(n50579), .Z(n50504) );
  XNOR U60095 ( .A(n50509), .B(n50513), .Z(n50579) );
  AND U60096 ( .A(n50580), .B(n50581), .Z(n50513) );
  NAND U60097 ( .A(n50582), .B(n50583), .Z(n50581) );
  NAND U60098 ( .A(n50584), .B(n50585), .Z(n50580) );
  AND U60099 ( .A(n50586), .B(n50587), .Z(n50509) );
  NAND U60100 ( .A(n50588), .B(n50589), .Z(n50587) );
  NAND U60101 ( .A(n50590), .B(n50591), .Z(n50586) );
  NANDN U60102 ( .A(n50592), .B(n50593), .Z(n50512) );
  ANDN U60103 ( .B(n50594), .A(n50595), .Z(n50506) );
  XNOR U60104 ( .A(n50497), .B(n50596), .Z(n50502) );
  XNOR U60105 ( .A(n50495), .B(n50499), .Z(n50596) );
  AND U60106 ( .A(n50597), .B(n50598), .Z(n50499) );
  NAND U60107 ( .A(n50599), .B(n50600), .Z(n50598) );
  NAND U60108 ( .A(n50601), .B(n50602), .Z(n50597) );
  AND U60109 ( .A(n50603), .B(n50604), .Z(n50495) );
  NAND U60110 ( .A(n50605), .B(n50606), .Z(n50604) );
  NAND U60111 ( .A(n50607), .B(n50608), .Z(n50603) );
  AND U60112 ( .A(n50609), .B(n50610), .Z(n50497) );
  XOR U60113 ( .A(n50577), .B(n50576), .Z(N60891) );
  XNOR U60114 ( .A(n50594), .B(n50595), .Z(n50576) );
  XNOR U60115 ( .A(n50609), .B(n50610), .Z(n50595) );
  XOR U60116 ( .A(n50606), .B(n50605), .Z(n50610) );
  XOR U60117 ( .A(y[564]), .B(x[564]), .Z(n50605) );
  XOR U60118 ( .A(n50608), .B(n50607), .Z(n50606) );
  XOR U60119 ( .A(y[566]), .B(x[566]), .Z(n50607) );
  XOR U60120 ( .A(y[565]), .B(x[565]), .Z(n50608) );
  XOR U60121 ( .A(n50600), .B(n50599), .Z(n50609) );
  XOR U60122 ( .A(n50602), .B(n50601), .Z(n50599) );
  XOR U60123 ( .A(y[563]), .B(x[563]), .Z(n50601) );
  XOR U60124 ( .A(y[562]), .B(x[562]), .Z(n50602) );
  XOR U60125 ( .A(y[561]), .B(x[561]), .Z(n50600) );
  XNOR U60126 ( .A(n50593), .B(n50592), .Z(n50594) );
  XNOR U60127 ( .A(n50589), .B(n50588), .Z(n50592) );
  XOR U60128 ( .A(n50591), .B(n50590), .Z(n50588) );
  XOR U60129 ( .A(y[560]), .B(x[560]), .Z(n50590) );
  XOR U60130 ( .A(y[559]), .B(x[559]), .Z(n50591) );
  XOR U60131 ( .A(y[558]), .B(x[558]), .Z(n50589) );
  XOR U60132 ( .A(n50583), .B(n50582), .Z(n50593) );
  XOR U60133 ( .A(n50585), .B(n50584), .Z(n50582) );
  XOR U60134 ( .A(y[557]), .B(x[557]), .Z(n50584) );
  XOR U60135 ( .A(y[556]), .B(x[556]), .Z(n50585) );
  XOR U60136 ( .A(y[555]), .B(x[555]), .Z(n50583) );
  XNOR U60137 ( .A(n50559), .B(n50560), .Z(n50577) );
  XNOR U60138 ( .A(n50574), .B(n50575), .Z(n50560) );
  XOR U60139 ( .A(n50571), .B(n50570), .Z(n50575) );
  XOR U60140 ( .A(y[552]), .B(x[552]), .Z(n50570) );
  XOR U60141 ( .A(n50573), .B(n50572), .Z(n50571) );
  XOR U60142 ( .A(y[554]), .B(x[554]), .Z(n50572) );
  XOR U60143 ( .A(y[553]), .B(x[553]), .Z(n50573) );
  XOR U60144 ( .A(n50565), .B(n50564), .Z(n50574) );
  XOR U60145 ( .A(n50567), .B(n50566), .Z(n50564) );
  XOR U60146 ( .A(y[551]), .B(x[551]), .Z(n50566) );
  XOR U60147 ( .A(y[550]), .B(x[550]), .Z(n50567) );
  XOR U60148 ( .A(y[549]), .B(x[549]), .Z(n50565) );
  XNOR U60149 ( .A(n50558), .B(n50557), .Z(n50559) );
  XNOR U60150 ( .A(n50554), .B(n50553), .Z(n50557) );
  XOR U60151 ( .A(n50556), .B(n50555), .Z(n50553) );
  XOR U60152 ( .A(y[548]), .B(x[548]), .Z(n50555) );
  XOR U60153 ( .A(y[547]), .B(x[547]), .Z(n50556) );
  XOR U60154 ( .A(y[546]), .B(x[546]), .Z(n50554) );
  XOR U60155 ( .A(n50548), .B(n50547), .Z(n50558) );
  XOR U60156 ( .A(n50550), .B(n50549), .Z(n50547) );
  XOR U60157 ( .A(y[545]), .B(x[545]), .Z(n50549) );
  XOR U60158 ( .A(y[544]), .B(x[544]), .Z(n50550) );
  XOR U60159 ( .A(y[543]), .B(x[543]), .Z(n50548) );
  NAND U60160 ( .A(n50611), .B(n50612), .Z(N60882) );
  NAND U60161 ( .A(n50613), .B(n50614), .Z(n50612) );
  NANDN U60162 ( .A(n50615), .B(n50616), .Z(n50614) );
  NANDN U60163 ( .A(n50616), .B(n50615), .Z(n50611) );
  XOR U60164 ( .A(n50615), .B(n50617), .Z(N60881) );
  XNOR U60165 ( .A(n50613), .B(n50616), .Z(n50617) );
  NAND U60166 ( .A(n50618), .B(n50619), .Z(n50616) );
  NAND U60167 ( .A(n50620), .B(n50621), .Z(n50619) );
  NANDN U60168 ( .A(n50622), .B(n50623), .Z(n50621) );
  NANDN U60169 ( .A(n50623), .B(n50622), .Z(n50618) );
  AND U60170 ( .A(n50624), .B(n50625), .Z(n50613) );
  NAND U60171 ( .A(n50626), .B(n50627), .Z(n50625) );
  NANDN U60172 ( .A(n50628), .B(n50629), .Z(n50627) );
  NANDN U60173 ( .A(n50629), .B(n50628), .Z(n50624) );
  IV U60174 ( .A(n50630), .Z(n50629) );
  AND U60175 ( .A(n50631), .B(n50632), .Z(n50615) );
  NAND U60176 ( .A(n50633), .B(n50634), .Z(n50632) );
  NANDN U60177 ( .A(n50635), .B(n50636), .Z(n50634) );
  NANDN U60178 ( .A(n50636), .B(n50635), .Z(n50631) );
  XOR U60179 ( .A(n50628), .B(n50637), .Z(N60880) );
  XNOR U60180 ( .A(n50626), .B(n50630), .Z(n50637) );
  XOR U60181 ( .A(n50623), .B(n50638), .Z(n50630) );
  XNOR U60182 ( .A(n50620), .B(n50622), .Z(n50638) );
  AND U60183 ( .A(n50639), .B(n50640), .Z(n50622) );
  NANDN U60184 ( .A(n50641), .B(n50642), .Z(n50640) );
  OR U60185 ( .A(n50643), .B(n50644), .Z(n50642) );
  IV U60186 ( .A(n50645), .Z(n50644) );
  NANDN U60187 ( .A(n50645), .B(n50643), .Z(n50639) );
  AND U60188 ( .A(n50646), .B(n50647), .Z(n50620) );
  NAND U60189 ( .A(n50648), .B(n50649), .Z(n50647) );
  NANDN U60190 ( .A(n50650), .B(n50651), .Z(n50649) );
  NANDN U60191 ( .A(n50651), .B(n50650), .Z(n50646) );
  IV U60192 ( .A(n50652), .Z(n50651) );
  NAND U60193 ( .A(n50653), .B(n50654), .Z(n50623) );
  NANDN U60194 ( .A(n50655), .B(n50656), .Z(n50654) );
  NANDN U60195 ( .A(n50657), .B(n50658), .Z(n50656) );
  NANDN U60196 ( .A(n50658), .B(n50657), .Z(n50653) );
  IV U60197 ( .A(n50659), .Z(n50657) );
  AND U60198 ( .A(n50660), .B(n50661), .Z(n50626) );
  NAND U60199 ( .A(n50662), .B(n50663), .Z(n50661) );
  NANDN U60200 ( .A(n50664), .B(n50665), .Z(n50663) );
  NANDN U60201 ( .A(n50665), .B(n50664), .Z(n50660) );
  XOR U60202 ( .A(n50636), .B(n50666), .Z(n50628) );
  XNOR U60203 ( .A(n50633), .B(n50635), .Z(n50666) );
  AND U60204 ( .A(n50667), .B(n50668), .Z(n50635) );
  NANDN U60205 ( .A(n50669), .B(n50670), .Z(n50668) );
  OR U60206 ( .A(n50671), .B(n50672), .Z(n50670) );
  IV U60207 ( .A(n50673), .Z(n50672) );
  NANDN U60208 ( .A(n50673), .B(n50671), .Z(n50667) );
  AND U60209 ( .A(n50674), .B(n50675), .Z(n50633) );
  NAND U60210 ( .A(n50676), .B(n50677), .Z(n50675) );
  NANDN U60211 ( .A(n50678), .B(n50679), .Z(n50677) );
  NANDN U60212 ( .A(n50679), .B(n50678), .Z(n50674) );
  IV U60213 ( .A(n50680), .Z(n50679) );
  NAND U60214 ( .A(n50681), .B(n50682), .Z(n50636) );
  NANDN U60215 ( .A(n50683), .B(n50684), .Z(n50682) );
  NANDN U60216 ( .A(n50685), .B(n50686), .Z(n50684) );
  NANDN U60217 ( .A(n50686), .B(n50685), .Z(n50681) );
  IV U60218 ( .A(n50687), .Z(n50685) );
  XOR U60219 ( .A(n50662), .B(n50688), .Z(N60879) );
  XNOR U60220 ( .A(n50665), .B(n50664), .Z(n50688) );
  XNOR U60221 ( .A(n50676), .B(n50689), .Z(n50664) );
  XNOR U60222 ( .A(n50680), .B(n50678), .Z(n50689) );
  XOR U60223 ( .A(n50686), .B(n50690), .Z(n50678) );
  XNOR U60224 ( .A(n50683), .B(n50687), .Z(n50690) );
  AND U60225 ( .A(n50691), .B(n50692), .Z(n50687) );
  NAND U60226 ( .A(n50693), .B(n50694), .Z(n50692) );
  NAND U60227 ( .A(n50695), .B(n50696), .Z(n50691) );
  AND U60228 ( .A(n50697), .B(n50698), .Z(n50683) );
  NAND U60229 ( .A(n50699), .B(n50700), .Z(n50698) );
  NAND U60230 ( .A(n50701), .B(n50702), .Z(n50697) );
  NANDN U60231 ( .A(n50703), .B(n50704), .Z(n50686) );
  ANDN U60232 ( .B(n50705), .A(n50706), .Z(n50680) );
  XNOR U60233 ( .A(n50671), .B(n50707), .Z(n50676) );
  XNOR U60234 ( .A(n50669), .B(n50673), .Z(n50707) );
  AND U60235 ( .A(n50708), .B(n50709), .Z(n50673) );
  NAND U60236 ( .A(n50710), .B(n50711), .Z(n50709) );
  NAND U60237 ( .A(n50712), .B(n50713), .Z(n50708) );
  AND U60238 ( .A(n50714), .B(n50715), .Z(n50669) );
  NAND U60239 ( .A(n50716), .B(n50717), .Z(n50715) );
  NAND U60240 ( .A(n50718), .B(n50719), .Z(n50714) );
  AND U60241 ( .A(n50720), .B(n50721), .Z(n50671) );
  NAND U60242 ( .A(n50722), .B(n50723), .Z(n50665) );
  XNOR U60243 ( .A(n50648), .B(n50724), .Z(n50662) );
  XNOR U60244 ( .A(n50652), .B(n50650), .Z(n50724) );
  XOR U60245 ( .A(n50658), .B(n50725), .Z(n50650) );
  XNOR U60246 ( .A(n50655), .B(n50659), .Z(n50725) );
  AND U60247 ( .A(n50726), .B(n50727), .Z(n50659) );
  NAND U60248 ( .A(n50728), .B(n50729), .Z(n50727) );
  NAND U60249 ( .A(n50730), .B(n50731), .Z(n50726) );
  AND U60250 ( .A(n50732), .B(n50733), .Z(n50655) );
  NAND U60251 ( .A(n50734), .B(n50735), .Z(n50733) );
  NAND U60252 ( .A(n50736), .B(n50737), .Z(n50732) );
  NANDN U60253 ( .A(n50738), .B(n50739), .Z(n50658) );
  ANDN U60254 ( .B(n50740), .A(n50741), .Z(n50652) );
  XNOR U60255 ( .A(n50643), .B(n50742), .Z(n50648) );
  XNOR U60256 ( .A(n50641), .B(n50645), .Z(n50742) );
  AND U60257 ( .A(n50743), .B(n50744), .Z(n50645) );
  NAND U60258 ( .A(n50745), .B(n50746), .Z(n50744) );
  NAND U60259 ( .A(n50747), .B(n50748), .Z(n50743) );
  AND U60260 ( .A(n50749), .B(n50750), .Z(n50641) );
  NAND U60261 ( .A(n50751), .B(n50752), .Z(n50750) );
  NAND U60262 ( .A(n50753), .B(n50754), .Z(n50749) );
  AND U60263 ( .A(n50755), .B(n50756), .Z(n50643) );
  XOR U60264 ( .A(n50723), .B(n50722), .Z(N60878) );
  XNOR U60265 ( .A(n50740), .B(n50741), .Z(n50722) );
  XNOR U60266 ( .A(n50755), .B(n50756), .Z(n50741) );
  XOR U60267 ( .A(n50752), .B(n50751), .Z(n50756) );
  XOR U60268 ( .A(y[540]), .B(x[540]), .Z(n50751) );
  XOR U60269 ( .A(n50754), .B(n50753), .Z(n50752) );
  XOR U60270 ( .A(y[542]), .B(x[542]), .Z(n50753) );
  XOR U60271 ( .A(y[541]), .B(x[541]), .Z(n50754) );
  XOR U60272 ( .A(n50746), .B(n50745), .Z(n50755) );
  XOR U60273 ( .A(n50748), .B(n50747), .Z(n50745) );
  XOR U60274 ( .A(y[539]), .B(x[539]), .Z(n50747) );
  XOR U60275 ( .A(y[538]), .B(x[538]), .Z(n50748) );
  XOR U60276 ( .A(y[537]), .B(x[537]), .Z(n50746) );
  XNOR U60277 ( .A(n50739), .B(n50738), .Z(n50740) );
  XNOR U60278 ( .A(n50735), .B(n50734), .Z(n50738) );
  XOR U60279 ( .A(n50737), .B(n50736), .Z(n50734) );
  XOR U60280 ( .A(y[536]), .B(x[536]), .Z(n50736) );
  XOR U60281 ( .A(y[535]), .B(x[535]), .Z(n50737) );
  XOR U60282 ( .A(y[534]), .B(x[534]), .Z(n50735) );
  XOR U60283 ( .A(n50729), .B(n50728), .Z(n50739) );
  XOR U60284 ( .A(n50731), .B(n50730), .Z(n50728) );
  XOR U60285 ( .A(y[533]), .B(x[533]), .Z(n50730) );
  XOR U60286 ( .A(y[532]), .B(x[532]), .Z(n50731) );
  XOR U60287 ( .A(y[531]), .B(x[531]), .Z(n50729) );
  XNOR U60288 ( .A(n50705), .B(n50706), .Z(n50723) );
  XNOR U60289 ( .A(n50720), .B(n50721), .Z(n50706) );
  XOR U60290 ( .A(n50717), .B(n50716), .Z(n50721) );
  XOR U60291 ( .A(y[528]), .B(x[528]), .Z(n50716) );
  XOR U60292 ( .A(n50719), .B(n50718), .Z(n50717) );
  XOR U60293 ( .A(y[530]), .B(x[530]), .Z(n50718) );
  XOR U60294 ( .A(y[529]), .B(x[529]), .Z(n50719) );
  XOR U60295 ( .A(n50711), .B(n50710), .Z(n50720) );
  XOR U60296 ( .A(n50713), .B(n50712), .Z(n50710) );
  XOR U60297 ( .A(y[527]), .B(x[527]), .Z(n50712) );
  XOR U60298 ( .A(y[526]), .B(x[526]), .Z(n50713) );
  XOR U60299 ( .A(y[525]), .B(x[525]), .Z(n50711) );
  XNOR U60300 ( .A(n50704), .B(n50703), .Z(n50705) );
  XNOR U60301 ( .A(n50700), .B(n50699), .Z(n50703) );
  XOR U60302 ( .A(n50702), .B(n50701), .Z(n50699) );
  XOR U60303 ( .A(y[524]), .B(x[524]), .Z(n50701) );
  XOR U60304 ( .A(y[523]), .B(x[523]), .Z(n50702) );
  XOR U60305 ( .A(y[522]), .B(x[522]), .Z(n50700) );
  XOR U60306 ( .A(n50694), .B(n50693), .Z(n50704) );
  XOR U60307 ( .A(n50696), .B(n50695), .Z(n50693) );
  XOR U60308 ( .A(y[521]), .B(x[521]), .Z(n50695) );
  XOR U60309 ( .A(y[520]), .B(x[520]), .Z(n50696) );
  XOR U60310 ( .A(y[519]), .B(x[519]), .Z(n50694) );
  NAND U60311 ( .A(n50757), .B(n50758), .Z(N60869) );
  NAND U60312 ( .A(n50759), .B(n50760), .Z(n50758) );
  NANDN U60313 ( .A(n50761), .B(n50762), .Z(n50760) );
  NANDN U60314 ( .A(n50762), .B(n50761), .Z(n50757) );
  XOR U60315 ( .A(n50761), .B(n50763), .Z(N60868) );
  XNOR U60316 ( .A(n50759), .B(n50762), .Z(n50763) );
  NAND U60317 ( .A(n50764), .B(n50765), .Z(n50762) );
  NAND U60318 ( .A(n50766), .B(n50767), .Z(n50765) );
  NANDN U60319 ( .A(n50768), .B(n50769), .Z(n50767) );
  NANDN U60320 ( .A(n50769), .B(n50768), .Z(n50764) );
  AND U60321 ( .A(n50770), .B(n50771), .Z(n50759) );
  NAND U60322 ( .A(n50772), .B(n50773), .Z(n50771) );
  NANDN U60323 ( .A(n50774), .B(n50775), .Z(n50773) );
  NANDN U60324 ( .A(n50775), .B(n50774), .Z(n50770) );
  IV U60325 ( .A(n50776), .Z(n50775) );
  AND U60326 ( .A(n50777), .B(n50778), .Z(n50761) );
  NAND U60327 ( .A(n50779), .B(n50780), .Z(n50778) );
  NANDN U60328 ( .A(n50781), .B(n50782), .Z(n50780) );
  NANDN U60329 ( .A(n50782), .B(n50781), .Z(n50777) );
  XOR U60330 ( .A(n50774), .B(n50783), .Z(N60867) );
  XNOR U60331 ( .A(n50772), .B(n50776), .Z(n50783) );
  XOR U60332 ( .A(n50769), .B(n50784), .Z(n50776) );
  XNOR U60333 ( .A(n50766), .B(n50768), .Z(n50784) );
  AND U60334 ( .A(n50785), .B(n50786), .Z(n50768) );
  NANDN U60335 ( .A(n50787), .B(n50788), .Z(n50786) );
  OR U60336 ( .A(n50789), .B(n50790), .Z(n50788) );
  IV U60337 ( .A(n50791), .Z(n50790) );
  NANDN U60338 ( .A(n50791), .B(n50789), .Z(n50785) );
  AND U60339 ( .A(n50792), .B(n50793), .Z(n50766) );
  NAND U60340 ( .A(n50794), .B(n50795), .Z(n50793) );
  NANDN U60341 ( .A(n50796), .B(n50797), .Z(n50795) );
  NANDN U60342 ( .A(n50797), .B(n50796), .Z(n50792) );
  IV U60343 ( .A(n50798), .Z(n50797) );
  NAND U60344 ( .A(n50799), .B(n50800), .Z(n50769) );
  NANDN U60345 ( .A(n50801), .B(n50802), .Z(n50800) );
  NANDN U60346 ( .A(n50803), .B(n50804), .Z(n50802) );
  NANDN U60347 ( .A(n50804), .B(n50803), .Z(n50799) );
  IV U60348 ( .A(n50805), .Z(n50803) );
  AND U60349 ( .A(n50806), .B(n50807), .Z(n50772) );
  NAND U60350 ( .A(n50808), .B(n50809), .Z(n50807) );
  NANDN U60351 ( .A(n50810), .B(n50811), .Z(n50809) );
  NANDN U60352 ( .A(n50811), .B(n50810), .Z(n50806) );
  XOR U60353 ( .A(n50782), .B(n50812), .Z(n50774) );
  XNOR U60354 ( .A(n50779), .B(n50781), .Z(n50812) );
  AND U60355 ( .A(n50813), .B(n50814), .Z(n50781) );
  NANDN U60356 ( .A(n50815), .B(n50816), .Z(n50814) );
  OR U60357 ( .A(n50817), .B(n50818), .Z(n50816) );
  IV U60358 ( .A(n50819), .Z(n50818) );
  NANDN U60359 ( .A(n50819), .B(n50817), .Z(n50813) );
  AND U60360 ( .A(n50820), .B(n50821), .Z(n50779) );
  NAND U60361 ( .A(n50822), .B(n50823), .Z(n50821) );
  NANDN U60362 ( .A(n50824), .B(n50825), .Z(n50823) );
  NANDN U60363 ( .A(n50825), .B(n50824), .Z(n50820) );
  IV U60364 ( .A(n50826), .Z(n50825) );
  NAND U60365 ( .A(n50827), .B(n50828), .Z(n50782) );
  NANDN U60366 ( .A(n50829), .B(n50830), .Z(n50828) );
  NANDN U60367 ( .A(n50831), .B(n50832), .Z(n50830) );
  NANDN U60368 ( .A(n50832), .B(n50831), .Z(n50827) );
  IV U60369 ( .A(n50833), .Z(n50831) );
  XOR U60370 ( .A(n50808), .B(n50834), .Z(N60866) );
  XNOR U60371 ( .A(n50811), .B(n50810), .Z(n50834) );
  XNOR U60372 ( .A(n50822), .B(n50835), .Z(n50810) );
  XNOR U60373 ( .A(n50826), .B(n50824), .Z(n50835) );
  XOR U60374 ( .A(n50832), .B(n50836), .Z(n50824) );
  XNOR U60375 ( .A(n50829), .B(n50833), .Z(n50836) );
  AND U60376 ( .A(n50837), .B(n50838), .Z(n50833) );
  NAND U60377 ( .A(n50839), .B(n50840), .Z(n50838) );
  NAND U60378 ( .A(n50841), .B(n50842), .Z(n50837) );
  AND U60379 ( .A(n50843), .B(n50844), .Z(n50829) );
  NAND U60380 ( .A(n50845), .B(n50846), .Z(n50844) );
  NAND U60381 ( .A(n50847), .B(n50848), .Z(n50843) );
  NANDN U60382 ( .A(n50849), .B(n50850), .Z(n50832) );
  ANDN U60383 ( .B(n50851), .A(n50852), .Z(n50826) );
  XNOR U60384 ( .A(n50817), .B(n50853), .Z(n50822) );
  XNOR U60385 ( .A(n50815), .B(n50819), .Z(n50853) );
  AND U60386 ( .A(n50854), .B(n50855), .Z(n50819) );
  NAND U60387 ( .A(n50856), .B(n50857), .Z(n50855) );
  NAND U60388 ( .A(n50858), .B(n50859), .Z(n50854) );
  AND U60389 ( .A(n50860), .B(n50861), .Z(n50815) );
  NAND U60390 ( .A(n50862), .B(n50863), .Z(n50861) );
  NAND U60391 ( .A(n50864), .B(n50865), .Z(n50860) );
  AND U60392 ( .A(n50866), .B(n50867), .Z(n50817) );
  NAND U60393 ( .A(n50868), .B(n50869), .Z(n50811) );
  XNOR U60394 ( .A(n50794), .B(n50870), .Z(n50808) );
  XNOR U60395 ( .A(n50798), .B(n50796), .Z(n50870) );
  XOR U60396 ( .A(n50804), .B(n50871), .Z(n50796) );
  XNOR U60397 ( .A(n50801), .B(n50805), .Z(n50871) );
  AND U60398 ( .A(n50872), .B(n50873), .Z(n50805) );
  NAND U60399 ( .A(n50874), .B(n50875), .Z(n50873) );
  NAND U60400 ( .A(n50876), .B(n50877), .Z(n50872) );
  AND U60401 ( .A(n50878), .B(n50879), .Z(n50801) );
  NAND U60402 ( .A(n50880), .B(n50881), .Z(n50879) );
  NAND U60403 ( .A(n50882), .B(n50883), .Z(n50878) );
  NANDN U60404 ( .A(n50884), .B(n50885), .Z(n50804) );
  ANDN U60405 ( .B(n50886), .A(n50887), .Z(n50798) );
  XNOR U60406 ( .A(n50789), .B(n50888), .Z(n50794) );
  XNOR U60407 ( .A(n50787), .B(n50791), .Z(n50888) );
  AND U60408 ( .A(n50889), .B(n50890), .Z(n50791) );
  NAND U60409 ( .A(n50891), .B(n50892), .Z(n50890) );
  NAND U60410 ( .A(n50893), .B(n50894), .Z(n50889) );
  AND U60411 ( .A(n50895), .B(n50896), .Z(n50787) );
  NAND U60412 ( .A(n50897), .B(n50898), .Z(n50896) );
  NAND U60413 ( .A(n50899), .B(n50900), .Z(n50895) );
  AND U60414 ( .A(n50901), .B(n50902), .Z(n50789) );
  XOR U60415 ( .A(n50869), .B(n50868), .Z(N60865) );
  XNOR U60416 ( .A(n50886), .B(n50887), .Z(n50868) );
  XNOR U60417 ( .A(n50901), .B(n50902), .Z(n50887) );
  XOR U60418 ( .A(n50898), .B(n50897), .Z(n50902) );
  XOR U60419 ( .A(y[516]), .B(x[516]), .Z(n50897) );
  XOR U60420 ( .A(n50900), .B(n50899), .Z(n50898) );
  XOR U60421 ( .A(y[518]), .B(x[518]), .Z(n50899) );
  XOR U60422 ( .A(y[517]), .B(x[517]), .Z(n50900) );
  XOR U60423 ( .A(n50892), .B(n50891), .Z(n50901) );
  XOR U60424 ( .A(n50894), .B(n50893), .Z(n50891) );
  XOR U60425 ( .A(y[515]), .B(x[515]), .Z(n50893) );
  XOR U60426 ( .A(y[514]), .B(x[514]), .Z(n50894) );
  XOR U60427 ( .A(y[513]), .B(x[513]), .Z(n50892) );
  XNOR U60428 ( .A(n50885), .B(n50884), .Z(n50886) );
  XNOR U60429 ( .A(n50881), .B(n50880), .Z(n50884) );
  XOR U60430 ( .A(n50883), .B(n50882), .Z(n50880) );
  XOR U60431 ( .A(y[512]), .B(x[512]), .Z(n50882) );
  XOR U60432 ( .A(y[511]), .B(x[511]), .Z(n50883) );
  XOR U60433 ( .A(y[510]), .B(x[510]), .Z(n50881) );
  XOR U60434 ( .A(n50875), .B(n50874), .Z(n50885) );
  XOR U60435 ( .A(n50877), .B(n50876), .Z(n50874) );
  XOR U60436 ( .A(y[509]), .B(x[509]), .Z(n50876) );
  XOR U60437 ( .A(y[508]), .B(x[508]), .Z(n50877) );
  XOR U60438 ( .A(y[507]), .B(x[507]), .Z(n50875) );
  XNOR U60439 ( .A(n50851), .B(n50852), .Z(n50869) );
  XNOR U60440 ( .A(n50866), .B(n50867), .Z(n50852) );
  XOR U60441 ( .A(n50863), .B(n50862), .Z(n50867) );
  XOR U60442 ( .A(y[504]), .B(x[504]), .Z(n50862) );
  XOR U60443 ( .A(n50865), .B(n50864), .Z(n50863) );
  XOR U60444 ( .A(y[506]), .B(x[506]), .Z(n50864) );
  XOR U60445 ( .A(y[505]), .B(x[505]), .Z(n50865) );
  XOR U60446 ( .A(n50857), .B(n50856), .Z(n50866) );
  XOR U60447 ( .A(n50859), .B(n50858), .Z(n50856) );
  XOR U60448 ( .A(y[503]), .B(x[503]), .Z(n50858) );
  XOR U60449 ( .A(y[502]), .B(x[502]), .Z(n50859) );
  XOR U60450 ( .A(y[501]), .B(x[501]), .Z(n50857) );
  XNOR U60451 ( .A(n50850), .B(n50849), .Z(n50851) );
  XNOR U60452 ( .A(n50846), .B(n50845), .Z(n50849) );
  XOR U60453 ( .A(n50848), .B(n50847), .Z(n50845) );
  XOR U60454 ( .A(y[500]), .B(x[500]), .Z(n50847) );
  XOR U60455 ( .A(y[499]), .B(x[499]), .Z(n50848) );
  XOR U60456 ( .A(y[498]), .B(x[498]), .Z(n50846) );
  XOR U60457 ( .A(n50840), .B(n50839), .Z(n50850) );
  XOR U60458 ( .A(n50842), .B(n50841), .Z(n50839) );
  XOR U60459 ( .A(y[497]), .B(x[497]), .Z(n50841) );
  XOR U60460 ( .A(y[496]), .B(x[496]), .Z(n50842) );
  XOR U60461 ( .A(y[495]), .B(x[495]), .Z(n50840) );
  NAND U60462 ( .A(n50903), .B(n50904), .Z(N60856) );
  NAND U60463 ( .A(n50905), .B(n50906), .Z(n50904) );
  NANDN U60464 ( .A(n50907), .B(n50908), .Z(n50906) );
  NANDN U60465 ( .A(n50908), .B(n50907), .Z(n50903) );
  XOR U60466 ( .A(n50907), .B(n50909), .Z(N60855) );
  XNOR U60467 ( .A(n50905), .B(n50908), .Z(n50909) );
  NAND U60468 ( .A(n50910), .B(n50911), .Z(n50908) );
  NAND U60469 ( .A(n50912), .B(n50913), .Z(n50911) );
  NANDN U60470 ( .A(n50914), .B(n50915), .Z(n50913) );
  NANDN U60471 ( .A(n50915), .B(n50914), .Z(n50910) );
  AND U60472 ( .A(n50916), .B(n50917), .Z(n50905) );
  NAND U60473 ( .A(n50918), .B(n50919), .Z(n50917) );
  NANDN U60474 ( .A(n50920), .B(n50921), .Z(n50919) );
  NANDN U60475 ( .A(n50921), .B(n50920), .Z(n50916) );
  IV U60476 ( .A(n50922), .Z(n50921) );
  AND U60477 ( .A(n50923), .B(n50924), .Z(n50907) );
  NAND U60478 ( .A(n50925), .B(n50926), .Z(n50924) );
  NANDN U60479 ( .A(n50927), .B(n50928), .Z(n50926) );
  NANDN U60480 ( .A(n50928), .B(n50927), .Z(n50923) );
  XOR U60481 ( .A(n50920), .B(n50929), .Z(N60854) );
  XNOR U60482 ( .A(n50918), .B(n50922), .Z(n50929) );
  XOR U60483 ( .A(n50915), .B(n50930), .Z(n50922) );
  XNOR U60484 ( .A(n50912), .B(n50914), .Z(n50930) );
  AND U60485 ( .A(n50931), .B(n50932), .Z(n50914) );
  NANDN U60486 ( .A(n50933), .B(n50934), .Z(n50932) );
  OR U60487 ( .A(n50935), .B(n50936), .Z(n50934) );
  IV U60488 ( .A(n50937), .Z(n50936) );
  NANDN U60489 ( .A(n50937), .B(n50935), .Z(n50931) );
  AND U60490 ( .A(n50938), .B(n50939), .Z(n50912) );
  NAND U60491 ( .A(n50940), .B(n50941), .Z(n50939) );
  NANDN U60492 ( .A(n50942), .B(n50943), .Z(n50941) );
  NANDN U60493 ( .A(n50943), .B(n50942), .Z(n50938) );
  IV U60494 ( .A(n50944), .Z(n50943) );
  NAND U60495 ( .A(n50945), .B(n50946), .Z(n50915) );
  NANDN U60496 ( .A(n50947), .B(n50948), .Z(n50946) );
  NANDN U60497 ( .A(n50949), .B(n50950), .Z(n50948) );
  NANDN U60498 ( .A(n50950), .B(n50949), .Z(n50945) );
  IV U60499 ( .A(n50951), .Z(n50949) );
  AND U60500 ( .A(n50952), .B(n50953), .Z(n50918) );
  NAND U60501 ( .A(n50954), .B(n50955), .Z(n50953) );
  NANDN U60502 ( .A(n50956), .B(n50957), .Z(n50955) );
  NANDN U60503 ( .A(n50957), .B(n50956), .Z(n50952) );
  XOR U60504 ( .A(n50928), .B(n50958), .Z(n50920) );
  XNOR U60505 ( .A(n50925), .B(n50927), .Z(n50958) );
  AND U60506 ( .A(n50959), .B(n50960), .Z(n50927) );
  NANDN U60507 ( .A(n50961), .B(n50962), .Z(n50960) );
  OR U60508 ( .A(n50963), .B(n50964), .Z(n50962) );
  IV U60509 ( .A(n50965), .Z(n50964) );
  NANDN U60510 ( .A(n50965), .B(n50963), .Z(n50959) );
  AND U60511 ( .A(n50966), .B(n50967), .Z(n50925) );
  NAND U60512 ( .A(n50968), .B(n50969), .Z(n50967) );
  NANDN U60513 ( .A(n50970), .B(n50971), .Z(n50969) );
  NANDN U60514 ( .A(n50971), .B(n50970), .Z(n50966) );
  IV U60515 ( .A(n50972), .Z(n50971) );
  NAND U60516 ( .A(n50973), .B(n50974), .Z(n50928) );
  NANDN U60517 ( .A(n50975), .B(n50976), .Z(n50974) );
  NANDN U60518 ( .A(n50977), .B(n50978), .Z(n50976) );
  NANDN U60519 ( .A(n50978), .B(n50977), .Z(n50973) );
  IV U60520 ( .A(n50979), .Z(n50977) );
  XOR U60521 ( .A(n50954), .B(n50980), .Z(N60853) );
  XNOR U60522 ( .A(n50957), .B(n50956), .Z(n50980) );
  XNOR U60523 ( .A(n50968), .B(n50981), .Z(n50956) );
  XNOR U60524 ( .A(n50972), .B(n50970), .Z(n50981) );
  XOR U60525 ( .A(n50978), .B(n50982), .Z(n50970) );
  XNOR U60526 ( .A(n50975), .B(n50979), .Z(n50982) );
  AND U60527 ( .A(n50983), .B(n50984), .Z(n50979) );
  NAND U60528 ( .A(n50985), .B(n50986), .Z(n50984) );
  NAND U60529 ( .A(n50987), .B(n50988), .Z(n50983) );
  AND U60530 ( .A(n50989), .B(n50990), .Z(n50975) );
  NAND U60531 ( .A(n50991), .B(n50992), .Z(n50990) );
  NAND U60532 ( .A(n50993), .B(n50994), .Z(n50989) );
  NANDN U60533 ( .A(n50995), .B(n50996), .Z(n50978) );
  ANDN U60534 ( .B(n50997), .A(n50998), .Z(n50972) );
  XNOR U60535 ( .A(n50963), .B(n50999), .Z(n50968) );
  XNOR U60536 ( .A(n50961), .B(n50965), .Z(n50999) );
  AND U60537 ( .A(n51000), .B(n51001), .Z(n50965) );
  NAND U60538 ( .A(n51002), .B(n51003), .Z(n51001) );
  NAND U60539 ( .A(n51004), .B(n51005), .Z(n51000) );
  AND U60540 ( .A(n51006), .B(n51007), .Z(n50961) );
  NAND U60541 ( .A(n51008), .B(n51009), .Z(n51007) );
  NAND U60542 ( .A(n51010), .B(n51011), .Z(n51006) );
  AND U60543 ( .A(n51012), .B(n51013), .Z(n50963) );
  NAND U60544 ( .A(n51014), .B(n51015), .Z(n50957) );
  XNOR U60545 ( .A(n50940), .B(n51016), .Z(n50954) );
  XNOR U60546 ( .A(n50944), .B(n50942), .Z(n51016) );
  XOR U60547 ( .A(n50950), .B(n51017), .Z(n50942) );
  XNOR U60548 ( .A(n50947), .B(n50951), .Z(n51017) );
  AND U60549 ( .A(n51018), .B(n51019), .Z(n50951) );
  NAND U60550 ( .A(n51020), .B(n51021), .Z(n51019) );
  NAND U60551 ( .A(n51022), .B(n51023), .Z(n51018) );
  AND U60552 ( .A(n51024), .B(n51025), .Z(n50947) );
  NAND U60553 ( .A(n51026), .B(n51027), .Z(n51025) );
  NAND U60554 ( .A(n51028), .B(n51029), .Z(n51024) );
  NANDN U60555 ( .A(n51030), .B(n51031), .Z(n50950) );
  ANDN U60556 ( .B(n51032), .A(n51033), .Z(n50944) );
  XNOR U60557 ( .A(n50935), .B(n51034), .Z(n50940) );
  XNOR U60558 ( .A(n50933), .B(n50937), .Z(n51034) );
  AND U60559 ( .A(n51035), .B(n51036), .Z(n50937) );
  NAND U60560 ( .A(n51037), .B(n51038), .Z(n51036) );
  NAND U60561 ( .A(n51039), .B(n51040), .Z(n51035) );
  AND U60562 ( .A(n51041), .B(n51042), .Z(n50933) );
  NAND U60563 ( .A(n51043), .B(n51044), .Z(n51042) );
  NAND U60564 ( .A(n51045), .B(n51046), .Z(n51041) );
  AND U60565 ( .A(n51047), .B(n51048), .Z(n50935) );
  XOR U60566 ( .A(n51015), .B(n51014), .Z(N60852) );
  XNOR U60567 ( .A(n51032), .B(n51033), .Z(n51014) );
  XNOR U60568 ( .A(n51047), .B(n51048), .Z(n51033) );
  XOR U60569 ( .A(n51044), .B(n51043), .Z(n51048) );
  XOR U60570 ( .A(y[492]), .B(x[492]), .Z(n51043) );
  XOR U60571 ( .A(n51046), .B(n51045), .Z(n51044) );
  XOR U60572 ( .A(y[494]), .B(x[494]), .Z(n51045) );
  XOR U60573 ( .A(y[493]), .B(x[493]), .Z(n51046) );
  XOR U60574 ( .A(n51038), .B(n51037), .Z(n51047) );
  XOR U60575 ( .A(n51040), .B(n51039), .Z(n51037) );
  XOR U60576 ( .A(y[491]), .B(x[491]), .Z(n51039) );
  XOR U60577 ( .A(y[490]), .B(x[490]), .Z(n51040) );
  XOR U60578 ( .A(y[489]), .B(x[489]), .Z(n51038) );
  XNOR U60579 ( .A(n51031), .B(n51030), .Z(n51032) );
  XNOR U60580 ( .A(n51027), .B(n51026), .Z(n51030) );
  XOR U60581 ( .A(n51029), .B(n51028), .Z(n51026) );
  XOR U60582 ( .A(y[488]), .B(x[488]), .Z(n51028) );
  XOR U60583 ( .A(y[487]), .B(x[487]), .Z(n51029) );
  XOR U60584 ( .A(y[486]), .B(x[486]), .Z(n51027) );
  XOR U60585 ( .A(n51021), .B(n51020), .Z(n51031) );
  XOR U60586 ( .A(n51023), .B(n51022), .Z(n51020) );
  XOR U60587 ( .A(y[485]), .B(x[485]), .Z(n51022) );
  XOR U60588 ( .A(y[484]), .B(x[484]), .Z(n51023) );
  XOR U60589 ( .A(y[483]), .B(x[483]), .Z(n51021) );
  XNOR U60590 ( .A(n50997), .B(n50998), .Z(n51015) );
  XNOR U60591 ( .A(n51012), .B(n51013), .Z(n50998) );
  XOR U60592 ( .A(n51009), .B(n51008), .Z(n51013) );
  XOR U60593 ( .A(y[480]), .B(x[480]), .Z(n51008) );
  XOR U60594 ( .A(n51011), .B(n51010), .Z(n51009) );
  XOR U60595 ( .A(y[482]), .B(x[482]), .Z(n51010) );
  XOR U60596 ( .A(y[481]), .B(x[481]), .Z(n51011) );
  XOR U60597 ( .A(n51003), .B(n51002), .Z(n51012) );
  XOR U60598 ( .A(n51005), .B(n51004), .Z(n51002) );
  XOR U60599 ( .A(y[479]), .B(x[479]), .Z(n51004) );
  XOR U60600 ( .A(y[478]), .B(x[478]), .Z(n51005) );
  XOR U60601 ( .A(y[477]), .B(x[477]), .Z(n51003) );
  XNOR U60602 ( .A(n50996), .B(n50995), .Z(n50997) );
  XNOR U60603 ( .A(n50992), .B(n50991), .Z(n50995) );
  XOR U60604 ( .A(n50994), .B(n50993), .Z(n50991) );
  XOR U60605 ( .A(y[476]), .B(x[476]), .Z(n50993) );
  XOR U60606 ( .A(y[475]), .B(x[475]), .Z(n50994) );
  XOR U60607 ( .A(y[474]), .B(x[474]), .Z(n50992) );
  XOR U60608 ( .A(n50986), .B(n50985), .Z(n50996) );
  XOR U60609 ( .A(n50988), .B(n50987), .Z(n50985) );
  XOR U60610 ( .A(y[473]), .B(x[473]), .Z(n50987) );
  XOR U60611 ( .A(y[472]), .B(x[472]), .Z(n50988) );
  XOR U60612 ( .A(y[471]), .B(x[471]), .Z(n50986) );
  NAND U60613 ( .A(n51049), .B(n51050), .Z(N60843) );
  NAND U60614 ( .A(n51051), .B(n51052), .Z(n51050) );
  NANDN U60615 ( .A(n51053), .B(n51054), .Z(n51052) );
  NANDN U60616 ( .A(n51054), .B(n51053), .Z(n51049) );
  XOR U60617 ( .A(n51053), .B(n51055), .Z(N60842) );
  XNOR U60618 ( .A(n51051), .B(n51054), .Z(n51055) );
  NAND U60619 ( .A(n51056), .B(n51057), .Z(n51054) );
  NAND U60620 ( .A(n51058), .B(n51059), .Z(n51057) );
  NANDN U60621 ( .A(n51060), .B(n51061), .Z(n51059) );
  NANDN U60622 ( .A(n51061), .B(n51060), .Z(n51056) );
  AND U60623 ( .A(n51062), .B(n51063), .Z(n51051) );
  NAND U60624 ( .A(n51064), .B(n51065), .Z(n51063) );
  NANDN U60625 ( .A(n51066), .B(n51067), .Z(n51065) );
  NANDN U60626 ( .A(n51067), .B(n51066), .Z(n51062) );
  IV U60627 ( .A(n51068), .Z(n51067) );
  AND U60628 ( .A(n51069), .B(n51070), .Z(n51053) );
  NAND U60629 ( .A(n51071), .B(n51072), .Z(n51070) );
  NANDN U60630 ( .A(n51073), .B(n51074), .Z(n51072) );
  NANDN U60631 ( .A(n51074), .B(n51073), .Z(n51069) );
  XOR U60632 ( .A(n51066), .B(n51075), .Z(N60841) );
  XNOR U60633 ( .A(n51064), .B(n51068), .Z(n51075) );
  XOR U60634 ( .A(n51061), .B(n51076), .Z(n51068) );
  XNOR U60635 ( .A(n51058), .B(n51060), .Z(n51076) );
  AND U60636 ( .A(n51077), .B(n51078), .Z(n51060) );
  NANDN U60637 ( .A(n51079), .B(n51080), .Z(n51078) );
  OR U60638 ( .A(n51081), .B(n51082), .Z(n51080) );
  IV U60639 ( .A(n51083), .Z(n51082) );
  NANDN U60640 ( .A(n51083), .B(n51081), .Z(n51077) );
  AND U60641 ( .A(n51084), .B(n51085), .Z(n51058) );
  NAND U60642 ( .A(n51086), .B(n51087), .Z(n51085) );
  NANDN U60643 ( .A(n51088), .B(n51089), .Z(n51087) );
  NANDN U60644 ( .A(n51089), .B(n51088), .Z(n51084) );
  IV U60645 ( .A(n51090), .Z(n51089) );
  NAND U60646 ( .A(n51091), .B(n51092), .Z(n51061) );
  NANDN U60647 ( .A(n51093), .B(n51094), .Z(n51092) );
  NANDN U60648 ( .A(n51095), .B(n51096), .Z(n51094) );
  NANDN U60649 ( .A(n51096), .B(n51095), .Z(n51091) );
  IV U60650 ( .A(n51097), .Z(n51095) );
  AND U60651 ( .A(n51098), .B(n51099), .Z(n51064) );
  NAND U60652 ( .A(n51100), .B(n51101), .Z(n51099) );
  NANDN U60653 ( .A(n51102), .B(n51103), .Z(n51101) );
  NANDN U60654 ( .A(n51103), .B(n51102), .Z(n51098) );
  XOR U60655 ( .A(n51074), .B(n51104), .Z(n51066) );
  XNOR U60656 ( .A(n51071), .B(n51073), .Z(n51104) );
  AND U60657 ( .A(n51105), .B(n51106), .Z(n51073) );
  NANDN U60658 ( .A(n51107), .B(n51108), .Z(n51106) );
  OR U60659 ( .A(n51109), .B(n51110), .Z(n51108) );
  IV U60660 ( .A(n51111), .Z(n51110) );
  NANDN U60661 ( .A(n51111), .B(n51109), .Z(n51105) );
  AND U60662 ( .A(n51112), .B(n51113), .Z(n51071) );
  NAND U60663 ( .A(n51114), .B(n51115), .Z(n51113) );
  NANDN U60664 ( .A(n51116), .B(n51117), .Z(n51115) );
  NANDN U60665 ( .A(n51117), .B(n51116), .Z(n51112) );
  IV U60666 ( .A(n51118), .Z(n51117) );
  NAND U60667 ( .A(n51119), .B(n51120), .Z(n51074) );
  NANDN U60668 ( .A(n51121), .B(n51122), .Z(n51120) );
  NANDN U60669 ( .A(n51123), .B(n51124), .Z(n51122) );
  NANDN U60670 ( .A(n51124), .B(n51123), .Z(n51119) );
  IV U60671 ( .A(n51125), .Z(n51123) );
  XOR U60672 ( .A(n51100), .B(n51126), .Z(N60840) );
  XNOR U60673 ( .A(n51103), .B(n51102), .Z(n51126) );
  XNOR U60674 ( .A(n51114), .B(n51127), .Z(n51102) );
  XNOR U60675 ( .A(n51118), .B(n51116), .Z(n51127) );
  XOR U60676 ( .A(n51124), .B(n51128), .Z(n51116) );
  XNOR U60677 ( .A(n51121), .B(n51125), .Z(n51128) );
  AND U60678 ( .A(n51129), .B(n51130), .Z(n51125) );
  NAND U60679 ( .A(n51131), .B(n51132), .Z(n51130) );
  NAND U60680 ( .A(n51133), .B(n51134), .Z(n51129) );
  AND U60681 ( .A(n51135), .B(n51136), .Z(n51121) );
  NAND U60682 ( .A(n51137), .B(n51138), .Z(n51136) );
  NAND U60683 ( .A(n51139), .B(n51140), .Z(n51135) );
  NANDN U60684 ( .A(n51141), .B(n51142), .Z(n51124) );
  ANDN U60685 ( .B(n51143), .A(n51144), .Z(n51118) );
  XNOR U60686 ( .A(n51109), .B(n51145), .Z(n51114) );
  XNOR U60687 ( .A(n51107), .B(n51111), .Z(n51145) );
  AND U60688 ( .A(n51146), .B(n51147), .Z(n51111) );
  NAND U60689 ( .A(n51148), .B(n51149), .Z(n51147) );
  NAND U60690 ( .A(n51150), .B(n51151), .Z(n51146) );
  AND U60691 ( .A(n51152), .B(n51153), .Z(n51107) );
  NAND U60692 ( .A(n51154), .B(n51155), .Z(n51153) );
  NAND U60693 ( .A(n51156), .B(n51157), .Z(n51152) );
  AND U60694 ( .A(n51158), .B(n51159), .Z(n51109) );
  NAND U60695 ( .A(n51160), .B(n51161), .Z(n51103) );
  XNOR U60696 ( .A(n51086), .B(n51162), .Z(n51100) );
  XNOR U60697 ( .A(n51090), .B(n51088), .Z(n51162) );
  XOR U60698 ( .A(n51096), .B(n51163), .Z(n51088) );
  XNOR U60699 ( .A(n51093), .B(n51097), .Z(n51163) );
  AND U60700 ( .A(n51164), .B(n51165), .Z(n51097) );
  NAND U60701 ( .A(n51166), .B(n51167), .Z(n51165) );
  NAND U60702 ( .A(n51168), .B(n51169), .Z(n51164) );
  AND U60703 ( .A(n51170), .B(n51171), .Z(n51093) );
  NAND U60704 ( .A(n51172), .B(n51173), .Z(n51171) );
  NAND U60705 ( .A(n51174), .B(n51175), .Z(n51170) );
  NANDN U60706 ( .A(n51176), .B(n51177), .Z(n51096) );
  ANDN U60707 ( .B(n51178), .A(n51179), .Z(n51090) );
  XNOR U60708 ( .A(n51081), .B(n51180), .Z(n51086) );
  XNOR U60709 ( .A(n51079), .B(n51083), .Z(n51180) );
  AND U60710 ( .A(n51181), .B(n51182), .Z(n51083) );
  NAND U60711 ( .A(n51183), .B(n51184), .Z(n51182) );
  NAND U60712 ( .A(n51185), .B(n51186), .Z(n51181) );
  AND U60713 ( .A(n51187), .B(n51188), .Z(n51079) );
  NAND U60714 ( .A(n51189), .B(n51190), .Z(n51188) );
  NAND U60715 ( .A(n51191), .B(n51192), .Z(n51187) );
  AND U60716 ( .A(n51193), .B(n51194), .Z(n51081) );
  XOR U60717 ( .A(n51161), .B(n51160), .Z(N60839) );
  XNOR U60718 ( .A(n51178), .B(n51179), .Z(n51160) );
  XNOR U60719 ( .A(n51193), .B(n51194), .Z(n51179) );
  XOR U60720 ( .A(n51190), .B(n51189), .Z(n51194) );
  XOR U60721 ( .A(y[468]), .B(x[468]), .Z(n51189) );
  XOR U60722 ( .A(n51192), .B(n51191), .Z(n51190) );
  XOR U60723 ( .A(y[470]), .B(x[470]), .Z(n51191) );
  XOR U60724 ( .A(y[469]), .B(x[469]), .Z(n51192) );
  XOR U60725 ( .A(n51184), .B(n51183), .Z(n51193) );
  XOR U60726 ( .A(n51186), .B(n51185), .Z(n51183) );
  XOR U60727 ( .A(y[467]), .B(x[467]), .Z(n51185) );
  XOR U60728 ( .A(y[466]), .B(x[466]), .Z(n51186) );
  XOR U60729 ( .A(y[465]), .B(x[465]), .Z(n51184) );
  XNOR U60730 ( .A(n51177), .B(n51176), .Z(n51178) );
  XNOR U60731 ( .A(n51173), .B(n51172), .Z(n51176) );
  XOR U60732 ( .A(n51175), .B(n51174), .Z(n51172) );
  XOR U60733 ( .A(y[464]), .B(x[464]), .Z(n51174) );
  XOR U60734 ( .A(y[463]), .B(x[463]), .Z(n51175) );
  XOR U60735 ( .A(y[462]), .B(x[462]), .Z(n51173) );
  XOR U60736 ( .A(n51167), .B(n51166), .Z(n51177) );
  XOR U60737 ( .A(n51169), .B(n51168), .Z(n51166) );
  XOR U60738 ( .A(y[461]), .B(x[461]), .Z(n51168) );
  XOR U60739 ( .A(y[460]), .B(x[460]), .Z(n51169) );
  XOR U60740 ( .A(y[459]), .B(x[459]), .Z(n51167) );
  XNOR U60741 ( .A(n51143), .B(n51144), .Z(n51161) );
  XNOR U60742 ( .A(n51158), .B(n51159), .Z(n51144) );
  XOR U60743 ( .A(n51155), .B(n51154), .Z(n51159) );
  XOR U60744 ( .A(y[456]), .B(x[456]), .Z(n51154) );
  XOR U60745 ( .A(n51157), .B(n51156), .Z(n51155) );
  XOR U60746 ( .A(y[458]), .B(x[458]), .Z(n51156) );
  XOR U60747 ( .A(y[457]), .B(x[457]), .Z(n51157) );
  XOR U60748 ( .A(n51149), .B(n51148), .Z(n51158) );
  XOR U60749 ( .A(n51151), .B(n51150), .Z(n51148) );
  XOR U60750 ( .A(y[455]), .B(x[455]), .Z(n51150) );
  XOR U60751 ( .A(y[454]), .B(x[454]), .Z(n51151) );
  XOR U60752 ( .A(y[453]), .B(x[453]), .Z(n51149) );
  XNOR U60753 ( .A(n51142), .B(n51141), .Z(n51143) );
  XNOR U60754 ( .A(n51138), .B(n51137), .Z(n51141) );
  XOR U60755 ( .A(n51140), .B(n51139), .Z(n51137) );
  XOR U60756 ( .A(y[452]), .B(x[452]), .Z(n51139) );
  XOR U60757 ( .A(y[451]), .B(x[451]), .Z(n51140) );
  XOR U60758 ( .A(y[450]), .B(x[450]), .Z(n51138) );
  XOR U60759 ( .A(n51132), .B(n51131), .Z(n51142) );
  XOR U60760 ( .A(n51134), .B(n51133), .Z(n51131) );
  XOR U60761 ( .A(y[449]), .B(x[449]), .Z(n51133) );
  XOR U60762 ( .A(y[448]), .B(x[448]), .Z(n51134) );
  XOR U60763 ( .A(y[447]), .B(x[447]), .Z(n51132) );
  NAND U60764 ( .A(n51195), .B(n51196), .Z(N60830) );
  NAND U60765 ( .A(n51197), .B(n51198), .Z(n51196) );
  NANDN U60766 ( .A(n51199), .B(n51200), .Z(n51198) );
  NANDN U60767 ( .A(n51200), .B(n51199), .Z(n51195) );
  XOR U60768 ( .A(n51199), .B(n51201), .Z(N60829) );
  XNOR U60769 ( .A(n51197), .B(n51200), .Z(n51201) );
  NAND U60770 ( .A(n51202), .B(n51203), .Z(n51200) );
  NAND U60771 ( .A(n51204), .B(n51205), .Z(n51203) );
  NANDN U60772 ( .A(n51206), .B(n51207), .Z(n51205) );
  NANDN U60773 ( .A(n51207), .B(n51206), .Z(n51202) );
  AND U60774 ( .A(n51208), .B(n51209), .Z(n51197) );
  NAND U60775 ( .A(n51210), .B(n51211), .Z(n51209) );
  NANDN U60776 ( .A(n51212), .B(n51213), .Z(n51211) );
  NANDN U60777 ( .A(n51213), .B(n51212), .Z(n51208) );
  IV U60778 ( .A(n51214), .Z(n51213) );
  AND U60779 ( .A(n51215), .B(n51216), .Z(n51199) );
  NAND U60780 ( .A(n51217), .B(n51218), .Z(n51216) );
  NANDN U60781 ( .A(n51219), .B(n51220), .Z(n51218) );
  NANDN U60782 ( .A(n51220), .B(n51219), .Z(n51215) );
  XOR U60783 ( .A(n51212), .B(n51221), .Z(N60828) );
  XNOR U60784 ( .A(n51210), .B(n51214), .Z(n51221) );
  XOR U60785 ( .A(n51207), .B(n51222), .Z(n51214) );
  XNOR U60786 ( .A(n51204), .B(n51206), .Z(n51222) );
  AND U60787 ( .A(n51223), .B(n51224), .Z(n51206) );
  NANDN U60788 ( .A(n51225), .B(n51226), .Z(n51224) );
  OR U60789 ( .A(n51227), .B(n51228), .Z(n51226) );
  IV U60790 ( .A(n51229), .Z(n51228) );
  NANDN U60791 ( .A(n51229), .B(n51227), .Z(n51223) );
  AND U60792 ( .A(n51230), .B(n51231), .Z(n51204) );
  NAND U60793 ( .A(n51232), .B(n51233), .Z(n51231) );
  NANDN U60794 ( .A(n51234), .B(n51235), .Z(n51233) );
  NANDN U60795 ( .A(n51235), .B(n51234), .Z(n51230) );
  IV U60796 ( .A(n51236), .Z(n51235) );
  NAND U60797 ( .A(n51237), .B(n51238), .Z(n51207) );
  NANDN U60798 ( .A(n51239), .B(n51240), .Z(n51238) );
  NANDN U60799 ( .A(n51241), .B(n51242), .Z(n51240) );
  NANDN U60800 ( .A(n51242), .B(n51241), .Z(n51237) );
  IV U60801 ( .A(n51243), .Z(n51241) );
  AND U60802 ( .A(n51244), .B(n51245), .Z(n51210) );
  NAND U60803 ( .A(n51246), .B(n51247), .Z(n51245) );
  NANDN U60804 ( .A(n51248), .B(n51249), .Z(n51247) );
  NANDN U60805 ( .A(n51249), .B(n51248), .Z(n51244) );
  XOR U60806 ( .A(n51220), .B(n51250), .Z(n51212) );
  XNOR U60807 ( .A(n51217), .B(n51219), .Z(n51250) );
  AND U60808 ( .A(n51251), .B(n51252), .Z(n51219) );
  NANDN U60809 ( .A(n51253), .B(n51254), .Z(n51252) );
  OR U60810 ( .A(n51255), .B(n51256), .Z(n51254) );
  IV U60811 ( .A(n51257), .Z(n51256) );
  NANDN U60812 ( .A(n51257), .B(n51255), .Z(n51251) );
  AND U60813 ( .A(n51258), .B(n51259), .Z(n51217) );
  NAND U60814 ( .A(n51260), .B(n51261), .Z(n51259) );
  NANDN U60815 ( .A(n51262), .B(n51263), .Z(n51261) );
  NANDN U60816 ( .A(n51263), .B(n51262), .Z(n51258) );
  IV U60817 ( .A(n51264), .Z(n51263) );
  NAND U60818 ( .A(n51265), .B(n51266), .Z(n51220) );
  NANDN U60819 ( .A(n51267), .B(n51268), .Z(n51266) );
  NANDN U60820 ( .A(n51269), .B(n51270), .Z(n51268) );
  NANDN U60821 ( .A(n51270), .B(n51269), .Z(n51265) );
  IV U60822 ( .A(n51271), .Z(n51269) );
  XOR U60823 ( .A(n51246), .B(n51272), .Z(N60827) );
  XNOR U60824 ( .A(n51249), .B(n51248), .Z(n51272) );
  XNOR U60825 ( .A(n51260), .B(n51273), .Z(n51248) );
  XNOR U60826 ( .A(n51264), .B(n51262), .Z(n51273) );
  XOR U60827 ( .A(n51270), .B(n51274), .Z(n51262) );
  XNOR U60828 ( .A(n51267), .B(n51271), .Z(n51274) );
  AND U60829 ( .A(n51275), .B(n51276), .Z(n51271) );
  NAND U60830 ( .A(n51277), .B(n51278), .Z(n51276) );
  NAND U60831 ( .A(n51279), .B(n51280), .Z(n51275) );
  AND U60832 ( .A(n51281), .B(n51282), .Z(n51267) );
  NAND U60833 ( .A(n51283), .B(n51284), .Z(n51282) );
  NAND U60834 ( .A(n51285), .B(n51286), .Z(n51281) );
  NANDN U60835 ( .A(n51287), .B(n51288), .Z(n51270) );
  ANDN U60836 ( .B(n51289), .A(n51290), .Z(n51264) );
  XNOR U60837 ( .A(n51255), .B(n51291), .Z(n51260) );
  XNOR U60838 ( .A(n51253), .B(n51257), .Z(n51291) );
  AND U60839 ( .A(n51292), .B(n51293), .Z(n51257) );
  NAND U60840 ( .A(n51294), .B(n51295), .Z(n51293) );
  NAND U60841 ( .A(n51296), .B(n51297), .Z(n51292) );
  AND U60842 ( .A(n51298), .B(n51299), .Z(n51253) );
  NAND U60843 ( .A(n51300), .B(n51301), .Z(n51299) );
  NAND U60844 ( .A(n51302), .B(n51303), .Z(n51298) );
  AND U60845 ( .A(n51304), .B(n51305), .Z(n51255) );
  NAND U60846 ( .A(n51306), .B(n51307), .Z(n51249) );
  XNOR U60847 ( .A(n51232), .B(n51308), .Z(n51246) );
  XNOR U60848 ( .A(n51236), .B(n51234), .Z(n51308) );
  XOR U60849 ( .A(n51242), .B(n51309), .Z(n51234) );
  XNOR U60850 ( .A(n51239), .B(n51243), .Z(n51309) );
  AND U60851 ( .A(n51310), .B(n51311), .Z(n51243) );
  NAND U60852 ( .A(n51312), .B(n51313), .Z(n51311) );
  NAND U60853 ( .A(n51314), .B(n51315), .Z(n51310) );
  AND U60854 ( .A(n51316), .B(n51317), .Z(n51239) );
  NAND U60855 ( .A(n51318), .B(n51319), .Z(n51317) );
  NAND U60856 ( .A(n51320), .B(n51321), .Z(n51316) );
  NANDN U60857 ( .A(n51322), .B(n51323), .Z(n51242) );
  ANDN U60858 ( .B(n51324), .A(n51325), .Z(n51236) );
  XNOR U60859 ( .A(n51227), .B(n51326), .Z(n51232) );
  XNOR U60860 ( .A(n51225), .B(n51229), .Z(n51326) );
  AND U60861 ( .A(n51327), .B(n51328), .Z(n51229) );
  NAND U60862 ( .A(n51329), .B(n51330), .Z(n51328) );
  NAND U60863 ( .A(n51331), .B(n51332), .Z(n51327) );
  AND U60864 ( .A(n51333), .B(n51334), .Z(n51225) );
  NAND U60865 ( .A(n51335), .B(n51336), .Z(n51334) );
  NAND U60866 ( .A(n51337), .B(n51338), .Z(n51333) );
  AND U60867 ( .A(n51339), .B(n51340), .Z(n51227) );
  XOR U60868 ( .A(n51307), .B(n51306), .Z(N60826) );
  XNOR U60869 ( .A(n51324), .B(n51325), .Z(n51306) );
  XNOR U60870 ( .A(n51339), .B(n51340), .Z(n51325) );
  XOR U60871 ( .A(n51336), .B(n51335), .Z(n51340) );
  XOR U60872 ( .A(y[444]), .B(x[444]), .Z(n51335) );
  XOR U60873 ( .A(n51338), .B(n51337), .Z(n51336) );
  XOR U60874 ( .A(y[446]), .B(x[446]), .Z(n51337) );
  XOR U60875 ( .A(y[445]), .B(x[445]), .Z(n51338) );
  XOR U60876 ( .A(n51330), .B(n51329), .Z(n51339) );
  XOR U60877 ( .A(n51332), .B(n51331), .Z(n51329) );
  XOR U60878 ( .A(y[443]), .B(x[443]), .Z(n51331) );
  XOR U60879 ( .A(y[442]), .B(x[442]), .Z(n51332) );
  XOR U60880 ( .A(y[441]), .B(x[441]), .Z(n51330) );
  XNOR U60881 ( .A(n51323), .B(n51322), .Z(n51324) );
  XNOR U60882 ( .A(n51319), .B(n51318), .Z(n51322) );
  XOR U60883 ( .A(n51321), .B(n51320), .Z(n51318) );
  XOR U60884 ( .A(y[440]), .B(x[440]), .Z(n51320) );
  XOR U60885 ( .A(y[439]), .B(x[439]), .Z(n51321) );
  XOR U60886 ( .A(y[438]), .B(x[438]), .Z(n51319) );
  XOR U60887 ( .A(n51313), .B(n51312), .Z(n51323) );
  XOR U60888 ( .A(n51315), .B(n51314), .Z(n51312) );
  XOR U60889 ( .A(y[437]), .B(x[437]), .Z(n51314) );
  XOR U60890 ( .A(y[436]), .B(x[436]), .Z(n51315) );
  XOR U60891 ( .A(y[435]), .B(x[435]), .Z(n51313) );
  XNOR U60892 ( .A(n51289), .B(n51290), .Z(n51307) );
  XNOR U60893 ( .A(n51304), .B(n51305), .Z(n51290) );
  XOR U60894 ( .A(n51301), .B(n51300), .Z(n51305) );
  XOR U60895 ( .A(y[432]), .B(x[432]), .Z(n51300) );
  XOR U60896 ( .A(n51303), .B(n51302), .Z(n51301) );
  XOR U60897 ( .A(y[434]), .B(x[434]), .Z(n51302) );
  XOR U60898 ( .A(y[433]), .B(x[433]), .Z(n51303) );
  XOR U60899 ( .A(n51295), .B(n51294), .Z(n51304) );
  XOR U60900 ( .A(n51297), .B(n51296), .Z(n51294) );
  XOR U60901 ( .A(y[431]), .B(x[431]), .Z(n51296) );
  XOR U60902 ( .A(y[430]), .B(x[430]), .Z(n51297) );
  XOR U60903 ( .A(y[429]), .B(x[429]), .Z(n51295) );
  XNOR U60904 ( .A(n51288), .B(n51287), .Z(n51289) );
  XNOR U60905 ( .A(n51284), .B(n51283), .Z(n51287) );
  XOR U60906 ( .A(n51286), .B(n51285), .Z(n51283) );
  XOR U60907 ( .A(y[428]), .B(x[428]), .Z(n51285) );
  XOR U60908 ( .A(y[427]), .B(x[427]), .Z(n51286) );
  XOR U60909 ( .A(y[426]), .B(x[426]), .Z(n51284) );
  XOR U60910 ( .A(n51278), .B(n51277), .Z(n51288) );
  XOR U60911 ( .A(n51280), .B(n51279), .Z(n51277) );
  XOR U60912 ( .A(y[425]), .B(x[425]), .Z(n51279) );
  XOR U60913 ( .A(y[424]), .B(x[424]), .Z(n51280) );
  XOR U60914 ( .A(y[423]), .B(x[423]), .Z(n51278) );
  NAND U60915 ( .A(n51341), .B(n51342), .Z(N60817) );
  NAND U60916 ( .A(n51343), .B(n51344), .Z(n51342) );
  NANDN U60917 ( .A(n51345), .B(n51346), .Z(n51344) );
  NANDN U60918 ( .A(n51346), .B(n51345), .Z(n51341) );
  XOR U60919 ( .A(n51345), .B(n51347), .Z(N60816) );
  XNOR U60920 ( .A(n51343), .B(n51346), .Z(n51347) );
  NAND U60921 ( .A(n51348), .B(n51349), .Z(n51346) );
  NAND U60922 ( .A(n51350), .B(n51351), .Z(n51349) );
  NANDN U60923 ( .A(n51352), .B(n51353), .Z(n51351) );
  NANDN U60924 ( .A(n51353), .B(n51352), .Z(n51348) );
  AND U60925 ( .A(n51354), .B(n51355), .Z(n51343) );
  NAND U60926 ( .A(n51356), .B(n51357), .Z(n51355) );
  NANDN U60927 ( .A(n51358), .B(n51359), .Z(n51357) );
  NANDN U60928 ( .A(n51359), .B(n51358), .Z(n51354) );
  IV U60929 ( .A(n51360), .Z(n51359) );
  AND U60930 ( .A(n51361), .B(n51362), .Z(n51345) );
  NAND U60931 ( .A(n51363), .B(n51364), .Z(n51362) );
  NANDN U60932 ( .A(n51365), .B(n51366), .Z(n51364) );
  NANDN U60933 ( .A(n51366), .B(n51365), .Z(n51361) );
  XOR U60934 ( .A(n51358), .B(n51367), .Z(N60815) );
  XNOR U60935 ( .A(n51356), .B(n51360), .Z(n51367) );
  XOR U60936 ( .A(n51353), .B(n51368), .Z(n51360) );
  XNOR U60937 ( .A(n51350), .B(n51352), .Z(n51368) );
  AND U60938 ( .A(n51369), .B(n51370), .Z(n51352) );
  NANDN U60939 ( .A(n51371), .B(n51372), .Z(n51370) );
  OR U60940 ( .A(n51373), .B(n51374), .Z(n51372) );
  IV U60941 ( .A(n51375), .Z(n51374) );
  NANDN U60942 ( .A(n51375), .B(n51373), .Z(n51369) );
  AND U60943 ( .A(n51376), .B(n51377), .Z(n51350) );
  NAND U60944 ( .A(n51378), .B(n51379), .Z(n51377) );
  NANDN U60945 ( .A(n51380), .B(n51381), .Z(n51379) );
  NANDN U60946 ( .A(n51381), .B(n51380), .Z(n51376) );
  IV U60947 ( .A(n51382), .Z(n51381) );
  NAND U60948 ( .A(n51383), .B(n51384), .Z(n51353) );
  NANDN U60949 ( .A(n51385), .B(n51386), .Z(n51384) );
  NANDN U60950 ( .A(n51387), .B(n51388), .Z(n51386) );
  NANDN U60951 ( .A(n51388), .B(n51387), .Z(n51383) );
  IV U60952 ( .A(n51389), .Z(n51387) );
  AND U60953 ( .A(n51390), .B(n51391), .Z(n51356) );
  NAND U60954 ( .A(n51392), .B(n51393), .Z(n51391) );
  NANDN U60955 ( .A(n51394), .B(n51395), .Z(n51393) );
  NANDN U60956 ( .A(n51395), .B(n51394), .Z(n51390) );
  XOR U60957 ( .A(n51366), .B(n51396), .Z(n51358) );
  XNOR U60958 ( .A(n51363), .B(n51365), .Z(n51396) );
  AND U60959 ( .A(n51397), .B(n51398), .Z(n51365) );
  NANDN U60960 ( .A(n51399), .B(n51400), .Z(n51398) );
  OR U60961 ( .A(n51401), .B(n51402), .Z(n51400) );
  IV U60962 ( .A(n51403), .Z(n51402) );
  NANDN U60963 ( .A(n51403), .B(n51401), .Z(n51397) );
  AND U60964 ( .A(n51404), .B(n51405), .Z(n51363) );
  NAND U60965 ( .A(n51406), .B(n51407), .Z(n51405) );
  NANDN U60966 ( .A(n51408), .B(n51409), .Z(n51407) );
  NANDN U60967 ( .A(n51409), .B(n51408), .Z(n51404) );
  IV U60968 ( .A(n51410), .Z(n51409) );
  NAND U60969 ( .A(n51411), .B(n51412), .Z(n51366) );
  NANDN U60970 ( .A(n51413), .B(n51414), .Z(n51412) );
  NANDN U60971 ( .A(n51415), .B(n51416), .Z(n51414) );
  NANDN U60972 ( .A(n51416), .B(n51415), .Z(n51411) );
  IV U60973 ( .A(n51417), .Z(n51415) );
  XOR U60974 ( .A(n51392), .B(n51418), .Z(N60814) );
  XNOR U60975 ( .A(n51395), .B(n51394), .Z(n51418) );
  XNOR U60976 ( .A(n51406), .B(n51419), .Z(n51394) );
  XNOR U60977 ( .A(n51410), .B(n51408), .Z(n51419) );
  XOR U60978 ( .A(n51416), .B(n51420), .Z(n51408) );
  XNOR U60979 ( .A(n51413), .B(n51417), .Z(n51420) );
  AND U60980 ( .A(n51421), .B(n51422), .Z(n51417) );
  NAND U60981 ( .A(n51423), .B(n51424), .Z(n51422) );
  NAND U60982 ( .A(n51425), .B(n51426), .Z(n51421) );
  AND U60983 ( .A(n51427), .B(n51428), .Z(n51413) );
  NAND U60984 ( .A(n51429), .B(n51430), .Z(n51428) );
  NAND U60985 ( .A(n51431), .B(n51432), .Z(n51427) );
  NANDN U60986 ( .A(n51433), .B(n51434), .Z(n51416) );
  ANDN U60987 ( .B(n51435), .A(n51436), .Z(n51410) );
  XNOR U60988 ( .A(n51401), .B(n51437), .Z(n51406) );
  XNOR U60989 ( .A(n51399), .B(n51403), .Z(n51437) );
  AND U60990 ( .A(n51438), .B(n51439), .Z(n51403) );
  NAND U60991 ( .A(n51440), .B(n51441), .Z(n51439) );
  NAND U60992 ( .A(n51442), .B(n51443), .Z(n51438) );
  AND U60993 ( .A(n51444), .B(n51445), .Z(n51399) );
  NAND U60994 ( .A(n51446), .B(n51447), .Z(n51445) );
  NAND U60995 ( .A(n51448), .B(n51449), .Z(n51444) );
  AND U60996 ( .A(n51450), .B(n51451), .Z(n51401) );
  NAND U60997 ( .A(n51452), .B(n51453), .Z(n51395) );
  XNOR U60998 ( .A(n51378), .B(n51454), .Z(n51392) );
  XNOR U60999 ( .A(n51382), .B(n51380), .Z(n51454) );
  XOR U61000 ( .A(n51388), .B(n51455), .Z(n51380) );
  XNOR U61001 ( .A(n51385), .B(n51389), .Z(n51455) );
  AND U61002 ( .A(n51456), .B(n51457), .Z(n51389) );
  NAND U61003 ( .A(n51458), .B(n51459), .Z(n51457) );
  NAND U61004 ( .A(n51460), .B(n51461), .Z(n51456) );
  AND U61005 ( .A(n51462), .B(n51463), .Z(n51385) );
  NAND U61006 ( .A(n51464), .B(n51465), .Z(n51463) );
  NAND U61007 ( .A(n51466), .B(n51467), .Z(n51462) );
  NANDN U61008 ( .A(n51468), .B(n51469), .Z(n51388) );
  ANDN U61009 ( .B(n51470), .A(n51471), .Z(n51382) );
  XNOR U61010 ( .A(n51373), .B(n51472), .Z(n51378) );
  XNOR U61011 ( .A(n51371), .B(n51375), .Z(n51472) );
  AND U61012 ( .A(n51473), .B(n51474), .Z(n51375) );
  NAND U61013 ( .A(n51475), .B(n51476), .Z(n51474) );
  NAND U61014 ( .A(n51477), .B(n51478), .Z(n51473) );
  AND U61015 ( .A(n51479), .B(n51480), .Z(n51371) );
  NAND U61016 ( .A(n51481), .B(n51482), .Z(n51480) );
  NAND U61017 ( .A(n51483), .B(n51484), .Z(n51479) );
  AND U61018 ( .A(n51485), .B(n51486), .Z(n51373) );
  XOR U61019 ( .A(n51453), .B(n51452), .Z(N60813) );
  XNOR U61020 ( .A(n51470), .B(n51471), .Z(n51452) );
  XNOR U61021 ( .A(n51485), .B(n51486), .Z(n51471) );
  XOR U61022 ( .A(n51482), .B(n51481), .Z(n51486) );
  XOR U61023 ( .A(y[420]), .B(x[420]), .Z(n51481) );
  XOR U61024 ( .A(n51484), .B(n51483), .Z(n51482) );
  XOR U61025 ( .A(y[422]), .B(x[422]), .Z(n51483) );
  XOR U61026 ( .A(y[421]), .B(x[421]), .Z(n51484) );
  XOR U61027 ( .A(n51476), .B(n51475), .Z(n51485) );
  XOR U61028 ( .A(n51478), .B(n51477), .Z(n51475) );
  XOR U61029 ( .A(y[419]), .B(x[419]), .Z(n51477) );
  XOR U61030 ( .A(y[418]), .B(x[418]), .Z(n51478) );
  XOR U61031 ( .A(y[417]), .B(x[417]), .Z(n51476) );
  XNOR U61032 ( .A(n51469), .B(n51468), .Z(n51470) );
  XNOR U61033 ( .A(n51465), .B(n51464), .Z(n51468) );
  XOR U61034 ( .A(n51467), .B(n51466), .Z(n51464) );
  XOR U61035 ( .A(y[416]), .B(x[416]), .Z(n51466) );
  XOR U61036 ( .A(y[415]), .B(x[415]), .Z(n51467) );
  XOR U61037 ( .A(y[414]), .B(x[414]), .Z(n51465) );
  XOR U61038 ( .A(n51459), .B(n51458), .Z(n51469) );
  XOR U61039 ( .A(n51461), .B(n51460), .Z(n51458) );
  XOR U61040 ( .A(y[413]), .B(x[413]), .Z(n51460) );
  XOR U61041 ( .A(y[412]), .B(x[412]), .Z(n51461) );
  XOR U61042 ( .A(y[411]), .B(x[411]), .Z(n51459) );
  XNOR U61043 ( .A(n51435), .B(n51436), .Z(n51453) );
  XNOR U61044 ( .A(n51450), .B(n51451), .Z(n51436) );
  XOR U61045 ( .A(n51447), .B(n51446), .Z(n51451) );
  XOR U61046 ( .A(y[408]), .B(x[408]), .Z(n51446) );
  XOR U61047 ( .A(n51449), .B(n51448), .Z(n51447) );
  XOR U61048 ( .A(y[410]), .B(x[410]), .Z(n51448) );
  XOR U61049 ( .A(y[409]), .B(x[409]), .Z(n51449) );
  XOR U61050 ( .A(n51441), .B(n51440), .Z(n51450) );
  XOR U61051 ( .A(n51443), .B(n51442), .Z(n51440) );
  XOR U61052 ( .A(y[407]), .B(x[407]), .Z(n51442) );
  XOR U61053 ( .A(y[406]), .B(x[406]), .Z(n51443) );
  XOR U61054 ( .A(y[405]), .B(x[405]), .Z(n51441) );
  XNOR U61055 ( .A(n51434), .B(n51433), .Z(n51435) );
  XNOR U61056 ( .A(n51430), .B(n51429), .Z(n51433) );
  XOR U61057 ( .A(n51432), .B(n51431), .Z(n51429) );
  XOR U61058 ( .A(y[404]), .B(x[404]), .Z(n51431) );
  XOR U61059 ( .A(y[403]), .B(x[403]), .Z(n51432) );
  XOR U61060 ( .A(y[402]), .B(x[402]), .Z(n51430) );
  XOR U61061 ( .A(n51424), .B(n51423), .Z(n51434) );
  XOR U61062 ( .A(n51426), .B(n51425), .Z(n51423) );
  XOR U61063 ( .A(y[401]), .B(x[401]), .Z(n51425) );
  XOR U61064 ( .A(y[400]), .B(x[400]), .Z(n51426) );
  XOR U61065 ( .A(y[399]), .B(x[399]), .Z(n51424) );
  NAND U61066 ( .A(n51487), .B(n51488), .Z(N60804) );
  NAND U61067 ( .A(n51489), .B(n51490), .Z(n51488) );
  NANDN U61068 ( .A(n51491), .B(n51492), .Z(n51490) );
  NANDN U61069 ( .A(n51492), .B(n51491), .Z(n51487) );
  XOR U61070 ( .A(n51491), .B(n51493), .Z(N60803) );
  XNOR U61071 ( .A(n51489), .B(n51492), .Z(n51493) );
  NAND U61072 ( .A(n51494), .B(n51495), .Z(n51492) );
  NAND U61073 ( .A(n51496), .B(n51497), .Z(n51495) );
  NANDN U61074 ( .A(n51498), .B(n51499), .Z(n51497) );
  NANDN U61075 ( .A(n51499), .B(n51498), .Z(n51494) );
  AND U61076 ( .A(n51500), .B(n51501), .Z(n51489) );
  NAND U61077 ( .A(n51502), .B(n51503), .Z(n51501) );
  NANDN U61078 ( .A(n51504), .B(n51505), .Z(n51503) );
  NANDN U61079 ( .A(n51505), .B(n51504), .Z(n51500) );
  IV U61080 ( .A(n51506), .Z(n51505) );
  AND U61081 ( .A(n51507), .B(n51508), .Z(n51491) );
  NAND U61082 ( .A(n51509), .B(n51510), .Z(n51508) );
  NANDN U61083 ( .A(n51511), .B(n51512), .Z(n51510) );
  NANDN U61084 ( .A(n51512), .B(n51511), .Z(n51507) );
  XOR U61085 ( .A(n51504), .B(n51513), .Z(N60802) );
  XNOR U61086 ( .A(n51502), .B(n51506), .Z(n51513) );
  XOR U61087 ( .A(n51499), .B(n51514), .Z(n51506) );
  XNOR U61088 ( .A(n51496), .B(n51498), .Z(n51514) );
  AND U61089 ( .A(n51515), .B(n51516), .Z(n51498) );
  NANDN U61090 ( .A(n51517), .B(n51518), .Z(n51516) );
  OR U61091 ( .A(n51519), .B(n51520), .Z(n51518) );
  IV U61092 ( .A(n51521), .Z(n51520) );
  NANDN U61093 ( .A(n51521), .B(n51519), .Z(n51515) );
  AND U61094 ( .A(n51522), .B(n51523), .Z(n51496) );
  NAND U61095 ( .A(n51524), .B(n51525), .Z(n51523) );
  NANDN U61096 ( .A(n51526), .B(n51527), .Z(n51525) );
  NANDN U61097 ( .A(n51527), .B(n51526), .Z(n51522) );
  IV U61098 ( .A(n51528), .Z(n51527) );
  NAND U61099 ( .A(n51529), .B(n51530), .Z(n51499) );
  NANDN U61100 ( .A(n51531), .B(n51532), .Z(n51530) );
  NANDN U61101 ( .A(n51533), .B(n51534), .Z(n51532) );
  NANDN U61102 ( .A(n51534), .B(n51533), .Z(n51529) );
  IV U61103 ( .A(n51535), .Z(n51533) );
  AND U61104 ( .A(n51536), .B(n51537), .Z(n51502) );
  NAND U61105 ( .A(n51538), .B(n51539), .Z(n51537) );
  NANDN U61106 ( .A(n51540), .B(n51541), .Z(n51539) );
  NANDN U61107 ( .A(n51541), .B(n51540), .Z(n51536) );
  XOR U61108 ( .A(n51512), .B(n51542), .Z(n51504) );
  XNOR U61109 ( .A(n51509), .B(n51511), .Z(n51542) );
  AND U61110 ( .A(n51543), .B(n51544), .Z(n51511) );
  NANDN U61111 ( .A(n51545), .B(n51546), .Z(n51544) );
  OR U61112 ( .A(n51547), .B(n51548), .Z(n51546) );
  IV U61113 ( .A(n51549), .Z(n51548) );
  NANDN U61114 ( .A(n51549), .B(n51547), .Z(n51543) );
  AND U61115 ( .A(n51550), .B(n51551), .Z(n51509) );
  NAND U61116 ( .A(n51552), .B(n51553), .Z(n51551) );
  NANDN U61117 ( .A(n51554), .B(n51555), .Z(n51553) );
  NANDN U61118 ( .A(n51555), .B(n51554), .Z(n51550) );
  IV U61119 ( .A(n51556), .Z(n51555) );
  NAND U61120 ( .A(n51557), .B(n51558), .Z(n51512) );
  NANDN U61121 ( .A(n51559), .B(n51560), .Z(n51558) );
  NANDN U61122 ( .A(n51561), .B(n51562), .Z(n51560) );
  NANDN U61123 ( .A(n51562), .B(n51561), .Z(n51557) );
  IV U61124 ( .A(n51563), .Z(n51561) );
  XOR U61125 ( .A(n51538), .B(n51564), .Z(N60801) );
  XNOR U61126 ( .A(n51541), .B(n51540), .Z(n51564) );
  XNOR U61127 ( .A(n51552), .B(n51565), .Z(n51540) );
  XNOR U61128 ( .A(n51556), .B(n51554), .Z(n51565) );
  XOR U61129 ( .A(n51562), .B(n51566), .Z(n51554) );
  XNOR U61130 ( .A(n51559), .B(n51563), .Z(n51566) );
  AND U61131 ( .A(n51567), .B(n51568), .Z(n51563) );
  NAND U61132 ( .A(n51569), .B(n51570), .Z(n51568) );
  NAND U61133 ( .A(n51571), .B(n51572), .Z(n51567) );
  AND U61134 ( .A(n51573), .B(n51574), .Z(n51559) );
  NAND U61135 ( .A(n51575), .B(n51576), .Z(n51574) );
  NAND U61136 ( .A(n51577), .B(n51578), .Z(n51573) );
  NANDN U61137 ( .A(n51579), .B(n51580), .Z(n51562) );
  ANDN U61138 ( .B(n51581), .A(n51582), .Z(n51556) );
  XNOR U61139 ( .A(n51547), .B(n51583), .Z(n51552) );
  XNOR U61140 ( .A(n51545), .B(n51549), .Z(n51583) );
  AND U61141 ( .A(n51584), .B(n51585), .Z(n51549) );
  NAND U61142 ( .A(n51586), .B(n51587), .Z(n51585) );
  NAND U61143 ( .A(n51588), .B(n51589), .Z(n51584) );
  AND U61144 ( .A(n51590), .B(n51591), .Z(n51545) );
  NAND U61145 ( .A(n51592), .B(n51593), .Z(n51591) );
  NAND U61146 ( .A(n51594), .B(n51595), .Z(n51590) );
  AND U61147 ( .A(n51596), .B(n51597), .Z(n51547) );
  NAND U61148 ( .A(n51598), .B(n51599), .Z(n51541) );
  XNOR U61149 ( .A(n51524), .B(n51600), .Z(n51538) );
  XNOR U61150 ( .A(n51528), .B(n51526), .Z(n51600) );
  XOR U61151 ( .A(n51534), .B(n51601), .Z(n51526) );
  XNOR U61152 ( .A(n51531), .B(n51535), .Z(n51601) );
  AND U61153 ( .A(n51602), .B(n51603), .Z(n51535) );
  NAND U61154 ( .A(n51604), .B(n51605), .Z(n51603) );
  NAND U61155 ( .A(n51606), .B(n51607), .Z(n51602) );
  AND U61156 ( .A(n51608), .B(n51609), .Z(n51531) );
  NAND U61157 ( .A(n51610), .B(n51611), .Z(n51609) );
  NAND U61158 ( .A(n51612), .B(n51613), .Z(n51608) );
  NANDN U61159 ( .A(n51614), .B(n51615), .Z(n51534) );
  ANDN U61160 ( .B(n51616), .A(n51617), .Z(n51528) );
  XNOR U61161 ( .A(n51519), .B(n51618), .Z(n51524) );
  XNOR U61162 ( .A(n51517), .B(n51521), .Z(n51618) );
  AND U61163 ( .A(n51619), .B(n51620), .Z(n51521) );
  NAND U61164 ( .A(n51621), .B(n51622), .Z(n51620) );
  NAND U61165 ( .A(n51623), .B(n51624), .Z(n51619) );
  AND U61166 ( .A(n51625), .B(n51626), .Z(n51517) );
  NAND U61167 ( .A(n51627), .B(n51628), .Z(n51626) );
  NAND U61168 ( .A(n51629), .B(n51630), .Z(n51625) );
  AND U61169 ( .A(n51631), .B(n51632), .Z(n51519) );
  XOR U61170 ( .A(n51599), .B(n51598), .Z(N60800) );
  XNOR U61171 ( .A(n51616), .B(n51617), .Z(n51598) );
  XNOR U61172 ( .A(n51631), .B(n51632), .Z(n51617) );
  XOR U61173 ( .A(n51628), .B(n51627), .Z(n51632) );
  XOR U61174 ( .A(y[396]), .B(x[396]), .Z(n51627) );
  XOR U61175 ( .A(n51630), .B(n51629), .Z(n51628) );
  XOR U61176 ( .A(y[398]), .B(x[398]), .Z(n51629) );
  XOR U61177 ( .A(y[397]), .B(x[397]), .Z(n51630) );
  XOR U61178 ( .A(n51622), .B(n51621), .Z(n51631) );
  XOR U61179 ( .A(n51624), .B(n51623), .Z(n51621) );
  XOR U61180 ( .A(y[395]), .B(x[395]), .Z(n51623) );
  XOR U61181 ( .A(y[394]), .B(x[394]), .Z(n51624) );
  XOR U61182 ( .A(y[393]), .B(x[393]), .Z(n51622) );
  XNOR U61183 ( .A(n51615), .B(n51614), .Z(n51616) );
  XNOR U61184 ( .A(n51611), .B(n51610), .Z(n51614) );
  XOR U61185 ( .A(n51613), .B(n51612), .Z(n51610) );
  XOR U61186 ( .A(y[392]), .B(x[392]), .Z(n51612) );
  XOR U61187 ( .A(y[391]), .B(x[391]), .Z(n51613) );
  XOR U61188 ( .A(y[390]), .B(x[390]), .Z(n51611) );
  XOR U61189 ( .A(n51605), .B(n51604), .Z(n51615) );
  XOR U61190 ( .A(n51607), .B(n51606), .Z(n51604) );
  XOR U61191 ( .A(y[389]), .B(x[389]), .Z(n51606) );
  XOR U61192 ( .A(y[388]), .B(x[388]), .Z(n51607) );
  XOR U61193 ( .A(y[387]), .B(x[387]), .Z(n51605) );
  XNOR U61194 ( .A(n51581), .B(n51582), .Z(n51599) );
  XNOR U61195 ( .A(n51596), .B(n51597), .Z(n51582) );
  XOR U61196 ( .A(n51593), .B(n51592), .Z(n51597) );
  XOR U61197 ( .A(y[384]), .B(x[384]), .Z(n51592) );
  XOR U61198 ( .A(n51595), .B(n51594), .Z(n51593) );
  XOR U61199 ( .A(y[386]), .B(x[386]), .Z(n51594) );
  XOR U61200 ( .A(y[385]), .B(x[385]), .Z(n51595) );
  XOR U61201 ( .A(n51587), .B(n51586), .Z(n51596) );
  XOR U61202 ( .A(n51589), .B(n51588), .Z(n51586) );
  XOR U61203 ( .A(y[383]), .B(x[383]), .Z(n51588) );
  XOR U61204 ( .A(y[382]), .B(x[382]), .Z(n51589) );
  XOR U61205 ( .A(y[381]), .B(x[381]), .Z(n51587) );
  XNOR U61206 ( .A(n51580), .B(n51579), .Z(n51581) );
  XNOR U61207 ( .A(n51576), .B(n51575), .Z(n51579) );
  XOR U61208 ( .A(n51578), .B(n51577), .Z(n51575) );
  XOR U61209 ( .A(y[380]), .B(x[380]), .Z(n51577) );
  XOR U61210 ( .A(y[379]), .B(x[379]), .Z(n51578) );
  XOR U61211 ( .A(y[378]), .B(x[378]), .Z(n51576) );
  XOR U61212 ( .A(n51570), .B(n51569), .Z(n51580) );
  XOR U61213 ( .A(n51572), .B(n51571), .Z(n51569) );
  XOR U61214 ( .A(y[377]), .B(x[377]), .Z(n51571) );
  XOR U61215 ( .A(y[376]), .B(x[376]), .Z(n51572) );
  XOR U61216 ( .A(y[375]), .B(x[375]), .Z(n51570) );
  NAND U61217 ( .A(n51633), .B(n51634), .Z(N60791) );
  NAND U61218 ( .A(n51635), .B(n51636), .Z(n51634) );
  NANDN U61219 ( .A(n51637), .B(n51638), .Z(n51636) );
  NANDN U61220 ( .A(n51638), .B(n51637), .Z(n51633) );
  XOR U61221 ( .A(n51637), .B(n51639), .Z(N60790) );
  XNOR U61222 ( .A(n51635), .B(n51638), .Z(n51639) );
  NAND U61223 ( .A(n51640), .B(n51641), .Z(n51638) );
  NAND U61224 ( .A(n51642), .B(n51643), .Z(n51641) );
  NANDN U61225 ( .A(n51644), .B(n51645), .Z(n51643) );
  NANDN U61226 ( .A(n51645), .B(n51644), .Z(n51640) );
  AND U61227 ( .A(n51646), .B(n51647), .Z(n51635) );
  NAND U61228 ( .A(n51648), .B(n51649), .Z(n51647) );
  NANDN U61229 ( .A(n51650), .B(n51651), .Z(n51649) );
  NANDN U61230 ( .A(n51651), .B(n51650), .Z(n51646) );
  IV U61231 ( .A(n51652), .Z(n51651) );
  AND U61232 ( .A(n51653), .B(n51654), .Z(n51637) );
  NAND U61233 ( .A(n51655), .B(n51656), .Z(n51654) );
  NANDN U61234 ( .A(n51657), .B(n51658), .Z(n51656) );
  NANDN U61235 ( .A(n51658), .B(n51657), .Z(n51653) );
  XOR U61236 ( .A(n51650), .B(n51659), .Z(N60789) );
  XNOR U61237 ( .A(n51648), .B(n51652), .Z(n51659) );
  XOR U61238 ( .A(n51645), .B(n51660), .Z(n51652) );
  XNOR U61239 ( .A(n51642), .B(n51644), .Z(n51660) );
  AND U61240 ( .A(n51661), .B(n51662), .Z(n51644) );
  NANDN U61241 ( .A(n51663), .B(n51664), .Z(n51662) );
  OR U61242 ( .A(n51665), .B(n51666), .Z(n51664) );
  IV U61243 ( .A(n51667), .Z(n51666) );
  NANDN U61244 ( .A(n51667), .B(n51665), .Z(n51661) );
  AND U61245 ( .A(n51668), .B(n51669), .Z(n51642) );
  NAND U61246 ( .A(n51670), .B(n51671), .Z(n51669) );
  NANDN U61247 ( .A(n51672), .B(n51673), .Z(n51671) );
  NANDN U61248 ( .A(n51673), .B(n51672), .Z(n51668) );
  IV U61249 ( .A(n51674), .Z(n51673) );
  NAND U61250 ( .A(n51675), .B(n51676), .Z(n51645) );
  NANDN U61251 ( .A(n51677), .B(n51678), .Z(n51676) );
  NANDN U61252 ( .A(n51679), .B(n51680), .Z(n51678) );
  NANDN U61253 ( .A(n51680), .B(n51679), .Z(n51675) );
  IV U61254 ( .A(n51681), .Z(n51679) );
  AND U61255 ( .A(n51682), .B(n51683), .Z(n51648) );
  NAND U61256 ( .A(n51684), .B(n51685), .Z(n51683) );
  NANDN U61257 ( .A(n51686), .B(n51687), .Z(n51685) );
  NANDN U61258 ( .A(n51687), .B(n51686), .Z(n51682) );
  XOR U61259 ( .A(n51658), .B(n51688), .Z(n51650) );
  XNOR U61260 ( .A(n51655), .B(n51657), .Z(n51688) );
  AND U61261 ( .A(n51689), .B(n51690), .Z(n51657) );
  NANDN U61262 ( .A(n51691), .B(n51692), .Z(n51690) );
  OR U61263 ( .A(n51693), .B(n51694), .Z(n51692) );
  IV U61264 ( .A(n51695), .Z(n51694) );
  NANDN U61265 ( .A(n51695), .B(n51693), .Z(n51689) );
  AND U61266 ( .A(n51696), .B(n51697), .Z(n51655) );
  NAND U61267 ( .A(n51698), .B(n51699), .Z(n51697) );
  NANDN U61268 ( .A(n51700), .B(n51701), .Z(n51699) );
  NANDN U61269 ( .A(n51701), .B(n51700), .Z(n51696) );
  IV U61270 ( .A(n51702), .Z(n51701) );
  NAND U61271 ( .A(n51703), .B(n51704), .Z(n51658) );
  NANDN U61272 ( .A(n51705), .B(n51706), .Z(n51704) );
  NANDN U61273 ( .A(n51707), .B(n51708), .Z(n51706) );
  NANDN U61274 ( .A(n51708), .B(n51707), .Z(n51703) );
  IV U61275 ( .A(n51709), .Z(n51707) );
  XOR U61276 ( .A(n51684), .B(n51710), .Z(N60788) );
  XNOR U61277 ( .A(n51687), .B(n51686), .Z(n51710) );
  XNOR U61278 ( .A(n51698), .B(n51711), .Z(n51686) );
  XNOR U61279 ( .A(n51702), .B(n51700), .Z(n51711) );
  XOR U61280 ( .A(n51708), .B(n51712), .Z(n51700) );
  XNOR U61281 ( .A(n51705), .B(n51709), .Z(n51712) );
  AND U61282 ( .A(n51713), .B(n51714), .Z(n51709) );
  NAND U61283 ( .A(n51715), .B(n51716), .Z(n51714) );
  NAND U61284 ( .A(n51717), .B(n51718), .Z(n51713) );
  AND U61285 ( .A(n51719), .B(n51720), .Z(n51705) );
  NAND U61286 ( .A(n51721), .B(n51722), .Z(n51720) );
  NAND U61287 ( .A(n51723), .B(n51724), .Z(n51719) );
  NANDN U61288 ( .A(n51725), .B(n51726), .Z(n51708) );
  ANDN U61289 ( .B(n51727), .A(n51728), .Z(n51702) );
  XNOR U61290 ( .A(n51693), .B(n51729), .Z(n51698) );
  XNOR U61291 ( .A(n51691), .B(n51695), .Z(n51729) );
  AND U61292 ( .A(n51730), .B(n51731), .Z(n51695) );
  NAND U61293 ( .A(n51732), .B(n51733), .Z(n51731) );
  NAND U61294 ( .A(n51734), .B(n51735), .Z(n51730) );
  AND U61295 ( .A(n51736), .B(n51737), .Z(n51691) );
  NAND U61296 ( .A(n51738), .B(n51739), .Z(n51737) );
  NAND U61297 ( .A(n51740), .B(n51741), .Z(n51736) );
  AND U61298 ( .A(n51742), .B(n51743), .Z(n51693) );
  NAND U61299 ( .A(n51744), .B(n51745), .Z(n51687) );
  XNOR U61300 ( .A(n51670), .B(n51746), .Z(n51684) );
  XNOR U61301 ( .A(n51674), .B(n51672), .Z(n51746) );
  XOR U61302 ( .A(n51680), .B(n51747), .Z(n51672) );
  XNOR U61303 ( .A(n51677), .B(n51681), .Z(n51747) );
  AND U61304 ( .A(n51748), .B(n51749), .Z(n51681) );
  NAND U61305 ( .A(n51750), .B(n51751), .Z(n51749) );
  NAND U61306 ( .A(n51752), .B(n51753), .Z(n51748) );
  AND U61307 ( .A(n51754), .B(n51755), .Z(n51677) );
  NAND U61308 ( .A(n51756), .B(n51757), .Z(n51755) );
  NAND U61309 ( .A(n51758), .B(n51759), .Z(n51754) );
  NANDN U61310 ( .A(n51760), .B(n51761), .Z(n51680) );
  ANDN U61311 ( .B(n51762), .A(n51763), .Z(n51674) );
  XNOR U61312 ( .A(n51665), .B(n51764), .Z(n51670) );
  XNOR U61313 ( .A(n51663), .B(n51667), .Z(n51764) );
  AND U61314 ( .A(n51765), .B(n51766), .Z(n51667) );
  NAND U61315 ( .A(n51767), .B(n51768), .Z(n51766) );
  NAND U61316 ( .A(n51769), .B(n51770), .Z(n51765) );
  AND U61317 ( .A(n51771), .B(n51772), .Z(n51663) );
  NAND U61318 ( .A(n51773), .B(n51774), .Z(n51772) );
  NAND U61319 ( .A(n51775), .B(n51776), .Z(n51771) );
  AND U61320 ( .A(n51777), .B(n51778), .Z(n51665) );
  XOR U61321 ( .A(n51745), .B(n51744), .Z(N60787) );
  XNOR U61322 ( .A(n51762), .B(n51763), .Z(n51744) );
  XNOR U61323 ( .A(n51777), .B(n51778), .Z(n51763) );
  XOR U61324 ( .A(n51774), .B(n51773), .Z(n51778) );
  XOR U61325 ( .A(y[372]), .B(x[372]), .Z(n51773) );
  XOR U61326 ( .A(n51776), .B(n51775), .Z(n51774) );
  XOR U61327 ( .A(y[374]), .B(x[374]), .Z(n51775) );
  XOR U61328 ( .A(y[373]), .B(x[373]), .Z(n51776) );
  XOR U61329 ( .A(n51768), .B(n51767), .Z(n51777) );
  XOR U61330 ( .A(n51770), .B(n51769), .Z(n51767) );
  XOR U61331 ( .A(y[371]), .B(x[371]), .Z(n51769) );
  XOR U61332 ( .A(y[370]), .B(x[370]), .Z(n51770) );
  XOR U61333 ( .A(y[369]), .B(x[369]), .Z(n51768) );
  XNOR U61334 ( .A(n51761), .B(n51760), .Z(n51762) );
  XNOR U61335 ( .A(n51757), .B(n51756), .Z(n51760) );
  XOR U61336 ( .A(n51759), .B(n51758), .Z(n51756) );
  XOR U61337 ( .A(y[368]), .B(x[368]), .Z(n51758) );
  XOR U61338 ( .A(y[367]), .B(x[367]), .Z(n51759) );
  XOR U61339 ( .A(y[366]), .B(x[366]), .Z(n51757) );
  XOR U61340 ( .A(n51751), .B(n51750), .Z(n51761) );
  XOR U61341 ( .A(n51753), .B(n51752), .Z(n51750) );
  XOR U61342 ( .A(y[365]), .B(x[365]), .Z(n51752) );
  XOR U61343 ( .A(y[364]), .B(x[364]), .Z(n51753) );
  XOR U61344 ( .A(y[363]), .B(x[363]), .Z(n51751) );
  XNOR U61345 ( .A(n51727), .B(n51728), .Z(n51745) );
  XNOR U61346 ( .A(n51742), .B(n51743), .Z(n51728) );
  XOR U61347 ( .A(n51739), .B(n51738), .Z(n51743) );
  XOR U61348 ( .A(y[360]), .B(x[360]), .Z(n51738) );
  XOR U61349 ( .A(n51741), .B(n51740), .Z(n51739) );
  XOR U61350 ( .A(y[362]), .B(x[362]), .Z(n51740) );
  XOR U61351 ( .A(y[361]), .B(x[361]), .Z(n51741) );
  XOR U61352 ( .A(n51733), .B(n51732), .Z(n51742) );
  XOR U61353 ( .A(n51735), .B(n51734), .Z(n51732) );
  XOR U61354 ( .A(y[359]), .B(x[359]), .Z(n51734) );
  XOR U61355 ( .A(y[358]), .B(x[358]), .Z(n51735) );
  XOR U61356 ( .A(y[357]), .B(x[357]), .Z(n51733) );
  XNOR U61357 ( .A(n51726), .B(n51725), .Z(n51727) );
  XNOR U61358 ( .A(n51722), .B(n51721), .Z(n51725) );
  XOR U61359 ( .A(n51724), .B(n51723), .Z(n51721) );
  XOR U61360 ( .A(y[356]), .B(x[356]), .Z(n51723) );
  XOR U61361 ( .A(y[355]), .B(x[355]), .Z(n51724) );
  XOR U61362 ( .A(y[354]), .B(x[354]), .Z(n51722) );
  XOR U61363 ( .A(n51716), .B(n51715), .Z(n51726) );
  XOR U61364 ( .A(n51718), .B(n51717), .Z(n51715) );
  XOR U61365 ( .A(y[353]), .B(x[353]), .Z(n51717) );
  XOR U61366 ( .A(y[352]), .B(x[352]), .Z(n51718) );
  XOR U61367 ( .A(y[351]), .B(x[351]), .Z(n51716) );
  NAND U61368 ( .A(n51779), .B(n51780), .Z(N60778) );
  NAND U61369 ( .A(n51781), .B(n51782), .Z(n51780) );
  NANDN U61370 ( .A(n51783), .B(n51784), .Z(n51782) );
  NANDN U61371 ( .A(n51784), .B(n51783), .Z(n51779) );
  XOR U61372 ( .A(n51783), .B(n51785), .Z(N60777) );
  XNOR U61373 ( .A(n51781), .B(n51784), .Z(n51785) );
  NAND U61374 ( .A(n51786), .B(n51787), .Z(n51784) );
  NAND U61375 ( .A(n51788), .B(n51789), .Z(n51787) );
  NANDN U61376 ( .A(n51790), .B(n51791), .Z(n51789) );
  NANDN U61377 ( .A(n51791), .B(n51790), .Z(n51786) );
  AND U61378 ( .A(n51792), .B(n51793), .Z(n51781) );
  NAND U61379 ( .A(n51794), .B(n51795), .Z(n51793) );
  NANDN U61380 ( .A(n51796), .B(n51797), .Z(n51795) );
  NANDN U61381 ( .A(n51797), .B(n51796), .Z(n51792) );
  IV U61382 ( .A(n51798), .Z(n51797) );
  AND U61383 ( .A(n51799), .B(n51800), .Z(n51783) );
  NAND U61384 ( .A(n51801), .B(n51802), .Z(n51800) );
  NANDN U61385 ( .A(n51803), .B(n51804), .Z(n51802) );
  NANDN U61386 ( .A(n51804), .B(n51803), .Z(n51799) );
  XOR U61387 ( .A(n51796), .B(n51805), .Z(N60776) );
  XNOR U61388 ( .A(n51794), .B(n51798), .Z(n51805) );
  XOR U61389 ( .A(n51791), .B(n51806), .Z(n51798) );
  XNOR U61390 ( .A(n51788), .B(n51790), .Z(n51806) );
  AND U61391 ( .A(n51807), .B(n51808), .Z(n51790) );
  NANDN U61392 ( .A(n51809), .B(n51810), .Z(n51808) );
  OR U61393 ( .A(n51811), .B(n51812), .Z(n51810) );
  IV U61394 ( .A(n51813), .Z(n51812) );
  NANDN U61395 ( .A(n51813), .B(n51811), .Z(n51807) );
  AND U61396 ( .A(n51814), .B(n51815), .Z(n51788) );
  NAND U61397 ( .A(n51816), .B(n51817), .Z(n51815) );
  NANDN U61398 ( .A(n51818), .B(n51819), .Z(n51817) );
  NANDN U61399 ( .A(n51819), .B(n51818), .Z(n51814) );
  IV U61400 ( .A(n51820), .Z(n51819) );
  NAND U61401 ( .A(n51821), .B(n51822), .Z(n51791) );
  NANDN U61402 ( .A(n51823), .B(n51824), .Z(n51822) );
  NANDN U61403 ( .A(n51825), .B(n51826), .Z(n51824) );
  NANDN U61404 ( .A(n51826), .B(n51825), .Z(n51821) );
  IV U61405 ( .A(n51827), .Z(n51825) );
  AND U61406 ( .A(n51828), .B(n51829), .Z(n51794) );
  NAND U61407 ( .A(n51830), .B(n51831), .Z(n51829) );
  NANDN U61408 ( .A(n51832), .B(n51833), .Z(n51831) );
  NANDN U61409 ( .A(n51833), .B(n51832), .Z(n51828) );
  XOR U61410 ( .A(n51804), .B(n51834), .Z(n51796) );
  XNOR U61411 ( .A(n51801), .B(n51803), .Z(n51834) );
  AND U61412 ( .A(n51835), .B(n51836), .Z(n51803) );
  NANDN U61413 ( .A(n51837), .B(n51838), .Z(n51836) );
  OR U61414 ( .A(n51839), .B(n51840), .Z(n51838) );
  IV U61415 ( .A(n51841), .Z(n51840) );
  NANDN U61416 ( .A(n51841), .B(n51839), .Z(n51835) );
  AND U61417 ( .A(n51842), .B(n51843), .Z(n51801) );
  NAND U61418 ( .A(n51844), .B(n51845), .Z(n51843) );
  NANDN U61419 ( .A(n51846), .B(n51847), .Z(n51845) );
  NANDN U61420 ( .A(n51847), .B(n51846), .Z(n51842) );
  IV U61421 ( .A(n51848), .Z(n51847) );
  NAND U61422 ( .A(n51849), .B(n51850), .Z(n51804) );
  NANDN U61423 ( .A(n51851), .B(n51852), .Z(n51850) );
  NANDN U61424 ( .A(n51853), .B(n51854), .Z(n51852) );
  NANDN U61425 ( .A(n51854), .B(n51853), .Z(n51849) );
  IV U61426 ( .A(n51855), .Z(n51853) );
  XOR U61427 ( .A(n51830), .B(n51856), .Z(N60775) );
  XNOR U61428 ( .A(n51833), .B(n51832), .Z(n51856) );
  XNOR U61429 ( .A(n51844), .B(n51857), .Z(n51832) );
  XNOR U61430 ( .A(n51848), .B(n51846), .Z(n51857) );
  XOR U61431 ( .A(n51854), .B(n51858), .Z(n51846) );
  XNOR U61432 ( .A(n51851), .B(n51855), .Z(n51858) );
  AND U61433 ( .A(n51859), .B(n51860), .Z(n51855) );
  NAND U61434 ( .A(n51861), .B(n51862), .Z(n51860) );
  NAND U61435 ( .A(n51863), .B(n51864), .Z(n51859) );
  AND U61436 ( .A(n51865), .B(n51866), .Z(n51851) );
  NAND U61437 ( .A(n51867), .B(n51868), .Z(n51866) );
  NAND U61438 ( .A(n51869), .B(n51870), .Z(n51865) );
  NANDN U61439 ( .A(n51871), .B(n51872), .Z(n51854) );
  ANDN U61440 ( .B(n51873), .A(n51874), .Z(n51848) );
  XNOR U61441 ( .A(n51839), .B(n51875), .Z(n51844) );
  XNOR U61442 ( .A(n51837), .B(n51841), .Z(n51875) );
  AND U61443 ( .A(n51876), .B(n51877), .Z(n51841) );
  NAND U61444 ( .A(n51878), .B(n51879), .Z(n51877) );
  NAND U61445 ( .A(n51880), .B(n51881), .Z(n51876) );
  AND U61446 ( .A(n51882), .B(n51883), .Z(n51837) );
  NAND U61447 ( .A(n51884), .B(n51885), .Z(n51883) );
  NAND U61448 ( .A(n51886), .B(n51887), .Z(n51882) );
  AND U61449 ( .A(n51888), .B(n51889), .Z(n51839) );
  NAND U61450 ( .A(n51890), .B(n51891), .Z(n51833) );
  XNOR U61451 ( .A(n51816), .B(n51892), .Z(n51830) );
  XNOR U61452 ( .A(n51820), .B(n51818), .Z(n51892) );
  XOR U61453 ( .A(n51826), .B(n51893), .Z(n51818) );
  XNOR U61454 ( .A(n51823), .B(n51827), .Z(n51893) );
  AND U61455 ( .A(n51894), .B(n51895), .Z(n51827) );
  NAND U61456 ( .A(n51896), .B(n51897), .Z(n51895) );
  NAND U61457 ( .A(n51898), .B(n51899), .Z(n51894) );
  AND U61458 ( .A(n51900), .B(n51901), .Z(n51823) );
  NAND U61459 ( .A(n51902), .B(n51903), .Z(n51901) );
  NAND U61460 ( .A(n51904), .B(n51905), .Z(n51900) );
  NANDN U61461 ( .A(n51906), .B(n51907), .Z(n51826) );
  ANDN U61462 ( .B(n51908), .A(n51909), .Z(n51820) );
  XNOR U61463 ( .A(n51811), .B(n51910), .Z(n51816) );
  XNOR U61464 ( .A(n51809), .B(n51813), .Z(n51910) );
  AND U61465 ( .A(n51911), .B(n51912), .Z(n51813) );
  NAND U61466 ( .A(n51913), .B(n51914), .Z(n51912) );
  NAND U61467 ( .A(n51915), .B(n51916), .Z(n51911) );
  AND U61468 ( .A(n51917), .B(n51918), .Z(n51809) );
  NAND U61469 ( .A(n51919), .B(n51920), .Z(n51918) );
  NAND U61470 ( .A(n51921), .B(n51922), .Z(n51917) );
  AND U61471 ( .A(n51923), .B(n51924), .Z(n51811) );
  XOR U61472 ( .A(n51891), .B(n51890), .Z(N60774) );
  XNOR U61473 ( .A(n51908), .B(n51909), .Z(n51890) );
  XNOR U61474 ( .A(n51923), .B(n51924), .Z(n51909) );
  XOR U61475 ( .A(n51920), .B(n51919), .Z(n51924) );
  XOR U61476 ( .A(y[348]), .B(x[348]), .Z(n51919) );
  XOR U61477 ( .A(n51922), .B(n51921), .Z(n51920) );
  XOR U61478 ( .A(y[350]), .B(x[350]), .Z(n51921) );
  XOR U61479 ( .A(y[349]), .B(x[349]), .Z(n51922) );
  XOR U61480 ( .A(n51914), .B(n51913), .Z(n51923) );
  XOR U61481 ( .A(n51916), .B(n51915), .Z(n51913) );
  XOR U61482 ( .A(y[347]), .B(x[347]), .Z(n51915) );
  XOR U61483 ( .A(y[346]), .B(x[346]), .Z(n51916) );
  XOR U61484 ( .A(y[345]), .B(x[345]), .Z(n51914) );
  XNOR U61485 ( .A(n51907), .B(n51906), .Z(n51908) );
  XNOR U61486 ( .A(n51903), .B(n51902), .Z(n51906) );
  XOR U61487 ( .A(n51905), .B(n51904), .Z(n51902) );
  XOR U61488 ( .A(y[344]), .B(x[344]), .Z(n51904) );
  XOR U61489 ( .A(y[343]), .B(x[343]), .Z(n51905) );
  XOR U61490 ( .A(y[342]), .B(x[342]), .Z(n51903) );
  XOR U61491 ( .A(n51897), .B(n51896), .Z(n51907) );
  XOR U61492 ( .A(n51899), .B(n51898), .Z(n51896) );
  XOR U61493 ( .A(y[341]), .B(x[341]), .Z(n51898) );
  XOR U61494 ( .A(y[340]), .B(x[340]), .Z(n51899) );
  XOR U61495 ( .A(y[339]), .B(x[339]), .Z(n51897) );
  XNOR U61496 ( .A(n51873), .B(n51874), .Z(n51891) );
  XNOR U61497 ( .A(n51888), .B(n51889), .Z(n51874) );
  XOR U61498 ( .A(n51885), .B(n51884), .Z(n51889) );
  XOR U61499 ( .A(y[336]), .B(x[336]), .Z(n51884) );
  XOR U61500 ( .A(n51887), .B(n51886), .Z(n51885) );
  XOR U61501 ( .A(y[338]), .B(x[338]), .Z(n51886) );
  XOR U61502 ( .A(y[337]), .B(x[337]), .Z(n51887) );
  XOR U61503 ( .A(n51879), .B(n51878), .Z(n51888) );
  XOR U61504 ( .A(n51881), .B(n51880), .Z(n51878) );
  XOR U61505 ( .A(y[335]), .B(x[335]), .Z(n51880) );
  XOR U61506 ( .A(y[334]), .B(x[334]), .Z(n51881) );
  XOR U61507 ( .A(y[333]), .B(x[333]), .Z(n51879) );
  XNOR U61508 ( .A(n51872), .B(n51871), .Z(n51873) );
  XNOR U61509 ( .A(n51868), .B(n51867), .Z(n51871) );
  XOR U61510 ( .A(n51870), .B(n51869), .Z(n51867) );
  XOR U61511 ( .A(y[332]), .B(x[332]), .Z(n51869) );
  XOR U61512 ( .A(y[331]), .B(x[331]), .Z(n51870) );
  XOR U61513 ( .A(y[330]), .B(x[330]), .Z(n51868) );
  XOR U61514 ( .A(n51862), .B(n51861), .Z(n51872) );
  XOR U61515 ( .A(n51864), .B(n51863), .Z(n51861) );
  XOR U61516 ( .A(y[329]), .B(x[329]), .Z(n51863) );
  XOR U61517 ( .A(y[328]), .B(x[328]), .Z(n51864) );
  XOR U61518 ( .A(y[327]), .B(x[327]), .Z(n51862) );
  NAND U61519 ( .A(n51925), .B(n51926), .Z(N60765) );
  NAND U61520 ( .A(n51927), .B(n51928), .Z(n51926) );
  NANDN U61521 ( .A(n51929), .B(n51930), .Z(n51928) );
  NANDN U61522 ( .A(n51930), .B(n51929), .Z(n51925) );
  XOR U61523 ( .A(n51929), .B(n51931), .Z(N60764) );
  XNOR U61524 ( .A(n51927), .B(n51930), .Z(n51931) );
  NAND U61525 ( .A(n51932), .B(n51933), .Z(n51930) );
  NAND U61526 ( .A(n51934), .B(n51935), .Z(n51933) );
  NANDN U61527 ( .A(n51936), .B(n51937), .Z(n51935) );
  NANDN U61528 ( .A(n51937), .B(n51936), .Z(n51932) );
  AND U61529 ( .A(n51938), .B(n51939), .Z(n51927) );
  NAND U61530 ( .A(n51940), .B(n51941), .Z(n51939) );
  NANDN U61531 ( .A(n51942), .B(n51943), .Z(n51941) );
  NANDN U61532 ( .A(n51943), .B(n51942), .Z(n51938) );
  IV U61533 ( .A(n51944), .Z(n51943) );
  AND U61534 ( .A(n51945), .B(n51946), .Z(n51929) );
  NAND U61535 ( .A(n51947), .B(n51948), .Z(n51946) );
  NANDN U61536 ( .A(n51949), .B(n51950), .Z(n51948) );
  NANDN U61537 ( .A(n51950), .B(n51949), .Z(n51945) );
  XOR U61538 ( .A(n51942), .B(n51951), .Z(N60763) );
  XNOR U61539 ( .A(n51940), .B(n51944), .Z(n51951) );
  XOR U61540 ( .A(n51937), .B(n51952), .Z(n51944) );
  XNOR U61541 ( .A(n51934), .B(n51936), .Z(n51952) );
  AND U61542 ( .A(n51953), .B(n51954), .Z(n51936) );
  NANDN U61543 ( .A(n51955), .B(n51956), .Z(n51954) );
  OR U61544 ( .A(n51957), .B(n51958), .Z(n51956) );
  IV U61545 ( .A(n51959), .Z(n51958) );
  NANDN U61546 ( .A(n51959), .B(n51957), .Z(n51953) );
  AND U61547 ( .A(n51960), .B(n51961), .Z(n51934) );
  NAND U61548 ( .A(n51962), .B(n51963), .Z(n51961) );
  NANDN U61549 ( .A(n51964), .B(n51965), .Z(n51963) );
  NANDN U61550 ( .A(n51965), .B(n51964), .Z(n51960) );
  IV U61551 ( .A(n51966), .Z(n51965) );
  NAND U61552 ( .A(n51967), .B(n51968), .Z(n51937) );
  NANDN U61553 ( .A(n51969), .B(n51970), .Z(n51968) );
  NANDN U61554 ( .A(n51971), .B(n51972), .Z(n51970) );
  NANDN U61555 ( .A(n51972), .B(n51971), .Z(n51967) );
  IV U61556 ( .A(n51973), .Z(n51971) );
  AND U61557 ( .A(n51974), .B(n51975), .Z(n51940) );
  NAND U61558 ( .A(n51976), .B(n51977), .Z(n51975) );
  NANDN U61559 ( .A(n51978), .B(n51979), .Z(n51977) );
  NANDN U61560 ( .A(n51979), .B(n51978), .Z(n51974) );
  XOR U61561 ( .A(n51950), .B(n51980), .Z(n51942) );
  XNOR U61562 ( .A(n51947), .B(n51949), .Z(n51980) );
  AND U61563 ( .A(n51981), .B(n51982), .Z(n51949) );
  NANDN U61564 ( .A(n51983), .B(n51984), .Z(n51982) );
  OR U61565 ( .A(n51985), .B(n51986), .Z(n51984) );
  IV U61566 ( .A(n51987), .Z(n51986) );
  NANDN U61567 ( .A(n51987), .B(n51985), .Z(n51981) );
  AND U61568 ( .A(n51988), .B(n51989), .Z(n51947) );
  NAND U61569 ( .A(n51990), .B(n51991), .Z(n51989) );
  NANDN U61570 ( .A(n51992), .B(n51993), .Z(n51991) );
  NANDN U61571 ( .A(n51993), .B(n51992), .Z(n51988) );
  IV U61572 ( .A(n51994), .Z(n51993) );
  NAND U61573 ( .A(n51995), .B(n51996), .Z(n51950) );
  NANDN U61574 ( .A(n51997), .B(n51998), .Z(n51996) );
  NANDN U61575 ( .A(n51999), .B(n52000), .Z(n51998) );
  NANDN U61576 ( .A(n52000), .B(n51999), .Z(n51995) );
  IV U61577 ( .A(n52001), .Z(n51999) );
  XOR U61578 ( .A(n51976), .B(n52002), .Z(N60762) );
  XNOR U61579 ( .A(n51979), .B(n51978), .Z(n52002) );
  XNOR U61580 ( .A(n51990), .B(n52003), .Z(n51978) );
  XNOR U61581 ( .A(n51994), .B(n51992), .Z(n52003) );
  XOR U61582 ( .A(n52000), .B(n52004), .Z(n51992) );
  XNOR U61583 ( .A(n51997), .B(n52001), .Z(n52004) );
  AND U61584 ( .A(n52005), .B(n52006), .Z(n52001) );
  NAND U61585 ( .A(n52007), .B(n52008), .Z(n52006) );
  NAND U61586 ( .A(n52009), .B(n52010), .Z(n52005) );
  AND U61587 ( .A(n52011), .B(n52012), .Z(n51997) );
  NAND U61588 ( .A(n52013), .B(n52014), .Z(n52012) );
  NAND U61589 ( .A(n52015), .B(n52016), .Z(n52011) );
  NANDN U61590 ( .A(n52017), .B(n52018), .Z(n52000) );
  ANDN U61591 ( .B(n52019), .A(n52020), .Z(n51994) );
  XNOR U61592 ( .A(n51985), .B(n52021), .Z(n51990) );
  XNOR U61593 ( .A(n51983), .B(n51987), .Z(n52021) );
  AND U61594 ( .A(n52022), .B(n52023), .Z(n51987) );
  NAND U61595 ( .A(n52024), .B(n52025), .Z(n52023) );
  NAND U61596 ( .A(n52026), .B(n52027), .Z(n52022) );
  AND U61597 ( .A(n52028), .B(n52029), .Z(n51983) );
  NAND U61598 ( .A(n52030), .B(n52031), .Z(n52029) );
  NAND U61599 ( .A(n52032), .B(n52033), .Z(n52028) );
  AND U61600 ( .A(n52034), .B(n52035), .Z(n51985) );
  NAND U61601 ( .A(n52036), .B(n52037), .Z(n51979) );
  XNOR U61602 ( .A(n51962), .B(n52038), .Z(n51976) );
  XNOR U61603 ( .A(n51966), .B(n51964), .Z(n52038) );
  XOR U61604 ( .A(n51972), .B(n52039), .Z(n51964) );
  XNOR U61605 ( .A(n51969), .B(n51973), .Z(n52039) );
  AND U61606 ( .A(n52040), .B(n52041), .Z(n51973) );
  NAND U61607 ( .A(n52042), .B(n52043), .Z(n52041) );
  NAND U61608 ( .A(n52044), .B(n52045), .Z(n52040) );
  AND U61609 ( .A(n52046), .B(n52047), .Z(n51969) );
  NAND U61610 ( .A(n52048), .B(n52049), .Z(n52047) );
  NAND U61611 ( .A(n52050), .B(n52051), .Z(n52046) );
  NANDN U61612 ( .A(n52052), .B(n52053), .Z(n51972) );
  ANDN U61613 ( .B(n52054), .A(n52055), .Z(n51966) );
  XNOR U61614 ( .A(n51957), .B(n52056), .Z(n51962) );
  XNOR U61615 ( .A(n51955), .B(n51959), .Z(n52056) );
  AND U61616 ( .A(n52057), .B(n52058), .Z(n51959) );
  NAND U61617 ( .A(n52059), .B(n52060), .Z(n52058) );
  NAND U61618 ( .A(n52061), .B(n52062), .Z(n52057) );
  AND U61619 ( .A(n52063), .B(n52064), .Z(n51955) );
  NAND U61620 ( .A(n52065), .B(n52066), .Z(n52064) );
  NAND U61621 ( .A(n52067), .B(n52068), .Z(n52063) );
  AND U61622 ( .A(n52069), .B(n52070), .Z(n51957) );
  XOR U61623 ( .A(n52037), .B(n52036), .Z(N60761) );
  XNOR U61624 ( .A(n52054), .B(n52055), .Z(n52036) );
  XNOR U61625 ( .A(n52069), .B(n52070), .Z(n52055) );
  XOR U61626 ( .A(n52066), .B(n52065), .Z(n52070) );
  XOR U61627 ( .A(y[324]), .B(x[324]), .Z(n52065) );
  XOR U61628 ( .A(n52068), .B(n52067), .Z(n52066) );
  XOR U61629 ( .A(y[326]), .B(x[326]), .Z(n52067) );
  XOR U61630 ( .A(y[325]), .B(x[325]), .Z(n52068) );
  XOR U61631 ( .A(n52060), .B(n52059), .Z(n52069) );
  XOR U61632 ( .A(n52062), .B(n52061), .Z(n52059) );
  XOR U61633 ( .A(y[323]), .B(x[323]), .Z(n52061) );
  XOR U61634 ( .A(y[322]), .B(x[322]), .Z(n52062) );
  XOR U61635 ( .A(y[321]), .B(x[321]), .Z(n52060) );
  XNOR U61636 ( .A(n52053), .B(n52052), .Z(n52054) );
  XNOR U61637 ( .A(n52049), .B(n52048), .Z(n52052) );
  XOR U61638 ( .A(n52051), .B(n52050), .Z(n52048) );
  XOR U61639 ( .A(y[320]), .B(x[320]), .Z(n52050) );
  XOR U61640 ( .A(y[319]), .B(x[319]), .Z(n52051) );
  XOR U61641 ( .A(y[318]), .B(x[318]), .Z(n52049) );
  XOR U61642 ( .A(n52043), .B(n52042), .Z(n52053) );
  XOR U61643 ( .A(n52045), .B(n52044), .Z(n52042) );
  XOR U61644 ( .A(y[317]), .B(x[317]), .Z(n52044) );
  XOR U61645 ( .A(y[316]), .B(x[316]), .Z(n52045) );
  XOR U61646 ( .A(y[315]), .B(x[315]), .Z(n52043) );
  XNOR U61647 ( .A(n52019), .B(n52020), .Z(n52037) );
  XNOR U61648 ( .A(n52034), .B(n52035), .Z(n52020) );
  XOR U61649 ( .A(n52031), .B(n52030), .Z(n52035) );
  XOR U61650 ( .A(y[312]), .B(x[312]), .Z(n52030) );
  XOR U61651 ( .A(n52033), .B(n52032), .Z(n52031) );
  XOR U61652 ( .A(y[314]), .B(x[314]), .Z(n52032) );
  XOR U61653 ( .A(y[313]), .B(x[313]), .Z(n52033) );
  XOR U61654 ( .A(n52025), .B(n52024), .Z(n52034) );
  XOR U61655 ( .A(n52027), .B(n52026), .Z(n52024) );
  XOR U61656 ( .A(y[311]), .B(x[311]), .Z(n52026) );
  XOR U61657 ( .A(y[310]), .B(x[310]), .Z(n52027) );
  XOR U61658 ( .A(y[309]), .B(x[309]), .Z(n52025) );
  XNOR U61659 ( .A(n52018), .B(n52017), .Z(n52019) );
  XNOR U61660 ( .A(n52014), .B(n52013), .Z(n52017) );
  XOR U61661 ( .A(n52016), .B(n52015), .Z(n52013) );
  XOR U61662 ( .A(y[308]), .B(x[308]), .Z(n52015) );
  XOR U61663 ( .A(y[307]), .B(x[307]), .Z(n52016) );
  XOR U61664 ( .A(y[306]), .B(x[306]), .Z(n52014) );
  XOR U61665 ( .A(n52008), .B(n52007), .Z(n52018) );
  XOR U61666 ( .A(n52010), .B(n52009), .Z(n52007) );
  XOR U61667 ( .A(y[305]), .B(x[305]), .Z(n52009) );
  XOR U61668 ( .A(y[304]), .B(x[304]), .Z(n52010) );
  XOR U61669 ( .A(y[303]), .B(x[303]), .Z(n52008) );
  NAND U61670 ( .A(n52071), .B(n52072), .Z(N60752) );
  NAND U61671 ( .A(n52073), .B(n52074), .Z(n52072) );
  NANDN U61672 ( .A(n52075), .B(n52076), .Z(n52074) );
  NANDN U61673 ( .A(n52076), .B(n52075), .Z(n52071) );
  XOR U61674 ( .A(n52075), .B(n52077), .Z(N60751) );
  XNOR U61675 ( .A(n52073), .B(n52076), .Z(n52077) );
  NAND U61676 ( .A(n52078), .B(n52079), .Z(n52076) );
  NAND U61677 ( .A(n52080), .B(n52081), .Z(n52079) );
  NANDN U61678 ( .A(n52082), .B(n52083), .Z(n52081) );
  NANDN U61679 ( .A(n52083), .B(n52082), .Z(n52078) );
  AND U61680 ( .A(n52084), .B(n52085), .Z(n52073) );
  NAND U61681 ( .A(n52086), .B(n52087), .Z(n52085) );
  NANDN U61682 ( .A(n52088), .B(n52089), .Z(n52087) );
  NANDN U61683 ( .A(n52089), .B(n52088), .Z(n52084) );
  IV U61684 ( .A(n52090), .Z(n52089) );
  AND U61685 ( .A(n52091), .B(n52092), .Z(n52075) );
  NAND U61686 ( .A(n52093), .B(n52094), .Z(n52092) );
  NANDN U61687 ( .A(n52095), .B(n52096), .Z(n52094) );
  NANDN U61688 ( .A(n52096), .B(n52095), .Z(n52091) );
  XOR U61689 ( .A(n52088), .B(n52097), .Z(N60750) );
  XNOR U61690 ( .A(n52086), .B(n52090), .Z(n52097) );
  XOR U61691 ( .A(n52083), .B(n52098), .Z(n52090) );
  XNOR U61692 ( .A(n52080), .B(n52082), .Z(n52098) );
  AND U61693 ( .A(n52099), .B(n52100), .Z(n52082) );
  NANDN U61694 ( .A(n52101), .B(n52102), .Z(n52100) );
  OR U61695 ( .A(n52103), .B(n52104), .Z(n52102) );
  IV U61696 ( .A(n52105), .Z(n52104) );
  NANDN U61697 ( .A(n52105), .B(n52103), .Z(n52099) );
  AND U61698 ( .A(n52106), .B(n52107), .Z(n52080) );
  NAND U61699 ( .A(n52108), .B(n52109), .Z(n52107) );
  NANDN U61700 ( .A(n52110), .B(n52111), .Z(n52109) );
  NANDN U61701 ( .A(n52111), .B(n52110), .Z(n52106) );
  IV U61702 ( .A(n52112), .Z(n52111) );
  NAND U61703 ( .A(n52113), .B(n52114), .Z(n52083) );
  NANDN U61704 ( .A(n52115), .B(n52116), .Z(n52114) );
  NANDN U61705 ( .A(n52117), .B(n52118), .Z(n52116) );
  NANDN U61706 ( .A(n52118), .B(n52117), .Z(n52113) );
  IV U61707 ( .A(n52119), .Z(n52117) );
  AND U61708 ( .A(n52120), .B(n52121), .Z(n52086) );
  NAND U61709 ( .A(n52122), .B(n52123), .Z(n52121) );
  NANDN U61710 ( .A(n52124), .B(n52125), .Z(n52123) );
  NANDN U61711 ( .A(n52125), .B(n52124), .Z(n52120) );
  XOR U61712 ( .A(n52096), .B(n52126), .Z(n52088) );
  XNOR U61713 ( .A(n52093), .B(n52095), .Z(n52126) );
  AND U61714 ( .A(n52127), .B(n52128), .Z(n52095) );
  NANDN U61715 ( .A(n52129), .B(n52130), .Z(n52128) );
  OR U61716 ( .A(n52131), .B(n52132), .Z(n52130) );
  IV U61717 ( .A(n52133), .Z(n52132) );
  NANDN U61718 ( .A(n52133), .B(n52131), .Z(n52127) );
  AND U61719 ( .A(n52134), .B(n52135), .Z(n52093) );
  NAND U61720 ( .A(n52136), .B(n52137), .Z(n52135) );
  NANDN U61721 ( .A(n52138), .B(n52139), .Z(n52137) );
  NANDN U61722 ( .A(n52139), .B(n52138), .Z(n52134) );
  IV U61723 ( .A(n52140), .Z(n52139) );
  NAND U61724 ( .A(n52141), .B(n52142), .Z(n52096) );
  NANDN U61725 ( .A(n52143), .B(n52144), .Z(n52142) );
  NANDN U61726 ( .A(n52145), .B(n52146), .Z(n52144) );
  NANDN U61727 ( .A(n52146), .B(n52145), .Z(n52141) );
  IV U61728 ( .A(n52147), .Z(n52145) );
  XOR U61729 ( .A(n52122), .B(n52148), .Z(N60749) );
  XNOR U61730 ( .A(n52125), .B(n52124), .Z(n52148) );
  XNOR U61731 ( .A(n52136), .B(n52149), .Z(n52124) );
  XNOR U61732 ( .A(n52140), .B(n52138), .Z(n52149) );
  XOR U61733 ( .A(n52146), .B(n52150), .Z(n52138) );
  XNOR U61734 ( .A(n52143), .B(n52147), .Z(n52150) );
  AND U61735 ( .A(n52151), .B(n52152), .Z(n52147) );
  NAND U61736 ( .A(n52153), .B(n52154), .Z(n52152) );
  NAND U61737 ( .A(n52155), .B(n52156), .Z(n52151) );
  AND U61738 ( .A(n52157), .B(n52158), .Z(n52143) );
  NAND U61739 ( .A(n52159), .B(n52160), .Z(n52158) );
  NAND U61740 ( .A(n52161), .B(n52162), .Z(n52157) );
  NANDN U61741 ( .A(n52163), .B(n52164), .Z(n52146) );
  ANDN U61742 ( .B(n52165), .A(n52166), .Z(n52140) );
  XNOR U61743 ( .A(n52131), .B(n52167), .Z(n52136) );
  XNOR U61744 ( .A(n52129), .B(n52133), .Z(n52167) );
  AND U61745 ( .A(n52168), .B(n52169), .Z(n52133) );
  NAND U61746 ( .A(n52170), .B(n52171), .Z(n52169) );
  NAND U61747 ( .A(n52172), .B(n52173), .Z(n52168) );
  AND U61748 ( .A(n52174), .B(n52175), .Z(n52129) );
  NAND U61749 ( .A(n52176), .B(n52177), .Z(n52175) );
  NAND U61750 ( .A(n52178), .B(n52179), .Z(n52174) );
  AND U61751 ( .A(n52180), .B(n52181), .Z(n52131) );
  NAND U61752 ( .A(n52182), .B(n52183), .Z(n52125) );
  XNOR U61753 ( .A(n52108), .B(n52184), .Z(n52122) );
  XNOR U61754 ( .A(n52112), .B(n52110), .Z(n52184) );
  XOR U61755 ( .A(n52118), .B(n52185), .Z(n52110) );
  XNOR U61756 ( .A(n52115), .B(n52119), .Z(n52185) );
  AND U61757 ( .A(n52186), .B(n52187), .Z(n52119) );
  NAND U61758 ( .A(n52188), .B(n52189), .Z(n52187) );
  NAND U61759 ( .A(n52190), .B(n52191), .Z(n52186) );
  AND U61760 ( .A(n52192), .B(n52193), .Z(n52115) );
  NAND U61761 ( .A(n52194), .B(n52195), .Z(n52193) );
  NAND U61762 ( .A(n52196), .B(n52197), .Z(n52192) );
  NANDN U61763 ( .A(n52198), .B(n52199), .Z(n52118) );
  ANDN U61764 ( .B(n52200), .A(n52201), .Z(n52112) );
  XNOR U61765 ( .A(n52103), .B(n52202), .Z(n52108) );
  XNOR U61766 ( .A(n52101), .B(n52105), .Z(n52202) );
  AND U61767 ( .A(n52203), .B(n52204), .Z(n52105) );
  NAND U61768 ( .A(n52205), .B(n52206), .Z(n52204) );
  NAND U61769 ( .A(n52207), .B(n52208), .Z(n52203) );
  AND U61770 ( .A(n52209), .B(n52210), .Z(n52101) );
  NAND U61771 ( .A(n52211), .B(n52212), .Z(n52210) );
  NAND U61772 ( .A(n52213), .B(n52214), .Z(n52209) );
  AND U61773 ( .A(n52215), .B(n52216), .Z(n52103) );
  XOR U61774 ( .A(n52183), .B(n52182), .Z(N60748) );
  XNOR U61775 ( .A(n52200), .B(n52201), .Z(n52182) );
  XNOR U61776 ( .A(n52215), .B(n52216), .Z(n52201) );
  XOR U61777 ( .A(n52212), .B(n52211), .Z(n52216) );
  XOR U61778 ( .A(y[300]), .B(x[300]), .Z(n52211) );
  XOR U61779 ( .A(n52214), .B(n52213), .Z(n52212) );
  XOR U61780 ( .A(y[302]), .B(x[302]), .Z(n52213) );
  XOR U61781 ( .A(y[301]), .B(x[301]), .Z(n52214) );
  XOR U61782 ( .A(n52206), .B(n52205), .Z(n52215) );
  XOR U61783 ( .A(n52208), .B(n52207), .Z(n52205) );
  XOR U61784 ( .A(y[299]), .B(x[299]), .Z(n52207) );
  XOR U61785 ( .A(y[298]), .B(x[298]), .Z(n52208) );
  XOR U61786 ( .A(y[297]), .B(x[297]), .Z(n52206) );
  XNOR U61787 ( .A(n52199), .B(n52198), .Z(n52200) );
  XNOR U61788 ( .A(n52195), .B(n52194), .Z(n52198) );
  XOR U61789 ( .A(n52197), .B(n52196), .Z(n52194) );
  XOR U61790 ( .A(y[296]), .B(x[296]), .Z(n52196) );
  XOR U61791 ( .A(y[295]), .B(x[295]), .Z(n52197) );
  XOR U61792 ( .A(y[294]), .B(x[294]), .Z(n52195) );
  XOR U61793 ( .A(n52189), .B(n52188), .Z(n52199) );
  XOR U61794 ( .A(n52191), .B(n52190), .Z(n52188) );
  XOR U61795 ( .A(y[293]), .B(x[293]), .Z(n52190) );
  XOR U61796 ( .A(y[292]), .B(x[292]), .Z(n52191) );
  XOR U61797 ( .A(y[291]), .B(x[291]), .Z(n52189) );
  XNOR U61798 ( .A(n52165), .B(n52166), .Z(n52183) );
  XNOR U61799 ( .A(n52180), .B(n52181), .Z(n52166) );
  XOR U61800 ( .A(n52177), .B(n52176), .Z(n52181) );
  XOR U61801 ( .A(y[288]), .B(x[288]), .Z(n52176) );
  XOR U61802 ( .A(n52179), .B(n52178), .Z(n52177) );
  XOR U61803 ( .A(y[290]), .B(x[290]), .Z(n52178) );
  XOR U61804 ( .A(y[289]), .B(x[289]), .Z(n52179) );
  XOR U61805 ( .A(n52171), .B(n52170), .Z(n52180) );
  XOR U61806 ( .A(n52173), .B(n52172), .Z(n52170) );
  XOR U61807 ( .A(y[287]), .B(x[287]), .Z(n52172) );
  XOR U61808 ( .A(y[286]), .B(x[286]), .Z(n52173) );
  XOR U61809 ( .A(y[285]), .B(x[285]), .Z(n52171) );
  XNOR U61810 ( .A(n52164), .B(n52163), .Z(n52165) );
  XNOR U61811 ( .A(n52160), .B(n52159), .Z(n52163) );
  XOR U61812 ( .A(n52162), .B(n52161), .Z(n52159) );
  XOR U61813 ( .A(y[284]), .B(x[284]), .Z(n52161) );
  XOR U61814 ( .A(y[283]), .B(x[283]), .Z(n52162) );
  XOR U61815 ( .A(y[282]), .B(x[282]), .Z(n52160) );
  XOR U61816 ( .A(n52154), .B(n52153), .Z(n52164) );
  XOR U61817 ( .A(n52156), .B(n52155), .Z(n52153) );
  XOR U61818 ( .A(y[281]), .B(x[281]), .Z(n52155) );
  XOR U61819 ( .A(y[280]), .B(x[280]), .Z(n52156) );
  XOR U61820 ( .A(y[279]), .B(x[279]), .Z(n52154) );
  NAND U61821 ( .A(n52217), .B(n52218), .Z(N60739) );
  NAND U61822 ( .A(n52219), .B(n52220), .Z(n52218) );
  NANDN U61823 ( .A(n52221), .B(n52222), .Z(n52220) );
  NANDN U61824 ( .A(n52222), .B(n52221), .Z(n52217) );
  XOR U61825 ( .A(n52221), .B(n52223), .Z(N60738) );
  XNOR U61826 ( .A(n52219), .B(n52222), .Z(n52223) );
  NAND U61827 ( .A(n52224), .B(n52225), .Z(n52222) );
  NAND U61828 ( .A(n52226), .B(n52227), .Z(n52225) );
  NANDN U61829 ( .A(n52228), .B(n52229), .Z(n52227) );
  NANDN U61830 ( .A(n52229), .B(n52228), .Z(n52224) );
  AND U61831 ( .A(n52230), .B(n52231), .Z(n52219) );
  NAND U61832 ( .A(n52232), .B(n52233), .Z(n52231) );
  NANDN U61833 ( .A(n52234), .B(n52235), .Z(n52233) );
  NANDN U61834 ( .A(n52235), .B(n52234), .Z(n52230) );
  IV U61835 ( .A(n52236), .Z(n52235) );
  AND U61836 ( .A(n52237), .B(n52238), .Z(n52221) );
  NAND U61837 ( .A(n52239), .B(n52240), .Z(n52238) );
  NANDN U61838 ( .A(n52241), .B(n52242), .Z(n52240) );
  NANDN U61839 ( .A(n52242), .B(n52241), .Z(n52237) );
  XOR U61840 ( .A(n52234), .B(n52243), .Z(N60737) );
  XNOR U61841 ( .A(n52232), .B(n52236), .Z(n52243) );
  XOR U61842 ( .A(n52229), .B(n52244), .Z(n52236) );
  XNOR U61843 ( .A(n52226), .B(n52228), .Z(n52244) );
  AND U61844 ( .A(n52245), .B(n52246), .Z(n52228) );
  NANDN U61845 ( .A(n52247), .B(n52248), .Z(n52246) );
  OR U61846 ( .A(n52249), .B(n52250), .Z(n52248) );
  IV U61847 ( .A(n52251), .Z(n52250) );
  NANDN U61848 ( .A(n52251), .B(n52249), .Z(n52245) );
  AND U61849 ( .A(n52252), .B(n52253), .Z(n52226) );
  NAND U61850 ( .A(n52254), .B(n52255), .Z(n52253) );
  NANDN U61851 ( .A(n52256), .B(n52257), .Z(n52255) );
  NANDN U61852 ( .A(n52257), .B(n52256), .Z(n52252) );
  IV U61853 ( .A(n52258), .Z(n52257) );
  NAND U61854 ( .A(n52259), .B(n52260), .Z(n52229) );
  NANDN U61855 ( .A(n52261), .B(n52262), .Z(n52260) );
  NANDN U61856 ( .A(n52263), .B(n52264), .Z(n52262) );
  NANDN U61857 ( .A(n52264), .B(n52263), .Z(n52259) );
  IV U61858 ( .A(n52265), .Z(n52263) );
  AND U61859 ( .A(n52266), .B(n52267), .Z(n52232) );
  NAND U61860 ( .A(n52268), .B(n52269), .Z(n52267) );
  NANDN U61861 ( .A(n52270), .B(n52271), .Z(n52269) );
  NANDN U61862 ( .A(n52271), .B(n52270), .Z(n52266) );
  XOR U61863 ( .A(n52242), .B(n52272), .Z(n52234) );
  XNOR U61864 ( .A(n52239), .B(n52241), .Z(n52272) );
  AND U61865 ( .A(n52273), .B(n52274), .Z(n52241) );
  NANDN U61866 ( .A(n52275), .B(n52276), .Z(n52274) );
  OR U61867 ( .A(n52277), .B(n52278), .Z(n52276) );
  IV U61868 ( .A(n52279), .Z(n52278) );
  NANDN U61869 ( .A(n52279), .B(n52277), .Z(n52273) );
  AND U61870 ( .A(n52280), .B(n52281), .Z(n52239) );
  NAND U61871 ( .A(n52282), .B(n52283), .Z(n52281) );
  NANDN U61872 ( .A(n52284), .B(n52285), .Z(n52283) );
  NANDN U61873 ( .A(n52285), .B(n52284), .Z(n52280) );
  IV U61874 ( .A(n52286), .Z(n52285) );
  NAND U61875 ( .A(n52287), .B(n52288), .Z(n52242) );
  NANDN U61876 ( .A(n52289), .B(n52290), .Z(n52288) );
  NANDN U61877 ( .A(n52291), .B(n52292), .Z(n52290) );
  NANDN U61878 ( .A(n52292), .B(n52291), .Z(n52287) );
  IV U61879 ( .A(n52293), .Z(n52291) );
  XOR U61880 ( .A(n52268), .B(n52294), .Z(N60736) );
  XNOR U61881 ( .A(n52271), .B(n52270), .Z(n52294) );
  XNOR U61882 ( .A(n52282), .B(n52295), .Z(n52270) );
  XNOR U61883 ( .A(n52286), .B(n52284), .Z(n52295) );
  XOR U61884 ( .A(n52292), .B(n52296), .Z(n52284) );
  XNOR U61885 ( .A(n52289), .B(n52293), .Z(n52296) );
  AND U61886 ( .A(n52297), .B(n52298), .Z(n52293) );
  NAND U61887 ( .A(n52299), .B(n52300), .Z(n52298) );
  NAND U61888 ( .A(n52301), .B(n52302), .Z(n52297) );
  AND U61889 ( .A(n52303), .B(n52304), .Z(n52289) );
  NAND U61890 ( .A(n52305), .B(n52306), .Z(n52304) );
  NAND U61891 ( .A(n52307), .B(n52308), .Z(n52303) );
  NANDN U61892 ( .A(n52309), .B(n52310), .Z(n52292) );
  ANDN U61893 ( .B(n52311), .A(n52312), .Z(n52286) );
  XNOR U61894 ( .A(n52277), .B(n52313), .Z(n52282) );
  XNOR U61895 ( .A(n52275), .B(n52279), .Z(n52313) );
  AND U61896 ( .A(n52314), .B(n52315), .Z(n52279) );
  NAND U61897 ( .A(n52316), .B(n52317), .Z(n52315) );
  NAND U61898 ( .A(n52318), .B(n52319), .Z(n52314) );
  AND U61899 ( .A(n52320), .B(n52321), .Z(n52275) );
  NAND U61900 ( .A(n52322), .B(n52323), .Z(n52321) );
  NAND U61901 ( .A(n52324), .B(n52325), .Z(n52320) );
  AND U61902 ( .A(n52326), .B(n52327), .Z(n52277) );
  NAND U61903 ( .A(n52328), .B(n52329), .Z(n52271) );
  XNOR U61904 ( .A(n52254), .B(n52330), .Z(n52268) );
  XNOR U61905 ( .A(n52258), .B(n52256), .Z(n52330) );
  XOR U61906 ( .A(n52264), .B(n52331), .Z(n52256) );
  XNOR U61907 ( .A(n52261), .B(n52265), .Z(n52331) );
  AND U61908 ( .A(n52332), .B(n52333), .Z(n52265) );
  NAND U61909 ( .A(n52334), .B(n52335), .Z(n52333) );
  NAND U61910 ( .A(n52336), .B(n52337), .Z(n52332) );
  AND U61911 ( .A(n52338), .B(n52339), .Z(n52261) );
  NAND U61912 ( .A(n52340), .B(n52341), .Z(n52339) );
  NAND U61913 ( .A(n52342), .B(n52343), .Z(n52338) );
  NANDN U61914 ( .A(n52344), .B(n52345), .Z(n52264) );
  ANDN U61915 ( .B(n52346), .A(n52347), .Z(n52258) );
  XNOR U61916 ( .A(n52249), .B(n52348), .Z(n52254) );
  XNOR U61917 ( .A(n52247), .B(n52251), .Z(n52348) );
  AND U61918 ( .A(n52349), .B(n52350), .Z(n52251) );
  NAND U61919 ( .A(n52351), .B(n52352), .Z(n52350) );
  NAND U61920 ( .A(n52353), .B(n52354), .Z(n52349) );
  AND U61921 ( .A(n52355), .B(n52356), .Z(n52247) );
  NAND U61922 ( .A(n52357), .B(n52358), .Z(n52356) );
  NAND U61923 ( .A(n52359), .B(n52360), .Z(n52355) );
  AND U61924 ( .A(n52361), .B(n52362), .Z(n52249) );
  XOR U61925 ( .A(n52329), .B(n52328), .Z(N60735) );
  XNOR U61926 ( .A(n52346), .B(n52347), .Z(n52328) );
  XNOR U61927 ( .A(n52361), .B(n52362), .Z(n52347) );
  XOR U61928 ( .A(n52358), .B(n52357), .Z(n52362) );
  XOR U61929 ( .A(y[276]), .B(x[276]), .Z(n52357) );
  XOR U61930 ( .A(n52360), .B(n52359), .Z(n52358) );
  XOR U61931 ( .A(y[278]), .B(x[278]), .Z(n52359) );
  XOR U61932 ( .A(y[277]), .B(x[277]), .Z(n52360) );
  XOR U61933 ( .A(n52352), .B(n52351), .Z(n52361) );
  XOR U61934 ( .A(n52354), .B(n52353), .Z(n52351) );
  XOR U61935 ( .A(y[275]), .B(x[275]), .Z(n52353) );
  XOR U61936 ( .A(y[274]), .B(x[274]), .Z(n52354) );
  XOR U61937 ( .A(y[273]), .B(x[273]), .Z(n52352) );
  XNOR U61938 ( .A(n52345), .B(n52344), .Z(n52346) );
  XNOR U61939 ( .A(n52341), .B(n52340), .Z(n52344) );
  XOR U61940 ( .A(n52343), .B(n52342), .Z(n52340) );
  XOR U61941 ( .A(y[272]), .B(x[272]), .Z(n52342) );
  XOR U61942 ( .A(y[271]), .B(x[271]), .Z(n52343) );
  XOR U61943 ( .A(y[270]), .B(x[270]), .Z(n52341) );
  XOR U61944 ( .A(n52335), .B(n52334), .Z(n52345) );
  XOR U61945 ( .A(n52337), .B(n52336), .Z(n52334) );
  XOR U61946 ( .A(y[269]), .B(x[269]), .Z(n52336) );
  XOR U61947 ( .A(y[268]), .B(x[268]), .Z(n52337) );
  XOR U61948 ( .A(y[267]), .B(x[267]), .Z(n52335) );
  XNOR U61949 ( .A(n52311), .B(n52312), .Z(n52329) );
  XNOR U61950 ( .A(n52326), .B(n52327), .Z(n52312) );
  XOR U61951 ( .A(n52323), .B(n52322), .Z(n52327) );
  XOR U61952 ( .A(y[264]), .B(x[264]), .Z(n52322) );
  XOR U61953 ( .A(n52325), .B(n52324), .Z(n52323) );
  XOR U61954 ( .A(y[266]), .B(x[266]), .Z(n52324) );
  XOR U61955 ( .A(y[265]), .B(x[265]), .Z(n52325) );
  XOR U61956 ( .A(n52317), .B(n52316), .Z(n52326) );
  XOR U61957 ( .A(n52319), .B(n52318), .Z(n52316) );
  XOR U61958 ( .A(y[263]), .B(x[263]), .Z(n52318) );
  XOR U61959 ( .A(y[262]), .B(x[262]), .Z(n52319) );
  XOR U61960 ( .A(y[261]), .B(x[261]), .Z(n52317) );
  XNOR U61961 ( .A(n52310), .B(n52309), .Z(n52311) );
  XNOR U61962 ( .A(n52306), .B(n52305), .Z(n52309) );
  XOR U61963 ( .A(n52308), .B(n52307), .Z(n52305) );
  XOR U61964 ( .A(y[260]), .B(x[260]), .Z(n52307) );
  XOR U61965 ( .A(y[259]), .B(x[259]), .Z(n52308) );
  XOR U61966 ( .A(y[258]), .B(x[258]), .Z(n52306) );
  XOR U61967 ( .A(n52300), .B(n52299), .Z(n52310) );
  XOR U61968 ( .A(n52302), .B(n52301), .Z(n52299) );
  XOR U61969 ( .A(y[257]), .B(x[257]), .Z(n52301) );
  XOR U61970 ( .A(y[256]), .B(x[256]), .Z(n52302) );
  XOR U61971 ( .A(y[255]), .B(x[255]), .Z(n52300) );
  NAND U61972 ( .A(n52363), .B(n52364), .Z(N60726) );
  NAND U61973 ( .A(n52365), .B(n52366), .Z(n52364) );
  NANDN U61974 ( .A(n52367), .B(n52368), .Z(n52366) );
  NANDN U61975 ( .A(n52368), .B(n52367), .Z(n52363) );
  XOR U61976 ( .A(n52367), .B(n52369), .Z(N60725) );
  XNOR U61977 ( .A(n52365), .B(n52368), .Z(n52369) );
  NAND U61978 ( .A(n52370), .B(n52371), .Z(n52368) );
  NAND U61979 ( .A(n52372), .B(n52373), .Z(n52371) );
  NANDN U61980 ( .A(n52374), .B(n52375), .Z(n52373) );
  NANDN U61981 ( .A(n52375), .B(n52374), .Z(n52370) );
  AND U61982 ( .A(n52376), .B(n52377), .Z(n52365) );
  NAND U61983 ( .A(n52378), .B(n52379), .Z(n52377) );
  NANDN U61984 ( .A(n52380), .B(n52381), .Z(n52379) );
  NANDN U61985 ( .A(n52381), .B(n52380), .Z(n52376) );
  IV U61986 ( .A(n52382), .Z(n52381) );
  AND U61987 ( .A(n52383), .B(n52384), .Z(n52367) );
  NAND U61988 ( .A(n52385), .B(n52386), .Z(n52384) );
  NANDN U61989 ( .A(n52387), .B(n52388), .Z(n52386) );
  NANDN U61990 ( .A(n52388), .B(n52387), .Z(n52383) );
  XOR U61991 ( .A(n52380), .B(n52389), .Z(N60724) );
  XNOR U61992 ( .A(n52378), .B(n52382), .Z(n52389) );
  XOR U61993 ( .A(n52375), .B(n52390), .Z(n52382) );
  XNOR U61994 ( .A(n52372), .B(n52374), .Z(n52390) );
  AND U61995 ( .A(n52391), .B(n52392), .Z(n52374) );
  NANDN U61996 ( .A(n52393), .B(n52394), .Z(n52392) );
  OR U61997 ( .A(n52395), .B(n52396), .Z(n52394) );
  IV U61998 ( .A(n52397), .Z(n52396) );
  NANDN U61999 ( .A(n52397), .B(n52395), .Z(n52391) );
  AND U62000 ( .A(n52398), .B(n52399), .Z(n52372) );
  NAND U62001 ( .A(n52400), .B(n52401), .Z(n52399) );
  NANDN U62002 ( .A(n52402), .B(n52403), .Z(n52401) );
  NANDN U62003 ( .A(n52403), .B(n52402), .Z(n52398) );
  IV U62004 ( .A(n52404), .Z(n52403) );
  NAND U62005 ( .A(n52405), .B(n52406), .Z(n52375) );
  NANDN U62006 ( .A(n52407), .B(n52408), .Z(n52406) );
  NANDN U62007 ( .A(n52409), .B(n52410), .Z(n52408) );
  NANDN U62008 ( .A(n52410), .B(n52409), .Z(n52405) );
  IV U62009 ( .A(n52411), .Z(n52409) );
  AND U62010 ( .A(n52412), .B(n52413), .Z(n52378) );
  NAND U62011 ( .A(n52414), .B(n52415), .Z(n52413) );
  NANDN U62012 ( .A(n52416), .B(n52417), .Z(n52415) );
  NANDN U62013 ( .A(n52417), .B(n52416), .Z(n52412) );
  XOR U62014 ( .A(n52388), .B(n52418), .Z(n52380) );
  XNOR U62015 ( .A(n52385), .B(n52387), .Z(n52418) );
  AND U62016 ( .A(n52419), .B(n52420), .Z(n52387) );
  NANDN U62017 ( .A(n52421), .B(n52422), .Z(n52420) );
  OR U62018 ( .A(n52423), .B(n52424), .Z(n52422) );
  IV U62019 ( .A(n52425), .Z(n52424) );
  NANDN U62020 ( .A(n52425), .B(n52423), .Z(n52419) );
  AND U62021 ( .A(n52426), .B(n52427), .Z(n52385) );
  NAND U62022 ( .A(n52428), .B(n52429), .Z(n52427) );
  NANDN U62023 ( .A(n52430), .B(n52431), .Z(n52429) );
  NANDN U62024 ( .A(n52431), .B(n52430), .Z(n52426) );
  IV U62025 ( .A(n52432), .Z(n52431) );
  NAND U62026 ( .A(n52433), .B(n52434), .Z(n52388) );
  NANDN U62027 ( .A(n52435), .B(n52436), .Z(n52434) );
  NANDN U62028 ( .A(n52437), .B(n52438), .Z(n52436) );
  NANDN U62029 ( .A(n52438), .B(n52437), .Z(n52433) );
  IV U62030 ( .A(n52439), .Z(n52437) );
  XOR U62031 ( .A(n52414), .B(n52440), .Z(N60723) );
  XNOR U62032 ( .A(n52417), .B(n52416), .Z(n52440) );
  XNOR U62033 ( .A(n52428), .B(n52441), .Z(n52416) );
  XNOR U62034 ( .A(n52432), .B(n52430), .Z(n52441) );
  XOR U62035 ( .A(n52438), .B(n52442), .Z(n52430) );
  XNOR U62036 ( .A(n52435), .B(n52439), .Z(n52442) );
  AND U62037 ( .A(n52443), .B(n52444), .Z(n52439) );
  NAND U62038 ( .A(n52445), .B(n52446), .Z(n52444) );
  NAND U62039 ( .A(n52447), .B(n52448), .Z(n52443) );
  AND U62040 ( .A(n52449), .B(n52450), .Z(n52435) );
  NAND U62041 ( .A(n52451), .B(n52452), .Z(n52450) );
  NAND U62042 ( .A(n52453), .B(n52454), .Z(n52449) );
  NANDN U62043 ( .A(n52455), .B(n52456), .Z(n52438) );
  ANDN U62044 ( .B(n52457), .A(n52458), .Z(n52432) );
  XNOR U62045 ( .A(n52423), .B(n52459), .Z(n52428) );
  XNOR U62046 ( .A(n52421), .B(n52425), .Z(n52459) );
  AND U62047 ( .A(n52460), .B(n52461), .Z(n52425) );
  NAND U62048 ( .A(n52462), .B(n52463), .Z(n52461) );
  NAND U62049 ( .A(n52464), .B(n52465), .Z(n52460) );
  AND U62050 ( .A(n52466), .B(n52467), .Z(n52421) );
  NAND U62051 ( .A(n52468), .B(n52469), .Z(n52467) );
  NAND U62052 ( .A(n52470), .B(n52471), .Z(n52466) );
  AND U62053 ( .A(n52472), .B(n52473), .Z(n52423) );
  NAND U62054 ( .A(n52474), .B(n52475), .Z(n52417) );
  XNOR U62055 ( .A(n52400), .B(n52476), .Z(n52414) );
  XNOR U62056 ( .A(n52404), .B(n52402), .Z(n52476) );
  XOR U62057 ( .A(n52410), .B(n52477), .Z(n52402) );
  XNOR U62058 ( .A(n52407), .B(n52411), .Z(n52477) );
  AND U62059 ( .A(n52478), .B(n52479), .Z(n52411) );
  NAND U62060 ( .A(n52480), .B(n52481), .Z(n52479) );
  NAND U62061 ( .A(n52482), .B(n52483), .Z(n52478) );
  AND U62062 ( .A(n52484), .B(n52485), .Z(n52407) );
  NAND U62063 ( .A(n52486), .B(n52487), .Z(n52485) );
  NAND U62064 ( .A(n52488), .B(n52489), .Z(n52484) );
  NANDN U62065 ( .A(n52490), .B(n52491), .Z(n52410) );
  ANDN U62066 ( .B(n52492), .A(n52493), .Z(n52404) );
  XNOR U62067 ( .A(n52395), .B(n52494), .Z(n52400) );
  XNOR U62068 ( .A(n52393), .B(n52397), .Z(n52494) );
  AND U62069 ( .A(n52495), .B(n52496), .Z(n52397) );
  NAND U62070 ( .A(n52497), .B(n52498), .Z(n52496) );
  NAND U62071 ( .A(n52499), .B(n52500), .Z(n52495) );
  AND U62072 ( .A(n52501), .B(n52502), .Z(n52393) );
  NAND U62073 ( .A(n52503), .B(n52504), .Z(n52502) );
  NAND U62074 ( .A(n52505), .B(n52506), .Z(n52501) );
  AND U62075 ( .A(n52507), .B(n52508), .Z(n52395) );
  XOR U62076 ( .A(n52475), .B(n52474), .Z(N60722) );
  XNOR U62077 ( .A(n52492), .B(n52493), .Z(n52474) );
  XNOR U62078 ( .A(n52507), .B(n52508), .Z(n52493) );
  XOR U62079 ( .A(n52504), .B(n52503), .Z(n52508) );
  XOR U62080 ( .A(y[252]), .B(x[252]), .Z(n52503) );
  XOR U62081 ( .A(n52506), .B(n52505), .Z(n52504) );
  XOR U62082 ( .A(y[254]), .B(x[254]), .Z(n52505) );
  XOR U62083 ( .A(y[253]), .B(x[253]), .Z(n52506) );
  XOR U62084 ( .A(n52498), .B(n52497), .Z(n52507) );
  XOR U62085 ( .A(n52500), .B(n52499), .Z(n52497) );
  XOR U62086 ( .A(y[251]), .B(x[251]), .Z(n52499) );
  XOR U62087 ( .A(y[250]), .B(x[250]), .Z(n52500) );
  XOR U62088 ( .A(y[249]), .B(x[249]), .Z(n52498) );
  XNOR U62089 ( .A(n52491), .B(n52490), .Z(n52492) );
  XNOR U62090 ( .A(n52487), .B(n52486), .Z(n52490) );
  XOR U62091 ( .A(n52489), .B(n52488), .Z(n52486) );
  XOR U62092 ( .A(y[248]), .B(x[248]), .Z(n52488) );
  XOR U62093 ( .A(y[247]), .B(x[247]), .Z(n52489) );
  XOR U62094 ( .A(y[246]), .B(x[246]), .Z(n52487) );
  XOR U62095 ( .A(n52481), .B(n52480), .Z(n52491) );
  XOR U62096 ( .A(n52483), .B(n52482), .Z(n52480) );
  XOR U62097 ( .A(y[245]), .B(x[245]), .Z(n52482) );
  XOR U62098 ( .A(y[244]), .B(x[244]), .Z(n52483) );
  XOR U62099 ( .A(y[243]), .B(x[243]), .Z(n52481) );
  XNOR U62100 ( .A(n52457), .B(n52458), .Z(n52475) );
  XNOR U62101 ( .A(n52472), .B(n52473), .Z(n52458) );
  XOR U62102 ( .A(n52469), .B(n52468), .Z(n52473) );
  XOR U62103 ( .A(y[240]), .B(x[240]), .Z(n52468) );
  XOR U62104 ( .A(n52471), .B(n52470), .Z(n52469) );
  XOR U62105 ( .A(y[242]), .B(x[242]), .Z(n52470) );
  XOR U62106 ( .A(y[241]), .B(x[241]), .Z(n52471) );
  XOR U62107 ( .A(n52463), .B(n52462), .Z(n52472) );
  XOR U62108 ( .A(n52465), .B(n52464), .Z(n52462) );
  XOR U62109 ( .A(y[239]), .B(x[239]), .Z(n52464) );
  XOR U62110 ( .A(y[238]), .B(x[238]), .Z(n52465) );
  XOR U62111 ( .A(y[237]), .B(x[237]), .Z(n52463) );
  XNOR U62112 ( .A(n52456), .B(n52455), .Z(n52457) );
  XNOR U62113 ( .A(n52452), .B(n52451), .Z(n52455) );
  XOR U62114 ( .A(n52454), .B(n52453), .Z(n52451) );
  XOR U62115 ( .A(y[236]), .B(x[236]), .Z(n52453) );
  XOR U62116 ( .A(y[235]), .B(x[235]), .Z(n52454) );
  XOR U62117 ( .A(y[234]), .B(x[234]), .Z(n52452) );
  XOR U62118 ( .A(n52446), .B(n52445), .Z(n52456) );
  XOR U62119 ( .A(n52448), .B(n52447), .Z(n52445) );
  XOR U62120 ( .A(y[233]), .B(x[233]), .Z(n52447) );
  XOR U62121 ( .A(y[232]), .B(x[232]), .Z(n52448) );
  XOR U62122 ( .A(y[231]), .B(x[231]), .Z(n52446) );
  NAND U62123 ( .A(n52509), .B(n52510), .Z(N60713) );
  NAND U62124 ( .A(n52511), .B(n52512), .Z(n52510) );
  NANDN U62125 ( .A(n52513), .B(n52514), .Z(n52512) );
  NANDN U62126 ( .A(n52514), .B(n52513), .Z(n52509) );
  XOR U62127 ( .A(n52513), .B(n52515), .Z(N60712) );
  XNOR U62128 ( .A(n52511), .B(n52514), .Z(n52515) );
  NAND U62129 ( .A(n52516), .B(n52517), .Z(n52514) );
  NAND U62130 ( .A(n52518), .B(n52519), .Z(n52517) );
  NANDN U62131 ( .A(n52520), .B(n52521), .Z(n52519) );
  NANDN U62132 ( .A(n52521), .B(n52520), .Z(n52516) );
  AND U62133 ( .A(n52522), .B(n52523), .Z(n52511) );
  NAND U62134 ( .A(n52524), .B(n52525), .Z(n52523) );
  NANDN U62135 ( .A(n52526), .B(n52527), .Z(n52525) );
  NANDN U62136 ( .A(n52527), .B(n52526), .Z(n52522) );
  IV U62137 ( .A(n52528), .Z(n52527) );
  AND U62138 ( .A(n52529), .B(n52530), .Z(n52513) );
  NAND U62139 ( .A(n52531), .B(n52532), .Z(n52530) );
  NANDN U62140 ( .A(n52533), .B(n52534), .Z(n52532) );
  NANDN U62141 ( .A(n52534), .B(n52533), .Z(n52529) );
  XOR U62142 ( .A(n52526), .B(n52535), .Z(N60711) );
  XNOR U62143 ( .A(n52524), .B(n52528), .Z(n52535) );
  XOR U62144 ( .A(n52521), .B(n52536), .Z(n52528) );
  XNOR U62145 ( .A(n52518), .B(n52520), .Z(n52536) );
  AND U62146 ( .A(n52537), .B(n52538), .Z(n52520) );
  NANDN U62147 ( .A(n52539), .B(n52540), .Z(n52538) );
  OR U62148 ( .A(n52541), .B(n52542), .Z(n52540) );
  IV U62149 ( .A(n52543), .Z(n52542) );
  NANDN U62150 ( .A(n52543), .B(n52541), .Z(n52537) );
  AND U62151 ( .A(n52544), .B(n52545), .Z(n52518) );
  NAND U62152 ( .A(n52546), .B(n52547), .Z(n52545) );
  NANDN U62153 ( .A(n52548), .B(n52549), .Z(n52547) );
  NANDN U62154 ( .A(n52549), .B(n52548), .Z(n52544) );
  IV U62155 ( .A(n52550), .Z(n52549) );
  NAND U62156 ( .A(n52551), .B(n52552), .Z(n52521) );
  NANDN U62157 ( .A(n52553), .B(n52554), .Z(n52552) );
  NANDN U62158 ( .A(n52555), .B(n52556), .Z(n52554) );
  NANDN U62159 ( .A(n52556), .B(n52555), .Z(n52551) );
  IV U62160 ( .A(n52557), .Z(n52555) );
  AND U62161 ( .A(n52558), .B(n52559), .Z(n52524) );
  NAND U62162 ( .A(n52560), .B(n52561), .Z(n52559) );
  NANDN U62163 ( .A(n52562), .B(n52563), .Z(n52561) );
  NANDN U62164 ( .A(n52563), .B(n52562), .Z(n52558) );
  XOR U62165 ( .A(n52534), .B(n52564), .Z(n52526) );
  XNOR U62166 ( .A(n52531), .B(n52533), .Z(n52564) );
  AND U62167 ( .A(n52565), .B(n52566), .Z(n52533) );
  NANDN U62168 ( .A(n52567), .B(n52568), .Z(n52566) );
  OR U62169 ( .A(n52569), .B(n52570), .Z(n52568) );
  IV U62170 ( .A(n52571), .Z(n52570) );
  NANDN U62171 ( .A(n52571), .B(n52569), .Z(n52565) );
  AND U62172 ( .A(n52572), .B(n52573), .Z(n52531) );
  NAND U62173 ( .A(n52574), .B(n52575), .Z(n52573) );
  NANDN U62174 ( .A(n52576), .B(n52577), .Z(n52575) );
  NANDN U62175 ( .A(n52577), .B(n52576), .Z(n52572) );
  IV U62176 ( .A(n52578), .Z(n52577) );
  NAND U62177 ( .A(n52579), .B(n52580), .Z(n52534) );
  NANDN U62178 ( .A(n52581), .B(n52582), .Z(n52580) );
  NANDN U62179 ( .A(n52583), .B(n52584), .Z(n52582) );
  NANDN U62180 ( .A(n52584), .B(n52583), .Z(n52579) );
  IV U62181 ( .A(n52585), .Z(n52583) );
  XOR U62182 ( .A(n52560), .B(n52586), .Z(N60710) );
  XNOR U62183 ( .A(n52563), .B(n52562), .Z(n52586) );
  XNOR U62184 ( .A(n52574), .B(n52587), .Z(n52562) );
  XNOR U62185 ( .A(n52578), .B(n52576), .Z(n52587) );
  XOR U62186 ( .A(n52584), .B(n52588), .Z(n52576) );
  XNOR U62187 ( .A(n52581), .B(n52585), .Z(n52588) );
  AND U62188 ( .A(n52589), .B(n52590), .Z(n52585) );
  NAND U62189 ( .A(n52591), .B(n52592), .Z(n52590) );
  NAND U62190 ( .A(n52593), .B(n52594), .Z(n52589) );
  AND U62191 ( .A(n52595), .B(n52596), .Z(n52581) );
  NAND U62192 ( .A(n52597), .B(n52598), .Z(n52596) );
  NAND U62193 ( .A(n52599), .B(n52600), .Z(n52595) );
  NANDN U62194 ( .A(n52601), .B(n52602), .Z(n52584) );
  ANDN U62195 ( .B(n52603), .A(n52604), .Z(n52578) );
  XNOR U62196 ( .A(n52569), .B(n52605), .Z(n52574) );
  XNOR U62197 ( .A(n52567), .B(n52571), .Z(n52605) );
  AND U62198 ( .A(n52606), .B(n52607), .Z(n52571) );
  NAND U62199 ( .A(n52608), .B(n52609), .Z(n52607) );
  NAND U62200 ( .A(n52610), .B(n52611), .Z(n52606) );
  AND U62201 ( .A(n52612), .B(n52613), .Z(n52567) );
  NAND U62202 ( .A(n52614), .B(n52615), .Z(n52613) );
  NAND U62203 ( .A(n52616), .B(n52617), .Z(n52612) );
  AND U62204 ( .A(n52618), .B(n52619), .Z(n52569) );
  NAND U62205 ( .A(n52620), .B(n52621), .Z(n52563) );
  XNOR U62206 ( .A(n52546), .B(n52622), .Z(n52560) );
  XNOR U62207 ( .A(n52550), .B(n52548), .Z(n52622) );
  XOR U62208 ( .A(n52556), .B(n52623), .Z(n52548) );
  XNOR U62209 ( .A(n52553), .B(n52557), .Z(n52623) );
  AND U62210 ( .A(n52624), .B(n52625), .Z(n52557) );
  NAND U62211 ( .A(n52626), .B(n52627), .Z(n52625) );
  NAND U62212 ( .A(n52628), .B(n52629), .Z(n52624) );
  AND U62213 ( .A(n52630), .B(n52631), .Z(n52553) );
  NAND U62214 ( .A(n52632), .B(n52633), .Z(n52631) );
  NAND U62215 ( .A(n52634), .B(n52635), .Z(n52630) );
  NANDN U62216 ( .A(n52636), .B(n52637), .Z(n52556) );
  ANDN U62217 ( .B(n52638), .A(n52639), .Z(n52550) );
  XNOR U62218 ( .A(n52541), .B(n52640), .Z(n52546) );
  XNOR U62219 ( .A(n52539), .B(n52543), .Z(n52640) );
  AND U62220 ( .A(n52641), .B(n52642), .Z(n52543) );
  NAND U62221 ( .A(n52643), .B(n52644), .Z(n52642) );
  NAND U62222 ( .A(n52645), .B(n52646), .Z(n52641) );
  AND U62223 ( .A(n52647), .B(n52648), .Z(n52539) );
  NAND U62224 ( .A(n52649), .B(n52650), .Z(n52648) );
  NAND U62225 ( .A(n52651), .B(n52652), .Z(n52647) );
  AND U62226 ( .A(n52653), .B(n52654), .Z(n52541) );
  XOR U62227 ( .A(n52621), .B(n52620), .Z(N60709) );
  XNOR U62228 ( .A(n52638), .B(n52639), .Z(n52620) );
  XNOR U62229 ( .A(n52653), .B(n52654), .Z(n52639) );
  XOR U62230 ( .A(n52650), .B(n52649), .Z(n52654) );
  XOR U62231 ( .A(y[228]), .B(x[228]), .Z(n52649) );
  XOR U62232 ( .A(n52652), .B(n52651), .Z(n52650) );
  XOR U62233 ( .A(y[230]), .B(x[230]), .Z(n52651) );
  XOR U62234 ( .A(y[229]), .B(x[229]), .Z(n52652) );
  XOR U62235 ( .A(n52644), .B(n52643), .Z(n52653) );
  XOR U62236 ( .A(n52646), .B(n52645), .Z(n52643) );
  XOR U62237 ( .A(y[227]), .B(x[227]), .Z(n52645) );
  XOR U62238 ( .A(y[226]), .B(x[226]), .Z(n52646) );
  XOR U62239 ( .A(y[225]), .B(x[225]), .Z(n52644) );
  XNOR U62240 ( .A(n52637), .B(n52636), .Z(n52638) );
  XNOR U62241 ( .A(n52633), .B(n52632), .Z(n52636) );
  XOR U62242 ( .A(n52635), .B(n52634), .Z(n52632) );
  XOR U62243 ( .A(y[224]), .B(x[224]), .Z(n52634) );
  XOR U62244 ( .A(y[223]), .B(x[223]), .Z(n52635) );
  XOR U62245 ( .A(y[222]), .B(x[222]), .Z(n52633) );
  XOR U62246 ( .A(n52627), .B(n52626), .Z(n52637) );
  XOR U62247 ( .A(n52629), .B(n52628), .Z(n52626) );
  XOR U62248 ( .A(y[221]), .B(x[221]), .Z(n52628) );
  XOR U62249 ( .A(y[220]), .B(x[220]), .Z(n52629) );
  XOR U62250 ( .A(y[219]), .B(x[219]), .Z(n52627) );
  XNOR U62251 ( .A(n52603), .B(n52604), .Z(n52621) );
  XNOR U62252 ( .A(n52618), .B(n52619), .Z(n52604) );
  XOR U62253 ( .A(n52615), .B(n52614), .Z(n52619) );
  XOR U62254 ( .A(y[216]), .B(x[216]), .Z(n52614) );
  XOR U62255 ( .A(n52617), .B(n52616), .Z(n52615) );
  XOR U62256 ( .A(y[218]), .B(x[218]), .Z(n52616) );
  XOR U62257 ( .A(y[217]), .B(x[217]), .Z(n52617) );
  XOR U62258 ( .A(n52609), .B(n52608), .Z(n52618) );
  XOR U62259 ( .A(n52611), .B(n52610), .Z(n52608) );
  XOR U62260 ( .A(y[215]), .B(x[215]), .Z(n52610) );
  XOR U62261 ( .A(y[214]), .B(x[214]), .Z(n52611) );
  XOR U62262 ( .A(y[213]), .B(x[213]), .Z(n52609) );
  XNOR U62263 ( .A(n52602), .B(n52601), .Z(n52603) );
  XNOR U62264 ( .A(n52598), .B(n52597), .Z(n52601) );
  XOR U62265 ( .A(n52600), .B(n52599), .Z(n52597) );
  XOR U62266 ( .A(y[212]), .B(x[212]), .Z(n52599) );
  XOR U62267 ( .A(y[211]), .B(x[211]), .Z(n52600) );
  XOR U62268 ( .A(y[210]), .B(x[210]), .Z(n52598) );
  XOR U62269 ( .A(n52592), .B(n52591), .Z(n52602) );
  XOR U62270 ( .A(n52594), .B(n52593), .Z(n52591) );
  XOR U62271 ( .A(y[209]), .B(x[209]), .Z(n52593) );
  XOR U62272 ( .A(y[208]), .B(x[208]), .Z(n52594) );
  XOR U62273 ( .A(y[207]), .B(x[207]), .Z(n52592) );
  NAND U62274 ( .A(n52655), .B(n52656), .Z(N60700) );
  NAND U62275 ( .A(n52657), .B(n52658), .Z(n52656) );
  NANDN U62276 ( .A(n52659), .B(n52660), .Z(n52658) );
  NANDN U62277 ( .A(n52660), .B(n52659), .Z(n52655) );
  XOR U62278 ( .A(n52659), .B(n52661), .Z(N60699) );
  XNOR U62279 ( .A(n52657), .B(n52660), .Z(n52661) );
  NAND U62280 ( .A(n52662), .B(n52663), .Z(n52660) );
  NAND U62281 ( .A(n52664), .B(n52665), .Z(n52663) );
  NANDN U62282 ( .A(n52666), .B(n52667), .Z(n52665) );
  NANDN U62283 ( .A(n52667), .B(n52666), .Z(n52662) );
  AND U62284 ( .A(n52668), .B(n52669), .Z(n52657) );
  NAND U62285 ( .A(n52670), .B(n52671), .Z(n52669) );
  NANDN U62286 ( .A(n52672), .B(n52673), .Z(n52671) );
  NANDN U62287 ( .A(n52673), .B(n52672), .Z(n52668) );
  IV U62288 ( .A(n52674), .Z(n52673) );
  AND U62289 ( .A(n52675), .B(n52676), .Z(n52659) );
  NAND U62290 ( .A(n52677), .B(n52678), .Z(n52676) );
  NANDN U62291 ( .A(n52679), .B(n52680), .Z(n52678) );
  NANDN U62292 ( .A(n52680), .B(n52679), .Z(n52675) );
  XOR U62293 ( .A(n52672), .B(n52681), .Z(N60698) );
  XNOR U62294 ( .A(n52670), .B(n52674), .Z(n52681) );
  XOR U62295 ( .A(n52667), .B(n52682), .Z(n52674) );
  XNOR U62296 ( .A(n52664), .B(n52666), .Z(n52682) );
  AND U62297 ( .A(n52683), .B(n52684), .Z(n52666) );
  NANDN U62298 ( .A(n52685), .B(n52686), .Z(n52684) );
  OR U62299 ( .A(n52687), .B(n52688), .Z(n52686) );
  IV U62300 ( .A(n52689), .Z(n52688) );
  NANDN U62301 ( .A(n52689), .B(n52687), .Z(n52683) );
  AND U62302 ( .A(n52690), .B(n52691), .Z(n52664) );
  NAND U62303 ( .A(n52692), .B(n52693), .Z(n52691) );
  NANDN U62304 ( .A(n52694), .B(n52695), .Z(n52693) );
  NANDN U62305 ( .A(n52695), .B(n52694), .Z(n52690) );
  IV U62306 ( .A(n52696), .Z(n52695) );
  NAND U62307 ( .A(n52697), .B(n52698), .Z(n52667) );
  NANDN U62308 ( .A(n52699), .B(n52700), .Z(n52698) );
  NANDN U62309 ( .A(n52701), .B(n52702), .Z(n52700) );
  NANDN U62310 ( .A(n52702), .B(n52701), .Z(n52697) );
  IV U62311 ( .A(n52703), .Z(n52701) );
  AND U62312 ( .A(n52704), .B(n52705), .Z(n52670) );
  NAND U62313 ( .A(n52706), .B(n52707), .Z(n52705) );
  NANDN U62314 ( .A(n52708), .B(n52709), .Z(n52707) );
  NANDN U62315 ( .A(n52709), .B(n52708), .Z(n52704) );
  XOR U62316 ( .A(n52680), .B(n52710), .Z(n52672) );
  XNOR U62317 ( .A(n52677), .B(n52679), .Z(n52710) );
  AND U62318 ( .A(n52711), .B(n52712), .Z(n52679) );
  NANDN U62319 ( .A(n52713), .B(n52714), .Z(n52712) );
  OR U62320 ( .A(n52715), .B(n52716), .Z(n52714) );
  IV U62321 ( .A(n52717), .Z(n52716) );
  NANDN U62322 ( .A(n52717), .B(n52715), .Z(n52711) );
  AND U62323 ( .A(n52718), .B(n52719), .Z(n52677) );
  NAND U62324 ( .A(n52720), .B(n52721), .Z(n52719) );
  NANDN U62325 ( .A(n52722), .B(n52723), .Z(n52721) );
  NANDN U62326 ( .A(n52723), .B(n52722), .Z(n52718) );
  IV U62327 ( .A(n52724), .Z(n52723) );
  NAND U62328 ( .A(n52725), .B(n52726), .Z(n52680) );
  NANDN U62329 ( .A(n52727), .B(n52728), .Z(n52726) );
  NANDN U62330 ( .A(n52729), .B(n52730), .Z(n52728) );
  NANDN U62331 ( .A(n52730), .B(n52729), .Z(n52725) );
  IV U62332 ( .A(n52731), .Z(n52729) );
  XOR U62333 ( .A(n52706), .B(n52732), .Z(N60697) );
  XNOR U62334 ( .A(n52709), .B(n52708), .Z(n52732) );
  XNOR U62335 ( .A(n52720), .B(n52733), .Z(n52708) );
  XNOR U62336 ( .A(n52724), .B(n52722), .Z(n52733) );
  XOR U62337 ( .A(n52730), .B(n52734), .Z(n52722) );
  XNOR U62338 ( .A(n52727), .B(n52731), .Z(n52734) );
  AND U62339 ( .A(n52735), .B(n52736), .Z(n52731) );
  NAND U62340 ( .A(n52737), .B(n52738), .Z(n52736) );
  NAND U62341 ( .A(n52739), .B(n52740), .Z(n52735) );
  AND U62342 ( .A(n52741), .B(n52742), .Z(n52727) );
  NAND U62343 ( .A(n52743), .B(n52744), .Z(n52742) );
  NAND U62344 ( .A(n52745), .B(n52746), .Z(n52741) );
  NANDN U62345 ( .A(n52747), .B(n52748), .Z(n52730) );
  ANDN U62346 ( .B(n52749), .A(n52750), .Z(n52724) );
  XNOR U62347 ( .A(n52715), .B(n52751), .Z(n52720) );
  XNOR U62348 ( .A(n52713), .B(n52717), .Z(n52751) );
  AND U62349 ( .A(n52752), .B(n52753), .Z(n52717) );
  NAND U62350 ( .A(n52754), .B(n52755), .Z(n52753) );
  NAND U62351 ( .A(n52756), .B(n52757), .Z(n52752) );
  AND U62352 ( .A(n52758), .B(n52759), .Z(n52713) );
  NAND U62353 ( .A(n52760), .B(n52761), .Z(n52759) );
  NAND U62354 ( .A(n52762), .B(n52763), .Z(n52758) );
  AND U62355 ( .A(n52764), .B(n52765), .Z(n52715) );
  NAND U62356 ( .A(n52766), .B(n52767), .Z(n52709) );
  XNOR U62357 ( .A(n52692), .B(n52768), .Z(n52706) );
  XNOR U62358 ( .A(n52696), .B(n52694), .Z(n52768) );
  XOR U62359 ( .A(n52702), .B(n52769), .Z(n52694) );
  XNOR U62360 ( .A(n52699), .B(n52703), .Z(n52769) );
  AND U62361 ( .A(n52770), .B(n52771), .Z(n52703) );
  NAND U62362 ( .A(n52772), .B(n52773), .Z(n52771) );
  NAND U62363 ( .A(n52774), .B(n52775), .Z(n52770) );
  AND U62364 ( .A(n52776), .B(n52777), .Z(n52699) );
  NAND U62365 ( .A(n52778), .B(n52779), .Z(n52777) );
  NAND U62366 ( .A(n52780), .B(n52781), .Z(n52776) );
  NANDN U62367 ( .A(n52782), .B(n52783), .Z(n52702) );
  ANDN U62368 ( .B(n52784), .A(n52785), .Z(n52696) );
  XNOR U62369 ( .A(n52687), .B(n52786), .Z(n52692) );
  XNOR U62370 ( .A(n52685), .B(n52689), .Z(n52786) );
  AND U62371 ( .A(n52787), .B(n52788), .Z(n52689) );
  NAND U62372 ( .A(n52789), .B(n52790), .Z(n52788) );
  NAND U62373 ( .A(n52791), .B(n52792), .Z(n52787) );
  AND U62374 ( .A(n52793), .B(n52794), .Z(n52685) );
  NAND U62375 ( .A(n52795), .B(n52796), .Z(n52794) );
  NAND U62376 ( .A(n52797), .B(n52798), .Z(n52793) );
  AND U62377 ( .A(n52799), .B(n52800), .Z(n52687) );
  XOR U62378 ( .A(n52767), .B(n52766), .Z(N60696) );
  XNOR U62379 ( .A(n52784), .B(n52785), .Z(n52766) );
  XNOR U62380 ( .A(n52799), .B(n52800), .Z(n52785) );
  XOR U62381 ( .A(n52796), .B(n52795), .Z(n52800) );
  XOR U62382 ( .A(y[204]), .B(x[204]), .Z(n52795) );
  XOR U62383 ( .A(n52798), .B(n52797), .Z(n52796) );
  XOR U62384 ( .A(y[206]), .B(x[206]), .Z(n52797) );
  XOR U62385 ( .A(y[205]), .B(x[205]), .Z(n52798) );
  XOR U62386 ( .A(n52790), .B(n52789), .Z(n52799) );
  XOR U62387 ( .A(n52792), .B(n52791), .Z(n52789) );
  XOR U62388 ( .A(y[203]), .B(x[203]), .Z(n52791) );
  XOR U62389 ( .A(y[202]), .B(x[202]), .Z(n52792) );
  XOR U62390 ( .A(y[201]), .B(x[201]), .Z(n52790) );
  XNOR U62391 ( .A(n52783), .B(n52782), .Z(n52784) );
  XNOR U62392 ( .A(n52779), .B(n52778), .Z(n52782) );
  XOR U62393 ( .A(n52781), .B(n52780), .Z(n52778) );
  XOR U62394 ( .A(y[200]), .B(x[200]), .Z(n52780) );
  XOR U62395 ( .A(y[199]), .B(x[199]), .Z(n52781) );
  XOR U62396 ( .A(y[198]), .B(x[198]), .Z(n52779) );
  XOR U62397 ( .A(n52773), .B(n52772), .Z(n52783) );
  XOR U62398 ( .A(n52775), .B(n52774), .Z(n52772) );
  XOR U62399 ( .A(y[197]), .B(x[197]), .Z(n52774) );
  XOR U62400 ( .A(y[196]), .B(x[196]), .Z(n52775) );
  XOR U62401 ( .A(y[195]), .B(x[195]), .Z(n52773) );
  XNOR U62402 ( .A(n52749), .B(n52750), .Z(n52767) );
  XNOR U62403 ( .A(n52764), .B(n52765), .Z(n52750) );
  XOR U62404 ( .A(n52761), .B(n52760), .Z(n52765) );
  XOR U62405 ( .A(y[192]), .B(x[192]), .Z(n52760) );
  XOR U62406 ( .A(n52763), .B(n52762), .Z(n52761) );
  XOR U62407 ( .A(y[194]), .B(x[194]), .Z(n52762) );
  XOR U62408 ( .A(y[193]), .B(x[193]), .Z(n52763) );
  XOR U62409 ( .A(n52755), .B(n52754), .Z(n52764) );
  XOR U62410 ( .A(n52757), .B(n52756), .Z(n52754) );
  XOR U62411 ( .A(y[191]), .B(x[191]), .Z(n52756) );
  XOR U62412 ( .A(y[190]), .B(x[190]), .Z(n52757) );
  XOR U62413 ( .A(y[189]), .B(x[189]), .Z(n52755) );
  XNOR U62414 ( .A(n52748), .B(n52747), .Z(n52749) );
  XNOR U62415 ( .A(n52744), .B(n52743), .Z(n52747) );
  XOR U62416 ( .A(n52746), .B(n52745), .Z(n52743) );
  XOR U62417 ( .A(y[188]), .B(x[188]), .Z(n52745) );
  XOR U62418 ( .A(y[187]), .B(x[187]), .Z(n52746) );
  XOR U62419 ( .A(y[186]), .B(x[186]), .Z(n52744) );
  XOR U62420 ( .A(n52738), .B(n52737), .Z(n52748) );
  XOR U62421 ( .A(n52740), .B(n52739), .Z(n52737) );
  XOR U62422 ( .A(y[185]), .B(x[185]), .Z(n52739) );
  XOR U62423 ( .A(y[184]), .B(x[184]), .Z(n52740) );
  XOR U62424 ( .A(y[183]), .B(x[183]), .Z(n52738) );
  NAND U62425 ( .A(n52801), .B(n52802), .Z(N60687) );
  NAND U62426 ( .A(n52803), .B(n52804), .Z(n52802) );
  NANDN U62427 ( .A(n52805), .B(n52806), .Z(n52804) );
  NANDN U62428 ( .A(n52806), .B(n52805), .Z(n52801) );
  XOR U62429 ( .A(n52805), .B(n52807), .Z(N60686) );
  XNOR U62430 ( .A(n52803), .B(n52806), .Z(n52807) );
  NAND U62431 ( .A(n52808), .B(n52809), .Z(n52806) );
  NAND U62432 ( .A(n52810), .B(n52811), .Z(n52809) );
  NANDN U62433 ( .A(n52812), .B(n52813), .Z(n52811) );
  NANDN U62434 ( .A(n52813), .B(n52812), .Z(n52808) );
  AND U62435 ( .A(n52814), .B(n52815), .Z(n52803) );
  NAND U62436 ( .A(n52816), .B(n52817), .Z(n52815) );
  NANDN U62437 ( .A(n52818), .B(n52819), .Z(n52817) );
  NANDN U62438 ( .A(n52819), .B(n52818), .Z(n52814) );
  IV U62439 ( .A(n52820), .Z(n52819) );
  AND U62440 ( .A(n52821), .B(n52822), .Z(n52805) );
  NAND U62441 ( .A(n52823), .B(n52824), .Z(n52822) );
  NANDN U62442 ( .A(n52825), .B(n52826), .Z(n52824) );
  NANDN U62443 ( .A(n52826), .B(n52825), .Z(n52821) );
  XOR U62444 ( .A(n52818), .B(n52827), .Z(N60685) );
  XNOR U62445 ( .A(n52816), .B(n52820), .Z(n52827) );
  XOR U62446 ( .A(n52813), .B(n52828), .Z(n52820) );
  XNOR U62447 ( .A(n52810), .B(n52812), .Z(n52828) );
  AND U62448 ( .A(n52829), .B(n52830), .Z(n52812) );
  NANDN U62449 ( .A(n52831), .B(n52832), .Z(n52830) );
  OR U62450 ( .A(n52833), .B(n52834), .Z(n52832) );
  IV U62451 ( .A(n52835), .Z(n52834) );
  NANDN U62452 ( .A(n52835), .B(n52833), .Z(n52829) );
  AND U62453 ( .A(n52836), .B(n52837), .Z(n52810) );
  NAND U62454 ( .A(n52838), .B(n52839), .Z(n52837) );
  NANDN U62455 ( .A(n52840), .B(n52841), .Z(n52839) );
  NANDN U62456 ( .A(n52841), .B(n52840), .Z(n52836) );
  IV U62457 ( .A(n52842), .Z(n52841) );
  NAND U62458 ( .A(n52843), .B(n52844), .Z(n52813) );
  NANDN U62459 ( .A(n52845), .B(n52846), .Z(n52844) );
  NANDN U62460 ( .A(n52847), .B(n52848), .Z(n52846) );
  NANDN U62461 ( .A(n52848), .B(n52847), .Z(n52843) );
  IV U62462 ( .A(n52849), .Z(n52847) );
  AND U62463 ( .A(n52850), .B(n52851), .Z(n52816) );
  NAND U62464 ( .A(n52852), .B(n52853), .Z(n52851) );
  NANDN U62465 ( .A(n52854), .B(n52855), .Z(n52853) );
  NANDN U62466 ( .A(n52855), .B(n52854), .Z(n52850) );
  XOR U62467 ( .A(n52826), .B(n52856), .Z(n52818) );
  XNOR U62468 ( .A(n52823), .B(n52825), .Z(n52856) );
  AND U62469 ( .A(n52857), .B(n52858), .Z(n52825) );
  NANDN U62470 ( .A(n52859), .B(n52860), .Z(n52858) );
  OR U62471 ( .A(n52861), .B(n52862), .Z(n52860) );
  IV U62472 ( .A(n52863), .Z(n52862) );
  NANDN U62473 ( .A(n52863), .B(n52861), .Z(n52857) );
  AND U62474 ( .A(n52864), .B(n52865), .Z(n52823) );
  NAND U62475 ( .A(n52866), .B(n52867), .Z(n52865) );
  NANDN U62476 ( .A(n52868), .B(n52869), .Z(n52867) );
  NANDN U62477 ( .A(n52869), .B(n52868), .Z(n52864) );
  IV U62478 ( .A(n52870), .Z(n52869) );
  NAND U62479 ( .A(n52871), .B(n52872), .Z(n52826) );
  NANDN U62480 ( .A(n52873), .B(n52874), .Z(n52872) );
  NANDN U62481 ( .A(n52875), .B(n52876), .Z(n52874) );
  NANDN U62482 ( .A(n52876), .B(n52875), .Z(n52871) );
  IV U62483 ( .A(n52877), .Z(n52875) );
  XOR U62484 ( .A(n52852), .B(n52878), .Z(N60684) );
  XNOR U62485 ( .A(n52855), .B(n52854), .Z(n52878) );
  XNOR U62486 ( .A(n52866), .B(n52879), .Z(n52854) );
  XNOR U62487 ( .A(n52870), .B(n52868), .Z(n52879) );
  XOR U62488 ( .A(n52876), .B(n52880), .Z(n52868) );
  XNOR U62489 ( .A(n52873), .B(n52877), .Z(n52880) );
  AND U62490 ( .A(n52881), .B(n52882), .Z(n52877) );
  NAND U62491 ( .A(n52883), .B(n52884), .Z(n52882) );
  NAND U62492 ( .A(n52885), .B(n52886), .Z(n52881) );
  AND U62493 ( .A(n52887), .B(n52888), .Z(n52873) );
  NAND U62494 ( .A(n52889), .B(n52890), .Z(n52888) );
  NAND U62495 ( .A(n52891), .B(n52892), .Z(n52887) );
  NANDN U62496 ( .A(n52893), .B(n52894), .Z(n52876) );
  ANDN U62497 ( .B(n52895), .A(n52896), .Z(n52870) );
  XNOR U62498 ( .A(n52861), .B(n52897), .Z(n52866) );
  XNOR U62499 ( .A(n52859), .B(n52863), .Z(n52897) );
  AND U62500 ( .A(n52898), .B(n52899), .Z(n52863) );
  NAND U62501 ( .A(n52900), .B(n52901), .Z(n52899) );
  NAND U62502 ( .A(n52902), .B(n52903), .Z(n52898) );
  AND U62503 ( .A(n52904), .B(n52905), .Z(n52859) );
  NAND U62504 ( .A(n52906), .B(n52907), .Z(n52905) );
  NAND U62505 ( .A(n52908), .B(n52909), .Z(n52904) );
  AND U62506 ( .A(n52910), .B(n52911), .Z(n52861) );
  NAND U62507 ( .A(n52912), .B(n52913), .Z(n52855) );
  XNOR U62508 ( .A(n52838), .B(n52914), .Z(n52852) );
  XNOR U62509 ( .A(n52842), .B(n52840), .Z(n52914) );
  XOR U62510 ( .A(n52848), .B(n52915), .Z(n52840) );
  XNOR U62511 ( .A(n52845), .B(n52849), .Z(n52915) );
  AND U62512 ( .A(n52916), .B(n52917), .Z(n52849) );
  NAND U62513 ( .A(n52918), .B(n52919), .Z(n52917) );
  NAND U62514 ( .A(n52920), .B(n52921), .Z(n52916) );
  AND U62515 ( .A(n52922), .B(n52923), .Z(n52845) );
  NAND U62516 ( .A(n52924), .B(n52925), .Z(n52923) );
  NAND U62517 ( .A(n52926), .B(n52927), .Z(n52922) );
  NANDN U62518 ( .A(n52928), .B(n52929), .Z(n52848) );
  ANDN U62519 ( .B(n52930), .A(n52931), .Z(n52842) );
  XNOR U62520 ( .A(n52833), .B(n52932), .Z(n52838) );
  XNOR U62521 ( .A(n52831), .B(n52835), .Z(n52932) );
  AND U62522 ( .A(n52933), .B(n52934), .Z(n52835) );
  NAND U62523 ( .A(n52935), .B(n52936), .Z(n52934) );
  NAND U62524 ( .A(n52937), .B(n52938), .Z(n52933) );
  AND U62525 ( .A(n52939), .B(n52940), .Z(n52831) );
  NAND U62526 ( .A(n52941), .B(n52942), .Z(n52940) );
  NAND U62527 ( .A(n52943), .B(n52944), .Z(n52939) );
  AND U62528 ( .A(n52945), .B(n52946), .Z(n52833) );
  XOR U62529 ( .A(n52913), .B(n52912), .Z(N60683) );
  XNOR U62530 ( .A(n52930), .B(n52931), .Z(n52912) );
  XNOR U62531 ( .A(n52945), .B(n52946), .Z(n52931) );
  XOR U62532 ( .A(n52942), .B(n52941), .Z(n52946) );
  XOR U62533 ( .A(y[180]), .B(x[180]), .Z(n52941) );
  XOR U62534 ( .A(n52944), .B(n52943), .Z(n52942) );
  XOR U62535 ( .A(y[182]), .B(x[182]), .Z(n52943) );
  XOR U62536 ( .A(y[181]), .B(x[181]), .Z(n52944) );
  XOR U62537 ( .A(n52936), .B(n52935), .Z(n52945) );
  XOR U62538 ( .A(n52938), .B(n52937), .Z(n52935) );
  XOR U62539 ( .A(y[179]), .B(x[179]), .Z(n52937) );
  XOR U62540 ( .A(y[178]), .B(x[178]), .Z(n52938) );
  XOR U62541 ( .A(y[177]), .B(x[177]), .Z(n52936) );
  XNOR U62542 ( .A(n52929), .B(n52928), .Z(n52930) );
  XNOR U62543 ( .A(n52925), .B(n52924), .Z(n52928) );
  XOR U62544 ( .A(n52927), .B(n52926), .Z(n52924) );
  XOR U62545 ( .A(y[176]), .B(x[176]), .Z(n52926) );
  XOR U62546 ( .A(y[175]), .B(x[175]), .Z(n52927) );
  XOR U62547 ( .A(y[174]), .B(x[174]), .Z(n52925) );
  XOR U62548 ( .A(n52919), .B(n52918), .Z(n52929) );
  XOR U62549 ( .A(n52921), .B(n52920), .Z(n52918) );
  XOR U62550 ( .A(y[173]), .B(x[173]), .Z(n52920) );
  XOR U62551 ( .A(y[172]), .B(x[172]), .Z(n52921) );
  XOR U62552 ( .A(y[171]), .B(x[171]), .Z(n52919) );
  XNOR U62553 ( .A(n52895), .B(n52896), .Z(n52913) );
  XNOR U62554 ( .A(n52910), .B(n52911), .Z(n52896) );
  XOR U62555 ( .A(n52907), .B(n52906), .Z(n52911) );
  XOR U62556 ( .A(y[168]), .B(x[168]), .Z(n52906) );
  XOR U62557 ( .A(n52909), .B(n52908), .Z(n52907) );
  XOR U62558 ( .A(y[170]), .B(x[170]), .Z(n52908) );
  XOR U62559 ( .A(y[169]), .B(x[169]), .Z(n52909) );
  XOR U62560 ( .A(n52901), .B(n52900), .Z(n52910) );
  XOR U62561 ( .A(n52903), .B(n52902), .Z(n52900) );
  XOR U62562 ( .A(y[167]), .B(x[167]), .Z(n52902) );
  XOR U62563 ( .A(y[166]), .B(x[166]), .Z(n52903) );
  XOR U62564 ( .A(y[165]), .B(x[165]), .Z(n52901) );
  XNOR U62565 ( .A(n52894), .B(n52893), .Z(n52895) );
  XNOR U62566 ( .A(n52890), .B(n52889), .Z(n52893) );
  XOR U62567 ( .A(n52892), .B(n52891), .Z(n52889) );
  XOR U62568 ( .A(y[164]), .B(x[164]), .Z(n52891) );
  XOR U62569 ( .A(y[163]), .B(x[163]), .Z(n52892) );
  XOR U62570 ( .A(y[162]), .B(x[162]), .Z(n52890) );
  XOR U62571 ( .A(n52884), .B(n52883), .Z(n52894) );
  XOR U62572 ( .A(n52886), .B(n52885), .Z(n52883) );
  XOR U62573 ( .A(y[161]), .B(x[161]), .Z(n52885) );
  XOR U62574 ( .A(y[160]), .B(x[160]), .Z(n52886) );
  XOR U62575 ( .A(y[159]), .B(x[159]), .Z(n52884) );
  NAND U62576 ( .A(n52947), .B(n52948), .Z(N60674) );
  NAND U62577 ( .A(n52949), .B(n52950), .Z(n52948) );
  NANDN U62578 ( .A(n52951), .B(n52952), .Z(n52950) );
  NANDN U62579 ( .A(n52952), .B(n52951), .Z(n52947) );
  XOR U62580 ( .A(n52951), .B(n52953), .Z(N60673) );
  XNOR U62581 ( .A(n52949), .B(n52952), .Z(n52953) );
  NAND U62582 ( .A(n52954), .B(n52955), .Z(n52952) );
  NAND U62583 ( .A(n52956), .B(n52957), .Z(n52955) );
  NANDN U62584 ( .A(n52958), .B(n52959), .Z(n52957) );
  NANDN U62585 ( .A(n52959), .B(n52958), .Z(n52954) );
  AND U62586 ( .A(n52960), .B(n52961), .Z(n52949) );
  NAND U62587 ( .A(n52962), .B(n52963), .Z(n52961) );
  NANDN U62588 ( .A(n52964), .B(n52965), .Z(n52963) );
  NANDN U62589 ( .A(n52965), .B(n52964), .Z(n52960) );
  IV U62590 ( .A(n52966), .Z(n52965) );
  AND U62591 ( .A(n52967), .B(n52968), .Z(n52951) );
  NAND U62592 ( .A(n52969), .B(n52970), .Z(n52968) );
  NANDN U62593 ( .A(n52971), .B(n52972), .Z(n52970) );
  NANDN U62594 ( .A(n52972), .B(n52971), .Z(n52967) );
  XOR U62595 ( .A(n52964), .B(n52973), .Z(N60672) );
  XNOR U62596 ( .A(n52962), .B(n52966), .Z(n52973) );
  XOR U62597 ( .A(n52959), .B(n52974), .Z(n52966) );
  XNOR U62598 ( .A(n52956), .B(n52958), .Z(n52974) );
  AND U62599 ( .A(n52975), .B(n52976), .Z(n52958) );
  NANDN U62600 ( .A(n52977), .B(n52978), .Z(n52976) );
  OR U62601 ( .A(n52979), .B(n52980), .Z(n52978) );
  IV U62602 ( .A(n52981), .Z(n52980) );
  NANDN U62603 ( .A(n52981), .B(n52979), .Z(n52975) );
  AND U62604 ( .A(n52982), .B(n52983), .Z(n52956) );
  NAND U62605 ( .A(n52984), .B(n52985), .Z(n52983) );
  NANDN U62606 ( .A(n52986), .B(n52987), .Z(n52985) );
  NANDN U62607 ( .A(n52987), .B(n52986), .Z(n52982) );
  IV U62608 ( .A(n52988), .Z(n52987) );
  NAND U62609 ( .A(n52989), .B(n52990), .Z(n52959) );
  NANDN U62610 ( .A(n52991), .B(n52992), .Z(n52990) );
  NANDN U62611 ( .A(n52993), .B(n52994), .Z(n52992) );
  NANDN U62612 ( .A(n52994), .B(n52993), .Z(n52989) );
  IV U62613 ( .A(n52995), .Z(n52993) );
  AND U62614 ( .A(n52996), .B(n52997), .Z(n52962) );
  NAND U62615 ( .A(n52998), .B(n52999), .Z(n52997) );
  NANDN U62616 ( .A(n53000), .B(n53001), .Z(n52999) );
  NANDN U62617 ( .A(n53001), .B(n53000), .Z(n52996) );
  XOR U62618 ( .A(n52972), .B(n53002), .Z(n52964) );
  XNOR U62619 ( .A(n52969), .B(n52971), .Z(n53002) );
  AND U62620 ( .A(n53003), .B(n53004), .Z(n52971) );
  NANDN U62621 ( .A(n53005), .B(n53006), .Z(n53004) );
  OR U62622 ( .A(n53007), .B(n53008), .Z(n53006) );
  IV U62623 ( .A(n53009), .Z(n53008) );
  NANDN U62624 ( .A(n53009), .B(n53007), .Z(n53003) );
  AND U62625 ( .A(n53010), .B(n53011), .Z(n52969) );
  NAND U62626 ( .A(n53012), .B(n53013), .Z(n53011) );
  NANDN U62627 ( .A(n53014), .B(n53015), .Z(n53013) );
  NANDN U62628 ( .A(n53015), .B(n53014), .Z(n53010) );
  IV U62629 ( .A(n53016), .Z(n53015) );
  NAND U62630 ( .A(n53017), .B(n53018), .Z(n52972) );
  NANDN U62631 ( .A(n53019), .B(n53020), .Z(n53018) );
  NANDN U62632 ( .A(n53021), .B(n53022), .Z(n53020) );
  NANDN U62633 ( .A(n53022), .B(n53021), .Z(n53017) );
  IV U62634 ( .A(n53023), .Z(n53021) );
  XOR U62635 ( .A(n52998), .B(n53024), .Z(N60671) );
  XNOR U62636 ( .A(n53001), .B(n53000), .Z(n53024) );
  XNOR U62637 ( .A(n53012), .B(n53025), .Z(n53000) );
  XNOR U62638 ( .A(n53016), .B(n53014), .Z(n53025) );
  XOR U62639 ( .A(n53022), .B(n53026), .Z(n53014) );
  XNOR U62640 ( .A(n53019), .B(n53023), .Z(n53026) );
  AND U62641 ( .A(n53027), .B(n53028), .Z(n53023) );
  NAND U62642 ( .A(n53029), .B(n53030), .Z(n53028) );
  NAND U62643 ( .A(n53031), .B(n53032), .Z(n53027) );
  AND U62644 ( .A(n53033), .B(n53034), .Z(n53019) );
  NAND U62645 ( .A(n53035), .B(n53036), .Z(n53034) );
  NAND U62646 ( .A(n53037), .B(n53038), .Z(n53033) );
  NANDN U62647 ( .A(n53039), .B(n53040), .Z(n53022) );
  ANDN U62648 ( .B(n53041), .A(n53042), .Z(n53016) );
  XNOR U62649 ( .A(n53007), .B(n53043), .Z(n53012) );
  XNOR U62650 ( .A(n53005), .B(n53009), .Z(n53043) );
  AND U62651 ( .A(n53044), .B(n53045), .Z(n53009) );
  NAND U62652 ( .A(n53046), .B(n53047), .Z(n53045) );
  NAND U62653 ( .A(n53048), .B(n53049), .Z(n53044) );
  AND U62654 ( .A(n53050), .B(n53051), .Z(n53005) );
  NAND U62655 ( .A(n53052), .B(n53053), .Z(n53051) );
  NAND U62656 ( .A(n53054), .B(n53055), .Z(n53050) );
  AND U62657 ( .A(n53056), .B(n53057), .Z(n53007) );
  NAND U62658 ( .A(n53058), .B(n53059), .Z(n53001) );
  XNOR U62659 ( .A(n52984), .B(n53060), .Z(n52998) );
  XNOR U62660 ( .A(n52988), .B(n52986), .Z(n53060) );
  XOR U62661 ( .A(n52994), .B(n53061), .Z(n52986) );
  XNOR U62662 ( .A(n52991), .B(n52995), .Z(n53061) );
  AND U62663 ( .A(n53062), .B(n53063), .Z(n52995) );
  NAND U62664 ( .A(n53064), .B(n53065), .Z(n53063) );
  NAND U62665 ( .A(n53066), .B(n53067), .Z(n53062) );
  AND U62666 ( .A(n53068), .B(n53069), .Z(n52991) );
  NAND U62667 ( .A(n53070), .B(n53071), .Z(n53069) );
  NAND U62668 ( .A(n53072), .B(n53073), .Z(n53068) );
  NANDN U62669 ( .A(n53074), .B(n53075), .Z(n52994) );
  ANDN U62670 ( .B(n53076), .A(n53077), .Z(n52988) );
  XNOR U62671 ( .A(n52979), .B(n53078), .Z(n52984) );
  XNOR U62672 ( .A(n52977), .B(n52981), .Z(n53078) );
  AND U62673 ( .A(n53079), .B(n53080), .Z(n52981) );
  NAND U62674 ( .A(n53081), .B(n53082), .Z(n53080) );
  NAND U62675 ( .A(n53083), .B(n53084), .Z(n53079) );
  AND U62676 ( .A(n53085), .B(n53086), .Z(n52977) );
  NAND U62677 ( .A(n53087), .B(n53088), .Z(n53086) );
  NAND U62678 ( .A(n53089), .B(n53090), .Z(n53085) );
  AND U62679 ( .A(n53091), .B(n53092), .Z(n52979) );
  XOR U62680 ( .A(n53059), .B(n53058), .Z(N60670) );
  XNOR U62681 ( .A(n53076), .B(n53077), .Z(n53058) );
  XNOR U62682 ( .A(n53091), .B(n53092), .Z(n53077) );
  XOR U62683 ( .A(n53088), .B(n53087), .Z(n53092) );
  XOR U62684 ( .A(y[156]), .B(x[156]), .Z(n53087) );
  XOR U62685 ( .A(n53090), .B(n53089), .Z(n53088) );
  XOR U62686 ( .A(y[158]), .B(x[158]), .Z(n53089) );
  XOR U62687 ( .A(y[157]), .B(x[157]), .Z(n53090) );
  XOR U62688 ( .A(n53082), .B(n53081), .Z(n53091) );
  XOR U62689 ( .A(n53084), .B(n53083), .Z(n53081) );
  XOR U62690 ( .A(y[155]), .B(x[155]), .Z(n53083) );
  XOR U62691 ( .A(y[154]), .B(x[154]), .Z(n53084) );
  XOR U62692 ( .A(y[153]), .B(x[153]), .Z(n53082) );
  XNOR U62693 ( .A(n53075), .B(n53074), .Z(n53076) );
  XNOR U62694 ( .A(n53071), .B(n53070), .Z(n53074) );
  XOR U62695 ( .A(n53073), .B(n53072), .Z(n53070) );
  XOR U62696 ( .A(y[152]), .B(x[152]), .Z(n53072) );
  XOR U62697 ( .A(y[151]), .B(x[151]), .Z(n53073) );
  XOR U62698 ( .A(y[150]), .B(x[150]), .Z(n53071) );
  XOR U62699 ( .A(n53065), .B(n53064), .Z(n53075) );
  XOR U62700 ( .A(n53067), .B(n53066), .Z(n53064) );
  XOR U62701 ( .A(y[149]), .B(x[149]), .Z(n53066) );
  XOR U62702 ( .A(y[148]), .B(x[148]), .Z(n53067) );
  XOR U62703 ( .A(y[147]), .B(x[147]), .Z(n53065) );
  XNOR U62704 ( .A(n53041), .B(n53042), .Z(n53059) );
  XNOR U62705 ( .A(n53056), .B(n53057), .Z(n53042) );
  XOR U62706 ( .A(n53053), .B(n53052), .Z(n53057) );
  XOR U62707 ( .A(y[144]), .B(x[144]), .Z(n53052) );
  XOR U62708 ( .A(n53055), .B(n53054), .Z(n53053) );
  XOR U62709 ( .A(y[146]), .B(x[146]), .Z(n53054) );
  XOR U62710 ( .A(y[145]), .B(x[145]), .Z(n53055) );
  XOR U62711 ( .A(n53047), .B(n53046), .Z(n53056) );
  XOR U62712 ( .A(n53049), .B(n53048), .Z(n53046) );
  XOR U62713 ( .A(y[143]), .B(x[143]), .Z(n53048) );
  XOR U62714 ( .A(y[142]), .B(x[142]), .Z(n53049) );
  XOR U62715 ( .A(y[141]), .B(x[141]), .Z(n53047) );
  XNOR U62716 ( .A(n53040), .B(n53039), .Z(n53041) );
  XNOR U62717 ( .A(n53036), .B(n53035), .Z(n53039) );
  XOR U62718 ( .A(n53038), .B(n53037), .Z(n53035) );
  XOR U62719 ( .A(y[140]), .B(x[140]), .Z(n53037) );
  XOR U62720 ( .A(y[139]), .B(x[139]), .Z(n53038) );
  XOR U62721 ( .A(y[138]), .B(x[138]), .Z(n53036) );
  XOR U62722 ( .A(n53030), .B(n53029), .Z(n53040) );
  XOR U62723 ( .A(n53032), .B(n53031), .Z(n53029) );
  XOR U62724 ( .A(y[137]), .B(x[137]), .Z(n53031) );
  XOR U62725 ( .A(y[136]), .B(x[136]), .Z(n53032) );
  XOR U62726 ( .A(y[135]), .B(x[135]), .Z(n53030) );
  NAND U62727 ( .A(n53093), .B(n53094), .Z(N60661) );
  NAND U62728 ( .A(n53095), .B(n53096), .Z(n53094) );
  NANDN U62729 ( .A(n53097), .B(n53098), .Z(n53096) );
  NANDN U62730 ( .A(n53098), .B(n53097), .Z(n53093) );
  XOR U62731 ( .A(n53097), .B(n53099), .Z(N60660) );
  XNOR U62732 ( .A(n53095), .B(n53098), .Z(n53099) );
  NAND U62733 ( .A(n53100), .B(n53101), .Z(n53098) );
  NAND U62734 ( .A(n53102), .B(n53103), .Z(n53101) );
  NANDN U62735 ( .A(n53104), .B(n53105), .Z(n53103) );
  NANDN U62736 ( .A(n53105), .B(n53104), .Z(n53100) );
  AND U62737 ( .A(n53106), .B(n53107), .Z(n53095) );
  NAND U62738 ( .A(n53108), .B(n53109), .Z(n53107) );
  NANDN U62739 ( .A(n53110), .B(n53111), .Z(n53109) );
  NANDN U62740 ( .A(n53111), .B(n53110), .Z(n53106) );
  IV U62741 ( .A(n53112), .Z(n53111) );
  AND U62742 ( .A(n53113), .B(n53114), .Z(n53097) );
  NAND U62743 ( .A(n53115), .B(n53116), .Z(n53114) );
  NANDN U62744 ( .A(n53117), .B(n53118), .Z(n53116) );
  NANDN U62745 ( .A(n53118), .B(n53117), .Z(n53113) );
  XOR U62746 ( .A(n53110), .B(n53119), .Z(N60659) );
  XNOR U62747 ( .A(n53108), .B(n53112), .Z(n53119) );
  XOR U62748 ( .A(n53105), .B(n53120), .Z(n53112) );
  XNOR U62749 ( .A(n53102), .B(n53104), .Z(n53120) );
  AND U62750 ( .A(n53121), .B(n53122), .Z(n53104) );
  NANDN U62751 ( .A(n53123), .B(n53124), .Z(n53122) );
  OR U62752 ( .A(n53125), .B(n53126), .Z(n53124) );
  IV U62753 ( .A(n53127), .Z(n53126) );
  NANDN U62754 ( .A(n53127), .B(n53125), .Z(n53121) );
  AND U62755 ( .A(n53128), .B(n53129), .Z(n53102) );
  NAND U62756 ( .A(n53130), .B(n53131), .Z(n53129) );
  NANDN U62757 ( .A(n53132), .B(n53133), .Z(n53131) );
  NANDN U62758 ( .A(n53133), .B(n53132), .Z(n53128) );
  IV U62759 ( .A(n53134), .Z(n53133) );
  NAND U62760 ( .A(n53135), .B(n53136), .Z(n53105) );
  NANDN U62761 ( .A(n53137), .B(n53138), .Z(n53136) );
  NANDN U62762 ( .A(n53139), .B(n53140), .Z(n53138) );
  NANDN U62763 ( .A(n53140), .B(n53139), .Z(n53135) );
  IV U62764 ( .A(n53141), .Z(n53139) );
  AND U62765 ( .A(n53142), .B(n53143), .Z(n53108) );
  NAND U62766 ( .A(n53144), .B(n53145), .Z(n53143) );
  NANDN U62767 ( .A(n53146), .B(n53147), .Z(n53145) );
  NANDN U62768 ( .A(n53147), .B(n53146), .Z(n53142) );
  XOR U62769 ( .A(n53118), .B(n53148), .Z(n53110) );
  XNOR U62770 ( .A(n53115), .B(n53117), .Z(n53148) );
  AND U62771 ( .A(n53149), .B(n53150), .Z(n53117) );
  NANDN U62772 ( .A(n53151), .B(n53152), .Z(n53150) );
  OR U62773 ( .A(n53153), .B(n53154), .Z(n53152) );
  IV U62774 ( .A(n53155), .Z(n53154) );
  NANDN U62775 ( .A(n53155), .B(n53153), .Z(n53149) );
  AND U62776 ( .A(n53156), .B(n53157), .Z(n53115) );
  NAND U62777 ( .A(n53158), .B(n53159), .Z(n53157) );
  NANDN U62778 ( .A(n53160), .B(n53161), .Z(n53159) );
  NANDN U62779 ( .A(n53161), .B(n53160), .Z(n53156) );
  IV U62780 ( .A(n53162), .Z(n53161) );
  NAND U62781 ( .A(n53163), .B(n53164), .Z(n53118) );
  NANDN U62782 ( .A(n53165), .B(n53166), .Z(n53164) );
  NANDN U62783 ( .A(n53167), .B(n53168), .Z(n53166) );
  NANDN U62784 ( .A(n53168), .B(n53167), .Z(n53163) );
  IV U62785 ( .A(n53169), .Z(n53167) );
  XOR U62786 ( .A(n53144), .B(n53170), .Z(N60658) );
  XNOR U62787 ( .A(n53147), .B(n53146), .Z(n53170) );
  XNOR U62788 ( .A(n53158), .B(n53171), .Z(n53146) );
  XNOR U62789 ( .A(n53162), .B(n53160), .Z(n53171) );
  XOR U62790 ( .A(n53168), .B(n53172), .Z(n53160) );
  XNOR U62791 ( .A(n53165), .B(n53169), .Z(n53172) );
  AND U62792 ( .A(n53173), .B(n53174), .Z(n53169) );
  NAND U62793 ( .A(n53175), .B(n53176), .Z(n53174) );
  NAND U62794 ( .A(n53177), .B(n53178), .Z(n53173) );
  AND U62795 ( .A(n53179), .B(n53180), .Z(n53165) );
  NAND U62796 ( .A(n53181), .B(n53182), .Z(n53180) );
  NAND U62797 ( .A(n53183), .B(n53184), .Z(n53179) );
  NANDN U62798 ( .A(n53185), .B(n53186), .Z(n53168) );
  ANDN U62799 ( .B(n53187), .A(n53188), .Z(n53162) );
  XNOR U62800 ( .A(n53153), .B(n53189), .Z(n53158) );
  XNOR U62801 ( .A(n53151), .B(n53155), .Z(n53189) );
  AND U62802 ( .A(n53190), .B(n53191), .Z(n53155) );
  NAND U62803 ( .A(n53192), .B(n53193), .Z(n53191) );
  NAND U62804 ( .A(n53194), .B(n53195), .Z(n53190) );
  AND U62805 ( .A(n53196), .B(n53197), .Z(n53151) );
  NAND U62806 ( .A(n53198), .B(n53199), .Z(n53197) );
  NAND U62807 ( .A(n53200), .B(n53201), .Z(n53196) );
  AND U62808 ( .A(n53202), .B(n53203), .Z(n53153) );
  NAND U62809 ( .A(n53204), .B(n53205), .Z(n53147) );
  XNOR U62810 ( .A(n53130), .B(n53206), .Z(n53144) );
  XNOR U62811 ( .A(n53134), .B(n53132), .Z(n53206) );
  XOR U62812 ( .A(n53140), .B(n53207), .Z(n53132) );
  XNOR U62813 ( .A(n53137), .B(n53141), .Z(n53207) );
  AND U62814 ( .A(n53208), .B(n53209), .Z(n53141) );
  NAND U62815 ( .A(n53210), .B(n53211), .Z(n53209) );
  NAND U62816 ( .A(n53212), .B(n53213), .Z(n53208) );
  AND U62817 ( .A(n53214), .B(n53215), .Z(n53137) );
  NAND U62818 ( .A(n53216), .B(n53217), .Z(n53215) );
  NAND U62819 ( .A(n53218), .B(n53219), .Z(n53214) );
  NANDN U62820 ( .A(n53220), .B(n53221), .Z(n53140) );
  ANDN U62821 ( .B(n53222), .A(n53223), .Z(n53134) );
  XNOR U62822 ( .A(n53125), .B(n53224), .Z(n53130) );
  XNOR U62823 ( .A(n53123), .B(n53127), .Z(n53224) );
  AND U62824 ( .A(n53225), .B(n53226), .Z(n53127) );
  NAND U62825 ( .A(n53227), .B(n53228), .Z(n53226) );
  NAND U62826 ( .A(n53229), .B(n53230), .Z(n53225) );
  AND U62827 ( .A(n53231), .B(n53232), .Z(n53123) );
  NAND U62828 ( .A(n53233), .B(n53234), .Z(n53232) );
  NAND U62829 ( .A(n53235), .B(n53236), .Z(n53231) );
  AND U62830 ( .A(n53237), .B(n53238), .Z(n53125) );
  XOR U62831 ( .A(n53205), .B(n53204), .Z(N60657) );
  XNOR U62832 ( .A(n53222), .B(n53223), .Z(n53204) );
  XNOR U62833 ( .A(n53237), .B(n53238), .Z(n53223) );
  XOR U62834 ( .A(n53234), .B(n53233), .Z(n53238) );
  XOR U62835 ( .A(y[132]), .B(x[132]), .Z(n53233) );
  XOR U62836 ( .A(n53236), .B(n53235), .Z(n53234) );
  XOR U62837 ( .A(y[134]), .B(x[134]), .Z(n53235) );
  XOR U62838 ( .A(y[133]), .B(x[133]), .Z(n53236) );
  XOR U62839 ( .A(n53228), .B(n53227), .Z(n53237) );
  XOR U62840 ( .A(n53230), .B(n53229), .Z(n53227) );
  XOR U62841 ( .A(y[131]), .B(x[131]), .Z(n53229) );
  XOR U62842 ( .A(y[130]), .B(x[130]), .Z(n53230) );
  XOR U62843 ( .A(y[129]), .B(x[129]), .Z(n53228) );
  XNOR U62844 ( .A(n53221), .B(n53220), .Z(n53222) );
  XNOR U62845 ( .A(n53217), .B(n53216), .Z(n53220) );
  XOR U62846 ( .A(n53219), .B(n53218), .Z(n53216) );
  XOR U62847 ( .A(y[128]), .B(x[128]), .Z(n53218) );
  XOR U62848 ( .A(y[127]), .B(x[127]), .Z(n53219) );
  XOR U62849 ( .A(y[126]), .B(x[126]), .Z(n53217) );
  XOR U62850 ( .A(n53211), .B(n53210), .Z(n53221) );
  XOR U62851 ( .A(n53213), .B(n53212), .Z(n53210) );
  XOR U62852 ( .A(y[125]), .B(x[125]), .Z(n53212) );
  XOR U62853 ( .A(y[124]), .B(x[124]), .Z(n53213) );
  XOR U62854 ( .A(y[123]), .B(x[123]), .Z(n53211) );
  XNOR U62855 ( .A(n53187), .B(n53188), .Z(n53205) );
  XNOR U62856 ( .A(n53202), .B(n53203), .Z(n53188) );
  XOR U62857 ( .A(n53199), .B(n53198), .Z(n53203) );
  XOR U62858 ( .A(y[120]), .B(x[120]), .Z(n53198) );
  XOR U62859 ( .A(n53201), .B(n53200), .Z(n53199) );
  XOR U62860 ( .A(y[122]), .B(x[122]), .Z(n53200) );
  XOR U62861 ( .A(y[121]), .B(x[121]), .Z(n53201) );
  XOR U62862 ( .A(n53193), .B(n53192), .Z(n53202) );
  XOR U62863 ( .A(n53195), .B(n53194), .Z(n53192) );
  XOR U62864 ( .A(y[119]), .B(x[119]), .Z(n53194) );
  XOR U62865 ( .A(y[118]), .B(x[118]), .Z(n53195) );
  XOR U62866 ( .A(y[117]), .B(x[117]), .Z(n53193) );
  XNOR U62867 ( .A(n53186), .B(n53185), .Z(n53187) );
  XNOR U62868 ( .A(n53182), .B(n53181), .Z(n53185) );
  XOR U62869 ( .A(n53184), .B(n53183), .Z(n53181) );
  XOR U62870 ( .A(y[116]), .B(x[116]), .Z(n53183) );
  XOR U62871 ( .A(y[115]), .B(x[115]), .Z(n53184) );
  XOR U62872 ( .A(y[114]), .B(x[114]), .Z(n53182) );
  XOR U62873 ( .A(n53176), .B(n53175), .Z(n53186) );
  XOR U62874 ( .A(n53178), .B(n53177), .Z(n53175) );
  XOR U62875 ( .A(y[113]), .B(x[113]), .Z(n53177) );
  XOR U62876 ( .A(y[112]), .B(x[112]), .Z(n53178) );
  XOR U62877 ( .A(y[111]), .B(x[111]), .Z(n53176) );
  NAND U62878 ( .A(n53239), .B(n53240), .Z(N60648) );
  NAND U62879 ( .A(n53241), .B(n53242), .Z(n53240) );
  NANDN U62880 ( .A(n53243), .B(n53244), .Z(n53242) );
  NANDN U62881 ( .A(n53244), .B(n53243), .Z(n53239) );
  XOR U62882 ( .A(n53243), .B(n53245), .Z(N60647) );
  XNOR U62883 ( .A(n53241), .B(n53244), .Z(n53245) );
  NAND U62884 ( .A(n53246), .B(n53247), .Z(n53244) );
  NAND U62885 ( .A(n53248), .B(n53249), .Z(n53247) );
  NANDN U62886 ( .A(n53250), .B(n53251), .Z(n53249) );
  NANDN U62887 ( .A(n53251), .B(n53250), .Z(n53246) );
  AND U62888 ( .A(n53252), .B(n53253), .Z(n53241) );
  NAND U62889 ( .A(n53254), .B(n53255), .Z(n53253) );
  NANDN U62890 ( .A(n53256), .B(n53257), .Z(n53255) );
  NANDN U62891 ( .A(n53257), .B(n53256), .Z(n53252) );
  IV U62892 ( .A(n53258), .Z(n53257) );
  AND U62893 ( .A(n53259), .B(n53260), .Z(n53243) );
  NAND U62894 ( .A(n53261), .B(n53262), .Z(n53260) );
  NANDN U62895 ( .A(n53263), .B(n53264), .Z(n53262) );
  NANDN U62896 ( .A(n53264), .B(n53263), .Z(n53259) );
  XOR U62897 ( .A(n53256), .B(n53265), .Z(N60646) );
  XNOR U62898 ( .A(n53254), .B(n53258), .Z(n53265) );
  XOR U62899 ( .A(n53251), .B(n53266), .Z(n53258) );
  XNOR U62900 ( .A(n53248), .B(n53250), .Z(n53266) );
  AND U62901 ( .A(n53267), .B(n53268), .Z(n53250) );
  NANDN U62902 ( .A(n53269), .B(n53270), .Z(n53268) );
  OR U62903 ( .A(n53271), .B(n53272), .Z(n53270) );
  IV U62904 ( .A(n53273), .Z(n53272) );
  NANDN U62905 ( .A(n53273), .B(n53271), .Z(n53267) );
  AND U62906 ( .A(n53274), .B(n53275), .Z(n53248) );
  NAND U62907 ( .A(n53276), .B(n53277), .Z(n53275) );
  NANDN U62908 ( .A(n53278), .B(n53279), .Z(n53277) );
  NANDN U62909 ( .A(n53279), .B(n53278), .Z(n53274) );
  IV U62910 ( .A(n53280), .Z(n53279) );
  NAND U62911 ( .A(n53281), .B(n53282), .Z(n53251) );
  NANDN U62912 ( .A(n53283), .B(n53284), .Z(n53282) );
  NANDN U62913 ( .A(n53285), .B(n53286), .Z(n53284) );
  NANDN U62914 ( .A(n53286), .B(n53285), .Z(n53281) );
  IV U62915 ( .A(n53287), .Z(n53285) );
  AND U62916 ( .A(n53288), .B(n53289), .Z(n53254) );
  NAND U62917 ( .A(n53290), .B(n53291), .Z(n53289) );
  NANDN U62918 ( .A(n53292), .B(n53293), .Z(n53291) );
  NANDN U62919 ( .A(n53293), .B(n53292), .Z(n53288) );
  XOR U62920 ( .A(n53264), .B(n53294), .Z(n53256) );
  XNOR U62921 ( .A(n53261), .B(n53263), .Z(n53294) );
  AND U62922 ( .A(n53295), .B(n53296), .Z(n53263) );
  NANDN U62923 ( .A(n53297), .B(n53298), .Z(n53296) );
  OR U62924 ( .A(n53299), .B(n53300), .Z(n53298) );
  IV U62925 ( .A(n53301), .Z(n53300) );
  NANDN U62926 ( .A(n53301), .B(n53299), .Z(n53295) );
  AND U62927 ( .A(n53302), .B(n53303), .Z(n53261) );
  NAND U62928 ( .A(n53304), .B(n53305), .Z(n53303) );
  NANDN U62929 ( .A(n53306), .B(n53307), .Z(n53305) );
  NANDN U62930 ( .A(n53307), .B(n53306), .Z(n53302) );
  IV U62931 ( .A(n53308), .Z(n53307) );
  NAND U62932 ( .A(n53309), .B(n53310), .Z(n53264) );
  NANDN U62933 ( .A(n53311), .B(n53312), .Z(n53310) );
  NANDN U62934 ( .A(n53313), .B(n53314), .Z(n53312) );
  NANDN U62935 ( .A(n53314), .B(n53313), .Z(n53309) );
  IV U62936 ( .A(n53315), .Z(n53313) );
  XOR U62937 ( .A(n53290), .B(n53316), .Z(N60645) );
  XNOR U62938 ( .A(n53293), .B(n53292), .Z(n53316) );
  XNOR U62939 ( .A(n53304), .B(n53317), .Z(n53292) );
  XNOR U62940 ( .A(n53308), .B(n53306), .Z(n53317) );
  XOR U62941 ( .A(n53314), .B(n53318), .Z(n53306) );
  XNOR U62942 ( .A(n53311), .B(n53315), .Z(n53318) );
  AND U62943 ( .A(n53319), .B(n53320), .Z(n53315) );
  NAND U62944 ( .A(n53321), .B(n53322), .Z(n53320) );
  NAND U62945 ( .A(n53323), .B(n53324), .Z(n53319) );
  AND U62946 ( .A(n53325), .B(n53326), .Z(n53311) );
  NAND U62947 ( .A(n53327), .B(n53328), .Z(n53326) );
  NAND U62948 ( .A(n53329), .B(n53330), .Z(n53325) );
  NANDN U62949 ( .A(n53331), .B(n53332), .Z(n53314) );
  ANDN U62950 ( .B(n53333), .A(n53334), .Z(n53308) );
  XNOR U62951 ( .A(n53299), .B(n53335), .Z(n53304) );
  XNOR U62952 ( .A(n53297), .B(n53301), .Z(n53335) );
  AND U62953 ( .A(n53336), .B(n53337), .Z(n53301) );
  NAND U62954 ( .A(n53338), .B(n53339), .Z(n53337) );
  NAND U62955 ( .A(n53340), .B(n53341), .Z(n53336) );
  AND U62956 ( .A(n53342), .B(n53343), .Z(n53297) );
  NAND U62957 ( .A(n53344), .B(n53345), .Z(n53343) );
  NAND U62958 ( .A(n53346), .B(n53347), .Z(n53342) );
  AND U62959 ( .A(n53348), .B(n53349), .Z(n53299) );
  NAND U62960 ( .A(n53350), .B(n53351), .Z(n53293) );
  XNOR U62961 ( .A(n53276), .B(n53352), .Z(n53290) );
  XNOR U62962 ( .A(n53280), .B(n53278), .Z(n53352) );
  XOR U62963 ( .A(n53286), .B(n53353), .Z(n53278) );
  XNOR U62964 ( .A(n53283), .B(n53287), .Z(n53353) );
  AND U62965 ( .A(n53354), .B(n53355), .Z(n53287) );
  NAND U62966 ( .A(n53356), .B(n53357), .Z(n53355) );
  NAND U62967 ( .A(n53358), .B(n53359), .Z(n53354) );
  AND U62968 ( .A(n53360), .B(n53361), .Z(n53283) );
  NAND U62969 ( .A(n53362), .B(n53363), .Z(n53361) );
  NAND U62970 ( .A(n53364), .B(n53365), .Z(n53360) );
  NANDN U62971 ( .A(n53366), .B(n53367), .Z(n53286) );
  ANDN U62972 ( .B(n53368), .A(n53369), .Z(n53280) );
  XNOR U62973 ( .A(n53271), .B(n53370), .Z(n53276) );
  XNOR U62974 ( .A(n53269), .B(n53273), .Z(n53370) );
  AND U62975 ( .A(n53371), .B(n53372), .Z(n53273) );
  NAND U62976 ( .A(n53373), .B(n53374), .Z(n53372) );
  NAND U62977 ( .A(n53375), .B(n53376), .Z(n53371) );
  AND U62978 ( .A(n53377), .B(n53378), .Z(n53269) );
  NAND U62979 ( .A(n53379), .B(n53380), .Z(n53378) );
  NAND U62980 ( .A(n53381), .B(n53382), .Z(n53377) );
  AND U62981 ( .A(n53383), .B(n53384), .Z(n53271) );
  XOR U62982 ( .A(n53351), .B(n53350), .Z(N60644) );
  XNOR U62983 ( .A(n53368), .B(n53369), .Z(n53350) );
  XNOR U62984 ( .A(n53383), .B(n53384), .Z(n53369) );
  XOR U62985 ( .A(n53380), .B(n53379), .Z(n53384) );
  XOR U62986 ( .A(y[108]), .B(x[108]), .Z(n53379) );
  XOR U62987 ( .A(n53382), .B(n53381), .Z(n53380) );
  XOR U62988 ( .A(y[110]), .B(x[110]), .Z(n53381) );
  XOR U62989 ( .A(y[109]), .B(x[109]), .Z(n53382) );
  XOR U62990 ( .A(n53374), .B(n53373), .Z(n53383) );
  XOR U62991 ( .A(n53376), .B(n53375), .Z(n53373) );
  XOR U62992 ( .A(y[107]), .B(x[107]), .Z(n53375) );
  XOR U62993 ( .A(y[106]), .B(x[106]), .Z(n53376) );
  XOR U62994 ( .A(y[105]), .B(x[105]), .Z(n53374) );
  XNOR U62995 ( .A(n53367), .B(n53366), .Z(n53368) );
  XNOR U62996 ( .A(n53363), .B(n53362), .Z(n53366) );
  XOR U62997 ( .A(n53365), .B(n53364), .Z(n53362) );
  XOR U62998 ( .A(y[104]), .B(x[104]), .Z(n53364) );
  XOR U62999 ( .A(y[103]), .B(x[103]), .Z(n53365) );
  XOR U63000 ( .A(y[102]), .B(x[102]), .Z(n53363) );
  XOR U63001 ( .A(n53357), .B(n53356), .Z(n53367) );
  XOR U63002 ( .A(n53359), .B(n53358), .Z(n53356) );
  XOR U63003 ( .A(y[101]), .B(x[101]), .Z(n53358) );
  XOR U63004 ( .A(y[100]), .B(x[100]), .Z(n53359) );
  XOR U63005 ( .A(y[99]), .B(x[99]), .Z(n53357) );
  XNOR U63006 ( .A(n53333), .B(n53334), .Z(n53351) );
  XNOR U63007 ( .A(n53348), .B(n53349), .Z(n53334) );
  XOR U63008 ( .A(n53345), .B(n53344), .Z(n53349) );
  XOR U63009 ( .A(y[96]), .B(x[96]), .Z(n53344) );
  XOR U63010 ( .A(n53347), .B(n53346), .Z(n53345) );
  XOR U63011 ( .A(y[98]), .B(x[98]), .Z(n53346) );
  XOR U63012 ( .A(y[97]), .B(x[97]), .Z(n53347) );
  XOR U63013 ( .A(n53339), .B(n53338), .Z(n53348) );
  XOR U63014 ( .A(n53341), .B(n53340), .Z(n53338) );
  XOR U63015 ( .A(y[95]), .B(x[95]), .Z(n53340) );
  XOR U63016 ( .A(y[94]), .B(x[94]), .Z(n53341) );
  XOR U63017 ( .A(y[93]), .B(x[93]), .Z(n53339) );
  XNOR U63018 ( .A(n53332), .B(n53331), .Z(n53333) );
  XNOR U63019 ( .A(n53328), .B(n53327), .Z(n53331) );
  XOR U63020 ( .A(n53330), .B(n53329), .Z(n53327) );
  XOR U63021 ( .A(y[92]), .B(x[92]), .Z(n53329) );
  XOR U63022 ( .A(y[91]), .B(x[91]), .Z(n53330) );
  XOR U63023 ( .A(y[90]), .B(x[90]), .Z(n53328) );
  XOR U63024 ( .A(n53322), .B(n53321), .Z(n53332) );
  XOR U63025 ( .A(n53324), .B(n53323), .Z(n53321) );
  XOR U63026 ( .A(y[89]), .B(x[89]), .Z(n53323) );
  XOR U63027 ( .A(y[88]), .B(x[88]), .Z(n53324) );
  XOR U63028 ( .A(y[87]), .B(x[87]), .Z(n53322) );
  NAND U63029 ( .A(n53385), .B(n53386), .Z(N60635) );
  NAND U63030 ( .A(n53387), .B(n53388), .Z(n53386) );
  NANDN U63031 ( .A(n53389), .B(n53390), .Z(n53388) );
  NANDN U63032 ( .A(n53390), .B(n53389), .Z(n53385) );
  XOR U63033 ( .A(n53389), .B(n53391), .Z(N60634) );
  XNOR U63034 ( .A(n53387), .B(n53390), .Z(n53391) );
  NAND U63035 ( .A(n53392), .B(n53393), .Z(n53390) );
  NAND U63036 ( .A(n53394), .B(n53395), .Z(n53393) );
  NANDN U63037 ( .A(n53396), .B(n53397), .Z(n53395) );
  NANDN U63038 ( .A(n53397), .B(n53396), .Z(n53392) );
  AND U63039 ( .A(n53398), .B(n53399), .Z(n53387) );
  NAND U63040 ( .A(n53400), .B(n53401), .Z(n53399) );
  NANDN U63041 ( .A(n53402), .B(n53403), .Z(n53401) );
  NANDN U63042 ( .A(n53403), .B(n53402), .Z(n53398) );
  IV U63043 ( .A(n53404), .Z(n53403) );
  AND U63044 ( .A(n53405), .B(n53406), .Z(n53389) );
  NAND U63045 ( .A(n53407), .B(n53408), .Z(n53406) );
  NANDN U63046 ( .A(n53409), .B(n53410), .Z(n53408) );
  NANDN U63047 ( .A(n53410), .B(n53409), .Z(n53405) );
  XOR U63048 ( .A(n53402), .B(n53411), .Z(N60633) );
  XNOR U63049 ( .A(n53400), .B(n53404), .Z(n53411) );
  XOR U63050 ( .A(n53397), .B(n53412), .Z(n53404) );
  XNOR U63051 ( .A(n53394), .B(n53396), .Z(n53412) );
  AND U63052 ( .A(n53413), .B(n53414), .Z(n53396) );
  NANDN U63053 ( .A(n53415), .B(n53416), .Z(n53414) );
  OR U63054 ( .A(n53417), .B(n53418), .Z(n53416) );
  IV U63055 ( .A(n53419), .Z(n53418) );
  NANDN U63056 ( .A(n53419), .B(n53417), .Z(n53413) );
  AND U63057 ( .A(n53420), .B(n53421), .Z(n53394) );
  NAND U63058 ( .A(n53422), .B(n53423), .Z(n53421) );
  NANDN U63059 ( .A(n53424), .B(n53425), .Z(n53423) );
  NANDN U63060 ( .A(n53425), .B(n53424), .Z(n53420) );
  IV U63061 ( .A(n53426), .Z(n53425) );
  NAND U63062 ( .A(n53427), .B(n53428), .Z(n53397) );
  NANDN U63063 ( .A(n53429), .B(n53430), .Z(n53428) );
  NANDN U63064 ( .A(n53431), .B(n53432), .Z(n53430) );
  NANDN U63065 ( .A(n53432), .B(n53431), .Z(n53427) );
  IV U63066 ( .A(n53433), .Z(n53431) );
  AND U63067 ( .A(n53434), .B(n53435), .Z(n53400) );
  NAND U63068 ( .A(n53436), .B(n53437), .Z(n53435) );
  NANDN U63069 ( .A(n53438), .B(n53439), .Z(n53437) );
  NANDN U63070 ( .A(n53439), .B(n53438), .Z(n53434) );
  XOR U63071 ( .A(n53410), .B(n53440), .Z(n53402) );
  XNOR U63072 ( .A(n53407), .B(n53409), .Z(n53440) );
  AND U63073 ( .A(n53441), .B(n53442), .Z(n53409) );
  NANDN U63074 ( .A(n53443), .B(n53444), .Z(n53442) );
  OR U63075 ( .A(n53445), .B(n53446), .Z(n53444) );
  IV U63076 ( .A(n53447), .Z(n53446) );
  NANDN U63077 ( .A(n53447), .B(n53445), .Z(n53441) );
  AND U63078 ( .A(n53448), .B(n53449), .Z(n53407) );
  NAND U63079 ( .A(n53450), .B(n53451), .Z(n53449) );
  NANDN U63080 ( .A(n53452), .B(n53453), .Z(n53451) );
  NANDN U63081 ( .A(n53453), .B(n53452), .Z(n53448) );
  IV U63082 ( .A(n53454), .Z(n53453) );
  NAND U63083 ( .A(n53455), .B(n53456), .Z(n53410) );
  NANDN U63084 ( .A(n53457), .B(n53458), .Z(n53456) );
  NANDN U63085 ( .A(n53459), .B(n53460), .Z(n53458) );
  NANDN U63086 ( .A(n53460), .B(n53459), .Z(n53455) );
  IV U63087 ( .A(n53461), .Z(n53459) );
  XOR U63088 ( .A(n53436), .B(n53462), .Z(N60632) );
  XNOR U63089 ( .A(n53439), .B(n53438), .Z(n53462) );
  XNOR U63090 ( .A(n53450), .B(n53463), .Z(n53438) );
  XNOR U63091 ( .A(n53454), .B(n53452), .Z(n53463) );
  XOR U63092 ( .A(n53460), .B(n53464), .Z(n53452) );
  XNOR U63093 ( .A(n53457), .B(n53461), .Z(n53464) );
  AND U63094 ( .A(n53465), .B(n53466), .Z(n53461) );
  NAND U63095 ( .A(n53467), .B(n53468), .Z(n53466) );
  NAND U63096 ( .A(n53469), .B(n53470), .Z(n53465) );
  AND U63097 ( .A(n53471), .B(n53472), .Z(n53457) );
  NAND U63098 ( .A(n53473), .B(n53474), .Z(n53472) );
  NAND U63099 ( .A(n53475), .B(n53476), .Z(n53471) );
  NANDN U63100 ( .A(n53477), .B(n53478), .Z(n53460) );
  ANDN U63101 ( .B(n53479), .A(n53480), .Z(n53454) );
  XNOR U63102 ( .A(n53445), .B(n53481), .Z(n53450) );
  XNOR U63103 ( .A(n53443), .B(n53447), .Z(n53481) );
  AND U63104 ( .A(n53482), .B(n53483), .Z(n53447) );
  NAND U63105 ( .A(n53484), .B(n53485), .Z(n53483) );
  NAND U63106 ( .A(n53486), .B(n53487), .Z(n53482) );
  AND U63107 ( .A(n53488), .B(n53489), .Z(n53443) );
  NAND U63108 ( .A(n53490), .B(n53491), .Z(n53489) );
  NAND U63109 ( .A(n53492), .B(n53493), .Z(n53488) );
  AND U63110 ( .A(n53494), .B(n53495), .Z(n53445) );
  NAND U63111 ( .A(n53496), .B(n53497), .Z(n53439) );
  XNOR U63112 ( .A(n53422), .B(n53498), .Z(n53436) );
  XNOR U63113 ( .A(n53426), .B(n53424), .Z(n53498) );
  XOR U63114 ( .A(n53432), .B(n53499), .Z(n53424) );
  XNOR U63115 ( .A(n53429), .B(n53433), .Z(n53499) );
  AND U63116 ( .A(n53500), .B(n53501), .Z(n53433) );
  NAND U63117 ( .A(n53502), .B(n53503), .Z(n53501) );
  NAND U63118 ( .A(n53504), .B(n53505), .Z(n53500) );
  AND U63119 ( .A(n53506), .B(n53507), .Z(n53429) );
  NAND U63120 ( .A(n53508), .B(n53509), .Z(n53507) );
  NAND U63121 ( .A(n53510), .B(n53511), .Z(n53506) );
  NANDN U63122 ( .A(n53512), .B(n53513), .Z(n53432) );
  ANDN U63123 ( .B(n53514), .A(n53515), .Z(n53426) );
  XNOR U63124 ( .A(n53417), .B(n53516), .Z(n53422) );
  XNOR U63125 ( .A(n53415), .B(n53419), .Z(n53516) );
  AND U63126 ( .A(n53517), .B(n53518), .Z(n53419) );
  NAND U63127 ( .A(n53519), .B(n53520), .Z(n53518) );
  NAND U63128 ( .A(n53521), .B(n53522), .Z(n53517) );
  AND U63129 ( .A(n53523), .B(n53524), .Z(n53415) );
  NAND U63130 ( .A(n53525), .B(n53526), .Z(n53524) );
  NAND U63131 ( .A(n53527), .B(n53528), .Z(n53523) );
  AND U63132 ( .A(n53529), .B(n53530), .Z(n53417) );
  XOR U63133 ( .A(n53497), .B(n53496), .Z(N60631) );
  XNOR U63134 ( .A(n53514), .B(n53515), .Z(n53496) );
  XNOR U63135 ( .A(n53529), .B(n53530), .Z(n53515) );
  XOR U63136 ( .A(n53526), .B(n53525), .Z(n53530) );
  XOR U63137 ( .A(y[84]), .B(x[84]), .Z(n53525) );
  XOR U63138 ( .A(n53528), .B(n53527), .Z(n53526) );
  XOR U63139 ( .A(y[86]), .B(x[86]), .Z(n53527) );
  XOR U63140 ( .A(y[85]), .B(x[85]), .Z(n53528) );
  XOR U63141 ( .A(n53520), .B(n53519), .Z(n53529) );
  XOR U63142 ( .A(n53522), .B(n53521), .Z(n53519) );
  XOR U63143 ( .A(y[83]), .B(x[83]), .Z(n53521) );
  XOR U63144 ( .A(y[82]), .B(x[82]), .Z(n53522) );
  XOR U63145 ( .A(y[81]), .B(x[81]), .Z(n53520) );
  XNOR U63146 ( .A(n53513), .B(n53512), .Z(n53514) );
  XNOR U63147 ( .A(n53509), .B(n53508), .Z(n53512) );
  XOR U63148 ( .A(n53511), .B(n53510), .Z(n53508) );
  XOR U63149 ( .A(y[80]), .B(x[80]), .Z(n53510) );
  XOR U63150 ( .A(y[79]), .B(x[79]), .Z(n53511) );
  XOR U63151 ( .A(y[78]), .B(x[78]), .Z(n53509) );
  XOR U63152 ( .A(n53503), .B(n53502), .Z(n53513) );
  XOR U63153 ( .A(n53505), .B(n53504), .Z(n53502) );
  XOR U63154 ( .A(y[77]), .B(x[77]), .Z(n53504) );
  XOR U63155 ( .A(y[76]), .B(x[76]), .Z(n53505) );
  XOR U63156 ( .A(y[75]), .B(x[75]), .Z(n53503) );
  XNOR U63157 ( .A(n53479), .B(n53480), .Z(n53497) );
  XNOR U63158 ( .A(n53494), .B(n53495), .Z(n53480) );
  XOR U63159 ( .A(n53491), .B(n53490), .Z(n53495) );
  XOR U63160 ( .A(y[72]), .B(x[72]), .Z(n53490) );
  XOR U63161 ( .A(n53493), .B(n53492), .Z(n53491) );
  XOR U63162 ( .A(y[74]), .B(x[74]), .Z(n53492) );
  XOR U63163 ( .A(y[73]), .B(x[73]), .Z(n53493) );
  XOR U63164 ( .A(n53485), .B(n53484), .Z(n53494) );
  XOR U63165 ( .A(n53487), .B(n53486), .Z(n53484) );
  XOR U63166 ( .A(y[71]), .B(x[71]), .Z(n53486) );
  XOR U63167 ( .A(y[70]), .B(x[70]), .Z(n53487) );
  XOR U63168 ( .A(y[69]), .B(x[69]), .Z(n53485) );
  XNOR U63169 ( .A(n53478), .B(n53477), .Z(n53479) );
  XNOR U63170 ( .A(n53474), .B(n53473), .Z(n53477) );
  XOR U63171 ( .A(n53476), .B(n53475), .Z(n53473) );
  XOR U63172 ( .A(y[68]), .B(x[68]), .Z(n53475) );
  XOR U63173 ( .A(y[67]), .B(x[67]), .Z(n53476) );
  XOR U63174 ( .A(y[66]), .B(x[66]), .Z(n53474) );
  XOR U63175 ( .A(n53468), .B(n53467), .Z(n53478) );
  XOR U63176 ( .A(n53470), .B(n53469), .Z(n53467) );
  XOR U63177 ( .A(y[65]), .B(x[65]), .Z(n53469) );
  XOR U63178 ( .A(y[64]), .B(x[64]), .Z(n53470) );
  XOR U63179 ( .A(y[63]), .B(x[63]), .Z(n53468) );
  NAND U63180 ( .A(n53531), .B(n53532), .Z(N60622) );
  NAND U63181 ( .A(n53533), .B(n53534), .Z(n53532) );
  NANDN U63182 ( .A(n53535), .B(n53536), .Z(n53534) );
  NANDN U63183 ( .A(n53536), .B(n53535), .Z(n53531) );
  XOR U63184 ( .A(n53535), .B(n53537), .Z(N60621) );
  XNOR U63185 ( .A(n53533), .B(n53536), .Z(n53537) );
  NAND U63186 ( .A(n53538), .B(n53539), .Z(n53536) );
  NAND U63187 ( .A(n53540), .B(n53541), .Z(n53539) );
  NANDN U63188 ( .A(n53542), .B(n53543), .Z(n53541) );
  NANDN U63189 ( .A(n53543), .B(n53542), .Z(n53538) );
  AND U63190 ( .A(n53544), .B(n53545), .Z(n53533) );
  NAND U63191 ( .A(n53546), .B(n53547), .Z(n53545) );
  NANDN U63192 ( .A(n53548), .B(n53549), .Z(n53547) );
  NANDN U63193 ( .A(n53549), .B(n53548), .Z(n53544) );
  IV U63194 ( .A(n53550), .Z(n53549) );
  AND U63195 ( .A(n53551), .B(n53552), .Z(n53535) );
  NAND U63196 ( .A(n53553), .B(n53554), .Z(n53552) );
  NANDN U63197 ( .A(n53555), .B(n53556), .Z(n53554) );
  NANDN U63198 ( .A(n53556), .B(n53555), .Z(n53551) );
  XOR U63199 ( .A(n53548), .B(n53557), .Z(N60620) );
  XNOR U63200 ( .A(n53546), .B(n53550), .Z(n53557) );
  XOR U63201 ( .A(n53543), .B(n53558), .Z(n53550) );
  XNOR U63202 ( .A(n53540), .B(n53542), .Z(n53558) );
  AND U63203 ( .A(n53559), .B(n53560), .Z(n53542) );
  NANDN U63204 ( .A(n53561), .B(n53562), .Z(n53560) );
  OR U63205 ( .A(n53563), .B(n53564), .Z(n53562) );
  IV U63206 ( .A(n53565), .Z(n53564) );
  NANDN U63207 ( .A(n53565), .B(n53563), .Z(n53559) );
  AND U63208 ( .A(n53566), .B(n53567), .Z(n53540) );
  NAND U63209 ( .A(n53568), .B(n53569), .Z(n53567) );
  NANDN U63210 ( .A(n53570), .B(n53571), .Z(n53569) );
  NANDN U63211 ( .A(n53571), .B(n53570), .Z(n53566) );
  IV U63212 ( .A(n53572), .Z(n53571) );
  NAND U63213 ( .A(n53573), .B(n53574), .Z(n53543) );
  NANDN U63214 ( .A(n53575), .B(n53576), .Z(n53574) );
  NANDN U63215 ( .A(n53577), .B(n53578), .Z(n53576) );
  NANDN U63216 ( .A(n53578), .B(n53577), .Z(n53573) );
  IV U63217 ( .A(n53579), .Z(n53577) );
  AND U63218 ( .A(n53580), .B(n53581), .Z(n53546) );
  NAND U63219 ( .A(n53582), .B(n53583), .Z(n53581) );
  NANDN U63220 ( .A(n53584), .B(n53585), .Z(n53583) );
  NANDN U63221 ( .A(n53585), .B(n53584), .Z(n53580) );
  XOR U63222 ( .A(n53556), .B(n53586), .Z(n53548) );
  XNOR U63223 ( .A(n53553), .B(n53555), .Z(n53586) );
  AND U63224 ( .A(n53587), .B(n53588), .Z(n53555) );
  NANDN U63225 ( .A(n53589), .B(n53590), .Z(n53588) );
  OR U63226 ( .A(n53591), .B(n53592), .Z(n53590) );
  IV U63227 ( .A(n53593), .Z(n53592) );
  NANDN U63228 ( .A(n53593), .B(n53591), .Z(n53587) );
  AND U63229 ( .A(n53594), .B(n53595), .Z(n53553) );
  NAND U63230 ( .A(n53596), .B(n53597), .Z(n53595) );
  NANDN U63231 ( .A(n53598), .B(n53599), .Z(n53597) );
  NANDN U63232 ( .A(n53599), .B(n53598), .Z(n53594) );
  IV U63233 ( .A(n53600), .Z(n53599) );
  NAND U63234 ( .A(n53601), .B(n53602), .Z(n53556) );
  NANDN U63235 ( .A(n53603), .B(n53604), .Z(n53602) );
  NANDN U63236 ( .A(n53605), .B(n53606), .Z(n53604) );
  NANDN U63237 ( .A(n53606), .B(n53605), .Z(n53601) );
  IV U63238 ( .A(n53607), .Z(n53605) );
  XOR U63239 ( .A(n53582), .B(n53608), .Z(N60619) );
  XNOR U63240 ( .A(n53585), .B(n53584), .Z(n53608) );
  XNOR U63241 ( .A(n53596), .B(n53609), .Z(n53584) );
  XNOR U63242 ( .A(n53600), .B(n53598), .Z(n53609) );
  XOR U63243 ( .A(n53606), .B(n53610), .Z(n53598) );
  XNOR U63244 ( .A(n53603), .B(n53607), .Z(n53610) );
  AND U63245 ( .A(n53611), .B(n53612), .Z(n53607) );
  NAND U63246 ( .A(n53613), .B(n53614), .Z(n53612) );
  NAND U63247 ( .A(n53615), .B(n53616), .Z(n53611) );
  AND U63248 ( .A(n53617), .B(n53618), .Z(n53603) );
  NAND U63249 ( .A(n53619), .B(n53620), .Z(n53618) );
  NAND U63250 ( .A(n53621), .B(n53622), .Z(n53617) );
  NANDN U63251 ( .A(n53623), .B(n53624), .Z(n53606) );
  ANDN U63252 ( .B(n53625), .A(n53626), .Z(n53600) );
  XNOR U63253 ( .A(n53591), .B(n53627), .Z(n53596) );
  XNOR U63254 ( .A(n53589), .B(n53593), .Z(n53627) );
  AND U63255 ( .A(n53628), .B(n53629), .Z(n53593) );
  NAND U63256 ( .A(n53630), .B(n53631), .Z(n53629) );
  NAND U63257 ( .A(n53632), .B(n53633), .Z(n53628) );
  AND U63258 ( .A(n53634), .B(n53635), .Z(n53589) );
  NAND U63259 ( .A(n53636), .B(n53637), .Z(n53635) );
  NAND U63260 ( .A(n53638), .B(n53639), .Z(n53634) );
  AND U63261 ( .A(n53640), .B(n53641), .Z(n53591) );
  NAND U63262 ( .A(n53642), .B(n53643), .Z(n53585) );
  XNOR U63263 ( .A(n53568), .B(n53644), .Z(n53582) );
  XNOR U63264 ( .A(n53572), .B(n53570), .Z(n53644) );
  XOR U63265 ( .A(n53578), .B(n53645), .Z(n53570) );
  XNOR U63266 ( .A(n53575), .B(n53579), .Z(n53645) );
  AND U63267 ( .A(n53646), .B(n53647), .Z(n53579) );
  NAND U63268 ( .A(n53648), .B(n53649), .Z(n53647) );
  NAND U63269 ( .A(n53650), .B(n53651), .Z(n53646) );
  AND U63270 ( .A(n53652), .B(n53653), .Z(n53575) );
  NAND U63271 ( .A(n53654), .B(n53655), .Z(n53653) );
  NAND U63272 ( .A(n53656), .B(n53657), .Z(n53652) );
  NANDN U63273 ( .A(n53658), .B(n53659), .Z(n53578) );
  ANDN U63274 ( .B(n53660), .A(n53661), .Z(n53572) );
  XNOR U63275 ( .A(n53563), .B(n53662), .Z(n53568) );
  XNOR U63276 ( .A(n53561), .B(n53565), .Z(n53662) );
  AND U63277 ( .A(n53663), .B(n53664), .Z(n53565) );
  NAND U63278 ( .A(n53665), .B(n53666), .Z(n53664) );
  NAND U63279 ( .A(n53667), .B(n53668), .Z(n53663) );
  AND U63280 ( .A(n53669), .B(n53670), .Z(n53561) );
  NAND U63281 ( .A(n53671), .B(n53672), .Z(n53670) );
  NAND U63282 ( .A(n53673), .B(n53674), .Z(n53669) );
  AND U63283 ( .A(n53675), .B(n53676), .Z(n53563) );
  XOR U63284 ( .A(n53643), .B(n53642), .Z(N60618) );
  XNOR U63285 ( .A(n53660), .B(n53661), .Z(n53642) );
  XNOR U63286 ( .A(n53675), .B(n53676), .Z(n53661) );
  XOR U63287 ( .A(n53672), .B(n53671), .Z(n53676) );
  XOR U63288 ( .A(y[60]), .B(x[60]), .Z(n53671) );
  XOR U63289 ( .A(n53674), .B(n53673), .Z(n53672) );
  XOR U63290 ( .A(y[62]), .B(x[62]), .Z(n53673) );
  XOR U63291 ( .A(y[61]), .B(x[61]), .Z(n53674) );
  XOR U63292 ( .A(n53666), .B(n53665), .Z(n53675) );
  XOR U63293 ( .A(n53668), .B(n53667), .Z(n53665) );
  XOR U63294 ( .A(y[59]), .B(x[59]), .Z(n53667) );
  XOR U63295 ( .A(y[58]), .B(x[58]), .Z(n53668) );
  XOR U63296 ( .A(y[57]), .B(x[57]), .Z(n53666) );
  XNOR U63297 ( .A(n53659), .B(n53658), .Z(n53660) );
  XNOR U63298 ( .A(n53655), .B(n53654), .Z(n53658) );
  XOR U63299 ( .A(n53657), .B(n53656), .Z(n53654) );
  XOR U63300 ( .A(y[56]), .B(x[56]), .Z(n53656) );
  XOR U63301 ( .A(y[55]), .B(x[55]), .Z(n53657) );
  XOR U63302 ( .A(y[54]), .B(x[54]), .Z(n53655) );
  XOR U63303 ( .A(n53649), .B(n53648), .Z(n53659) );
  XOR U63304 ( .A(n53651), .B(n53650), .Z(n53648) );
  XOR U63305 ( .A(y[53]), .B(x[53]), .Z(n53650) );
  XOR U63306 ( .A(y[52]), .B(x[52]), .Z(n53651) );
  XOR U63307 ( .A(y[51]), .B(x[51]), .Z(n53649) );
  XNOR U63308 ( .A(n53625), .B(n53626), .Z(n53643) );
  XNOR U63309 ( .A(n53640), .B(n53641), .Z(n53626) );
  XOR U63310 ( .A(n53637), .B(n53636), .Z(n53641) );
  XOR U63311 ( .A(y[48]), .B(x[48]), .Z(n53636) );
  XOR U63312 ( .A(n53639), .B(n53638), .Z(n53637) );
  XOR U63313 ( .A(y[50]), .B(x[50]), .Z(n53638) );
  XOR U63314 ( .A(y[49]), .B(x[49]), .Z(n53639) );
  XOR U63315 ( .A(n53631), .B(n53630), .Z(n53640) );
  XOR U63316 ( .A(n53633), .B(n53632), .Z(n53630) );
  XOR U63317 ( .A(y[47]), .B(x[47]), .Z(n53632) );
  XOR U63318 ( .A(y[46]), .B(x[46]), .Z(n53633) );
  XOR U63319 ( .A(y[45]), .B(x[45]), .Z(n53631) );
  XNOR U63320 ( .A(n53624), .B(n53623), .Z(n53625) );
  XNOR U63321 ( .A(n53620), .B(n53619), .Z(n53623) );
  XOR U63322 ( .A(n53622), .B(n53621), .Z(n53619) );
  XOR U63323 ( .A(y[44]), .B(x[44]), .Z(n53621) );
  XOR U63324 ( .A(y[43]), .B(x[43]), .Z(n53622) );
  XOR U63325 ( .A(y[42]), .B(x[42]), .Z(n53620) );
  XOR U63326 ( .A(n53614), .B(n53613), .Z(n53624) );
  XOR U63327 ( .A(n53616), .B(n53615), .Z(n53613) );
  XOR U63328 ( .A(y[41]), .B(x[41]), .Z(n53615) );
  XOR U63329 ( .A(y[40]), .B(x[40]), .Z(n53616) );
  XOR U63330 ( .A(y[39]), .B(x[39]), .Z(n53614) );
  NAND U63331 ( .A(n53677), .B(n53678), .Z(N60609) );
  NAND U63332 ( .A(n53679), .B(n53680), .Z(n53678) );
  NANDN U63333 ( .A(n53681), .B(n53682), .Z(n53680) );
  NANDN U63334 ( .A(n53682), .B(n53681), .Z(n53677) );
  XOR U63335 ( .A(n53681), .B(n53683), .Z(N60608) );
  XNOR U63336 ( .A(n53679), .B(n53682), .Z(n53683) );
  NAND U63337 ( .A(n53684), .B(n53685), .Z(n53682) );
  NAND U63338 ( .A(n53686), .B(n53687), .Z(n53685) );
  NANDN U63339 ( .A(n53688), .B(n53689), .Z(n53687) );
  NANDN U63340 ( .A(n53689), .B(n53688), .Z(n53684) );
  AND U63341 ( .A(n53690), .B(n53691), .Z(n53679) );
  NAND U63342 ( .A(n53692), .B(n53693), .Z(n53691) );
  NANDN U63343 ( .A(n53694), .B(n53695), .Z(n53693) );
  NANDN U63344 ( .A(n53695), .B(n53694), .Z(n53690) );
  IV U63345 ( .A(n53696), .Z(n53695) );
  AND U63346 ( .A(n53697), .B(n53698), .Z(n53681) );
  NAND U63347 ( .A(n53699), .B(n53700), .Z(n53698) );
  NANDN U63348 ( .A(n53701), .B(n53702), .Z(n53700) );
  NANDN U63349 ( .A(n53702), .B(n53701), .Z(n53697) );
  XOR U63350 ( .A(n53694), .B(n53703), .Z(N60607) );
  XNOR U63351 ( .A(n53692), .B(n53696), .Z(n53703) );
  XOR U63352 ( .A(n53689), .B(n53704), .Z(n53696) );
  XNOR U63353 ( .A(n53686), .B(n53688), .Z(n53704) );
  AND U63354 ( .A(n53705), .B(n53706), .Z(n53688) );
  NANDN U63355 ( .A(n53707), .B(n53708), .Z(n53706) );
  OR U63356 ( .A(n53709), .B(n53710), .Z(n53708) );
  IV U63357 ( .A(n53711), .Z(n53710) );
  NANDN U63358 ( .A(n53711), .B(n53709), .Z(n53705) );
  AND U63359 ( .A(n53712), .B(n53713), .Z(n53686) );
  NAND U63360 ( .A(n53714), .B(n53715), .Z(n53713) );
  NANDN U63361 ( .A(n53716), .B(n53717), .Z(n53715) );
  NANDN U63362 ( .A(n53717), .B(n53716), .Z(n53712) );
  IV U63363 ( .A(n53718), .Z(n53717) );
  NAND U63364 ( .A(n53719), .B(n53720), .Z(n53689) );
  NANDN U63365 ( .A(n53721), .B(n53722), .Z(n53720) );
  NANDN U63366 ( .A(n53723), .B(n53724), .Z(n53722) );
  NANDN U63367 ( .A(n53724), .B(n53723), .Z(n53719) );
  IV U63368 ( .A(n53725), .Z(n53723) );
  AND U63369 ( .A(n53726), .B(n53727), .Z(n53692) );
  NAND U63370 ( .A(n53728), .B(n53729), .Z(n53727) );
  NANDN U63371 ( .A(n53730), .B(n53731), .Z(n53729) );
  NANDN U63372 ( .A(n53731), .B(n53730), .Z(n53726) );
  XOR U63373 ( .A(n53702), .B(n53732), .Z(n53694) );
  XNOR U63374 ( .A(n53699), .B(n53701), .Z(n53732) );
  AND U63375 ( .A(n53733), .B(n53734), .Z(n53701) );
  NANDN U63376 ( .A(n53735), .B(n53736), .Z(n53734) );
  OR U63377 ( .A(n53737), .B(n53738), .Z(n53736) );
  IV U63378 ( .A(n53739), .Z(n53738) );
  NANDN U63379 ( .A(n53739), .B(n53737), .Z(n53733) );
  AND U63380 ( .A(n53740), .B(n53741), .Z(n53699) );
  NAND U63381 ( .A(n53742), .B(n53743), .Z(n53741) );
  NANDN U63382 ( .A(n53744), .B(n53745), .Z(n53743) );
  NANDN U63383 ( .A(n53745), .B(n53744), .Z(n53740) );
  IV U63384 ( .A(n53746), .Z(n53745) );
  NAND U63385 ( .A(n53747), .B(n53748), .Z(n53702) );
  NANDN U63386 ( .A(n53749), .B(n53750), .Z(n53748) );
  NANDN U63387 ( .A(n53751), .B(n53752), .Z(n53750) );
  NANDN U63388 ( .A(n53752), .B(n53751), .Z(n53747) );
  IV U63389 ( .A(n53753), .Z(n53751) );
  XOR U63390 ( .A(n53728), .B(n53754), .Z(N60606) );
  XNOR U63391 ( .A(n53731), .B(n53730), .Z(n53754) );
  XNOR U63392 ( .A(n53742), .B(n53755), .Z(n53730) );
  XNOR U63393 ( .A(n53746), .B(n53744), .Z(n53755) );
  XOR U63394 ( .A(n53752), .B(n53756), .Z(n53744) );
  XNOR U63395 ( .A(n53749), .B(n53753), .Z(n53756) );
  AND U63396 ( .A(n53757), .B(n53758), .Z(n53753) );
  NAND U63397 ( .A(n53759), .B(n53760), .Z(n53758) );
  NAND U63398 ( .A(n53761), .B(n53762), .Z(n53757) );
  AND U63399 ( .A(n53763), .B(n53764), .Z(n53749) );
  NAND U63400 ( .A(n53765), .B(n53766), .Z(n53764) );
  NAND U63401 ( .A(n53767), .B(n53768), .Z(n53763) );
  NANDN U63402 ( .A(n53769), .B(n53770), .Z(n53752) );
  ANDN U63403 ( .B(n53771), .A(n53772), .Z(n53746) );
  XNOR U63404 ( .A(n53737), .B(n53773), .Z(n53742) );
  XNOR U63405 ( .A(n53735), .B(n53739), .Z(n53773) );
  AND U63406 ( .A(n53774), .B(n53775), .Z(n53739) );
  NAND U63407 ( .A(n53776), .B(n53777), .Z(n53775) );
  NAND U63408 ( .A(n53778), .B(n53779), .Z(n53774) );
  AND U63409 ( .A(n53780), .B(n53781), .Z(n53735) );
  NAND U63410 ( .A(n53782), .B(n53783), .Z(n53781) );
  NAND U63411 ( .A(n53784), .B(n53785), .Z(n53780) );
  AND U63412 ( .A(n53786), .B(n53787), .Z(n53737) );
  NAND U63413 ( .A(n53788), .B(n53789), .Z(n53731) );
  XNOR U63414 ( .A(n53714), .B(n53790), .Z(n53728) );
  XNOR U63415 ( .A(n53718), .B(n53716), .Z(n53790) );
  XOR U63416 ( .A(n53724), .B(n53791), .Z(n53716) );
  XNOR U63417 ( .A(n53721), .B(n53725), .Z(n53791) );
  AND U63418 ( .A(n53792), .B(n53793), .Z(n53725) );
  NAND U63419 ( .A(n53794), .B(n53795), .Z(n53793) );
  NAND U63420 ( .A(n53796), .B(n53797), .Z(n53792) );
  AND U63421 ( .A(n53798), .B(n53799), .Z(n53721) );
  NAND U63422 ( .A(n53800), .B(n53801), .Z(n53799) );
  NAND U63423 ( .A(n53802), .B(n53803), .Z(n53798) );
  NANDN U63424 ( .A(n53804), .B(n53805), .Z(n53724) );
  ANDN U63425 ( .B(n53806), .A(n53807), .Z(n53718) );
  XNOR U63426 ( .A(n53709), .B(n53808), .Z(n53714) );
  XNOR U63427 ( .A(n53707), .B(n53711), .Z(n53808) );
  AND U63428 ( .A(n53809), .B(n53810), .Z(n53711) );
  NAND U63429 ( .A(n53811), .B(n53812), .Z(n53810) );
  NAND U63430 ( .A(n53813), .B(n53814), .Z(n53809) );
  AND U63431 ( .A(n53815), .B(n53816), .Z(n53707) );
  NAND U63432 ( .A(n53817), .B(n53818), .Z(n53816) );
  NAND U63433 ( .A(n53819), .B(n53820), .Z(n53815) );
  AND U63434 ( .A(n53821), .B(n53822), .Z(n53709) );
  XOR U63435 ( .A(n53789), .B(n53788), .Z(N60605) );
  XNOR U63436 ( .A(n53806), .B(n53807), .Z(n53788) );
  XNOR U63437 ( .A(n53821), .B(n53822), .Z(n53807) );
  XOR U63438 ( .A(n53818), .B(n53817), .Z(n53822) );
  XOR U63439 ( .A(y[36]), .B(x[36]), .Z(n53817) );
  XOR U63440 ( .A(n53820), .B(n53819), .Z(n53818) );
  XOR U63441 ( .A(y[38]), .B(x[38]), .Z(n53819) );
  XOR U63442 ( .A(y[37]), .B(x[37]), .Z(n53820) );
  XOR U63443 ( .A(n53812), .B(n53811), .Z(n53821) );
  XOR U63444 ( .A(n53814), .B(n53813), .Z(n53811) );
  XOR U63445 ( .A(y[35]), .B(x[35]), .Z(n53813) );
  XOR U63446 ( .A(y[34]), .B(x[34]), .Z(n53814) );
  XOR U63447 ( .A(y[33]), .B(x[33]), .Z(n53812) );
  XNOR U63448 ( .A(n53805), .B(n53804), .Z(n53806) );
  XNOR U63449 ( .A(n53801), .B(n53800), .Z(n53804) );
  XOR U63450 ( .A(n53803), .B(n53802), .Z(n53800) );
  XOR U63451 ( .A(y[32]), .B(x[32]), .Z(n53802) );
  XOR U63452 ( .A(y[31]), .B(x[31]), .Z(n53803) );
  XOR U63453 ( .A(y[30]), .B(x[30]), .Z(n53801) );
  XOR U63454 ( .A(n53795), .B(n53794), .Z(n53805) );
  XOR U63455 ( .A(n53797), .B(n53796), .Z(n53794) );
  XOR U63456 ( .A(y[29]), .B(x[29]), .Z(n53796) );
  XOR U63457 ( .A(y[28]), .B(x[28]), .Z(n53797) );
  XOR U63458 ( .A(y[27]), .B(x[27]), .Z(n53795) );
  XNOR U63459 ( .A(n53771), .B(n53772), .Z(n53789) );
  XNOR U63460 ( .A(n53786), .B(n53787), .Z(n53772) );
  XOR U63461 ( .A(n53783), .B(n53782), .Z(n53787) );
  XOR U63462 ( .A(y[24]), .B(x[24]), .Z(n53782) );
  XOR U63463 ( .A(n53785), .B(n53784), .Z(n53783) );
  XOR U63464 ( .A(y[26]), .B(x[26]), .Z(n53784) );
  XOR U63465 ( .A(y[25]), .B(x[25]), .Z(n53785) );
  XOR U63466 ( .A(n53777), .B(n53776), .Z(n53786) );
  XOR U63467 ( .A(n53779), .B(n53778), .Z(n53776) );
  XOR U63468 ( .A(y[23]), .B(x[23]), .Z(n53778) );
  XOR U63469 ( .A(y[22]), .B(x[22]), .Z(n53779) );
  XOR U63470 ( .A(y[21]), .B(x[21]), .Z(n53777) );
  XNOR U63471 ( .A(n53770), .B(n53769), .Z(n53771) );
  XNOR U63472 ( .A(n53766), .B(n53765), .Z(n53769) );
  XOR U63473 ( .A(n53768), .B(n53767), .Z(n53765) );
  XOR U63474 ( .A(y[20]), .B(x[20]), .Z(n53767) );
  XOR U63475 ( .A(y[19]), .B(x[19]), .Z(n53768) );
  XOR U63476 ( .A(y[18]), .B(x[18]), .Z(n53766) );
  XOR U63477 ( .A(n53760), .B(n53759), .Z(n53770) );
  XOR U63478 ( .A(n53762), .B(n53761), .Z(n53759) );
  XOR U63479 ( .A(y[17]), .B(x[17]), .Z(n53761) );
  XOR U63480 ( .A(y[16]), .B(x[16]), .Z(n53762) );
  XOR U63481 ( .A(y[15]), .B(x[15]), .Z(n53760) );
  NAND U63482 ( .A(n53823), .B(n53824), .Z(N60596) );
  NAND U63483 ( .A(n53825), .B(n53826), .Z(n53824) );
  NAND U63484 ( .A(n53827), .B(n53826), .Z(n53823) );
  XOR U63485 ( .A(n53827), .B(n53828), .Z(N60595) );
  XOR U63486 ( .A(n53825), .B(n53826), .Z(n53828) );
  AND U63487 ( .A(n53829), .B(n53830), .Z(n53826) );
  NAND U63488 ( .A(n53831), .B(n53832), .Z(n53830) );
  NANDN U63489 ( .A(n53833), .B(n53834), .Z(n53832) );
  NANDN U63490 ( .A(n53834), .B(n53833), .Z(n53829) );
  AND U63491 ( .A(n53835), .B(n53836), .Z(n53825) );
  NAND U63492 ( .A(n53837), .B(n53838), .Z(n53836) );
  NANDN U63493 ( .A(n53839), .B(n53840), .Z(n53838) );
  NANDN U63494 ( .A(n53840), .B(n53839), .Z(n53835) );
  IV U63495 ( .A(n53841), .Z(n53840) );
  ANDN U63496 ( .B(n53842), .A(n53843), .Z(n53827) );
  XOR U63497 ( .A(n53839), .B(n53844), .Z(N60594) );
  XNOR U63498 ( .A(n53837), .B(n53841), .Z(n53844) );
  XOR U63499 ( .A(n53834), .B(n53845), .Z(n53841) );
  XNOR U63500 ( .A(n53831), .B(n53833), .Z(n53845) );
  AND U63501 ( .A(n53846), .B(n53847), .Z(n53833) );
  NANDN U63502 ( .A(n53848), .B(n53849), .Z(n53847) );
  OR U63503 ( .A(n53850), .B(n53851), .Z(n53849) );
  IV U63504 ( .A(n53852), .Z(n53851) );
  NANDN U63505 ( .A(n53852), .B(n53850), .Z(n53846) );
  AND U63506 ( .A(n53853), .B(n53854), .Z(n53831) );
  NAND U63507 ( .A(n53855), .B(n53856), .Z(n53854) );
  NANDN U63508 ( .A(n53857), .B(n53858), .Z(n53856) );
  NANDN U63509 ( .A(n53858), .B(n53857), .Z(n53853) );
  IV U63510 ( .A(n53859), .Z(n53858) );
  NAND U63511 ( .A(n53860), .B(n53861), .Z(n53834) );
  NANDN U63512 ( .A(n53862), .B(n53863), .Z(n53861) );
  IV U63513 ( .A(n53864), .Z(n53862) );
  NANDN U63514 ( .A(n53865), .B(n53866), .Z(n53860) );
  AND U63515 ( .A(n53867), .B(n53868), .Z(n53837) );
  NAND U63516 ( .A(n53869), .B(n53870), .Z(n53868) );
  NANDN U63517 ( .A(n53871), .B(n53872), .Z(n53870) );
  NANDN U63518 ( .A(n53872), .B(n53871), .Z(n53867) );
  XOR U63519 ( .A(n53843), .B(n53842), .Z(n53839) );
  ANDN U63520 ( .B(n53873), .A(n53874), .Z(n53842) );
  AND U63521 ( .A(n53875), .B(n53876), .Z(n53843) );
  NAND U63522 ( .A(n53877), .B(n53878), .Z(n53876) );
  NANDN U63523 ( .A(n53879), .B(n53880), .Z(n53878) );
  NANDN U63524 ( .A(n53880), .B(n53879), .Z(n53875) );
  XOR U63525 ( .A(n53869), .B(n53881), .Z(N60593) );
  XNOR U63526 ( .A(n53872), .B(n53871), .Z(n53881) );
  XOR U63527 ( .A(n53877), .B(n53882), .Z(n53871) );
  XNOR U63528 ( .A(n53880), .B(n53879), .Z(n53882) );
  ANDN U63529 ( .B(n53883), .A(n53884), .Z(n53879) );
  AND U63530 ( .A(n53885), .B(n53886), .Z(n53880) );
  NAND U63531 ( .A(n53887), .B(n53888), .Z(n53886) );
  NAND U63532 ( .A(n53889), .B(n53890), .Z(n53885) );
  XNOR U63533 ( .A(n53874), .B(n53873), .Z(n53877) );
  NAND U63534 ( .A(n53891), .B(n53892), .Z(n53873) );
  NAND U63535 ( .A(n53893), .B(n53894), .Z(n53892) );
  NANDN U63536 ( .A(n53895), .B(n53896), .Z(n53891) );
  AND U63537 ( .A(n53897), .B(n53898), .Z(n53874) );
  NAND U63538 ( .A(n53899), .B(n53900), .Z(n53898) );
  NANDN U63539 ( .A(n53901), .B(n53902), .Z(n53897) );
  NAND U63540 ( .A(n53903), .B(n53904), .Z(n53872) );
  XNOR U63541 ( .A(n53855), .B(n53905), .Z(n53869) );
  XNOR U63542 ( .A(n53859), .B(n53857), .Z(n53905) );
  XOR U63543 ( .A(n53863), .B(n53864), .Z(n53857) );
  XNOR U63544 ( .A(n53865), .B(n53866), .Z(n53864) );
  NAND U63545 ( .A(n53906), .B(n53907), .Z(n53866) );
  NAND U63546 ( .A(n53908), .B(n53909), .Z(n53907) );
  NANDN U63547 ( .A(n53910), .B(n53911), .Z(n53906) );
  AND U63548 ( .A(n53912), .B(n53913), .Z(n53865) );
  NANDN U63549 ( .A(n53914), .B(n53915), .Z(n53913) );
  NAND U63550 ( .A(n53916), .B(n53917), .Z(n53912) );
  ANDN U63551 ( .B(n53918), .A(n53919), .Z(n53863) );
  ANDN U63552 ( .B(n53920), .A(n53921), .Z(n53859) );
  XNOR U63553 ( .A(n53850), .B(n53922), .Z(n53855) );
  XNOR U63554 ( .A(n53848), .B(n53852), .Z(n53922) );
  AND U63555 ( .A(n53923), .B(n53924), .Z(n53852) );
  NAND U63556 ( .A(n53925), .B(n53926), .Z(n53924) );
  NAND U63557 ( .A(n53927), .B(n53928), .Z(n53923) );
  AND U63558 ( .A(n53929), .B(n53930), .Z(n53848) );
  NAND U63559 ( .A(n53931), .B(n53932), .Z(n53930) );
  NAND U63560 ( .A(n53933), .B(n53934), .Z(n53929) );
  AND U63561 ( .A(n53935), .B(n53936), .Z(n53850) );
  XOR U63562 ( .A(n53904), .B(n53903), .Z(N60592) );
  XNOR U63563 ( .A(n53920), .B(n53921), .Z(n53903) );
  XNOR U63564 ( .A(n53935), .B(n53936), .Z(n53921) );
  XOR U63565 ( .A(n53932), .B(n53931), .Z(n53936) );
  XOR U63566 ( .A(y[12]), .B(x[12]), .Z(n53931) );
  XOR U63567 ( .A(n53934), .B(n53933), .Z(n53932) );
  XOR U63568 ( .A(y[14]), .B(x[14]), .Z(n53933) );
  XOR U63569 ( .A(y[13]), .B(x[13]), .Z(n53934) );
  XOR U63570 ( .A(n53926), .B(n53925), .Z(n53935) );
  XOR U63571 ( .A(n53928), .B(n53927), .Z(n53925) );
  XOR U63572 ( .A(y[11]), .B(x[11]), .Z(n53927) );
  XOR U63573 ( .A(y[10]), .B(x[10]), .Z(n53928) );
  XOR U63574 ( .A(y[9]), .B(x[9]), .Z(n53926) );
  XNOR U63575 ( .A(n53918), .B(n53919), .Z(n53920) );
  XNOR U63576 ( .A(n53909), .B(n53908), .Z(n53919) );
  XNOR U63577 ( .A(n53911), .B(n53910), .Z(n53908) );
  XNOR U63578 ( .A(y[5]), .B(x[5]), .Z(n53910) );
  XOR U63579 ( .A(y[4]), .B(x[4]), .Z(n53911) );
  XOR U63580 ( .A(y[3]), .B(x[3]), .Z(n53909) );
  XNOR U63581 ( .A(n53915), .B(n53914), .Z(n53918) );
  XNOR U63582 ( .A(n53917), .B(n53916), .Z(n53914) );
  XOR U63583 ( .A(y[8]), .B(x[8]), .Z(n53916) );
  XOR U63584 ( .A(y[7]), .B(x[7]), .Z(n53917) );
  XOR U63585 ( .A(y[6]), .B(x[6]), .Z(n53915) );
  XNOR U63586 ( .A(n53883), .B(n53884), .Z(n53904) );
  XNOR U63587 ( .A(n53894), .B(n53893), .Z(n53884) );
  XNOR U63588 ( .A(n53896), .B(n53895), .Z(n53893) );
  XNOR U63589 ( .A(n53900), .B(n53899), .Z(n53895) );
  XOR U63590 ( .A(y[0]), .B(x[0]), .Z(n53899) );
  XNOR U63591 ( .A(n53902), .B(n53901), .Z(n53900) );
  XNOR U63592 ( .A(y[2]), .B(x[2]), .Z(n53901) );
  XOR U63593 ( .A(y[1]), .B(x[1]), .Z(n53902) );
  XOR U63594 ( .A(y[7999]), .B(x[7999]), .Z(n53896) );
  XOR U63595 ( .A(y[7998]), .B(x[7998]), .Z(n53894) );
  XOR U63596 ( .A(n53888), .B(n53887), .Z(n53883) );
  XOR U63597 ( .A(n53890), .B(n53889), .Z(n53887) );
  XOR U63598 ( .A(y[7997]), .B(x[7997]), .Z(n53889) );
  XOR U63599 ( .A(y[7996]), .B(x[7996]), .Z(n53890) );
  XOR U63600 ( .A(y[7995]), .B(x[7995]), .Z(n53888) );
  NAND U63601 ( .A(n53937), .B(n53938), .Z(N60582) );
  NANDN U63602 ( .A(n53939), .B(n53940), .Z(n53938) );
  NANDN U63603 ( .A(n53941), .B(n53942), .Z(n53940) );
  NANDN U63604 ( .A(n53942), .B(n53941), .Z(n53937) );
  IV U63605 ( .A(n53943), .Z(n53941) );
  XOR U63606 ( .A(n53942), .B(n53944), .Z(N60581) );
  XNOR U63607 ( .A(n53939), .B(n53943), .Z(n53944) );
  AND U63608 ( .A(n53945), .B(n53946), .Z(n53943) );
  NANDN U63609 ( .A(n53947), .B(n53948), .Z(n53946) );
  NANDN U63610 ( .A(n53949), .B(n53950), .Z(n53948) );
  NANDN U63611 ( .A(n53950), .B(n53949), .Z(n53945) );
  IV U63612 ( .A(n53951), .Z(n53949) );
  IV U63613 ( .A(n53952), .Z(n53950) );
  AND U63614 ( .A(n53953), .B(n53954), .Z(n53939) );
  NAND U63615 ( .A(n53955), .B(n53956), .Z(n53954) );
  NANDN U63616 ( .A(n53957), .B(n53958), .Z(n53956) );
  NANDN U63617 ( .A(n53958), .B(n53957), .Z(n53953) );
  AND U63618 ( .A(n53959), .B(n53960), .Z(n53942) );
  NANDN U63619 ( .A(n53961), .B(n53962), .Z(n53960) );
  NANDN U63620 ( .A(n53963), .B(n53964), .Z(n53962) );
  NANDN U63621 ( .A(n53964), .B(n53963), .Z(n53959) );
  IV U63622 ( .A(n53965), .Z(n53963) );
  XOR U63623 ( .A(n53955), .B(n53966), .Z(N60580) );
  XNOR U63624 ( .A(n53958), .B(n53957), .Z(n53966) );
  XOR U63625 ( .A(n53964), .B(n53967), .Z(n53957) );
  XNOR U63626 ( .A(n53961), .B(n53965), .Z(n53967) );
  AND U63627 ( .A(n53968), .B(n53969), .Z(n53965) );
  NAND U63628 ( .A(n53970), .B(n53971), .Z(n53969) );
  NAND U63629 ( .A(n53972), .B(n53973), .Z(n53968) );
  AND U63630 ( .A(n53974), .B(n53975), .Z(n53961) );
  NAND U63631 ( .A(n53976), .B(n53977), .Z(n53975) );
  NAND U63632 ( .A(n53978), .B(n53979), .Z(n53974) );
  NANDN U63633 ( .A(n53980), .B(n53981), .Z(n53964) );
  NAND U63634 ( .A(n53982), .B(n53983), .Z(n53958) );
  XNOR U63635 ( .A(n53952), .B(n53984), .Z(n53955) );
  XNOR U63636 ( .A(n53947), .B(n53951), .Z(n53984) );
  AND U63637 ( .A(n53985), .B(n53986), .Z(n53951) );
  NAND U63638 ( .A(n53987), .B(n53988), .Z(n53986) );
  NAND U63639 ( .A(n53989), .B(n53990), .Z(n53985) );
  AND U63640 ( .A(n53991), .B(n53992), .Z(n53947) );
  NAND U63641 ( .A(n53993), .B(n53994), .Z(n53992) );
  NAND U63642 ( .A(n53995), .B(n53996), .Z(n53991) );
  ANDN U63643 ( .B(n53997), .A(n53998), .Z(n53952) );
  XOR U63644 ( .A(n53983), .B(n53982), .Z(N60579) );
  XNOR U63645 ( .A(n53997), .B(n53998), .Z(n53982) );
  XNOR U63646 ( .A(n53994), .B(n53993), .Z(n53998) );
  XOR U63647 ( .A(y[7992]), .B(x[7992]), .Z(n53993) );
  XOR U63648 ( .A(n53996), .B(n53995), .Z(n53994) );
  XOR U63649 ( .A(y[7994]), .B(x[7994]), .Z(n53995) );
  XOR U63650 ( .A(y[7993]), .B(x[7993]), .Z(n53996) );
  XOR U63651 ( .A(n53988), .B(n53987), .Z(n53997) );
  XOR U63652 ( .A(y[7989]), .B(x[7989]), .Z(n53987) );
  XOR U63653 ( .A(n53990), .B(n53989), .Z(n53988) );
  XOR U63654 ( .A(y[7991]), .B(x[7991]), .Z(n53989) );
  XOR U63655 ( .A(y[7990]), .B(x[7990]), .Z(n53990) );
  XNOR U63656 ( .A(n53981), .B(n53980), .Z(n53983) );
  XNOR U63657 ( .A(n53977), .B(n53976), .Z(n53980) );
  XOR U63658 ( .A(n53979), .B(n53978), .Z(n53976) );
  XOR U63659 ( .A(y[7988]), .B(x[7988]), .Z(n53978) );
  XOR U63660 ( .A(y[7987]), .B(x[7987]), .Z(n53979) );
  XOR U63661 ( .A(y[7986]), .B(x[7986]), .Z(n53977) );
  XOR U63662 ( .A(n53971), .B(n53970), .Z(n53981) );
  XOR U63663 ( .A(n53973), .B(n53972), .Z(n53970) );
  XOR U63664 ( .A(y[7985]), .B(x[7985]), .Z(n53972) );
  XOR U63665 ( .A(y[7984]), .B(x[7984]), .Z(n53973) );
  XOR U63666 ( .A(y[7983]), .B(x[7983]), .Z(n53971) );
endmodule

