
module compare_N16384_CC64 ( clk, rst, x, y, g );
  input [255:0] x;
  input [255:0] y;
  input clk, rst;
  output g;
  wire   ci, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280;

  DFF ci_reg ( .D(g), .CLK(clk), .RST(rst), .I(1'b1), .Q(ci) );
  XOR U260 ( .A(y[3]), .B(n1267), .Z(n1268) );
  XOR U261 ( .A(y[7]), .B(n1251), .Z(n1252) );
  XOR U262 ( .A(y[11]), .B(n1235), .Z(n1236) );
  XOR U263 ( .A(y[15]), .B(n1219), .Z(n1220) );
  XOR U264 ( .A(y[19]), .B(n1203), .Z(n1204) );
  XOR U265 ( .A(y[23]), .B(n1187), .Z(n1188) );
  XOR U266 ( .A(y[27]), .B(n1171), .Z(n1172) );
  XOR U267 ( .A(y[31]), .B(n1155), .Z(n1156) );
  XOR U268 ( .A(y[35]), .B(n1139), .Z(n1140) );
  XOR U269 ( .A(y[39]), .B(n1123), .Z(n1124) );
  XOR U270 ( .A(y[43]), .B(n1107), .Z(n1108) );
  XOR U271 ( .A(y[47]), .B(n1091), .Z(n1092) );
  XOR U272 ( .A(y[51]), .B(n1075), .Z(n1076) );
  XOR U273 ( .A(y[55]), .B(n1059), .Z(n1060) );
  XOR U274 ( .A(y[59]), .B(n1043), .Z(n1044) );
  XOR U275 ( .A(y[63]), .B(n1027), .Z(n1028) );
  XOR U276 ( .A(y[67]), .B(n1011), .Z(n1012) );
  XOR U277 ( .A(y[71]), .B(n995), .Z(n996) );
  XOR U278 ( .A(y[75]), .B(n979), .Z(n980) );
  XOR U279 ( .A(y[79]), .B(n963), .Z(n964) );
  XOR U280 ( .A(y[83]), .B(n947), .Z(n948) );
  XOR U281 ( .A(y[87]), .B(n931), .Z(n932) );
  XOR U282 ( .A(y[91]), .B(n915), .Z(n916) );
  XOR U283 ( .A(y[95]), .B(n899), .Z(n900) );
  XOR U284 ( .A(y[99]), .B(n883), .Z(n884) );
  XOR U285 ( .A(y[103]), .B(n867), .Z(n868) );
  XOR U286 ( .A(y[107]), .B(n851), .Z(n852) );
  XOR U287 ( .A(y[111]), .B(n835), .Z(n836) );
  XOR U288 ( .A(y[115]), .B(n819), .Z(n820) );
  XOR U289 ( .A(y[119]), .B(n803), .Z(n804) );
  XOR U290 ( .A(y[123]), .B(n787), .Z(n788) );
  XOR U291 ( .A(y[127]), .B(n771), .Z(n772) );
  XOR U292 ( .A(y[131]), .B(n755), .Z(n756) );
  XOR U293 ( .A(y[135]), .B(n739), .Z(n740) );
  XOR U294 ( .A(y[139]), .B(n723), .Z(n724) );
  XOR U295 ( .A(y[143]), .B(n707), .Z(n708) );
  XOR U296 ( .A(y[147]), .B(n691), .Z(n692) );
  XOR U297 ( .A(y[151]), .B(n675), .Z(n676) );
  XOR U298 ( .A(y[155]), .B(n659), .Z(n660) );
  XOR U299 ( .A(y[159]), .B(n643), .Z(n644) );
  XOR U300 ( .A(y[163]), .B(n627), .Z(n628) );
  XOR U301 ( .A(y[167]), .B(n611), .Z(n612) );
  XOR U302 ( .A(y[171]), .B(n595), .Z(n596) );
  XOR U303 ( .A(y[175]), .B(n579), .Z(n580) );
  XOR U304 ( .A(y[179]), .B(n563), .Z(n564) );
  XOR U305 ( .A(y[183]), .B(n547), .Z(n548) );
  XOR U306 ( .A(y[187]), .B(n531), .Z(n532) );
  XOR U307 ( .A(y[191]), .B(n515), .Z(n516) );
  XOR U308 ( .A(y[195]), .B(n499), .Z(n500) );
  XOR U309 ( .A(y[199]), .B(n483), .Z(n484) );
  XOR U310 ( .A(y[203]), .B(n467), .Z(n468) );
  XOR U311 ( .A(y[207]), .B(n451), .Z(n452) );
  XOR U312 ( .A(y[211]), .B(n435), .Z(n436) );
  XOR U313 ( .A(y[215]), .B(n419), .Z(n420) );
  XOR U314 ( .A(y[219]), .B(n403), .Z(n404) );
  XOR U315 ( .A(y[223]), .B(n387), .Z(n388) );
  XOR U316 ( .A(y[227]), .B(n371), .Z(n372) );
  XOR U317 ( .A(y[231]), .B(n355), .Z(n356) );
  XOR U318 ( .A(y[235]), .B(n339), .Z(n340) );
  XOR U319 ( .A(y[239]), .B(n323), .Z(n324) );
  XOR U320 ( .A(y[243]), .B(n307), .Z(n308) );
  XOR U321 ( .A(y[247]), .B(n291), .Z(n292) );
  XOR U322 ( .A(y[251]), .B(n275), .Z(n276) );
  XOR U323 ( .A(y[4]), .B(n1263), .Z(n1264) );
  XOR U324 ( .A(y[8]), .B(n1247), .Z(n1248) );
  XOR U325 ( .A(y[12]), .B(n1231), .Z(n1232) );
  XOR U326 ( .A(y[16]), .B(n1215), .Z(n1216) );
  XOR U327 ( .A(y[20]), .B(n1199), .Z(n1200) );
  XOR U328 ( .A(y[24]), .B(n1183), .Z(n1184) );
  XOR U329 ( .A(y[28]), .B(n1167), .Z(n1168) );
  XOR U330 ( .A(y[32]), .B(n1151), .Z(n1152) );
  XOR U331 ( .A(y[36]), .B(n1135), .Z(n1136) );
  XOR U332 ( .A(y[40]), .B(n1119), .Z(n1120) );
  XOR U333 ( .A(y[44]), .B(n1103), .Z(n1104) );
  XOR U334 ( .A(y[48]), .B(n1087), .Z(n1088) );
  XOR U335 ( .A(y[52]), .B(n1071), .Z(n1072) );
  XOR U336 ( .A(y[56]), .B(n1055), .Z(n1056) );
  XOR U337 ( .A(y[60]), .B(n1039), .Z(n1040) );
  XOR U338 ( .A(y[64]), .B(n1023), .Z(n1024) );
  XOR U339 ( .A(y[68]), .B(n1007), .Z(n1008) );
  XOR U340 ( .A(y[72]), .B(n991), .Z(n992) );
  XOR U341 ( .A(y[76]), .B(n975), .Z(n976) );
  XOR U342 ( .A(y[80]), .B(n959), .Z(n960) );
  XOR U343 ( .A(y[84]), .B(n943), .Z(n944) );
  XOR U344 ( .A(y[88]), .B(n927), .Z(n928) );
  XOR U345 ( .A(y[92]), .B(n911), .Z(n912) );
  XOR U346 ( .A(y[96]), .B(n895), .Z(n896) );
  XOR U347 ( .A(y[100]), .B(n879), .Z(n880) );
  XOR U348 ( .A(y[104]), .B(n863), .Z(n864) );
  XOR U349 ( .A(y[108]), .B(n847), .Z(n848) );
  XOR U350 ( .A(y[112]), .B(n831), .Z(n832) );
  XOR U351 ( .A(y[116]), .B(n815), .Z(n816) );
  XOR U352 ( .A(y[120]), .B(n799), .Z(n800) );
  XOR U353 ( .A(y[124]), .B(n783), .Z(n784) );
  XOR U354 ( .A(y[128]), .B(n767), .Z(n768) );
  XOR U355 ( .A(y[132]), .B(n751), .Z(n752) );
  XOR U356 ( .A(y[136]), .B(n735), .Z(n736) );
  XOR U357 ( .A(y[140]), .B(n719), .Z(n720) );
  XOR U358 ( .A(y[144]), .B(n703), .Z(n704) );
  XOR U359 ( .A(y[148]), .B(n687), .Z(n688) );
  XOR U360 ( .A(y[152]), .B(n671), .Z(n672) );
  XOR U361 ( .A(y[156]), .B(n655), .Z(n656) );
  XOR U362 ( .A(y[160]), .B(n639), .Z(n640) );
  XOR U363 ( .A(y[164]), .B(n623), .Z(n624) );
  XOR U364 ( .A(y[168]), .B(n607), .Z(n608) );
  XOR U365 ( .A(y[172]), .B(n591), .Z(n592) );
  XOR U366 ( .A(y[176]), .B(n575), .Z(n576) );
  XOR U367 ( .A(y[180]), .B(n559), .Z(n560) );
  XOR U368 ( .A(y[184]), .B(n543), .Z(n544) );
  XOR U369 ( .A(y[188]), .B(n527), .Z(n528) );
  XOR U370 ( .A(y[192]), .B(n511), .Z(n512) );
  XOR U371 ( .A(y[196]), .B(n495), .Z(n496) );
  XOR U372 ( .A(y[200]), .B(n479), .Z(n480) );
  XOR U373 ( .A(y[204]), .B(n463), .Z(n464) );
  XOR U374 ( .A(y[208]), .B(n447), .Z(n448) );
  XOR U375 ( .A(y[212]), .B(n431), .Z(n432) );
  XOR U376 ( .A(y[216]), .B(n415), .Z(n416) );
  XOR U377 ( .A(y[220]), .B(n399), .Z(n400) );
  XOR U378 ( .A(y[224]), .B(n383), .Z(n384) );
  XOR U379 ( .A(y[228]), .B(n367), .Z(n368) );
  XOR U380 ( .A(y[232]), .B(n351), .Z(n352) );
  XOR U381 ( .A(y[236]), .B(n335), .Z(n336) );
  XOR U382 ( .A(y[240]), .B(n319), .Z(n320) );
  XOR U383 ( .A(y[244]), .B(n303), .Z(n304) );
  XOR U384 ( .A(y[248]), .B(n287), .Z(n288) );
  XOR U385 ( .A(y[252]), .B(n271), .Z(n272) );
  XOR U386 ( .A(y[5]), .B(n1259), .Z(n1260) );
  XOR U387 ( .A(y[9]), .B(n1243), .Z(n1244) );
  XOR U388 ( .A(y[13]), .B(n1227), .Z(n1228) );
  XOR U389 ( .A(y[17]), .B(n1211), .Z(n1212) );
  XOR U390 ( .A(y[21]), .B(n1195), .Z(n1196) );
  XOR U391 ( .A(y[25]), .B(n1179), .Z(n1180) );
  XOR U392 ( .A(y[29]), .B(n1163), .Z(n1164) );
  XOR U393 ( .A(y[33]), .B(n1147), .Z(n1148) );
  XOR U394 ( .A(y[37]), .B(n1131), .Z(n1132) );
  XOR U395 ( .A(y[41]), .B(n1115), .Z(n1116) );
  XOR U396 ( .A(y[45]), .B(n1099), .Z(n1100) );
  XOR U397 ( .A(y[49]), .B(n1083), .Z(n1084) );
  XOR U398 ( .A(y[53]), .B(n1067), .Z(n1068) );
  XOR U399 ( .A(y[57]), .B(n1051), .Z(n1052) );
  XOR U400 ( .A(y[61]), .B(n1035), .Z(n1036) );
  XOR U401 ( .A(y[65]), .B(n1019), .Z(n1020) );
  XOR U402 ( .A(y[69]), .B(n1003), .Z(n1004) );
  XOR U403 ( .A(y[73]), .B(n987), .Z(n988) );
  XOR U404 ( .A(y[77]), .B(n971), .Z(n972) );
  XOR U405 ( .A(y[81]), .B(n955), .Z(n956) );
  XOR U406 ( .A(y[85]), .B(n939), .Z(n940) );
  XOR U407 ( .A(y[89]), .B(n923), .Z(n924) );
  XOR U408 ( .A(y[93]), .B(n907), .Z(n908) );
  XOR U409 ( .A(y[97]), .B(n891), .Z(n892) );
  XOR U410 ( .A(y[101]), .B(n875), .Z(n876) );
  XOR U411 ( .A(y[105]), .B(n859), .Z(n860) );
  XOR U412 ( .A(y[109]), .B(n843), .Z(n844) );
  XOR U413 ( .A(y[113]), .B(n827), .Z(n828) );
  XOR U414 ( .A(y[117]), .B(n811), .Z(n812) );
  XOR U415 ( .A(y[121]), .B(n795), .Z(n796) );
  XOR U416 ( .A(y[125]), .B(n779), .Z(n780) );
  XOR U417 ( .A(y[129]), .B(n763), .Z(n764) );
  XOR U418 ( .A(y[133]), .B(n747), .Z(n748) );
  XOR U419 ( .A(y[137]), .B(n731), .Z(n732) );
  XOR U420 ( .A(y[141]), .B(n715), .Z(n716) );
  XOR U421 ( .A(y[145]), .B(n699), .Z(n700) );
  XOR U422 ( .A(y[149]), .B(n683), .Z(n684) );
  XOR U423 ( .A(y[153]), .B(n667), .Z(n668) );
  XOR U424 ( .A(y[157]), .B(n651), .Z(n652) );
  XOR U425 ( .A(y[161]), .B(n635), .Z(n636) );
  XOR U426 ( .A(y[165]), .B(n619), .Z(n620) );
  XOR U427 ( .A(y[169]), .B(n603), .Z(n604) );
  XOR U428 ( .A(y[173]), .B(n587), .Z(n588) );
  XOR U429 ( .A(y[177]), .B(n571), .Z(n572) );
  XOR U430 ( .A(y[181]), .B(n555), .Z(n556) );
  XOR U431 ( .A(y[185]), .B(n539), .Z(n540) );
  XOR U432 ( .A(y[189]), .B(n523), .Z(n524) );
  XOR U433 ( .A(y[193]), .B(n507), .Z(n508) );
  XOR U434 ( .A(y[197]), .B(n491), .Z(n492) );
  XOR U435 ( .A(y[201]), .B(n475), .Z(n476) );
  XOR U436 ( .A(y[205]), .B(n459), .Z(n460) );
  XOR U437 ( .A(y[209]), .B(n443), .Z(n444) );
  XOR U438 ( .A(y[213]), .B(n427), .Z(n428) );
  XOR U439 ( .A(y[217]), .B(n411), .Z(n412) );
  XOR U440 ( .A(y[221]), .B(n395), .Z(n396) );
  XOR U441 ( .A(y[225]), .B(n379), .Z(n380) );
  XOR U442 ( .A(y[229]), .B(n363), .Z(n364) );
  XOR U443 ( .A(y[233]), .B(n347), .Z(n348) );
  XOR U444 ( .A(y[237]), .B(n331), .Z(n332) );
  XOR U445 ( .A(y[241]), .B(n315), .Z(n316) );
  XOR U446 ( .A(y[245]), .B(n299), .Z(n300) );
  XOR U447 ( .A(y[249]), .B(n283), .Z(n284) );
  XOR U448 ( .A(y[253]), .B(n267), .Z(n268) );
  XOR U449 ( .A(y[2]), .B(n1271), .Z(n1272) );
  XOR U450 ( .A(y[6]), .B(n1255), .Z(n1256) );
  XOR U451 ( .A(y[10]), .B(n1239), .Z(n1240) );
  XOR U452 ( .A(y[14]), .B(n1223), .Z(n1224) );
  XOR U453 ( .A(y[18]), .B(n1207), .Z(n1208) );
  XOR U454 ( .A(y[22]), .B(n1191), .Z(n1192) );
  XOR U455 ( .A(y[26]), .B(n1175), .Z(n1176) );
  XOR U456 ( .A(y[30]), .B(n1159), .Z(n1160) );
  XOR U457 ( .A(y[34]), .B(n1143), .Z(n1144) );
  XOR U458 ( .A(y[38]), .B(n1127), .Z(n1128) );
  XOR U459 ( .A(y[42]), .B(n1111), .Z(n1112) );
  XOR U460 ( .A(y[46]), .B(n1095), .Z(n1096) );
  XOR U461 ( .A(y[50]), .B(n1079), .Z(n1080) );
  XOR U462 ( .A(y[54]), .B(n1063), .Z(n1064) );
  XOR U463 ( .A(y[58]), .B(n1047), .Z(n1048) );
  XOR U464 ( .A(y[62]), .B(n1031), .Z(n1032) );
  XOR U465 ( .A(y[66]), .B(n1015), .Z(n1016) );
  XOR U466 ( .A(y[70]), .B(n999), .Z(n1000) );
  XOR U467 ( .A(y[74]), .B(n983), .Z(n984) );
  XOR U468 ( .A(y[78]), .B(n967), .Z(n968) );
  XOR U469 ( .A(y[82]), .B(n951), .Z(n952) );
  XOR U470 ( .A(y[86]), .B(n935), .Z(n936) );
  XOR U471 ( .A(y[90]), .B(n919), .Z(n920) );
  XOR U472 ( .A(y[94]), .B(n903), .Z(n904) );
  XOR U473 ( .A(y[98]), .B(n887), .Z(n888) );
  XOR U474 ( .A(y[102]), .B(n871), .Z(n872) );
  XOR U475 ( .A(y[106]), .B(n855), .Z(n856) );
  XOR U476 ( .A(y[110]), .B(n839), .Z(n840) );
  XOR U477 ( .A(y[114]), .B(n823), .Z(n824) );
  XOR U478 ( .A(y[118]), .B(n807), .Z(n808) );
  XOR U479 ( .A(y[122]), .B(n791), .Z(n792) );
  XOR U480 ( .A(y[126]), .B(n775), .Z(n776) );
  XOR U481 ( .A(y[130]), .B(n759), .Z(n760) );
  XOR U482 ( .A(y[134]), .B(n743), .Z(n744) );
  XOR U483 ( .A(y[138]), .B(n727), .Z(n728) );
  XOR U484 ( .A(y[142]), .B(n711), .Z(n712) );
  XOR U485 ( .A(y[146]), .B(n695), .Z(n696) );
  XOR U486 ( .A(y[150]), .B(n679), .Z(n680) );
  XOR U487 ( .A(y[154]), .B(n663), .Z(n664) );
  XOR U488 ( .A(y[158]), .B(n647), .Z(n648) );
  XOR U489 ( .A(y[162]), .B(n631), .Z(n632) );
  XOR U490 ( .A(y[166]), .B(n615), .Z(n616) );
  XOR U491 ( .A(y[170]), .B(n599), .Z(n600) );
  XOR U492 ( .A(y[174]), .B(n583), .Z(n584) );
  XOR U493 ( .A(y[178]), .B(n567), .Z(n568) );
  XOR U494 ( .A(y[182]), .B(n551), .Z(n552) );
  XOR U495 ( .A(y[186]), .B(n535), .Z(n536) );
  XOR U496 ( .A(y[190]), .B(n519), .Z(n520) );
  XOR U497 ( .A(y[194]), .B(n503), .Z(n504) );
  XOR U498 ( .A(y[198]), .B(n487), .Z(n488) );
  XOR U499 ( .A(y[202]), .B(n471), .Z(n472) );
  XOR U500 ( .A(y[206]), .B(n455), .Z(n456) );
  XOR U501 ( .A(y[210]), .B(n439), .Z(n440) );
  XOR U502 ( .A(y[214]), .B(n423), .Z(n424) );
  XOR U503 ( .A(y[218]), .B(n407), .Z(n408) );
  XOR U504 ( .A(y[222]), .B(n391), .Z(n392) );
  XOR U505 ( .A(y[226]), .B(n375), .Z(n376) );
  XOR U506 ( .A(y[230]), .B(n359), .Z(n360) );
  XOR U507 ( .A(y[234]), .B(n343), .Z(n344) );
  XOR U508 ( .A(y[238]), .B(n327), .Z(n328) );
  XOR U509 ( .A(y[242]), .B(n311), .Z(n312) );
  XOR U510 ( .A(y[246]), .B(n295), .Z(n296) );
  XOR U511 ( .A(y[250]), .B(n279), .Z(n280) );
  XOR U512 ( .A(y[254]), .B(n263), .Z(n264) );
  XOR U513 ( .A(n258), .B(n259), .Z(g) );
  AND U514 ( .A(n260), .B(n261), .Z(n258) );
  XOR U515 ( .A(x[255]), .B(n259), .Z(n261) );
  XNOR U516 ( .A(y[255]), .B(n259), .Z(n260) );
  XNOR U517 ( .A(n262), .B(n263), .Z(n259) );
  AND U518 ( .A(n264), .B(n265), .Z(n262) );
  XNOR U519 ( .A(x[254]), .B(n263), .Z(n265) );
  XOR U520 ( .A(n266), .B(n267), .Z(n263) );
  AND U521 ( .A(n268), .B(n269), .Z(n266) );
  XNOR U522 ( .A(x[253]), .B(n267), .Z(n269) );
  XOR U523 ( .A(n270), .B(n271), .Z(n267) );
  AND U524 ( .A(n272), .B(n273), .Z(n270) );
  XNOR U525 ( .A(x[252]), .B(n271), .Z(n273) );
  XOR U526 ( .A(n274), .B(n275), .Z(n271) );
  AND U527 ( .A(n276), .B(n277), .Z(n274) );
  XNOR U528 ( .A(x[251]), .B(n275), .Z(n277) );
  XOR U529 ( .A(n278), .B(n279), .Z(n275) );
  AND U530 ( .A(n280), .B(n281), .Z(n278) );
  XNOR U531 ( .A(x[250]), .B(n279), .Z(n281) );
  XOR U532 ( .A(n282), .B(n283), .Z(n279) );
  AND U533 ( .A(n284), .B(n285), .Z(n282) );
  XNOR U534 ( .A(x[249]), .B(n283), .Z(n285) );
  XOR U535 ( .A(n286), .B(n287), .Z(n283) );
  AND U536 ( .A(n288), .B(n289), .Z(n286) );
  XNOR U537 ( .A(x[248]), .B(n287), .Z(n289) );
  XOR U538 ( .A(n290), .B(n291), .Z(n287) );
  AND U539 ( .A(n292), .B(n293), .Z(n290) );
  XNOR U540 ( .A(x[247]), .B(n291), .Z(n293) );
  XOR U541 ( .A(n294), .B(n295), .Z(n291) );
  AND U542 ( .A(n296), .B(n297), .Z(n294) );
  XNOR U543 ( .A(x[246]), .B(n295), .Z(n297) );
  XOR U544 ( .A(n298), .B(n299), .Z(n295) );
  AND U545 ( .A(n300), .B(n301), .Z(n298) );
  XNOR U546 ( .A(x[245]), .B(n299), .Z(n301) );
  XOR U547 ( .A(n302), .B(n303), .Z(n299) );
  AND U548 ( .A(n304), .B(n305), .Z(n302) );
  XNOR U549 ( .A(x[244]), .B(n303), .Z(n305) );
  XOR U550 ( .A(n306), .B(n307), .Z(n303) );
  AND U551 ( .A(n308), .B(n309), .Z(n306) );
  XNOR U552 ( .A(x[243]), .B(n307), .Z(n309) );
  XOR U553 ( .A(n310), .B(n311), .Z(n307) );
  AND U554 ( .A(n312), .B(n313), .Z(n310) );
  XNOR U555 ( .A(x[242]), .B(n311), .Z(n313) );
  XOR U556 ( .A(n314), .B(n315), .Z(n311) );
  AND U557 ( .A(n316), .B(n317), .Z(n314) );
  XNOR U558 ( .A(x[241]), .B(n315), .Z(n317) );
  XOR U559 ( .A(n318), .B(n319), .Z(n315) );
  AND U560 ( .A(n320), .B(n321), .Z(n318) );
  XNOR U561 ( .A(x[240]), .B(n319), .Z(n321) );
  XOR U562 ( .A(n322), .B(n323), .Z(n319) );
  AND U563 ( .A(n324), .B(n325), .Z(n322) );
  XNOR U564 ( .A(x[239]), .B(n323), .Z(n325) );
  XOR U565 ( .A(n326), .B(n327), .Z(n323) );
  AND U566 ( .A(n328), .B(n329), .Z(n326) );
  XNOR U567 ( .A(x[238]), .B(n327), .Z(n329) );
  XOR U568 ( .A(n330), .B(n331), .Z(n327) );
  AND U569 ( .A(n332), .B(n333), .Z(n330) );
  XNOR U570 ( .A(x[237]), .B(n331), .Z(n333) );
  XOR U571 ( .A(n334), .B(n335), .Z(n331) );
  AND U572 ( .A(n336), .B(n337), .Z(n334) );
  XNOR U573 ( .A(x[236]), .B(n335), .Z(n337) );
  XOR U574 ( .A(n338), .B(n339), .Z(n335) );
  AND U575 ( .A(n340), .B(n341), .Z(n338) );
  XNOR U576 ( .A(x[235]), .B(n339), .Z(n341) );
  XOR U577 ( .A(n342), .B(n343), .Z(n339) );
  AND U578 ( .A(n344), .B(n345), .Z(n342) );
  XNOR U579 ( .A(x[234]), .B(n343), .Z(n345) );
  XOR U580 ( .A(n346), .B(n347), .Z(n343) );
  AND U581 ( .A(n348), .B(n349), .Z(n346) );
  XNOR U582 ( .A(x[233]), .B(n347), .Z(n349) );
  XOR U583 ( .A(n350), .B(n351), .Z(n347) );
  AND U584 ( .A(n352), .B(n353), .Z(n350) );
  XNOR U585 ( .A(x[232]), .B(n351), .Z(n353) );
  XOR U586 ( .A(n354), .B(n355), .Z(n351) );
  AND U587 ( .A(n356), .B(n357), .Z(n354) );
  XNOR U588 ( .A(x[231]), .B(n355), .Z(n357) );
  XOR U589 ( .A(n358), .B(n359), .Z(n355) );
  AND U590 ( .A(n360), .B(n361), .Z(n358) );
  XNOR U591 ( .A(x[230]), .B(n359), .Z(n361) );
  XOR U592 ( .A(n362), .B(n363), .Z(n359) );
  AND U593 ( .A(n364), .B(n365), .Z(n362) );
  XNOR U594 ( .A(x[229]), .B(n363), .Z(n365) );
  XOR U595 ( .A(n366), .B(n367), .Z(n363) );
  AND U596 ( .A(n368), .B(n369), .Z(n366) );
  XNOR U597 ( .A(x[228]), .B(n367), .Z(n369) );
  XOR U598 ( .A(n370), .B(n371), .Z(n367) );
  AND U599 ( .A(n372), .B(n373), .Z(n370) );
  XNOR U600 ( .A(x[227]), .B(n371), .Z(n373) );
  XOR U601 ( .A(n374), .B(n375), .Z(n371) );
  AND U602 ( .A(n376), .B(n377), .Z(n374) );
  XNOR U603 ( .A(x[226]), .B(n375), .Z(n377) );
  XOR U604 ( .A(n378), .B(n379), .Z(n375) );
  AND U605 ( .A(n380), .B(n381), .Z(n378) );
  XNOR U606 ( .A(x[225]), .B(n379), .Z(n381) );
  XOR U607 ( .A(n382), .B(n383), .Z(n379) );
  AND U608 ( .A(n384), .B(n385), .Z(n382) );
  XNOR U609 ( .A(x[224]), .B(n383), .Z(n385) );
  XOR U610 ( .A(n386), .B(n387), .Z(n383) );
  AND U611 ( .A(n388), .B(n389), .Z(n386) );
  XNOR U612 ( .A(x[223]), .B(n387), .Z(n389) );
  XOR U613 ( .A(n390), .B(n391), .Z(n387) );
  AND U614 ( .A(n392), .B(n393), .Z(n390) );
  XNOR U615 ( .A(x[222]), .B(n391), .Z(n393) );
  XOR U616 ( .A(n394), .B(n395), .Z(n391) );
  AND U617 ( .A(n396), .B(n397), .Z(n394) );
  XNOR U618 ( .A(x[221]), .B(n395), .Z(n397) );
  XOR U619 ( .A(n398), .B(n399), .Z(n395) );
  AND U620 ( .A(n400), .B(n401), .Z(n398) );
  XNOR U621 ( .A(x[220]), .B(n399), .Z(n401) );
  XOR U622 ( .A(n402), .B(n403), .Z(n399) );
  AND U623 ( .A(n404), .B(n405), .Z(n402) );
  XNOR U624 ( .A(x[219]), .B(n403), .Z(n405) );
  XOR U625 ( .A(n406), .B(n407), .Z(n403) );
  AND U626 ( .A(n408), .B(n409), .Z(n406) );
  XNOR U627 ( .A(x[218]), .B(n407), .Z(n409) );
  XOR U628 ( .A(n410), .B(n411), .Z(n407) );
  AND U629 ( .A(n412), .B(n413), .Z(n410) );
  XNOR U630 ( .A(x[217]), .B(n411), .Z(n413) );
  XOR U631 ( .A(n414), .B(n415), .Z(n411) );
  AND U632 ( .A(n416), .B(n417), .Z(n414) );
  XNOR U633 ( .A(x[216]), .B(n415), .Z(n417) );
  XOR U634 ( .A(n418), .B(n419), .Z(n415) );
  AND U635 ( .A(n420), .B(n421), .Z(n418) );
  XNOR U636 ( .A(x[215]), .B(n419), .Z(n421) );
  XOR U637 ( .A(n422), .B(n423), .Z(n419) );
  AND U638 ( .A(n424), .B(n425), .Z(n422) );
  XNOR U639 ( .A(x[214]), .B(n423), .Z(n425) );
  XOR U640 ( .A(n426), .B(n427), .Z(n423) );
  AND U641 ( .A(n428), .B(n429), .Z(n426) );
  XNOR U642 ( .A(x[213]), .B(n427), .Z(n429) );
  XOR U643 ( .A(n430), .B(n431), .Z(n427) );
  AND U644 ( .A(n432), .B(n433), .Z(n430) );
  XNOR U645 ( .A(x[212]), .B(n431), .Z(n433) );
  XOR U646 ( .A(n434), .B(n435), .Z(n431) );
  AND U647 ( .A(n436), .B(n437), .Z(n434) );
  XNOR U648 ( .A(x[211]), .B(n435), .Z(n437) );
  XOR U649 ( .A(n438), .B(n439), .Z(n435) );
  AND U650 ( .A(n440), .B(n441), .Z(n438) );
  XNOR U651 ( .A(x[210]), .B(n439), .Z(n441) );
  XOR U652 ( .A(n442), .B(n443), .Z(n439) );
  AND U653 ( .A(n444), .B(n445), .Z(n442) );
  XNOR U654 ( .A(x[209]), .B(n443), .Z(n445) );
  XOR U655 ( .A(n446), .B(n447), .Z(n443) );
  AND U656 ( .A(n448), .B(n449), .Z(n446) );
  XNOR U657 ( .A(x[208]), .B(n447), .Z(n449) );
  XOR U658 ( .A(n450), .B(n451), .Z(n447) );
  AND U659 ( .A(n452), .B(n453), .Z(n450) );
  XNOR U660 ( .A(x[207]), .B(n451), .Z(n453) );
  XOR U661 ( .A(n454), .B(n455), .Z(n451) );
  AND U662 ( .A(n456), .B(n457), .Z(n454) );
  XNOR U663 ( .A(x[206]), .B(n455), .Z(n457) );
  XOR U664 ( .A(n458), .B(n459), .Z(n455) );
  AND U665 ( .A(n460), .B(n461), .Z(n458) );
  XNOR U666 ( .A(x[205]), .B(n459), .Z(n461) );
  XOR U667 ( .A(n462), .B(n463), .Z(n459) );
  AND U668 ( .A(n464), .B(n465), .Z(n462) );
  XNOR U669 ( .A(x[204]), .B(n463), .Z(n465) );
  XOR U670 ( .A(n466), .B(n467), .Z(n463) );
  AND U671 ( .A(n468), .B(n469), .Z(n466) );
  XNOR U672 ( .A(x[203]), .B(n467), .Z(n469) );
  XOR U673 ( .A(n470), .B(n471), .Z(n467) );
  AND U674 ( .A(n472), .B(n473), .Z(n470) );
  XNOR U675 ( .A(x[202]), .B(n471), .Z(n473) );
  XOR U676 ( .A(n474), .B(n475), .Z(n471) );
  AND U677 ( .A(n476), .B(n477), .Z(n474) );
  XNOR U678 ( .A(x[201]), .B(n475), .Z(n477) );
  XOR U679 ( .A(n478), .B(n479), .Z(n475) );
  AND U680 ( .A(n480), .B(n481), .Z(n478) );
  XNOR U681 ( .A(x[200]), .B(n479), .Z(n481) );
  XOR U682 ( .A(n482), .B(n483), .Z(n479) );
  AND U683 ( .A(n484), .B(n485), .Z(n482) );
  XNOR U684 ( .A(x[199]), .B(n483), .Z(n485) );
  XOR U685 ( .A(n486), .B(n487), .Z(n483) );
  AND U686 ( .A(n488), .B(n489), .Z(n486) );
  XNOR U687 ( .A(x[198]), .B(n487), .Z(n489) );
  XOR U688 ( .A(n490), .B(n491), .Z(n487) );
  AND U689 ( .A(n492), .B(n493), .Z(n490) );
  XNOR U690 ( .A(x[197]), .B(n491), .Z(n493) );
  XOR U691 ( .A(n494), .B(n495), .Z(n491) );
  AND U692 ( .A(n496), .B(n497), .Z(n494) );
  XNOR U693 ( .A(x[196]), .B(n495), .Z(n497) );
  XOR U694 ( .A(n498), .B(n499), .Z(n495) );
  AND U695 ( .A(n500), .B(n501), .Z(n498) );
  XNOR U696 ( .A(x[195]), .B(n499), .Z(n501) );
  XOR U697 ( .A(n502), .B(n503), .Z(n499) );
  AND U698 ( .A(n504), .B(n505), .Z(n502) );
  XNOR U699 ( .A(x[194]), .B(n503), .Z(n505) );
  XOR U700 ( .A(n506), .B(n507), .Z(n503) );
  AND U701 ( .A(n508), .B(n509), .Z(n506) );
  XNOR U702 ( .A(x[193]), .B(n507), .Z(n509) );
  XOR U703 ( .A(n510), .B(n511), .Z(n507) );
  AND U704 ( .A(n512), .B(n513), .Z(n510) );
  XNOR U705 ( .A(x[192]), .B(n511), .Z(n513) );
  XOR U706 ( .A(n514), .B(n515), .Z(n511) );
  AND U707 ( .A(n516), .B(n517), .Z(n514) );
  XNOR U708 ( .A(x[191]), .B(n515), .Z(n517) );
  XOR U709 ( .A(n518), .B(n519), .Z(n515) );
  AND U710 ( .A(n520), .B(n521), .Z(n518) );
  XNOR U711 ( .A(x[190]), .B(n519), .Z(n521) );
  XOR U712 ( .A(n522), .B(n523), .Z(n519) );
  AND U713 ( .A(n524), .B(n525), .Z(n522) );
  XNOR U714 ( .A(x[189]), .B(n523), .Z(n525) );
  XOR U715 ( .A(n526), .B(n527), .Z(n523) );
  AND U716 ( .A(n528), .B(n529), .Z(n526) );
  XNOR U717 ( .A(x[188]), .B(n527), .Z(n529) );
  XOR U718 ( .A(n530), .B(n531), .Z(n527) );
  AND U719 ( .A(n532), .B(n533), .Z(n530) );
  XNOR U720 ( .A(x[187]), .B(n531), .Z(n533) );
  XOR U721 ( .A(n534), .B(n535), .Z(n531) );
  AND U722 ( .A(n536), .B(n537), .Z(n534) );
  XNOR U723 ( .A(x[186]), .B(n535), .Z(n537) );
  XOR U724 ( .A(n538), .B(n539), .Z(n535) );
  AND U725 ( .A(n540), .B(n541), .Z(n538) );
  XNOR U726 ( .A(x[185]), .B(n539), .Z(n541) );
  XOR U727 ( .A(n542), .B(n543), .Z(n539) );
  AND U728 ( .A(n544), .B(n545), .Z(n542) );
  XNOR U729 ( .A(x[184]), .B(n543), .Z(n545) );
  XOR U730 ( .A(n546), .B(n547), .Z(n543) );
  AND U731 ( .A(n548), .B(n549), .Z(n546) );
  XNOR U732 ( .A(x[183]), .B(n547), .Z(n549) );
  XOR U733 ( .A(n550), .B(n551), .Z(n547) );
  AND U734 ( .A(n552), .B(n553), .Z(n550) );
  XNOR U735 ( .A(x[182]), .B(n551), .Z(n553) );
  XOR U736 ( .A(n554), .B(n555), .Z(n551) );
  AND U737 ( .A(n556), .B(n557), .Z(n554) );
  XNOR U738 ( .A(x[181]), .B(n555), .Z(n557) );
  XOR U739 ( .A(n558), .B(n559), .Z(n555) );
  AND U740 ( .A(n560), .B(n561), .Z(n558) );
  XNOR U741 ( .A(x[180]), .B(n559), .Z(n561) );
  XOR U742 ( .A(n562), .B(n563), .Z(n559) );
  AND U743 ( .A(n564), .B(n565), .Z(n562) );
  XNOR U744 ( .A(x[179]), .B(n563), .Z(n565) );
  XOR U745 ( .A(n566), .B(n567), .Z(n563) );
  AND U746 ( .A(n568), .B(n569), .Z(n566) );
  XNOR U747 ( .A(x[178]), .B(n567), .Z(n569) );
  XOR U748 ( .A(n570), .B(n571), .Z(n567) );
  AND U749 ( .A(n572), .B(n573), .Z(n570) );
  XNOR U750 ( .A(x[177]), .B(n571), .Z(n573) );
  XOR U751 ( .A(n574), .B(n575), .Z(n571) );
  AND U752 ( .A(n576), .B(n577), .Z(n574) );
  XNOR U753 ( .A(x[176]), .B(n575), .Z(n577) );
  XOR U754 ( .A(n578), .B(n579), .Z(n575) );
  AND U755 ( .A(n580), .B(n581), .Z(n578) );
  XNOR U756 ( .A(x[175]), .B(n579), .Z(n581) );
  XOR U757 ( .A(n582), .B(n583), .Z(n579) );
  AND U758 ( .A(n584), .B(n585), .Z(n582) );
  XNOR U759 ( .A(x[174]), .B(n583), .Z(n585) );
  XOR U760 ( .A(n586), .B(n587), .Z(n583) );
  AND U761 ( .A(n588), .B(n589), .Z(n586) );
  XNOR U762 ( .A(x[173]), .B(n587), .Z(n589) );
  XOR U763 ( .A(n590), .B(n591), .Z(n587) );
  AND U764 ( .A(n592), .B(n593), .Z(n590) );
  XNOR U765 ( .A(x[172]), .B(n591), .Z(n593) );
  XOR U766 ( .A(n594), .B(n595), .Z(n591) );
  AND U767 ( .A(n596), .B(n597), .Z(n594) );
  XNOR U768 ( .A(x[171]), .B(n595), .Z(n597) );
  XOR U769 ( .A(n598), .B(n599), .Z(n595) );
  AND U770 ( .A(n600), .B(n601), .Z(n598) );
  XNOR U771 ( .A(x[170]), .B(n599), .Z(n601) );
  XOR U772 ( .A(n602), .B(n603), .Z(n599) );
  AND U773 ( .A(n604), .B(n605), .Z(n602) );
  XNOR U774 ( .A(x[169]), .B(n603), .Z(n605) );
  XOR U775 ( .A(n606), .B(n607), .Z(n603) );
  AND U776 ( .A(n608), .B(n609), .Z(n606) );
  XNOR U777 ( .A(x[168]), .B(n607), .Z(n609) );
  XOR U778 ( .A(n610), .B(n611), .Z(n607) );
  AND U779 ( .A(n612), .B(n613), .Z(n610) );
  XNOR U780 ( .A(x[167]), .B(n611), .Z(n613) );
  XOR U781 ( .A(n614), .B(n615), .Z(n611) );
  AND U782 ( .A(n616), .B(n617), .Z(n614) );
  XNOR U783 ( .A(x[166]), .B(n615), .Z(n617) );
  XOR U784 ( .A(n618), .B(n619), .Z(n615) );
  AND U785 ( .A(n620), .B(n621), .Z(n618) );
  XNOR U786 ( .A(x[165]), .B(n619), .Z(n621) );
  XOR U787 ( .A(n622), .B(n623), .Z(n619) );
  AND U788 ( .A(n624), .B(n625), .Z(n622) );
  XNOR U789 ( .A(x[164]), .B(n623), .Z(n625) );
  XOR U790 ( .A(n626), .B(n627), .Z(n623) );
  AND U791 ( .A(n628), .B(n629), .Z(n626) );
  XNOR U792 ( .A(x[163]), .B(n627), .Z(n629) );
  XOR U793 ( .A(n630), .B(n631), .Z(n627) );
  AND U794 ( .A(n632), .B(n633), .Z(n630) );
  XNOR U795 ( .A(x[162]), .B(n631), .Z(n633) );
  XOR U796 ( .A(n634), .B(n635), .Z(n631) );
  AND U797 ( .A(n636), .B(n637), .Z(n634) );
  XNOR U798 ( .A(x[161]), .B(n635), .Z(n637) );
  XOR U799 ( .A(n638), .B(n639), .Z(n635) );
  AND U800 ( .A(n640), .B(n641), .Z(n638) );
  XNOR U801 ( .A(x[160]), .B(n639), .Z(n641) );
  XOR U802 ( .A(n642), .B(n643), .Z(n639) );
  AND U803 ( .A(n644), .B(n645), .Z(n642) );
  XNOR U804 ( .A(x[159]), .B(n643), .Z(n645) );
  XOR U805 ( .A(n646), .B(n647), .Z(n643) );
  AND U806 ( .A(n648), .B(n649), .Z(n646) );
  XNOR U807 ( .A(x[158]), .B(n647), .Z(n649) );
  XOR U808 ( .A(n650), .B(n651), .Z(n647) );
  AND U809 ( .A(n652), .B(n653), .Z(n650) );
  XNOR U810 ( .A(x[157]), .B(n651), .Z(n653) );
  XOR U811 ( .A(n654), .B(n655), .Z(n651) );
  AND U812 ( .A(n656), .B(n657), .Z(n654) );
  XNOR U813 ( .A(x[156]), .B(n655), .Z(n657) );
  XOR U814 ( .A(n658), .B(n659), .Z(n655) );
  AND U815 ( .A(n660), .B(n661), .Z(n658) );
  XNOR U816 ( .A(x[155]), .B(n659), .Z(n661) );
  XOR U817 ( .A(n662), .B(n663), .Z(n659) );
  AND U818 ( .A(n664), .B(n665), .Z(n662) );
  XNOR U819 ( .A(x[154]), .B(n663), .Z(n665) );
  XOR U820 ( .A(n666), .B(n667), .Z(n663) );
  AND U821 ( .A(n668), .B(n669), .Z(n666) );
  XNOR U822 ( .A(x[153]), .B(n667), .Z(n669) );
  XOR U823 ( .A(n670), .B(n671), .Z(n667) );
  AND U824 ( .A(n672), .B(n673), .Z(n670) );
  XNOR U825 ( .A(x[152]), .B(n671), .Z(n673) );
  XOR U826 ( .A(n674), .B(n675), .Z(n671) );
  AND U827 ( .A(n676), .B(n677), .Z(n674) );
  XNOR U828 ( .A(x[151]), .B(n675), .Z(n677) );
  XOR U829 ( .A(n678), .B(n679), .Z(n675) );
  AND U830 ( .A(n680), .B(n681), .Z(n678) );
  XNOR U831 ( .A(x[150]), .B(n679), .Z(n681) );
  XOR U832 ( .A(n682), .B(n683), .Z(n679) );
  AND U833 ( .A(n684), .B(n685), .Z(n682) );
  XNOR U834 ( .A(x[149]), .B(n683), .Z(n685) );
  XOR U835 ( .A(n686), .B(n687), .Z(n683) );
  AND U836 ( .A(n688), .B(n689), .Z(n686) );
  XNOR U837 ( .A(x[148]), .B(n687), .Z(n689) );
  XOR U838 ( .A(n690), .B(n691), .Z(n687) );
  AND U839 ( .A(n692), .B(n693), .Z(n690) );
  XNOR U840 ( .A(x[147]), .B(n691), .Z(n693) );
  XOR U841 ( .A(n694), .B(n695), .Z(n691) );
  AND U842 ( .A(n696), .B(n697), .Z(n694) );
  XNOR U843 ( .A(x[146]), .B(n695), .Z(n697) );
  XOR U844 ( .A(n698), .B(n699), .Z(n695) );
  AND U845 ( .A(n700), .B(n701), .Z(n698) );
  XNOR U846 ( .A(x[145]), .B(n699), .Z(n701) );
  XOR U847 ( .A(n702), .B(n703), .Z(n699) );
  AND U848 ( .A(n704), .B(n705), .Z(n702) );
  XNOR U849 ( .A(x[144]), .B(n703), .Z(n705) );
  XOR U850 ( .A(n706), .B(n707), .Z(n703) );
  AND U851 ( .A(n708), .B(n709), .Z(n706) );
  XNOR U852 ( .A(x[143]), .B(n707), .Z(n709) );
  XOR U853 ( .A(n710), .B(n711), .Z(n707) );
  AND U854 ( .A(n712), .B(n713), .Z(n710) );
  XNOR U855 ( .A(x[142]), .B(n711), .Z(n713) );
  XOR U856 ( .A(n714), .B(n715), .Z(n711) );
  AND U857 ( .A(n716), .B(n717), .Z(n714) );
  XNOR U858 ( .A(x[141]), .B(n715), .Z(n717) );
  XOR U859 ( .A(n718), .B(n719), .Z(n715) );
  AND U860 ( .A(n720), .B(n721), .Z(n718) );
  XNOR U861 ( .A(x[140]), .B(n719), .Z(n721) );
  XOR U862 ( .A(n722), .B(n723), .Z(n719) );
  AND U863 ( .A(n724), .B(n725), .Z(n722) );
  XNOR U864 ( .A(x[139]), .B(n723), .Z(n725) );
  XOR U865 ( .A(n726), .B(n727), .Z(n723) );
  AND U866 ( .A(n728), .B(n729), .Z(n726) );
  XNOR U867 ( .A(x[138]), .B(n727), .Z(n729) );
  XOR U868 ( .A(n730), .B(n731), .Z(n727) );
  AND U869 ( .A(n732), .B(n733), .Z(n730) );
  XNOR U870 ( .A(x[137]), .B(n731), .Z(n733) );
  XOR U871 ( .A(n734), .B(n735), .Z(n731) );
  AND U872 ( .A(n736), .B(n737), .Z(n734) );
  XNOR U873 ( .A(x[136]), .B(n735), .Z(n737) );
  XOR U874 ( .A(n738), .B(n739), .Z(n735) );
  AND U875 ( .A(n740), .B(n741), .Z(n738) );
  XNOR U876 ( .A(x[135]), .B(n739), .Z(n741) );
  XOR U877 ( .A(n742), .B(n743), .Z(n739) );
  AND U878 ( .A(n744), .B(n745), .Z(n742) );
  XNOR U879 ( .A(x[134]), .B(n743), .Z(n745) );
  XOR U880 ( .A(n746), .B(n747), .Z(n743) );
  AND U881 ( .A(n748), .B(n749), .Z(n746) );
  XNOR U882 ( .A(x[133]), .B(n747), .Z(n749) );
  XOR U883 ( .A(n750), .B(n751), .Z(n747) );
  AND U884 ( .A(n752), .B(n753), .Z(n750) );
  XNOR U885 ( .A(x[132]), .B(n751), .Z(n753) );
  XOR U886 ( .A(n754), .B(n755), .Z(n751) );
  AND U887 ( .A(n756), .B(n757), .Z(n754) );
  XNOR U888 ( .A(x[131]), .B(n755), .Z(n757) );
  XOR U889 ( .A(n758), .B(n759), .Z(n755) );
  AND U890 ( .A(n760), .B(n761), .Z(n758) );
  XNOR U891 ( .A(x[130]), .B(n759), .Z(n761) );
  XOR U892 ( .A(n762), .B(n763), .Z(n759) );
  AND U893 ( .A(n764), .B(n765), .Z(n762) );
  XNOR U894 ( .A(x[129]), .B(n763), .Z(n765) );
  XOR U895 ( .A(n766), .B(n767), .Z(n763) );
  AND U896 ( .A(n768), .B(n769), .Z(n766) );
  XNOR U897 ( .A(x[128]), .B(n767), .Z(n769) );
  XOR U898 ( .A(n770), .B(n771), .Z(n767) );
  AND U899 ( .A(n772), .B(n773), .Z(n770) );
  XNOR U900 ( .A(x[127]), .B(n771), .Z(n773) );
  XOR U901 ( .A(n774), .B(n775), .Z(n771) );
  AND U902 ( .A(n776), .B(n777), .Z(n774) );
  XNOR U903 ( .A(x[126]), .B(n775), .Z(n777) );
  XOR U904 ( .A(n778), .B(n779), .Z(n775) );
  AND U905 ( .A(n780), .B(n781), .Z(n778) );
  XNOR U906 ( .A(x[125]), .B(n779), .Z(n781) );
  XOR U907 ( .A(n782), .B(n783), .Z(n779) );
  AND U908 ( .A(n784), .B(n785), .Z(n782) );
  XNOR U909 ( .A(x[124]), .B(n783), .Z(n785) );
  XOR U910 ( .A(n786), .B(n787), .Z(n783) );
  AND U911 ( .A(n788), .B(n789), .Z(n786) );
  XNOR U912 ( .A(x[123]), .B(n787), .Z(n789) );
  XOR U913 ( .A(n790), .B(n791), .Z(n787) );
  AND U914 ( .A(n792), .B(n793), .Z(n790) );
  XNOR U915 ( .A(x[122]), .B(n791), .Z(n793) );
  XOR U916 ( .A(n794), .B(n795), .Z(n791) );
  AND U917 ( .A(n796), .B(n797), .Z(n794) );
  XNOR U918 ( .A(x[121]), .B(n795), .Z(n797) );
  XOR U919 ( .A(n798), .B(n799), .Z(n795) );
  AND U920 ( .A(n800), .B(n801), .Z(n798) );
  XNOR U921 ( .A(x[120]), .B(n799), .Z(n801) );
  XOR U922 ( .A(n802), .B(n803), .Z(n799) );
  AND U923 ( .A(n804), .B(n805), .Z(n802) );
  XNOR U924 ( .A(x[119]), .B(n803), .Z(n805) );
  XOR U925 ( .A(n806), .B(n807), .Z(n803) );
  AND U926 ( .A(n808), .B(n809), .Z(n806) );
  XNOR U927 ( .A(x[118]), .B(n807), .Z(n809) );
  XOR U928 ( .A(n810), .B(n811), .Z(n807) );
  AND U929 ( .A(n812), .B(n813), .Z(n810) );
  XNOR U930 ( .A(x[117]), .B(n811), .Z(n813) );
  XOR U931 ( .A(n814), .B(n815), .Z(n811) );
  AND U932 ( .A(n816), .B(n817), .Z(n814) );
  XNOR U933 ( .A(x[116]), .B(n815), .Z(n817) );
  XOR U934 ( .A(n818), .B(n819), .Z(n815) );
  AND U935 ( .A(n820), .B(n821), .Z(n818) );
  XNOR U936 ( .A(x[115]), .B(n819), .Z(n821) );
  XOR U937 ( .A(n822), .B(n823), .Z(n819) );
  AND U938 ( .A(n824), .B(n825), .Z(n822) );
  XNOR U939 ( .A(x[114]), .B(n823), .Z(n825) );
  XOR U940 ( .A(n826), .B(n827), .Z(n823) );
  AND U941 ( .A(n828), .B(n829), .Z(n826) );
  XNOR U942 ( .A(x[113]), .B(n827), .Z(n829) );
  XOR U943 ( .A(n830), .B(n831), .Z(n827) );
  AND U944 ( .A(n832), .B(n833), .Z(n830) );
  XNOR U945 ( .A(x[112]), .B(n831), .Z(n833) );
  XOR U946 ( .A(n834), .B(n835), .Z(n831) );
  AND U947 ( .A(n836), .B(n837), .Z(n834) );
  XNOR U948 ( .A(x[111]), .B(n835), .Z(n837) );
  XOR U949 ( .A(n838), .B(n839), .Z(n835) );
  AND U950 ( .A(n840), .B(n841), .Z(n838) );
  XNOR U951 ( .A(x[110]), .B(n839), .Z(n841) );
  XOR U952 ( .A(n842), .B(n843), .Z(n839) );
  AND U953 ( .A(n844), .B(n845), .Z(n842) );
  XNOR U954 ( .A(x[109]), .B(n843), .Z(n845) );
  XOR U955 ( .A(n846), .B(n847), .Z(n843) );
  AND U956 ( .A(n848), .B(n849), .Z(n846) );
  XNOR U957 ( .A(x[108]), .B(n847), .Z(n849) );
  XOR U958 ( .A(n850), .B(n851), .Z(n847) );
  AND U959 ( .A(n852), .B(n853), .Z(n850) );
  XNOR U960 ( .A(x[107]), .B(n851), .Z(n853) );
  XOR U961 ( .A(n854), .B(n855), .Z(n851) );
  AND U962 ( .A(n856), .B(n857), .Z(n854) );
  XNOR U963 ( .A(x[106]), .B(n855), .Z(n857) );
  XOR U964 ( .A(n858), .B(n859), .Z(n855) );
  AND U965 ( .A(n860), .B(n861), .Z(n858) );
  XNOR U966 ( .A(x[105]), .B(n859), .Z(n861) );
  XOR U967 ( .A(n862), .B(n863), .Z(n859) );
  AND U968 ( .A(n864), .B(n865), .Z(n862) );
  XNOR U969 ( .A(x[104]), .B(n863), .Z(n865) );
  XOR U970 ( .A(n866), .B(n867), .Z(n863) );
  AND U971 ( .A(n868), .B(n869), .Z(n866) );
  XNOR U972 ( .A(x[103]), .B(n867), .Z(n869) );
  XOR U973 ( .A(n870), .B(n871), .Z(n867) );
  AND U974 ( .A(n872), .B(n873), .Z(n870) );
  XNOR U975 ( .A(x[102]), .B(n871), .Z(n873) );
  XOR U976 ( .A(n874), .B(n875), .Z(n871) );
  AND U977 ( .A(n876), .B(n877), .Z(n874) );
  XNOR U978 ( .A(x[101]), .B(n875), .Z(n877) );
  XOR U979 ( .A(n878), .B(n879), .Z(n875) );
  AND U980 ( .A(n880), .B(n881), .Z(n878) );
  XNOR U981 ( .A(x[100]), .B(n879), .Z(n881) );
  XOR U982 ( .A(n882), .B(n883), .Z(n879) );
  AND U983 ( .A(n884), .B(n885), .Z(n882) );
  XNOR U984 ( .A(x[99]), .B(n883), .Z(n885) );
  XOR U985 ( .A(n886), .B(n887), .Z(n883) );
  AND U986 ( .A(n888), .B(n889), .Z(n886) );
  XNOR U987 ( .A(x[98]), .B(n887), .Z(n889) );
  XOR U988 ( .A(n890), .B(n891), .Z(n887) );
  AND U989 ( .A(n892), .B(n893), .Z(n890) );
  XNOR U990 ( .A(x[97]), .B(n891), .Z(n893) );
  XOR U991 ( .A(n894), .B(n895), .Z(n891) );
  AND U992 ( .A(n896), .B(n897), .Z(n894) );
  XNOR U993 ( .A(x[96]), .B(n895), .Z(n897) );
  XOR U994 ( .A(n898), .B(n899), .Z(n895) );
  AND U995 ( .A(n900), .B(n901), .Z(n898) );
  XNOR U996 ( .A(x[95]), .B(n899), .Z(n901) );
  XOR U997 ( .A(n902), .B(n903), .Z(n899) );
  AND U998 ( .A(n904), .B(n905), .Z(n902) );
  XNOR U999 ( .A(x[94]), .B(n903), .Z(n905) );
  XOR U1000 ( .A(n906), .B(n907), .Z(n903) );
  AND U1001 ( .A(n908), .B(n909), .Z(n906) );
  XNOR U1002 ( .A(x[93]), .B(n907), .Z(n909) );
  XOR U1003 ( .A(n910), .B(n911), .Z(n907) );
  AND U1004 ( .A(n912), .B(n913), .Z(n910) );
  XNOR U1005 ( .A(x[92]), .B(n911), .Z(n913) );
  XOR U1006 ( .A(n914), .B(n915), .Z(n911) );
  AND U1007 ( .A(n916), .B(n917), .Z(n914) );
  XNOR U1008 ( .A(x[91]), .B(n915), .Z(n917) );
  XOR U1009 ( .A(n918), .B(n919), .Z(n915) );
  AND U1010 ( .A(n920), .B(n921), .Z(n918) );
  XNOR U1011 ( .A(x[90]), .B(n919), .Z(n921) );
  XOR U1012 ( .A(n922), .B(n923), .Z(n919) );
  AND U1013 ( .A(n924), .B(n925), .Z(n922) );
  XNOR U1014 ( .A(x[89]), .B(n923), .Z(n925) );
  XOR U1015 ( .A(n926), .B(n927), .Z(n923) );
  AND U1016 ( .A(n928), .B(n929), .Z(n926) );
  XNOR U1017 ( .A(x[88]), .B(n927), .Z(n929) );
  XOR U1018 ( .A(n930), .B(n931), .Z(n927) );
  AND U1019 ( .A(n932), .B(n933), .Z(n930) );
  XNOR U1020 ( .A(x[87]), .B(n931), .Z(n933) );
  XOR U1021 ( .A(n934), .B(n935), .Z(n931) );
  AND U1022 ( .A(n936), .B(n937), .Z(n934) );
  XNOR U1023 ( .A(x[86]), .B(n935), .Z(n937) );
  XOR U1024 ( .A(n938), .B(n939), .Z(n935) );
  AND U1025 ( .A(n940), .B(n941), .Z(n938) );
  XNOR U1026 ( .A(x[85]), .B(n939), .Z(n941) );
  XOR U1027 ( .A(n942), .B(n943), .Z(n939) );
  AND U1028 ( .A(n944), .B(n945), .Z(n942) );
  XNOR U1029 ( .A(x[84]), .B(n943), .Z(n945) );
  XOR U1030 ( .A(n946), .B(n947), .Z(n943) );
  AND U1031 ( .A(n948), .B(n949), .Z(n946) );
  XNOR U1032 ( .A(x[83]), .B(n947), .Z(n949) );
  XOR U1033 ( .A(n950), .B(n951), .Z(n947) );
  AND U1034 ( .A(n952), .B(n953), .Z(n950) );
  XNOR U1035 ( .A(x[82]), .B(n951), .Z(n953) );
  XOR U1036 ( .A(n954), .B(n955), .Z(n951) );
  AND U1037 ( .A(n956), .B(n957), .Z(n954) );
  XNOR U1038 ( .A(x[81]), .B(n955), .Z(n957) );
  XOR U1039 ( .A(n958), .B(n959), .Z(n955) );
  AND U1040 ( .A(n960), .B(n961), .Z(n958) );
  XNOR U1041 ( .A(x[80]), .B(n959), .Z(n961) );
  XOR U1042 ( .A(n962), .B(n963), .Z(n959) );
  AND U1043 ( .A(n964), .B(n965), .Z(n962) );
  XNOR U1044 ( .A(x[79]), .B(n963), .Z(n965) );
  XOR U1045 ( .A(n966), .B(n967), .Z(n963) );
  AND U1046 ( .A(n968), .B(n969), .Z(n966) );
  XNOR U1047 ( .A(x[78]), .B(n967), .Z(n969) );
  XOR U1048 ( .A(n970), .B(n971), .Z(n967) );
  AND U1049 ( .A(n972), .B(n973), .Z(n970) );
  XNOR U1050 ( .A(x[77]), .B(n971), .Z(n973) );
  XOR U1051 ( .A(n974), .B(n975), .Z(n971) );
  AND U1052 ( .A(n976), .B(n977), .Z(n974) );
  XNOR U1053 ( .A(x[76]), .B(n975), .Z(n977) );
  XOR U1054 ( .A(n978), .B(n979), .Z(n975) );
  AND U1055 ( .A(n980), .B(n981), .Z(n978) );
  XNOR U1056 ( .A(x[75]), .B(n979), .Z(n981) );
  XOR U1057 ( .A(n982), .B(n983), .Z(n979) );
  AND U1058 ( .A(n984), .B(n985), .Z(n982) );
  XNOR U1059 ( .A(x[74]), .B(n983), .Z(n985) );
  XOR U1060 ( .A(n986), .B(n987), .Z(n983) );
  AND U1061 ( .A(n988), .B(n989), .Z(n986) );
  XNOR U1062 ( .A(x[73]), .B(n987), .Z(n989) );
  XOR U1063 ( .A(n990), .B(n991), .Z(n987) );
  AND U1064 ( .A(n992), .B(n993), .Z(n990) );
  XNOR U1065 ( .A(x[72]), .B(n991), .Z(n993) );
  XOR U1066 ( .A(n994), .B(n995), .Z(n991) );
  AND U1067 ( .A(n996), .B(n997), .Z(n994) );
  XNOR U1068 ( .A(x[71]), .B(n995), .Z(n997) );
  XOR U1069 ( .A(n998), .B(n999), .Z(n995) );
  AND U1070 ( .A(n1000), .B(n1001), .Z(n998) );
  XNOR U1071 ( .A(x[70]), .B(n999), .Z(n1001) );
  XOR U1072 ( .A(n1002), .B(n1003), .Z(n999) );
  AND U1073 ( .A(n1004), .B(n1005), .Z(n1002) );
  XNOR U1074 ( .A(x[69]), .B(n1003), .Z(n1005) );
  XOR U1075 ( .A(n1006), .B(n1007), .Z(n1003) );
  AND U1076 ( .A(n1008), .B(n1009), .Z(n1006) );
  XNOR U1077 ( .A(x[68]), .B(n1007), .Z(n1009) );
  XOR U1078 ( .A(n1010), .B(n1011), .Z(n1007) );
  AND U1079 ( .A(n1012), .B(n1013), .Z(n1010) );
  XNOR U1080 ( .A(x[67]), .B(n1011), .Z(n1013) );
  XOR U1081 ( .A(n1014), .B(n1015), .Z(n1011) );
  AND U1082 ( .A(n1016), .B(n1017), .Z(n1014) );
  XNOR U1083 ( .A(x[66]), .B(n1015), .Z(n1017) );
  XOR U1084 ( .A(n1018), .B(n1019), .Z(n1015) );
  AND U1085 ( .A(n1020), .B(n1021), .Z(n1018) );
  XNOR U1086 ( .A(x[65]), .B(n1019), .Z(n1021) );
  XOR U1087 ( .A(n1022), .B(n1023), .Z(n1019) );
  AND U1088 ( .A(n1024), .B(n1025), .Z(n1022) );
  XNOR U1089 ( .A(x[64]), .B(n1023), .Z(n1025) );
  XOR U1090 ( .A(n1026), .B(n1027), .Z(n1023) );
  AND U1091 ( .A(n1028), .B(n1029), .Z(n1026) );
  XNOR U1092 ( .A(x[63]), .B(n1027), .Z(n1029) );
  XOR U1093 ( .A(n1030), .B(n1031), .Z(n1027) );
  AND U1094 ( .A(n1032), .B(n1033), .Z(n1030) );
  XNOR U1095 ( .A(x[62]), .B(n1031), .Z(n1033) );
  XOR U1096 ( .A(n1034), .B(n1035), .Z(n1031) );
  AND U1097 ( .A(n1036), .B(n1037), .Z(n1034) );
  XNOR U1098 ( .A(x[61]), .B(n1035), .Z(n1037) );
  XOR U1099 ( .A(n1038), .B(n1039), .Z(n1035) );
  AND U1100 ( .A(n1040), .B(n1041), .Z(n1038) );
  XNOR U1101 ( .A(x[60]), .B(n1039), .Z(n1041) );
  XOR U1102 ( .A(n1042), .B(n1043), .Z(n1039) );
  AND U1103 ( .A(n1044), .B(n1045), .Z(n1042) );
  XNOR U1104 ( .A(x[59]), .B(n1043), .Z(n1045) );
  XOR U1105 ( .A(n1046), .B(n1047), .Z(n1043) );
  AND U1106 ( .A(n1048), .B(n1049), .Z(n1046) );
  XNOR U1107 ( .A(x[58]), .B(n1047), .Z(n1049) );
  XOR U1108 ( .A(n1050), .B(n1051), .Z(n1047) );
  AND U1109 ( .A(n1052), .B(n1053), .Z(n1050) );
  XNOR U1110 ( .A(x[57]), .B(n1051), .Z(n1053) );
  XOR U1111 ( .A(n1054), .B(n1055), .Z(n1051) );
  AND U1112 ( .A(n1056), .B(n1057), .Z(n1054) );
  XNOR U1113 ( .A(x[56]), .B(n1055), .Z(n1057) );
  XOR U1114 ( .A(n1058), .B(n1059), .Z(n1055) );
  AND U1115 ( .A(n1060), .B(n1061), .Z(n1058) );
  XNOR U1116 ( .A(x[55]), .B(n1059), .Z(n1061) );
  XOR U1117 ( .A(n1062), .B(n1063), .Z(n1059) );
  AND U1118 ( .A(n1064), .B(n1065), .Z(n1062) );
  XNOR U1119 ( .A(x[54]), .B(n1063), .Z(n1065) );
  XOR U1120 ( .A(n1066), .B(n1067), .Z(n1063) );
  AND U1121 ( .A(n1068), .B(n1069), .Z(n1066) );
  XNOR U1122 ( .A(x[53]), .B(n1067), .Z(n1069) );
  XOR U1123 ( .A(n1070), .B(n1071), .Z(n1067) );
  AND U1124 ( .A(n1072), .B(n1073), .Z(n1070) );
  XNOR U1125 ( .A(x[52]), .B(n1071), .Z(n1073) );
  XOR U1126 ( .A(n1074), .B(n1075), .Z(n1071) );
  AND U1127 ( .A(n1076), .B(n1077), .Z(n1074) );
  XNOR U1128 ( .A(x[51]), .B(n1075), .Z(n1077) );
  XOR U1129 ( .A(n1078), .B(n1079), .Z(n1075) );
  AND U1130 ( .A(n1080), .B(n1081), .Z(n1078) );
  XNOR U1131 ( .A(x[50]), .B(n1079), .Z(n1081) );
  XOR U1132 ( .A(n1082), .B(n1083), .Z(n1079) );
  AND U1133 ( .A(n1084), .B(n1085), .Z(n1082) );
  XNOR U1134 ( .A(x[49]), .B(n1083), .Z(n1085) );
  XOR U1135 ( .A(n1086), .B(n1087), .Z(n1083) );
  AND U1136 ( .A(n1088), .B(n1089), .Z(n1086) );
  XNOR U1137 ( .A(x[48]), .B(n1087), .Z(n1089) );
  XOR U1138 ( .A(n1090), .B(n1091), .Z(n1087) );
  AND U1139 ( .A(n1092), .B(n1093), .Z(n1090) );
  XNOR U1140 ( .A(x[47]), .B(n1091), .Z(n1093) );
  XOR U1141 ( .A(n1094), .B(n1095), .Z(n1091) );
  AND U1142 ( .A(n1096), .B(n1097), .Z(n1094) );
  XNOR U1143 ( .A(x[46]), .B(n1095), .Z(n1097) );
  XOR U1144 ( .A(n1098), .B(n1099), .Z(n1095) );
  AND U1145 ( .A(n1100), .B(n1101), .Z(n1098) );
  XNOR U1146 ( .A(x[45]), .B(n1099), .Z(n1101) );
  XOR U1147 ( .A(n1102), .B(n1103), .Z(n1099) );
  AND U1148 ( .A(n1104), .B(n1105), .Z(n1102) );
  XNOR U1149 ( .A(x[44]), .B(n1103), .Z(n1105) );
  XOR U1150 ( .A(n1106), .B(n1107), .Z(n1103) );
  AND U1151 ( .A(n1108), .B(n1109), .Z(n1106) );
  XNOR U1152 ( .A(x[43]), .B(n1107), .Z(n1109) );
  XOR U1153 ( .A(n1110), .B(n1111), .Z(n1107) );
  AND U1154 ( .A(n1112), .B(n1113), .Z(n1110) );
  XNOR U1155 ( .A(x[42]), .B(n1111), .Z(n1113) );
  XOR U1156 ( .A(n1114), .B(n1115), .Z(n1111) );
  AND U1157 ( .A(n1116), .B(n1117), .Z(n1114) );
  XNOR U1158 ( .A(x[41]), .B(n1115), .Z(n1117) );
  XOR U1159 ( .A(n1118), .B(n1119), .Z(n1115) );
  AND U1160 ( .A(n1120), .B(n1121), .Z(n1118) );
  XNOR U1161 ( .A(x[40]), .B(n1119), .Z(n1121) );
  XOR U1162 ( .A(n1122), .B(n1123), .Z(n1119) );
  AND U1163 ( .A(n1124), .B(n1125), .Z(n1122) );
  XNOR U1164 ( .A(x[39]), .B(n1123), .Z(n1125) );
  XOR U1165 ( .A(n1126), .B(n1127), .Z(n1123) );
  AND U1166 ( .A(n1128), .B(n1129), .Z(n1126) );
  XNOR U1167 ( .A(x[38]), .B(n1127), .Z(n1129) );
  XOR U1168 ( .A(n1130), .B(n1131), .Z(n1127) );
  AND U1169 ( .A(n1132), .B(n1133), .Z(n1130) );
  XNOR U1170 ( .A(x[37]), .B(n1131), .Z(n1133) );
  XOR U1171 ( .A(n1134), .B(n1135), .Z(n1131) );
  AND U1172 ( .A(n1136), .B(n1137), .Z(n1134) );
  XNOR U1173 ( .A(x[36]), .B(n1135), .Z(n1137) );
  XOR U1174 ( .A(n1138), .B(n1139), .Z(n1135) );
  AND U1175 ( .A(n1140), .B(n1141), .Z(n1138) );
  XNOR U1176 ( .A(x[35]), .B(n1139), .Z(n1141) );
  XOR U1177 ( .A(n1142), .B(n1143), .Z(n1139) );
  AND U1178 ( .A(n1144), .B(n1145), .Z(n1142) );
  XNOR U1179 ( .A(x[34]), .B(n1143), .Z(n1145) );
  XOR U1180 ( .A(n1146), .B(n1147), .Z(n1143) );
  AND U1181 ( .A(n1148), .B(n1149), .Z(n1146) );
  XNOR U1182 ( .A(x[33]), .B(n1147), .Z(n1149) );
  XOR U1183 ( .A(n1150), .B(n1151), .Z(n1147) );
  AND U1184 ( .A(n1152), .B(n1153), .Z(n1150) );
  XNOR U1185 ( .A(x[32]), .B(n1151), .Z(n1153) );
  XOR U1186 ( .A(n1154), .B(n1155), .Z(n1151) );
  AND U1187 ( .A(n1156), .B(n1157), .Z(n1154) );
  XNOR U1188 ( .A(x[31]), .B(n1155), .Z(n1157) );
  XOR U1189 ( .A(n1158), .B(n1159), .Z(n1155) );
  AND U1190 ( .A(n1160), .B(n1161), .Z(n1158) );
  XNOR U1191 ( .A(x[30]), .B(n1159), .Z(n1161) );
  XOR U1192 ( .A(n1162), .B(n1163), .Z(n1159) );
  AND U1193 ( .A(n1164), .B(n1165), .Z(n1162) );
  XNOR U1194 ( .A(x[29]), .B(n1163), .Z(n1165) );
  XOR U1195 ( .A(n1166), .B(n1167), .Z(n1163) );
  AND U1196 ( .A(n1168), .B(n1169), .Z(n1166) );
  XNOR U1197 ( .A(x[28]), .B(n1167), .Z(n1169) );
  XOR U1198 ( .A(n1170), .B(n1171), .Z(n1167) );
  AND U1199 ( .A(n1172), .B(n1173), .Z(n1170) );
  XNOR U1200 ( .A(x[27]), .B(n1171), .Z(n1173) );
  XOR U1201 ( .A(n1174), .B(n1175), .Z(n1171) );
  AND U1202 ( .A(n1176), .B(n1177), .Z(n1174) );
  XNOR U1203 ( .A(x[26]), .B(n1175), .Z(n1177) );
  XOR U1204 ( .A(n1178), .B(n1179), .Z(n1175) );
  AND U1205 ( .A(n1180), .B(n1181), .Z(n1178) );
  XNOR U1206 ( .A(x[25]), .B(n1179), .Z(n1181) );
  XOR U1207 ( .A(n1182), .B(n1183), .Z(n1179) );
  AND U1208 ( .A(n1184), .B(n1185), .Z(n1182) );
  XNOR U1209 ( .A(x[24]), .B(n1183), .Z(n1185) );
  XOR U1210 ( .A(n1186), .B(n1187), .Z(n1183) );
  AND U1211 ( .A(n1188), .B(n1189), .Z(n1186) );
  XNOR U1212 ( .A(x[23]), .B(n1187), .Z(n1189) );
  XOR U1213 ( .A(n1190), .B(n1191), .Z(n1187) );
  AND U1214 ( .A(n1192), .B(n1193), .Z(n1190) );
  XNOR U1215 ( .A(x[22]), .B(n1191), .Z(n1193) );
  XOR U1216 ( .A(n1194), .B(n1195), .Z(n1191) );
  AND U1217 ( .A(n1196), .B(n1197), .Z(n1194) );
  XNOR U1218 ( .A(x[21]), .B(n1195), .Z(n1197) );
  XOR U1219 ( .A(n1198), .B(n1199), .Z(n1195) );
  AND U1220 ( .A(n1200), .B(n1201), .Z(n1198) );
  XNOR U1221 ( .A(x[20]), .B(n1199), .Z(n1201) );
  XOR U1222 ( .A(n1202), .B(n1203), .Z(n1199) );
  AND U1223 ( .A(n1204), .B(n1205), .Z(n1202) );
  XNOR U1224 ( .A(x[19]), .B(n1203), .Z(n1205) );
  XOR U1225 ( .A(n1206), .B(n1207), .Z(n1203) );
  AND U1226 ( .A(n1208), .B(n1209), .Z(n1206) );
  XNOR U1227 ( .A(x[18]), .B(n1207), .Z(n1209) );
  XOR U1228 ( .A(n1210), .B(n1211), .Z(n1207) );
  AND U1229 ( .A(n1212), .B(n1213), .Z(n1210) );
  XNOR U1230 ( .A(x[17]), .B(n1211), .Z(n1213) );
  XOR U1231 ( .A(n1214), .B(n1215), .Z(n1211) );
  AND U1232 ( .A(n1216), .B(n1217), .Z(n1214) );
  XNOR U1233 ( .A(x[16]), .B(n1215), .Z(n1217) );
  XOR U1234 ( .A(n1218), .B(n1219), .Z(n1215) );
  AND U1235 ( .A(n1220), .B(n1221), .Z(n1218) );
  XNOR U1236 ( .A(x[15]), .B(n1219), .Z(n1221) );
  XOR U1237 ( .A(n1222), .B(n1223), .Z(n1219) );
  AND U1238 ( .A(n1224), .B(n1225), .Z(n1222) );
  XNOR U1239 ( .A(x[14]), .B(n1223), .Z(n1225) );
  XOR U1240 ( .A(n1226), .B(n1227), .Z(n1223) );
  AND U1241 ( .A(n1228), .B(n1229), .Z(n1226) );
  XNOR U1242 ( .A(x[13]), .B(n1227), .Z(n1229) );
  XOR U1243 ( .A(n1230), .B(n1231), .Z(n1227) );
  AND U1244 ( .A(n1232), .B(n1233), .Z(n1230) );
  XNOR U1245 ( .A(x[12]), .B(n1231), .Z(n1233) );
  XOR U1246 ( .A(n1234), .B(n1235), .Z(n1231) );
  AND U1247 ( .A(n1236), .B(n1237), .Z(n1234) );
  XNOR U1248 ( .A(x[11]), .B(n1235), .Z(n1237) );
  XOR U1249 ( .A(n1238), .B(n1239), .Z(n1235) );
  AND U1250 ( .A(n1240), .B(n1241), .Z(n1238) );
  XNOR U1251 ( .A(x[10]), .B(n1239), .Z(n1241) );
  XOR U1252 ( .A(n1242), .B(n1243), .Z(n1239) );
  AND U1253 ( .A(n1244), .B(n1245), .Z(n1242) );
  XNOR U1254 ( .A(x[9]), .B(n1243), .Z(n1245) );
  XOR U1255 ( .A(n1246), .B(n1247), .Z(n1243) );
  AND U1256 ( .A(n1248), .B(n1249), .Z(n1246) );
  XNOR U1257 ( .A(x[8]), .B(n1247), .Z(n1249) );
  XOR U1258 ( .A(n1250), .B(n1251), .Z(n1247) );
  AND U1259 ( .A(n1252), .B(n1253), .Z(n1250) );
  XNOR U1260 ( .A(x[7]), .B(n1251), .Z(n1253) );
  XOR U1261 ( .A(n1254), .B(n1255), .Z(n1251) );
  AND U1262 ( .A(n1256), .B(n1257), .Z(n1254) );
  XNOR U1263 ( .A(x[6]), .B(n1255), .Z(n1257) );
  XOR U1264 ( .A(n1258), .B(n1259), .Z(n1255) );
  AND U1265 ( .A(n1260), .B(n1261), .Z(n1258) );
  XNOR U1266 ( .A(x[5]), .B(n1259), .Z(n1261) );
  XOR U1267 ( .A(n1262), .B(n1263), .Z(n1259) );
  AND U1268 ( .A(n1264), .B(n1265), .Z(n1262) );
  XNOR U1269 ( .A(x[4]), .B(n1263), .Z(n1265) );
  XOR U1270 ( .A(n1266), .B(n1267), .Z(n1263) );
  AND U1271 ( .A(n1268), .B(n1269), .Z(n1266) );
  XNOR U1272 ( .A(x[3]), .B(n1267), .Z(n1269) );
  XOR U1273 ( .A(n1270), .B(n1271), .Z(n1267) );
  AND U1274 ( .A(n1272), .B(n1273), .Z(n1270) );
  XNOR U1275 ( .A(x[2]), .B(n1271), .Z(n1273) );
  XOR U1276 ( .A(n1274), .B(n1275), .Z(n1271) );
  AND U1277 ( .A(n1276), .B(n1277), .Z(n1274) );
  XNOR U1278 ( .A(x[1]), .B(n1275), .Z(n1277) );
  XOR U1279 ( .A(y[1]), .B(n1275), .Z(n1276) );
  XOR U1280 ( .A(ci), .B(n1278), .Z(n1275) );
  NANDN U1281 ( .A(n1279), .B(n1280), .Z(n1278) );
  XOR U1282 ( .A(x[0]), .B(ci), .Z(n1280) );
  XOR U1283 ( .A(y[0]), .B(ci), .Z(n1279) );
endmodule

